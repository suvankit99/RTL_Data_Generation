
module dec(\count[0] , \count[1] , \count[2] , \count[3] , \count[4] ,
     \count[5] , \count[6] , \count[7] , \selectp1[0] , \selectp1[1] ,
     \selectp1[2] , \selectp1[3] , \selectp1[4] , \selectp1[5] ,
     \selectp1[6] , \selectp1[7] , \selectp1[8] , \selectp1[9] ,
     \selectp1[10] , \selectp1[11] , \selectp1[12] , \selectp1[13] ,
     \selectp1[14] , \selectp1[15] , \selectp1[16] , \selectp1[17] ,
     \selectp1[18] , \selectp1[19] , \selectp1[20] , \selectp1[21] ,
     \selectp1[22] , \selectp1[23] , \selectp1[24] , \selectp1[25] ,
     \selectp1[26] , \selectp1[27] , \selectp1[28] , \selectp1[29] ,
     \selectp1[30] , \selectp1[31] , \selectp1[32] , \selectp1[33] ,
     \selectp1[34] , \selectp1[35] , \selectp1[36] , \selectp1[37] ,
     \selectp1[38] , \selectp1[39] , \selectp1[40] , \selectp1[41] ,
     \selectp1[42] , \selectp1[43] , \selectp1[44] , \selectp1[45] ,
     \selectp1[46] , \selectp1[47] , \selectp1[48] , \selectp1[49] ,
     \selectp1[50] , \selectp1[51] , \selectp1[52] , \selectp1[53] ,
     \selectp1[54] , \selectp1[55] , \selectp1[56] , \selectp1[57] ,
     \selectp1[58] , \selectp1[59] , \selectp1[60] , \selectp1[61] ,
     \selectp1[62] , \selectp1[63] , \selectp1[64] , \selectp1[65] ,
     \selectp1[66] , \selectp1[67] , \selectp1[68] , \selectp1[69] ,
     \selectp1[70] , \selectp1[71] , \selectp1[72] , \selectp1[73] ,
     \selectp1[74] , \selectp1[75] , \selectp1[76] , \selectp1[77] ,
     \selectp1[78] , \selectp1[79] , \selectp1[80] , \selectp1[81] ,
     \selectp1[82] , \selectp1[83] , \selectp1[84] , \selectp1[85] ,
     \selectp1[86] , \selectp1[87] , \selectp1[88] , \selectp1[89] ,
     \selectp1[90] , \selectp1[91] , \selectp1[92] , \selectp1[93] ,
     \selectp1[94] , \selectp1[95] , \selectp1[96] , \selectp1[97] ,
     \selectp1[98] , \selectp1[99] , \selectp1[100] , \selectp1[101] ,
     \selectp1[102] , \selectp1[103] , \selectp1[104] , \selectp1[105]
     , \selectp1[106] , \selectp1[107] , \selectp1[108] ,
     \selectp1[109] , \selectp1[110] , \selectp1[111] , \selectp1[112]
     , \selectp1[113] , \selectp1[114] , \selectp1[115] ,
     \selectp1[116] , \selectp1[117] , \selectp1[118] , \selectp1[119]
     , \selectp1[120] , \selectp1[121] , \selectp1[122] ,
     \selectp1[123] , \selectp1[124] , \selectp1[125] , \selectp1[126]
     , \selectp1[127] , \selectp2[0] , \selectp2[1] , \selectp2[2] ,
     \selectp2[3] , \selectp2[4] , \selectp2[5] , \selectp2[6] ,
     \selectp2[7] , \selectp2[8] , \selectp2[9] , \selectp2[10] ,
     \selectp2[11] , \selectp2[12] , \selectp2[13] , \selectp2[14] ,
     \selectp2[15] , \selectp2[16] , \selectp2[17] , \selectp2[18] ,
     \selectp2[19] , \selectp2[20] , \selectp2[21] , \selectp2[22] ,
     \selectp2[23] , \selectp2[24] , \selectp2[25] , \selectp2[26] ,
     \selectp2[27] , \selectp2[28] , \selectp2[29] , \selectp2[30] ,
     \selectp2[31] , \selectp2[32] , \selectp2[33] , \selectp2[34] ,
     \selectp2[35] , \selectp2[36] , \selectp2[37] , \selectp2[38] ,
     \selectp2[39] , \selectp2[40] , \selectp2[41] , \selectp2[42] ,
     \selectp2[43] , \selectp2[44] , \selectp2[45] , \selectp2[46] ,
     \selectp2[47] , \selectp2[48] , \selectp2[49] , \selectp2[50] ,
     \selectp2[51] , \selectp2[52] , \selectp2[53] , \selectp2[54] ,
     \selectp2[55] , \selectp2[56] , \selectp2[57] , \selectp2[58] ,
     \selectp2[59] , \selectp2[60] , \selectp2[61] , \selectp2[62] ,
     \selectp2[63] , \selectp2[64] , \selectp2[65] , \selectp2[66] ,
     \selectp2[67] , \selectp2[68] , \selectp2[69] , \selectp2[70] ,
     \selectp2[71] , \selectp2[72] , \selectp2[73] , \selectp2[74] ,
     \selectp2[75] , \selectp2[76] , \selectp2[77] , \selectp2[78] ,
     \selectp2[79] , \selectp2[80] , \selectp2[81] , \selectp2[82] ,
     \selectp2[83] , \selectp2[84] , \selectp2[85] , \selectp2[86] ,
     \selectp2[87] , \selectp2[88] , \selectp2[89] , \selectp2[90] ,
     \selectp2[91] , \selectp2[92] , \selectp2[93] , \selectp2[94] ,
     \selectp2[95] , \selectp2[96] , \selectp2[97] , \selectp2[98] ,
     \selectp2[99] , \selectp2[100] , \selectp2[101] , \selectp2[102] ,
     \selectp2[103] , \selectp2[104] , \selectp2[105] , \selectp2[106]
     , \selectp2[107] , \selectp2[108] , \selectp2[109] ,
     \selectp2[110] , \selectp2[111] , \selectp2[112] , \selectp2[113]
     , \selectp2[114] , \selectp2[115] , \selectp2[116] ,
     \selectp2[117] , \selectp2[118] , \selectp2[119] , \selectp2[120]
     , \selectp2[121] , \selectp2[122] , \selectp2[123] ,
     \selectp2[124] , \selectp2[125] , \selectp2[126] , \selectp2[127]
     );
//   input \count[0] , \count[1] , \count[2] , \count[3] , \count[4] ,
       \count[5] , \count[6] , \count[7] ;
//   output \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
       \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
       \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
       \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
       \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
       \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
       \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
       \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
       \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
       \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
       \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
       \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
       \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
       \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
       \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
       \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
       \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
       \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
       \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
       \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
       \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
       \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
       \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
       \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
       \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
       \selectp1[100] , \selectp1[101] , \selectp1[102] ,
       \selectp1[103] , \selectp1[104] , \selectp1[105] ,
       \selectp1[106] , \selectp1[107] , \selectp1[108] ,
       \selectp1[109] , \selectp1[110] , \selectp1[111] ,
       \selectp1[112] , \selectp1[113] , \selectp1[114] ,
       \selectp1[115] , \selectp1[116] , \selectp1[117] ,
       \selectp1[118] , \selectp1[119] , \selectp1[120] ,
       \selectp1[121] , \selectp1[122] , \selectp1[123] ,
       \selectp1[124] , \selectp1[125] , \selectp1[126] ,
       \selectp1[127] , \selectp2[0] , \selectp2[1] , \selectp2[2] ,
       \selectp2[3] , \selectp2[4] , \selectp2[5] , \selectp2[6] ,
       \selectp2[7] , \selectp2[8] , \selectp2[9] , \selectp2[10] ,
       \selectp2[11] , \selectp2[12] , \selectp2[13] , \selectp2[14] ,
       \selectp2[15] , \selectp2[16] , \selectp2[17] , \selectp2[18] ,
       \selectp2[19] , \selectp2[20] , \selectp2[21] , \selectp2[22] ,
       \selectp2[23] , \selectp2[24] , \selectp2[25] , \selectp2[26] ,
       \selectp2[27] , \selectp2[28] , \selectp2[29] , \selectp2[30] ,
       \selectp2[31] , \selectp2[32] , \selectp2[33] , \selectp2[34] ,
       \selectp2[35] , \selectp2[36] , \selectp2[37] , \selectp2[38] ,
       \selectp2[39] , \selectp2[40] , \selectp2[41] , \selectp2[42] ,
       \selectp2[43] , \selectp2[44] , \selectp2[45] , \selectp2[46] ,
       \selectp2[47] , \selectp2[48] , \selectp2[49] , \selectp2[50] ,
       \selectp2[51] , \selectp2[52] , \selectp2[53] , \selectp2[54] ,
       \selectp2[55] , \selectp2[56] , \selectp2[57] , \selectp2[58] ,
       \selectp2[59] , \selectp2[60] , \selectp2[61] , \selectp2[62] ,
       \selectp2[63] , \selectp2[64] , \selectp2[65] , \selectp2[66] ,
       \selectp2[67] , \selectp2[68] , \selectp2[69] , \selectp2[70] ,
       \selectp2[71] , \selectp2[72] , \selectp2[73] , \selectp2[74] ,
       \selectp2[75] , \selectp2[76] , \selectp2[77] , \selectp2[78] ,
       \selectp2[79] , \selectp2[80] , \selectp2[81] , \selectp2[82] ,
       \selectp2[83] , \selectp2[84] , \selectp2[85] , \selectp2[86] ,
       \selectp2[87] , \selectp2[88] , \selectp2[89] , \selectp2[90] ,
       \selectp2[91] , \selectp2[92] , \selectp2[93] , \selectp2[94] ,
       \selectp2[95] , \selectp2[96] , \selectp2[97] , \selectp2[98] ,
       \selectp2[99] , \selectp2[100] , \selectp2[101] , \selectp2[102]
       , \selectp2[103] , \selectp2[104] , \selectp2[105] ,
       \selectp2[106] , \selectp2[107] , \selectp2[108] ,
       \selectp2[109] , \selectp2[110] , \selectp2[111] ,
       \selectp2[112] , \selectp2[113] , \selectp2[114] ,
       \selectp2[115] , \selectp2[116] , \selectp2[117] ,
       \selectp2[118] , \selectp2[119] , \selectp2[120] ,
       \selectp2[121] , \selectp2[122] , \selectp2[123] ,
       \selectp2[124] , \selectp2[125] , \selectp2[126] ,
       \selectp2[127] ;
  wire \count[0] , \count[1] , \count[2] , \count[3] , \count[4] ,
       \count[5] , \count[6] , \count[7] ;
  wire \selectp1[0] , \selectp1[1] , \selectp1[2] , \selectp1[3] ,
       \selectp1[4] , \selectp1[5] , \selectp1[6] , \selectp1[7] ,
       \selectp1[8] , \selectp1[9] , \selectp1[10] , \selectp1[11] ,
       \selectp1[12] , \selectp1[13] , \selectp1[14] , \selectp1[15] ,
       \selectp1[16] , \selectp1[17] , \selectp1[18] , \selectp1[19] ,
       \selectp1[20] , \selectp1[21] , \selectp1[22] , \selectp1[23] ,
       \selectp1[24] , \selectp1[25] , \selectp1[26] , \selectp1[27] ,
       \selectp1[28] , \selectp1[29] , \selectp1[30] , \selectp1[31] ,
       \selectp1[32] , \selectp1[33] , \selectp1[34] , \selectp1[35] ,
       \selectp1[36] , \selectp1[37] , \selectp1[38] , \selectp1[39] ,
       \selectp1[40] , \selectp1[41] , \selectp1[42] , \selectp1[43] ,
       \selectp1[44] , \selectp1[45] , \selectp1[46] , \selectp1[47] ,
       \selectp1[48] , \selectp1[49] , \selectp1[50] , \selectp1[51] ,
       \selectp1[52] , \selectp1[53] , \selectp1[54] , \selectp1[55] ,
       \selectp1[56] , \selectp1[57] , \selectp1[58] , \selectp1[59] ,
       \selectp1[60] , \selectp1[61] , \selectp1[62] , \selectp1[63] ,
       \selectp1[64] , \selectp1[65] , \selectp1[66] , \selectp1[67] ,
       \selectp1[68] , \selectp1[69] , \selectp1[70] , \selectp1[71] ,
       \selectp1[72] , \selectp1[73] , \selectp1[74] , \selectp1[75] ,
       \selectp1[76] , \selectp1[77] , \selectp1[78] , \selectp1[79] ,
       \selectp1[80] , \selectp1[81] , \selectp1[82] , \selectp1[83] ,
       \selectp1[84] , \selectp1[85] , \selectp1[86] , \selectp1[87] ,
       \selectp1[88] , \selectp1[89] , \selectp1[90] , \selectp1[91] ,
       \selectp1[92] , \selectp1[93] , \selectp1[94] , \selectp1[95] ,
       \selectp1[96] , \selectp1[97] , \selectp1[98] , \selectp1[99] ,
       \selectp1[100] , \selectp1[101] , \selectp1[102] ,
       \selectp1[103] , \selectp1[104] , \selectp1[105] ,
       \selectp1[106] , \selectp1[107] , \selectp1[108] ,
       \selectp1[109] , \selectp1[110] , \selectp1[111] ,
       \selectp1[112] , \selectp1[113] , \selectp1[114] ,
       \selectp1[115] , \selectp1[116] , \selectp1[117] ,
       \selectp1[118] , \selectp1[119] , \selectp1[120] ,
       \selectp1[121] , \selectp1[122] , \selectp1[123] ,
       \selectp1[124] , \selectp1[125] , \selectp1[126] ,
       \selectp1[127] , \selectp2[0] , \selectp2[1] , \selectp2[2] ,
       \selectp2[3] , \selectp2[4] , \selectp2[5] , \selectp2[6] ,
       \selectp2[7] , \selectp2[8] , \selectp2[9] , \selectp2[10] ,
       \selectp2[11] , \selectp2[12] , \selectp2[13] , \selectp2[14] ,
       \selectp2[15] , \selectp2[16] , \selectp2[17] , \selectp2[18] ,
       \selectp2[19] , \selectp2[20] , \selectp2[21] , \selectp2[22] ,
       \selectp2[23] , \selectp2[24] , \selectp2[25] , \selectp2[26] ,
       \selectp2[27] , \selectp2[28] , \selectp2[29] , \selectp2[30] ,
       \selectp2[31] , \selectp2[32] , \selectp2[33] , \selectp2[34] ,
       \selectp2[35] , \selectp2[36] , \selectp2[37] , \selectp2[38] ,
       \selectp2[39] , \selectp2[40] , \selectp2[41] , \selectp2[42] ,
       \selectp2[43] , \selectp2[44] , \selectp2[45] , \selectp2[46] ,
       \selectp2[47] , \selectp2[48] , \selectp2[49] , \selectp2[50] ,
       \selectp2[51] , \selectp2[52] , \selectp2[53] , \selectp2[54] ,
       \selectp2[55] , \selectp2[56] , \selectp2[57] , \selectp2[58] ,
       \selectp2[59] , \selectp2[60] , \selectp2[61] , \selectp2[62] ,
       \selectp2[63] , \selectp2[64] , \selectp2[65] , \selectp2[66] ,
       \selectp2[67] , \selectp2[68] , \selectp2[69] , \selectp2[70] ,
       \selectp2[71] , \selectp2[72] , \selectp2[73] , \selectp2[74] ,
       \selectp2[75] , \selectp2[76] , \selectp2[77] , \selectp2[78] ,
       \selectp2[79] , \selectp2[80] , \selectp2[81] , \selectp2[82] ,
       \selectp2[83] , \selectp2[84] , \selectp2[85] , \selectp2[86] ,
       \selectp2[87] , \selectp2[88] , \selectp2[89] , \selectp2[90] ,
       \selectp2[91] , \selectp2[92] , \selectp2[93] , \selectp2[94] ,
       \selectp2[95] , \selectp2[96] , \selectp2[97] , \selectp2[98] ,
       \selectp2[99] , \selectp2[100] , \selectp2[101] , \selectp2[102]
       , \selectp2[103] , \selectp2[104] , \selectp2[105] ,
       \selectp2[106] , \selectp2[107] , \selectp2[108] ,
       \selectp2[109] , \selectp2[110] , \selectp2[111] ,
       \selectp2[112] , \selectp2[113] , \selectp2[114] ,
       \selectp2[115] , \selectp2[116] , \selectp2[117] ,
       \selectp2[118] , \selectp2[119] , \selectp2[120] ,
       \selectp2[121] , \selectp2[122] , \selectp2[123] ,
       \selectp2[124] , \selectp2[125] , \selectp2[126] ,
       \selectp2[127] ;
  wire n265, n266, n267, n268, n269, n270, n272, n273;
  wire n275, n276, n278, n280, n281, n283, n284, n286;
  wire n288, n290, n291, n293, n295, n296, n298, n300;
  wire n302, n304, n306, n308, n309, n326, n327, n344;
  wire n345, n362, n363, n380, n397, n414, n431, n432;
  wire n449, n466, n483, n500, n501, n518, n535, n552;
  wire n_3, n_4, n_6, n_10, n_11, n_14, n_15, n_16;
  not g1 (n_3, \count[4] );
  not g2 (n_4, \count[5] );
  and g3 (n265, n_3, n_4);
  not g4 (n_6, \count[6] );
  and g5 (n266, n_6, \count[7] );
  and g6 (n267, n265, n266);
  not g7 (n_10, \count[0] );
  not g8 (n_11, \count[2] );
  and g9 (n268, n_10, n_11);
  not g10 (n_14, \count[1] );
  not g11 (n_15, \count[3] );
  and g12 (n269, n_14, n_15);
  and g13 (n270, n268, n269);
  and g14 (\selectp1[0] , n267, n270);
  and g15 (n272, \count[0] , n_11);
  and g16 (n273, n269, n272);
  and g17 (\selectp1[1] , n267, n273);
  and g18 (n275, \count[1] , n_15);
  and g19 (n276, n268, n275);
  and g20 (\selectp1[2] , n267, n276);
  and g21 (n278, n272, n275);
  and g22 (\selectp1[3] , n267, n278);
  and g23 (n280, n_10, \count[2] );
  and g24 (n281, n269, n280);
  and g25 (\selectp1[4] , n267, n281);
  and g26 (n283, \count[0] , \count[2] );
  and g27 (n284, n269, n283);
  and g28 (\selectp1[5] , n267, n284);
  and g29 (n286, n275, n280);
  and g30 (\selectp1[6] , n267, n286);
  and g31 (n288, n275, n283);
  and g32 (\selectp1[7] , n267, n288);
  and g33 (n290, n_14, \count[3] );
  and g34 (n291, n268, n290);
  and g35 (\selectp1[8] , n267, n291);
  and g36 (n293, n272, n290);
  and g37 (\selectp1[9] , n267, n293);
  and g38 (n295, \count[1] , \count[3] );
  and g39 (n296, n268, n295);
  and g40 (\selectp1[10] , n267, n296);
  and g41 (n298, n272, n295);
  and g42 (\selectp1[11] , n267, n298);
  and g43 (n300, n280, n290);
  and g44 (\selectp1[12] , n267, n300);
  and g45 (n302, n283, n290);
  and g46 (\selectp1[13] , n267, n302);
  and g47 (n304, n280, n295);
  and g48 (\selectp1[14] , n267, n304);
  and g49 (n306, n283, n295);
  and g50 (\selectp1[15] , n267, n306);
  and g51 (n308, \count[4] , n_4);
  and g52 (n309, n266, n308);
  and g53 (\selectp1[16] , n270, n309);
  and g54 (\selectp1[17] , n273, n309);
  and g55 (\selectp1[18] , n276, n309);
  and g56 (\selectp1[19] , n278, n309);
  and g57 (\selectp1[20] , n281, n309);
  and g58 (\selectp1[21] , n284, n309);
  and g59 (\selectp1[22] , n286, n309);
  and g60 (\selectp1[23] , n288, n309);
  and g61 (\selectp1[24] , n291, n309);
  and g62 (\selectp1[25] , n293, n309);
  and g63 (\selectp1[26] , n296, n309);
  and g64 (\selectp1[27] , n298, n309);
  and g65 (\selectp1[28] , n300, n309);
  and g66 (\selectp1[29] , n302, n309);
  and g67 (\selectp1[30] , n304, n309);
  and g68 (\selectp1[31] , n306, n309);
  and g69 (n326, n_3, \count[5] );
  and g70 (n327, n266, n326);
  and g71 (\selectp1[32] , n270, n327);
  and g72 (\selectp1[33] , n273, n327);
  and g73 (\selectp1[34] , n276, n327);
  and g74 (\selectp1[35] , n278, n327);
  and g75 (\selectp1[36] , n281, n327);
  and g76 (\selectp1[37] , n284, n327);
  and g77 (\selectp1[38] , n286, n327);
  and g78 (\selectp1[39] , n288, n327);
  and g79 (\selectp1[40] , n291, n327);
  and g80 (\selectp1[41] , n293, n327);
  and g81 (\selectp1[42] , n296, n327);
  and g82 (\selectp1[43] , n298, n327);
  and g83 (\selectp1[44] , n300, n327);
  and g84 (\selectp1[45] , n302, n327);
  and g85 (\selectp1[46] , n304, n327);
  and g86 (\selectp1[47] , n306, n327);
  and g87 (n344, \count[4] , \count[5] );
  and g88 (n345, n266, n344);
  and g89 (\selectp1[48] , n270, n345);
  and g90 (\selectp1[49] , n273, n345);
  and g91 (\selectp1[50] , n276, n345);
  and g92 (\selectp1[51] , n278, n345);
  and g93 (\selectp1[52] , n281, n345);
  and g94 (\selectp1[53] , n284, n345);
  and g95 (\selectp1[54] , n286, n345);
  and g96 (\selectp1[55] , n288, n345);
  and g97 (\selectp1[56] , n291, n345);
  and g98 (\selectp1[57] , n293, n345);
  and g99 (\selectp1[58] , n296, n345);
  and g100 (\selectp1[59] , n298, n345);
  and g101 (\selectp1[60] , n300, n345);
  and g102 (\selectp1[61] , n302, n345);
  and g103 (\selectp1[62] , n304, n345);
  and g104 (\selectp1[63] , n306, n345);
  and g105 (n362, \count[6] , \count[7] );
  and g106 (n363, n265, n362);
  and g107 (\selectp1[64] , n270, n363);
  and g108 (\selectp1[65] , n273, n363);
  and g109 (\selectp1[66] , n276, n363);
  and g110 (\selectp1[67] , n278, n363);
  and g111 (\selectp1[68] , n281, n363);
  and g112 (\selectp1[69] , n284, n363);
  and g113 (\selectp1[70] , n286, n363);
  and g114 (\selectp1[71] , n288, n363);
  and g115 (\selectp1[72] , n291, n363);
  and g116 (\selectp1[73] , n293, n363);
  and g117 (\selectp1[74] , n296, n363);
  and g118 (\selectp1[75] , n298, n363);
  and g119 (\selectp1[76] , n300, n363);
  and g120 (\selectp1[77] , n302, n363);
  and g121 (\selectp1[78] , n304, n363);
  and g122 (\selectp1[79] , n306, n363);
  and g123 (n380, n308, n362);
  and g124 (\selectp1[80] , n270, n380);
  and g125 (\selectp1[81] , n273, n380);
  and g126 (\selectp1[82] , n276, n380);
  and g127 (\selectp1[83] , n278, n380);
  and g128 (\selectp1[84] , n281, n380);
  and g129 (\selectp1[85] , n284, n380);
  and g130 (\selectp1[86] , n286, n380);
  and g131 (\selectp1[87] , n288, n380);
  and g132 (\selectp1[88] , n291, n380);
  and g133 (\selectp1[89] , n293, n380);
  and g134 (\selectp1[90] , n296, n380);
  and g135 (\selectp1[91] , n298, n380);
  and g136 (\selectp1[92] , n300, n380);
  and g137 (\selectp1[93] , n302, n380);
  and g138 (\selectp1[94] , n304, n380);
  and g139 (\selectp1[95] , n306, n380);
  and g140 (n397, n326, n362);
  and g141 (\selectp1[96] , n270, n397);
  and g142 (\selectp1[97] , n273, n397);
  and g143 (\selectp1[98] , n276, n397);
  and g144 (\selectp1[99] , n278, n397);
  and g145 (\selectp1[100] , n281, n397);
  and g146 (\selectp1[101] , n284, n397);
  and g147 (\selectp1[102] , n286, n397);
  and g148 (\selectp1[103] , n288, n397);
  and g149 (\selectp1[104] , n291, n397);
  and g150 (\selectp1[105] , n293, n397);
  and g151 (\selectp1[106] , n296, n397);
  and g152 (\selectp1[107] , n298, n397);
  and g153 (\selectp1[108] , n300, n397);
  and g154 (\selectp1[109] , n302, n397);
  and g155 (\selectp1[110] , n304, n397);
  and g156 (\selectp1[111] , n306, n397);
  and g157 (n414, n344, n362);
  and g158 (\selectp1[112] , n270, n414);
  and g159 (\selectp1[113] , n273, n414);
  and g160 (\selectp1[114] , n276, n414);
  and g161 (\selectp1[115] , n278, n414);
  and g162 (\selectp1[116] , n281, n414);
  and g163 (\selectp1[117] , n284, n414);
  and g164 (\selectp1[118] , n286, n414);
  and g165 (\selectp1[119] , n288, n414);
  and g166 (\selectp1[120] , n291, n414);
  and g167 (\selectp1[121] , n293, n414);
  and g168 (\selectp1[122] , n296, n414);
  and g169 (\selectp1[123] , n298, n414);
  and g170 (\selectp1[124] , n300, n414);
  and g171 (\selectp1[125] , n302, n414);
  and g172 (\selectp1[126] , n304, n414);
  and g173 (\selectp1[127] , n306, n414);
  not g174 (n_16, \count[7] );
  and g175 (n431, n_6, n_16);
  and g176 (n432, n265, n431);
  and g177 (\selectp2[0] , n270, n432);
  and g178 (\selectp2[1] , n273, n432);
  and g179 (\selectp2[2] , n276, n432);
  and g180 (\selectp2[3] , n278, n432);
  and g181 (\selectp2[4] , n281, n432);
  and g182 (\selectp2[5] , n284, n432);
  and g183 (\selectp2[6] , n286, n432);
  and g184 (\selectp2[7] , n288, n432);
  and g185 (\selectp2[8] , n291, n432);
  and g186 (\selectp2[9] , n293, n432);
  and g187 (\selectp2[10] , n296, n432);
  and g188 (\selectp2[11] , n298, n432);
  and g189 (\selectp2[12] , n300, n432);
  and g190 (\selectp2[13] , n302, n432);
  and g191 (\selectp2[14] , n304, n432);
  and g192 (\selectp2[15] , n306, n432);
  and g193 (n449, n308, n431);
  and g194 (\selectp2[16] , n270, n449);
  and g195 (\selectp2[17] , n273, n449);
  and g196 (\selectp2[18] , n276, n449);
  and g197 (\selectp2[19] , n278, n449);
  and g198 (\selectp2[20] , n281, n449);
  and g199 (\selectp2[21] , n284, n449);
  and g200 (\selectp2[22] , n286, n449);
  and g201 (\selectp2[23] , n288, n449);
  and g202 (\selectp2[24] , n291, n449);
  and g203 (\selectp2[25] , n293, n449);
  and g204 (\selectp2[26] , n296, n449);
  and g205 (\selectp2[27] , n298, n449);
  and g206 (\selectp2[28] , n300, n449);
  and g207 (\selectp2[29] , n302, n449);
  and g208 (\selectp2[30] , n304, n449);
  and g209 (\selectp2[31] , n306, n449);
  and g210 (n466, n326, n431);
  and g211 (\selectp2[32] , n270, n466);
  and g212 (\selectp2[33] , n273, n466);
  and g213 (\selectp2[34] , n276, n466);
  and g214 (\selectp2[35] , n278, n466);
  and g215 (\selectp2[36] , n281, n466);
  and g216 (\selectp2[37] , n284, n466);
  and g217 (\selectp2[38] , n286, n466);
  and g218 (\selectp2[39] , n288, n466);
  and g219 (\selectp2[40] , n291, n466);
  and g220 (\selectp2[41] , n293, n466);
  and g221 (\selectp2[42] , n296, n466);
  and g222 (\selectp2[43] , n298, n466);
  and g223 (\selectp2[44] , n300, n466);
  and g224 (\selectp2[45] , n302, n466);
  and g225 (\selectp2[46] , n304, n466);
  and g226 (\selectp2[47] , n306, n466);
  and g227 (n483, n344, n431);
  and g228 (\selectp2[48] , n270, n483);
  and g229 (\selectp2[49] , n273, n483);
  and g230 (\selectp2[50] , n276, n483);
  and g231 (\selectp2[51] , n278, n483);
  and g232 (\selectp2[52] , n281, n483);
  and g233 (\selectp2[53] , n284, n483);
  and g234 (\selectp2[54] , n286, n483);
  and g235 (\selectp2[55] , n288, n483);
  and g236 (\selectp2[56] , n291, n483);
  and g237 (\selectp2[57] , n293, n483);
  and g238 (\selectp2[58] , n296, n483);
  and g239 (\selectp2[59] , n298, n483);
  and g240 (\selectp2[60] , n300, n483);
  and g241 (\selectp2[61] , n302, n483);
  and g242 (\selectp2[62] , n304, n483);
  and g243 (\selectp2[63] , n306, n483);
  and g244 (n500, \count[6] , n_16);
  and g245 (n501, n265, n500);
  and g246 (\selectp2[64] , n270, n501);
  and g247 (\selectp2[65] , n273, n501);
  and g248 (\selectp2[66] , n276, n501);
  and g249 (\selectp2[67] , n278, n501);
  and g250 (\selectp2[68] , n281, n501);
  and g251 (\selectp2[69] , n284, n501);
  and g252 (\selectp2[70] , n286, n501);
  and g253 (\selectp2[71] , n288, n501);
  and g254 (\selectp2[72] , n291, n501);
  and g255 (\selectp2[73] , n293, n501);
  and g256 (\selectp2[74] , n296, n501);
  and g257 (\selectp2[75] , n298, n501);
  and g258 (\selectp2[76] , n300, n501);
  and g259 (\selectp2[77] , n302, n501);
  and g260 (\selectp2[78] , n304, n501);
  and g261 (\selectp2[79] , n306, n501);
  and g262 (n518, n308, n500);
  and g263 (\selectp2[80] , n270, n518);
  and g264 (\selectp2[81] , n273, n518);
  and g265 (\selectp2[82] , n276, n518);
  and g266 (\selectp2[83] , n278, n518);
  and g267 (\selectp2[84] , n281, n518);
  and g268 (\selectp2[85] , n284, n518);
  and g269 (\selectp2[86] , n286, n518);
  and g270 (\selectp2[87] , n288, n518);
  and g271 (\selectp2[88] , n291, n518);
  and g272 (\selectp2[89] , n293, n518);
  and g273 (\selectp2[90] , n296, n518);
  and g274 (\selectp2[91] , n298, n518);
  and g275 (\selectp2[92] , n300, n518);
  and g276 (\selectp2[93] , n302, n518);
  and g277 (\selectp2[94] , n304, n518);
  and g278 (\selectp2[95] , n306, n518);
  and g279 (n535, n326, n500);
  and g280 (\selectp2[96] , n270, n535);
  and g281 (\selectp2[97] , n273, n535);
  and g282 (\selectp2[98] , n276, n535);
  and g283 (\selectp2[99] , n278, n535);
  and g284 (\selectp2[100] , n281, n535);
  and g285 (\selectp2[101] , n284, n535);
  and g286 (\selectp2[102] , n286, n535);
  and g287 (\selectp2[103] , n288, n535);
  and g288 (\selectp2[104] , n291, n535);
  and g289 (\selectp2[105] , n293, n535);
  and g290 (\selectp2[106] , n296, n535);
  and g291 (\selectp2[107] , n298, n535);
  and g292 (\selectp2[108] , n300, n535);
  and g293 (\selectp2[109] , n302, n535);
  and g294 (\selectp2[110] , n304, n535);
  and g295 (\selectp2[111] , n306, n535);
  and g296 (n552, n344, n500);
  and g297 (\selectp2[112] , n270, n552);
  and g298 (\selectp2[113] , n273, n552);
  and g299 (\selectp2[114] , n276, n552);
  and g300 (\selectp2[115] , n278, n552);
  and g301 (\selectp2[116] , n281, n552);
  and g302 (\selectp2[117] , n284, n552);
  and g303 (\selectp2[118] , n286, n552);
  and g304 (\selectp2[119] , n288, n552);
  and g305 (\selectp2[120] , n291, n552);
  and g306 (\selectp2[121] , n293, n552);
  and g307 (\selectp2[122] , n296, n552);
  and g308 (\selectp2[123] , n298, n552);
  and g309 (\selectp2[124] , n300, n552);
  and g310 (\selectp2[125] , n302, n552);
  and g311 (\selectp2[126] , n304, n552);
  and g312 (\selectp2[127] , n306, n552);
endmodule

