
module c3540(N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97,
     N107, N116, N124, N125, N128, N132, N137, N143, N150, N159, N169,
     N179, N190, N200, N213, N222, N223, N226, N232, N238, N244, N250,
     N257, N264, N270, N274, N283, N294, N303, N311, N317, N322, N326,
     N329, N330, N343, N349, N350, N1713, N1947, N3195, N3833, N3987,
     N4028, N4145, N4589, N4667, N4815, N4944, N5002, N5045, N5047,
     N5078, N5102, N5120, N5121, N5192, N5231, N5360, N5361);
//   input N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97,
       N107, N116, N124, N125, N128, N132, N137, N143, N150, N159,
       N169, N179, N190, N200, N213, N222, N223, N226, N232, N238,
       N244, N250, N257, N264, N270, N274, N283, N294, N303, N311,
       N317, N322, N326, N329, N330, N343, N349, N350;
//   output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667,
       N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121,
       N5192, N5231, N5360, N5361;
  wire N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107,
       N116, N124, N125, N128, N132, N137, N143, N150, N159, N169,
       N179, N190, N200, N213, N222, N223, N226, N232, N238, N244,
       N250, N257, N264, N270, N274, N283, N294, N303, N311, N317,
       N322, N326, N329, N330, N343, N349, N350;
  wire N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667,
       N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121,
       N5192, N5231, N5360, N5361;
  wire N665, N679, N686, N702, N724, N736, N749, N763;
  wire N768, N769, N786, N793, N794, N820, N829, N832;
  wire N835, N839, N889, N890, N891, N892, N896, N913;
  wire N914, N920, N1067, N1117, N1179, N1196, N1197, N1202;
  wire N1219, N1250, N1251, N1252, N1253, N1254, N1255, N1256;
  wire N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264;
  wire N1267, N1306, N1315, N1322, N1325, N1328, N1331, N1337;
  wire N1338, N1340, N1343, N1353, N1358, N1366, N1401, N1409;
  wire N1426, N1452, N1460, N1461, N1464, N1467, N1468, N1469;
  wire N1470, N1505, N1507, N1508, N1509, N1510, N1511, N1512;
  wire N1520, N1562, N1579, N1580, N1581, N1586, N1589, N1592;
  wire N1597, N1600, N1643, N1644, N1645, N1646, N1647, N1648;
  wire N1649, N1650, N1667, N1673, N1691, N1692, N1693, N1694;
  wire N1714, N1715, N1718, N1721, N1722, N1725, N1727, N1729;
  wire N1730, N1738, N1747, N1756, N1761, N1770, N1787, N1788;
  wire N1789, N1790, N1791, N1792, N1793, N1794, N1795, N1796;
  wire N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1806;
  wire N1809, N1812, N1815, N1818, N1821, N1824, N1833, N1850;
  wire N1869, N1870, N1873, N1875, N1880, N1885, N1890, N1893;
  wire N1895, N1898, N1900, N1905, N1909, N1912, N1913, N1917;
  wire N1933, N1936, N1940, N1960, N1961, N1966, N1983, N1986;
  wire N1987, N1988, N1989, N1990, N1991, N2022, N2023, N2024;
  wire N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2032;
  wire N2033, N2034, N2035, N2036, N2037, N2043, N2068, N2073;
  wire N2078, N2083, N2088, N2093, N2098, N2103, N2121, N2133;
  wire N2134, N2135, N2136, N2137, N2138, N2139, N2141, N2142;
  wire N2143, N2144, N2145, N2146, N2147, N2148, N2180, N2181;
  wire N2184, N2185, N2188, N2191, N2194, N2197, N2200, N2203;
  wire N2206, N2211, N2230, N2234, N2238, N2239, N2240, N2241;
  wire N2242, N2243, N2244, N2245, N2270, N2277, N2282, N2287;
  wire N2294, N2299, N2307, N2310, N2325, N2328, N2331, N2334;
  wire N2341, N2342, N2347, N2348, N2349, N2350, N2351, N2352;
  wire N2353, N2354, N2355, N2374, N2375, N2376, N2379, N2398;
  wire N2417, N2418, N2419, N2420, N2422, N2425, N2427, N2430;
  wire N2432, N2435, N2436, N2437, N2438, N2439, N2440, N2443;
  wire N2445, N2448, N2450, N2467, N2468, N2471, N2474, N2475;
  wire N2476, N2477, N2478, N2481, N2482, N2483, N2486, N2487;
  wire N2632, N2633, N2641, N2648, N2652, N2656, N2659, N2662;
  wire N2666, N2670, N2673, N2677, N2681, N2684, N2688, N2692;
  wire N2697, N2702, N2706, N2710, N2715, N2719, N2723, N2730;
  wire N2748, N2749, N2754, N2755, N2756, N2757, N2758, N2761;
  wire N2764, N2768, N2769, N2898, N2899, N2900, N2901, N2966;
  wire N2973, N2977, N2980, N2984, N2985, N2986, N2987, N2988;
  wire N2989, N2990, N2991, N3115, N3119, N3125, N3131, N3138;
  wire N3145, N3149, N3155, N3161, N3168, N3172, N3175, N3178;
  wire N3181, N3184, N3187, N3194, N3196, N3206, N3207, N3208;
  wire N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216;
  wire N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224;
  wire N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232;
  wire N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240;
  wire N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248;
  wire N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256;
  wire N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264;
  wire N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3275;
  wire N3276, N3277, N3278, N3279, N3283, N3284, N3285, N3286;
  wire N3287, N3290, N3291, N3292, N3293, N3294, N3295, N3298;
  wire N3299, N3300, N3301, N3302, N3303, N3305, N3306, N3307;
  wire N3308, N3309, N3310, N3311, N3313, N3314, N3315, N3316;
  wire N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324;
  wire N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332;
  wire N3333, N3334, N3383, N3387, N3388, N3389, N3406, N3407;
  wire N3410, N3413, N3414, N3415, N3419, N3423, N3426, N3429;
  wire N3430, N3431, N3434, N3437, N3438, N3439, N3442, N3445;
  wire N3446, N3447, N3451, N3455, N3458, N3461, N3462, N3463;
  wire N3466, N3469, N3470, N3471, N3534, N3535, N3536, N3537;
  wire N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545;
  wire N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3557;
  wire N3568, N3573, N3578, N3589, N3594, N3605, N3627, N3628;
  wire N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639;
  wire N3640, N3641, N3642, N3644, N3645, N3648, N3651, N3652;
  wire N3654, N3657, N3658, N3661, N3663, N3664, N3667, N3670;
  wire N3671, N3673, N3676, N3677, N3680, N3681, N3682, N3685;
  wire N3687, N3689, N3690, N3693, N3694, N3705, N3706, N3711;
  wire N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719;
  wire N3720, N3721, N3731, N3734, N3740, N3743, N3753, N3756;
  wire N3762, N3773, N3775, N3776, N3779, N3780, N3786, N3789;
  wire N3800, N3803, N3809, N3812, N3815, N3818, N3834, N3838;
  wire N3845, N3894, N3895, N3898, N3906, N3912, N3916, N3920;
  wire N3926, N3930, N3931, N3932, N3935, N3936, N3947, N3948;
  wire N3992, N3996, N4013, N4029, N4030, N4031, N4032, N4033;
  wire N4034, N4042, N4043, N4046, N4049, N4050, N4051, N4056;
  wire N4073, N4074, N4075, N4076, N4077, N4078, N4079, N4080;
  wire N4091, N4094, N4104, N4105, N4106, N4107, N4108, N4109;
  wire N4110, N4111, N4112, N4113, N4122, N4146, N4147, N4148;
  wire N4149, N4150, N4151, N4152, N4153, N4186, N4189, N4190;
  wire N4191, N4192, N4193, N4194, N4195, N4196, N4238, N4242;
  wire N4252, N4256, N4283, N4284, N4287, N4291, N4295, N4303;
  wire N4304, N4310, N4317, N4319, N4322, N4325, N4326, N4327;
  wire N4328, N4329, N4331, N4335, N4338, N4341, N4344, N4347;
  wire N4350, N4387, N4390, N4393, N4416, N4421, N4427, N4435;
  wire N4442, N4443, N4446, N4447, N4448, N4458, N4461, N4463;
  wire N4468, N4472, N4475, N4487, N4493, N4496, N4498, N4503;
  wire N4506, N4507, N4508, N4509, N4510, N4511, N4515, N4526;
  wire N4527, N4528, N4530, N4545, N4549, N4552, N4555, N4558;
  wire N4559, N4562, N4572, N4573, N4576, N4588, N4593, N4596;
  wire N4599, N4602, N4608, N4619, N4623, N4629, N4630, N4635;
  wire N4636, N4640, N4641, N4644, N4647, N4650, N4668, N4669;
  wire N4670, N4673, N4674, N4675, N4676, N4677, N4678, N4688;
  wire N4704, N4705, N4706, N4708, N4711, N4716, N4717, N4730;
  wire N4733, N4740, N4743, N4747, N4748, N4753, N4754, N4757;
  wire N4769, N4772, N4775, N4786, N4788, N4794, N4797, N4800;
  wire N4808, N4816, N4817, N4818, N4823, N4829, N4831, N4838;
  wire N4859, N4860, N4868, N4870, N4872, N4880, N4889, N4895;
  wire N4896, N4897, N4900, N4901, N4902, N4904, N4905, N4906;
  wire N4907, N4913, N4916, N4921, N4924, N4926, N4928, N4930;
  wire N4931, N4946, N4950, N4951, N4953, N4954, N4957, N4965;
  wire N4968, N4969, N4970, N4973, N4981, N4982, N4983, N4984;
  wire N4985, N4991, N4999, N5007, N5010, N5013, N5021, N5030;
  wire N5055, N5061, N5066, N5085, N5094, N5108, N5110, N5114;
  wire N5122, N5125, N5128, N5133, N5136, N5145, N5166, N5183;
  wire N5193, N5196, N5201, N5212, N5215, N5217, N5220, N5222;
  wire N5223, N5228, N5232, N5233, N5236, N5242, N5245, N5250;
  wire N5253, N5254, N5258, N5266, N5277, N5278, N5279, N5284;
  wire N5285, N5286, N5295, N5298, N5309, N5340, N5344, N5348;
  wire N5350, N5352, N5354, N5358, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177;
  and AND2_25 (N793, N13, N20);
  and AND2_32 (N829, N33, N41);
  and AND2_53 (N890, N20, N200);
  and AND2_55 (N892, N20, N179);
  and AND2_79 (N1067, N250, N768);
  and AND2_84 (N1202, N913, N914);
  and AND2_110 (N1306, N769, N835);
  and AND2_112 (N1322, N769, N45);
  and AND2_176 (N1520, N50, N1263);
  and AND2_177 (N1562, N1, N1337);
  and AND2_179 (N1580, N794, N1117);
  and AND2_180 (N1581, N1338, N20);
  and AND2_185 (N1586, N686, N20);
  and AND2_188 (N1589, N77, N20);
  and AND2_191 (N1592, N1343, N20);
  and AND2_196 (N1597, N749, N20);
  and AND2_199 (N1600, N116, N20);
  and AND2_200 (N1643, N222, N1401);
  and AND2_201 (N1644, N223, N1401);
  and AND2_202 (N1645, N226, N1401);
  and AND2_203 (N1646, N232, N1401);
  and AND2_204 (N1647, N238, N1401);
  and AND2_205 (N1648, N244, N1401);
  and AND2_206 (N1649, N250, N1401);
  and AND2_207 (N1650, N257, N1401);
  and AND2_223 (N1714, N87, N1264);
  and AND2_227 (N1722, N763, N1340);
  and AND2_232 (N1729, N68, N665);
  and AND2_249 (N1787, N58, N1579);
  and AND2_250 (N1788, N150, N1580);
  and AND2_251 (N1789, N68, N1579);
  and AND2_252 (N1790, N159, N1580);
  and AND2_253 (N1791, N77, N1579);
  and AND2_254 (N1792, N50, N1580);
  and AND2_255 (N1793, N87, N1579);
  and AND2_256 (N1794, N58, N1580);
  and AND2_257 (N1795, N97, N1579);
  and AND2_258 (N1796, N68, N1580);
  and AND2_259 (N1797, N107, N1579);
  and AND2_260 (N1798, N77, N1580);
  and AND2_261 (N1799, N116, N1579);
  and AND2_262 (N1800, N87, N1580);
  and AND2_263 (N1801, N283, N1579);
  and AND2_264 (N1802, N97, N1580);
  and AND2_265 (N1803, N200, N892);
  and AND2_266 (N1806, N889, N892);
  and AND2_267 (N1809, N890, N1366);
  and AND2_268 (N1812, N891, N1366);
  and AND2_282 (N1850, N820, N896);
  and AND2_297 (N1869, N1202, N1409);
  and AND2_321 (N1909, N1452, N213);
  and AND2_341 (N1966, N1520, N839);
  and AND2_344 (N1983, N1067, N1325);
  and AND2_351 (N2022, N77, N33);
  and AND2_352 (N2023, N223, N1850);
  and AND2_353 (N2024, N87, N33);
  and AND2_354 (N2025, N226, N1850);
  and AND2_355 (N2026, N97, N33);
  and AND2_356 (N2027, N232, N1850);
  and AND2_357 (N2028, N107, N33);
  and AND2_358 (N2029, N238, N1850);
  and AND2_359 (N2030, N116, N33);
  and AND2_360 (N2031, N244, N1850);
  and AND2_361 (N2032, N283, N33);
  and AND2_362 (N2033, N250, N1850);
  and AND2_363 (N2034, N294, N33);
  and AND2_364 (N2035, N257, N1850);
  and AND2_365 (N2036, N303, N33);
  and AND2_366 (N2037, N264, N1850);
  and AND2_397 (N2144, N1738, N1747);
  and AND2_416 (N2181, N1756, N1328);
  and AND2_418 (N2184, N1331, N1756);
  and AND2_429 (N2211, N1815, N1818);
  and AND2_448 (N2270, N1986, N1673);
  and AND2_449 (N2277, N1987, N1673);
  and AND2_450 (N2282, N1988, N1673);
  and AND2_451 (N2287, N1989, N1673);
  and AND2_452 (N2294, N1990, N1673);
  and AND2_453 (N2299, N1991, N1673);
  and AND2_455 (N2307, N1464, N350);
  and AND2_467 (N2347, N724, N2144);
  and AND2_469 (N2349, N116, N2147);
  and AND2_470 (N2350, N2148, N839);
  and AND2_471 (N2351, N736, N2144);
  and AND2_472 (N2352, N1947, N2145);
  and AND2_473 (N2353, N763, N2144);
  and AND2_474 (N2354, N1725, N2145);
  and AND2_475 (N2355, N749, N2144);
  and AND2_478 (N2376, N1520, N2180);
  and AND2_479 (N2379, N1721, N2181);
  and AND2_480 (N2398, N665, N2211);
  and AND2_483 (N2419, N1667, N2238);
  and AND2_486 (N2422, N1667, N2239);
  and AND2_489 (N2427, N1667, N2240);
  and AND2_492 (N2432, N1667, N2241);
  and AND2_495 (N2437, N1667, N2242);
  and AND2_498 (N2440, N1667, N2243);
  and AND2_501 (N2445, N1667, N2244);
  and AND2_504 (N2450, N1667, N2245);
  and AND2_516 (N2482, N1761, N1);
  and AND2_517 (N2483, N2349, N2180);
  and AND2_518 (N2486, N2374, N20);
  and AND2_519 (N2487, N2375, N20);
  and AND2_537 (N2633, N1821, N1833);
  and AND2_545 (N2641, N1821, N1824);
  and AND2_574 (N2730, N1562, N1761);
  and AND2_599 (N2758, N1520, N2481);
  and AND2_600 (N2761, N1722, N2482);
  and AND2_601 (N2764, N2478, N1770);
  and AND2_604 (N2898, N665, N2633);
  and AND2_605 (N2899, N679, N2633);
  and AND2_606 (N2900, N686, N2633);
  and AND2_607 (N2901, N702, N2633);
  and AND2_614 (N2980, N2471, N2143);
  and AND2_746 (N3119, N2768, N1673);
  and AND2_758 (N3149, N2769, N1673);
  and AND2_767 (N3172, N1909, N2648);
  and AND2_768 (N3175, N1913, N2662);
  and AND2_769 (N3178, N1913, N2673);
  and AND2_770 (N3181, N1913, N2684);
  and AND2_771 (N3184, N1913, N2702);
  and AND2_772 (N3187, N1913, N2715);
  and AND2_781 (N3207, N124, N2984);
  and AND2_782 (N3208, N159, N2985);
  and AND2_783 (N3209, N150, N2986);
  and AND2_784 (N3210, N143, N2987);
  and AND2_785 (N3211, N137, N2988);
  and AND2_786 (N3212, N132, N2989);
  and AND2_787 (N3213, N128, N2990);
  and AND2_788 (N3214, N125, N2991);
  and AND2_789 (N3215, N125, N2984);
  and AND2_790 (N3216, N50, N2985);
  and AND2_791 (N3217, N159, N2986);
  and AND2_792 (N3218, N150, N2987);
  and AND2_793 (N3219, N143, N2988);
  and AND2_794 (N3220, N137, N2989);
  and AND2_795 (N3221, N132, N2990);
  and AND2_796 (N3222, N128, N2991);
  and AND2_797 (N3223, N128, N2984);
  and AND2_798 (N3224, N58, N2985);
  and AND2_799 (N3225, N50, N2986);
  and AND2_800 (N3226, N159, N2987);
  and AND2_801 (N3227, N150, N2988);
  and AND2_802 (N3228, N143, N2989);
  and AND2_803 (N3229, N137, N2990);
  and AND2_804 (N3230, N132, N2991);
  and AND2_805 (N3231, N132, N2984);
  and AND2_806 (N3232, N68, N2985);
  and AND2_807 (N3233, N58, N2986);
  and AND2_808 (N3234, N50, N2987);
  and AND2_809 (N3235, N159, N2988);
  and AND2_810 (N3236, N150, N2989);
  and AND2_811 (N3237, N143, N2990);
  and AND2_812 (N3238, N137, N2991);
  and AND2_813 (N3239, N137, N2984);
  and AND2_814 (N3240, N77, N2985);
  and AND2_815 (N3241, N68, N2986);
  and AND2_816 (N3242, N58, N2987);
  and AND2_817 (N3243, N50, N2988);
  and AND2_818 (N3244, N159, N2989);
  and AND2_819 (N3245, N150, N2990);
  and AND2_820 (N3246, N143, N2991);
  and AND2_821 (N3247, N143, N2984);
  and AND2_822 (N3248, N87, N2985);
  and AND2_823 (N3249, N77, N2986);
  and AND2_824 (N3250, N68, N2987);
  and AND2_825 (N3251, N58, N2988);
  and AND2_826 (N3252, N50, N2989);
  and AND2_827 (N3253, N159, N2990);
  and AND2_828 (N3254, N150, N2991);
  and AND2_829 (N3255, N150, N2984);
  and AND2_830 (N3256, N97, N2985);
  and AND2_831 (N3257, N87, N2986);
  and AND2_832 (N3258, N77, N2987);
  and AND2_833 (N3259, N68, N2988);
  and AND2_834 (N3260, N58, N2989);
  and AND2_835 (N3261, N50, N2990);
  and AND2_836 (N3262, N159, N2991);
  and AND2_837 (N3263, N159, N2984);
  and AND2_838 (N3264, N107, N2985);
  and AND2_839 (N3265, N97, N2986);
  and AND2_840 (N3266, N87, N2987);
  and AND2_841 (N3267, N77, N2988);
  and AND2_842 (N3268, N68, N2989);
  and AND2_843 (N3269, N58, N2990);
  and AND2_844 (N3270, N50, N2991);
  and AND2_845 (N3271, N283, N2984);
  and AND2_849 (N3275, N87, N2988);
  and AND2_850 (N3276, N97, N2989);
  and AND2_851 (N3277, N107, N2990);
  and AND2_852 (N3278, N116, N2991);
  and AND2_853 (N3279, N294, N2984);
  and AND2_857 (N3283, N97, N2988);
  and AND2_858 (N3284, N107, N2989);
  and AND2_859 (N3285, N116, N2990);
  and AND2_860 (N3286, N283, N2991);
  and AND2_861 (N3287, N303, N2984);
  and AND2_864 (N3290, N97, N2987);
  and AND2_865 (N3291, N107, N2988);
  and AND2_866 (N3292, N116, N2989);
  and AND2_867 (N3293, N283, N2990);
  and AND2_868 (N3294, N294, N2991);
  and AND2_869 (N3295, N311, N2984);
  and AND2_872 (N3298, N107, N2987);
  and AND2_873 (N3299, N116, N2988);
  and AND2_874 (N3300, N283, N2989);
  and AND2_875 (N3301, N294, N2990);
  and AND2_876 (N3302, N303, N2991);
  and AND2_877 (N3303, N317, N2984);
  and AND2_879 (N3305, N107, N2986);
  and AND2_880 (N3306, N116, N2987);
  and AND2_881 (N3307, N283, N2988);
  and AND2_882 (N3308, N294, N2989);
  and AND2_883 (N3309, N303, N2990);
  and AND2_884 (N3310, N311, N2991);
  and AND2_885 (N3311, N322, N2984);
  and AND2_887 (N3313, N116, N2986);
  and AND2_888 (N3314, N283, N2987);
  and AND2_889 (N3315, N294, N2988);
  and AND2_890 (N3316, N303, N2989);
  and AND2_891 (N3317, N311, N2990);
  and AND2_892 (N3318, N317, N2991);
  and AND2_893 (N3319, N326, N2984);
  and AND2_894 (N3320, N116, N2985);
  and AND2_895 (N3321, N283, N2986);
  and AND2_896 (N3322, N294, N2987);
  and AND2_897 (N3323, N303, N2988);
  and AND2_898 (N3324, N311, N2989);
  and AND2_899 (N3325, N317, N2990);
  and AND2_900 (N3326, N322, N2991);
  and AND2_901 (N3327, N329, N2984);
  and AND2_902 (N3328, N283, N2985);
  and AND2_903 (N3329, N294, N2986);
  and AND2_904 (N3330, N303, N2987);
  and AND2_905 (N3331, N311, N2988);
  and AND2_906 (N3332, N317, N2989);
  and AND2_907 (N3333, N322, N2990);
  and AND2_908 (N3334, N326, N2991);
  and AND2_911 (N3387, N3196, N45);
  and AND2_912 (N3388, N2977, N2143);
  and AND2_913 (N3389, N2973, N45);
  and AND2_930 (N3406, N3206, N2641);
  and AND2_1003 (N3605, N3471, N1913);
  and AND2_1010 (N3632, N3536, N2143);
  and AND2_1011 (N3633, N3534, N2143);
  and AND2_1020 (N3642, N3535, N2641);
  and AND2_1044 (N3682, N1909, N3415);
  and AND2_1050 (N3690, N1913, N3447);
  and AND2_1065 (N3713, N3634, N2632);
  and AND2_1066 (N3714, N3635, N2632);
  and AND2_1067 (N3715, N3636, N2632);
  and AND2_1068 (N3716, N3637, N2632);
  and AND2_1069 (N3717, N3638, N2632);
  and AND2_1070 (N3718, N3639, N2632);
  and AND2_1071 (N3719, N3640, N2632);
  and AND2_1072 (N3720, N3641, N2632);
  and AND2_1073 (N3721, N3644, N3557);
  and AND2_1075 (N3734, N3657, N3568);
  and AND2_1076 (N3740, N3661, N3573);
  and AND2_1077 (N3743, N3663, N3578);
  and AND2_1079 (N3756, N3676, N3589);
  and AND2_1080 (N3762, N3680, N3594);
  and AND2_1089 (N3779, N3712, N2641);
  and AND2_1090 (N3780, N3711, N2641);
  and AND2_1095 (N3809, N3654, N1917);
  and AND2_1096 (N3812, N3658, N1917);
  and AND2_1097 (N3815, N3673, N1917);
  and AND2_1098 (N3818, N3677, N1917);
  and AND2_1106 (N3838, N3789, N3731);
  and AND2_1107 (N3845, N3803, N3753);
  and AND2_1122 (N3912, N3786, N1912);
  and AND2_1124 (N3916, N3800, N1917);
  and AND2_1156 (N4028, N3932, N3926);
  and AND2_1178 (N4056, N3932, N1917);
  and AND2_1199 (N4091, N3996, N1917);
  and AND2_1203 (N4104, N4073, N4074);
  and AND2_1238 (N4186, N330, N4094);
  and AND2_1239 (N4189, N4146, N2230);
  and AND2_1241 (N4191, N4148, N2230);
  and AND2_1242 (N4192, N4149, N2230);
  and AND2_1243 (N4193, N4150, N2234);
  and AND2_1245 (N4195, N4152, N2234);
  and AND2_1246 (N4196, N4153, N2234);
  and AND2_1254 (N4238, N4111, N3818);
  and AND2_1257 (N4242, N330, N4112);
  and AND2_1267 (N4283, N4091, N3926);
  and AND2_1268 (N4284, N4094, N3926);
  and AND2_1274 (N4303, N4252, N2230);
  and AND2_1275 (N4304, N4256, N2234);
  and AND2_1279 (N4317, N4094, N4108);
  and AND2_1281 (N4319, N4112, N4111);
  and AND2_1282 (N4322, N4091, N4108);
  and AND2_1305 (N4387, N330, N4317);
  and AND2_1335 (N4493, N330, N4319);
  and AND2_1338 (N4498, N4442, N769);
  and AND2_1357 (N4549, N330, N4443);
  and AND2_1396 (N4647, N4559, N2121);
  and AND2_1397 (N4650, N4559, N2481);
  and AND2_1444 (N4772, N330, N4704);
  and AND2_1451 (N4794, N4711, N2121);
  and AND2_1452 (N4797, N4711, N2481);
  and AND2_1453 (N4800, N4717, N2121);
  and AND2_1455 (N4808, N4717, N4468);
  and AND2_1466 (N4831, N4743, N2121);
  and AND2_1467 (N4838, N4757, N2121);
  and AND2_1493 (N4907, N4818, N2121);
  and AND2_1494 (N4913, N4823, N2121);
  and AND2_1495 (N4916, N4818, N4644);
  and AND2_1497 (N4921, N4895, N2184);
  and AND2_1514 (N4954, N4926, N2481);
  and AND2_1515 (N4957, N4931, N2481);
  and AND2_1521 (N4973, N4953, N2481);
  and AND2_1529 (N4985, N4946, N2121);
  and AND2_1536 (N5010, N4983, N2481);
  and AND2_1537 (N5013, N4984, N2481);
  and AND2_1542 (N5030, N5007, N2481);
  and AND2_1566 (N5114, N5102, N1461);
  and AND2_1572 (N5128, N1461, N5120);
  and AND2_1582 (N5166, N5066, N5133);
  and AND2_1601 (N5215, N213, N5193);
  and AND3_86 (N1250, N665, N679, N686);
  and AND3_111 (N1315, N769, N45, N832);
  and AND3_113 (N1325, N1, N786, N20);
  and AND3_120 (N1340, N724, N736, N749);
  and AND3_148 (N1452, N769, N13, N794);
  and AND3_208 (N1667, N1, N13, N1426);
  and AND3_323 (N1913, N1452, N213, N343);
  and AND3_371 (N2068, N50, N1197, N1869);
  and AND3_372 (N2073, N58, N1197, N1869);
  and AND3_373 (N2078, N68, N1197, N1869);
  and AND3_374 (N2083, N77, N1197, N1869);
  and AND3_375 (N2088, N87, N1219, N1869);
  and AND3_376 (N2093, N97, N1219, N1869);
  and AND3_377 (N2098, N107, N1219, N1869);
  and AND3_378 (N2103, N116, N1219, N1869);
  and AND3_468 (N2348, N2146, N77, N50);
  and AND3_481 (N2417, N2043, N226, N1873);
  and AND3_482 (N2418, N2043, N274, N1306);
  and AND3_484 (N2420, N2043, N232, N1873);
  and AND3_487 (N2425, N2043, N238, N1873);
  and AND3_490 (N2430, N2043, N244, N1873);
  and AND3_493 (N2435, N2043, N250, N1893);
  and AND3_494 (N2436, N2043, N274, N1322);
  and AND3_496 (N2438, N2043, N257, N1898);
  and AND3_497 (N2439, N2043, N274, N1315);
  and AND3_499 (N2443, N2043, N264, N1898);
  and AND3_502 (N2448, N2043, N270, N1898);
  and AND3_931 (N3407, N169, N2648, N2656);
  and AND3_932 (N3410, N179, N2648, N3115);
  and AND3_933 (N3413, N190, N2652, N3115);
  and AND3_934 (N3414, N200, N2652, N2656);
  and AND3_937 (N3423, N169, N2662, N2670);
  and AND3_938 (N3426, N179, N2662, N3131);
  and AND3_939 (N3429, N190, N2666, N3131);
  and AND3_940 (N3430, N200, N2666, N2670);
  and AND3_941 (N3431, N169, N2673, N2681);
  and AND3_942 (N3434, N179, N2673, N3138);
  and AND3_943 (N3437, N190, N2677, N3138);
  and AND3_944 (N3438, N200, N2677, N2681);
  and AND3_945 (N3439, N169, N2684, N2692);
  and AND3_946 (N3442, N179, N2684, N3145);
  and AND3_947 (N3445, N190, N2688, N3145);
  and AND3_948 (N3446, N200, N2688, N2692);
  and AND3_951 (N3455, N169, N2702, N2710);
  and AND3_952 (N3458, N179, N2702, N3161);
  and AND3_953 (N3461, N190, N2706, N3161);
  and AND3_954 (N3462, N200, N2706, N2710);
  and AND3_955 (N3463, N169, N2715, N2723);
  and AND3_956 (N3466, N179, N2715, N3168);
  and AND3_957 (N3469, N190, N2719, N3168);
  and AND3_958 (N3470, N200, N2719, N2723);
  and AND3_1023 (N3645, N169, N3415, N2659);
  and AND3_1024 (N3648, N179, N3415, N3125);
  and AND3_1025 (N3651, N190, N3419, N3125);
  and AND3_1026 (N3652, N200, N3419, N2659);
  and AND3_1034 (N3664, N169, N3447, N2697);
  and AND3_1035 (N3667, N179, N3447, N3155);
  and AND3_1036 (N3670, N190, N3451, N3155);
  and AND3_1037 (N3671, N200, N3451, N2697);
  and AND3_1289 (N4331, N330, N4094, N4295);
  and AND3_1356 (N4545, N330, N4319, N4496);
  and AND3_1381 (N4608, N330, N4284, N4562);
  and AND3_1574 (N5136, N5055, N5085, N1464);
  and AND3_1630 (N5277, N5236, N5254, N2307);
  and AND3_1631 (N5278, N5250, N5254, N2310);
  and AND3_1635 (N5285, N5236, N5266, N2310);
  and AND3_1636 (N5286, N5250, N5266, N2307);
  and AND4_170 (N1507, N1251, N1252, N1253, N1254);
  and AND4_171 (N1508, N1255, N1256, N1257, N1258);
  and AND4_401 (N2148, N1722, N1267, N665, N58);
  and AND4_1130 (N3926, N3721, N3838, N3734, N3740);
  and AND4_1133 (N3932, N3743, N3845, N3756, N3762);
  and AND4_1316 (N4443, N4094, N4190, N4107, N4108);
  and AND4_1488 (N4901, N4717, N4757, N4823, N4468);
  and AND4_1526 (N4982, N4818, N4743, N4946, N4644);
  and AND4_1552 (N5066, N4730, N4999, N5021, N4991);
  and AND4_1573 (N5133, N4880, N5061, N5055, N5085);
  nand NAND2_58 (N913, N1, N13);
  nand NAND2_87 (N1251, N226, N50);
  nand NAND2_88 (N1252, N232, N58);
  nand NAND2_89 (N1253, N238, N68);
  nand NAND2_90 (N1254, N244, N77);
  nand NAND2_91 (N1255, N250, N87);
  nand NAND2_92 (N1256, N257, N97);
  nand NAND2_93 (N1257, N264, N107);
  nand NAND2_94 (N1258, N270, N116);
  nand NAND2_99 (N1263, N679, N686);
  nand NAND2_100 (N1264, N736, N749);
  nand NAND2_101 (N1267, N68, N77);
  nand NAND2_115 (N1331, N1, N786);
  nand NAND2_169 (N1505, N702, N1250);
  nand NAND2_172 (N1509, N232, N1259);
  nand NAND2_173 (N1510, N226, N1260);
  nand NAND2_174 (N1511, N244, N1261);
  nand NAND2_175 (N1512, N238, N1262);
  nand NAND2_218 (N1691, N257, N1467);
  nand NAND2_219 (N1692, N250, N1468);
  nand NAND2_220 (N1693, N270, N1469);
  nand NAND2_221 (N1694, N264, N1470);
  nand NAND2_224 (N1715, N1509, N1510);
  nand NAND2_225 (N1718, N1511, N1512);
  nand NAND2_226 (N1721, N1507, N1508);
  nand NAND2_230 (N1727, N68, N679);
  nand NAND2_233 (N1730, N107, N736);
  nand NAND2_238 (N1738, N1325, N33);
  nand NAND2_239 (N1747, N1325, N820);
  nand NAND2_269 (N1815, N820, N832);
  nand NAND2_270 (N1818, N33, N832);
  nand NAND2_273 (N1833, N786, N820);
  nand NAND2_328 (N1933, N1691, N1692);
  nand NAND2_329 (N1936, N1693, N1694);
  nand NAND2_331 (N1940, N679, N665);
  nand NAND2_339 (N1960, N58, N686);
  nand NAND2_340 (N1961, N97, N749);
  nand NAND2_387 (N2133, N50, N58);
  nand NAND2_388 (N2134, N702, N68);
  nand NAND2_389 (N2135, N686, N77);
  nand NAND2_390 (N2136, N736, N87);
  nand NAND2_391 (N2137, N724, N97);
  nand NAND2_392 (N2138, N763, N107);
  nand NAND2_393 (N2139, N749, N116);
  nand NAND2_399 (N2146, N1727, N1960);
  nand NAND2_400 (N2147, N1730, N1961);
  nand NAND2_419 (N2185, N1358, N1812);
  nand NAND2_420 (N2188, N1358, N1809);
  nand NAND2_421 (N2191, N1353, N1812);
  nand NAND2_422 (N2194, N1353, N1809);
  nand NAND2_423 (N2197, N1358, N1806);
  nand NAND2_424 (N2200, N1358, N1803);
  nand NAND2_425 (N2203, N1353, N1806);
  nand NAND2_426 (N2206, N1353, N1803);
  nand NAND2_461 (N2325, N1940, N2133);
  nand NAND2_462 (N2328, N2134, N2135);
  nand NAND2_463 (N2331, N2136, N2137);
  nand NAND2_464 (N2334, N2138, N2139);
  nand NAND2_465 (N2341, N1936, N2141);
  nand NAND2_466 (N2342, N1933, N2142);
  nand NAND2_509 (N2471, N2341, N2342);
  nand NAND2_591 (N2748, N1718, N2467);
  nand NAND2_592 (N2749, N1715, N2468);
  nand NAND2_595 (N2754, N2328, N2474);
  nand NAND2_596 (N2755, N2325, N2475);
  nand NAND2_597 (N2756, N2334, N2476);
  nand NAND2_598 (N2757, N2331, N2477);
  nand NAND2_609 (N2966, N2748, N2749);
  nand NAND2_612 (N2973, N2754, N2755);
  nand NAND2_613 (N2977, N2756, N2757);
  nand NAND2_1059 (N3705, N2471, N3196);
  nand NAND2_1060 (N3706, N2966, N3627);
  nand NAND2_1083 (N3773, N3705, N3706);
  nand NAND2_1085 (N3775, N2977, N3628);
  nand NAND2_1104 (N3834, N2973, N3776);
  nand NAND2_1114 (N3987, N3775, N3834);
  nand NAND2_1116 (N3894, N3721, N3786);
  nand NAND2_1117 (N3895, N3743, N3800);
  nand NAND2_1157 (N4029, N3721, N3681);
  nand NAND2_1158 (N4030, N3734, N3685);
  nand NAND2_1159 (N4031, N3740, N3687);
  nand NAND2_1160 (N4032, N3743, N3689);
  nand NAND2_1161 (N4033, N3756, N3693);
  nand NAND2_1162 (N4034, N3762, N3694);
  nand NAND2_1187 (N4073, N3926, N3996);
  nand NAND2_1189 (N4075, N3172, N4042);
  nand NAND2_1190 (N4076, N3175, N4043);
  nand NAND2_1191 (N4077, N3178, N4046);
  nand NAND2_1192 (N4078, N3181, N4049);
  nand NAND2_1193 (N4079, N3184, N4050);
  nand NAND2_1194 (N4080, N3187, N4051);
  nand NAND2_1204 (N4105, N4075, N4029);
  nand NAND2_1205 (N4106, N3838, N3898);
  nand NAND2_1206 (N4107, N4076, N4030);
  nand NAND2_1207 (N4108, N4077, N4031);
  nand NAND2_1208 (N4109, N4078, N4032);
  nand NAND2_1209 (N4110, N3845, N3906);
  nand NAND2_1210 (N4111, N4079, N4033);
  nand NAND2_1211 (N4112, N4080, N4034);
  nand NAND2_1226 (N4147, N3682, N4113);
  nand NAND2_1230 (N4151, N3690, N4122);
  nand NAND2_1240 (N4190, N4147, N4106);
  nand NAND2_1244 (N4194, N4151, N4110);
  nand NAND2_1283 (N4325, N4107, N3812);
  nand NAND2_1285 (N4327, N4194, N3815);
  nand NAND2_1287 (N4329, N4111, N4013);
  nand NAND2_1307 (N4393, N3818, N4152);
  nand NAND2_1317 (N4446, N4190, N3809);
  nand NAND2_1321 (N4458, N4329, N4393);
  nand NAND2_1324 (N4463, N4112, N1460);
  nand NAND2_1333 (N4487, N4108, N4295);
  nand NAND2_1343 (N4509, N4421, N4148);
  nand NAND2_1345 (N4511, N4427, N4150);
  nand NAND2_1346 (N4515, N330, N4153);
  nand NAND2_1348 (N4527, N4416, N4252);
  nand NAND2_1349 (N4528, N4091, N4149);
  nand NAND2_1351 (N4530, N4287, N4256);
  nand NAND2_1358 (N4552, N4107, N4508);
  nand NAND2_1359 (N4555, N4109, N4510);
  nand NAND2_1361 (N4559, N4463, N4515);
  nand NAND2_1367 (N4572, N4190, N4526);
  nand NAND2_1368 (N4573, N4194, N4496);
  nand NAND2_1369 (N4576, N4487, N4528);
  nand NAND2_1375 (N4593, N4552, N4509);
  nand NAND2_1378 (N4599, N4555, N4511);
  nand NAND2_1384 (N4619, N4572, N4527);
  nand NAND2_1385 (N4623, N4573, N4530);
  nand NAND2_1387 (N4629, N4443, N4506);
  nand NAND2_1390 (N4636, N4576, N4291);
  nand NAND2_1392 (N4641, N4458, N4461);
  nand NAND2_1402 (N4668, N4284, N4630);
  nand NAND2_1404 (N4670, N4503, N4146);
  nand NAND2_1406 (N4674, N4619, N4507);
  nand NAND2_1407 (N4675, N4186, N4635);
  nand NAND2_1409 (N4677, N4623, N4558);
  nand NAND2_1410 (N4678, N4242, N4640);
  nand NAND2_1413 (N4688, N4503, N4562);
  nand NAND2_1418 (N4704, N4629, N4668);
  nand NAND2_1419 (N4705, N4105, N4669);
  nand NAND2_1422 (N4708, N4435, N4673);
  nand NAND2_1423 (N4711, N4675, N4636);
  nand NAND2_1424 (N4716, N4493, N4676);
  nand NAND2_1425 (N4717, N4678, N4641);
  nand NAND2_1431 (N4733, N4310, N4669);
  nand NAND2_1432 (N4740, N4705, N4670);
  nand NAND2_1433 (N4743, N4708, N4674);
  nand NAND2_1435 (N4748, N4593, N4596);
  nand NAND2_1439 (N4754, N4599, N4602);
  nand NAND2_1442 (N4757, N4716, N4677);
  nand NAND2_1443 (N4769, N4733, N4688);
  nand NAND2_1447 (N4786, N4387, N4747);
  nand NAND2_1449 (N4788, N4390, N4753);
  nand NAND2_1460 (N4818, N4786, N4748);
  nand NAND2_1462 (N4823, N4788, N4754);
  nand NAND2_1464 (N4829, N4775, N4442);
  nand NAND2_1472 (N4859, N4772, N4816);
  nand NAND2_1473 (N4860, N4769, N4817);
  nand NAND2_1482 (N4895, N4859, N4860);
  nand NAND2_1484 (N4897, N4740, N4706);
  nand NAND2_1491 (N4905, N4757, N4872);
  nand NAND2_1492 (N4906, N4872, N4829);
  nand NAND2_1498 (N4924, N4549, N4896);
  nand NAND2_1501 (N4928, N4889, N4870);
  nand NAND2_1503 (N4930, N4808, N4904);
  nand NAND2_1508 (N4946, N4924, N4897);
  nand NAND2_1510 (N4950, N4916, N4902);
  nand NAND2_1513 (N4953, N4930, N4905);
  nand NAND2_1519 (N4969, N4743, N4951);
  nand NAND2_1520 (N4970, N4951, N4928);
  nand NAND2_1527 (N4983, N4950, N4969);
  nand NAND2_1557 (N5094, N5047, N4730);
  nand NAND2_1562 (N5108, N4815, N4999);
  nand NAND2_1564 (N5110, N5078, N4991);
  nand NAND2_1570 (N5122, N5094, N5108);
  nand NAND2_1571 (N5125, N5045, N5021);
  nand NAND2_1576 (N5145, N5125, N5110);
  nand NAND2_1587 (N5183, N5120, N5055);
  nand NAND2_1592 (N5196, N5121, N4880);
  nand NAND2_1600 (N5212, N5102, N5085);
  nand NAND2_1604 (N5220, N4944, N5061);
  nand NAND2_1607 (N5223, N5128, N5201);
  nand NAND2_1610 (N5228, N5183, N5212);
  nand NAND2_1612 (N5232, N5145, N5217);
  nand NAND2_1616 (N5236, N5196, N5220);
  nand NAND2_1618 (N5242, N5114, N5222);
  nand NAND2_1620 (N5245, N5122, N5233);
  nand NAND2_1624 (N5254, N5242, N5223);
  nand NAND2_1626 (N5258, N5232, N5245);
  nand NAND2_1634 (N5284, N5236, N5253);
  nand NAND2_1639 (N5295, N5228, N5250);
  nand NAND2_1643 (N5309, N5295, N5284);
  nand NAND2_1652 (N5340, N5298, N5258);
  nand NAND2_1656 (N5348, N5309, N5279);
  nand NAND2_1658 (N5350, N5279, N5344);
  nand NAND2_1662 (N5354, N5258, N5352);
  nand NAND2_1664 (N5360, N5350, N5340);
  nand NAND2_1666 (N5358, N5348, N5354);
  nand NAND3_59 (N914, N1, N20, N33);
  nand NAND3_117 (N1337, N13, N794, N45);
  nand NAND3_240 (N1756, N1, N13, N20);
  nand NAND3_271 (N1821, N1, N13, N1179);
  nand NAND3_272 (N1824, N786, N794, N820);
  nand NAND3_1131 (N3930, N3721, N3838, N3654);
  nand NAND3_1134 (N3935, N3743, N3845, N3673);
  nand NAND3_1284 (N4326, N4107, N4108, N4091);
  nand NAND3_1286 (N4328, N4194, N4111, N3818);
  nand NAND3_1310 (N4416, N3920, N4325, N4326);
  nand NAND3_1312 (N4427, N3948, N4327, N4328);
  nand NAND3_1318 (N4447, N4190, N4107, N3812);
  nand NAND4_241 (N1761, N1, N786, N20, N832);
  nand NAND4_1132 (N3931, N3658, N3838, N3734, N3721);
  nand NAND4_1135 (N3936, N3677, N3845, N3756, N3743);
  nand NAND4_1153 (N3992, N3644, N3894, N3930, N3931);
  nand NAND4_1154 (N3996, N3663, N3895, N3935, N3936);
  nand NAND4_1319 (N4448, N4190, N4107, N4108, N4091);
  nand NAND4_1339 (N4503, N3947, N4446, N4447, N4448);
  nor NOR2_132 (N1358, N794, N190);
  nor NOR2_152 (N1464, N920, N343);
  nor NOR2_298 (N1870, N50, N1409);
  nor NOR2_301 (N1875, N58, N1409);
  nor NOR2_304 (N1880, N68, N1409);
  nor NOR2_307 (N1885, N77, N1409);
  nor NOR2_310 (N1890, N87, N1409);
  nor NOR2_313 (N1895, N97, N1409);
  nor NOR2_316 (N1900, N107, N1409);
  nor NOR2_319 (N1905, N116, N1409);
  nor NOR2_978 (N3534, N3387, N2350);
  nor NOR2_980 (N3536, N3389, N1966);
  nor NOR2_1022 (N3644, N3407, N3410);
  nor NOR2_1029 (N3657, N3423, N3426);
  nor NOR2_1031 (N3661, N3431, N3434);
  nor NOR2_1033 (N3663, N3439, N3442);
  nor NOR2_1040 (N3676, N3455, N3458);
  nor NOR2_1042 (N3680, N3463, N3466);
  nor NOR2_1092 (N3789, N3645, N3648);
  nor NOR2_1094 (N3803, N3664, N3667);
  nor NOR2_1327 (N4468, N4331, N4091);
  nor NOR2_1395 (N4644, N4608, N4310);
  nor NOR2_1487 (N4900, N4868, N4468);
  nor NOR2_1525 (N4981, N4968, N4644);
  nor NOR2_1591 (N5193, N5136, N5166);
  nor NOR3_553 (N2652, N2270, N1870, N2068);
  nor NOR3_557 (N2666, N2277, N1880, N2078);
  nor NOR3_560 (N2677, N2282, N1885, N2083);
  nor NOR3_563 (N2688, N2287, N1890, N2088);
  nor NOR3_567 (N2706, N2294, N1900, N2098);
  nor NOR3_570 (N2719, N2299, N1905, N2103);
  nor NOR3_590 (N3195, N2376, N1983, N2379);
  nor NOR3_936 (N3419, N3119, N1875, N2073);
  nor NOR3_950 (N3451, N3149, N1895, N2093);
  nor NOR3_1373 (N4588, N2758, N4498, N2761);
  nor NOR3_1430 (N4730, N4647, N4650, N4350);
  nor NOR3_1479 (N4880, N4794, N4797, N4341);
  nor NOR3_1517 (N4965, N2764, N2483, N4921);
  nor NOR3_1531 (N4991, N4913, N4954, N4344);
  nor NOR3_1533 (N4999, N4800, N4957, N4347);
  nor NOR3_1539 (N5021, N4838, N4973, N4475);
  nor NOR3_1549 (N5055, N4831, N5010, N4472);
  nor NOR3_1551 (N5061, N4907, N5013, N4338);
  nor NOR3_1556 (N5085, N4985, N5030, N4335);
  not NOT1_2 (N665, N50);
  not NOT1_4 (N679, N58);
  not NOT1_6 (N686, N68);
  not NOT1_9 (N702, N77);
  not NOT1_12 (N724, N87);
  not NOT1_14 (N736, N97);
  not NOT1_16 (N749, N107);
  not NOT1_18 (N763, N116);
  not NOT1_20 (N769, N1);
  not NOT1_24 (N786, N13);
  not NOT1_26 (N794, N20);
  not NOT1_29 (N820, N33);
  not NOT1_33 (N832, N41);
  not NOT1_36 (N839, N45);
  not NOT1_52 (N889, N200);
  not NOT1_63 (N920, N213);
  not NOT1_82 (N1196, N793);
  not NOT1_95 (N1259, N226);
  not NOT1_96 (N1260, N232);
  not NOT1_97 (N1261, N238);
  not NOT1_98 (N1262, N244);
  not NOT1_134 (N1366, N892);
  not NOT1_137 (N1401, N896);
  not NOT1_146 (N1426, N829);
  not NOT1_150 (N1460, N330);
  not NOT1_153 (N1467, N250);
  not NOT1_154 (N1468, N257);
  not NOT1_155 (N1469, N264);
  not NOT1_156 (N1470, N270);
  not NOT1_178 (N1579, N1117);
  not NOT1_210 (N1673, N1202);
  not NOT1_222 (N1713, N1505);
  not NOT1_248 (N1770, N1331);
  not NOT1_299 (N1873, N1306);
  not NOT1_311 (N1893, N1322);
  not NOT1_314 (N1898, N1315);
  not NOT1_338 (N1947, N1714);
  not NOT1_368 (N2043, N1667);
  not NOT1_379 (N2121, N1562);
  not NOT1_394 (N2141, N1933);
  not NOT1_395 (N2142, N1936);
  not NOT1_396 (N2143, N1738);
  not NOT1_398 (N2145, N1747);
  not NOT1_415 (N2180, N1756);
  not NOT1_432 (N2230, N1833);
  not NOT1_436 (N2234, N1824);
  not NOT1_476 (N2374, N2146);
  not NOT1_477 (N2375, N2147);
  not NOT1_505 (N2467, N1715);
  not NOT1_506 (N2468, N1718);
  not NOT1_510 (N2474, N2325);
  not NOT1_511 (N2475, N2328);
  not NOT1_512 (N2476, N2331);
  not NOT1_513 (N2477, N2334);
  not NOT1_515 (N2481, N1761);
  not NOT1_536 (N2632, N1821);
  not NOT1_615 (N2984, N2185);
  not NOT1_616 (N2985, N2188);
  not NOT1_617 (N2986, N2191);
  not NOT1_618 (N2987, N2194);
  not NOT1_619 (N2988, N2197);
  not NOT1_620 (N2989, N2200);
  not NOT1_621 (N2990, N2203);
  not NOT1_622 (N2991, N2206);
  not NOT1_744 (N3115, N2656);
  not NOT1_745 (N2648, N2652);
  not NOT1_748 (N3125, N2659);
  not NOT1_750 (N3131, N2670);
  not NOT1_751 (N2662, N2666);
  not NOT1_753 (N3138, N2681);
  not NOT1_754 (N2673, N2677);
  not NOT1_756 (N3145, N2692);
  not NOT1_757 (N2684, N2688);
  not NOT1_760 (N3155, N2697);
  not NOT1_762 (N3161, N2710);
  not NOT1_763 (N2702, N2706);
  not NOT1_765 (N3168, N2723);
  not NOT1_766 (N2715, N2719);
  not NOT1_779 (N3196, N2966);
  not NOT1_1005 (N3627, N2471);
  not NOT1_1006 (N3628, N2973);
  not NOT1_1027 (N3415, N3419);
  not NOT1_1038 (N3447, N3451);
  not NOT1_1043 (N3681, N3172);
  not NOT1_1045 (N3685, N3175);
  not NOT1_1047 (N3687, N3178);
  not NOT1_1049 (N3689, N3181);
  not NOT1_1051 (N3693, N3184);
  not NOT1_1052 (N3694, N3187);
  not NOT1_1086 (N3776, N2977);
  not NOT1_1118 (N3898, N3682);
  not NOT1_1120 (N3906, N3690);
  not NOT1_1126 (N3920, N3809);
  not NOT1_1138 (N3947, N3912);
  not NOT1_1139 (N3948, N3916);
  not NOT1_1155 (N4013, N3818);
  not NOT1_1164 (N4042, N3721);
  not NOT1_1165 (N4043, N3734);
  not NOT1_1168 (N4046, N3740);
  not NOT1_1171 (N4049, N3743);
  not NOT1_1172 (N4050, N3756);
  not NOT1_1173 (N4051, N3762);
  not NOT1_1188 (N4074, N3992);
  not NOT1_1212 (N4113, N3838);
  not NOT1_1217 (N4122, N3845);
  not NOT1_1224 (N4145, N4104);
  not NOT1_1225 (N4146, N4105);
  not NOT1_1227 (N4148, N4107);
  not NOT1_1228 (N4149, N4108);
  not NOT1_1229 (N4150, N4109);
  not NOT1_1231 (N4152, N4111);
  not NOT1_1232 (N4153, N4112);
  not NOT1_1260 (N4252, N4190);
  not NOT1_1264 (N4256, N4194);
  not NOT1_1270 (N4291, N4186);
  not NOT1_1271 (N4295, N4091);
  not NOT1_1322 (N4461, N4242);
  not NOT1_1336 (N4496, N4287);
  not NOT1_1340 (N4506, N4284);
  not NOT1_1341 (N4507, N4435);
  not NOT1_1342 (N4508, N4421);
  not NOT1_1344 (N4510, N4427);
  not NOT1_1347 (N4526, N4416);
  not NOT1_1360 (N4558, N4493);
  not NOT1_1362 (N4562, N4310);
  not NOT1_1376 (N4596, N4387);
  not NOT1_1379 (N4602, N4390);
  not NOT1_1386 (N4667, N4588);
  not NOT1_1388 (N4630, N4443);
  not NOT1_1389 (N4635, N4576);
  not NOT1_1391 (N4640, N4458);
  not NOT1_1403 (N4669, N4503);
  not NOT1_1405 (N4673, N4619);
  not NOT1_1408 (N4676, N4623);
  not NOT1_1420 (N4706, N4549);
  not NOT1_1428 (N4442, N4468);
  not NOT1_1434 (N4747, N4593);
  not NOT1_1438 (N4753, N4599);
  not NOT1_1445 (N4775, N4717);
  not NOT1_1446 (N4815, N4730);
  not NOT1_1458 (N4816, N4769);
  not NOT1_1459 (N4817, N4772);
  not NOT1_1474 (N4868, N4823);
  not NOT1_1475 (N4870, N4644);
  not NOT1_1476 (N4872, N4808);
  not NOT1_1481 (N4889, N4818);
  not NOT1_1483 (N4896, N4740);
  not NOT1_1489 (N4902, N4743);
  not NOT1_1490 (N4904, N4757);
  not NOT1_1496 (N4944, N4880);
  not NOT1_1504 (N4931, N4906);
  not NOT1_1511 (N4951, N4916);
  not NOT1_1518 (N4968, N4946);
  not NOT1_1524 (N5002, N4965);
  not NOT1_1528 (N4984, N4970);
  not NOT1_1540 (N5045, N4991);
  not NOT1_1541 (N5047, N4999);
  not NOT1_1546 (N5078, N5021);
  not NOT1_1561 (N5121, N5061);
  not NOT1_1590 (N5192, N5166);
  not NOT1_1596 (N5201, N5114);
  not NOT1_1602 (N5217, N5122);
  not NOT1_1606 (N5222, N5128);
  not NOT1_1611 (N5231, N5215);
  not NOT1_1613 (N5233, N5145);
  not NOT1_1622 (N5250, N5236);
  not NOT1_1623 (N5253, N5228);
  not NOT1_1628 (N5266, N5254);
  not NOT1_1632 (N5279, N5258);
  not NOT1_1654 (N5344, N5298);
  not NOT1_1660 (N5352, N5309);
  or OR2_19 (N768, N257, N264);
  or OR2_34 (N835, N41, N45);
  or OR2_57 (N896, N349, N33);
  or OR2_80 (N1117, N820, N20);
  or OR2_81 (N1179, N794, N169);
  or OR2_83 (N1197, N794, N1);
  or OR2_85 (N1219, N820, N1);
  or OR2_145 (N1409, N1, N1196);
  or OR2_514 (N2478, N2348, N1729);
  or OR2_959 (N3471, N3194, N3383);
  or OR2_1013 (N3635, N3539, N3540);
  or OR2_1014 (N3636, N3541, N3542);
  or OR2_1015 (N3637, N3543, N3544);
  or OR2_1016 (N3638, N3545, N3546);
  or OR2_1017 (N3639, N3547, N3548);
  or OR2_1018 (N3640, N3549, N3550);
  or OR2_1019 (N3641, N3551, N3552);
  or OR2_1200 (N4094, N3605, N4056);
  or OR2_1269 (N4287, N3815, N4238);
  or OR2_1277 (N4310, N3992, N4283);
  or OR2_1311 (N4421, N3812, N4322);
  or OR2_1374 (N4589, N4545, N4287);
  or OR2_1500 (N4926, N4900, N4901);
  or OR2_1535 (N5007, N4981, N4982);
  or OR3_345 (N1986, N1581, N1787, N1788);
  or OR3_346 (N1987, N1586, N1791, N1792);
  or OR3_347 (N1988, N1589, N1793, N1794);
  or OR3_348 (N1989, N1592, N1795, N1796);
  or OR3_349 (N1990, N1597, N1799, N1800);
  or OR3_350 (N1991, N1600, N1801, N1802);
  or OR3_440 (N2238, N2022, N1643, N2023);
  or OR3_441 (N2239, N2024, N1644, N2025);
  or OR3_442 (N2240, N2026, N1645, N2027);
  or OR3_443 (N2241, N2028, N1646, N2029);
  or OR3_444 (N2242, N2030, N1647, N2031);
  or OR3_445 (N2243, N2032, N1648, N2033);
  or OR3_446 (N2244, N2034, N1649, N2035);
  or OR3_447 (N2245, N2036, N1650, N2037);
  or OR3_554 (N2656, N2417, N2418, N2419);
  or OR3_555 (N2659, N2420, N2418, N2422);
  or OR3_558 (N2670, N2425, N2418, N2427);
  or OR3_561 (N2681, N2430, N2418, N2432);
  or OR3_564 (N2692, N2435, N2436, N2437);
  or OR3_565 (N2697, N2438, N2439, N2440);
  or OR3_568 (N2710, N2443, N2439, N2445);
  or OR3_571 (N2723, N2448, N2439, N2450);
  or OR3_602 (N2768, N2486, N1789, N1790);
  or OR3_603 (N2769, N2487, N1797, N1798);
  or OR3_780 (N3206, N2980, N2145, N2347);
  or OR3_979 (N3535, N3388, N2145, N2351);
  or OR3_997 (N3557, N3413, N3414, N2648);
  or OR3_998 (N3568, N3429, N3430, N2662);
  or OR3_999 (N3573, N3437, N3438, N2673);
  or OR3_1000 (N3578, N3445, N3446, N2684);
  or OR3_1001 (N3589, N3461, N3462, N2702);
  or OR3_1002 (N3594, N3469, N3470, N2715);
  or OR3_1012 (N3634, N3537, N3538, N2398);
  or OR3_1063 (N3711, N3632, N2352, N2353);
  or OR3_1064 (N3712, N3633, N2354, N2355);
  or OR3_1074 (N3731, N3651, N3652, N3415);
  or OR3_1078 (N3753, N3670, N3671, N3447);
  or OR4_1640 (N5298, N5277, N5285, N5278, N5286);
  not g1 (N3833, N3773);
  not g2 (N5361, N5358);
  and g3 (n_74, n_73, N2692);
  not g4 (n_73, N179);
  and g5 (N3194, N2697, N2710, N2723, n_74);
  and g6 (n_75, N3145, N3155);
  and g7 (N3383, N3161, N3168, N179, n_75);
  and g8 (N4350, n_76, n_77, n_78, N2730);
  not g9 (n_76, N3720);
  not g10 (n_77, N4196);
  not g11 (n_78, N3780);
  nor g12 (n_80, N3263, N3264, N3265);
  nor g13 (n_81, N3266, N3267);
  nor g14 (n_82, N3268, N3269);
  and g15 (n_83, n_79, N820);
  not g16 (n_79, N3270);
  and g17 (N3551, n_80, n_81, n_82, n_83);
  nor g18 (n_85, N3327, N3328, N3329);
  nor g19 (n_86, N3330, N3331);
  nor g20 (n_87, N3332, N3333);
  and g21 (n_88, n_84, N33);
  not g22 (n_84, N3334);
  and g23 (N3552, n_85, n_86, n_87, n_88);
  and g24 (N4341, n_89, n_90, n_91, N2730);
  not g25 (n_89, N3716);
  not g26 (n_90, N4192);
  not g27 (n_91, N2901);
  nor g28 (n_93, N3231, N3232, N3233);
  nor g29 (n_94, N3234, N3235);
  nor g30 (n_95, N3236, N3237);
  and g31 (n_96, n_92, N820);
  not g32 (n_92, N3238);
  and g33 (N3543, n_93, n_94, n_95, n_96);
  nor g34 (n_98, N3295, N3248, N3265);
  nor g35 (n_99, N3298, N3299);
  nor g36 (n_100, N3300, N3301);
  and g37 (n_101, n_97, N33);
  not g38 (n_97, N3302);
  and g39 (N3544, n_98, n_99, n_100, n_101);
  and g40 (N4344, n_102, n_103, n_104, N2730);
  not g41 (n_102, N3717);
  not g42 (n_103, N4193);
  not g43 (n_104, N3406);
  and g44 (N4390, N330, N4112, N4111, N4194);
  nor g45 (n_106, N3239, N3240, N3241);
  nor g46 (n_107, N3242, N3243);
  nor g47 (n_108, N3244, N3245);
  and g48 (n_109, n_105, N820);
  not g49 (n_105, N3246);
  and g50 (N3545, n_106, n_107, n_108, n_109);
  nor g51 (n_111, N3303, N3256, N3305);
  nor g52 (n_112, N3306, N3307);
  nor g53 (n_113, N3308, N3309);
  and g54 (n_114, n_110, N33);
  not g55 (n_110, N3310);
  and g56 (N3546, n_111, n_112, n_113, n_114);
  and g57 (N4347, n_115, n_116, n_117, N2730);
  not g58 (n_115, N3719);
  not g59 (n_116, N4195);
  not g60 (n_117, N3779);
  nor g61 (n_119, N3255, N3256, N3257);
  nor g62 (n_120, N3258, N3259);
  nor g63 (n_121, N3260, N3261);
  and g64 (n_122, n_118, N820);
  not g65 (n_118, N3262);
  and g66 (N3549, n_119, n_120, n_121, n_122);
  nor g67 (n_124, N3319, N3320, N3321);
  nor g68 (n_125, N3322, N3323);
  nor g69 (n_126, N3324, N3325);
  and g70 (n_127, n_123, N33);
  not g71 (n_123, N3326);
  and g72 (N3550, n_124, n_125, n_126, n_127);
  and g73 (N4475, n_128, n_129, n_130, N2730);
  not g74 (n_128, N3718);
  not g75 (n_129, N4304);
  not g76 (n_130, N3642);
  nor g77 (n_132, N3247, N3248, N3249);
  nor g78 (n_133, N3250, N3251);
  nor g79 (n_134, N3252, N3253);
  and g80 (n_135, n_131, N820);
  not g81 (n_131, N3254);
  and g82 (N3547, n_132, n_133, n_134, n_135);
  nor g83 (n_137, N3311, N3264, N3313);
  nor g84 (n_138, N3314, N3315);
  nor g85 (n_139, N3316, N3317);
  and g86 (n_140, n_136, N33);
  not g87 (n_136, N3318);
  and g88 (N3548, n_137, n_138, n_139, n_140);
  and g89 (N4472, n_141, n_142, n_143, N2730);
  not g90 (n_141, N3714);
  not g91 (n_142, N4303);
  not g92 (n_143, N2899);
  and g93 (N4435, N330, N4094, N4108, N4107);
  nor g94 (n_145, N3215, N3216, N3217);
  nor g95 (n_146, N3218, N3219);
  nor g96 (n_147, N3220, N3221);
  and g97 (n_148, n_144, N820);
  not g98 (n_144, N3222);
  and g99 (N3539, n_145, n_146, n_147, n_148);
  nor g100 (n_150, N3279, N3232, N3249);
  nor g101 (n_151, N3266, N3283);
  nor g102 (n_152, N3284, N3285);
  and g103 (n_153, n_149, N33);
  not g104 (n_149, N3286);
  and g105 (N3540, n_150, n_151, n_152, n_153);
  and g106 (N4335, n_154, n_155, n_156, N2730);
  not g107 (n_154, N3713);
  not g108 (n_155, N4189);
  not g109 (n_156, N2898);
  nor g110 (n_157, N3207, N3208, N3209);
  nor g111 (n_158, N3210, N3211);
  nor g112 (n_159, N3212, N3213);
  nor g113 (n_160, N3214, N1815);
  and g114 (N3537, n_157, n_158, n_159, n_160);
  nor g115 (n_161, N3271, N3224, N3241);
  nor g116 (n_162, N3258, N3275);
  nor g117 (n_163, N3276, N3277);
  nor g118 (n_164, N3278, N1818);
  and g119 (N3538, n_161, n_162, n_163, n_164);
  and g120 (N4338, n_165, n_166, n_167, N2730);
  not g121 (n_165, N3715);
  not g122 (n_166, N4191);
  not g123 (n_167, N2900);
  nor g124 (n_169, N3223, N3224, N3225);
  nor g125 (n_170, N3226, N3227);
  nor g126 (n_171, N3228, N3229);
  and g127 (n_172, n_168, N820);
  not g128 (n_168, N3230);
  and g129 (N3541, n_169, n_170, n_171, n_172);
  nor g130 (n_174, N3287, N3240, N3257);
  nor g131 (n_175, N3290, N3291);
  nor g132 (n_176, N3292, N3293);
  and g133 (n_177, n_173, N33);
  not g134 (n_173, N3294);
  and g135 (N3542, n_174, n_175, n_176, n_177);
  not g136 (N891, N890);
  not g138 (N1725, N1722);
  not g139 (N1912, N1909);
  not g140 (N2310, N2307);
  not g143 (N1338, N1250);
  not g144 (N1328, N1325);
  not g145 (N1343, N1340);
  not g146 (N1917, N1913);
  not g147 (N1353, N1358);
  not g148 (N1461, N1464);
  not g150 (N3654, N3657);
  not g151 (N3658, N3661);
  not g153 (N3673, N3676);
  not g154 (N3677, N3680);
  not g155 (N3786, N3789);
  not g156 (N3800, N3803);
  not g174 (N5102, N5055);
  not g176 (N5120, N5085);
endmodule

