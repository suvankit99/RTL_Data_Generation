
module sin(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] ,
     \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14]
     , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
     \a[22] , \a[23] , \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4]
     , \sin[5] , \sin[6] , \sin[7] , \sin[8] , \sin[9] , \sin[10] ,
     \sin[11] , \sin[12] , \sin[13] , \sin[14] , \sin[15] , \sin[16] ,
     \sin[17] , \sin[18] , \sin[19] , \sin[20] , \sin[21] , \sin[22] ,
     \sin[23] , \sin[24] );
  input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] ,
       \sin[6] , \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] ,
       \sin[12] , \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17]
       , \sin[18] , \sin[19] , \sin[20] , \sin[21] , \sin[22] ,
       \sin[23] , \sin[24] ;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] ;
  wire \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] ,
       \sin[6] , \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] ,
       \sin[12] , \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17]
       , \sin[18] , \sin[19] , \sin[20] , \sin[21] , \sin[22] ,
       \sin[23] , \sin[24] ;
  wire n50, n51, n52, n53, n54, n55, n56, n57;
  wire n58, n59, n60, n61, n62, n63, n64, n65;
  wire n66, n67, n68, n69, n70, n71, n72, n73;
  wire n74, n75, n76, n77, n78, n79, n80, n81;
  wire n82, n83, n84, n85, n86, n87, n88, n89;
  wire n90, n91, n92, n93, n94, n95, n96, n97;
  wire n98, n99, n100, n101, n102, n103, n104, n105;
  wire n106, n107, n108, n109, n110, n111, n112, n113;
  wire n114, n115, n116, n117, n118, n119, n120, n121;
  wire n122, n123, n124, n125, n126, n127, n128, n129;
  wire n130, n131, n132, n133, n134, n135, n136, n137;
  wire n138, n139, n140, n141, n142, n143, n144, n145;
  wire n146, n147, n148, n149, n150, n151, n152, n153;
  wire n154, n155, n156, n157, n158, n165, n166, n167;
  wire n168, n169, n170, n171, n172, n173, n174, n175;
  wire n176, n177, n178, n179, n185, n186, n187, n188;
  wire n189, n190, n191, n192, n193, n194, n195, n196;
  wire n200, n204, n205, n206, n207, n208, n209, n210;
  wire n211, n212, n213, n214, n215, n216, n217, n218;
  wire n219, n220, n221, n222, n223, n224, n225, n226;
  wire n227, n228, n233, n234, n235, n236, n237, n238;
  wire n239, n249, n253, n254, n255, n256, n257, n258;
  wire n259, n271, n272, n273, n274, n275, n276, n277;
  wire n278, n279, n280, n281, n282, n283, n284, n285;
  wire n286, n287, n288, n289, n290, n291, n292, n293;
  wire n294, n295, n296, n297, n298, n299, n300, n301;
  wire n302, n303, n311, n312, n313, n314, n315, n316;
  wire n317, n318, n319, n323, n324, n325, n326, n327;
  wire n328, n329, n330, n331, n334, n335, n336, n337;
  wire n341, n342, n343, n344, n345, n346, n347, n348;
  wire n349, n350, n351, n352, n353, n354, n355, n356;
  wire n357, n358, n359, n360, n361, n362, n366, n367;
  wire n368, n369, n370, n371, n372, n373, n380, n381;
  wire n382, n393, n394, n395, n396, n397, n404, n405;
  wire n406, n407, n408, n411, n414, n415, n416, n417;
  wire n421, n422, n423, n431, n432, n437, n444, n445;
  wire n446, n447, n448, n449, n450, n451, n452, n453;
  wire n457, n458, n459, n460, n467, n468, n469, n470;
  wire n471, n472, n473, n474, n475, n476, n477, n478;
  wire n485, n489, n494, n495, n496, n499, n502, n503;
  wire n504, n505, n506, n507, n508, n514, n517, n518;
  wire n519, n520, n521, n522, n523, n524, n525, n526;
  wire n527, n528, n529, n530, n531, n532, n533, n534;
  wire n535, n536, n537, n538, n539, n540, n541, n542;
  wire n543, n544, n545, n546, n547, n548, n549, n550;
  wire n551, n552, n553, n554, n555, n558, n559, n560;
  wire n561, n562, n563, n564, n571, n572, n573, n577;
  wire n578, n581, n584, n585, n586, n587, n588, n589;
  wire n590, n598, n599, n606, n607, n608, n609, n614;
  wire n623, n624, n625, n626, n627, n628, n636, n637;
  wire n638, n643, n644, n645, n646, n647, n648, n653;
  wire n654, n655, n663, n664, n665, n666, n667, n668;
  wire n669, n670, n671, n672, n673, n674, n675, n676;
  wire n677, n678, n679, n680, n681, n682, n683, n684;
  wire n685, n686, n687, n688, n689, n692, n693, n694;
  wire n695, n696, n697, n698, n699, n700, n701, n702;
  wire n703, n704, n705, n706, n707, n708, n711, n712;
  wire n713, n714, n715, n716, n717, n718, n719, n720;
  wire n721, n722, n723, n724, n725, n726, n727, n728;
  wire n735, n736, n739, n744, n752, n753, n757, n758;
  wire n759, n760, n768, n773, n774, n775, n776, n777;
  wire n786, n787, n788, n789, n792, n793, n794, n795;
  wire n796, n805, n806, n807, n808, n809, n813, n814;
  wire n815, n826, n827, n828, n829, n830, n831, n832;
  wire n833, n834, n835, n836, n837, n838, n839, n840;
  wire n841, n842, n843, n844, n845, n846, n847, n848;
  wire n849, n852, n853, n854, n855, n856, n859, n860;
  wire n861, n862, n863, n864, n865, n866, n867, n868;
  wire n869, n870, n871, n872, n873, n874, n875, n876;
  wire n879, n880, n881, n882, n883, n884, n885, n886;
  wire n887, n888, n889, n890, n891, n892, n893, n894;
  wire n895, n896, n897, n898, n899, n900, n901, n902;
  wire n905, n906, n910, n911, n914, n923, n926, n930;
  wire n931, n938, n944, n945, n946, n947, n948, n959;
  wire n960, n961, n967, n968, n969, n970, n975, n976;
  wire n977, n978, n979, n980, n983, n986, n995, n999;
  wire n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014;
  wire n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  wire n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1032;
  wire n1033, n1034, n1035, n1036, n1037, n1038, n1041, n1042;
  wire n1043, n1044, n1045, n1048, n1049, n1050, n1051, n1052;
  wire n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060;
  wire n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068;
  wire n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076;
  wire n1077, n1078, n1081, n1082, n1083, n1084, n1085, n1088;
  wire n1089, n1090, n1091, n1092, n1093, n1096, n1104, n1105;
  wire n1106, n1107, n1108, n1115, n1116, n1117, n1130, n1134;
  wire n1145, n1152, n1162, n1165, n1175, n1176, n1177, n1178;
  wire n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186;
  wire n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194;
  wire n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202;
  wire n1203, n1204, n1205, n1206, n1207, n1210, n1211, n1212;
  wire n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220;
  wire n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228;
  wire n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236;
  wire n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244;
  wire n1245, n1246, n1249, n1250, n1251, n1252, n1253, n1256;
  wire n1257, n1258, n1259, n1260, n1263, n1264, n1265, n1266;
  wire n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274;
  wire n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282;
  wire n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;
  wire n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298;
  wire n1299, n1302, n1303, n1304, n1305, n1306, n1307, n1308;
  wire n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316;
  wire n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324;
  wire n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1334;
  wire n1335, n1336, n1337, n1338, n1341, n1342, n1343, n1344;
  wire n1345, n1346, n1349, n1350, n1351, n1352, n1353, n1354;
  wire n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1364;
  wire n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372;
  wire n1373, n1376, n1377, n1378, n1379, n1380, n1381, n1382;
  wire n1383, n1384, n1385, n1386, n1389, n1390, n1391, n1392;
  wire n1393, n1396, n1397, n1398, n1399, n1400, n1401, n1404;
  wire n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412;
  wire n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420;
  wire n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428;
  wire n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436;
  wire n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444;
  wire n1445, n1448, n1449, n1457, n1458, n1459, n1468, n1476;
  wire n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494;
  wire n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504;
  wire n1505, n1506, n1507, n1508, n1511, n1512, n1513, n1514;
  wire n1515, n1518, n1519, n1520, n1521, n1522, n1523, n1526;
  wire n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534;
  wire n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542;
  wire n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;
  wire n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
  wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
  wire n1569, n1570, n1571, n1572, n1573, n1574, n1577, n1578;
  wire n1579, n1580, n1581, n1584, n1585, n1586, n1587, n1588;
  wire n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598;
  wire n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606;
  wire n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614;
  wire n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622;
  wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
  wire n1633, n1634, n1635, n1636, n1637, n1640, n1641, n1642;
  wire n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650;
  wire n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658;
  wire n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666;
  wire n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674;
  wire n1675, n1676, n1677, n1680, n1681, n1682, n1683, n1684;
  wire n1685, n1688, n1689, n1690, n1691, n1692, n1695, n1696;
  wire n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704;
  wire n1705, n1708, n1709, n1710, n1711, n1712, n1713, n1714;
  wire n1715, n1716, n1717, n1718, n1721, n1722, n1723, n1724;
  wire n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732;
  wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
  wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
  wire n1749, n1750, n1751, n1752, n1753, n1754, n1757, n1758;
  wire n1759, n1760, n1761, n1764, n1765, n1766, n1767, n1768;
  wire n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778;
  wire n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786;
  wire n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794;
  wire n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802;
  wire n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810;
  wire n1811, n1812, n1815, n1816, n1817, n1818, n1819, n1820;
  wire n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
  wire n1831, n1832, n1835, n1836, n1837, n1838, n1839, n1840;
  wire n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848;
  wire n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856;
  wire n1857, n1858, n1859, n1862, n1863, n1864, n1865, n1866;
  wire n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874;
  wire n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882;
  wire n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890;
  wire n1891, n1892, n1893, n1894, n1897, n1898, n1899, n1900;
  wire n1901, n1904, n1905, n1906, n1907, n1908, n1911, n1912;
  wire n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920;
  wire n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928;
  wire n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936;
  wire n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946;
  wire n1949, n1950, n1951, n1952, n1953, n1956, n1957, n1958;
  wire n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966;
  wire n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1976;
  wire n1977, n1978, n1979, n1980, n1983, n1984, n1985, n1986;
  wire n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994;
  wire n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002;
  wire n2003, n2004, n2007, n2008, n2009, n2010, n2011, n2012;
  wire n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020;
  wire n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;
  wire n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036;
  wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
  wire n2045, n2046, n2047, n2051, n2052, n2053, n2054, n2055;
  wire n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063;
  wire n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071;
  wire n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079;
  wire n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087;
  wire n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095;
  wire n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103;
  wire n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111;
  wire n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119;
  wire n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127;
  wire n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135;
  wire n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143;
  wire n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151;
  wire n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159;
  wire n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2170;
  wire n2178, n2181, n2182, n2183, n2190, n2196, n2209, n2210;
  wire n2211, n2212, n2225, n2226, n2227, n2228, n2229, n2239;
  wire n2244, n2250, n2251, n2252, n2253, n2254, n2264, n2265;
  wire n2266, n2267, n2276, n2277, n2278, n2281, n2292, n2293;
  wire n2294, n2295, n2296, n2303, n2311, n2312, n2313, n2317;
  wire n2327, n2328, n2329, n2330, n2333, n2339, n2340, n2341;
  wire n2342, n2354, n2355, n2356, n2357, n2358, n2364, n2365;
  wire n2366, n2367, n2375, n2385, n2386, n2387, n2388, n2395;
  wire n2400, n2414, n2415, n2416, n2417, n2418, n2421, n2422;
  wire n2432, n2433, n2446, n2447, n2448, n2449, n2450, n2454;
  wire n2458, n2464, n2477, n2478, n2479, n2480, n2481, n2482;
  wire n2483, n2484, n2495, n2496, n2497, n2498, n2499, n2500;
  wire n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508;
  wire n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516;
  wire n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524;
  wire n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532;
  wire n2533, n2534, n2535, n2540, n2551, n2552, n2553, n2554;
  wire n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562;
  wire n2563, n2564, n2565, n2566, n2567, n2568, n2571, n2572;
  wire n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580;
  wire n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588;
  wire n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596;
  wire n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604;
  wire n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612;
  wire n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620;
  wire n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628;
  wire n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636;
  wire n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644;
  wire n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652;
  wire n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660;
  wire n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668;
  wire n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676;
  wire n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684;
  wire n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692;
  wire n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700;
  wire n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708;
  wire n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716;
  wire n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724;
  wire n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732;
  wire n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740;
  wire n2741, n2742, n2743, n2744, n2745, n2748, n2749, n2750;
  wire n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758;
  wire n2759, n2760, n2761, n2762, n2763, n2764, n2767, n2768;
  wire n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776;
  wire n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784;
  wire n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792;
  wire n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800;
  wire n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808;
  wire n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816;
  wire n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824;
  wire n2825, n2826, n2829, n2830, n2831, n2832, n2833, n2834;
  wire n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842;
  wire n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850;
  wire n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858;
  wire n2859, n2862, n2863, n2864, n2865, n2866, n2867, n2868;
  wire n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876;
  wire n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884;
  wire n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892;
  wire n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900;
  wire n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908;
  wire n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2918;
  wire n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926;
  wire n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934;
  wire n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942;
  wire n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950;
  wire n2951, n2952, n2955, n2956, n2957, n2958, n2959, n2960;
  wire n2961, n2962, n2965, n2966, n2967, n2968, n2969, n2970;
  wire n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978;
  wire n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986;
  wire n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994;
  wire n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002;
  wire n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010;
  wire n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018;
  wire n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028;
  wire n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036;
  wire n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044;
  wire n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052;
  wire n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060;
  wire n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068;
  wire n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076;
  wire n3077, n3078, n3079, n3080, n3081, n3084, n3085, n3086;
  wire n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094;
  wire n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102;
  wire n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3112;
  wire n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120;
  wire n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128;
  wire n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136;
  wire n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144;
  wire n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152;
  wire n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160;
  wire n3161, n3162, n3163, n3166, n3167, n3168, n3169, n3170;
  wire n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178;
  wire n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186;
  wire n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194;
  wire n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202;
  wire n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210;
  wire n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3229;
  wire n3230, n3231, n3243, n3256, n3257, n3258, n3259, n3269;
  wire n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277;
  wire n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285;
  wire n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293;
  wire n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301;
  wire n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309;
  wire n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317;
  wire n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325;
  wire n3326, n3327, n3328, n3331, n3332, n3333, n3334, n3335;
  wire n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343;
  wire n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351;
  wire n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359;
  wire n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367;
  wire n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375;
  wire n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383;
  wire n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391;
  wire n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399;
  wire n3400, n3401, n3402, n3408, n3409, n3410, n3411, n3412;
  wire n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422;
  wire n3423, n3424, n3425, n3428, n3429, n3430, n3431, n3432;
  wire n3433, n3436, n3437, n3438, n3439, n3440, n3441, n3442;
  wire n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450;
  wire n3453, n3454, n3455, n3456, n3457, n3458, n3461, n3462;
  wire n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470;
  wire n3471, n3472, n3473, n3474, n3477, n3478, n3479, n3480;
  wire n3481, n3482, n3483, n3486, n3487, n3488, n3489, n3490;
  wire n3491, n3494, n3495, n3496, n3497, n3498, n3499, n3500;
  wire n3501, n3502, n3505, n3506, n3507, n3508, n3509, n3510;
  wire n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518;
  wire n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528;
  wire n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536;
  wire n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544;
  wire n3545, n3546, n3547, n3550, n3551, n3552, n3553, n3554;
  wire n3555, n3556, n3557, n3558, n3559, n3562, n3563, n3564;
  wire n3565, n3566, n3567, n3568, n3569, n3570, n3573, n3574;
  wire n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582;
  wire n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590;
  wire n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598;
  wire n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606;
  wire n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614;
  wire n3615, n3616, n3617, n3624, n3625, n3626, n3627, n3628;
  wire n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636;
  wire n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644;
  wire n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652;
  wire n3653, n3657, n3666, n3675, n3678, n3690, n3691, n3692;
  wire n3693, n3699, n3702, n3715, n3716, n3717, n3718, n3719;
  wire n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727;
  wire n3734, n3747, n3748, n3749, n3750, n3751, n3752, n3753;
  wire n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763;
  wire n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771;
  wire n3772, n3775, n3776, n3777, n3778, n3779, n3780, n3781;
  wire n3782, n3783, n3784, n3785, n3786, n3789, n3790, n3791;
  wire n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799;
  wire n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807;
  wire n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815;
  wire n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823;
  wire n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831;
  wire n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839;
  wire n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847;
  wire n3848, n3849, n3850, n3851, n3861, n3862, n3863, n3864;
  wire n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872;
  wire n3873, n3875, n3876, n3883, n3893, n3894, n3895, n3896;
  wire n3897, n3898, n3899, n3902, n3903, n3904, n3905, n3906;
  wire n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914;
  wire n3915, n3916, n3917, n3918, n3921, n3922, n3923, n3924;
  wire n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932;
  wire n3933, n3936, n3937, n3938, n3939, n3940, n3941, n3942;
  wire n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950;
  wire n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958;
  wire n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966;
  wire n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974;
  wire n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982;
  wire n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990;
  wire n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998;
  wire n3999, n4002, n4015, n4016, n4017, n4018, n4019, n4020;
  wire n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028;
  wire n4029, n4030, n4032, n4037, n4048, n4049, n4050, n4051;
  wire n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059;
  wire n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4069;
  wire n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077;
  wire n4078, n4079, n4080, n4081, n4084, n4085, n4086, n4087;
  wire n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095;
  wire n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103;
  wire n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111;
  wire n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119;
  wire n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127;
  wire n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135;
  wire n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143;
  wire n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151;
  wire n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159;
  wire n4160, n4161, n4175, n4176, n4177, n4178, n4179, n4180;
  wire n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188;
  wire n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198;
  wire n4199, n4200, n4201, n4202, n4203, n4206, n4207, n4208;
  wire n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216;
  wire n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224;
  wire n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232;
  wire n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240;
  wire n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248;
  wire n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256;
  wire n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264;
  wire n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272;
  wire n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4281;
  wire n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298;
  wire n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308;
  wire n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316;
  wire n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324;
  wire n4325, n4328, n4329, n4330, n4331, n4332, n4333, n4334;
  wire n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342;
  wire n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352;
  wire n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4362;
  wire n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370;
  wire n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378;
  wire n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386;
  wire n4387, n4388, n4390, n4391, n4392, n4404, n4405, n4406;
  wire n4407, n4408, n4409, n4410, n4411, n4414, n4415, n4416;
  wire n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424;
  wire n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432;
  wire n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440;
  wire n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448;
  wire n4449, n4452, n4453, n4454, n4455, n4456, n4457, n4458;
  wire n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466;
  wire n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474;
  wire n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482;
  wire n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490;
  wire n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498;
  wire n4499, n4500, n4501, n4502, n4503, n4505, n4513, n4523;
  wire n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531;
  wire n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4541;
  wire n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549;
  wire n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557;
  wire n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565;
  wire n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573;
  wire n4574, n4575, n4578, n4579, n4580, n4581, n4582, n4583;
  wire n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591;
  wire n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599;
  wire n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607;
  wire n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615;
  wire n4616, n4618, n4619, n4620, n4621, n4622, n4623, n4624;
  wire n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632;
  wire n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4642;
  wire n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650;
  wire n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658;
  wire n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666;
  wire n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674;
  wire n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682;
  wire n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690;
  wire n4691, n4702, n4703, n4704, n4705, n4706, n4707, n4708;
  wire n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4717;
  wire n4726, n4737, n4738, n4739, n4740, n4741, n4742, n4743;
  wire n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751;
  wire n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759;
  wire n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767;
  wire n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775;
  wire n4776, n4777, n4778, n4779, n4782, n4783, n4784, n4785;
  wire n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793;
  wire n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801;
  wire n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809;
  wire n4810, n4811, n4812, n4813, n4814, n4815, n4817, n4829;
  wire n4830, n4831, n4832, n4833, n4834, n4837, n4838, n4839;
  wire n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847;
  wire n4848, n4849, n4850, n4851, n4852, n4853, n4856, n4857;
  wire n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865;
  wire n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873;
  wire n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881;
  wire n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889;
  wire n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897;
  wire n4898, n4900, n4911, n4912, n4913, n4914, n4915, n4916;
  wire n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924;
  wire n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932;
  wire n4933, n4936, n4937, n4938, n4939, n4940, n4941, n4942;
  wire n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950;
  wire n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958;
  wire n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966;
  wire n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974;
  wire n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982;
  wire n4983, n4984, n4985, n4987, n4993, n4994, n4995, n4996;
  wire n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004;
  wire n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012;
  wire n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020;
  wire n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028;
  wire n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036;
  wire n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044;
  wire n5045, n5046, n5047, n5048, n5049, n5051, n5055, n5063;
  wire n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071;
  wire n5072, n5073, n5074, n5077, n5078, n5079, n5080, n5081;
  wire n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089;
  wire n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097;
  wire n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105;
  wire n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113;
  wire n5114, n5115, n5116, n5117, n5118, n5119, n5121, n5125;
  wire n5138, n5139, n5140, n5141, n5142, n5145, n5146, n5147;
  wire n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155;
  wire n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163;
  wire n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171;
  wire n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179;
  wire n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187;
  wire n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209;
  wire n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217;
  wire n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225;
  wire n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233;
  wire n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241;
  wire n5242, n5244, n5247, n5258, n5259, n5260, n5261, n5262;
  wire n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270;
  wire n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278;
  wire n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286;
  wire n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5303;
  wire n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311;
  wire n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319;
  wire n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327;
  wire n5328, n5329, n5330, n5331, n5332, n5344, n5345, n5346;
  wire n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354;
  wire n5356, n5367, n5368, n5369, n5370, n5371, n5372, n5373;
  wire n5374, n5375, n5376, n5377, n5389, n5390, n5391, n5392;
  wire n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5412;
  wire n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420;
  wire n5421, n5422, n5427, n5428, n5429, n5430, n5431, n5432;
  wire n5433, n5434, n5435, n5436, n5437, n5439, n5440, n5441;
  wire n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449;
  wire n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458;
  wire n5459, n5461, n5462, n5463, n5464, n_5, n_6, n_8;
  wire n_10, n_12, n_14, n_16, n_18, n_20, n_22, n_24;
  wire n_26, n_28, n_30, n_32, n_34, n_36, n_38, n_40;
  wire n_42, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_614, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_638, n_639, n_640, n_641, n_642;
  wire n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_681, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718;
  wire n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
  wire n_735, n_736, n_737, n_738, n_739, n_740, n_757, n_758;
  wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
  wire n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790;
  wire n_791, n_792, n_793, n_794, n_795, n_804, n_805, n_806;
  wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814;
  wire n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822;
  wire n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830;
  wire n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_860, n_861;
  wire n_862, n_863, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_912, n_913, n_914, n_915, n_916, n_917;
  wire n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925;
  wire n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933;
  wire n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941;
  wire n_942, n_943, n_944, n_945, n_946, n_955, n_956, n_957;
  wire n_958, n_959, n_960, n_961, n_966, n_967, n_968, n_969;
  wire n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977;
  wire n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
  wire n_986, n_987, n_988, n_993, n_994, n_995, n_996, n_997;
  wire n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005;
  wire n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013;
  wire n_1014, n_1015, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049;
  wire n_1053, n_1054, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
  wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1104;
  wire n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112;
  wire n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120;
  wire n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128;
  wire n_1129, n_1130, n_1131, n_1132, n_1133, n_1139, n_1140, n_1141;
  wire n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149;
  wire n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157;
  wire n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165;
  wire n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
  wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189;
  wire n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197;
  wire n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213;
  wire n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
  wire n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261;
  wire n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293;
  wire n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317;
  wire n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325;
  wire n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1372, n_1373, n_1374, n_1375, n_1376;
  wire n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408;
  wire n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416;
  wire n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424;
  wire n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432;
  wire n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440;
  wire n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465;
  wire n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473;
  wire n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481;
  wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505;
  wire n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1516;
  wire n_1517, n_1518, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1534, n_1535, n_1537;
  wire n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545;
  wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553;
  wire n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561;
  wire n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569;
  wire n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577;
  wire n_1578, n_1579, n_1580, n_1584, n_1585, n_1587, n_1588, n_1589;
  wire n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597;
  wire n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605;
  wire n_1606, n_1607, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633;
  wire n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641;
  wire n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1651, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1697;
  wire n_1698, n_1699, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1751, n_1752;
  wire n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761;
  wire n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769;
  wire n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777;
  wire n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785;
  wire n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793;
  wire n_1794, n_1795, n_1796, n_1797, n_1802, n_1803, n_1804, n_1805;
  wire n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813;
  wire n_1814, n_1815, n_1816, n_1817, n_1822, n_1823, n_1824, n_1825;
  wire n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833;
  wire n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841;
  wire n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849;
  wire n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1861;
  wire n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869;
  wire n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877;
  wire n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885;
  wire n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893;
  wire n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901;
  wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909;
  wire n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917;
  wire n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925;
  wire n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933;
  wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957;
  wire n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965;
  wire n_1966, n_1967, n_1968, n_1969, n_1970, n_1974, n_1975, n_1977;
  wire n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985;
  wire n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993;
  wire n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001;
  wire n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009;
  wire n_2010, n_2011, n_2012, n_2013, n_2020, n_2025, n_2026, n_2027;
  wire n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2039;
  wire n_2040, n_2041, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051;
  wire n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2063;
  wire n_2064, n_2065, n_2066, n_2071, n_2072, n_2073, n_2074, n_2075;
  wire n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083;
  wire n_2088, n_2089, n_2090, n_2091, n_2092, n_2097, n_2098, n_2099;
  wire n_2100, n_2101, n_2102, n_2103, n_2108, n_2109, n_2110, n_2111;
  wire n_2112, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123;
  wire n_2124, n_2125, n_2126, n_2131, n_2132, n_2133, n_2134, n_2135;
  wire n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143;
  wire n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151;
  wire n_2152, n_2153, n_2154, n_2159, n_2160, n_2161, n_2166, n_2167;
  wire n_2168, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179;
  wire n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203;
  wire n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211;
  wire n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219;
  wire n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227;
  wire n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235;
  wire n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243;
  wire n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251;
  wire n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259;
  wire n_2260, n_2261, n_2262, n_2266, n_2267, n_2268, n_2269, n_2270;
  wire n_2271, n_2272, n_2274, n_2275, n_2276, n_2277, n_2282, n_2283;
  wire n_2284, n_2285, n_2286, n_2291, n_2292, n_2293, n_2294, n_2295;
  wire n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303;
  wire n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311;
  wire n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319;
  wire n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327;
  wire n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335;
  wire n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343;
  wire n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351;
  wire n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359;
  wire n_2360, n_2361, n_2362, n_2363, n_2364, n_2368, n_2369, n_2370;
  wire n_2371, n_2372, n_2373, n_2374, n_2376, n_2377, n_2378, n_2379;
  wire n_2384, n_2385, n_2386, n_2387, n_2388, n_2393, n_2394, n_2395;
  wire n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403;
  wire n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411;
  wire n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419;
  wire n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435;
  wire n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443;
  wire n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451;
  wire n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459;
  wire n_2460, n_2461, n_2462, n_2464, n_2465, n_2466, n_2468, n_2469;
  wire n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477;
  wire n_2478, n_2479, n_2480, n_2485, n_2486, n_2487, n_2488, n_2489;
  wire n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517;
  wire n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525;
  wire n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533;
  wire n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541;
  wire n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549;
  wire n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557;
  wire n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565;
  wire n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573;
  wire n_2574, n_2579, n_2580, n_2581, n_2582, n_2583, n_2588, n_2589;
  wire n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597;
  wire n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605;
  wire n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613;
  wire n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621;
  wire n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629;
  wire n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637;
  wire n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645;
  wire n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653;
  wire n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661;
  wire n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673;
  wire n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681;
  wire n_2682, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693;
  wire n_2694, n_2695, n_2696, n_2697, n_2702, n_2703, n_2704, n_2705;
  wire n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713;
  wire n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725;
  wire n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733;
  wire n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741;
  wire n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2752, n_2753;
  wire n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761;
  wire n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769;
  wire n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2781;
  wire n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789;
  wire n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797;
  wire n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805;
  wire n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813;
  wire n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821;
  wire n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829;
  wire n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837;
  wire n_2838, n_2839, n_2840, n_2845, n_2846, n_2847, n_2848, n_2849;
  wire n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857;
  wire n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865;
  wire n_2866, n_2867, n_2868, n_2873, n_2874, n_2875, n_2876, n_2877;
  wire n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885;
  wire n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893;
  wire n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901;
  wire n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909;
  wire n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917;
  wire n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925;
  wire n_2926, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937;
  wire n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945;
  wire n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953;
  wire n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961;
  wire n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969;
  wire n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977;
  wire n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985;
  wire n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993;
  wire n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001;
  wire n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009;
  wire n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017;
  wire n_3018, n_3019, n_3020, n_3021, n_3022, n_3027, n_3028, n_3029;
  wire n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037;
  wire n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045;
  wire n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053;
  wire n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061;
  wire n_3062, n_3063, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073;
  wire n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3085;
  wire n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093;
  wire n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101;
  wire n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109;
  wire n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117;
  wire n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125;
  wire n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133;
  wire n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3144, n_3145;
  wire n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153;
  wire n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161;
  wire n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169;
  wire n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177;
  wire n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185;
  wire n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193;
  wire n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201;
  wire n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209;
  wire n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217;
  wire n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225;
  wire n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233;
  wire n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241;
  wire n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3253;
  wire n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261;
  wire n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269;
  wire n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277;
  wire n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285;
  wire n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293;
  wire n_3294, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305;
  wire n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313;
  wire n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321;
  wire n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329;
  wire n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337;
  wire n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345;
  wire n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353;
  wire n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361;
  wire n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369;
  wire n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377;
  wire n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385;
  wire n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393;
  wire n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401;
  wire n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409;
  wire n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417;
  wire n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425;
  wire n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433;
  wire n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441;
  wire n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449;
  wire n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457;
  wire n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465;
  wire n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473;
  wire n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481;
  wire n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489;
  wire n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497;
  wire n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505;
  wire n_3506, n_3507, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537;
  wire n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545;
  wire n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553;
  wire n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561;
  wire n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569;
  wire n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577;
  wire n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585;
  wire n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593;
  wire n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609;
  wire n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617;
  wire n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625;
  wire n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633;
  wire n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641;
  wire n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649;
  wire n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657;
  wire n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665;
  wire n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673;
  wire n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681;
  wire n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689;
  wire n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697;
  wire n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705;
  wire n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713;
  wire n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721;
  wire n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729;
  wire n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737;
  wire n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745;
  wire n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753;
  wire n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761;
  wire n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769;
  wire n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777;
  wire n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785;
  wire n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793;
  wire n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801;
  wire n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809;
  wire n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817;
  wire n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825;
  wire n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833;
  wire n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841;
  wire n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849;
  wire n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857;
  wire n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865;
  wire n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873;
  wire n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881;
  wire n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889;
  wire n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897;
  wire n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905;
  wire n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913;
  wire n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921;
  wire n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929;
  wire n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937;
  wire n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945;
  wire n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953;
  wire n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961;
  wire n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969;
  wire n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977;
  wire n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985;
  wire n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993;
  wire n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001;
  wire n_4002, n_4003, n_4004, n_4005, n_4006, n_4007;
  and g1 (n50, \a[21] , \a[22] );
  not g2 (n_5, \a[1] );
  not g3 (n_6, \a[2] );
  and g4 (n51, n_5, n_6);
  not g5 (n_8, \a[0] );
  and g6 (n52, n_8, n51);
  not g7 (n_10, \a[3] );
  and g8 (n53, n_10, n52);
  not g9 (n_12, \a[4] );
  and g10 (n54, n_12, n53);
  not g11 (n_14, \a[5] );
  and g12 (n55, n_14, n54);
  not g13 (n_16, \a[6] );
  and g14 (n56, n_16, n55);
  not g15 (n_18, \a[7] );
  and g16 (n57, n_18, n56);
  not g17 (n_20, \a[8] );
  and g18 (n58, n_20, n57);
  not g19 (n_22, \a[9] );
  and g20 (n59, n_22, n58);
  not g21 (n_24, \a[10] );
  and g22 (n60, n_24, n59);
  not g23 (n_26, \a[11] );
  and g24 (n61, n_26, n60);
  not g25 (n_28, \a[12] );
  and g26 (n62, n_28, n61);
  not g27 (n_30, \a[13] );
  and g28 (n63, n_30, n62);
  not g29 (n_32, \a[14] );
  and g30 (n64, n_32, n63);
  not g31 (n_34, \a[15] );
  and g32 (n65, n_34, n64);
  not g33 (n_36, \a[16] );
  and g34 (n66, n_36, n65);
  not g35 (n_38, \a[17] );
  and g36 (n67, n_38, n66);
  not g37 (n_40, \a[18] );
  and g38 (n68, n_40, n67);
  not g39 (n_42, \a[19] );
  and g40 (n69, n_42, n68);
  not g41 (n_44, \a[20] );
  and g42 (n70, n_44, n69);
  not g43 (n_45, \a[21] );
  and g44 (n71, n_45, n70);
  not g45 (n_46, n70);
  and g46 (n72, \a[21] , n_46);
  not g47 (n_47, n71);
  not g48 (n_48, n72);
  and g49 (n73, n_47, n_48);
  not g50 (n_49, \a[22] );
  and g51 (n74, n_49, n73);
  not g52 (n_50, n50);
  not g53 (n_51, n74);
  and g54 (n75, n_50, n_51);
  and g55 (n76, \a[20] , \a[22] );
  not g56 (n_52, n69);
  and g57 (n77, \a[20] , n_52);
  not g58 (n_53, n77);
  and g59 (n78, n_46, n_53);
  and g60 (n79, n_49, n78);
  not g61 (n_54, n76);
  not g62 (n_55, n79);
  and g63 (n80, n_54, n_55);
  and g64 (n81, n75, n80);
  and g65 (n82, \a[15] , \a[22] );
  not g66 (n_56, n65);
  and g67 (n83, n_49, n_56);
  not g68 (n_57, n64);
  and g69 (n84, \a[15] , n_57);
  not g70 (n_58, n84);
  and g71 (n85, n83, n_58);
  not g72 (n_59, n82);
  not g73 (n_60, n85);
  and g74 (n86, n_59, n_60);
  and g75 (n87, n81, n86);
  not g76 (n_61, n68);
  and g77 (n88, n_49, n_61);
  not g78 (n_62, n88);
  and g79 (n89, \a[19] , n_62);
  and g80 (n90, n_42, n88);
  not g81 (n_63, n89);
  not g82 (n_64, n90);
  and g83 (n91, n_63, n_64);
  and g84 (n92, \a[18] , \a[22] );
  not g85 (n_65, n67);
  and g86 (n93, \a[18] , n_65);
  not g87 (n_66, n93);
  and g88 (n94, n88, n_66);
  not g89 (n_67, n92);
  not g90 (n_68, n94);
  and g91 (n95, n_67, n_68);
  not g92 (n_69, n91);
  not g93 (n_70, n95);
  and g94 (n96, n_69, n_70);
  not g95 (n_71, n66);
  and g96 (n97, n_49, n_71);
  not g97 (n_72, n97);
  and g98 (n98, \a[17] , n_72);
  and g99 (n99, n_38, n97);
  not g100 (n_73, n98);
  not g101 (n_74, n99);
  and g102 (n100, n_73, n_74);
  not g103 (n_75, n83);
  and g104 (n101, \a[16] , n_75);
  and g105 (n102, n_36, n83);
  not g106 (n_76, n101);
  not g107 (n_77, n102);
  and g108 (n103, n_76, n_77);
  not g109 (n_78, n100);
  and g110 (n104, n_78, n103);
  and g111 (n105, n96, n104);
  and g112 (n106, n87, n105);
  and g113 (n107, n100, n103);
  and g114 (n108, n96, n107);
  not g115 (n_79, n80);
  and g116 (n109, n75, n_79);
  and g117 (n110, n86, n109);
  and g118 (n111, n108, n110);
  and g119 (n112, n_69, n95);
  and g120 (n113, n107, n112);
  and g121 (n114, n110, n113);
  not g122 (n_80, n86);
  and g123 (n115, n_80, n109);
  and g124 (n116, n91, n_70);
  and g125 (n117, n107, n116);
  and g126 (n118, n115, n117);
  not g127 (n_81, n75);
  and g128 (n119, n_81, n80);
  and g129 (n120, n_80, n119);
  not g130 (n_82, n103);
  and g131 (n121, n100, n_82);
  and g132 (n122, n112, n121);
  and g133 (n123, n120, n122);
  and g134 (n124, n_81, n_79);
  and g135 (n125, n_80, n124);
  and g136 (n126, n104, n112);
  and g137 (n127, n125, n126);
  and g138 (n128, n86, n124);
  and g139 (n129, n105, n128);
  and g140 (n130, n81, n_80);
  and g141 (n131, n104, n116);
  and g142 (n132, n130, n131);
  and g143 (n133, n105, n120);
  and g144 (n134, n122, n125);
  and g145 (n135, n_78, n_82);
  and g146 (n136, n116, n135);
  and g147 (n137, n125, n136);
  and g148 (n138, n128, n136);
  and g149 (n139, n122, n128);
  and g150 (n140, n128, n131);
  not g151 (n_83, n139);
  not g152 (n_84, n140);
  and g153 (n141, n_83, n_84);
  and g154 (n142, n105, n110);
  and g155 (n143, n96, n121);
  and g156 (n144, n128, n143);
  not g157 (n_85, n142);
  not g158 (n_86, n144);
  and g159 (n145, n_85, n_86);
  and g160 (n146, n105, n115);
  and g161 (n147, n116, n121);
  and g162 (n148, n110, n147);
  not g163 (n_87, n146);
  not g164 (n_88, n148);
  and g165 (n149, n_87, n_88);
  and g166 (n150, n126, n128);
  and g167 (n151, n112, n135);
  and g168 (n152, n128, n151);
  not g169 (n_89, n150);
  not g170 (n_90, n152);
  and g171 (n153, n_89, n_90);
  and g172 (n154, n130, n136);
  and g173 (n155, n105, n125);
  not g174 (n_91, n154);
  not g175 (n_92, n155);
  and g176 (n156, n_91, n_92);
  and g177 (n157, n153, n156);
  and g178 (n158, n149, n157);
  not g181 (n_93, n138);
  not g183 (n_94, n137);
  not g185 (n_95, n134);
  not g187 (n_96, n133);
  not g189 (n_97, n132);
  and g191 (n166, n110, n143);
  and g192 (n167, n120, n151);
  and g193 (n168, n87, n151);
  and g194 (n169, n115, n122);
  and g195 (n170, n91, n95);
  and g196 (n171, n107, n170);
  and g197 (n172, n115, n171);
  and g198 (n173, n86, n119);
  and g199 (n174, n151, n173);
  and g200 (n175, n108, n125);
  and g201 (n176, n125, n143);
  and g202 (n177, n117, n173);
  and g203 (n178, n108, n128);
  not g204 (n_98, n177);
  not g205 (n_99, n178);
  and g206 (n179, n_98, n_99);
  not g207 (n_100, n176);
  not g209 (n_101, n175);
  not g211 (n_102, n174);
  not g213 (n_103, n172);
  not g215 (n_104, n169);
  not g217 (n_105, n168);
  and g219 (n186, n108, n120);
  and g220 (n187, n135, n170);
  and g221 (n188, n128, n187);
  not g222 (n_106, n186);
  not g223 (n_107, n188);
  and g224 (n189, n_106, n_107);
  and g225 (n190, n110, n151);
  and g226 (n191, n117, n120);
  and g227 (n192, n120, n126);
  and g228 (n193, n121, n170);
  and g229 (n194, n125, n193);
  and g230 (n195, n96, n135);
  and g231 (n196, n128, n195);
  not g232 (n_108, n194);
  not g233 (n_109, n196);
  not g235 (n_110, n192);
  not g237 (n_111, n191);
  not g239 (n_112, n190);
  not g243 (n_113, n167);
  not g245 (n_114, n166);
  and g247 (n205, n104, n170);
  and g248 (n206, n115, n205);
  and g249 (n207, n120, n131);
  and g250 (n208, n128, n147);
  not g251 (n_115, n207);
  not g252 (n_116, n208);
  and g253 (n209, n_115, n_116);
  not g254 (n_117, n206);
  and g255 (n210, n_117, n209);
  and g256 (n211, n130, n147);
  and g257 (n212, n115, n195);
  and g258 (n213, n171, n173);
  and g259 (n214, n125, n171);
  and g260 (n215, n117, n130);
  and g261 (n216, n110, n126);
  and g262 (n217, n120, n147);
  and g263 (n218, n108, n173);
  and g264 (n219, n125, n187);
  and g265 (n220, n125, n131);
  and g266 (n221, n125, n147);
  and g267 (n222, n128, n193);
  and g268 (n223, n122, n130);
  and g269 (n224, n115, n126);
  and g270 (n225, n120, n143);
  and g271 (n226, n105, n173);
  and g272 (n227, n125, n151);
  and g273 (n228, n113, n125);
  not g274 (n_118, n227);
  not g275 (n_119, n228);
  not g277 (n_120, n226);
  not g279 (n_121, n225);
  not g281 (n_122, n224);
  not g283 (n_123, n223);
  and g285 (n234, n115, n187);
  and g286 (n235, n105, n130);
  not g287 (n_124, n234);
  not g288 (n_125, n235);
  and g289 (n236, n_124, n_125);
  and g290 (n237, n130, n187);
  and g291 (n238, n130, n205);
  not g292 (n_126, n237);
  not g293 (n_127, n238);
  and g294 (n239, n_126, n_127);
  not g297 (n_128, n222);
  not g299 (n_129, n221);
  not g301 (n_130, n220);
  not g303 (n_131, n219);
  not g305 (n_132, n218);
  not g307 (n_133, n217);
  not g309 (n_134, n216);
  not g311 (n_135, n215);
  not g313 (n_136, n214);
  not g315 (n_137, n213);
  not g317 (n_138, n212);
  not g319 (n_139, n211);
  and g321 (n254, n173, n193);
  and g322 (n255, n120, n195);
  not g323 (n_140, n254);
  not g324 (n_141, n255);
  and g325 (n256, n_140, n_141);
  and g326 (n257, n113, n173);
  and g327 (n258, n87, n193);
  not g328 (n_142, n257);
  not g329 (n_143, n258);
  and g330 (n259, n_142, n_143);
  not g336 (n_144, n129);
  not g338 (n_145, n127);
  not g340 (n_146, n123);
  not g342 (n_147, n118);
  not g344 (n_148, n114);
  not g346 (n_149, n111);
  not g348 (n_150, n106);
  not g350 (n_151, n54);
  and g351 (n272, n_49, n_151);
  not g352 (n_152, n272);
  and g353 (n273, \a[5] , n_152);
  and g354 (n274, n_14, n272);
  not g355 (n_153, n273);
  not g356 (n_154, n274);
  and g357 (n275, n_153, n_154);
  and g358 (n276, \a[4] , \a[22] );
  not g359 (n_155, n53);
  and g360 (n277, \a[4] , n_155);
  not g361 (n_156, n277);
  and g362 (n278, n272, n_156);
  not g363 (n_157, n276);
  not g364 (n_158, n278);
  and g365 (n279, n_157, n_158);
  not g366 (n_159, n279);
  and g367 (n280, n275, n_159);
  not g368 (n_160, n275);
  and g369 (n281, n_160, n279);
  not g370 (n_161, n280);
  not g371 (n_162, n281);
  and g372 (n282, n_161, n_162);
  not g373 (n_163, n52);
  and g374 (n283, n_49, n_163);
  not g375 (n_164, n283);
  and g376 (n284, \a[3] , n_164);
  and g377 (n285, n_10, n283);
  not g378 (n_165, n284);
  not g379 (n_166, n285);
  and g380 (n286, n_165, n_166);
  and g381 (n287, \a[2] , \a[22] );
  and g382 (n288, n_8, n_5);
  not g383 (n_167, n288);
  and g384 (n289, \a[2] , n_167);
  not g385 (n_168, n289);
  and g386 (n290, n283, n_168);
  not g387 (n_169, n287);
  not g388 (n_170, n290);
  and g389 (n291, n_169, n_170);
  not g390 (n_171, n291);
  and g391 (n292, n286, n_171);
  not g392 (n_172, n286);
  and g393 (n293, n_172, n291);
  not g394 (n_173, n292);
  not g395 (n_174, n293);
  and g396 (n294, n_173, n_174);
  not g397 (n_175, n294);
  and g398 (n295, n282, n_175);
  and g399 (n296, n130, n151);
  and g400 (n297, n108, n115);
  and g401 (n298, n113, n115);
  and g402 (n299, n122, n173);
  and g403 (n300, n120, n205);
  not g404 (n_176, n300);
  and g405 (n301, n_139, n_176);
  and g406 (n302, n115, n131);
  not g407 (n_177, n302);
  and g408 (n303, n_149, n_177);
  not g412 (n_178, n299);
  not g415 (n_179, n298);
  not g417 (n_180, n297);
  not g419 (n_181, n296);
  and g421 (n312, n173, n195);
  and g422 (n313, n120, n136);
  not g423 (n_182, n313);
  and g424 (n314, n_129, n_182);
  and g425 (n315, n110, n187);
  not g426 (n_183, n315);
  and g427 (n316, n_148, n_183);
  and g428 (n317, n125, n205);
  not g429 (n_184, n317);
  and g430 (n318, n_144, n_184);
  and g431 (n319, n_115, n318);
  not g434 (n_185, n312);
  and g437 (n324, n87, n171);
  not g438 (n_186, n324);
  and g439 (n325, n_146, n_186);
  and g440 (n326, n87, n147);
  and g441 (n327, n136, n173);
  and g442 (n328, n128, n205);
  and g443 (n329, n147, n173);
  not g444 (n_187, n328);
  not g445 (n_188, n329);
  and g446 (n330, n_187, n_188);
  and g447 (n331, n_141, n330);
  not g448 (n_189, n327);
  not g451 (n_190, n326);
  and g453 (n335, n110, n193);
  and g454 (n336, n113, n120);
  and g455 (n337, n113, n128);
  not g456 (n_191, n337);
  not g459 (n_192, n336);
  not g461 (n_193, n335);
  and g463 (n342, n108, n130);
  and g464 (n343, n173, n187);
  not g465 (n_194, n342);
  not g466 (n_195, n343);
  and g467 (n344, n_194, n_195);
  and g468 (n345, n130, n171);
  not g469 (n_196, n345);
  and g470 (n346, n_89, n_196);
  and g471 (n347, n110, n195);
  and g472 (n348, n131, n173);
  not g473 (n_197, n347);
  not g474 (n_198, n348);
  and g475 (n349, n_197, n_198);
  and g476 (n350, n126, n173);
  and g477 (n351, n87, n113);
  and g478 (n352, n_110, n_120);
  not g479 (n_199, n351);
  and g480 (n353, n_199, n352);
  and g481 (n354, n_133, n353);
  and g482 (n355, n_134, n354);
  and g483 (n356, n110, n171);
  and g484 (n357, n110, n136);
  and g485 (n358, n110, n205);
  and g486 (n359, n110, n117);
  and g487 (n360, n120, n187);
  and g488 (n361, n115, n147);
  not g489 (n_200, n360);
  not g490 (n_201, n361);
  and g491 (n362, n_200, n_201);
  not g492 (n_202, n359);
  not g494 (n_203, n358);
  not g496 (n_204, n357);
  not g498 (n_205, n356);
  and g500 (n367, n87, n195);
  and g501 (n368, n87, n126);
  not g502 (n_206, n368);
  and g503 (n369, n_145, n_206);
  and g504 (n370, n173, n205);
  not g505 (n_207, n370);
  and g506 (n371, n369, n_207);
  not g507 (n_208, n367);
  and g508 (n372, n_208, n371);
  and g509 (n373, n_150, n_135);
  and g517 (n381, n156, n380);
  not g518 (n_209, n350);
  and g519 (n382, n_209, n381);
  and g531 (n394, n125, n195);
  and g532 (n395, n_110, n_209);
  and g533 (n396, n_102, n_191);
  and g534 (n397, n_115, n_189);
  and g542 (n405, n117, n125);
  and g543 (n406, n_94, n_142);
  and g544 (n407, n_192, n406);
  and g545 (n408, n117, n128);
  not g546 (n_210, n408);
  not g551 (n_211, n405);
  and g554 (n415, n128, n171);
  not g555 (n_212, n415);
  and g556 (n416, n_141, n_212);
  and g557 (n417, n143, n173);
  not g562 (n_213, n417);
  and g563 (n422, n_213, n421);
  and g564 (n423, n_132, n422);
  and g573 (n432, n_92, n_108);
  not g585 (n_214, n394);
  and g587 (n445, n87, n122);
  and g588 (n446, n120, n171);
  and g589 (n447, n115, n151);
  not g590 (n_215, n447);
  and g591 (n448, n_112, n_215);
  and g592 (n449, n115, n143);
  not g593 (n_216, n449);
  and g594 (n450, n_180, n_216);
  and g595 (n451, n_114, n450);
  and g596 (n452, n448, n451);
  and g597 (n453, n_87, n452);
  and g602 (n458, n120, n193);
  not g603 (n_217, n458);
  and g604 (n459, n_176, n_217);
  and g605 (n460, n_200, n_207);
  not g611 (n_218, n446);
  and g614 (n468, n113, n130);
  and g615 (n469, n126, n130);
  and g616 (n470, n87, n108);
  and g617 (n471, n130, n195);
  and g618 (n472, n87, n143);
  and g619 (n473, n_98, n_188);
  and g620 (n474, n_125, n_205);
  and g621 (n475, n_111, n_133);
  and g622 (n476, n_103, n475);
  and g623 (n477, n130, n143);
  not g624 (n_219, n477);
  and g625 (n478, n_194, n_219);
  not g631 (n_220, n472);
  not g633 (n_221, n471);
  not g635 (n_222, n470);
  not g639 (n_223, n469);
  not g641 (n_224, n468);
  not g645 (n_225, n445);
  and g648 (n495, n115, n193);
  and g649 (n496, n_147, n_193);
  not g650 (n_226, n495);
  and g657 (n503, n110, n122);
  and g658 (n504, n115, n136);
  not g659 (n_227, n504);
  and g660 (n505, n_134, n_227);
  and g661 (n506, n110, n131);
  and g662 (n507, n_204, n_201);
  not g663 (n_228, n506);
  and g664 (n508, n_228, n507);
  not g670 (n_229, n503);
  and g675 (n518, n502, n517);
  and g676 (n519, n_88, n518);
  not g677 (n_230, n494);
  not g678 (n_231, n519);
  and g679 (n520, n_230, n_231);
  and g680 (n521, \a[14] , \a[22] );
  not g681 (n_232, n63);
  and g682 (n522, \a[14] , n_232);
  not g683 (n_233, n522);
  and g684 (n523, n_57, n_233);
  and g685 (n524, n_49, n523);
  not g686 (n_234, n521);
  not g687 (n_235, n524);
  and g688 (n525, n_234, n_235);
  not g689 (n_236, n62);
  and g690 (n526, n_49, n_236);
  not g691 (n_237, n526);
  and g692 (n527, \a[13] , n_237);
  and g693 (n528, n_30, n526);
  not g694 (n_238, n527);
  not g695 (n_239, n528);
  and g696 (n529, n_238, n_239);
  not g697 (n_240, n525);
  and g698 (n530, n_240, n529);
  not g699 (n_241, n529);
  and g700 (n531, n525, n_241);
  not g701 (n_242, n530);
  not g702 (n_243, n531);
  and g703 (n532, n_242, n_243);
  and g704 (n533, n520, n532);
  not g705 (n_244, n520);
  not g706 (n_245, n532);
  and g707 (n534, n_244, n_245);
  not g708 (n_246, n533);
  not g709 (n_247, n534);
  and g710 (n535, n_246, n_247);
  not g711 (n_248, n444);
  and g712 (n536, n_248, n535);
  and g713 (n537, n494, n_231);
  and g714 (n538, n_230, n519);
  not g715 (n_249, n537);
  not g716 (n_250, n538);
  and g717 (n539, n_249, n_250);
  and g718 (n540, n494, n519);
  not g719 (n_251, n540);
  and g720 (n541, n444, n_251);
  not g721 (n_252, n541);
  and g722 (n542, n539, n_252);
  and g723 (n543, n_240, n542);
  and g724 (n544, n_248, n_244);
  not g725 (n_253, n539);
  not g726 (n_254, n544);
  and g727 (n545, n_253, n_254);
  and g728 (n546, n525, n_254);
  not g729 (n_255, n545);
  not g730 (n_256, n546);
  and g731 (n547, n_255, n_256);
  not g732 (n_257, n543);
  and g733 (n548, n_257, n547);
  and g734 (n549, n_248, n_241);
  not g735 (n_258, n549);
  and g736 (n550, n548, n_258);
  not g737 (n_259, n548);
  and g738 (n551, n_259, n549);
  and g739 (n552, n87, n136);
  and g740 (n553, n87, n205);
  and g741 (n554, n87, n131);
  not g742 (n_260, n554);
  and g743 (n555, n_127, n_260);
  and g747 (n559, n_121, n_213);
  and g748 (n560, n_181, n559);
  and g749 (n561, n_124, n_221);
  and g750 (n562, n_126, n561);
  and g751 (n563, n_118, n_214);
  and g752 (n564, n_145, n563);
  not g759 (n_261, n553);
  and g761 (n572, n_113, n_130);
  and g762 (n573, n_111, n572);
  and g767 (n578, n_147, n_109);
  and g774 (n585, n_179, n_197);
  and g775 (n586, n_205, n585);
  and g776 (n587, n165, n_119);
  and g777 (n588, n_202, n587);
  and g778 (n589, n87, n187);
  not g779 (n_262, n589);
  and g780 (n590, n_106, n_262);
  not g788 (n_263, n552);
  and g790 (n599, n87, n117);
  and g798 (n607, n_128, n_191);
  and g799 (n608, n_148, n607);
  and g800 (n609, n_184, n_211);
  and g815 (n624, n_214, n623);
  and g816 (n625, n_199, n624);
  and g817 (n626, n_116, n_136);
  and g818 (n627, n_94, n626);
  and g819 (n628, n_104, n627);
  not g826 (n_264, n599);
  and g829 (n637, n_185, n_212);
  and g830 (n638, n_100, n_229);
  and g836 (n644, n_137, n_220);
  and g837 (n645, n_93, n_119);
  and g838 (n646, n_219, n645);
  and g839 (n647, n_145, n_187);
  and g840 (n648, n_207, n647);
  and g846 (n654, n_131, n653);
  and g847 (n655, n_217, n654);
  not g856 (n_265, n598);
  not g857 (n_266, n663);
  and g858 (n664, n_265, n_266);
  not g859 (n_267, n664);
  and g860 (n665, n_230, n_267);
  not g861 (n_268, n60);
  and g862 (n666, n_49, n_268);
  not g863 (n_269, n666);
  and g864 (n667, \a[11] , n_269);
  and g865 (n668, n_26, n666);
  not g866 (n_270, n667);
  not g867 (n_271, n668);
  and g868 (n669, n_270, n_271);
  not g869 (n_272, n669);
  and g870 (n670, n_248, n_272);
  not g871 (n_273, n665);
  and g872 (n671, n_273, n670);
  not g873 (n_274, n670);
  and g874 (n672, n665, n_274);
  not g875 (n_275, n671);
  not g876 (n_276, n672);
  and g877 (n673, n_275, n_276);
  and g878 (n674, \a[12] , \a[22] );
  not g879 (n_277, n61);
  and g880 (n675, \a[12] , n_277);
  not g881 (n_278, n675);
  and g882 (n676, n526, n_278);
  not g883 (n_279, n674);
  not g884 (n_280, n676);
  and g885 (n677, n_279, n_280);
  not g886 (n_281, n677);
  and g887 (n678, n_248, n_281);
  and g888 (n679, n673, n678);
  not g889 (n_282, n679);
  and g890 (n680, n_275, n_282);
  not g891 (n_283, n550);
  not g892 (n_284, n680);
  and g893 (n681, n_283, n_284);
  not g894 (n_285, n551);
  and g895 (n682, n_285, n681);
  not g896 (n_286, n682);
  and g897 (n683, n_283, n_286);
  and g898 (n684, n_253, n_252);
  and g899 (n685, n_240, n684);
  and g900 (n686, n525, n545);
  and g901 (n687, n539, n_254);
  and g902 (n688, n529, n687);
  and g903 (n689, n_241, n542);
  and g911 (n693, n598, n_266);
  and g912 (n694, n_265, n663);
  not g913 (n_291, n693);
  not g914 (n_292, n694);
  and g915 (n695, n_291, n_292);
  and g916 (n696, n598, n663);
  not g917 (n_293, n696);
  and g918 (n697, n494, n_293);
  not g919 (n_294, n697);
  and g920 (n698, n695, n_294);
  and g921 (n699, n_240, n698);
  not g922 (n_295, n695);
  and g923 (n700, n_273, n_295);
  and g924 (n701, n525, n_273);
  not g925 (n_296, n700);
  not g926 (n_297, n701);
  and g927 (n702, n_296, n_297);
  not g928 (n_298, n699);
  and g929 (n703, n_298, n702);
  and g930 (n704, n_274, n703);
  and g931 (n705, n_241, n684);
  and g932 (n706, n529, n545);
  and g933 (n707, n677, n687);
  and g934 (n708, n542, n_281);
  not g942 (n_303, n703);
  and g943 (n712, n670, n_303);
  not g944 (n_304, n704);
  not g945 (n_305, n712);
  and g946 (n713, n_304, n_305);
  and g947 (n714, n711, n713);
  not g948 (n_306, n714);
  and g949 (n715, n_304, n_306);
  not g950 (n_307, n715);
  and g951 (n716, n692, n_307);
  not g952 (n_308, n692);
  and g953 (n717, n_308, n715);
  not g954 (n_309, n716);
  not g955 (n_310, n717);
  and g956 (n718, n_309, n_310);
  not g957 (n_311, n673);
  not g958 (n_312, n678);
  and g959 (n719, n_311, n_312);
  not g960 (n_313, n719);
  and g961 (n720, n_282, n_313);
  and g962 (n721, n718, n720);
  not g963 (n_314, n721);
  and g964 (n722, n_309, n_314);
  and g965 (n723, n_284, n_286);
  and g966 (n724, n_285, n683);
  not g967 (n_315, n723);
  not g968 (n_316, n724);
  and g969 (n725, n_315, n_316);
  not g970 (n_317, n722);
  and g971 (n726, n_317, n725);
  not g972 (n_318, n725);
  and g973 (n727, n722, n_318);
  not g974 (n_319, n726);
  not g975 (n_320, n727);
  and g976 (n728, n_319, n_320);
  and g984 (n736, n130, n193);
  not g987 (n_321, n736);
  and g1002 (n753, n_97, n_179);
  and g1007 (n758, n_98, n_139);
  and g1008 (n759, n_135, n758);
  and g1009 (n760, n_138, n_220);
  and g1023 (n774, n_136, n_211);
  and g1024 (n775, n_177, n774);
  and g1025 (n776, n_140, n_176);
  and g1026 (n777, n_121, n776);
  and g1036 (n787, n_114, n_120);
  and g1037 (n788, n_126, n787);
  and g1038 (n789, n_219, n788);
  and g1042 (n793, n_149, n_100);
  and g1043 (n794, n_222, n793);
  and g1044 (n795, n_95, n_99);
  and g1045 (n796, n_138, n795);
  and g1055 (n806, n_121, n_178);
  and g1056 (n807, n_146, n_101);
  and g1057 (n808, n_86, n_192);
  and g1058 (n809, n_217, n_262);
  and g1063 (n814, n_180, n813);
  and g1064 (n815, n_117, n814);
  not g1076 (n_322, n786);
  not g1077 (n_323, n826);
  and g1078 (n827, n_322, n_323);
  not g1079 (n_324, n827);
  and g1080 (n828, n_265, n_324);
  not g1081 (n_325, n58);
  and g1082 (n829, n_49, n_325);
  not g1083 (n_326, n829);
  and g1084 (n830, \a[9] , n_326);
  and g1085 (n831, n_22, n829);
  not g1086 (n_327, n830);
  not g1087 (n_328, n831);
  and g1088 (n832, n_327, n_328);
  not g1089 (n_329, n832);
  and g1090 (n833, n_248, n_329);
  not g1091 (n_330, n828);
  and g1092 (n834, n_330, n833);
  not g1093 (n_331, n833);
  and g1094 (n835, n828, n_331);
  not g1095 (n_332, n834);
  not g1096 (n_333, n835);
  and g1097 (n836, n_332, n_333);
  and g1098 (n837, \a[10] , \a[22] );
  not g1099 (n_334, n59);
  and g1100 (n838, \a[10] , n_334);
  not g1101 (n_335, n838);
  and g1102 (n839, n666, n_335);
  not g1103 (n_336, n837);
  not g1104 (n_337, n839);
  and g1105 (n840, n_336, n_337);
  not g1106 (n_338, n840);
  and g1107 (n841, n_248, n_338);
  and g1108 (n842, n836, n841);
  not g1109 (n_339, n842);
  and g1110 (n843, n_332, n_339);
  and g1111 (n844, n_295, n_294);
  and g1112 (n845, n_240, n844);
  and g1113 (n846, n525, n700);
  and g1114 (n847, n_273, n695);
  and g1115 (n848, n529, n847);
  and g1116 (n849, n_241, n698);
  and g1124 (n853, n_281, n684);
  and g1125 (n854, n545, n677);
  and g1126 (n855, n669, n687);
  and g1127 (n856, n542, n_272);
  and g1135 (n860, n852, n859);
  and g1136 (n861, n786, n_323);
  and g1137 (n862, n_322, n826);
  not g1138 (n_348, n861);
  not g1139 (n_349, n862);
  and g1140 (n863, n_348, n_349);
  and g1141 (n864, n786, n826);
  not g1142 (n_350, n864);
  and g1143 (n865, n598, n_350);
  not g1144 (n_351, n865);
  and g1145 (n866, n863, n_351);
  and g1146 (n867, n_240, n866);
  not g1147 (n_352, n863);
  and g1148 (n868, n_330, n_352);
  and g1149 (n869, n525, n_330);
  not g1150 (n_353, n868);
  not g1151 (n_354, n869);
  and g1152 (n870, n_353, n_354);
  not g1153 (n_355, n867);
  and g1154 (n871, n_355, n870);
  and g1155 (n872, n_331, n871);
  and g1156 (n873, n_241, n844);
  and g1157 (n874, n529, n700);
  and g1158 (n875, n677, n847);
  and g1159 (n876, n_281, n698);
  not g1167 (n_360, n871);
  and g1168 (n880, n833, n_360);
  not g1169 (n_361, n872);
  not g1170 (n_362, n880);
  and g1171 (n881, n_361, n_362);
  and g1172 (n882, n879, n881);
  not g1173 (n_363, n882);
  and g1174 (n883, n_361, n_363);
  not g1175 (n_364, n852);
  not g1176 (n_365, n859);
  and g1177 (n884, n_364, n_365);
  not g1178 (n_366, n860);
  not g1179 (n_367, n884);
  and g1180 (n885, n_366, n_367);
  not g1181 (n_368, n883);
  and g1182 (n886, n_368, n885);
  not g1183 (n_369, n886);
  and g1184 (n887, n_366, n_369);
  not g1185 (n_370, n843);
  not g1186 (n_371, n887);
  and g1187 (n888, n_370, n_371);
  not g1188 (n_372, n888);
  and g1189 (n889, n_370, n_372);
  and g1190 (n890, n_371, n_372);
  not g1191 (n_373, n889);
  not g1192 (n_374, n890);
  and g1193 (n891, n_373, n_374);
  not g1194 (n_375, n711);
  not g1195 (n_376, n713);
  and g1196 (n892, n_375, n_376);
  not g1197 (n_377, n892);
  and g1198 (n893, n_306, n_377);
  not g1199 (n_378, n891);
  and g1200 (n894, n_378, n893);
  not g1201 (n_379, n894);
  and g1202 (n895, n_372, n_379);
  not g1203 (n_380, n718);
  not g1204 (n_381, n720);
  and g1205 (n896, n_380, n_381);
  not g1206 (n_382, n896);
  and g1207 (n897, n_314, n_382);
  not g1208 (n_383, n895);
  and g1209 (n898, n_383, n897);
  and g1210 (n899, n_272, n684);
  and g1211 (n900, n545, n669);
  and g1212 (n901, n687, n840);
  and g1213 (n902, n542, n_338);
  and g1221 (n906, n_114, n_218);
  and g1226 (n911, n_102, n_222);
  and g1246 (n931, n_83, n_189);
  and g1260 (n945, n_112, n_214);
  and g1261 (n946, n_125, n945);
  and g1262 (n947, n_92, n_211);
  and g1263 (n948, n_199, n947);
  and g1275 (n960, n_104, n_200);
  and g1276 (n961, n_215, n960);
  and g1283 (n968, n_96, n_142);
  and g1284 (n969, n_206, n968);
  and g1285 (n970, n_223, n_221);
  and g1291 (n976, n_112, n_177);
  and g1292 (n977, n_102, n976);
  and g1293 (n978, n_111, n977);
  and g1294 (n979, n_105, n978);
  and g1295 (n980, n_128, n_210);
  not g1323 (n_388, n959);
  not g1324 (n_389, n1007);
  and g1325 (n1008, n_388, n_389);
  not g1326 (n_390, n1008);
  and g1327 (n1009, n_322, n_390);
  not g1328 (n_391, n56);
  and g1329 (n1010, n_49, n_391);
  not g1330 (n_392, n1010);
  and g1331 (n1011, \a[7] , n_392);
  and g1332 (n1012, n_18, n1010);
  not g1333 (n_393, n1011);
  not g1334 (n_394, n1012);
  and g1335 (n1013, n_393, n_394);
  not g1336 (n_395, n1013);
  and g1337 (n1014, n_248, n_395);
  not g1338 (n_396, n1009);
  and g1339 (n1015, n_396, n1014);
  not g1340 (n_397, n1014);
  and g1341 (n1016, n1009, n_397);
  not g1342 (n_398, n1015);
  not g1343 (n_399, n1016);
  and g1344 (n1017, n_398, n_399);
  and g1345 (n1018, \a[8] , \a[22] );
  not g1346 (n_400, n57);
  and g1347 (n1019, \a[8] , n_400);
  not g1348 (n_401, n1019);
  and g1349 (n1020, n829, n_401);
  not g1350 (n_402, n1018);
  not g1351 (n_403, n1020);
  and g1352 (n1021, n_402, n_403);
  not g1353 (n_404, n1021);
  and g1354 (n1022, n1017, n_404);
  and g1355 (n1023, n_248, n1022);
  not g1356 (n_405, n1023);
  and g1357 (n1024, n_398, n_405);
  not g1358 (n_406, n1024);
  and g1359 (n1025, n905, n_406);
  and g1360 (n1026, n684, n_338);
  and g1361 (n1027, n545, n840);
  and g1362 (n1028, n687, n832);
  and g1363 (n1029, n542, n_329);
  and g1371 (n1033, n_352, n_351);
  and g1372 (n1034, n_240, n1033);
  and g1373 (n1035, n525, n868);
  and g1374 (n1036, n_330, n863);
  and g1375 (n1037, n529, n1036);
  and g1376 (n1038, n_241, n866);
  and g1384 (n1042, n_281, n844);
  and g1385 (n1043, n677, n700);
  and g1386 (n1044, n669, n847);
  and g1387 (n1045, n_272, n698);
  not g1395 (n_419, n1048);
  and g1396 (n1049, n1041, n_419);
  not g1397 (n_420, n1041);
  and g1398 (n1050, n_420, n1048);
  not g1399 (n_421, n1049);
  not g1400 (n_422, n1050);
  and g1401 (n1051, n_421, n_422);
  not g1402 (n_423, n1051);
  and g1403 (n1052, n1032, n_423);
  and g1404 (n1053, n1041, n1048);
  not g1405 (n_424, n1052);
  not g1406 (n_425, n1053);
  and g1407 (n1054, n_424, n_425);
  not g1408 (n_426, n1025);
  and g1409 (n1055, n905, n_426);
  and g1410 (n1056, n_406, n_426);
  not g1411 (n_427, n1055);
  not g1412 (n_428, n1056);
  and g1413 (n1057, n_427, n_428);
  not g1414 (n_429, n1054);
  not g1415 (n_430, n1057);
  and g1416 (n1058, n_429, n_430);
  not g1417 (n_431, n1058);
  and g1418 (n1059, n_426, n_431);
  not g1419 (n_432, n836);
  not g1420 (n_433, n841);
  and g1421 (n1060, n_432, n_433);
  not g1422 (n_434, n1060);
  and g1423 (n1061, n_339, n_434);
  not g1424 (n_435, n1059);
  and g1425 (n1062, n_435, n1061);
  not g1426 (n_436, n1061);
  and g1427 (n1063, n1059, n_436);
  not g1428 (n_437, n1062);
  not g1429 (n_438, n1063);
  and g1430 (n1064, n_437, n_438);
  not g1431 (n_439, n885);
  and g1432 (n1065, n883, n_439);
  not g1433 (n_440, n1065);
  and g1434 (n1066, n_369, n_440);
  and g1435 (n1067, n1064, n1066);
  not g1436 (n_441, n1067);
  and g1437 (n1068, n_437, n_441);
  and g1438 (n1069, n_378, n_379);
  and g1439 (n1070, n893, n_379);
  not g1440 (n_442, n1069);
  not g1441 (n_443, n1070);
  and g1442 (n1071, n_442, n_443);
  not g1443 (n_444, n1068);
  and g1444 (n1072, n_444, n1071);
  not g1445 (n_445, n1071);
  and g1446 (n1073, n1068, n_445);
  not g1447 (n_446, n1072);
  not g1448 (n_447, n1073);
  and g1449 (n1074, n_446, n_447);
  and g1450 (n1075, n_272, n844);
  and g1451 (n1076, n669, n700);
  and g1452 (n1077, n840, n847);
  and g1453 (n1078, n698, n_338);
  and g1461 (n1082, n684, n_329);
  and g1462 (n1083, n545, n832);
  and g1463 (n1084, n687, n1021);
  and g1464 (n1085, n542, n_404);
  and g1472 (n1089, n1081, n1088);
  and g1473 (n1090, n_198, n_226);
  and g1474 (n1091, n_193, n1090);
  and g1475 (n1092, n_120, n_218);
  and g1476 (n1093, n_261, n1092);
  and g1488 (n1105, n_147, n395);
  and g1489 (n1106, n_125, n1105);
  and g1490 (n1107, n448, n1106);
  and g1491 (n1108, n_122, n1107);
  and g1499 (n1116, n_123, n_264);
  and g1500 (n1117, n_84, n_192);
  not g1559 (n_456, n1130);
  not g1560 (n_457, n1175);
  and g1561 (n1176, n_456, n_457);
  not g1562 (n_458, n1176);
  and g1563 (n1177, n_388, n_458);
  not g1564 (n_459, n1177);
  and g1565 (n1178, n1130, n_459);
  and g1566 (n1179, n_456, n1177);
  and g1567 (n1180, \a[6] , \a[22] );
  not g1568 (n_460, n55);
  and g1569 (n1181, \a[6] , n_460);
  not g1570 (n_461, n1181);
  and g1571 (n1182, n1010, n_461);
  not g1572 (n_462, n1180);
  not g1573 (n_463, n1182);
  and g1574 (n1183, n_462, n_463);
  not g1575 (n_464, n1183);
  and g1576 (n1184, n_248, n_464);
  not g1577 (n_465, n1178);
  and g1578 (n1185, n_465, n1184);
  not g1579 (n_466, n1179);
  and g1580 (n1186, n_466, n1185);
  not g1581 (n_467, n1186);
  and g1582 (n1187, n_465, n_467);
  not g1583 (n_468, n1081);
  not g1584 (n_469, n1088);
  and g1585 (n1188, n_468, n_469);
  not g1586 (n_470, n1089);
  not g1587 (n_471, n1188);
  and g1588 (n1189, n_470, n_471);
  not g1589 (n_472, n1187);
  and g1590 (n1190, n_472, n1189);
  not g1591 (n_473, n1190);
  and g1592 (n1191, n_470, n_473);
  and g1593 (n1192, n959, n_389);
  and g1594 (n1193, n_388, n1007);
  not g1595 (n_474, n1192);
  not g1596 (n_475, n1193);
  and g1597 (n1194, n_474, n_475);
  and g1598 (n1195, n959, n1007);
  not g1599 (n_476, n1195);
  and g1600 (n1196, n786, n_476);
  not g1601 (n_477, n1196);
  and g1602 (n1197, n1194, n_477);
  and g1603 (n1198, n_240, n1197);
  not g1604 (n_478, n1194);
  and g1605 (n1199, n_396, n_478);
  and g1606 (n1200, n525, n_396);
  not g1607 (n_479, n1199);
  not g1608 (n_480, n1200);
  and g1609 (n1201, n_479, n_480);
  not g1610 (n_481, n1198);
  and g1611 (n1202, n_481, n1201);
  and g1612 (n1203, n_397, n1202);
  and g1613 (n1204, n_241, n1033);
  and g1614 (n1205, n529, n868);
  and g1615 (n1206, n677, n1036);
  and g1616 (n1207, n_281, n866);
  not g1624 (n_486, n1202);
  and g1625 (n1211, n1014, n_486);
  not g1626 (n_487, n1203);
  not g1627 (n_488, n1211);
  and g1628 (n1212, n_487, n_488);
  and g1629 (n1213, n1210, n1212);
  not g1630 (n_489, n1213);
  and g1631 (n1214, n_487, n_489);
  not g1632 (n_490, n1191);
  not g1633 (n_491, n1214);
  and g1634 (n1215, n_490, n_491);
  not g1635 (n_492, n1215);
  and g1636 (n1216, n_490, n_492);
  and g1637 (n1217, n_491, n_492);
  not g1638 (n_493, n1216);
  not g1639 (n_494, n1217);
  and g1640 (n1218, n_493, n_494);
  and g1641 (n1219, n_248, n_405);
  and g1642 (n1220, n_404, n1219);
  and g1643 (n1221, n1017, n_405);
  not g1644 (n_495, n1220);
  not g1645 (n_496, n1221);
  and g1646 (n1222, n_495, n_496);
  not g1647 (n_497, n1218);
  not g1648 (n_498, n1222);
  and g1649 (n1223, n_497, n_498);
  not g1650 (n_499, n1223);
  and g1651 (n1224, n_492, n_499);
  not g1652 (n_500, n879);
  not g1653 (n_501, n881);
  and g1654 (n1225, n_500, n_501);
  not g1655 (n_502, n1225);
  and g1656 (n1226, n_363, n_502);
  not g1657 (n_503, n1224);
  and g1658 (n1227, n_503, n1226);
  and g1659 (n1228, n_429, n_431);
  and g1660 (n1229, n_430, n_431);
  not g1661 (n_504, n1228);
  not g1662 (n_505, n1229);
  and g1663 (n1230, n_504, n_505);
  not g1664 (n_506, n1226);
  and g1665 (n1231, n1224, n_506);
  not g1666 (n_507, n1227);
  not g1667 (n_508, n1231);
  and g1668 (n1232, n_507, n_508);
  not g1669 (n_509, n1230);
  and g1670 (n1233, n_509, n1232);
  not g1671 (n_510, n1233);
  and g1672 (n1234, n_507, n_510);
  not g1673 (n_511, n1064);
  not g1674 (n_512, n1066);
  and g1675 (n1235, n_511, n_512);
  not g1676 (n_513, n1235);
  and g1677 (n1236, n_441, n_513);
  not g1678 (n_514, n1234);
  and g1679 (n1237, n_514, n1236);
  and g1680 (n1238, n1232, n_510);
  and g1681 (n1239, n_509, n_510);
  not g1682 (n_515, n1238);
  not g1683 (n_516, n1239);
  and g1684 (n1240, n_515, n_516);
  and g1685 (n1241, n_478, n_477);
  and g1686 (n1242, n_240, n1241);
  and g1687 (n1243, n525, n1199);
  and g1688 (n1244, n_396, n1194);
  and g1689 (n1245, n529, n1244);
  and g1690 (n1246, n_241, n1197);
  and g1698 (n1250, n_338, n844);
  and g1699 (n1251, n700, n840);
  and g1700 (n1252, n832, n847);
  and g1701 (n1253, n698, n_329);
  and g1709 (n1257, n684, n_404);
  and g1710 (n1258, n545, n1021);
  and g1711 (n1259, n687, n1013);
  and g1712 (n1260, n542, n_395);
  not g1720 (n_529, n1263);
  and g1721 (n1264, n1256, n_529);
  not g1722 (n_530, n1256);
  and g1723 (n1265, n_530, n1263);
  not g1724 (n_531, n1264);
  not g1725 (n_532, n1265);
  and g1726 (n1266, n_531, n_532);
  not g1727 (n_533, n1266);
  and g1728 (n1267, n1249, n_533);
  and g1729 (n1268, n1256, n1263);
  not g1730 (n_534, n1267);
  not g1731 (n_535, n1268);
  and g1732 (n1269, n_534, n_535);
  not g1733 (n_536, n1210);
  not g1734 (n_537, n1212);
  and g1735 (n1270, n_536, n_537);
  not g1736 (n_538, n1270);
  and g1737 (n1271, n_489, n_538);
  not g1738 (n_539, n1269);
  and g1739 (n1272, n_539, n1271);
  not g1740 (n_540, n1272);
  and g1741 (n1273, n_539, n_540);
  and g1742 (n1274, n1271, n_540);
  not g1743 (n_541, n1273);
  not g1744 (n_542, n1274);
  and g1745 (n1275, n_541, n_542);
  not g1746 (n_543, n1189);
  and g1747 (n1276, n1187, n_543);
  not g1748 (n_544, n1276);
  and g1749 (n1277, n_473, n_544);
  not g1750 (n_545, n1275);
  and g1751 (n1278, n_545, n1277);
  not g1752 (n_546, n1278);
  and g1753 (n1279, n_540, n_546);
  and g1754 (n1280, n1032, n_424);
  and g1755 (n1281, n_423, n_424);
  not g1756 (n_547, n1280);
  not g1757 (n_548, n1281);
  and g1758 (n1282, n_547, n_548);
  not g1759 (n_549, n1279);
  not g1760 (n_550, n1282);
  and g1761 (n1283, n_549, n_550);
  not g1762 (n_551, n1283);
  and g1763 (n1284, n_549, n_551);
  and g1764 (n1285, n_550, n_551);
  not g1765 (n_552, n1284);
  not g1766 (n_553, n1285);
  and g1767 (n1286, n_552, n_553);
  and g1768 (n1287, n_497, n_499);
  and g1769 (n1288, n_498, n_499);
  not g1770 (n_554, n1287);
  not g1771 (n_555, n1288);
  and g1772 (n1289, n_554, n_555);
  not g1773 (n_556, n1286);
  not g1774 (n_557, n1289);
  and g1775 (n1290, n_556, n_557);
  not g1776 (n_558, n1290);
  and g1777 (n1291, n_551, n_558);
  not g1778 (n_559, n1240);
  not g1779 (n_560, n1291);
  and g1780 (n1292, n_559, n_560);
  not g1781 (n_561, n1292);
  and g1782 (n1293, n_559, n_561);
  and g1783 (n1294, n_560, n_561);
  not g1784 (n_562, n1293);
  not g1785 (n_563, n1294);
  and g1786 (n1295, n_562, n_563);
  and g1787 (n1296, n_281, n1033);
  and g1788 (n1297, n677, n868);
  and g1789 (n1298, n669, n1036);
  and g1790 (n1299, n_272, n866);
  and g1798 (n1303, n_466, n1187);
  and g1799 (n1304, n1184, n_467);
  not g1800 (n_568, n1303);
  not g1801 (n_569, n1304);
  and g1802 (n1305, n_568, n_569);
  not g1803 (n_570, n1305);
  and g1804 (n1306, n1302, n_570);
  and g1805 (n1307, n_160, n_248);
  and g1806 (n1308, n_456, n1307);
  not g1807 (n_571, n1307);
  and g1808 (n1309, n1130, n_571);
  and g1809 (n1310, n1130, n_457);
  and g1810 (n1311, n_456, n1175);
  not g1811 (n_572, n1310);
  not g1812 (n_573, n1311);
  and g1813 (n1312, n_572, n_573);
  and g1814 (n1313, n1130, n1175);
  not g1815 (n_574, n1313);
  and g1816 (n1314, n959, n_574);
  not g1817 (n_575, n1314);
  and g1818 (n1315, n1312, n_575);
  and g1819 (n1316, n_240, n1315);
  not g1820 (n_576, n1312);
  and g1821 (n1317, n_459, n_576);
  and g1822 (n1318, n525, n_459);
  not g1823 (n_577, n1317);
  not g1824 (n_578, n1318);
  and g1825 (n1319, n_577, n_578);
  not g1826 (n_579, n1316);
  and g1827 (n1320, n_579, n1319);
  not g1828 (n_580, n1308);
  and g1829 (n1321, n_580, n1320);
  not g1830 (n_581, n1309);
  and g1831 (n1322, n_581, n1321);
  not g1832 (n_582, n1322);
  and g1833 (n1323, n_580, n_582);
  not g1834 (n_583, n1302);
  and g1835 (n1324, n_583, n1305);
  not g1836 (n_584, n1306);
  not g1837 (n_585, n1324);
  and g1838 (n1325, n_584, n_585);
  not g1839 (n_586, n1323);
  and g1840 (n1326, n_586, n1325);
  not g1841 (n_587, n1326);
  and g1842 (n1327, n_584, n_587);
  and g1843 (n1328, n_241, n1241);
  and g1844 (n1329, n529, n1199);
  and g1845 (n1330, n677, n1244);
  and g1846 (n1331, n_281, n1197);
  and g1854 (n1335, n_272, n1033);
  and g1855 (n1336, n669, n868);
  and g1856 (n1337, n840, n1036);
  and g1857 (n1338, n_338, n866);
  and g1865 (n1342, n1334, n1341);
  and g1866 (n1343, n_329, n844);
  and g1867 (n1344, n700, n832);
  and g1868 (n1345, n847, n1021);
  and g1869 (n1346, n698, n_404);
  not g1877 (n_600, n1341);
  and g1878 (n1350, n1334, n_600);
  not g1879 (n_601, n1334);
  and g1880 (n1351, n_601, n1341);
  not g1881 (n_602, n1350);
  not g1882 (n_603, n1351);
  and g1883 (n1352, n_602, n_603);
  not g1884 (n_604, n1352);
  and g1885 (n1353, n1349, n_604);
  not g1886 (n_605, n1342);
  not g1887 (n_606, n1353);
  and g1888 (n1354, n_605, n_606);
  not g1889 (n_607, n1249);
  and g1890 (n1355, n_607, n1266);
  not g1891 (n_608, n1355);
  and g1892 (n1356, n_534, n_608);
  not g1893 (n_609, n1354);
  and g1894 (n1357, n_609, n1356);
  and g1895 (n1358, n684, n_395);
  and g1896 (n1359, n545, n1013);
  and g1897 (n1360, n687, n1183);
  and g1898 (n1361, n542, n_464);
  and g1906 (n1365, n_159, n_248);
  and g1907 (n1366, n_456, n1365);
  not g1908 (n_614, n1365);
  and g1909 (n1367, n1130, n_614);
  and g1910 (n1368, n_576, n_575);
  and g1911 (n1369, n_240, n1368);
  and g1912 (n1370, n525, n1317);
  and g1913 (n1371, n_459, n1312);
  and g1914 (n1372, n529, n1371);
  and g1915 (n1373, n_241, n1315);
  not g1923 (n_619, n1366);
  and g1924 (n1377, n_619, n1376);
  not g1925 (n_620, n1367);
  and g1926 (n1378, n_620, n1377);
  not g1927 (n_621, n1378);
  and g1928 (n1379, n_619, n_621);
  not g1929 (n_622, n1379);
  and g1930 (n1380, n1364, n_622);
  not g1931 (n_623, n1364);
  and g1932 (n1381, n_623, n1379);
  not g1933 (n_624, n1380);
  not g1934 (n_625, n1381);
  and g1935 (n1382, n_624, n_625);
  and g1936 (n1383, n_338, n1033);
  and g1937 (n1384, n840, n868);
  and g1938 (n1385, n832, n1036);
  and g1939 (n1386, n_329, n866);
  and g1947 (n1390, n_281, n1241);
  and g1948 (n1391, n677, n1199);
  and g1949 (n1392, n669, n1244);
  and g1950 (n1393, n_272, n1197);
  and g1958 (n1397, n1389, n1396);
  and g1959 (n1398, n844, n_404);
  and g1960 (n1399, n700, n1021);
  and g1961 (n1400, n847, n1013);
  and g1962 (n1401, n698, n_395);
  not g1970 (n_638, n1389);
  and g1971 (n1405, n_638, n1396);
  not g1972 (n_639, n1396);
  and g1973 (n1406, n1389, n_639);
  not g1974 (n_640, n1405);
  not g1975 (n_641, n1406);
  and g1976 (n1407, n_640, n_641);
  not g1977 (n_642, n1407);
  and g1978 (n1408, n1404, n_642);
  not g1979 (n_643, n1397);
  not g1980 (n_644, n1408);
  and g1981 (n1409, n_643, n_644);
  not g1982 (n_645, n1409);
  and g1983 (n1410, n1382, n_645);
  not g1984 (n_646, n1410);
  and g1985 (n1411, n_624, n_646);
  not g1986 (n_647, n1356);
  and g1987 (n1412, n1354, n_647);
  not g1988 (n_648, n1357);
  not g1989 (n_649, n1412);
  and g1990 (n1413, n_648, n_649);
  not g1991 (n_650, n1411);
  and g1992 (n1414, n_650, n1413);
  not g1993 (n_651, n1414);
  and g1994 (n1415, n_648, n_651);
  not g1995 (n_652, n1327);
  not g1996 (n_653, n1415);
  and g1997 (n1416, n_652, n_653);
  not g1998 (n_654, n1416);
  and g1999 (n1417, n_652, n_654);
  and g2000 (n1418, n_653, n_654);
  not g2001 (n_655, n1417);
  not g2002 (n_656, n1418);
  and g2003 (n1419, n_655, n_656);
  and g2004 (n1420, n1277, n_546);
  and g2005 (n1421, n_545, n_546);
  not g2006 (n_657, n1420);
  not g2007 (n_658, n1421);
  and g2008 (n1422, n_657, n_658);
  not g2009 (n_659, n1419);
  not g2010 (n_660, n1422);
  and g2011 (n1423, n_659, n_660);
  not g2012 (n_661, n1423);
  and g2013 (n1424, n_654, n_661);
  and g2014 (n1425, n_556, n1289);
  and g2015 (n1426, n1286, n_557);
  not g2016 (n_662, n1425);
  not g2017 (n_663, n1426);
  and g2018 (n1427, n_662, n_663);
  not g2019 (n_664, n1424);
  not g2020 (n_665, n1427);
  and g2021 (n1428, n_664, n_665);
  and g2022 (n1429, n_659, n_661);
  and g2023 (n1430, n_660, n_661);
  not g2024 (n_666, n1429);
  not g2025 (n_667, n1430);
  and g2026 (n1431, n_666, n_667);
  and g2027 (n1432, n_581, n1323);
  and g2028 (n1433, n1320, n_582);
  not g2029 (n_668, n1432);
  not g2030 (n_669, n1433);
  and g2031 (n1434, n_668, n_669);
  and g2032 (n1435, n1349, n_606);
  and g2033 (n1436, n_604, n_606);
  not g2034 (n_670, n1435);
  not g2035 (n_671, n1436);
  and g2036 (n1437, n_670, n_671);
  not g2037 (n_672, n1434);
  not g2038 (n_673, n1437);
  and g2039 (n1438, n_672, n_673);
  not g2040 (n_674, n1438);
  and g2041 (n1439, n_672, n_674);
  and g2042 (n1440, n_673, n_674);
  not g2043 (n_675, n1439);
  not g2044 (n_676, n1440);
  and g2045 (n1441, n_675, n_676);
  and g2046 (n1442, n684, n_464);
  and g2047 (n1443, n545, n1183);
  and g2048 (n1444, n275, n687);
  and g2049 (n1445, n_160, n542);
  and g2057 (n1449, n_172, n_248);
  and g2066 (n1458, n_130, n_209);
  and g2067 (n1459, n_183, n1458);
  and g2096 (n1488, n_240, n1487);
  not g2097 (n_681, n1488);
  and g2098 (n1489, n_456, n_681);
  and g2099 (n1490, n1449, n1489);
  and g2100 (n1491, n_241, n1368);
  and g2101 (n1492, n529, n1317);
  and g2102 (n1493, n677, n1371);
  and g2103 (n1494, n_281, n1315);
  not g2111 (n_686, n1449);
  not g2112 (n_687, n1489);
  and g2113 (n1498, n_686, n_687);
  not g2114 (n_688, n1490);
  not g2115 (n_689, n1498);
  and g2116 (n1499, n_688, n_689);
  and g2117 (n1500, n1497, n1499);
  not g2118 (n_690, n1500);
  and g2119 (n1501, n_688, n_690);
  not g2120 (n_691, n1501);
  and g2121 (n1502, n1448, n_691);
  not g2122 (n_692, n1448);
  and g2123 (n1503, n_692, n1501);
  not g2124 (n_693, n1502);
  not g2125 (n_694, n1503);
  and g2126 (n1504, n_693, n_694);
  and g2127 (n1505, n_329, n1033);
  and g2128 (n1506, n832, n868);
  and g2129 (n1507, n1021, n1036);
  and g2130 (n1508, n866, n_404);
  and g2138 (n1512, n_272, n1241);
  and g2139 (n1513, n669, n1199);
  and g2140 (n1514, n840, n1244);
  and g2141 (n1515, n_338, n1197);
  and g2149 (n1519, n1511, n1518);
  and g2150 (n1520, n844, n_395);
  and g2151 (n1521, n700, n1013);
  and g2152 (n1522, n847, n1183);
  and g2153 (n1523, n698, n_464);
  not g2161 (n_707, n1511);
  and g2162 (n1527, n_707, n1518);
  not g2163 (n_708, n1518);
  and g2164 (n1528, n1511, n_708);
  not g2165 (n_709, n1527);
  not g2166 (n_710, n1528);
  and g2167 (n1529, n_709, n_710);
  not g2168 (n_711, n1529);
  and g2169 (n1530, n1526, n_711);
  not g2170 (n_712, n1519);
  not g2171 (n_713, n1530);
  and g2172 (n1531, n_712, n_713);
  not g2173 (n_714, n1531);
  and g2174 (n1532, n1504, n_714);
  not g2175 (n_715, n1532);
  and g2176 (n1533, n_693, n_715);
  not g2177 (n_716, n1441);
  not g2178 (n_717, n1533);
  and g2179 (n1534, n_716, n_717);
  not g2180 (n_718, n1534);
  and g2181 (n1535, n_674, n_718);
  not g2182 (n_719, n1325);
  and g2183 (n1536, n1323, n_719);
  not g2184 (n_720, n1536);
  and g2185 (n1537, n_587, n_720);
  not g2186 (n_721, n1535);
  and g2187 (n1538, n_721, n1537);
  not g2188 (n_722, n1537);
  and g2189 (n1539, n1535, n_722);
  not g2190 (n_723, n1538);
  not g2191 (n_724, n1539);
  and g2192 (n1540, n_723, n_724);
  not g2193 (n_725, n1413);
  and g2194 (n1541, n1411, n_725);
  not g2195 (n_726, n1541);
  and g2196 (n1542, n_651, n_726);
  and g2197 (n1543, n1540, n1542);
  not g2198 (n_727, n1543);
  and g2199 (n1544, n_723, n_727);
  not g2200 (n_728, n1431);
  not g2201 (n_729, n1544);
  and g2202 (n1545, n_728, n_729);
  and g2203 (n1546, n1431, n_729);
  and g2204 (n1547, n_728, n1544);
  not g2205 (n_730, n1546);
  not g2206 (n_731, n1547);
  and g2207 (n1548, n_730, n_731);
  not g2208 (n_732, n1487);
  and g2209 (n1549, n1130, n_732);
  not g2210 (n_733, n1549);
  and g2211 (n1550, n_732, n_733);
  and g2212 (n1551, n_240, n1550);
  and g2213 (n1552, n525, n1549);
  and g2214 (n1553, n529, n_456);
  not g2215 (n_734, n1553);
  and g2216 (n1554, n1487, n_734);
  not g2217 (n_735, n1552);
  not g2218 (n_736, n1554);
  and g2219 (n1555, n_735, n_736);
  not g2220 (n_737, n1551);
  and g2221 (n1556, n_737, n1555);
  and g2222 (n1557, n_172, n684);
  and g2223 (n1558, n286, n_254);
  not g2224 (n_738, n687);
  not g2225 (n_739, n1558);
  and g2226 (n1559, n_738, n_739);
  not g2227 (n_740, n1557);
  and g2228 (n1560, n_740, n1559);
  and g2229 (n1561, n544, n1560);
  and g2230 (n1562, n1556, n1561);
  and g2231 (n1563, n_160, n684);
  and g2232 (n1564, n275, n545);
  and g2233 (n1565, n279, n687);
  and g2234 (n1566, n_159, n542);
  and g2242 (n1570, n1562, n1569);
  and g2243 (n1571, n_338, n1241);
  and g2244 (n1572, n840, n1199);
  and g2245 (n1573, n832, n1244);
  and g2246 (n1574, n_329, n1197);
  and g2254 (n1578, n_404, n1033);
  and g2255 (n1579, n868, n1021);
  and g2256 (n1580, n1013, n1036);
  and g2257 (n1581, n866, n_395);
  and g2265 (n1585, n844, n_464);
  and g2266 (n1586, n700, n1183);
  and g2267 (n1587, n275, n847);
  and g2268 (n1588, n_160, n698);
  not g2276 (n_757, n1591);
  and g2277 (n1592, n1584, n_757);
  not g2278 (n_758, n1584);
  and g2279 (n1593, n_758, n1591);
  not g2280 (n_759, n1592);
  not g2281 (n_760, n1593);
  and g2282 (n1594, n_759, n_760);
  not g2283 (n_761, n1594);
  and g2284 (n1595, n1577, n_761);
  and g2285 (n1596, n1584, n1591);
  not g2286 (n_762, n1595);
  not g2287 (n_763, n1596);
  and g2288 (n1597, n_762, n_763);
  not g2289 (n_764, n1562);
  not g2290 (n_765, n1569);
  and g2291 (n1598, n_764, n_765);
  not g2292 (n_766, n1570);
  not g2293 (n_767, n1598);
  and g2294 (n1599, n_766, n_767);
  not g2295 (n_768, n1597);
  and g2296 (n1600, n_768, n1599);
  not g2297 (n_769, n1600);
  and g2298 (n1601, n_766, n_769);
  and g2299 (n1602, n_620, n1379);
  and g2300 (n1603, n1376, n_621);
  not g2301 (n_770, n1602);
  not g2302 (n_771, n1603);
  and g2303 (n1604, n_770, n_771);
  not g2304 (n_772, n1604);
  and g2305 (n1605, n1601, n_772);
  not g2306 (n_773, n1601);
  and g2307 (n1606, n_773, n1604);
  not g2308 (n_774, n1605);
  not g2309 (n_775, n1606);
  and g2310 (n1607, n_774, n_775);
  and g2311 (n1608, n1404, n_644);
  and g2312 (n1609, n_642, n_644);
  not g2313 (n_776, n1608);
  not g2314 (n_777, n1609);
  and g2315 (n1610, n_776, n_777);
  not g2316 (n_778, n1607);
  not g2317 (n_779, n1610);
  and g2318 (n1611, n_778, n_779);
  and g2319 (n1612, n_773, n_772);
  not g2320 (n_780, n1611);
  not g2321 (n_781, n1612);
  and g2322 (n1613, n_780, n_781);
  not g2323 (n_782, n1382);
  and g2324 (n1614, n_782, n1409);
  not g2325 (n_783, n1614);
  and g2326 (n1615, n_646, n_783);
  not g2327 (n_784, n1613);
  and g2328 (n1616, n_784, n1615);
  and g2329 (n1617, n1441, n_717);
  and g2330 (n1618, n_716, n1533);
  not g2331 (n_785, n1617);
  not g2332 (n_786, n1618);
  and g2333 (n1619, n_785, n_786);
  not g2334 (n_787, n1615);
  and g2335 (n1620, n1613, n_787);
  not g2336 (n_788, n1616);
  not g2337 (n_789, n1620);
  and g2338 (n1621, n_788, n_789);
  not g2339 (n_790, n1619);
  and g2340 (n1622, n_790, n1621);
  not g2341 (n_791, n1622);
  and g2342 (n1623, n_788, n_791);
  not g2343 (n_792, n1540);
  not g2344 (n_793, n1542);
  and g2345 (n1624, n_792, n_793);
  not g2346 (n_794, n1624);
  and g2347 (n1625, n_727, n_794);
  not g2348 (n_795, n1623);
  and g2349 (n1626, n_795, n1625);
  and g2350 (n1627, n_281, n1368);
  and g2351 (n1628, n677, n1317);
  and g2352 (n1629, n669, n1371);
  and g2353 (n1630, n_272, n1315);
  and g2361 (n1634, n_159, n684);
  and g2362 (n1635, n279, n545);
  and g2363 (n1636, n286, n687);
  and g2364 (n1637, n_172, n542);
  and g2372 (n1641, n1633, n1640);
  not g2373 (n_804, n1556);
  not g2374 (n_805, n1561);
  and g2375 (n1642, n_804, n_805);
  not g2376 (n_806, n1642);
  and g2377 (n1643, n_764, n_806);
  not g2378 (n_807, n1633);
  not g2379 (n_808, n1640);
  and g2380 (n1644, n_807, n_808);
  not g2381 (n_809, n1641);
  not g2382 (n_810, n1644);
  and g2383 (n1645, n_809, n_810);
  and g2384 (n1646, n1643, n1645);
  not g2385 (n_811, n1646);
  and g2386 (n1647, n_809, n_811);
  not g2387 (n_812, n1497);
  not g2388 (n_813, n1499);
  and g2389 (n1648, n_812, n_813);
  not g2390 (n_814, n1648);
  and g2391 (n1649, n_690, n_814);
  not g2392 (n_815, n1647);
  and g2393 (n1650, n_815, n1649);
  not g2394 (n_816, n1649);
  and g2395 (n1651, n1647, n_816);
  not g2396 (n_817, n1650);
  not g2397 (n_818, n1651);
  and g2398 (n1652, n_817, n_818);
  and g2399 (n1653, n1526, n_713);
  and g2400 (n1654, n_711, n_713);
  not g2401 (n_819, n1653);
  not g2402 (n_820, n1654);
  and g2403 (n1655, n_819, n_820);
  not g2404 (n_821, n1655);
  and g2405 (n1656, n1652, n_821);
  not g2406 (n_822, n1656);
  and g2407 (n1657, n_817, n_822);
  not g2408 (n_823, n1504);
  and g2409 (n1658, n_823, n1531);
  not g2410 (n_824, n1658);
  and g2411 (n1659, n_715, n_824);
  not g2412 (n_825, n1657);
  and g2413 (n1660, n_825, n1659);
  not g2414 (n_826, n1659);
  and g2415 (n1661, n1657, n_826);
  not g2416 (n_827, n1660);
  not g2417 (n_828, n1661);
  and g2418 (n1662, n_827, n_828);
  and g2419 (n1663, n1607, n1610);
  not g2420 (n_829, n1663);
  and g2421 (n1664, n_780, n_829);
  and g2422 (n1665, n1662, n1664);
  not g2423 (n_830, n1665);
  and g2424 (n1666, n_827, n_830);
  not g2425 (n_831, n1621);
  and g2426 (n1667, n1619, n_831);
  not g2427 (n_832, n1667);
  and g2428 (n1668, n_791, n_832);
  not g2429 (n_833, n1666);
  and g2430 (n1669, n_833, n1668);
  and g2431 (n1670, n_281, n1550);
  and g2432 (n1671, n677, n1549);
  and g2433 (n1672, n669, n_456);
  not g2434 (n_834, n1672);
  and g2435 (n1673, n1487, n_834);
  not g2436 (n_835, n1671);
  not g2437 (n_836, n1673);
  and g2438 (n1674, n_835, n_836);
  not g2439 (n_837, n1670);
  and g2440 (n1675, n_837, n1674);
  and g2441 (n1676, n_172, n844);
  and g2442 (n1677, n286, n_273);
  and g2449 (n1681, n1675, n1680);
  and g2450 (n1682, n_329, n1241);
  and g2451 (n1683, n832, n1199);
  and g2452 (n1684, n1021, n1244);
  and g2453 (n1685, n_404, n1197);
  and g2461 (n1689, n_395, n1033);
  and g2462 (n1690, n868, n1013);
  and g2463 (n1691, n1036, n1183);
  and g2464 (n1692, n866, n_464);
  not g2472 (n_849, n1695);
  and g2473 (n1696, n1688, n_849);
  not g2474 (n_850, n1688);
  and g2475 (n1697, n_850, n1695);
  not g2476 (n_851, n1696);
  not g2477 (n_852, n1697);
  and g2478 (n1698, n_851, n_852);
  not g2479 (n_853, n1698);
  and g2480 (n1699, n1681, n_853);
  and g2481 (n1700, n1688, n1695);
  not g2482 (n_854, n1699);
  not g2483 (n_855, n1700);
  and g2484 (n1701, n_854, n_855);
  and g2485 (n1702, n_160, n844);
  and g2486 (n1703, n275, n700);
  and g2487 (n1704, n279, n847);
  and g2488 (n1705, n_159, n698);
  and g2496 (n1709, n_241, n1550);
  and g2497 (n1710, n529, n1549);
  and g2498 (n1711, n677, n_456);
  not g2499 (n_860, n1711);
  and g2500 (n1712, n1487, n_860);
  not g2501 (n_861, n1710);
  not g2502 (n_862, n1712);
  and g2503 (n1713, n_861, n_862);
  not g2504 (n_863, n1709);
  and g2505 (n1714, n_863, n1713);
  and g2506 (n1715, n_272, n1368);
  and g2507 (n1716, n669, n1317);
  and g2508 (n1717, n840, n1371);
  and g2509 (n1718, n_338, n1315);
  not g2517 (n_868, n1721);
  and g2518 (n1722, n1714, n_868);
  not g2519 (n_869, n1714);
  and g2520 (n1723, n_869, n1721);
  not g2521 (n_870, n1722);
  not g2522 (n_871, n1723);
  and g2523 (n1724, n_870, n_871);
  not g2524 (n_872, n1724);
  and g2525 (n1725, n1708, n_872);
  and g2526 (n1726, n1714, n1721);
  not g2527 (n_873, n1725);
  not g2528 (n_874, n1726);
  and g2529 (n1727, n_873, n_874);
  not g2530 (n_875, n1701);
  not g2531 (n_876, n1727);
  and g2532 (n1728, n_875, n_876);
  not g2533 (n_877, n1728);
  and g2534 (n1729, n_875, n_877);
  and g2535 (n1730, n_876, n_877);
  not g2536 (n_878, n1729);
  not g2537 (n_879, n1730);
  and g2538 (n1731, n_878, n_879);
  and g2539 (n1732, n1577, n_762);
  and g2540 (n1733, n_761, n_762);
  not g2541 (n_880, n1732);
  not g2542 (n_881, n1733);
  and g2543 (n1734, n_880, n_881);
  not g2544 (n_882, n1731);
  not g2545 (n_883, n1734);
  and g2546 (n1735, n_882, n_883);
  not g2547 (n_884, n1735);
  and g2548 (n1736, n_877, n_884);
  not g2549 (n_885, n1599);
  and g2550 (n1737, n1597, n_885);
  not g2551 (n_886, n1737);
  and g2552 (n1738, n_769, n_886);
  not g2553 (n_887, n1736);
  and g2554 (n1739, n_887, n1738);
  and g2555 (n1740, n1652, n_822);
  and g2556 (n1741, n_821, n_822);
  not g2557 (n_888, n1740);
  not g2558 (n_889, n1741);
  and g2559 (n1742, n_888, n_889);
  not g2560 (n_890, n1738);
  and g2561 (n1743, n1736, n_890);
  not g2562 (n_891, n1739);
  not g2563 (n_892, n1743);
  and g2564 (n1744, n_891, n_892);
  not g2565 (n_893, n1742);
  and g2566 (n1745, n_893, n1744);
  not g2567 (n_894, n1745);
  and g2568 (n1746, n_891, n_894);
  not g2569 (n_895, n1662);
  not g2570 (n_896, n1664);
  and g2571 (n1747, n_895, n_896);
  not g2572 (n_897, n1747);
  and g2573 (n1748, n_830, n_897);
  not g2574 (n_898, n1746);
  and g2575 (n1749, n_898, n1748);
  not g2576 (n_899, n1560);
  and g2577 (n1750, n_254, n_899);
  and g2578 (n1751, n_404, n1241);
  and g2579 (n1752, n1021, n1199);
  and g2580 (n1753, n1013, n1244);
  and g2581 (n1754, n_395, n1197);
  and g2589 (n1758, n_338, n1368);
  and g2590 (n1759, n840, n1317);
  and g2591 (n1760, n832, n1371);
  and g2592 (n1761, n_329, n1315);
  and g2600 (n1765, n1033, n_464);
  and g2601 (n1766, n868, n1183);
  and g2602 (n1767, n275, n1036);
  and g2603 (n1768, n_160, n866);
  not g2611 (n_912, n1771);
  and g2612 (n1772, n1764, n_912);
  not g2613 (n_913, n1764);
  and g2614 (n1773, n_913, n1771);
  not g2615 (n_914, n1772);
  not g2616 (n_915, n1773);
  and g2617 (n1774, n_914, n_915);
  not g2618 (n_916, n1774);
  and g2619 (n1775, n1757, n_916);
  and g2620 (n1776, n1764, n1771);
  not g2621 (n_917, n1775);
  not g2622 (n_918, n1776);
  and g2623 (n1777, n_917, n_918);
  not g2624 (n_919, n1777);
  and g2625 (n1778, n_805, n_919);
  not g2626 (n_920, n1750);
  and g2627 (n1779, n_920, n1778);
  not g2628 (n_921, n1779);
  and g2629 (n1780, n_805, n_921);
  and g2630 (n1781, n_920, n1780);
  and g2631 (n1782, n_919, n_921);
  not g2632 (n_922, n1781);
  not g2633 (n_923, n1782);
  and g2634 (n1783, n_922, n_923);
  not g2635 (n_924, n1681);
  and g2636 (n1784, n_924, n1698);
  not g2637 (n_925, n1784);
  and g2638 (n1785, n_854, n_925);
  not g2639 (n_926, n1783);
  and g2640 (n1786, n_926, n1785);
  not g2641 (n_927, n1786);
  and g2642 (n1787, n_921, n_927);
  and g2643 (n1788, n1643, n_811);
  and g2644 (n1789, n_810, n1647);
  not g2645 (n_928, n1788);
  not g2646 (n_929, n1789);
  and g2647 (n1790, n_928, n_929);
  not g2648 (n_930, n1787);
  and g2649 (n1791, n_930, n1790);
  not g2650 (n_931, n1790);
  and g2651 (n1792, n1787, n_931);
  not g2652 (n_932, n1791);
  not g2653 (n_933, n1792);
  and g2654 (n1793, n_932, n_933);
  and g2655 (n1794, n_882, n_884);
  and g2656 (n1795, n_883, n_884);
  not g2657 (n_934, n1794);
  not g2658 (n_935, n1795);
  and g2659 (n1796, n_934, n_935);
  not g2660 (n_936, n1793);
  not g2661 (n_937, n1796);
  and g2662 (n1797, n_936, n_937);
  and g2663 (n1798, n_930, n_931);
  not g2664 (n_938, n1797);
  not g2665 (n_939, n1798);
  and g2666 (n1799, n_938, n_939);
  not g2667 (n_940, n1744);
  and g2668 (n1800, n1742, n_940);
  not g2669 (n_941, n1800);
  and g2670 (n1801, n_894, n_941);
  not g2671 (n_942, n1799);
  and g2672 (n1802, n_942, n1801);
  and g2673 (n1803, n_272, n1550);
  and g2674 (n1804, n669, n1549);
  and g2675 (n1805, n840, n_456);
  not g2676 (n_943, n1805);
  and g2677 (n1806, n1487, n_943);
  not g2678 (n_944, n1804);
  not g2679 (n_945, n1806);
  and g2680 (n1807, n_944, n_945);
  not g2681 (n_946, n1803);
  and g2682 (n1808, n_946, n1807);
  and g2683 (n1809, n_329, n1368);
  and g2684 (n1810, n832, n1317);
  and g2685 (n1811, n1021, n1371);
  and g2686 (n1812, n_404, n1315);
  and g2694 (n1816, n1808, n1815);
  and g2695 (n1817, n_395, n1241);
  and g2696 (n1818, n1013, n1199);
  and g2697 (n1819, n1183, n1244);
  and g2698 (n1820, n_464, n1197);
  not g2706 (n_955, n1815);
  and g2707 (n1824, n1808, n_955);
  not g2708 (n_956, n1808);
  and g2709 (n1825, n_956, n1815);
  not g2710 (n_957, n1824);
  not g2711 (n_958, n1825);
  and g2712 (n1826, n_957, n_958);
  not g2713 (n_959, n1826);
  and g2714 (n1827, n1823, n_959);
  not g2715 (n_960, n1816);
  not g2716 (n_961, n1827);
  and g2717 (n1828, n_960, n_961);
  and g2718 (n1829, n_159, n844);
  and g2719 (n1830, n279, n700);
  and g2720 (n1831, n286, n847);
  and g2721 (n1832, n_172, n698);
  not g2729 (n_966, n1675);
  not g2730 (n_967, n1680);
  and g2731 (n1836, n_966, n_967);
  not g2732 (n_968, n1836);
  and g2733 (n1837, n_924, n_968);
  not g2734 (n_969, n1837);
  and g2735 (n1838, n1835, n_969);
  not g2736 (n_970, n1835);
  and g2737 (n1839, n_970, n1837);
  not g2738 (n_971, n1838);
  not g2739 (n_972, n1839);
  and g2740 (n1840, n_971, n_972);
  not g2741 (n_973, n1828);
  not g2742 (n_974, n1840);
  and g2743 (n1841, n_973, n_974);
  and g2744 (n1842, n1835, n1837);
  not g2745 (n_975, n1841);
  not g2746 (n_976, n1842);
  and g2747 (n1843, n_975, n_976);
  and g2748 (n1844, n1708, n_873);
  and g2749 (n1845, n_872, n_873);
  not g2750 (n_977, n1844);
  not g2751 (n_978, n1845);
  and g2752 (n1846, n_977, n_978);
  not g2753 (n_979, n1843);
  not g2754 (n_980, n1846);
  and g2755 (n1847, n_979, n_980);
  and g2756 (n1848, n_926, n_927);
  and g2757 (n1849, n1785, n_927);
  not g2758 (n_981, n1848);
  not g2759 (n_982, n1849);
  and g2760 (n1850, n_981, n_982);
  not g2761 (n_983, n1847);
  and g2762 (n1851, n_979, n_983);
  and g2763 (n1852, n_980, n_983);
  not g2764 (n_984, n1851);
  not g2765 (n_985, n1852);
  and g2766 (n1853, n_984, n_985);
  not g2767 (n_986, n1850);
  not g2768 (n_987, n1853);
  and g2769 (n1854, n_986, n_987);
  not g2770 (n_988, n1854);
  and g2771 (n1855, n_983, n_988);
  and g2772 (n1856, n_160, n1033);
  and g2773 (n1857, n275, n868);
  and g2774 (n1858, n279, n1036);
  and g2775 (n1859, n_159, n866);
  and g2783 (n1863, n_338, n1550);
  and g2784 (n1864, n840, n1549);
  and g2785 (n1865, n832, n_456);
  not g2786 (n_993, n1865);
  and g2787 (n1866, n1487, n_993);
  not g2788 (n_994, n1864);
  not g2789 (n_995, n1866);
  and g2790 (n1867, n_994, n_995);
  not g2791 (n_996, n1863);
  and g2792 (n1868, n_996, n1867);
  and g2793 (n1869, n_172, n1033);
  and g2794 (n1870, n286, n_330);
  not g2795 (n_997, n1036);
  not g2796 (n_998, n1870);
  and g2797 (n1871, n_997, n_998);
  not g2798 (n_999, n1869);
  and g2799 (n1872, n_999, n1871);
  and g2800 (n1873, n828, n1872);
  and g2801 (n1874, n1868, n1873);
  and g2802 (n1875, n1862, n1874);
  not g2803 (n_1000, n1862);
  and g2804 (n1876, n_1000, n1874);
  not g2805 (n_1001, n1874);
  and g2806 (n1877, n1862, n_1001);
  not g2807 (n_1002, n1876);
  not g2808 (n_1003, n1877);
  and g2809 (n1878, n_1002, n_1003);
  and g2810 (n1879, n_172, n_295);
  not g2811 (n_1004, n1878);
  and g2812 (n1880, n_1004, n1879);
  not g2813 (n_1005, n1875);
  not g2814 (n_1006, n1880);
  and g2815 (n1881, n_1005, n_1006);
  not g2816 (n_1007, n1757);
  and g2817 (n1882, n_1007, n1774);
  not g2818 (n_1008, n1882);
  and g2819 (n1883, n_917, n_1008);
  not g2820 (n_1009, n1881);
  and g2821 (n1884, n_1009, n1883);
  not g2822 (n_1010, n1883);
  and g2823 (n1885, n1881, n_1010);
  not g2824 (n_1011, n1884);
  not g2825 (n_1012, n1885);
  and g2826 (n1886, n_1011, n_1012);
  and g2827 (n1887, n1828, n1840);
  not g2828 (n_1013, n1887);
  and g2829 (n1888, n_975, n_1013);
  not g2830 (n_1014, n1886);
  not g2831 (n_1015, n1888);
  and g2832 (n1889, n_1014, n_1015);
  and g2833 (n1890, n1886, n1888);
  and g2834 (n1891, n_159, n1033);
  and g2835 (n1892, n279, n868);
  and g2836 (n1893, n286, n1036);
  and g2837 (n1894, n_172, n866);
  and g2845 (n1898, n_404, n1368);
  and g2846 (n1899, n1021, n1317);
  and g2847 (n1900, n1013, n1371);
  and g2848 (n1901, n_395, n1315);
  and g2856 (n1905, n_464, n1241);
  and g2857 (n1906, n1183, n1199);
  and g2858 (n1907, n275, n1244);
  and g2859 (n1908, n_160, n1197);
  not g2867 (n_1028, n1911);
  and g2868 (n1912, n1904, n_1028);
  not g2869 (n_1029, n1904);
  and g2870 (n1913, n_1029, n1911);
  not g2871 (n_1030, n1912);
  not g2872 (n_1031, n1913);
  and g2873 (n1914, n_1030, n_1031);
  not g2874 (n_1032, n1914);
  and g2875 (n1915, n1897, n_1032);
  and g2876 (n1916, n1904, n1911);
  not g2877 (n_1033, n1915);
  not g2878 (n_1034, n1916);
  and g2879 (n1917, n_1033, n_1034);
  not g2880 (n_1035, n1823);
  and g2881 (n1918, n_1035, n1826);
  not g2882 (n_1036, n1918);
  and g2883 (n1919, n_961, n_1036);
  not g2884 (n_1037, n1917);
  and g2885 (n1920, n_1037, n1919);
  not g2886 (n_1038, n1879);
  and g2887 (n1921, n1878, n_1038);
  not g2888 (n_1039, n1921);
  and g2889 (n1922, n_1006, n_1039);
  not g2890 (n_1040, n1920);
  and g2891 (n1923, n_1037, n_1040);
  and g2892 (n1924, n1919, n_1040);
  not g2893 (n_1041, n1923);
  not g2894 (n_1042, n1924);
  and g2895 (n1925, n_1041, n_1042);
  not g2896 (n_1043, n1925);
  and g2897 (n1926, n1922, n_1043);
  not g2898 (n_1044, n1926);
  and g2899 (n1927, n_1040, n_1044);
  not g2900 (n_1045, n1872);
  and g2901 (n1928, n_330, n_1045);
  and g2902 (n1929, n_404, n1550);
  and g2903 (n1930, n1021, n1549);
  and g2904 (n1931, n1013, n_456);
  not g2905 (n_1046, n1931);
  and g2906 (n1932, n1487, n_1046);
  not g2907 (n_1047, n1930);
  not g2908 (n_1048, n1932);
  and g2909 (n1933, n_1047, n_1048);
  not g2910 (n_1049, n1929);
  and g2911 (n1934, n_1049, n1933);
  and g2912 (n1935, n_172, n1241);
  and g2913 (n1936, n286, n_396);
  and g2920 (n1940, n1934, n1939);
  not g2921 (n_1053, n1873);
  and g2922 (n1941, n_1053, n1940);
  not g2923 (n_1054, n1928);
  and g2924 (n1942, n_1054, n1941);
  and g2925 (n1943, n_464, n1368);
  and g2926 (n1944, n1183, n1317);
  and g2927 (n1945, n275, n1371);
  and g2928 (n1946, n_160, n1315);
  and g2936 (n1950, n_159, n1241);
  and g2937 (n1951, n279, n1199);
  and g2938 (n1952, n286, n1244);
  and g2939 (n1953, n_172, n1197);
  and g2947 (n1957, n1949, n1956);
  not g2948 (n_1063, n1934);
  not g2949 (n_1064, n1939);
  and g2950 (n1958, n_1063, n_1064);
  not g2951 (n_1065, n1940);
  not g2952 (n_1066, n1958);
  and g2953 (n1959, n_1065, n_1066);
  not g2954 (n_1067, n1949);
  not g2955 (n_1068, n1956);
  and g2956 (n1960, n_1067, n_1068);
  not g2957 (n_1069, n1957);
  not g2958 (n_1070, n1960);
  and g2959 (n1961, n_1069, n_1070);
  and g2960 (n1962, n1959, n1961);
  not g2961 (n_1071, n1962);
  and g2962 (n1963, n_1069, n_1071);
  not g2963 (n_1072, n1942);
  and g2964 (n1964, n1940, n_1072);
  and g2965 (n1965, n_1053, n_1072);
  and g2966 (n1966, n_1054, n1965);
  not g2967 (n_1073, n1964);
  not g2968 (n_1074, n1966);
  and g2969 (n1967, n_1073, n_1074);
  not g2970 (n_1075, n1963);
  not g2971 (n_1076, n1967);
  and g2972 (n1968, n_1075, n_1076);
  not g2973 (n_1077, n1968);
  and g2974 (n1969, n_1072, n_1077);
  and g2975 (n1970, n_160, n1241);
  and g2976 (n1971, n275, n1199);
  and g2977 (n1972, n279, n1244);
  and g2978 (n1973, n_159, n1197);
  and g2986 (n1977, n_395, n1368);
  and g2987 (n1978, n1013, n1317);
  and g2988 (n1979, n1183, n1371);
  and g2989 (n1980, n_464, n1315);
  and g2997 (n1984, n_329, n1550);
  and g2998 (n1985, n832, n1549);
  and g2999 (n1986, n1021, n_456);
  not g3000 (n_1086, n1986);
  and g3001 (n1987, n1487, n_1086);
  not g3002 (n_1087, n1985);
  not g3003 (n_1088, n1987);
  and g3004 (n1988, n_1087, n_1088);
  not g3005 (n_1089, n1984);
  and g3006 (n1989, n_1089, n1988);
  not g3007 (n_1090, n1983);
  and g3008 (n1990, n_1090, n1989);
  not g3009 (n_1091, n1989);
  and g3010 (n1991, n1983, n_1091);
  not g3011 (n_1092, n1990);
  not g3012 (n_1093, n1991);
  and g3013 (n1992, n_1092, n_1093);
  not g3014 (n_1094, n1976);
  and g3015 (n1993, n_1094, n1992);
  not g3016 (n_1095, n1992);
  and g3017 (n1994, n1976, n_1095);
  and g3018 (n1995, n_395, n1550);
  and g3019 (n1996, n1013, n1549);
  and g3020 (n1997, n_456, n1183);
  not g3021 (n_1096, n1997);
  and g3022 (n1998, n1487, n_1096);
  not g3023 (n_1097, n1996);
  not g3024 (n_1098, n1998);
  and g3025 (n1999, n_1097, n_1098);
  not g3026 (n_1099, n1995);
  and g3027 (n2000, n_1099, n1999);
  and g3028 (n2001, n_160, n1368);
  and g3029 (n2002, n275, n1317);
  and g3030 (n2003, n279, n1371);
  and g3031 (n2004, n_159, n1315);
  not g3039 (n_1104, n2007);
  and g3040 (n2008, n2000, n_1104);
  not g3041 (n_1105, n2000);
  and g3042 (n2009, n_1105, n2007);
  not g3043 (n_1106, n2008);
  not g3044 (n_1107, n2009);
  and g3045 (n2010, n_1106, n_1107);
  and g3046 (n2011, n_464, n1550);
  and g3047 (n2012, n1183, n1549);
  and g3048 (n2013, n275, n_456);
  not g3049 (n_1108, n2013);
  and g3050 (n2014, n1487, n_1108);
  not g3051 (n_1109, n2012);
  not g3052 (n_1110, n2014);
  and g3053 (n2015, n_1109, n_1110);
  not g3054 (n_1111, n2011);
  and g3055 (n2016, n_1111, n2015);
  and g3056 (n2017, n_172, n1368);
  and g3057 (n2018, n286, n_459);
  not g3058 (n_1112, n1371);
  not g3059 (n_1113, n2018);
  and g3060 (n2019, n_1112, n_1113);
  not g3061 (n_1114, n2017);
  and g3062 (n2020, n_1114, n2019);
  and g3063 (n2021, n1177, n2020);
  and g3064 (n2022, n2016, n2021);
  not g3065 (n_1115, n2022);
  and g3066 (n2023, n2010, n_1115);
  not g3067 (n_1116, n2010);
  and g3068 (n2024, n_1116, n2022);
  and g3069 (n2025, n_159, n1368);
  and g3070 (n2026, n279, n1317);
  and g3071 (n2027, n_172, n1315);
  not g3072 (n_1117, n2020);
  and g3073 (n2028, n_459, n_1117);
  and g3074 (n2029, n_160, n1550);
  and g3075 (n2030, n275, n1549);
  and g3076 (n2031, n_159, n_732);
  and g3077 (n2032, n1130, n1487);
  not g3078 (n_1118, n2032);
  and g3079 (n2033, n279, n_1118);
  not g3080 (n_1119, n2031);
  not g3081 (n_1120, n2033);
  and g3082 (n2034, n_1119, n_1120);
  not g3083 (n_1121, n2030);
  not g3084 (n_1122, n2034);
  and g3085 (n2035, n_1121, n_1122);
  not g3086 (n_1123, n2029);
  and g3087 (n2036, n_1123, n2035);
  and g3088 (n2037, n286, n_456);
  and g3089 (n2038, n_1119, n2037);
  not g3090 (n_1124, n2036);
  not g3091 (n_1125, n2038);
  and g3092 (n2039, n_1124, n_1125);
  not g3093 (n_1126, n2021);
  not g3094 (n_1127, n2039);
  and g3095 (n2040, n_1126, n_1127);
  not g3096 (n_1128, n2028);
  and g3097 (n2041, n_1128, n2040);
  and g3098 (n2042, n2036, n2038);
  not g3099 (n_1129, n2041);
  not g3100 (n_1130, n2042);
  and g3101 (n2043, n_1129, n_1130);
  not g3102 (n_1131, n2016);
  and g3103 (n2044, n_1131, n_1126);
  not g3104 (n_1132, n2044);
  and g3105 (n2045, n_1115, n_1132);
  not g3106 (n_1133, n2045);
  and g3107 (n2046, n2043, n_1133);
  and g3108 (n2047, n286, n1371);
  not g3118 (n_1139, n2043);
  and g3119 (n2052, n_1139, n2045);
  not g3120 (n_1140, n2051);
  not g3121 (n_1141, n2052);
  and g3122 (n2053, n_1140, n_1141);
  and g3123 (n2054, n_172, n_478);
  not g3124 (n_1142, n2054);
  and g3125 (n2055, n2053, n_1142);
  not g3126 (n_1143, n2024);
  not g3127 (n_1144, n2055);
  and g3128 (n2056, n_1143, n_1144);
  not g3129 (n_1145, n2023);
  and g3130 (n2057, n_1145, n2056);
  not g3131 (n_1146, n2053);
  and g3132 (n2058, n_1146, n2054);
  not g3133 (n_1147, n2057);
  not g3134 (n_1148, n2058);
  and g3135 (n2059, n_1147, n_1148);
  and g3136 (n2060, n1959, n_1071);
  and g3137 (n2061, n_1070, n1963);
  not g3138 (n_1149, n2060);
  not g3139 (n_1150, n2061);
  and g3140 (n2062, n_1149, n_1150);
  and g3141 (n2063, n2059, n2062);
  and g3142 (n2064, n2000, n2007);
  not g3143 (n_1151, n2064);
  and g3144 (n2065, n_1143, n_1151);
  not g3145 (n_1152, n2063);
  not g3146 (n_1153, n2065);
  and g3147 (n2066, n_1152, n_1153);
  not g3148 (n_1154, n2059);
  not g3149 (n_1155, n2062);
  and g3150 (n2067, n_1154, n_1155);
  not g3151 (n_1156, n2066);
  not g3152 (n_1157, n2067);
  and g3153 (n2068, n_1156, n_1157);
  and g3154 (n2069, n_1075, n_1077);
  and g3155 (n2070, n_1076, n_1077);
  not g3156 (n_1158, n2069);
  not g3157 (n_1159, n2070);
  and g3158 (n2071, n_1158, n_1159);
  and g3159 (n2072, n2068, n2071);
  not g3160 (n_1160, n1994);
  not g3161 (n_1161, n2072);
  and g3162 (n2073, n_1160, n_1161);
  not g3163 (n_1162, n1993);
  and g3164 (n2074, n_1162, n2073);
  not g3165 (n_1163, n2068);
  not g3166 (n_1164, n2071);
  and g3167 (n2075, n_1163, n_1164);
  not g3168 (n_1165, n2074);
  not g3169 (n_1166, n2075);
  and g3170 (n2076, n_1165, n_1166);
  not g3171 (n_1167, n1969);
  not g3172 (n_1168, n2076);
  and g3173 (n2077, n_1167, n_1168);
  and g3174 (n2078, n1969, n2076);
  and g3175 (n2079, n1897, n_1033);
  and g3176 (n2080, n_1032, n_1033);
  not g3177 (n_1169, n2079);
  not g3178 (n_1170, n2080);
  and g3179 (n2081, n_1169, n_1170);
  not g3180 (n_1171, n1868);
  and g3181 (n2082, n_1171, n_1053);
  not g3182 (n_1172, n2082);
  and g3183 (n2083, n_1001, n_1172);
  and g3184 (n2084, n1983, n1989);
  not g3185 (n_1173, n2084);
  and g3186 (n2085, n_1160, n_1173);
  not g3187 (n_1174, n2085);
  and g3188 (n2086, n2083, n_1174);
  not g3189 (n_1175, n2083);
  and g3190 (n2087, n_1175, n2085);
  not g3191 (n_1176, n2086);
  not g3192 (n_1177, n2087);
  and g3193 (n2088, n_1176, n_1177);
  not g3194 (n_1178, n2081);
  and g3195 (n2089, n_1178, n2088);
  not g3196 (n_1179, n2088);
  and g3197 (n2090, n2081, n_1179);
  not g3198 (n_1180, n2089);
  not g3199 (n_1181, n2090);
  and g3200 (n2091, n_1180, n_1181);
  not g3201 (n_1182, n2078);
  and g3202 (n2092, n_1182, n2091);
  not g3203 (n_1183, n2077);
  not g3204 (n_1184, n2092);
  and g3205 (n2093, n_1183, n_1184);
  and g3206 (n2094, n_1176, n_1180);
  not g3207 (n_1185, n2093);
  not g3208 (n_1186, n2094);
  and g3209 (n2095, n_1185, n_1186);
  and g3210 (n2096, n2093, n2094);
  not g3211 (n_1187, n1922);
  and g3212 (n2097, n_1187, n1925);
  not g3213 (n_1188, n2097);
  and g3214 (n2098, n_1044, n_1188);
  not g3215 (n_1189, n2096);
  and g3216 (n2099, n_1189, n2098);
  not g3217 (n_1190, n2095);
  not g3218 (n_1191, n2099);
  and g3219 (n2100, n_1190, n_1191);
  and g3220 (n2101, n1927, n2100);
  not g3221 (n_1192, n1890);
  not g3222 (n_1193, n2101);
  and g3223 (n2102, n_1192, n_1193);
  not g3224 (n_1194, n1889);
  and g3225 (n2103, n_1194, n2102);
  not g3226 (n_1195, n1927);
  not g3227 (n_1196, n2100);
  and g3228 (n2104, n_1195, n_1196);
  not g3229 (n_1197, n2103);
  not g3230 (n_1198, n2104);
  and g3231 (n2105, n_1197, n_1198);
  and g3232 (n2106, n_1011, n_1192);
  not g3233 (n_1199, n2105);
  not g3234 (n_1200, n2106);
  and g3235 (n2107, n_1199, n_1200);
  and g3236 (n2108, n2105, n2106);
  and g3237 (n2109, n1850, n1853);
  not g3238 (n_1201, n2109);
  and g3239 (n2110, n_988, n_1201);
  not g3240 (n_1202, n2108);
  and g3241 (n2111, n_1202, n2110);
  not g3242 (n_1203, n2107);
  not g3243 (n_1204, n2111);
  and g3244 (n2112, n_1203, n_1204);
  and g3245 (n2113, n1855, n2112);
  and g3246 (n2114, n1793, n1796);
  not g3247 (n_1205, n2113);
  not g3248 (n_1206, n2114);
  and g3249 (n2115, n_1205, n_1206);
  and g3250 (n2116, n_938, n2115);
  not g3251 (n_1207, n1855);
  not g3252 (n_1208, n2112);
  and g3253 (n2117, n_1207, n_1208);
  not g3254 (n_1209, n2116);
  not g3255 (n_1210, n2117);
  and g3256 (n2118, n_1209, n_1210);
  not g3257 (n_1211, n1801);
  and g3258 (n2119, n1799, n_1211);
  not g3259 (n_1212, n1802);
  not g3260 (n_1213, n2119);
  and g3261 (n2120, n_1212, n_1213);
  not g3262 (n_1214, n2118);
  and g3263 (n2121, n_1214, n2120);
  not g3264 (n_1215, n2121);
  and g3265 (n2122, n_1212, n_1215);
  not g3266 (n_1216, n1748);
  and g3267 (n2123, n1746, n_1216);
  not g3268 (n_1217, n1749);
  not g3269 (n_1218, n2123);
  and g3270 (n2124, n_1217, n_1218);
  not g3271 (n_1219, n2122);
  and g3272 (n2125, n_1219, n2124);
  not g3273 (n_1220, n2125);
  and g3274 (n2126, n_1217, n_1220);
  not g3275 (n_1221, n1668);
  and g3276 (n2127, n1666, n_1221);
  not g3277 (n_1222, n1669);
  not g3278 (n_1223, n2127);
  and g3279 (n2128, n_1222, n_1223);
  not g3280 (n_1224, n2126);
  and g3281 (n2129, n_1224, n2128);
  not g3282 (n_1225, n2129);
  and g3283 (n2130, n_1222, n_1225);
  not g3284 (n_1226, n1625);
  and g3285 (n2131, n1623, n_1226);
  not g3286 (n_1227, n1626);
  not g3287 (n_1228, n2131);
  and g3288 (n2132, n_1227, n_1228);
  not g3289 (n_1229, n2130);
  and g3290 (n2133, n_1229, n2132);
  not g3291 (n_1230, n2133);
  and g3292 (n2134, n_1227, n_1230);
  not g3293 (n_1231, n1548);
  not g3294 (n_1232, n2134);
  and g3295 (n2135, n_1231, n_1232);
  not g3296 (n_1233, n1545);
  not g3297 (n_1234, n2135);
  and g3298 (n2136, n_1233, n_1234);
  and g3299 (n2137, n1424, n1427);
  not g3300 (n_1235, n1428);
  not g3301 (n_1236, n2137);
  and g3302 (n2138, n_1235, n_1236);
  not g3303 (n_1237, n2136);
  and g3304 (n2139, n_1237, n2138);
  not g3305 (n_1238, n2139);
  and g3306 (n2140, n_1235, n_1238);
  not g3307 (n_1239, n1295);
  not g3308 (n_1240, n2140);
  and g3309 (n2141, n_1239, n_1240);
  not g3310 (n_1241, n2141);
  and g3311 (n2142, n_561, n_1241);
  not g3312 (n_1242, n1236);
  and g3313 (n2143, n1234, n_1242);
  not g3314 (n_1243, n1237);
  not g3315 (n_1244, n2143);
  and g3316 (n2144, n_1243, n_1244);
  not g3317 (n_1245, n2142);
  and g3318 (n2145, n_1245, n2144);
  not g3319 (n_1246, n2145);
  and g3320 (n2146, n_1243, n_1246);
  not g3321 (n_1247, n1074);
  not g3322 (n_1248, n2146);
  and g3323 (n2147, n_1247, n_1248);
  and g3324 (n2148, n_444, n_445);
  not g3325 (n_1249, n2147);
  not g3326 (n_1250, n2148);
  and g3327 (n2149, n_1249, n_1250);
  not g3328 (n_1251, n897);
  and g3329 (n2150, n895, n_1251);
  not g3330 (n_1252, n898);
  not g3331 (n_1253, n2150);
  and g3332 (n2151, n_1252, n_1253);
  not g3333 (n_1254, n2149);
  and g3334 (n2152, n_1254, n2151);
  not g3335 (n_1255, n2152);
  and g3336 (n2153, n_1252, n_1255);
  not g3337 (n_1256, n728);
  not g3338 (n_1257, n2153);
  and g3339 (n2154, n_1256, n_1257);
  and g3340 (n2155, n_317, n_318);
  not g3341 (n_1258, n2154);
  not g3342 (n_1259, n2155);
  and g3343 (n2156, n_1258, n_1259);
  not g3344 (n_1260, n2156);
  and g3345 (n2157, n683, n_1260);
  not g3346 (n_1261, n683);
  and g3347 (n2158, n_1261, n2156);
  not g3348 (n_1262, n2157);
  not g3349 (n_1263, n2158);
  and g3350 (n2159, n_1262, n_1263);
  and g3351 (n2160, n536, n2159);
  not g3352 (n_1264, n536);
  not g3353 (n_1265, n2159);
  and g3354 (n2161, n_1264, n_1265);
  not g3355 (n_1266, n2160);
  not g3356 (n_1267, n2161);
  and g3357 (n2162, n_1266, n_1267);
  not g3358 (n_1268, n393);
  not g3359 (n_1269, n2162);
  and g3360 (n2163, n_1268, n_1269);
  and g3361 (n2164, n393, n2162);
  and g3362 (n2165, n_95, n_224);
  and g3363 (n2166, n_131, n2165);
  and g3379 (n2182, n_201, n968);
  and g3380 (n2183, n_85, n2182);
  and g3407 (n2210, n728, n2153);
  not g3408 (n_1270, n2210);
  and g3409 (n2211, n_1258, n_1270);
  not g3410 (n_1271, n2209);
  not g3411 (n_1272, n2211);
  and g3412 (n2212, n_1271, n_1272);
  not g3426 (n_1273, n2151);
  and g3427 (n2226, n2149, n_1273);
  not g3428 (n_1274, n2226);
  and g3429 (n2227, n_1255, n_1274);
  not g3430 (n_1275, n2225);
  not g3431 (n_1276, n2227);
  and g3432 (n2228, n_1275, n_1276);
  and g3433 (n2229, n2225, n2227);
  and g3455 (n2251, n_99, n_228);
  and g3456 (n2252, n_221, n2251);
  and g3457 (n2253, n_177, n_182);
  and g3458 (n2254, n_225, n2253);
  and g3469 (n2265, n1074, n2146);
  not g3470 (n_1277, n2265);
  and g3471 (n2266, n_1249, n_1277);
  not g3472 (n_1278, n2264);
  not g3473 (n_1279, n2266);
  and g3474 (n2267, n_1278, n_1279);
  and g3484 (n2277, n_215, n_263);
  and g3485 (n2278, n_126, n2277);
  not g3500 (n_1280, n2144);
  and g3501 (n2293, n2142, n_1280);
  not g3502 (n_1281, n2293);
  and g3503 (n2294, n_1246, n_1281);
  not g3504 (n_1282, n2292);
  not g3505 (n_1283, n2294);
  and g3506 (n2295, n_1282, n_1283);
  and g3507 (n2296, n2292, n2294);
  and g3523 (n2312, n_150, n923);
  and g3524 (n2313, n_190, n2312);
  and g3539 (n2328, n1295, n2140);
  not g3540 (n_1284, n2328);
  and g3541 (n2329, n_1241, n_1284);
  not g3542 (n_1285, n2327);
  not g3543 (n_1286, n2329);
  and g3544 (n2330, n_1285, n_1286);
  and g3554 (n2340, n_93, n_87);
  and g3555 (n2341, n_150, n_198);
  and g3556 (n2342, n_127, n2341);
  not g3569 (n_1287, n2138);
  and g3570 (n2355, n2136, n_1287);
  not g3571 (n_1288, n2355);
  and g3572 (n2356, n_1238, n_1288);
  not g3573 (n_1289, n2354);
  not g3574 (n_1290, n2356);
  and g3575 (n2357, n_1289, n_1290);
  and g3576 (n2358, n2354, n2356);
  and g3583 (n2365, n_141, n_216);
  and g3584 (n2366, n_260, n2365);
  and g3585 (n2367, n_108, n_126);
  and g3604 (n2386, n1548, n2134);
  not g3605 (n_1291, n2386);
  and g3606 (n2387, n_1234, n_1291);
  not g3607 (n_1292, n2385);
  not g3608 (n_1293, n2387);
  and g3609 (n2388, n_1292, n_1293);
  not g3636 (n_1294, n2132);
  and g3637 (n2415, n2130, n_1294);
  not g3638 (n_1295, n2415);
  and g3639 (n2416, n_1230, n_1295);
  not g3640 (n_1296, n2414);
  not g3641 (n_1297, n2416);
  and g3642 (n2417, n_1296, n_1297);
  and g3643 (n2418, n_261, n_264);
  and g3647 (n2422, n_181, n_216);
  and g3658 (n2433, n_199, n_227);
  not g3672 (n_1298, n2128);
  and g3673 (n2447, n2126, n_1298);
  not g3674 (n_1299, n2447);
  and g3675 (n2448, n_1225, n_1299);
  not g3676 (n_1300, n2446);
  not g3677 (n_1301, n2448);
  and g3678 (n2449, n_1300, n_1301);
  and g3679 (n2450, n2446, n2448);
  not g3707 (n_1302, n2124);
  and g3708 (n2478, n2122, n_1302);
  not g3709 (n_1303, n2478);
  and g3710 (n2479, n_1220, n_1303);
  not g3711 (n_1304, n2477);
  not g3712 (n_1305, n2479);
  and g3713 (n2480, n_1304, n_1305);
  and g3714 (n2481, n2477, n2479);
  and g3715 (n2482, n_1214, n_1215);
  and g3716 (n2483, n2120, n_1215);
  not g3717 (n_1306, n2482);
  not g3718 (n_1307, n2483);
  and g3719 (n2484, n_1306, n_1307);
  not g3731 (n_1308, n2484);
  and g3732 (n2496, n_1308, n2495);
  not g3733 (n_1309, n2480);
  not g3734 (n_1310, n2496);
  and g3735 (n2497, n_1309, n_1310);
  not g3736 (n_1311, n2481);
  and g3737 (n2498, n_1311, n2497);
  not g3738 (n_1312, n2498);
  and g3739 (n2499, n_1309, n_1312);
  not g3740 (n_1313, n2449);
  not g3741 (n_1314, n2499);
  and g3742 (n2500, n_1313, n_1314);
  not g3743 (n_1315, n2450);
  and g3744 (n2501, n_1315, n2500);
  not g3745 (n_1316, n2501);
  and g3746 (n2502, n_1313, n_1316);
  and g3747 (n2503, n2414, n2416);
  not g3748 (n_1317, n2417);
  not g3749 (n_1318, n2503);
  and g3750 (n2504, n_1317, n_1318);
  not g3751 (n_1319, n2502);
  and g3752 (n2505, n_1319, n2504);
  not g3753 (n_1320, n2505);
  and g3754 (n2506, n_1317, n_1320);
  and g3755 (n2507, n2385, n2387);
  not g3756 (n_1321, n2388);
  not g3757 (n_1322, n2507);
  and g3758 (n2508, n_1321, n_1322);
  not g3759 (n_1323, n2506);
  and g3760 (n2509, n_1323, n2508);
  not g3761 (n_1324, n2509);
  and g3762 (n2510, n_1321, n_1324);
  not g3763 (n_1325, n2357);
  not g3764 (n_1326, n2510);
  and g3765 (n2511, n_1325, n_1326);
  not g3766 (n_1327, n2358);
  and g3767 (n2512, n_1327, n2511);
  not g3768 (n_1328, n2512);
  and g3769 (n2513, n_1325, n_1328);
  not g3770 (n_1329, n2330);
  and g3771 (n2514, n_1285, n_1329);
  and g3772 (n2515, n_1286, n_1329);
  not g3773 (n_1330, n2514);
  not g3774 (n_1331, n2515);
  and g3775 (n2516, n_1330, n_1331);
  not g3776 (n_1332, n2513);
  not g3777 (n_1333, n2516);
  and g3778 (n2517, n_1332, n_1333);
  not g3779 (n_1334, n2517);
  and g3780 (n2518, n_1329, n_1334);
  not g3781 (n_1335, n2295);
  not g3782 (n_1336, n2518);
  and g3783 (n2519, n_1335, n_1336);
  not g3784 (n_1337, n2296);
  and g3785 (n2520, n_1337, n2519);
  not g3786 (n_1338, n2520);
  and g3787 (n2521, n_1335, n_1338);
  and g3788 (n2522, n2264, n2266);
  not g3789 (n_1339, n2267);
  not g3790 (n_1340, n2522);
  and g3791 (n2523, n_1339, n_1340);
  not g3792 (n_1341, n2521);
  and g3793 (n2524, n_1341, n2523);
  not g3794 (n_1342, n2524);
  and g3795 (n2525, n_1339, n_1342);
  not g3796 (n_1343, n2228);
  not g3797 (n_1344, n2525);
  and g3798 (n2526, n_1343, n_1344);
  not g3799 (n_1345, n2229);
  and g3800 (n2527, n_1345, n2526);
  not g3801 (n_1346, n2527);
  and g3802 (n2528, n_1343, n_1346);
  and g3803 (n2529, n2209, n2211);
  not g3804 (n_1347, n2212);
  not g3805 (n_1348, n2529);
  and g3806 (n2530, n_1347, n_1348);
  not g3807 (n_1349, n2528);
  and g3808 (n2531, n_1349, n2530);
  not g3809 (n_1350, n2531);
  and g3810 (n2532, n_1347, n_1350);
  not g3811 (n_1351, n2163);
  not g3812 (n_1352, n2532);
  and g3813 (n2533, n_1351, n_1352);
  not g3814 (n_1353, n2164);
  and g3815 (n2534, n_1353, n2533);
  not g3816 (n_1354, n2534);
  and g3817 (n2535, n_1351, n_1354);
  and g3834 (n2552, n2535, n2551);
  not g3835 (n_1355, n2535);
  not g3836 (n_1356, n2551);
  and g3837 (n2553, n_1355, n_1356);
  not g3838 (n_1357, n2552);
  not g3839 (n_1358, n2553);
  and g3840 (n2554, n_1357, n_1358);
  not g3841 (n_1359, n2554);
  and g3842 (n2555, n295, n_1359);
  and g3843 (n2556, n_159, n286);
  and g3844 (n2557, n279, n_172);
  not g3845 (n_1360, n2556);
  not g3846 (n_1361, n2557);
  and g3847 (n2558, n_1360, n_1361);
  not g3848 (n_1362, n282);
  and g3849 (n2559, n_1362, n294);
  and g3850 (n2560, n2558, n2559);
  not g3851 (n_1363, n2530);
  and g3852 (n2561, n2528, n_1363);
  not g3853 (n_1364, n2561);
  and g3854 (n2562, n_1350, n_1364);
  and g3855 (n2563, n2560, n2562);
  and g3856 (n2564, n_1352, n_1354);
  and g3857 (n2565, n_1353, n2535);
  not g3858 (n_1365, n2564);
  not g3859 (n_1366, n2565);
  and g3860 (n2566, n_1365, n_1366);
  not g3861 (n_1367, n2558);
  and g3862 (n2567, n294, n_1367);
  not g3863 (n_1368, n2566);
  and g3864 (n2568, n_1368, n2567);
  and g3870 (n2571, n_1362, n_175);
  and g3871 (n2572, n2562, n_1368);
  and g3872 (n2573, n_1344, n_1346);
  and g3873 (n2574, n_1345, n2528);
  not g3874 (n_1372, n2573);
  not g3875 (n_1373, n2574);
  and g3876 (n2575, n_1372, n_1373);
  not g3877 (n_1374, n2575);
  and g3878 (n2576, n2562, n_1374);
  not g3879 (n_1375, n2523);
  and g3880 (n2577, n2521, n_1375);
  not g3881 (n_1376, n2577);
  and g3882 (n2578, n_1342, n_1376);
  and g3883 (n2579, n_1374, n2578);
  and g3884 (n2580, n_1336, n_1338);
  and g3885 (n2581, n_1337, n2521);
  not g3886 (n_1377, n2580);
  not g3887 (n_1378, n2581);
  and g3888 (n2582, n_1377, n_1378);
  not g3889 (n_1379, n2582);
  and g3890 (n2583, n2578, n_1379);
  and g3891 (n2584, n_1332, n_1334);
  and g3892 (n2585, n_1333, n_1334);
  not g3893 (n_1380, n2584);
  not g3894 (n_1381, n2585);
  and g3895 (n2586, n_1380, n_1381);
  not g3896 (n_1382, n2586);
  and g3897 (n2587, n_1379, n_1382);
  and g3898 (n2588, n_1326, n_1328);
  and g3899 (n2589, n_1327, n2513);
  not g3900 (n_1383, n2588);
  not g3901 (n_1384, n2589);
  and g3902 (n2590, n_1383, n_1384);
  not g3903 (n_1385, n2590);
  and g3904 (n2591, n_1382, n_1385);
  not g3905 (n_1386, n2508);
  and g3906 (n2592, n2506, n_1386);
  not g3907 (n_1387, n2592);
  and g3908 (n2593, n_1324, n_1387);
  and g3909 (n2594, n_1385, n2593);
  not g3910 (n_1388, n2504);
  and g3911 (n2595, n2502, n_1388);
  not g3912 (n_1389, n2595);
  and g3913 (n2596, n_1320, n_1389);
  and g3914 (n2597, n2593, n2596);
  and g3915 (n2598, n_1314, n_1316);
  and g3916 (n2599, n_1315, n2502);
  not g3917 (n_1390, n2598);
  not g3918 (n_1391, n2599);
  and g3919 (n2600, n_1390, n_1391);
  not g3920 (n_1392, n2600);
  and g3921 (n2601, n2596, n_1392);
  and g3922 (n2602, n_1310, n_1312);
  and g3923 (n2603, n_1311, n2499);
  not g3924 (n_1393, n2602);
  not g3925 (n_1394, n2603);
  and g3926 (n2604, n_1393, n_1394);
  not g3927 (n_1395, n2604);
  and g3928 (n2605, n_1392, n_1395);
  not g3929 (n_1396, n2495);
  and g3930 (n2606, n2484, n_1396);
  not g3931 (n_1397, n2606);
  and g3932 (n2607, n_1310, n_1397);
  not g3933 (n_1398, n2607);
  and g3934 (n2608, n_1395, n_1398);
  and g3935 (n2609, n2600, n2608);
  not g3936 (n_1399, n2605);
  not g3937 (n_1400, n2609);
  and g3938 (n2610, n_1399, n_1400);
  not g3939 (n_1401, n2596);
  and g3940 (n2611, n_1401, n2600);
  not g3941 (n_1402, n2610);
  not g3942 (n_1403, n2611);
  and g3943 (n2612, n_1402, n_1403);
  not g3944 (n_1404, n2601);
  and g3945 (n2613, n_1404, n2612);
  not g3946 (n_1405, n2613);
  and g3947 (n2614, n_1404, n_1405);
  not g3948 (n_1406, n2593);
  and g3949 (n2615, n_1406, n_1401);
  not g3950 (n_1407, n2614);
  not g3951 (n_1408, n2615);
  and g3952 (n2616, n_1407, n_1408);
  not g3953 (n_1409, n2597);
  and g3954 (n2617, n_1409, n2616);
  not g3955 (n_1410, n2617);
  and g3956 (n2618, n_1409, n_1410);
  and g3957 (n2619, n2590, n_1406);
  not g3958 (n_1411, n2594);
  not g3959 (n_1412, n2619);
  and g3960 (n2620, n_1411, n_1412);
  not g3961 (n_1413, n2618);
  and g3962 (n2621, n_1413, n2620);
  not g3963 (n_1414, n2621);
  and g3964 (n2622, n_1411, n_1414);
  and g3965 (n2623, n2586, n2590);
  not g3966 (n_1415, n2591);
  not g3967 (n_1416, n2623);
  and g3968 (n2624, n_1415, n_1416);
  not g3969 (n_1417, n2622);
  and g3970 (n2625, n_1417, n2624);
  not g3971 (n_1418, n2625);
  and g3972 (n2626, n_1415, n_1418);
  and g3973 (n2627, n2582, n2586);
  not g3974 (n_1419, n2587);
  not g3975 (n_1420, n2627);
  and g3976 (n2628, n_1419, n_1420);
  not g3977 (n_1421, n2626);
  and g3978 (n2629, n_1421, n2628);
  not g3979 (n_1422, n2629);
  and g3980 (n2630, n_1419, n_1422);
  not g3981 (n_1423, n2578);
  and g3982 (n2631, n_1423, n2582);
  not g3983 (n_1424, n2583);
  not g3984 (n_1425, n2631);
  and g3985 (n2632, n_1424, n_1425);
  not g3986 (n_1426, n2630);
  and g3987 (n2633, n_1426, n2632);
  not g3988 (n_1427, n2633);
  and g3989 (n2634, n_1424, n_1427);
  and g3990 (n2635, n2575, n_1423);
  not g3991 (n_1428, n2579);
  not g3992 (n_1429, n2635);
  and g3993 (n2636, n_1428, n_1429);
  not g3994 (n_1430, n2634);
  and g3995 (n2637, n_1430, n2636);
  not g3996 (n_1431, n2637);
  and g3997 (n2638, n_1428, n_1431);
  not g3998 (n_1432, n2562);
  and g3999 (n2639, n_1432, n2575);
  not g4000 (n_1433, n2576);
  not g4001 (n_1434, n2639);
  and g4002 (n2640, n_1433, n_1434);
  not g4003 (n_1435, n2638);
  and g4004 (n2641, n_1435, n2640);
  not g4005 (n_1436, n2641);
  and g4006 (n2642, n_1433, n_1436);
  and g4007 (n2643, n_1432, n2566);
  not g4008 (n_1437, n2572);
  not g4009 (n_1438, n2643);
  and g4010 (n2644, n_1437, n_1438);
  not g4011 (n_1439, n2642);
  and g4012 (n2645, n_1439, n2644);
  not g4013 (n_1440, n2645);
  and g4014 (n2646, n_1437, n_1440);
  and g4015 (n2647, n_1359, n_1368);
  and g4016 (n2648, n2554, n2566);
  not g4017 (n_1441, n2647);
  not g4018 (n_1442, n2648);
  and g4019 (n2649, n_1441, n_1442);
  not g4020 (n_1443, n2646);
  and g4021 (n2650, n_1443, n2649);
  not g4022 (n_1444, n2649);
  and g4023 (n2651, n2646, n_1444);
  not g4024 (n_1445, n2650);
  not g4025 (n_1446, n2651);
  and g4026 (n2652, n_1445, n_1446);
  and g4027 (n2653, n2571, n2652);
  not g4030 (n_1448, n2654);
  and g4031 (n2655, n_160, n_1448);
  and g4032 (n2656, n275, n2654);
  not g4033 (n_1449, n2655);
  not g4034 (n_1450, n2656);
  and g4035 (n2657, n_1449, n_1450);
  and g4036 (n2658, n669, n_281);
  and g4037 (n2659, n_272, n677);
  not g4038 (n_1451, n2658);
  not g4039 (n_1452, n2659);
  and g4040 (n2660, n_1451, n_1452);
  not g4041 (n_1453, n2660);
  and g4042 (n2661, n_1398, n_1453);
  not g4043 (n_1454, n2661);
  and g4044 (n2662, n_240, n_1454);
  and g4045 (n2663, n529, n_281);
  and g4046 (n2664, n_241, n677);
  not g4047 (n_1455, n2663);
  not g4048 (n_1456, n2664);
  and g4049 (n2665, n_1455, n_1456);
  not g4050 (n_1457, n2665);
  and g4051 (n2666, n2660, n_1457);
  and g4052 (n2667, n_1398, n2666);
  and g4053 (n2668, n532, n_1453);
  and g4054 (n2669, n_1395, n2668);
  not g4055 (n_1458, n2667);
  not g4056 (n_1459, n2669);
  and g4057 (n2670, n_1458, n_1459);
  and g4058 (n2671, n2604, n_1398);
  and g4059 (n2672, n_1395, n2607);
  not g4060 (n_1460, n2671);
  not g4061 (n_1461, n2672);
  and g4062 (n2673, n_1460, n_1461);
  and g4063 (n2674, n_245, n_1453);
  not g4064 (n_1462, n2673);
  and g4065 (n2675, n_1462, n2674);
  not g4066 (n_1463, n2675);
  and g4067 (n2676, n2670, n_1463);
  not g4068 (n_1464, n2676);
  and g4069 (n2677, n_240, n_1464);
  not g4070 (n_1465, n2677);
  and g4071 (n2678, n_240, n_1465);
  and g4072 (n2679, n_1464, n_1465);
  not g4073 (n_1466, n2678);
  not g4074 (n_1467, n2679);
  and g4075 (n2680, n_1466, n_1467);
  not g4076 (n_1468, n2680);
  and g4077 (n2681, n2662, n_1468);
  not g4078 (n_1469, n2662);
  and g4079 (n2682, n_1469, n2680);
  not g4080 (n_1470, n2681);
  not g4081 (n_1471, n2682);
  and g4082 (n2683, n_1470, n_1471);
  and g4083 (n2684, n832, n_404);
  and g4084 (n2685, n_329, n1021);
  not g4085 (n_1472, n2684);
  not g4086 (n_1473, n2685);
  and g4087 (n2686, n_1472, n_1473);
  and g4088 (n2687, n669, n_338);
  and g4089 (n2688, n_272, n840);
  not g4090 (n_1474, n2687);
  not g4091 (n_1475, n2688);
  and g4092 (n2689, n_1474, n_1475);
  not g4093 (n_1476, n2686);
  not g4094 (n_1477, n2689);
  and g4095 (n2690, n_1476, n_1477);
  and g4096 (n2691, n832, n_338);
  and g4097 (n2692, n_329, n840);
  not g4098 (n_1478, n2691);
  not g4099 (n_1479, n2692);
  and g4100 (n2693, n_1478, n_1479);
  and g4101 (n2694, n2686, n_1477);
  and g4102 (n2695, n2693, n2694);
  and g4103 (n2696, n_1392, n2695);
  not g4104 (n_1480, n2693);
  and g4105 (n2697, n2686, n_1480);
  and g4106 (n2698, n2596, n2697);
  and g4107 (n2699, n_1476, n2689);
  and g4108 (n2700, n2593, n2699);
  not g4109 (n_1481, n2698);
  not g4110 (n_1482, n2700);
  and g4111 (n2701, n_1481, n_1482);
  not g4112 (n_1483, n2696);
  and g4113 (n2702, n_1483, n2701);
  not g4114 (n_1484, n2690);
  and g4115 (n2703, n_1484, n2702);
  and g4116 (n2704, n_1407, n_1410);
  and g4117 (n2705, n_1408, n2618);
  not g4118 (n_1485, n2704);
  not g4119 (n_1486, n2705);
  and g4120 (n2706, n_1485, n_1486);
  and g4121 (n2707, n2702, n2706);
  not g4122 (n_1487, n2703);
  not g4123 (n_1488, n2707);
  and g4124 (n2708, n_1487, n_1488);
  not g4125 (n_1489, n2708);
  and g4126 (n2709, n669, n_1489);
  and g4127 (n2710, n_272, n2708);
  not g4128 (n_1490, n2709);
  not g4129 (n_1491, n2710);
  and g4130 (n2711, n_1490, n_1491);
  and g4131 (n2712, n2683, n2711);
  and g4132 (n2713, n_1398, n_1476);
  not g4133 (n_1492, n2713);
  and g4134 (n2714, n_272, n_1492);
  and g4135 (n2715, n_1398, n2697);
  and g4136 (n2716, n_1395, n2699);
  not g4137 (n_1493, n2715);
  not g4138 (n_1494, n2716);
  and g4139 (n2717, n_1493, n_1494);
  and g4140 (n2718, n_1462, n2690);
  not g4141 (n_1495, n2718);
  and g4142 (n2719, n2717, n_1495);
  not g4143 (n_1496, n2719);
  and g4144 (n2720, n_272, n_1496);
  and g4145 (n2721, n669, n2719);
  not g4146 (n_1497, n2720);
  not g4147 (n_1498, n2721);
  and g4148 (n2722, n_1497, n_1498);
  and g4149 (n2723, n2714, n2722);
  and g4150 (n2724, n_1392, n2699);
  and g4151 (n2725, n_1398, n2695);
  and g4152 (n2726, n_1395, n2697);
  not g4153 (n_1499, n2725);
  not g4154 (n_1500, n2726);
  and g4155 (n2727, n_1499, n_1500);
  not g4156 (n_1501, n2724);
  and g4157 (n2728, n_1501, n2727);
  and g4158 (n2729, n_1484, n2728);
  and g4159 (n2730, n2600, n_1461);
  and g4160 (n2731, n_1392, n2672);
  not g4161 (n_1502, n2730);
  not g4162 (n_1503, n2731);
  and g4163 (n2732, n_1502, n_1503);
  not g4164 (n_1504, n2732);
  and g4165 (n2733, n2728, n_1504);
  not g4166 (n_1505, n2729);
  not g4167 (n_1506, n2733);
  and g4168 (n2734, n_1505, n_1506);
  not g4169 (n_1507, n2734);
  and g4170 (n2735, n669, n_1507);
  and g4171 (n2736, n_272, n2734);
  not g4172 (n_1508, n2735);
  not g4173 (n_1509, n2736);
  and g4174 (n2737, n_1508, n_1509);
  and g4175 (n2738, n2723, n2737);
  and g4176 (n2739, n2661, n2738);
  not g4177 (n_1510, n2739);
  and g4178 (n2740, n2738, n_1510);
  and g4179 (n2741, n2661, n_1510);
  not g4180 (n_1511, n2740);
  not g4181 (n_1512, n2741);
  and g4182 (n2742, n_1511, n_1512);
  and g4183 (n2743, n_1392, n2697);
  and g4184 (n2744, n2596, n2699);
  and g4185 (n2745, n_1395, n2695);
  and g4191 (n2748, n_1402, n_1405);
  and g4192 (n2749, n_1403, n2614);
  not g4193 (n_1516, n2748);
  not g4194 (n_1517, n2749);
  and g4195 (n2750, n_1516, n_1517);
  not g4196 (n_1518, n2750);
  and g4197 (n2751, n2690, n_1518);
  not g4200 (n_1520, n2752);
  and g4201 (n2753, n_272, n_1520);
  and g4202 (n2754, n669, n2752);
  not g4203 (n_1521, n2753);
  not g4204 (n_1522, n2754);
  and g4205 (n2755, n_1521, n_1522);
  not g4206 (n_1523, n2742);
  and g4207 (n2756, n_1523, n2755);
  not g4208 (n_1524, n2756);
  and g4209 (n2757, n_1510, n_1524);
  not g4210 (n_1525, n2683);
  not g4211 (n_1526, n2711);
  and g4212 (n2758, n_1525, n_1526);
  not g4213 (n_1527, n2712);
  not g4214 (n_1528, n2758);
  and g4215 (n2759, n_1527, n_1528);
  not g4216 (n_1529, n2757);
  and g4217 (n2760, n_1529, n2759);
  not g4218 (n_1530, n2760);
  and g4219 (n2761, n_1527, n_1530);
  and g4220 (n2762, n_1385, n2699);
  and g4221 (n2763, n2596, n2695);
  and g4222 (n2764, n2593, n2697);
  not g4228 (n_1534, n2620);
  and g4229 (n2767, n2618, n_1534);
  not g4230 (n_1535, n2767);
  and g4231 (n2768, n_1414, n_1535);
  and g4232 (n2769, n2690, n2768);
  not g4235 (n_1537, n2770);
  and g4236 (n2771, n_272, n_1537);
  and g4237 (n2772, n669, n2770);
  not g4238 (n_1538, n2771);
  not g4239 (n_1539, n2772);
  and g4240 (n2773, n_1538, n_1539);
  and g4241 (n2774, n_1392, n2668);
  and g4242 (n2775, n_245, n2660);
  and g4243 (n2776, n2665, n2775);
  and g4244 (n2777, n_1398, n2776);
  and g4245 (n2778, n_1395, n2666);
  not g4246 (n_1540, n2777);
  not g4247 (n_1541, n2778);
  and g4248 (n2779, n_1540, n_1541);
  not g4249 (n_1542, n2774);
  and g4250 (n2780, n_1542, n2779);
  not g4251 (n_1543, n2674);
  and g4252 (n2781, n_1543, n2780);
  and g4253 (n2782, n_1504, n2780);
  not g4254 (n_1544, n2781);
  not g4255 (n_1545, n2782);
  and g4256 (n2783, n_1544, n_1545);
  not g4257 (n_1546, n2783);
  and g4258 (n2784, n525, n_1546);
  and g4259 (n2785, n_240, n2783);
  not g4260 (n_1547, n2784);
  not g4261 (n_1548, n2785);
  and g4262 (n2786, n_1547, n_1548);
  and g4263 (n2787, n2681, n2786);
  not g4264 (n_1549, n2786);
  and g4265 (n2788, n_1470, n_1549);
  not g4266 (n_1550, n2787);
  not g4267 (n_1551, n2788);
  and g4268 (n2789, n_1550, n_1551);
  and g4269 (n2790, n2773, n2789);
  not g4270 (n_1552, n2773);
  not g4271 (n_1553, n2789);
  and g4272 (n2791, n_1552, n_1553);
  not g4273 (n_1554, n2790);
  not g4274 (n_1555, n2791);
  and g4275 (n2792, n_1554, n_1555);
  not g4276 (n_1556, n2792);
  and g4277 (n2793, n2761, n_1556);
  not g4278 (n_1557, n2761);
  and g4279 (n2794, n_1557, n2792);
  not g4280 (n_1558, n2793);
  not g4281 (n_1559, n2794);
  and g4282 (n2795, n_1558, n_1559);
  and g4283 (n2796, n1013, n_404);
  and g4284 (n2797, n_395, n1021);
  not g4285 (n_1560, n2796);
  not g4286 (n_1561, n2797);
  and g4287 (n2798, n_1560, n_1561);
  and g4288 (n2799, n275, n_464);
  and g4289 (n2800, n_160, n1183);
  not g4290 (n_1562, n2799);
  not g4291 (n_1563, n2800);
  and g4292 (n2801, n_1562, n_1563);
  not g4293 (n_1564, n2801);
  and g4294 (n2802, n2798, n_1564);
  and g4295 (n2803, n2578, n2802);
  and g4296 (n2804, n1013, n_464);
  and g4297 (n2805, n_395, n1183);
  not g4298 (n_1565, n2804);
  not g4299 (n_1566, n2805);
  and g4300 (n2806, n_1565, n_1566);
  not g4301 (n_1567, n2798);
  and g4302 (n2807, n_1567, n2801);
  and g4303 (n2808, n2806, n2807);
  and g4304 (n2809, n_1382, n2808);
  not g4305 (n_1568, n2806);
  and g4306 (n2810, n2801, n_1568);
  and g4307 (n2811, n_1379, n2810);
  not g4308 (n_1569, n2809);
  not g4309 (n_1570, n2811);
  and g4310 (n2812, n_1569, n_1570);
  not g4311 (n_1571, n2803);
  and g4312 (n2813, n_1571, n2812);
  not g4313 (n_1572, n2632);
  and g4314 (n2814, n2630, n_1572);
  not g4315 (n_1573, n2814);
  and g4316 (n2815, n_1427, n_1573);
  not g4317 (n_1574, n2815);
  and g4318 (n2816, n2813, n_1574);
  and g4319 (n2817, n_1567, n_1564);
  not g4320 (n_1575, n2817);
  and g4321 (n2818, n2813, n_1575);
  not g4322 (n_1576, n2816);
  not g4323 (n_1577, n2818);
  and g4324 (n2819, n_1576, n_1577);
  not g4325 (n_1578, n2819);
  and g4326 (n2820, n1021, n_1578);
  and g4327 (n2821, n_404, n2819);
  not g4328 (n_1579, n2820);
  not g4329 (n_1580, n2821);
  and g4330 (n2822, n_1579, n_1580);
  and g4331 (n2823, n2795, n2822);
  and g4332 (n2824, n_1379, n2802);
  and g4333 (n2825, n_1385, n2808);
  and g4334 (n2826, n_1382, n2810);
  not g4340 (n_1584, n2628);
  and g4341 (n2829, n2626, n_1584);
  not g4342 (n_1585, n2829);
  and g4343 (n2830, n_1422, n_1585);
  and g4344 (n2831, n2817, n2830);
  not g4347 (n_1587, n2832);
  and g4348 (n2833, n_404, n_1587);
  not g4349 (n_1588, n2833);
  and g4350 (n2834, n_1587, n_1588);
  and g4351 (n2835, n_404, n_1588);
  not g4352 (n_1589, n2834);
  not g4353 (n_1590, n2835);
  and g4354 (n2836, n_1589, n_1590);
  not g4355 (n_1591, n2759);
  and g4356 (n2837, n2757, n_1591);
  not g4357 (n_1592, n2837);
  and g4358 (n2838, n_1530, n_1592);
  not g4359 (n_1593, n2836);
  and g4360 (n2839, n_1593, n2838);
  and g4361 (n2840, n_1523, n_1524);
  and g4362 (n2841, n2755, n_1524);
  not g4363 (n_1594, n2840);
  not g4364 (n_1595, n2841);
  and g4365 (n2842, n_1594, n_1595);
  and g4366 (n2843, n_1382, n2802);
  and g4367 (n2844, n2593, n2808);
  and g4368 (n2845, n_1385, n2810);
  not g4369 (n_1596, n2844);
  not g4370 (n_1597, n2845);
  and g4371 (n2846, n_1596, n_1597);
  not g4372 (n_1598, n2843);
  and g4373 (n2847, n_1598, n2846);
  not g4374 (n_1599, n2624);
  and g4375 (n2848, n2622, n_1599);
  not g4376 (n_1600, n2848);
  and g4377 (n2849, n_1418, n_1600);
  not g4378 (n_1601, n2849);
  and g4379 (n2850, n2847, n_1601);
  and g4380 (n2851, n_1575, n2847);
  not g4381 (n_1602, n2850);
  not g4382 (n_1603, n2851);
  and g4383 (n2852, n_1602, n_1603);
  not g4384 (n_1604, n2852);
  and g4385 (n2853, n1021, n_1604);
  and g4386 (n2854, n_404, n2852);
  not g4387 (n_1605, n2853);
  not g4388 (n_1606, n2854);
  and g4389 (n2855, n_1605, n_1606);
  not g4390 (n_1607, n2842);
  and g4391 (n2856, n_1607, n2855);
  and g4392 (n2857, n_1385, n2802);
  and g4393 (n2858, n2596, n2808);
  and g4394 (n2859, n2593, n2810);
  and g4400 (n2862, n2768, n2817);
  not g4403 (n_1612, n2863);
  and g4404 (n2864, n_404, n_1612);
  not g4405 (n_1613, n2864);
  and g4406 (n2865, n_1612, n_1613);
  and g4407 (n2866, n_404, n_1613);
  not g4408 (n_1614, n2865);
  not g4409 (n_1615, n2866);
  and g4410 (n2867, n_1614, n_1615);
  not g4411 (n_1616, n2723);
  not g4412 (n_1617, n2737);
  and g4413 (n2868, n_1616, n_1617);
  not g4414 (n_1618, n2738);
  not g4415 (n_1619, n2868);
  and g4416 (n2869, n_1618, n_1619);
  not g4417 (n_1620, n2867);
  and g4418 (n2870, n_1620, n2869);
  not g4419 (n_1621, n2714);
  not g4420 (n_1622, n2722);
  and g4421 (n2871, n_1621, n_1622);
  not g4422 (n_1623, n2871);
  and g4423 (n2872, n_1616, n_1623);
  and g4424 (n2873, n_1392, n2808);
  and g4425 (n2874, n2596, n2810);
  and g4426 (n2875, n2593, n2802);
  not g4427 (n_1624, n2874);
  not g4428 (n_1625, n2875);
  and g4429 (n2876, n_1624, n_1625);
  not g4430 (n_1626, n2873);
  and g4431 (n2877, n_1626, n2876);
  and g4432 (n2878, n_1575, n2877);
  and g4433 (n2879, n2706, n2877);
  not g4434 (n_1627, n2878);
  not g4435 (n_1628, n2879);
  and g4436 (n2880, n_1627, n_1628);
  not g4437 (n_1629, n2880);
  and g4438 (n2881, n1021, n_1629);
  and g4439 (n2882, n_404, n2880);
  not g4440 (n_1630, n2881);
  not g4441 (n_1631, n2882);
  and g4442 (n2883, n_1630, n_1631);
  and g4443 (n2884, n2872, n2883);
  and g4444 (n2885, n_1398, n2810);
  and g4445 (n2886, n_1395, n2802);
  not g4446 (n_1632, n2885);
  not g4447 (n_1633, n2886);
  and g4448 (n2887, n_1632, n_1633);
  and g4449 (n2888, n_1462, n2817);
  not g4450 (n_1634, n2888);
  and g4451 (n2889, n2887, n_1634);
  not g4452 (n_1635, n2889);
  and g4453 (n2890, n_404, n_1635);
  not g4454 (n_1636, n2890);
  and g4455 (n2891, n_404, n_1636);
  and g4456 (n2892, n_1635, n_1636);
  not g4457 (n_1637, n2891);
  not g4458 (n_1638, n2892);
  and g4459 (n2893, n_1637, n_1638);
  and g4460 (n2894, n_1398, n_1564);
  not g4461 (n_1639, n2894);
  and g4462 (n2895, n_404, n_1639);
  not g4463 (n_1640, n2893);
  and g4464 (n2896, n_1640, n2895);
  and g4465 (n2897, n_1392, n2802);
  and g4466 (n2898, n_1398, n2808);
  and g4467 (n2899, n_1395, n2810);
  not g4468 (n_1641, n2898);
  not g4469 (n_1642, n2899);
  and g4470 (n2900, n_1641, n_1642);
  not g4471 (n_1643, n2897);
  and g4472 (n2901, n_1643, n2900);
  and g4473 (n2902, n_1504, n2901);
  and g4474 (n2903, n_1575, n2901);
  not g4475 (n_1644, n2902);
  not g4476 (n_1645, n2903);
  and g4477 (n2904, n_1644, n_1645);
  not g4478 (n_1646, n2904);
  and g4479 (n2905, n1021, n_1646);
  and g4480 (n2906, n_404, n2904);
  not g4481 (n_1647, n2905);
  not g4482 (n_1648, n2906);
  and g4483 (n2907, n_1647, n_1648);
  and g4484 (n2908, n2896, n2907);
  and g4485 (n2909, n2713, n2908);
  not g4486 (n_1649, n2909);
  and g4487 (n2910, n2908, n_1649);
  and g4488 (n2911, n2713, n_1649);
  not g4489 (n_1650, n2910);
  not g4490 (n_1651, n2911);
  and g4491 (n2912, n_1650, n_1651);
  and g4492 (n2913, n_1392, n2810);
  and g4493 (n2914, n2596, n2802);
  and g4494 (n2915, n_1395, n2808);
  and g4500 (n2918, n_1518, n2817);
  not g4503 (n_1656, n2919);
  and g4504 (n2920, n_404, n_1656);
  not g4505 (n_1657, n2920);
  and g4506 (n2921, n_404, n_1657);
  and g4507 (n2922, n_1656, n_1657);
  not g4508 (n_1658, n2921);
  not g4509 (n_1659, n2922);
  and g4510 (n2923, n_1658, n_1659);
  not g4511 (n_1660, n2912);
  not g4512 (n_1661, n2923);
  and g4513 (n2924, n_1660, n_1661);
  not g4514 (n_1662, n2924);
  and g4515 (n2925, n_1649, n_1662);
  not g4516 (n_1663, n2872);
  not g4517 (n_1664, n2883);
  and g4518 (n2926, n_1663, n_1664);
  not g4519 (n_1665, n2884);
  not g4520 (n_1666, n2926);
  and g4521 (n2927, n_1665, n_1666);
  not g4522 (n_1667, n2925);
  and g4523 (n2928, n_1667, n2927);
  not g4524 (n_1668, n2928);
  and g4525 (n2929, n_1665, n_1668);
  not g4526 (n_1669, n2870);
  and g4527 (n2930, n_1620, n_1669);
  and g4528 (n2931, n2869, n_1669);
  not g4529 (n_1670, n2930);
  not g4530 (n_1671, n2931);
  and g4531 (n2932, n_1670, n_1671);
  not g4532 (n_1672, n2929);
  not g4533 (n_1673, n2932);
  and g4534 (n2933, n_1672, n_1673);
  not g4535 (n_1674, n2933);
  and g4536 (n2934, n_1669, n_1674);
  not g4537 (n_1675, n2856);
  and g4538 (n2935, n_1607, n_1675);
  and g4539 (n2936, n2855, n_1675);
  not g4540 (n_1676, n2935);
  not g4541 (n_1677, n2936);
  and g4542 (n2937, n_1676, n_1677);
  not g4543 (n_1678, n2934);
  not g4544 (n_1679, n2937);
  and g4545 (n2938, n_1678, n_1679);
  not g4546 (n_1680, n2938);
  and g4547 (n2939, n_1675, n_1680);
  not g4548 (n_1681, n2839);
  and g4549 (n2940, n_1593, n_1681);
  and g4550 (n2941, n2838, n_1681);
  not g4551 (n_1682, n2940);
  not g4552 (n_1683, n2941);
  and g4553 (n2942, n_1682, n_1683);
  not g4554 (n_1684, n2939);
  not g4555 (n_1685, n2942);
  and g4556 (n2943, n_1684, n_1685);
  not g4557 (n_1686, n2943);
  and g4558 (n2944, n_1681, n_1686);
  not g4559 (n_1687, n2823);
  and g4560 (n2945, n2795, n_1687);
  and g4561 (n2946, n2822, n_1687);
  not g4562 (n_1688, n2945);
  not g4563 (n_1689, n2946);
  and g4564 (n2947, n_1688, n_1689);
  not g4565 (n_1690, n2944);
  not g4566 (n_1691, n2947);
  and g4567 (n2948, n_1690, n_1691);
  not g4568 (n_1692, n2948);
  and g4569 (n2949, n_1687, n_1692);
  and g4570 (n2950, n_1382, n2699);
  and g4571 (n2951, n2593, n2695);
  and g4572 (n2952, n_1385, n2697);
  and g4578 (n2955, n2690, n2849);
  not g4581 (n_1697, n2956);
  and g4582 (n2957, n_272, n_1697);
  and g4583 (n2958, n669, n2956);
  not g4584 (n_1698, n2957);
  not g4585 (n_1699, n2958);
  and g4586 (n2959, n_1698, n_1699);
  and g4587 (n2960, n_1392, n2666);
  and g4588 (n2961, n2596, n2668);
  and g4589 (n2962, n_1395, n2776);
  and g4595 (n2965, n2674, n_1518);
  not g4598 (n_1704, n2966);
  and g4599 (n2967, n_240, n_1704);
  not g4600 (n_1705, n2967);
  and g4601 (n2968, n_1704, n_1705);
  and g4602 (n2969, n_240, n_1705);
  not g4603 (n_1706, n2968);
  not g4604 (n_1707, n2969);
  and g4605 (n2970, n_1706, n_1707);
  and g4606 (n2971, n_240, n_1398);
  not g4607 (n_1708, n2971);
  and g4608 (n2972, n_1550, n_1708);
  and g4609 (n2973, n2787, n2971);
  not g4610 (n_1709, n2970);
  not g4611 (n_1710, n2973);
  and g4612 (n2974, n_1709, n_1710);
  not g4613 (n_1711, n2972);
  and g4614 (n2975, n_1711, n2974);
  not g4615 (n_1712, n2975);
  and g4616 (n2976, n_1709, n_1712);
  and g4617 (n2977, n_1710, n_1712);
  and g4618 (n2978, n_1711, n2977);
  not g4619 (n_1713, n2976);
  not g4620 (n_1714, n2978);
  and g4621 (n2979, n_1713, n_1714);
  not g4622 (n_1715, n2979);
  and g4623 (n2980, n2959, n_1715);
  not g4624 (n_1716, n2980);
  and g4625 (n2981, n2959, n_1716);
  and g4626 (n2982, n_1715, n_1716);
  not g4627 (n_1717, n2981);
  not g4628 (n_1718, n2982);
  and g4629 (n2983, n_1717, n_1718);
  and g4630 (n2984, n_1554, n_1559);
  and g4631 (n2985, n2983, n2984);
  not g4632 (n_1719, n2983);
  not g4633 (n_1720, n2984);
  and g4634 (n2986, n_1719, n_1720);
  not g4635 (n_1721, n2985);
  not g4636 (n_1722, n2986);
  and g4637 (n2987, n_1721, n_1722);
  not g4638 (n_1723, n2636);
  and g4639 (n2988, n2634, n_1723);
  not g4640 (n_1724, n2988);
  and g4641 (n2989, n_1431, n_1724);
  and g4642 (n2990, n_1374, n2802);
  and g4643 (n2991, n_1379, n2808);
  and g4644 (n2992, n2578, n2810);
  not g4645 (n_1725, n2991);
  not g4646 (n_1726, n2992);
  and g4647 (n2993, n_1725, n_1726);
  not g4648 (n_1727, n2990);
  and g4649 (n2994, n_1727, n2993);
  not g4650 (n_1728, n2989);
  and g4651 (n2995, n_1728, n2994);
  and g4652 (n2996, n_1575, n2994);
  not g4653 (n_1729, n2995);
  not g4654 (n_1730, n2996);
  and g4655 (n2997, n_1729, n_1730);
  not g4656 (n_1731, n2997);
  and g4657 (n2998, n1021, n_1731);
  and g4658 (n2999, n_404, n2997);
  not g4659 (n_1732, n2998);
  not g4660 (n_1733, n2999);
  and g4661 (n3000, n_1732, n_1733);
  and g4662 (n3001, n2987, n3000);
  not g4663 (n_1734, n3001);
  and g4664 (n3002, n2987, n_1734);
  and g4665 (n3003, n3000, n_1734);
  not g4666 (n_1735, n3002);
  not g4667 (n_1736, n3003);
  and g4668 (n3004, n_1735, n_1736);
  not g4669 (n_1737, n2949);
  not g4670 (n_1738, n3004);
  and g4671 (n3005, n_1737, n_1738);
  not g4672 (n_1739, n3005);
  and g4673 (n3006, n_1737, n_1739);
  and g4674 (n3007, n_1738, n_1739);
  not g4675 (n_1740, n3006);
  not g4676 (n_1741, n3007);
  and g4677 (n3008, n_1740, n_1741);
  not g4678 (n_1742, n3008);
  and g4679 (n3009, n2657, n_1742);
  not g4680 (n_1743, n3009);
  and g4681 (n3010, n2657, n_1743);
  and g4682 (n3011, n_1742, n_1743);
  not g4683 (n_1744, n3010);
  not g4684 (n_1745, n3011);
  and g4685 (n3012, n_1744, n_1745);
  and g4686 (n3013, n_1690, n_1692);
  and g4687 (n3014, n_1691, n_1692);
  not g4688 (n_1746, n3013);
  not g4689 (n_1747, n3014);
  and g4690 (n3015, n_1746, n_1747);
  and g4691 (n3016, n295, n_1368);
  and g4692 (n3017, n2560, n_1374);
  and g4693 (n3018, n2562, n2567);
  not g4699 (n_1751, n2644);
  and g4700 (n3021, n2642, n_1751);
  not g4701 (n_1752, n3021);
  and g4702 (n3022, n_1440, n_1752);
  and g4703 (n3023, n2571, n3022);
  not g4706 (n_1754, n3024);
  and g4707 (n3025, n_160, n_1754);
  and g4708 (n3026, n275, n3024);
  not g4709 (n_1755, n3025);
  not g4710 (n_1756, n3026);
  and g4711 (n3027, n_1755, n_1756);
  not g4712 (n_1757, n3015);
  and g4713 (n3028, n_1757, n3027);
  not g4714 (n_1758, n3028);
  and g4715 (n3029, n3027, n_1758);
  and g4716 (n3030, n_1757, n_1758);
  not g4717 (n_1759, n3029);
  not g4718 (n_1760, n3030);
  and g4719 (n3031, n_1759, n_1760);
  and g4720 (n3032, n_1684, n2942);
  and g4721 (n3033, n2939, n_1685);
  not g4722 (n_1761, n3032);
  not g4723 (n_1762, n3033);
  and g4724 (n3034, n_1761, n_1762);
  and g4725 (n3035, n295, n2562);
  and g4726 (n3036, n2560, n2578);
  and g4727 (n3037, n2567, n_1374);
  not g4728 (n_1763, n3036);
  not g4729 (n_1764, n3037);
  and g4730 (n3038, n_1763, n_1764);
  not g4731 (n_1765, n3035);
  and g4732 (n3039, n_1765, n3038);
  not g4733 (n_1766, n2571);
  and g4734 (n3040, n_1766, n3039);
  not g4735 (n_1767, n2640);
  and g4736 (n3041, n2638, n_1767);
  not g4737 (n_1768, n3041);
  and g4738 (n3042, n_1436, n_1768);
  not g4739 (n_1769, n3042);
  and g4740 (n3043, n3039, n_1769);
  not g4741 (n_1770, n3040);
  not g4742 (n_1771, n3043);
  and g4743 (n3044, n_1770, n_1771);
  not g4744 (n_1772, n3044);
  and g4745 (n3045, n275, n_1772);
  and g4746 (n3046, n_160, n3044);
  not g4747 (n_1773, n3045);
  not g4748 (n_1774, n3046);
  and g4749 (n3047, n_1773, n_1774);
  not g4750 (n_1775, n3034);
  and g4751 (n3048, n_1775, n3047);
  and g4752 (n3049, n_1678, n_1680);
  and g4753 (n3050, n_1679, n_1680);
  not g4754 (n_1776, n3049);
  not g4755 (n_1777, n3050);
  and g4756 (n3051, n_1776, n_1777);
  and g4757 (n3052, n295, n_1374);
  and g4758 (n3053, n2560, n_1379);
  and g4759 (n3054, n2567, n2578);
  not g4760 (n_1778, n3053);
  not g4761 (n_1779, n3054);
  and g4762 (n3055, n_1778, n_1779);
  not g4763 (n_1780, n3052);
  and g4764 (n3056, n_1780, n3055);
  and g4765 (n3057, n_1766, n3056);
  and g4766 (n3058, n_1728, n3056);
  not g4767 (n_1781, n3057);
  not g4768 (n_1782, n3058);
  and g4769 (n3059, n_1781, n_1782);
  not g4770 (n_1783, n3059);
  and g4771 (n3060, n275, n_1783);
  and g4772 (n3061, n_160, n3059);
  not g4773 (n_1784, n3060);
  not g4774 (n_1785, n3061);
  and g4775 (n3062, n_1784, n_1785);
  not g4776 (n_1786, n3051);
  and g4777 (n3063, n_1786, n3062);
  and g4778 (n3064, n_1672, n2932);
  and g4779 (n3065, n2929, n_1673);
  not g4780 (n_1787, n3064);
  not g4781 (n_1788, n3065);
  and g4782 (n3066, n_1787, n_1788);
  and g4783 (n3067, n295, n2578);
  and g4784 (n3068, n2560, n_1382);
  and g4785 (n3069, n2567, n_1379);
  not g4786 (n_1789, n3068);
  not g4787 (n_1790, n3069);
  and g4788 (n3070, n_1789, n_1790);
  not g4789 (n_1791, n3067);
  and g4790 (n3071, n_1791, n3070);
  and g4791 (n3072, n_1766, n3071);
  and g4792 (n3073, n_1574, n3071);
  not g4793 (n_1792, n3072);
  not g4794 (n_1793, n3073);
  and g4795 (n3074, n_1792, n_1793);
  not g4796 (n_1794, n3074);
  and g4797 (n3075, n275, n_1794);
  and g4798 (n3076, n_160, n3074);
  not g4799 (n_1795, n3075);
  not g4800 (n_1796, n3076);
  and g4801 (n3077, n_1795, n_1796);
  not g4802 (n_1797, n3066);
  and g4803 (n3078, n_1797, n3077);
  and g4804 (n3079, n295, n_1379);
  and g4805 (n3080, n2560, n_1385);
  and g4806 (n3081, n2567, n_1382);
  and g4812 (n3084, n2571, n2830);
  not g4815 (n_1802, n3085);
  and g4816 (n3086, n_160, n_1802);
  and g4817 (n3087, n275, n3085);
  not g4818 (n_1803, n3086);
  not g4819 (n_1804, n3087);
  and g4820 (n3088, n_1803, n_1804);
  not g4821 (n_1805, n2927);
  and g4822 (n3089, n2925, n_1805);
  not g4823 (n_1806, n3089);
  and g4824 (n3090, n_1668, n_1806);
  and g4825 (n3091, n3088, n3090);
  and g4826 (n3092, n_1660, n_1662);
  and g4827 (n3093, n_1661, n_1662);
  not g4828 (n_1807, n3092);
  not g4829 (n_1808, n3093);
  and g4830 (n3094, n_1807, n_1808);
  and g4831 (n3095, n295, n_1382);
  and g4832 (n3096, n2560, n2593);
  and g4833 (n3097, n2567, n_1385);
  not g4834 (n_1809, n3096);
  not g4835 (n_1810, n3097);
  and g4836 (n3098, n_1809, n_1810);
  not g4837 (n_1811, n3095);
  and g4838 (n3099, n_1811, n3098);
  and g4839 (n3100, n_1766, n3099);
  and g4840 (n3101, n_1601, n3099);
  not g4841 (n_1812, n3100);
  not g4842 (n_1813, n3101);
  and g4843 (n3102, n_1812, n_1813);
  not g4844 (n_1814, n3102);
  and g4845 (n3103, n275, n_1814);
  and g4846 (n3104, n_160, n3102);
  not g4847 (n_1815, n3103);
  not g4848 (n_1816, n3104);
  and g4849 (n3105, n_1815, n_1816);
  not g4850 (n_1817, n3094);
  and g4851 (n3106, n_1817, n3105);
  and g4852 (n3107, n295, n_1385);
  and g4853 (n3108, n2560, n2596);
  and g4854 (n3109, n2567, n2593);
  and g4860 (n3112, n2571, n2768);
  not g4863 (n_1822, n3113);
  and g4864 (n3114, n_160, n_1822);
  and g4865 (n3115, n275, n3113);
  not g4866 (n_1823, n3114);
  not g4867 (n_1824, n3115);
  and g4868 (n3116, n_1823, n_1824);
  not g4869 (n_1825, n2896);
  not g4870 (n_1826, n2907);
  and g4871 (n3117, n_1825, n_1826);
  not g4872 (n_1827, n2908);
  not g4873 (n_1828, n3117);
  and g4874 (n3118, n_1827, n_1828);
  and g4875 (n3119, n3116, n3118);
  not g4876 (n_1829, n2895);
  and g4877 (n3120, n2893, n_1829);
  not g4878 (n_1830, n3120);
  and g4879 (n3121, n_1825, n_1830);
  and g4880 (n3122, n2560, n_1392);
  and g4881 (n3123, n2567, n2596);
  and g4882 (n3124, n295, n2593);
  not g4883 (n_1831, n3123);
  not g4884 (n_1832, n3124);
  and g4885 (n3125, n_1831, n_1832);
  not g4886 (n_1833, n3122);
  and g4887 (n3126, n_1833, n3125);
  and g4888 (n3127, n_1766, n3126);
  and g4889 (n3128, n2706, n3126);
  not g4890 (n_1834, n3127);
  not g4891 (n_1835, n3128);
  and g4892 (n3129, n_1834, n_1835);
  not g4893 (n_1836, n3129);
  and g4894 (n3130, n275, n_1836);
  and g4895 (n3131, n_160, n3129);
  not g4896 (n_1837, n3130);
  not g4897 (n_1838, n3131);
  and g4898 (n3132, n_1837, n_1838);
  and g4899 (n3133, n3121, n3132);
  and g4900 (n3134, n_175, n_1398);
  not g4901 (n_1839, n3134);
  and g4902 (n3135, n_160, n_1839);
  and g4903 (n3136, n2567, n_1398);
  and g4904 (n3137, n295, n_1395);
  not g4905 (n_1840, n3136);
  not g4906 (n_1841, n3137);
  and g4907 (n3138, n_1840, n_1841);
  and g4908 (n3139, n2571, n_1462);
  not g4909 (n_1842, n3139);
  and g4910 (n3140, n3138, n_1842);
  not g4911 (n_1843, n3140);
  and g4912 (n3141, n_160, n_1843);
  and g4913 (n3142, n275, n3140);
  not g4914 (n_1844, n3141);
  not g4915 (n_1845, n3142);
  and g4916 (n3143, n_1844, n_1845);
  and g4917 (n3144, n3135, n3143);
  and g4918 (n3145, n295, n_1392);
  and g4919 (n3146, n2560, n_1398);
  and g4920 (n3147, n2567, n_1395);
  not g4921 (n_1846, n3146);
  not g4922 (n_1847, n3147);
  and g4923 (n3148, n_1846, n_1847);
  not g4924 (n_1848, n3145);
  and g4925 (n3149, n_1848, n3148);
  and g4926 (n3150, n_1766, n3149);
  and g4927 (n3151, n_1504, n3149);
  not g4928 (n_1849, n3150);
  not g4929 (n_1850, n3151);
  and g4930 (n3152, n_1849, n_1850);
  not g4931 (n_1851, n3152);
  and g4932 (n3153, n275, n_1851);
  and g4933 (n3154, n_160, n3152);
  not g4934 (n_1852, n3153);
  not g4935 (n_1853, n3154);
  and g4936 (n3155, n_1852, n_1853);
  and g4937 (n3156, n3144, n3155);
  and g4938 (n3157, n2894, n3156);
  not g4939 (n_1854, n3157);
  and g4940 (n3158, n3156, n_1854);
  and g4941 (n3159, n2894, n_1854);
  not g4942 (n_1855, n3158);
  not g4943 (n_1856, n3159);
  and g4944 (n3160, n_1855, n_1856);
  and g4945 (n3161, n2567, n_1392);
  and g4946 (n3162, n295, n2596);
  and g4947 (n3163, n2560, n_1395);
  and g4953 (n3166, n2571, n_1518);
  not g4956 (n_1861, n3167);
  and g4957 (n3168, n_160, n_1861);
  and g4958 (n3169, n275, n3167);
  not g4959 (n_1862, n3168);
  not g4960 (n_1863, n3169);
  and g4961 (n3170, n_1862, n_1863);
  not g4962 (n_1864, n3160);
  and g4963 (n3171, n_1864, n3170);
  not g4964 (n_1865, n3171);
  and g4965 (n3172, n_1854, n_1865);
  not g4966 (n_1866, n3121);
  not g4967 (n_1867, n3132);
  and g4968 (n3173, n_1866, n_1867);
  not g4969 (n_1868, n3133);
  not g4970 (n_1869, n3173);
  and g4971 (n3174, n_1868, n_1869);
  not g4972 (n_1870, n3172);
  and g4973 (n3175, n_1870, n3174);
  not g4974 (n_1871, n3175);
  and g4975 (n3176, n_1868, n_1871);
  not g4976 (n_1872, n3116);
  not g4977 (n_1873, n3118);
  and g4978 (n3177, n_1872, n_1873);
  not g4979 (n_1874, n3119);
  not g4980 (n_1875, n3177);
  and g4981 (n3178, n_1874, n_1875);
  not g4982 (n_1876, n3176);
  and g4983 (n3179, n_1876, n3178);
  not g4984 (n_1877, n3179);
  and g4985 (n3180, n_1874, n_1877);
  not g4986 (n_1878, n3106);
  and g4987 (n3181, n_1817, n_1878);
  and g4988 (n3182, n3105, n_1878);
  not g4989 (n_1879, n3181);
  not g4990 (n_1880, n3182);
  and g4991 (n3183, n_1879, n_1880);
  not g4992 (n_1881, n3180);
  not g4993 (n_1882, n3183);
  and g4994 (n3184, n_1881, n_1882);
  not g4995 (n_1883, n3184);
  and g4996 (n3185, n_1878, n_1883);
  not g4997 (n_1884, n3088);
  not g4998 (n_1885, n3090);
  and g4999 (n3186, n_1884, n_1885);
  not g5000 (n_1886, n3091);
  not g5001 (n_1887, n3186);
  and g5002 (n3187, n_1886, n_1887);
  not g5003 (n_1888, n3185);
  and g5004 (n3188, n_1888, n3187);
  not g5005 (n_1889, n3188);
  and g5006 (n3189, n_1886, n_1889);
  not g5007 (n_1890, n3078);
  and g5008 (n3190, n_1797, n_1890);
  and g5009 (n3191, n3077, n_1890);
  not g5010 (n_1891, n3190);
  not g5011 (n_1892, n3191);
  and g5012 (n3192, n_1891, n_1892);
  not g5013 (n_1893, n3189);
  not g5014 (n_1894, n3192);
  and g5015 (n3193, n_1893, n_1894);
  not g5016 (n_1895, n3193);
  and g5017 (n3194, n_1890, n_1895);
  not g5018 (n_1896, n3063);
  and g5019 (n3195, n_1786, n_1896);
  and g5020 (n3196, n3062, n_1896);
  not g5021 (n_1897, n3195);
  not g5022 (n_1898, n3196);
  and g5023 (n3197, n_1897, n_1898);
  not g5024 (n_1899, n3194);
  not g5025 (n_1900, n3197);
  and g5026 (n3198, n_1899, n_1900);
  not g5027 (n_1901, n3198);
  and g5028 (n3199, n_1896, n_1901);
  not g5029 (n_1902, n3047);
  and g5030 (n3200, n3034, n_1902);
  not g5031 (n_1903, n3048);
  not g5032 (n_1904, n3200);
  and g5033 (n3201, n_1903, n_1904);
  not g5034 (n_1905, n3199);
  and g5035 (n3202, n_1905, n3201);
  not g5036 (n_1906, n3202);
  and g5037 (n3203, n_1903, n_1906);
  not g5038 (n_1907, n3031);
  not g5039 (n_1908, n3203);
  and g5040 (n3204, n_1907, n_1908);
  not g5041 (n_1909, n3204);
  and g5042 (n3205, n_1758, n_1909);
  and g5043 (n3206, n3012, n3205);
  not g5044 (n_1910, n3012);
  not g5045 (n_1911, n3205);
  and g5046 (n3207, n_1910, n_1911);
  not g5047 (n_1912, n3206);
  not g5048 (n_1913, n3207);
  and g5049 (n3208, n_1912, n_1913);
  and g5050 (n3209, \a[0] , n_49);
  not g5051 (n_1914, n3209);
  and g5052 (n3210, \a[1] , n_1914);
  and g5053 (n3211, n_5, n3209);
  not g5054 (n_1915, n3210);
  not g5055 (n_1916, n3211);
  and g5056 (n3212, n_1915, n_1916);
  and g5057 (n3213, n_171, n3212);
  not g5058 (n_1917, n3212);
  and g5059 (n3214, n291, n_1917);
  not g5060 (n_1918, n3213);
  not g5061 (n_1919, n3214);
  and g5062 (n3215, n_1918, n_1919);
  not g5063 (n_1920, n3215);
  and g5064 (n3216, \a[0] , n_1920);
  and g5065 (n3217, \a[0] , n3215);
  and g5078 (n3230, n_176, n808);
  and g5079 (n3231, n_190, n3230);
  and g5105 (n3257, n2552, n3256);
  and g5106 (n3258, n3229, n3257);
  and g5107 (n3259, n_95, n_211);
  not g5118 (n_1921, n3258);
  and g5119 (n3270, n_1921, n3269);
  not g5120 (n_1922, n3269);
  and g5121 (n3271, n3258, n_1922);
  not g5122 (n_1923, n3270);
  not g5123 (n_1924, n3271);
  and g5124 (n3272, n_1923, n_1924);
  and g5125 (n3273, n3217, n3272);
  and g5126 (n3274, n288, n_1920);
  and g5127 (n3275, n_1357, n3256);
  not g5128 (n_1925, n3256);
  and g5129 (n3276, n2552, n_1925);
  not g5130 (n_1926, n3275);
  not g5131 (n_1927, n3276);
  and g5132 (n3277, n_1926, n_1927);
  and g5133 (n3278, n3274, n3277);
  not g5134 (n_1928, n3229);
  not g5135 (n_1929, n3257);
  and g5136 (n3279, n_1928, n_1929);
  not g5137 (n_1930, n3279);
  and g5138 (n3280, n_1921, n_1930);
  and g5139 (n3281, n_8, n_1917);
  not g5140 (n_1931, n3280);
  and g5141 (n3282, n_1931, n3281);
  not g5142 (n_1932, n3278);
  not g5143 (n_1933, n3282);
  and g5144 (n3283, n_1932, n_1933);
  not g5145 (n_1934, n3273);
  and g5146 (n3284, n_1934, n3283);
  not g5147 (n_1935, n3216);
  and g5148 (n3285, n_1935, n3284);
  and g5149 (n3286, n3277, n_1931);
  and g5150 (n3287, n_1359, n3277);
  and g5151 (n3288, n_1441, n_1445);
  not g5152 (n_1936, n3277);
  and g5153 (n3289, n2554, n_1936);
  not g5154 (n_1937, n3287);
  not g5155 (n_1938, n3289);
  and g5156 (n3290, n_1937, n_1938);
  not g5157 (n_1939, n3288);
  and g5158 (n3291, n_1939, n3290);
  not g5159 (n_1940, n3291);
  and g5160 (n3292, n_1937, n_1940);
  and g5161 (n3293, n_1936, n3280);
  not g5162 (n_1941, n3286);
  not g5163 (n_1942, n3293);
  and g5164 (n3294, n_1941, n_1942);
  not g5165 (n_1943, n3292);
  and g5166 (n3295, n_1943, n3294);
  not g5167 (n_1944, n3295);
  and g5168 (n3296, n_1941, n_1944);
  not g5169 (n_1945, n3272);
  and g5170 (n3297, n_1945, n3280);
  and g5171 (n3298, n3272, n_1931);
  not g5172 (n_1946, n3297);
  not g5173 (n_1947, n3298);
  and g5174 (n3299, n_1946, n_1947);
  not g5175 (n_1948, n3296);
  and g5176 (n3300, n_1948, n3299);
  not g5177 (n_1949, n3299);
  and g5178 (n3301, n3296, n_1949);
  not g5179 (n_1950, n3300);
  not g5180 (n_1951, n3301);
  and g5181 (n3302, n_1950, n_1951);
  not g5182 (n_1952, n3302);
  and g5183 (n3303, n3284, n_1952);
  not g5184 (n_1953, n3285);
  not g5185 (n_1954, n3303);
  and g5186 (n3304, n_1953, n_1954);
  not g5187 (n_1955, n3304);
  and g5188 (n3305, n291, n_1955);
  and g5189 (n3306, n_171, n3304);
  not g5190 (n_1956, n3305);
  not g5191 (n_1957, n3306);
  and g5192 (n3307, n_1956, n_1957);
  and g5193 (n3308, n3208, n3307);
  and g5194 (n3309, n3031, n3203);
  not g5195 (n_1958, n3309);
  and g5196 (n3310, n_1909, n_1958);
  and g5197 (n3311, n3217, n_1931);
  and g5198 (n3312, n_1359, n3274);
  and g5199 (n3313, n3277, n3281);
  not g5200 (n_1959, n3312);
  not g5201 (n_1960, n3313);
  and g5202 (n3314, n_1959, n_1960);
  not g5203 (n_1961, n3311);
  and g5204 (n3315, n_1961, n3314);
  and g5205 (n3316, n_1935, n3315);
  not g5206 (n_1962, n3294);
  and g5207 (n3317, n3292, n_1962);
  not g5208 (n_1963, n3317);
  and g5209 (n3318, n_1944, n_1963);
  not g5210 (n_1964, n3318);
  and g5211 (n3319, n3315, n_1964);
  not g5212 (n_1965, n3316);
  not g5213 (n_1966, n3319);
  and g5214 (n3320, n_1965, n_1966);
  not g5215 (n_1967, n3320);
  and g5216 (n3321, n291, n_1967);
  and g5217 (n3322, n_171, n3320);
  not g5218 (n_1968, n3321);
  not g5219 (n_1969, n3322);
  and g5220 (n3323, n_1968, n_1969);
  and g5221 (n3324, n3310, n3323);
  not g5222 (n_1970, n3201);
  and g5223 (n3325, n3199, n_1970);
  and g5224 (n3326, n3217, n3277);
  and g5225 (n3327, n_1368, n3274);
  and g5226 (n3328, n_1359, n3281);
  not g5232 (n_1974, n3290);
  and g5233 (n3331, n3288, n_1974);
  not g5234 (n_1975, n3331);
  and g5235 (n3332, n_1940, n_1975);
  and g5236 (n3333, n3216, n3332);
  not g5239 (n_1977, n3334);
  and g5240 (n3335, n_171, n_1977);
  not g5241 (n_1978, n3335);
  and g5242 (n3336, n_1977, n_1978);
  and g5243 (n3337, n_171, n_1978);
  not g5244 (n_1979, n3336);
  not g5245 (n_1980, n3337);
  and g5246 (n3338, n_1979, n_1980);
  and g5247 (n3339, n2562, n3217);
  and g5248 (n3340, n2578, n3274);
  and g5249 (n3341, n_1374, n3281);
  not g5250 (n_1981, n3340);
  not g5251 (n_1982, n3341);
  and g5252 (n3342, n_1981, n_1982);
  not g5253 (n_1983, n3339);
  and g5254 (n3343, n_1983, n3342);
  not g5255 (n_1984, n3343);
  and g5256 (n3344, n_171, n_1984);
  and g5257 (n3345, n3042, n3216);
  not g5258 (n_1985, n3345);
  and g5259 (n3346, n3343, n_1985);
  and g5260 (n3347, n291, n3346);
  and g5261 (n3348, n_171, n3216);
  and g5262 (n3349, n3042, n3348);
  and g5263 (n3350, n_1374, n3217);
  and g5264 (n3351, n_1379, n3274);
  and g5265 (n3352, n2578, n3281);
  not g5266 (n_1986, n3351);
  not g5267 (n_1987, n3352);
  and g5268 (n3353, n_1986, n_1987);
  not g5269 (n_1988, n3350);
  and g5270 (n3354, n_1988, n3353);
  not g5271 (n_1989, n3354);
  and g5272 (n3355, n_171, n_1989);
  and g5273 (n3356, n2989, n3216);
  not g5274 (n_1990, n3356);
  and g5275 (n3357, n3354, n_1990);
  and g5276 (n3358, n291, n3357);
  and g5277 (n3359, n2989, n3348);
  and g5278 (n3360, n2578, n3217);
  and g5279 (n3361, n_1382, n3274);
  and g5280 (n3362, n_1379, n3281);
  not g5281 (n_1991, n3361);
  not g5282 (n_1992, n3362);
  and g5283 (n3363, n_1991, n_1992);
  not g5284 (n_1993, n3360);
  and g5285 (n3364, n_1993, n3363);
  not g5286 (n_1994, n3364);
  and g5287 (n3365, n_171, n_1994);
  and g5288 (n3366, n2815, n3216);
  not g5289 (n_1995, n3366);
  and g5290 (n3367, n3364, n_1995);
  and g5291 (n3368, n291, n3367);
  and g5292 (n3369, n2815, n3348);
  not g5293 (n_1996, n3174);
  and g5294 (n3370, n3172, n_1996);
  and g5295 (n3371, n_1382, n3217);
  and g5296 (n3372, n2593, n3274);
  and g5297 (n3373, n_1385, n3281);
  not g5298 (n_1997, n3372);
  not g5299 (n_1998, n3373);
  and g5300 (n3374, n_1997, n_1998);
  not g5301 (n_1999, n3371);
  and g5302 (n3375, n_1999, n3374);
  not g5303 (n_2000, n3375);
  and g5304 (n3376, n_171, n_2000);
  and g5305 (n3377, n2849, n3216);
  not g5306 (n_2001, n3377);
  and g5307 (n3378, n3375, n_2001);
  and g5308 (n3379, n291, n3378);
  and g5309 (n3380, n2849, n3348);
  not g5310 (n_2002, n3144);
  not g5311 (n_2003, n3155);
  and g5312 (n3381, n_2002, n_2003);
  and g5313 (n3382, n_1392, n3274);
  and g5314 (n3383, n2596, n3281);
  and g5315 (n3384, n2593, n3217);
  not g5316 (n_2004, n3383);
  not g5317 (n_2005, n3384);
  and g5318 (n3385, n_2004, n_2005);
  not g5319 (n_2006, n3382);
  and g5320 (n3386, n_2006, n3385);
  not g5321 (n_2007, n3386);
  and g5322 (n3387, n_171, n_2007);
  not g5323 (n_2008, n2706);
  and g5324 (n3388, n_2008, n3216);
  not g5325 (n_2009, n3388);
  and g5326 (n3389, n3386, n_2009);
  and g5327 (n3390, n291, n3389);
  and g5328 (n3391, n_2008, n3348);
  and g5329 (n3392, \a[0] , n_1398);
  and g5330 (n3393, n2732, n3348);
  and g5331 (n3394, n_1392, n3217);
  and g5332 (n3395, n_1398, n3274);
  and g5333 (n3396, n_1395, n3281);
  not g5334 (n_2010, n3395);
  not g5335 (n_2011, n3396);
  and g5336 (n3397, n_2010, n_2011);
  not g5337 (n_2012, n3394);
  and g5338 (n3398, n_2012, n3397);
  not g5339 (n_2013, n3398);
  and g5340 (n3399, n_171, n_2013);
  and g5341 (n3400, n_1462, n3348);
  and g5342 (n3401, n_1395, n3217);
  and g5343 (n3402, n_1398, n3281);
  not g5356 (n_2020, n3408);
  and g5357 (n3409, n_1839, n_2020);
  and g5358 (n3410, n_1392, n3281);
  and g5359 (n3411, n2596, n3217);
  and g5360 (n3412, n_1395, n3274);
  and g5366 (n3415, n_1518, n3216);
  not g5369 (n_2025, n3416);
  and g5370 (n3417, n_171, n_2025);
  and g5371 (n3418, n291, n3416);
  not g5372 (n_2026, n3417);
  not g5373 (n_2027, n3418);
  and g5374 (n3419, n_2026, n_2027);
  not g5375 (n_2028, n3409);
  and g5376 (n3420, n_2028, n3419);
  and g5377 (n3421, n3134, n3408);
  not g5378 (n_2029, n3420);
  not g5379 (n_2030, n3421);
  and g5380 (n3422, n_2029, n_2030);
  not g5381 (n_2031, n3135);
  not g5382 (n_2032, n3143);
  and g5383 (n3423, n_2031, n_2032);
  not g5384 (n_2033, n3423);
  and g5385 (n3424, n_2002, n_2033);
  not g5386 (n_2034, n3424);
  and g5387 (n3425, n3422, n_2034);
  not g5395 (n_2039, n3422);
  and g5396 (n3429, n_2039, n3424);
  not g5397 (n_2040, n3428);
  not g5398 (n_2041, n3429);
  and g5399 (n3430, n_2040, n_2041);
  and g5400 (n3431, n_1385, n3217);
  and g5401 (n3432, n2596, n3274);
  and g5402 (n3433, n2593, n3281);
  and g5408 (n3436, n2768, n3216);
  not g5411 (n_2046, n3437);
  and g5412 (n3438, n_171, n_2046);
  not g5413 (n_2047, n3438);
  and g5414 (n3439, n_2046, n_2047);
  and g5415 (n3440, n_171, n_2047);
  not g5416 (n_2048, n3439);
  not g5417 (n_2049, n3440);
  and g5418 (n3441, n_2048, n_2049);
  and g5419 (n3442, n3430, n3441);
  not g5420 (n_2050, n3156);
  not g5421 (n_2051, n3442);
  and g5422 (n3443, n_2050, n_2051);
  not g5423 (n_2052, n3381);
  and g5424 (n3444, n_2052, n3443);
  not g5425 (n_2053, n3430);
  not g5426 (n_2054, n3441);
  and g5427 (n3445, n_2053, n_2054);
  not g5428 (n_2055, n3444);
  not g5429 (n_2056, n3445);
  and g5430 (n3446, n_2055, n_2056);
  and g5431 (n3447, n_1864, n_1865);
  and g5432 (n3448, n3170, n_1865);
  not g5433 (n_2057, n3447);
  not g5434 (n_2058, n3448);
  and g5435 (n3449, n_2057, n_2058);
  and g5436 (n3450, n3446, n3449);
  not g5444 (n_2063, n3446);
  not g5445 (n_2064, n3449);
  and g5446 (n3454, n_2063, n_2064);
  not g5447 (n_2065, n3453);
  not g5448 (n_2066, n3454);
  and g5449 (n3455, n_2065, n_2066);
  and g5450 (n3456, n_1379, n3217);
  and g5451 (n3457, n_1385, n3274);
  and g5452 (n3458, n_1382, n3281);
  and g5458 (n3461, n2830, n3216);
  not g5461 (n_2071, n3462);
  and g5462 (n3463, n_171, n_2071);
  not g5463 (n_2072, n3463);
  and g5464 (n3464, n_2071, n_2072);
  and g5465 (n3465, n_171, n_2072);
  not g5466 (n_2073, n3464);
  not g5467 (n_2074, n3465);
  and g5468 (n3466, n_2073, n_2074);
  and g5469 (n3467, n3455, n3466);
  not g5470 (n_2075, n3467);
  and g5471 (n3468, n_1871, n_2075);
  not g5472 (n_2076, n3370);
  and g5473 (n3469, n_2076, n3468);
  not g5474 (n_2077, n3455);
  not g5475 (n_2078, n3466);
  and g5476 (n3470, n_2077, n_2078);
  not g5477 (n_2079, n3469);
  not g5478 (n_2080, n3470);
  and g5479 (n3471, n_2079, n_2080);
  not g5480 (n_2081, n3178);
  and g5481 (n3472, n3176, n_2081);
  not g5482 (n_2082, n3472);
  and g5483 (n3473, n_1877, n_2082);
  not g5484 (n_2083, n3473);
  and g5485 (n3474, n3471, n_2083);
  not g5493 (n_2088, n3471);
  and g5494 (n3478, n_2088, n3473);
  not g5495 (n_2089, n3477);
  not g5496 (n_2090, n3478);
  and g5497 (n3479, n_2089, n_2090);
  and g5498 (n3480, n_1881, n_1883);
  and g5499 (n3481, n_1882, n_1883);
  not g5500 (n_2091, n3480);
  not g5501 (n_2092, n3481);
  and g5502 (n3482, n_2091, n_2092);
  and g5503 (n3483, n3479, n3482);
  not g5511 (n_2097, n3479);
  not g5512 (n_2098, n3482);
  and g5513 (n3487, n_2097, n_2098);
  not g5514 (n_2099, n3486);
  not g5515 (n_2100, n3487);
  and g5516 (n3488, n_2099, n_2100);
  not g5517 (n_2101, n3187);
  and g5518 (n3489, n3185, n_2101);
  not g5519 (n_2102, n3489);
  and g5520 (n3490, n_1889, n_2102);
  not g5521 (n_2103, n3490);
  and g5522 (n3491, n3488, n_2103);
  not g5530 (n_2108, n3488);
  and g5531 (n3495, n_2108, n3490);
  not g5532 (n_2109, n3494);
  not g5533 (n_2110, n3495);
  and g5534 (n3496, n_2109, n_2110);
  and g5535 (n3497, n3189, n3192);
  not g5536 (n_2111, n3497);
  and g5537 (n3498, n_1895, n_2111);
  not g5538 (n_2112, n3496);
  and g5539 (n3499, n_2112, n3498);
  and g5540 (n3500, n_1368, n3217);
  and g5541 (n3501, n_1374, n3274);
  and g5542 (n3502, n2562, n3281);
  and g5548 (n3505, n3022, n3216);
  not g5551 (n_2117, n3506);
  and g5552 (n3507, n291, n_2117);
  and g5553 (n3508, n_171, n3506);
  not g5554 (n_2118, n3507);
  not g5555 (n_2119, n3508);
  and g5556 (n3509, n_2118, n_2119);
  not g5557 (n_2120, n3499);
  and g5558 (n3510, n_2120, n3509);
  not g5559 (n_2121, n3498);
  and g5560 (n3511, n3496, n_2121);
  not g5561 (n_2122, n3510);
  not g5562 (n_2123, n3511);
  and g5563 (n3512, n_2122, n_2123);
  and g5564 (n3513, n3194, n3197);
  not g5565 (n_2124, n3513);
  and g5566 (n3514, n_1901, n_2124);
  not g5567 (n_2125, n3512);
  not g5568 (n_2126, n3514);
  and g5569 (n3515, n_2125, n_2126);
  and g5570 (n3516, n_1359, n3217);
  and g5571 (n3517, n2562, n3274);
  and g5572 (n3518, n_1368, n3281);
  and g5578 (n3521, n2652, n3216);
  not g5581 (n_2131, n3522);
  and g5582 (n3523, n_171, n_2131);
  and g5583 (n3524, n291, n3522);
  not g5584 (n_2132, n3523);
  not g5585 (n_2133, n3524);
  and g5586 (n3525, n_2132, n_2133);
  not g5587 (n_2134, n3515);
  and g5588 (n3526, n_2134, n3525);
  and g5589 (n3527, n3512, n3514);
  not g5590 (n_2135, n3526);
  not g5591 (n_2136, n3527);
  and g5592 (n3528, n_2135, n_2136);
  and g5593 (n3529, n3338, n3528);
  not g5594 (n_2137, n3529);
  and g5595 (n3530, n_1906, n_2137);
  not g5596 (n_2138, n3325);
  and g5597 (n3531, n_2138, n3530);
  not g5598 (n_2139, n3338);
  not g5599 (n_2140, n3528);
  and g5600 (n3532, n_2139, n_2140);
  not g5601 (n_2141, n3531);
  not g5602 (n_2142, n3532);
  and g5603 (n3533, n_2141, n_2142);
  not g5604 (n_2143, n3324);
  and g5605 (n3534, n3310, n_2143);
  and g5606 (n3535, n3323, n_2143);
  not g5607 (n_2144, n3534);
  not g5608 (n_2145, n3535);
  and g5609 (n3536, n_2144, n_2145);
  not g5610 (n_2146, n3533);
  not g5611 (n_2147, n3536);
  and g5612 (n3537, n_2146, n_2147);
  not g5613 (n_2148, n3537);
  and g5614 (n3538, n_2143, n_2148);
  not g5615 (n_2149, n3308);
  and g5616 (n3539, n3208, n_2149);
  and g5617 (n3540, n3307, n_2149);
  not g5618 (n_2150, n3539);
  not g5619 (n_2151, n3540);
  and g5620 (n3541, n_2150, n_2151);
  not g5621 (n_2152, n3538);
  not g5622 (n_2153, n3541);
  and g5623 (n3542, n_2152, n_2153);
  not g5624 (n_2154, n3542);
  and g5625 (n3543, n_2149, n_2154);
  and g5626 (n3544, n_1743, n_1913);
  and g5627 (n3545, n295, n3277);
  and g5628 (n3546, n2560, n_1368);
  and g5629 (n3547, n_1359, n2567);
  and g5635 (n3550, n2571, n3332);
  not g5638 (n_2159, n3551);
  and g5639 (n3552, n_160, n_2159);
  and g5640 (n3553, n275, n3551);
  not g5641 (n_2160, n3552);
  not g5642 (n_2161, n3553);
  and g5643 (n3554, n_2160, n_2161);
  and g5644 (n3555, n_1734, n_1739);
  and g5645 (n3556, n_1716, n_1722);
  and g5646 (n3557, n_1379, n2699);
  and g5647 (n3558, n_1385, n2695);
  and g5648 (n3559, n_1382, n2697);
  and g5654 (n3562, n2690, n2830);
  not g5657 (n_2166, n3563);
  and g5658 (n3564, n_272, n_2166);
  and g5659 (n3565, n669, n3563);
  not g5660 (n_2167, n3564);
  not g5661 (n_2168, n3565);
  and g5662 (n3566, n_2167, n_2168);
  and g5663 (n3567, n_240, n_1395);
  and g5664 (n3568, n_1392, n2776);
  and g5665 (n3569, n2596, n2666);
  and g5666 (n3570, n2593, n2668);
  and g5672 (n3573, n2674, n_2008);
  not g5675 (n_2173, n3574);
  and g5676 (n3575, n_240, n_2173);
  not g5677 (n_2174, n3575);
  and g5678 (n3576, n3567, n_2174);
  not g5679 (n_2175, n3576);
  and g5680 (n3577, n3567, n_2175);
  and g5681 (n3578, n525, n3574);
  not g5682 (n_2176, n3578);
  and g5683 (n3579, n_2174, n_2176);
  and g5684 (n3580, n_2175, n3579);
  not g5685 (n_2177, n3577);
  not g5686 (n_2178, n3580);
  and g5687 (n3581, n_2177, n_2178);
  not g5688 (n_2179, n2977);
  not g5689 (n_2180, n3581);
  and g5690 (n3582, n_2179, n_2180);
  not g5691 (n_2181, n3582);
  and g5692 (n3583, n_2179, n_2181);
  and g5693 (n3584, n_2180, n_2181);
  not g5694 (n_2182, n3583);
  not g5695 (n_2183, n3584);
  and g5696 (n3585, n_2182, n_2183);
  not g5697 (n_2184, n3585);
  and g5698 (n3586, n3566, n_2184);
  not g5699 (n_2185, n3586);
  and g5700 (n3587, n3566, n_2185);
  and g5701 (n3588, n_2184, n_2185);
  not g5702 (n_2186, n3587);
  not g5703 (n_2187, n3588);
  and g5704 (n3589, n_2186, n_2187);
  not g5705 (n_2188, n3556);
  and g5706 (n3590, n_2188, n3589);
  not g5707 (n_2189, n3589);
  and g5708 (n3591, n3556, n_2189);
  not g5709 (n_2190, n3590);
  not g5710 (n_2191, n3591);
  and g5711 (n3592, n_2190, n_2191);
  and g5712 (n3593, n2562, n2802);
  and g5713 (n3594, n2578, n2808);
  and g5714 (n3595, n_1374, n2810);
  not g5715 (n_2192, n3594);
  not g5716 (n_2193, n3595);
  and g5717 (n3596, n_2192, n_2193);
  not g5718 (n_2194, n3593);
  and g5719 (n3597, n_2194, n3596);
  and g5720 (n3598, n_1769, n3597);
  and g5721 (n3599, n_1575, n3597);
  not g5722 (n_2195, n3598);
  not g5723 (n_2196, n3599);
  and g5724 (n3600, n_2195, n_2196);
  not g5725 (n_2197, n3600);
  and g5726 (n3601, n1021, n_2197);
  and g5727 (n3602, n_404, n3600);
  not g5728 (n_2198, n3601);
  not g5729 (n_2199, n3602);
  and g5730 (n3603, n_2198, n_2199);
  not g5731 (n_2200, n3592);
  and g5732 (n3604, n_2200, n3603);
  not g5733 (n_2201, n3603);
  and g5734 (n3605, n3592, n_2201);
  not g5735 (n_2202, n3604);
  not g5736 (n_2203, n3605);
  and g5737 (n3606, n_2202, n_2203);
  not g5738 (n_2204, n3555);
  and g5739 (n3607, n_2204, n3606);
  not g5740 (n_2205, n3606);
  and g5741 (n3608, n3555, n_2205);
  not g5742 (n_2206, n3607);
  not g5743 (n_2207, n3608);
  and g5744 (n3609, n_2206, n_2207);
  and g5745 (n3610, n3554, n3609);
  not g5746 (n_2208, n3554);
  not g5747 (n_2209, n3609);
  and g5748 (n3611, n_2208, n_2209);
  not g5749 (n_2210, n3610);
  not g5750 (n_2211, n3611);
  and g5751 (n3612, n_2210, n_2211);
  not g5752 (n_2212, n3544);
  and g5753 (n3613, n_2212, n3612);
  not g5754 (n_2213, n3612);
  and g5755 (n3614, n3544, n_2213);
  not g5756 (n_2214, n3613);
  not g5757 (n_2215, n3614);
  and g5758 (n3615, n_2214, n_2215);
  and g5759 (n3616, n_198, n502);
  and g5760 (n3617, n_88, n3616);
  and g5768 (n3625, n3258, n3269);
  not g5769 (n_2216, n3624);
  not g5770 (n_2217, n3625);
  and g5771 (n3626, n_2216, n_2217);
  and g5772 (n3627, n3624, n3625);
  not g5773 (n_2218, n3626);
  not g5774 (n_2219, n3627);
  and g5775 (n3628, n_2218, n_2219);
  not g5776 (n_2220, n3628);
  and g5777 (n3629, n3217, n_2220);
  and g5778 (n3630, n3274, n_1931);
  and g5779 (n3631, n3272, n3281);
  not g5780 (n_2221, n3630);
  not g5781 (n_2222, n3631);
  and g5782 (n3632, n_2221, n_2222);
  not g5783 (n_2223, n3629);
  and g5784 (n3633, n_2223, n3632);
  and g5785 (n3634, n_1935, n3633);
  and g5786 (n3635, n_1947, n_1950);
  and g5787 (n3636, n_1945, n3628);
  and g5788 (n3637, n3272, n_2220);
  not g5789 (n_2224, n3636);
  not g5790 (n_2225, n3637);
  and g5791 (n3638, n_2224, n_2225);
  not g5792 (n_2226, n3635);
  and g5793 (n3639, n_2226, n3638);
  not g5794 (n_2227, n3638);
  and g5795 (n3640, n3635, n_2227);
  not g5796 (n_2228, n3639);
  not g5797 (n_2229, n3640);
  and g5798 (n3641, n_2228, n_2229);
  not g5799 (n_2230, n3641);
  and g5800 (n3642, n3633, n_2230);
  not g5801 (n_2231, n3634);
  not g5802 (n_2232, n3642);
  and g5803 (n3643, n_2231, n_2232);
  not g5804 (n_2233, n3643);
  and g5805 (n3644, n291, n_2233);
  and g5806 (n3645, n_171, n3643);
  not g5807 (n_2234, n3644);
  not g5808 (n_2235, n3645);
  and g5809 (n3646, n_2234, n_2235);
  and g5810 (n3647, n3615, n3646);
  not g5811 (n_2236, n3615);
  not g5812 (n_2237, n3646);
  and g5813 (n3648, n_2236, n_2237);
  not g5814 (n_2238, n3647);
  not g5815 (n_2239, n3648);
  and g5816 (n3649, n_2238, n_2239);
  not g5817 (n_2240, n3543);
  and g5818 (n3650, n_2240, n3649);
  not g5819 (n_2241, n3649);
  and g5820 (n3651, n3543, n_2241);
  not g5821 (n_2242, n3650);
  not g5822 (n_2243, n3651);
  and g5823 (n3652, n_2242, n_2243);
  not g5824 (n_2244, n271);
  and g5825 (n3653, n_2244, n3652);
  and g5863 (n3691, n3538, n_2151);
  and g5864 (n3692, n_2150, n3691);
  not g5865 (n_2245, n3692);
  and g5866 (n3693, n_2154, n_2245);
  and g5889 (n3716, n3533, n3536);
  not g5890 (n_2246, n3716);
  and g5891 (n3717, n_2148, n_2246);
  not g5892 (n_2247, n3715);
  and g5893 (n3718, n_2247, n3717);
  not g5894 (n_2248, n3693);
  not g5895 (n_2249, n3718);
  and g5896 (n3719, n_2248, n_2249);
  not g5897 (n_2250, n3690);
  not g5898 (n_2251, n3719);
  and g5899 (n3720, n_2250, n_2251);
  and g5900 (n3721, n3693, n3718);
  not g5901 (n_2252, n3720);
  not g5902 (n_2253, n3721);
  and g5903 (n3722, n_2252, n_2253);
  not g5904 (n_2254, n3653);
  and g5905 (n3723, n_2244, n_2254);
  and g5906 (n3724, n3652, n_2254);
  not g5907 (n_2255, n3723);
  not g5908 (n_2256, n3724);
  and g5909 (n3725, n_2255, n_2256);
  not g5910 (n_2257, n3722);
  not g5911 (n_2258, n3725);
  and g5912 (n3726, n_2257, n_2258);
  not g5913 (n_2259, n3726);
  and g5914 (n3727, n_2254, n_2259);
  and g5935 (n3748, n_2219, n3747);
  not g5936 (n_2260, n3747);
  and g5937 (n3749, n3627, n_2260);
  not g5938 (n_2261, n3748);
  not g5939 (n_2262, n3749);
  and g5940 (n3750, n_2261, n_2262);
  and g5941 (n3751, n3217, n3750);
  and g5942 (n3752, n3272, n3274);
  and g5943 (n3753, n3281, n_2220);
  and g5949 (n3756, n_2225, n_2228);
  not g5950 (n_2266, n3750);
  and g5951 (n3757, n3628, n_2266);
  and g5952 (n3758, n_2220, n3750);
  not g5953 (n_2267, n3757);
  not g5954 (n_2268, n3758);
  and g5955 (n3759, n_2267, n_2268);
  not g5956 (n_2269, n3756);
  and g5957 (n3760, n_2269, n3759);
  not g5958 (n_2270, n3759);
  and g5959 (n3761, n3756, n_2270);
  not g5960 (n_2271, n3760);
  not g5961 (n_2272, n3761);
  and g5962 (n3762, n_2271, n_2272);
  and g5963 (n3763, n3216, n3762);
  not g5966 (n_2274, n3764);
  and g5967 (n3765, n_171, n_2274);
  not g5968 (n_2275, n3765);
  and g5969 (n3766, n_2274, n_2275);
  and g5970 (n3767, n_171, n_2275);
  not g5971 (n_2276, n3766);
  not g5972 (n_2277, n3767);
  and g5973 (n3768, n_2276, n_2277);
  and g5974 (n3769, n_2210, n_2214);
  and g5975 (n3770, n_1368, n2802);
  and g5976 (n3771, n_1374, n2808);
  and g5977 (n3772, n2562, n2810);
  and g5983 (n3775, n2817, n3022);
  not g5986 (n_2282, n3776);
  and g5987 (n3777, n_404, n_2282);
  not g5988 (n_2283, n3777);
  and g5989 (n3778, n_2282, n_2283);
  and g5990 (n3779, n_404, n_2283);
  not g5991 (n_2284, n3778);
  not g5992 (n_2285, n3779);
  and g5993 (n3780, n_2284, n_2285);
  and g5994 (n3781, n_2188, n_2189);
  not g5995 (n_2286, n3781);
  and g5996 (n3782, n_2185, n_2286);
  and g5997 (n3783, n_2175, n_2181);
  and g5998 (n3784, n_1385, n2668);
  and g5999 (n3785, n2596, n2776);
  and g6000 (n3786, n2593, n2666);
  and g6006 (n3789, n2674, n2768);
  and g6009 (n3791, n_240, n2600);
  not g6010 (n_2291, n3790);
  and g6011 (n3792, n_2291, n3791);
  not g6012 (n_2292, n3791);
  and g6013 (n3793, n3790, n_2292);
  not g6014 (n_2293, n3792);
  not g6015 (n_2294, n3793);
  and g6016 (n3794, n_2293, n_2294);
  not g6017 (n_2295, n3783);
  and g6018 (n3795, n_2295, n3794);
  not g6019 (n_2296, n3794);
  and g6020 (n3796, n3783, n_2296);
  not g6021 (n_2297, n3795);
  not g6022 (n_2298, n3796);
  and g6023 (n3797, n_2297, n_2298);
  and g6024 (n3798, n2578, n2699);
  and g6025 (n3799, n_1382, n2695);
  and g6026 (n3800, n_1379, n2697);
  not g6027 (n_2299, n3799);
  not g6028 (n_2300, n3800);
  and g6029 (n3801, n_2299, n_2300);
  not g6030 (n_2301, n3798);
  and g6031 (n3802, n_2301, n3801);
  and g6032 (n3803, n_1484, n3802);
  and g6033 (n3804, n_1574, n3802);
  not g6034 (n_2302, n3803);
  not g6035 (n_2303, n3804);
  and g6036 (n3805, n_2302, n_2303);
  not g6037 (n_2304, n3805);
  and g6038 (n3806, n669, n_2304);
  and g6039 (n3807, n_272, n3805);
  not g6040 (n_2305, n3806);
  not g6041 (n_2306, n3807);
  and g6042 (n3808, n_2305, n_2306);
  and g6043 (n3809, n3797, n3808);
  not g6044 (n_2307, n3809);
  and g6045 (n3810, n3797, n_2307);
  and g6046 (n3811, n3808, n_2307);
  not g6047 (n_2308, n3810);
  not g6048 (n_2309, n3811);
  and g6049 (n3812, n_2308, n_2309);
  not g6050 (n_2310, n3782);
  not g6051 (n_2311, n3812);
  and g6052 (n3813, n_2310, n_2311);
  not g6053 (n_2312, n3813);
  and g6054 (n3814, n_2310, n_2312);
  and g6055 (n3815, n_2311, n_2312);
  not g6056 (n_2313, n3814);
  not g6057 (n_2314, n3815);
  and g6058 (n3816, n_2313, n_2314);
  not g6059 (n_2315, n3780);
  not g6060 (n_2316, n3816);
  and g6061 (n3817, n_2315, n_2316);
  not g6062 (n_2317, n3817);
  and g6063 (n3818, n_2315, n_2317);
  and g6064 (n3819, n_2316, n_2317);
  not g6065 (n_2318, n3818);
  not g6066 (n_2319, n3819);
  and g6067 (n3820, n_2318, n_2319);
  and g6068 (n3821, n_2202, n_2206);
  and g6069 (n3822, n3820, n3821);
  not g6070 (n_2320, n3820);
  not g6071 (n_2321, n3821);
  and g6072 (n3823, n_2320, n_2321);
  not g6073 (n_2322, n3822);
  not g6074 (n_2323, n3823);
  and g6075 (n3824, n_2322, n_2323);
  and g6076 (n3825, n295, n_1931);
  and g6077 (n3826, n_1359, n2560);
  and g6078 (n3827, n2567, n3277);
  not g6079 (n_2324, n3826);
  not g6080 (n_2325, n3827);
  and g6081 (n3828, n_2324, n_2325);
  not g6082 (n_2326, n3825);
  and g6083 (n3829, n_2326, n3828);
  and g6084 (n3830, n_1766, n3829);
  and g6085 (n3831, n_1964, n3829);
  not g6086 (n_2327, n3830);
  not g6087 (n_2328, n3831);
  and g6088 (n3832, n_2327, n_2328);
  not g6089 (n_2329, n3832);
  and g6090 (n3833, n275, n_2329);
  and g6091 (n3834, n_160, n3832);
  not g6092 (n_2330, n3833);
  not g6093 (n_2331, n3834);
  and g6094 (n3835, n_2330, n_2331);
  and g6095 (n3836, n3824, n3835);
  not g6096 (n_2332, n3836);
  and g6097 (n3837, n3824, n_2332);
  and g6098 (n3838, n3835, n_2332);
  not g6099 (n_2333, n3837);
  not g6100 (n_2334, n3838);
  and g6101 (n3839, n_2333, n_2334);
  not g6102 (n_2335, n3769);
  not g6103 (n_2336, n3839);
  and g6104 (n3840, n_2335, n_2336);
  not g6105 (n_2337, n3840);
  and g6106 (n3841, n_2335, n_2337);
  and g6107 (n3842, n_2336, n_2337);
  not g6108 (n_2338, n3841);
  not g6109 (n_2339, n3842);
  and g6110 (n3843, n_2338, n_2339);
  not g6111 (n_2340, n3768);
  not g6112 (n_2341, n3843);
  and g6113 (n3844, n_2340, n_2341);
  not g6114 (n_2342, n3844);
  and g6115 (n3845, n_2340, n_2342);
  and g6116 (n3846, n_2341, n_2342);
  not g6117 (n_2343, n3845);
  not g6118 (n_2344, n3846);
  and g6119 (n3847, n_2343, n_2344);
  and g6120 (n3848, n_2238, n_2242);
  and g6121 (n3849, n3847, n3848);
  not g6122 (n_2345, n3847);
  not g6123 (n_2346, n3848);
  and g6124 (n3850, n_2345, n_2346);
  not g6125 (n_2347, n3849);
  not g6126 (n_2348, n3850);
  and g6127 (n3851, n_2347, n_2348);
  not g6138 (n_2349, n3851);
  and g6139 (n3862, n_2349, n3861);
  not g6140 (n_2350, n3861);
  and g6141 (n3863, n3851, n_2350);
  not g6142 (n_2351, n3862);
  not g6143 (n_2352, n3863);
  and g6144 (n3864, n_2351, n_2352);
  not g6145 (n_2353, n3727);
  and g6146 (n3865, n_2353, n3864);
  not g6147 (n_2354, n3864);
  and g6148 (n3866, n3727, n_2354);
  not g6149 (n_2355, n3865);
  not g6150 (n_2356, n3866);
  and g6151 (n3867, n_2355, n_2356);
  and g6152 (n3868, n_2257, n_2259);
  and g6153 (n3869, n_2258, n_2259);
  not g6154 (n_2357, n3868);
  not g6155 (n_2358, n3869);
  and g6156 (n3870, n_2357, n_2358);
  not g6157 (n_2359, n3870);
  and g6158 (n3871, n3867, n_2359);
  not g6159 (n_2360, n3871);
  and g6160 (n3872, n3867, n_2360);
  and g6161 (n3873, n_2359, n_2360);
  or g6162 (\sin[0] , n3872, n3873);
  and g6163 (n3875, n_2352, n_2355);
  and g6164 (n3876, n3627, n3747);
  not g6182 (n_2361, n3876);
  and g6183 (n3894, n_2361, n3893);
  not g6184 (n_2362, n3893);
  and g6185 (n3895, n3876, n_2362);
  not g6186 (n_2363, n3894);
  not g6187 (n_2364, n3895);
  and g6188 (n3896, n_2363, n_2364);
  and g6189 (n3897, n3217, n3896);
  and g6190 (n3898, n3274, n_2220);
  and g6191 (n3899, n3281, n3750);
  and g6197 (n3902, n_2268, n_2271);
  not g6198 (n_2368, n3896);
  and g6199 (n3903, n_2266, n_2368);
  and g6200 (n3904, n3750, n3896);
  not g6201 (n_2369, n3903);
  not g6202 (n_2370, n3904);
  and g6203 (n3905, n_2369, n_2370);
  not g6204 (n_2371, n3902);
  and g6205 (n3906, n_2371, n3905);
  not g6206 (n_2372, n3905);
  and g6207 (n3907, n3902, n_2372);
  not g6208 (n_2373, n3906);
  not g6209 (n_2374, n3907);
  and g6210 (n3908, n_2373, n_2374);
  and g6211 (n3909, n3216, n3908);
  not g6214 (n_2376, n3910);
  and g6215 (n3911, n_171, n_2376);
  not g6216 (n_2377, n3911);
  and g6217 (n3912, n_2376, n_2377);
  and g6218 (n3913, n_171, n_2377);
  not g6219 (n_2378, n3912);
  not g6220 (n_2379, n3913);
  and g6221 (n3914, n_2378, n_2379);
  and g6222 (n3915, n_2332, n_2337);
  and g6223 (n3916, n_1359, n2802);
  and g6224 (n3917, n2562, n2808);
  and g6225 (n3918, n_1368, n2810);
  and g6231 (n3921, n2652, n2817);
  not g6234 (n_2384, n3922);
  and g6235 (n3923, n_404, n_2384);
  not g6236 (n_2385, n3923);
  and g6237 (n3924, n_2384, n_2385);
  and g6238 (n3925, n_404, n_2385);
  not g6239 (n_2386, n3924);
  not g6240 (n_2387, n3925);
  and g6241 (n3926, n_2386, n_2387);
  and g6242 (n3927, n_2307, n_2312);
  and g6243 (n3928, n_240, n_1392);
  and g6244 (n3929, n3790, n3928);
  not g6245 (n_2388, n3929);
  and g6246 (n3930, n_2297, n_2388);
  and g6247 (n3931, n_1382, n2668);
  and g6248 (n3932, n2593, n2776);
  and g6249 (n3933, n_1385, n2666);
  and g6255 (n3936, n2674, n2849);
  and g6258 (n3938, n_240, n_1401);
  not g6259 (n_2393, n3937);
  and g6260 (n3939, n_2393, n3938);
  not g6261 (n_2394, n3938);
  and g6262 (n3940, n3937, n_2394);
  not g6263 (n_2395, n3939);
  not g6264 (n_2396, n3940);
  and g6265 (n3941, n_2395, n_2396);
  not g6266 (n_2397, n3930);
  and g6267 (n3942, n_2397, n3941);
  not g6268 (n_2398, n3942);
  and g6269 (n3943, n_2397, n_2398);
  and g6270 (n3944, n3941, n_2398);
  not g6271 (n_2399, n3943);
  not g6272 (n_2400, n3944);
  and g6273 (n3945, n_2399, n_2400);
  and g6274 (n3946, n_1374, n2699);
  and g6275 (n3947, n_1379, n2695);
  and g6276 (n3948, n2578, n2697);
  not g6277 (n_2401, n3947);
  not g6278 (n_2402, n3948);
  and g6279 (n3949, n_2401, n_2402);
  not g6280 (n_2403, n3946);
  and g6281 (n3950, n_2403, n3949);
  and g6282 (n3951, n_1484, n3950);
  and g6283 (n3952, n_1728, n3950);
  not g6284 (n_2404, n3951);
  not g6285 (n_2405, n3952);
  and g6286 (n3953, n_2404, n_2405);
  not g6287 (n_2406, n3953);
  and g6288 (n3954, n669, n_2406);
  and g6289 (n3955, n_272, n3953);
  not g6290 (n_2407, n3954);
  not g6291 (n_2408, n3955);
  and g6292 (n3956, n_2407, n_2408);
  not g6293 (n_2409, n3945);
  and g6294 (n3957, n_2409, n3956);
  not g6295 (n_2410, n3957);
  and g6296 (n3958, n_2409, n_2410);
  and g6297 (n3959, n3956, n_2410);
  not g6298 (n_2411, n3958);
  not g6299 (n_2412, n3959);
  and g6300 (n3960, n_2411, n_2412);
  not g6301 (n_2413, n3927);
  not g6302 (n_2414, n3960);
  and g6303 (n3961, n_2413, n_2414);
  not g6304 (n_2415, n3961);
  and g6305 (n3962, n_2413, n_2415);
  and g6306 (n3963, n_2414, n_2415);
  not g6307 (n_2416, n3962);
  not g6308 (n_2417, n3963);
  and g6309 (n3964, n_2416, n_2417);
  not g6310 (n_2418, n3926);
  not g6311 (n_2419, n3964);
  and g6312 (n3965, n_2418, n_2419);
  not g6313 (n_2420, n3965);
  and g6314 (n3966, n_2418, n_2420);
  and g6315 (n3967, n_2419, n_2420);
  not g6316 (n_2421, n3966);
  not g6317 (n_2422, n3967);
  and g6318 (n3968, n_2421, n_2422);
  and g6319 (n3969, n_2317, n_2323);
  and g6320 (n3970, n3968, n3969);
  not g6321 (n_2423, n3968);
  not g6322 (n_2424, n3969);
  and g6323 (n3971, n_2423, n_2424);
  not g6324 (n_2425, n3970);
  not g6325 (n_2426, n3971);
  and g6326 (n3972, n_2425, n_2426);
  and g6327 (n3973, n295, n3272);
  and g6328 (n3974, n2560, n3277);
  and g6329 (n3975, n2567, n_1931);
  not g6330 (n_2427, n3974);
  not g6331 (n_2428, n3975);
  and g6332 (n3976, n_2427, n_2428);
  not g6333 (n_2429, n3973);
  and g6334 (n3977, n_2429, n3976);
  and g6335 (n3978, n_1766, n3977);
  and g6336 (n3979, n_1952, n3977);
  not g6337 (n_2430, n3978);
  not g6338 (n_2431, n3979);
  and g6339 (n3980, n_2430, n_2431);
  not g6340 (n_2432, n3980);
  and g6341 (n3981, n275, n_2432);
  and g6342 (n3982, n_160, n3980);
  not g6343 (n_2433, n3981);
  not g6344 (n_2434, n3982);
  and g6345 (n3983, n_2433, n_2434);
  and g6346 (n3984, n3972, n3983);
  not g6347 (n_2435, n3984);
  and g6348 (n3985, n3972, n_2435);
  and g6349 (n3986, n3983, n_2435);
  not g6350 (n_2436, n3985);
  not g6351 (n_2437, n3986);
  and g6352 (n3987, n_2436, n_2437);
  not g6353 (n_2438, n3915);
  not g6354 (n_2439, n3987);
  and g6355 (n3988, n_2438, n_2439);
  not g6356 (n_2440, n3988);
  and g6357 (n3989, n_2438, n_2440);
  and g6358 (n3990, n_2439, n_2440);
  not g6359 (n_2441, n3989);
  not g6360 (n_2442, n3990);
  and g6361 (n3991, n_2441, n_2442);
  not g6362 (n_2443, n3914);
  not g6363 (n_2444, n3991);
  and g6364 (n3992, n_2443, n_2444);
  not g6365 (n_2445, n3992);
  and g6366 (n3993, n_2443, n_2445);
  and g6367 (n3994, n_2444, n_2445);
  not g6368 (n_2446, n3993);
  not g6369 (n_2447, n3994);
  and g6370 (n3995, n_2446, n_2447);
  and g6371 (n3996, n_2342, n_2348);
  and g6372 (n3997, n3995, n3996);
  not g6373 (n_2448, n3995);
  not g6374 (n_2449, n3996);
  and g6375 (n3998, n_2448, n_2449);
  not g6376 (n_2450, n3997);
  not g6377 (n_2451, n3998);
  and g6378 (n3999, n_2450, n_2451);
  not g6395 (n_2452, n3999);
  and g6396 (n4016, n_2452, n4015);
  not g6397 (n_2453, n4015);
  and g6398 (n4017, n3999, n_2453);
  not g6399 (n_2454, n4016);
  not g6400 (n_2455, n4017);
  and g6401 (n4018, n_2454, n_2455);
  not g6402 (n_2456, n3875);
  and g6403 (n4019, n_2456, n4018);
  not g6404 (n_2457, n4018);
  and g6405 (n4020, n3875, n_2457);
  not g6406 (n_2458, n4019);
  not g6407 (n_2459, n4020);
  and g6408 (n4021, n_2458, n_2459);
  and g6409 (n4022, n3871, n4021);
  not g6410 (n_2460, n4021);
  and g6411 (n4023, n_2360, n_2460);
  not g6412 (n_2461, n4022);
  not g6413 (n_2462, n4023);
  and g6414 (n4024, n_2461, n_2462);
  not g6415 (n_2464, \a[23] );
  and g6416 (n4025, \a[22] , n_2464);
  and g6417 (n4026, n_49, \a[23] );
  not g6418 (n_2465, n4025);
  not g6419 (n_2466, n4026);
  and g6420 (n4027, n_2465, n_2466);
  not g6421 (n_2468, n4027);
  and g6422 (n4028, \sin[0] , n_2468);
  not g6423 (n_2469, n4024);
  and g6424 (n4029, n_2469, n4028);
  not g6425 (n_2470, n4028);
  and g6426 (n4030, n4024, n_2470);
  or g6427 (\sin[1] , n4029, n4030);
  and g6428 (n4032, n_2455, n_2458);
  and g6445 (n4049, n_2445, n_2451);
  and g6446 (n4050, n3274, n3750);
  and g6447 (n4051, n3281, n3896);
  not g6448 (n_2471, n4050);
  not g6449 (n_2472, n4051);
  and g6450 (n4052, n_2471, n_2472);
  and g6451 (n4053, n_2266, n_2373);
  not g6452 (n_2473, n4053);
  and g6453 (n4054, n3896, n_2473);
  and g6454 (n4055, n_2368, n_2373);
  not g6455 (n_2474, n4054);
  not g6456 (n_2475, n4055);
  and g6457 (n4056, n_2474, n_2475);
  and g6458 (n4057, n3216, n4056);
  not g6459 (n_2476, n4057);
  and g6460 (n4058, n4052, n_2476);
  not g6461 (n_2477, n4058);
  and g6462 (n4059, n_171, n_2477);
  not g6463 (n_2478, n4059);
  and g6464 (n4060, n_2477, n_2478);
  and g6465 (n4061, n_171, n_2478);
  not g6466 (n_2479, n4060);
  not g6467 (n_2480, n4061);
  and g6468 (n4062, n_2479, n_2480);
  and g6469 (n4063, n_2435, n_2440);
  and g6470 (n4064, n2802, n3277);
  and g6471 (n4065, n_1368, n2808);
  and g6472 (n4066, n_1359, n2810);
  and g6478 (n4069, n2817, n3332);
  not g6481 (n_2485, n4070);
  and g6482 (n4071, n_404, n_2485);
  not g6483 (n_2486, n4071);
  and g6484 (n4072, n_2485, n_2486);
  and g6485 (n4073, n_404, n_2486);
  not g6486 (n_2487, n4072);
  not g6487 (n_2488, n4073);
  and g6488 (n4074, n_2487, n_2488);
  and g6489 (n4075, n_2410, n_2415);
  and g6490 (n4076, n_240, n3937);
  and g6491 (n4077, n2596, n4076);
  not g6492 (n_2489, n4077);
  and g6493 (n4078, n_2398, n_2489);
  and g6494 (n4079, n_1379, n2668);
  and g6495 (n4080, n_1385, n2776);
  and g6496 (n4081, n_1382, n2666);
  and g6502 (n4084, n2674, n2830);
  and g6505 (n4086, n_240, n_1406);
  not g6506 (n_2494, n4085);
  and g6507 (n4087, n_2494, n4086);
  not g6508 (n_2495, n4086);
  and g6509 (n4088, n4085, n_2495);
  not g6510 (n_2496, n4087);
  not g6511 (n_2497, n4088);
  and g6512 (n4089, n_2496, n_2497);
  not g6513 (n_2498, n4078);
  and g6514 (n4090, n_2498, n4089);
  not g6515 (n_2499, n4090);
  and g6516 (n4091, n_2498, n_2499);
  and g6517 (n4092, n4089, n_2499);
  not g6518 (n_2500, n4091);
  not g6519 (n_2501, n4092);
  and g6520 (n4093, n_2500, n_2501);
  and g6521 (n4094, n2562, n2699);
  and g6522 (n4095, n2578, n2695);
  and g6523 (n4096, n_1374, n2697);
  not g6524 (n_2502, n4095);
  not g6525 (n_2503, n4096);
  and g6526 (n4097, n_2502, n_2503);
  not g6527 (n_2504, n4094);
  and g6528 (n4098, n_2504, n4097);
  and g6529 (n4099, n_1484, n4098);
  and g6530 (n4100, n_1769, n4098);
  not g6531 (n_2505, n4099);
  not g6532 (n_2506, n4100);
  and g6533 (n4101, n_2505, n_2506);
  not g6534 (n_2507, n4101);
  and g6535 (n4102, n669, n_2507);
  and g6536 (n4103, n_272, n4101);
  not g6537 (n_2508, n4102);
  not g6538 (n_2509, n4103);
  and g6539 (n4104, n_2508, n_2509);
  not g6540 (n_2510, n4093);
  and g6541 (n4105, n_2510, n4104);
  not g6542 (n_2511, n4105);
  and g6543 (n4106, n_2510, n_2511);
  and g6544 (n4107, n4104, n_2511);
  not g6545 (n_2512, n4106);
  not g6546 (n_2513, n4107);
  and g6547 (n4108, n_2512, n_2513);
  not g6548 (n_2514, n4075);
  not g6549 (n_2515, n4108);
  and g6550 (n4109, n_2514, n_2515);
  not g6551 (n_2516, n4109);
  and g6552 (n4110, n_2514, n_2516);
  and g6553 (n4111, n_2515, n_2516);
  not g6554 (n_2517, n4110);
  not g6555 (n_2518, n4111);
  and g6556 (n4112, n_2517, n_2518);
  not g6557 (n_2519, n4074);
  not g6558 (n_2520, n4112);
  and g6559 (n4113, n_2519, n_2520);
  not g6560 (n_2521, n4113);
  and g6561 (n4114, n_2519, n_2521);
  and g6562 (n4115, n_2520, n_2521);
  not g6563 (n_2522, n4114);
  not g6564 (n_2523, n4115);
  and g6565 (n4116, n_2522, n_2523);
  and g6566 (n4117, n_2420, n_2426);
  and g6567 (n4118, n4116, n4117);
  not g6568 (n_2524, n4116);
  not g6569 (n_2525, n4117);
  and g6570 (n4119, n_2524, n_2525);
  not g6571 (n_2526, n4118);
  not g6572 (n_2527, n4119);
  and g6573 (n4120, n_2526, n_2527);
  and g6574 (n4121, n295, n_2220);
  and g6575 (n4122, n2560, n_1931);
  and g6576 (n4123, n2567, n3272);
  not g6577 (n_2528, n4122);
  not g6578 (n_2529, n4123);
  and g6579 (n4124, n_2528, n_2529);
  not g6580 (n_2530, n4121);
  and g6581 (n4125, n_2530, n4124);
  and g6582 (n4126, n_1766, n4125);
  and g6583 (n4127, n_2230, n4125);
  not g6584 (n_2531, n4126);
  not g6585 (n_2532, n4127);
  and g6586 (n4128, n_2531, n_2532);
  not g6587 (n_2533, n4128);
  and g6588 (n4129, n275, n_2533);
  and g6589 (n4130, n_160, n4128);
  not g6590 (n_2534, n4129);
  not g6591 (n_2535, n4130);
  and g6592 (n4131, n_2534, n_2535);
  and g6593 (n4132, n4120, n4131);
  not g6594 (n_2536, n4132);
  and g6595 (n4133, n4120, n_2536);
  and g6596 (n4134, n4131, n_2536);
  not g6597 (n_2537, n4133);
  not g6598 (n_2538, n4134);
  and g6599 (n4135, n_2537, n_2538);
  not g6600 (n_2539, n4063);
  not g6601 (n_2540, n4135);
  and g6602 (n4136, n_2539, n_2540);
  not g6603 (n_2541, n4136);
  and g6604 (n4137, n_2539, n_2541);
  and g6605 (n4138, n_2540, n_2541);
  not g6606 (n_2542, n4137);
  not g6607 (n_2543, n4138);
  and g6608 (n4139, n_2542, n_2543);
  not g6609 (n_2544, n4062);
  not g6610 (n_2545, n4139);
  and g6611 (n4140, n_2544, n_2545);
  not g6612 (n_2546, n4140);
  and g6613 (n4141, n_2544, n_2546);
  and g6614 (n4142, n_2545, n_2546);
  not g6615 (n_2547, n4141);
  not g6616 (n_2548, n4142);
  and g6617 (n4143, n_2547, n_2548);
  not g6618 (n_2549, n4049);
  and g6619 (n4144, n_2549, n4143);
  not g6620 (n_2550, n4143);
  and g6621 (n4145, n4049, n_2550);
  not g6622 (n_2551, n4144);
  not g6623 (n_2552, n4145);
  and g6624 (n4146, n_2551, n_2552);
  not g6625 (n_2553, n4048);
  not g6626 (n_2554, n4146);
  and g6627 (n4147, n_2553, n_2554);
  and g6628 (n4148, n4048, n4146);
  not g6629 (n_2555, n4032);
  not g6630 (n_2556, n4148);
  and g6631 (n4149, n_2555, n_2556);
  not g6632 (n_2557, n4147);
  and g6633 (n4150, n_2557, n4149);
  not g6634 (n_2558, n4150);
  and g6635 (n4151, n_2555, n_2558);
  and g6636 (n4152, n_2557, n_2558);
  and g6637 (n4153, n_2556, n4152);
  not g6638 (n_2559, n4151);
  not g6639 (n_2560, n4153);
  and g6640 (n4154, n_2559, n_2560);
  and g6641 (n4155, n_2461, n4154);
  not g6642 (n_2561, n4154);
  and g6643 (n4156, n4022, n_2561);
  not g6644 (n_2562, n4155);
  not g6645 (n_2563, n4156);
  and g6646 (n4157, n_2562, n_2563);
  not g6647 (n_2564, \sin[0] );
  and g6648 (n4158, n_2564, n_2469);
  not g6649 (n_2565, n4158);
  and g6650 (n4159, n_2468, n_2565);
  not g6651 (n_2566, n4157);
  and g6652 (n4160, n_2566, n4159);
  not g6653 (n_2567, n4159);
  and g6654 (n4161, n4157, n_2567);
  or g6655 (\sin[2] , n4160, n4161);
  and g6669 (n4176, n_2549, n_2550);
  not g6670 (n_2568, n4176);
  and g6671 (n4177, n_2546, n_2568);
  and g6672 (n4178, n_2536, n_2541);
  and g6673 (n4179, n3274, n3896);
  and g6674 (n4180, n3216, n4054);
  not g6675 (n_2569, n4179);
  not g6676 (n_2570, n4180);
  and g6677 (n4181, n_2569, n_2570);
  not g6678 (n_2571, n4181);
  and g6679 (n4182, n_171, n_2571);
  not g6680 (n_2572, n4182);
  and g6681 (n4183, n_2571, n_2572);
  and g6682 (n4184, n_171, n_2572);
  not g6683 (n_2573, n4183);
  not g6684 (n_2574, n4184);
  and g6685 (n4185, n_2573, n_2574);
  and g6686 (n4186, n2802, n_1931);
  and g6687 (n4187, n_1359, n2808);
  and g6688 (n4188, n2810, n3277);
  and g6694 (n4191, n2817, n3318);
  not g6697 (n_2579, n4192);
  and g6698 (n4193, n_404, n_2579);
  not g6699 (n_2580, n4193);
  and g6700 (n4194, n_2579, n_2580);
  and g6701 (n4195, n_404, n_2580);
  not g6702 (n_2581, n4194);
  not g6703 (n_2582, n4195);
  and g6704 (n4196, n_2581, n_2582);
  and g6705 (n4197, n_2511, n_2516);
  and g6706 (n4198, n_240, n4085);
  and g6707 (n4199, n2593, n4198);
  not g6708 (n_2583, n4199);
  and g6709 (n4200, n_2499, n_2583);
  and g6710 (n4201, n2578, n2668);
  and g6711 (n4202, n_1382, n2776);
  and g6712 (n4203, n_1379, n2666);
  and g6718 (n4206, n2674, n2815);
  and g6721 (n4208, n_240, n2590);
  not g6722 (n_2588, n4207);
  and g6723 (n4209, n_2588, n4208);
  not g6724 (n_2589, n4208);
  and g6725 (n4210, n4207, n_2589);
  not g6726 (n_2590, n4209);
  not g6727 (n_2591, n4210);
  and g6728 (n4211, n_2590, n_2591);
  not g6729 (n_2592, n4200);
  and g6730 (n4212, n_2592, n4211);
  not g6731 (n_2593, n4212);
  and g6732 (n4213, n_2592, n_2593);
  and g6733 (n4214, n4211, n_2593);
  not g6734 (n_2594, n4213);
  not g6735 (n_2595, n4214);
  and g6736 (n4215, n_2594, n_2595);
  and g6737 (n4216, n_1368, n2699);
  and g6738 (n4217, n_1374, n2695);
  and g6739 (n4218, n2562, n2697);
  not g6740 (n_2596, n4217);
  not g6741 (n_2597, n4218);
  and g6742 (n4219, n_2596, n_2597);
  not g6743 (n_2598, n4216);
  and g6744 (n4220, n_2598, n4219);
  and g6745 (n4221, n_1484, n4220);
  not g6746 (n_2599, n3022);
  and g6747 (n4222, n_2599, n4220);
  not g6748 (n_2600, n4221);
  not g6749 (n_2601, n4222);
  and g6750 (n4223, n_2600, n_2601);
  not g6751 (n_2602, n4223);
  and g6752 (n4224, n669, n_2602);
  and g6753 (n4225, n_272, n4223);
  not g6754 (n_2603, n4224);
  not g6755 (n_2604, n4225);
  and g6756 (n4226, n_2603, n_2604);
  not g6757 (n_2605, n4215);
  and g6758 (n4227, n_2605, n4226);
  not g6759 (n_2606, n4226);
  and g6760 (n4228, n4215, n_2606);
  not g6761 (n_2607, n4227);
  not g6762 (n_2608, n4228);
  and g6763 (n4229, n_2607, n_2608);
  not g6764 (n_2609, n4197);
  and g6765 (n4230, n_2609, n4229);
  not g6766 (n_2610, n4229);
  and g6767 (n4231, n4197, n_2610);
  not g6768 (n_2611, n4230);
  not g6769 (n_2612, n4231);
  and g6770 (n4232, n_2611, n_2612);
  not g6771 (n_2613, n4196);
  and g6772 (n4233, n_2613, n4232);
  not g6773 (n_2614, n4233);
  and g6774 (n4234, n_2613, n_2614);
  and g6775 (n4235, n4232, n_2614);
  not g6776 (n_2615, n4234);
  not g6777 (n_2616, n4235);
  and g6778 (n4236, n_2615, n_2616);
  and g6779 (n4237, n_2521, n_2527);
  and g6780 (n4238, n4236, n4237);
  not g6781 (n_2617, n4236);
  not g6782 (n_2618, n4237);
  and g6783 (n4239, n_2617, n_2618);
  not g6784 (n_2619, n4238);
  not g6785 (n_2620, n4239);
  and g6786 (n4240, n_2619, n_2620);
  and g6787 (n4241, n295, n3750);
  and g6788 (n4242, n2560, n3272);
  and g6789 (n4243, n2567, n_2220);
  not g6790 (n_2621, n4242);
  not g6791 (n_2622, n4243);
  and g6792 (n4244, n_2621, n_2622);
  not g6793 (n_2623, n4241);
  and g6794 (n4245, n_2623, n4244);
  and g6795 (n4246, n_1766, n4245);
  not g6796 (n_2624, n3762);
  and g6797 (n4247, n_2624, n4245);
  not g6798 (n_2625, n4246);
  not g6799 (n_2626, n4247);
  and g6800 (n4248, n_2625, n_2626);
  not g6801 (n_2627, n4248);
  and g6802 (n4249, n275, n_2627);
  and g6803 (n4250, n_160, n4248);
  not g6804 (n_2628, n4249);
  not g6805 (n_2629, n4250);
  and g6806 (n4251, n_2628, n_2629);
  and g6807 (n4252, n4240, n4251);
  not g6808 (n_2630, n4240);
  not g6809 (n_2631, n4251);
  and g6810 (n4253, n_2630, n_2631);
  not g6811 (n_2632, n4252);
  not g6812 (n_2633, n4253);
  and g6813 (n4254, n_2632, n_2633);
  not g6814 (n_2634, n4185);
  and g6815 (n4255, n_2634, n4254);
  not g6816 (n_2635, n4254);
  and g6817 (n4256, n4185, n_2635);
  not g6818 (n_2636, n4255);
  not g6819 (n_2637, n4256);
  and g6820 (n4257, n_2636, n_2637);
  not g6821 (n_2638, n4178);
  and g6822 (n4258, n_2638, n4257);
  not g6823 (n_2639, n4257);
  and g6824 (n4259, n4178, n_2639);
  not g6825 (n_2640, n4258);
  not g6826 (n_2641, n4259);
  and g6827 (n4260, n_2640, n_2641);
  not g6828 (n_2642, n4177);
  and g6829 (n4261, n_2642, n4260);
  not g6830 (n_2643, n4260);
  and g6831 (n4262, n4177, n_2643);
  not g6832 (n_2644, n4261);
  not g6833 (n_2645, n4262);
  and g6834 (n4263, n_2644, n_2645);
  not g6835 (n_2646, n4175);
  and g6836 (n4264, n_2646, n4263);
  not g6837 (n_2647, n4264);
  and g6838 (n4265, n_2646, n_2647);
  and g6839 (n4266, n4263, n_2647);
  not g6840 (n_2648, n4265);
  not g6841 (n_2649, n4266);
  and g6842 (n4267, n_2648, n_2649);
  not g6843 (n_2650, n4152);
  not g6844 (n_2651, n4267);
  and g6845 (n4268, n_2650, n_2651);
  and g6846 (n4269, n4152, n_2649);
  and g6847 (n4270, n_2648, n4269);
  not g6848 (n_2652, n4268);
  not g6849 (n_2653, n4270);
  and g6850 (n4271, n_2652, n_2653);
  and g6851 (n4272, n4156, n4271);
  not g6852 (n_2654, n4272);
  and g6853 (n4273, n4271, n_2654);
  and g6854 (n4274, n4156, n_2654);
  not g6855 (n_2655, n4273);
  not g6856 (n_2656, n4274);
  and g6857 (n4275, n_2655, n_2656);
  and g6858 (n4276, n_2566, n4158);
  not g6859 (n_2657, n4276);
  and g6860 (n4277, n_2468, n_2657);
  not g6861 (n_2658, n4275);
  and g6862 (n4278, n_2658, n4277);
  not g6863 (n_2659, n4277);
  and g6864 (n4279, n4275, n_2659);
  not g6865 (n_2660, n4278);
  not g6866 (n_2661, n4279);
  and g6867 (\sin[3] , n_2660, n_2661);
  and g6868 (n4281, n_2647, n_2652);
  and g6879 (n4292, n_2640, n_2644);
  and g6880 (n4293, n_2632, n_2636);
  and g6881 (n4294, n_2614, n_2620);
  and g6882 (n4295, n_2607, n_2611);
  and g6883 (n4296, n_1374, n2668);
  and g6884 (n4297, n_1379, n2776);
  and g6885 (n4298, n2578, n2666);
  and g6891 (n4301, n2674, n2989);
  not g6894 (n_2666, n4302);
  and g6895 (n4303, n_240, n_2666);
  not g6896 (n_2667, n4303);
  and g6897 (n4304, n_2666, n_2667);
  and g6898 (n4305, n_240, n_2667);
  not g6899 (n_2668, n4304);
  not g6900 (n_2669, n4305);
  and g6901 (n4306, n_2668, n_2669);
  and g6902 (n4307, n_171, n_240);
  and g6903 (n4308, n_1382, n4307);
  not g6904 (n_2670, n4308);
  and g6905 (n4309, n_171, n_2670);
  and g6906 (n4310, n_1382, n_2670);
  and g6907 (n4311, n_240, n4310);
  not g6908 (n_2671, n4309);
  not g6909 (n_2672, n4311);
  and g6910 (n4312, n_2671, n_2672);
  not g6911 (n_2673, n4306);
  not g6912 (n_2674, n4312);
  and g6913 (n4313, n_2673, n_2674);
  not g6914 (n_2675, n4313);
  and g6915 (n4314, n_2673, n_2675);
  and g6916 (n4315, n_2674, n_2675);
  not g6917 (n_2676, n4314);
  not g6918 (n_2677, n4315);
  and g6919 (n4316, n_2676, n_2677);
  and g6920 (n4317, n_240, n_1385);
  and g6921 (n4318, n4207, n4317);
  not g6922 (n_2678, n4318);
  and g6923 (n4319, n_2593, n_2678);
  not g6924 (n_2679, n4319);
  and g6925 (n4320, n4316, n_2679);
  not g6926 (n_2680, n4316);
  and g6927 (n4321, n_2680, n4319);
  not g6928 (n_2681, n4320);
  not g6929 (n_2682, n4321);
  and g6930 (n4322, n_2681, n_2682);
  and g6931 (n4323, n_1359, n2699);
  and g6932 (n4324, n2562, n2695);
  and g6933 (n4325, n_1368, n2697);
  and g6939 (n4328, n2652, n2690);
  not g6942 (n_2687, n4329);
  and g6943 (n4330, n_272, n_2687);
  and g6944 (n4331, n669, n4329);
  not g6945 (n_2688, n4330);
  not g6946 (n_2689, n4331);
  and g6947 (n4332, n_2688, n_2689);
  not g6948 (n_2690, n4322);
  and g6949 (n4333, n_2690, n4332);
  not g6950 (n_2691, n4333);
  and g6951 (n4334, n_2690, n_2691);
  and g6952 (n4335, n4332, n_2691);
  not g6953 (n_2692, n4334);
  not g6954 (n_2693, n4335);
  and g6955 (n4336, n_2692, n_2693);
  not g6956 (n_2694, n4295);
  and g6957 (n4337, n_2694, n4336);
  not g6958 (n_2695, n4336);
  and g6959 (n4338, n4295, n_2695);
  not g6960 (n_2696, n4337);
  not g6961 (n_2697, n4338);
  and g6962 (n4339, n_2696, n_2697);
  and g6963 (n4340, n2802, n3272);
  and g6964 (n4341, n2808, n3277);
  and g6965 (n4342, n2810, n_1931);
  and g6971 (n4345, n2817, n3302);
  not g6974 (n_2702, n4346);
  and g6975 (n4347, n_404, n_2702);
  not g6976 (n_2703, n4347);
  and g6977 (n4348, n_404, n_2703);
  and g6978 (n4349, n_2702, n_2703);
  not g6979 (n_2704, n4348);
  not g6980 (n_2705, n4349);
  and g6981 (n4350, n_2704, n_2705);
  not g6982 (n_2706, n4339);
  not g6983 (n_2707, n4350);
  and g6984 (n4351, n_2706, n_2707);
  and g6985 (n4352, n4339, n4350);
  not g6986 (n_2708, n4351);
  not g6987 (n_2709, n4352);
  and g6988 (n4353, n_2708, n_2709);
  not g6989 (n_2710, n4294);
  and g6990 (n4354, n_2710, n4353);
  not g6991 (n_2711, n4353);
  and g6992 (n4355, n4294, n_2711);
  not g6993 (n_2712, n4354);
  not g6994 (n_2713, n4355);
  and g6995 (n4356, n_2712, n_2713);
  and g6996 (n4357, n295, n3896);
  and g6997 (n4358, n2560, n_2220);
  and g6998 (n4359, n2567, n3750);
  and g7004 (n4362, n2571, n3908);
  not g7007 (n_2718, n4363);
  and g7008 (n4364, n_160, n_2718);
  and g7009 (n4365, n275, n4363);
  not g7010 (n_2719, n4364);
  not g7011 (n_2720, n4365);
  and g7012 (n4366, n_2719, n_2720);
  and g7013 (n4367, n4356, n4366);
  not g7014 (n_2721, n4356);
  not g7015 (n_2722, n4366);
  and g7016 (n4368, n_2721, n_2722);
  not g7017 (n_2723, n4367);
  not g7018 (n_2724, n4368);
  and g7019 (n4369, n_2723, n_2724);
  not g7020 (n_2725, n4293);
  and g7021 (n4370, n_2725, n4369);
  not g7022 (n_2726, n4369);
  and g7023 (n4371, n4293, n_2726);
  not g7024 (n_2727, n4370);
  not g7025 (n_2728, n4371);
  and g7026 (n4372, n_2727, n_2728);
  not g7027 (n_2729, n4372);
  and g7028 (n4373, n4292, n_2729);
  not g7029 (n_2730, n4292);
  and g7030 (n4374, n_2730, n4372);
  not g7031 (n_2731, n4373);
  not g7032 (n_2732, n4374);
  and g7033 (n4375, n_2731, n_2732);
  not g7034 (n_2733, n4375);
  and g7035 (n4376, n4291, n_2733);
  not g7036 (n_2734, n4291);
  and g7037 (n4377, n_2734, n4375);
  not g7038 (n_2735, n4376);
  not g7039 (n_2736, n4377);
  and g7040 (n4378, n_2735, n_2736);
  not g7041 (n_2737, n4281);
  and g7042 (n4379, n_2737, n4378);
  not g7043 (n_2738, n4378);
  and g7044 (n4380, n4281, n_2738);
  not g7045 (n_2739, n4379);
  not g7046 (n_2740, n4380);
  and g7047 (n4381, n_2739, n_2740);
  not g7048 (n_2741, n4381);
  and g7049 (n4382, n_2654, n_2741);
  and g7050 (n4383, n4272, n4381);
  not g7051 (n_2742, n4382);
  not g7052 (n_2743, n4383);
  and g7053 (n4384, n_2742, n_2743);
  and g7054 (n4385, n4275, n4276);
  not g7055 (n_2744, n4385);
  and g7056 (n4386, n_2468, n_2744);
  not g7057 (n_2745, n4384);
  and g7058 (n4387, n_2745, n4386);
  not g7059 (n_2746, n4386);
  and g7060 (n4388, n4384, n_2746);
  or g7061 (\sin[4] , n4387, n4388);
  and g7062 (n4390, n_2736, n_2739);
  and g7063 (n4391, n_184, n_202);
  and g7064 (n4392, n_220, n4391);
  and g7077 (n4405, n_2727, n_2732);
  and g7078 (n4406, n_2712, n_2723);
  and g7079 (n4407, n_2694, n_2695);
  not g7080 (n_2747, n4407);
  and g7081 (n4408, n_2708, n_2747);
  and g7082 (n4409, n2802, n_2220);
  and g7083 (n4410, n2808, n_1931);
  and g7084 (n4411, n2810, n3272);
  and g7090 (n4414, n2817, n3641);
  not g7093 (n_2752, n4415);
  and g7094 (n4416, n_404, n_2752);
  not g7095 (n_2753, n4416);
  and g7096 (n4417, n_2752, n_2753);
  and g7097 (n4418, n_404, n_2753);
  not g7098 (n_2754, n4417);
  not g7099 (n_2755, n4418);
  and g7100 (n4419, n_2754, n_2755);
  and g7101 (n4420, n_2680, n_2679);
  not g7102 (n_2756, n4420);
  and g7103 (n4421, n_2691, n_2756);
  and g7104 (n4422, n_2670, n_2675);
  and g7105 (n4423, n_1379, n4307);
  not g7106 (n_2757, n4423);
  and g7107 (n4424, n_171, n_2757);
  and g7108 (n4425, n_1379, n_2757);
  and g7109 (n4426, n_240, n4425);
  not g7110 (n_2758, n4424);
  not g7111 (n_2759, n4426);
  and g7112 (n4427, n_2758, n_2759);
  not g7113 (n_2760, n4422);
  not g7114 (n_2761, n4427);
  and g7115 (n4428, n_2760, n_2761);
  not g7116 (n_2762, n4428);
  and g7117 (n4429, n_2760, n_2762);
  and g7118 (n4430, n_2761, n_2762);
  not g7119 (n_2763, n4429);
  not g7120 (n_2764, n4430);
  and g7121 (n4431, n_2763, n_2764);
  and g7122 (n4432, n2562, n2668);
  and g7123 (n4433, n2578, n2776);
  and g7124 (n4434, n_1374, n2666);
  not g7125 (n_2765, n4433);
  not g7126 (n_2766, n4434);
  and g7127 (n4435, n_2765, n_2766);
  not g7128 (n_2767, n4432);
  and g7129 (n4436, n_2767, n4435);
  and g7130 (n4437, n_1543, n4436);
  and g7131 (n4438, n_1769, n4436);
  not g7132 (n_2768, n4437);
  not g7133 (n_2769, n4438);
  and g7134 (n4439, n_2768, n_2769);
  not g7135 (n_2770, n4439);
  and g7136 (n4440, n525, n_2770);
  and g7137 (n4441, n_240, n4439);
  not g7138 (n_2771, n4440);
  not g7139 (n_2772, n4441);
  and g7140 (n4442, n_2771, n_2772);
  not g7141 (n_2773, n4431);
  and g7142 (n4443, n_2773, n4442);
  not g7143 (n_2774, n4443);
  and g7144 (n4444, n_2773, n_2774);
  and g7145 (n4445, n4442, n_2774);
  not g7146 (n_2775, n4444);
  not g7147 (n_2776, n4445);
  and g7148 (n4446, n_2775, n_2776);
  and g7149 (n4447, n2699, n3277);
  and g7150 (n4448, n_1368, n2695);
  and g7151 (n4449, n_1359, n2697);
  and g7157 (n4452, n2690, n3332);
  not g7160 (n_2781, n4453);
  and g7161 (n4454, n_272, n_2781);
  and g7162 (n4455, n669, n4453);
  not g7163 (n_2782, n4454);
  not g7164 (n_2783, n4455);
  and g7165 (n4456, n_2782, n_2783);
  not g7166 (n_2784, n4446);
  and g7167 (n4457, n_2784, n4456);
  not g7168 (n_2785, n4456);
  and g7169 (n4458, n_2776, n_2785);
  and g7170 (n4459, n_2775, n4458);
  not g7171 (n_2786, n4457);
  not g7172 (n_2787, n4459);
  and g7173 (n4460, n_2786, n_2787);
  not g7174 (n_2788, n4421);
  and g7175 (n4461, n_2788, n4460);
  not g7176 (n_2789, n4461);
  and g7177 (n4462, n_2788, n_2789);
  and g7178 (n4463, n4460, n_2789);
  not g7179 (n_2790, n4462);
  not g7180 (n_2791, n4463);
  and g7181 (n4464, n_2790, n_2791);
  not g7182 (n_2792, n4419);
  not g7183 (n_2793, n4464);
  and g7184 (n4465, n_2792, n_2793);
  and g7185 (n4466, n4419, n_2791);
  and g7186 (n4467, n_2790, n4466);
  not g7187 (n_2794, n4465);
  not g7188 (n_2795, n4467);
  and g7189 (n4468, n_2794, n_2795);
  not g7190 (n_2796, n4408);
  and g7191 (n4469, n_2796, n4468);
  not g7192 (n_2797, n4469);
  and g7193 (n4470, n_2796, n_2797);
  and g7194 (n4471, n4468, n_2797);
  not g7195 (n_2798, n4470);
  not g7196 (n_2799, n4471);
  and g7197 (n4472, n_2798, n_2799);
  and g7198 (n4473, n2560, n3750);
  and g7199 (n4474, n2567, n3896);
  not g7200 (n_2800, n4473);
  not g7201 (n_2801, n4474);
  and g7202 (n4475, n_2800, n_2801);
  and g7203 (n4476, n2571, n4056);
  not g7204 (n_2802, n4476);
  and g7205 (n4477, n4475, n_2802);
  not g7206 (n_2803, n4477);
  and g7207 (n4478, n_160, n_2803);
  and g7208 (n4479, n275, n4477);
  not g7209 (n_2804, n4478);
  not g7210 (n_2805, n4479);
  and g7211 (n4480, n_2804, n_2805);
  not g7212 (n_2806, n4472);
  and g7213 (n4481, n_2806, n4480);
  not g7214 (n_2807, n4480);
  and g7215 (n4482, n_2799, n_2807);
  and g7216 (n4483, n_2798, n4482);
  not g7217 (n_2808, n4481);
  not g7218 (n_2809, n4483);
  and g7219 (n4484, n_2808, n_2809);
  not g7220 (n_2810, n4406);
  and g7221 (n4485, n_2810, n4484);
  not g7222 (n_2811, n4484);
  and g7223 (n4486, n4406, n_2811);
  not g7224 (n_2812, n4485);
  not g7225 (n_2813, n4486);
  and g7226 (n4487, n_2812, n_2813);
  not g7227 (n_2814, n4405);
  and g7228 (n4488, n_2814, n4487);
  not g7229 (n_2815, n4487);
  and g7230 (n4489, n4405, n_2815);
  not g7231 (n_2816, n4488);
  not g7232 (n_2817, n4489);
  and g7233 (n4490, n_2816, n_2817);
  not g7234 (n_2818, n4490);
  and g7235 (n4491, n4404, n_2818);
  not g7236 (n_2819, n4404);
  and g7237 (n4492, n_2819, n4490);
  not g7238 (n_2820, n4491);
  not g7239 (n_2821, n4492);
  and g7240 (n4493, n_2820, n_2821);
  not g7241 (n_2822, n4390);
  and g7242 (n4494, n_2822, n4493);
  not g7243 (n_2823, n4493);
  and g7244 (n4495, n4390, n_2823);
  not g7245 (n_2824, n4494);
  not g7246 (n_2825, n4495);
  and g7247 (n4496, n_2824, n_2825);
  not g7248 (n_2826, n4496);
  and g7249 (n4497, n_2743, n_2826);
  and g7250 (n4498, n4383, n4496);
  not g7251 (n_2827, n4497);
  not g7252 (n_2828, n4498);
  and g7253 (n4499, n_2827, n_2828);
  and g7254 (n4500, n_2745, n4385);
  not g7255 (n_2829, n4500);
  and g7256 (n4501, n_2468, n_2829);
  not g7257 (n_2830, n4499);
  and g7258 (n4502, n_2830, n4501);
  not g7259 (n_2831, n4501);
  and g7260 (n4503, n4499, n_2831);
  or g7261 (\sin[5] , n4502, n4503);
  and g7262 (n4505, n_2821, n_2824);
  and g7281 (n4524, n_2812, n_2816);
  and g7282 (n4525, n_2797, n_2808);
  and g7283 (n4526, n_2789, n_2794);
  and g7284 (n4527, n2560, n3896);
  and g7285 (n4528, n2571, n4054);
  not g7286 (n_2832, n4527);
  not g7287 (n_2833, n4528);
  and g7288 (n4529, n_2832, n_2833);
  not g7289 (n_2834, n4529);
  and g7290 (n4530, n275, n_2834);
  and g7291 (n4531, n_160, n4529);
  not g7292 (n_2835, n4530);
  not g7293 (n_2836, n4531);
  and g7294 (n4532, n_2835, n_2836);
  not g7295 (n_2837, n4526);
  not g7296 (n_2838, n4532);
  and g7297 (n4533, n_2837, n_2838);
  and g7298 (n4534, n4526, n4532);
  not g7299 (n_2839, n4533);
  not g7300 (n_2840, n4534);
  and g7301 (n4535, n_2839, n_2840);
  and g7302 (n4536, n2802, n3750);
  and g7303 (n4537, n2808, n3272);
  and g7304 (n4538, n2810, n_2220);
  and g7310 (n4541, n2817, n3762);
  not g7313 (n_2845, n4542);
  and g7314 (n4543, n_404, n_2845);
  not g7315 (n_2846, n4543);
  and g7316 (n4544, n_2845, n_2846);
  and g7317 (n4545, n_404, n_2846);
  not g7318 (n_2847, n4544);
  not g7319 (n_2848, n4545);
  and g7320 (n4546, n_2847, n_2848);
  and g7321 (n4547, n_2774, n_2786);
  and g7322 (n4548, n_2757, n_2762);
  and g7323 (n4549, n2578, n4307);
  not g7324 (n_2849, n4549);
  and g7325 (n4550, n_171, n_2849);
  and g7326 (n4551, n2578, n_2849);
  and g7327 (n4552, n_240, n4551);
  not g7328 (n_2850, n4550);
  not g7329 (n_2851, n4552);
  and g7330 (n4553, n_2850, n_2851);
  not g7331 (n_2852, n4548);
  not g7332 (n_2853, n4553);
  and g7333 (n4554, n_2852, n_2853);
  not g7334 (n_2854, n4554);
  and g7335 (n4555, n_2852, n_2854);
  and g7336 (n4556, n_2853, n_2854);
  not g7337 (n_2855, n4555);
  not g7338 (n_2856, n4556);
  and g7339 (n4557, n_2855, n_2856);
  and g7340 (n4558, n_1368, n2668);
  and g7341 (n4559, n_1374, n2776);
  and g7342 (n4560, n2562, n2666);
  not g7343 (n_2857, n4559);
  not g7344 (n_2858, n4560);
  and g7345 (n4561, n_2857, n_2858);
  not g7346 (n_2859, n4558);
  and g7347 (n4562, n_2859, n4561);
  and g7348 (n4563, n_1543, n4562);
  and g7349 (n4564, n_2599, n4562);
  not g7350 (n_2860, n4563);
  not g7351 (n_2861, n4564);
  and g7352 (n4565, n_2860, n_2861);
  not g7353 (n_2862, n4565);
  and g7354 (n4566, n525, n_2862);
  and g7355 (n4567, n_240, n4565);
  not g7356 (n_2863, n4566);
  not g7357 (n_2864, n4567);
  and g7358 (n4568, n_2863, n_2864);
  not g7359 (n_2865, n4557);
  and g7360 (n4569, n_2865, n4568);
  not g7361 (n_2866, n4569);
  and g7362 (n4570, n_2865, n_2866);
  and g7363 (n4571, n4568, n_2866);
  not g7364 (n_2867, n4570);
  not g7365 (n_2868, n4571);
  and g7366 (n4572, n_2867, n_2868);
  and g7367 (n4573, n2699, n_1931);
  and g7368 (n4574, n_1359, n2695);
  and g7369 (n4575, n2697, n3277);
  and g7375 (n4578, n2690, n3318);
  not g7378 (n_2873, n4579);
  and g7379 (n4580, n_272, n_2873);
  and g7380 (n4581, n669, n4579);
  not g7381 (n_2874, n4580);
  not g7382 (n_2875, n4581);
  and g7383 (n4582, n_2874, n_2875);
  not g7384 (n_2876, n4572);
  and g7385 (n4583, n_2876, n4582);
  not g7386 (n_2877, n4582);
  and g7387 (n4584, n_2868, n_2877);
  and g7388 (n4585, n_2867, n4584);
  not g7389 (n_2878, n4583);
  not g7390 (n_2879, n4585);
  and g7391 (n4586, n_2878, n_2879);
  not g7392 (n_2880, n4547);
  and g7393 (n4587, n_2880, n4586);
  not g7394 (n_2881, n4587);
  and g7395 (n4588, n_2880, n_2881);
  and g7396 (n4589, n4586, n_2881);
  not g7397 (n_2882, n4588);
  not g7398 (n_2883, n4589);
  and g7399 (n4590, n_2882, n_2883);
  not g7400 (n_2884, n4546);
  not g7401 (n_2885, n4590);
  and g7402 (n4591, n_2884, n_2885);
  and g7403 (n4592, n4546, n_2883);
  and g7404 (n4593, n_2882, n4592);
  not g7405 (n_2886, n4591);
  not g7406 (n_2887, n4593);
  and g7407 (n4594, n_2886, n_2887);
  and g7408 (n4595, n4535, n4594);
  not g7409 (n_2888, n4535);
  not g7410 (n_2889, n4594);
  and g7411 (n4596, n_2888, n_2889);
  not g7412 (n_2890, n4595);
  not g7413 (n_2891, n4596);
  and g7414 (n4597, n_2890, n_2891);
  not g7415 (n_2892, n4525);
  and g7416 (n4598, n_2892, n4597);
  not g7417 (n_2893, n4597);
  and g7418 (n4599, n4525, n_2893);
  not g7419 (n_2894, n4598);
  not g7420 (n_2895, n4599);
  and g7421 (n4600, n_2894, n_2895);
  not g7422 (n_2896, n4524);
  and g7423 (n4601, n_2896, n4600);
  not g7424 (n_2897, n4600);
  and g7425 (n4602, n4524, n_2897);
  not g7426 (n_2898, n4601);
  not g7427 (n_2899, n4602);
  and g7428 (n4603, n_2898, n_2899);
  not g7429 (n_2900, n4603);
  and g7430 (n4604, n4523, n_2900);
  not g7431 (n_2901, n4523);
  and g7432 (n4605, n_2901, n4603);
  not g7433 (n_2902, n4604);
  not g7434 (n_2903, n4605);
  and g7435 (n4606, n_2902, n_2903);
  not g7436 (n_2904, n4505);
  and g7437 (n4607, n_2904, n4606);
  not g7438 (n_2905, n4606);
  and g7439 (n4608, n4505, n_2905);
  not g7440 (n_2906, n4607);
  not g7441 (n_2907, n4608);
  and g7442 (n4609, n_2906, n_2907);
  not g7443 (n_2908, n4609);
  and g7444 (n4610, n_2828, n_2908);
  and g7445 (n4611, n4498, n4609);
  not g7446 (n_2909, n4610);
  not g7447 (n_2910, n4611);
  and g7448 (n4612, n_2909, n_2910);
  and g7449 (n4613, n_2830, n4500);
  not g7450 (n_2911, n4613);
  and g7451 (n4614, n_2468, n_2911);
  not g7452 (n_2912, n4612);
  and g7453 (n4615, n_2912, n4614);
  not g7454 (n_2913, n4614);
  and g7455 (n4616, n4612, n_2913);
  or g7456 (\sin[6] , n4615, n4616);
  and g7457 (n4618, n_2903, n_2906);
  and g7458 (n4619, n_2839, n_2890);
  and g7459 (n4620, n_2881, n_2886);
  and g7460 (n4621, n2802, n3896);
  and g7461 (n4622, n2808, n_2220);
  and g7462 (n4623, n2810, n3750);
  not g7463 (n_2914, n4622);
  not g7464 (n_2915, n4623);
  and g7465 (n4624, n_2914, n_2915);
  not g7466 (n_2916, n4621);
  and g7467 (n4625, n_2916, n4624);
  not g7468 (n_2917, n3908);
  and g7469 (n4626, n_2917, n4625);
  and g7470 (n4627, n_1575, n4625);
  not g7471 (n_2918, n4626);
  not g7472 (n_2919, n4627);
  and g7473 (n4628, n_2918, n_2919);
  not g7474 (n_2920, n4628);
  and g7475 (n4629, n1021, n_2920);
  and g7476 (n4630, n_404, n4628);
  not g7477 (n_2921, n4629);
  not g7478 (n_2922, n4630);
  and g7479 (n4631, n_2921, n_2922);
  not g7480 (n_2923, n4620);
  and g7481 (n4632, n_2923, n4631);
  not g7482 (n_2924, n4631);
  and g7483 (n4633, n4620, n_2924);
  not g7484 (n_2925, n4632);
  not g7485 (n_2926, n4633);
  and g7486 (n4634, n_2925, n_2926);
  and g7487 (n4635, n_2866, n_2878);
  and g7488 (n4636, n_2849, n_2854);
  and g7489 (n4637, n_1359, n2668);
  and g7490 (n4638, n2562, n2776);
  and g7491 (n4639, n_1368, n2666);
  and g7497 (n4642, n2652, n2674);
  not g7500 (n_2931, n4643);
  and g7501 (n4644, n_240, n_2931);
  not g7502 (n_2932, n4644);
  and g7503 (n4645, n_2931, n_2932);
  and g7504 (n4646, n_240, n_2932);
  not g7505 (n_2933, n4645);
  not g7506 (n_2934, n4646);
  and g7507 (n4647, n_2933, n_2934);
  and g7508 (n4648, n_240, n_1374);
  and g7509 (n4649, n275, n291);
  and g7510 (n4650, n_160, n_171);
  not g7511 (n_2935, n4649);
  not g7512 (n_2936, n4650);
  and g7513 (n4651, n_2935, n_2936);
  and g7514 (n4652, n4648, n4651);
  not g7515 (n_2937, n4648);
  not g7516 (n_2938, n4651);
  and g7517 (n4653, n_2937, n_2938);
  not g7518 (n_2939, n4652);
  not g7519 (n_2940, n4653);
  and g7520 (n4654, n_2939, n_2940);
  not g7521 (n_2941, n4647);
  and g7522 (n4655, n_2941, n4654);
  not g7523 (n_2942, n4655);
  and g7524 (n4656, n_2941, n_2942);
  and g7525 (n4657, n4654, n_2942);
  not g7526 (n_2943, n4656);
  not g7527 (n_2944, n4657);
  and g7528 (n4658, n_2943, n_2944);
  not g7529 (n_2945, n4636);
  and g7530 (n4659, n_2945, n4658);
  not g7531 (n_2946, n4658);
  and g7532 (n4660, n4636, n_2946);
  not g7533 (n_2947, n4659);
  not g7534 (n_2948, n4660);
  and g7535 (n4661, n_2947, n_2948);
  and g7536 (n4662, n2699, n3272);
  and g7537 (n4663, n2695, n3277);
  and g7538 (n4664, n2697, n_1931);
  not g7539 (n_2949, n4663);
  not g7540 (n_2950, n4664);
  and g7541 (n4665, n_2949, n_2950);
  not g7542 (n_2951, n4662);
  and g7543 (n4666, n_2951, n4665);
  and g7544 (n4667, n_1484, n4666);
  and g7545 (n4668, n_1952, n4666);
  not g7546 (n_2952, n4667);
  not g7547 (n_2953, n4668);
  and g7548 (n4669, n_2952, n_2953);
  not g7549 (n_2954, n4669);
  and g7550 (n4670, n669, n_2954);
  and g7551 (n4671, n_272, n4669);
  not g7552 (n_2955, n4670);
  not g7553 (n_2956, n4671);
  and g7554 (n4672, n_2955, n_2956);
  not g7555 (n_2957, n4661);
  and g7556 (n4673, n_2957, n4672);
  not g7557 (n_2958, n4673);
  and g7558 (n4674, n_2957, n_2958);
  and g7559 (n4675, n4672, n_2958);
  not g7560 (n_2959, n4674);
  not g7561 (n_2960, n4675);
  and g7562 (n4676, n_2959, n_2960);
  not g7563 (n_2961, n4635);
  not g7564 (n_2962, n4676);
  and g7565 (n4677, n_2961, n_2962);
  not g7566 (n_2963, n4677);
  and g7567 (n4678, n_2961, n_2963);
  and g7568 (n4679, n_2962, n_2963);
  not g7569 (n_2964, n4678);
  not g7570 (n_2965, n4679);
  and g7571 (n4680, n_2964, n_2965);
  not g7572 (n_2966, n4680);
  and g7573 (n4681, n4634, n_2966);
  not g7574 (n_2967, n4681);
  and g7575 (n4682, n4634, n_2967);
  and g7576 (n4683, n_2966, n_2967);
  not g7577 (n_2968, n4682);
  not g7578 (n_2969, n4683);
  and g7579 (n4684, n_2968, n_2969);
  not g7580 (n_2970, n4619);
  and g7581 (n4685, n_2970, n4684);
  not g7582 (n_2971, n4684);
  and g7583 (n4686, n4619, n_2971);
  not g7584 (n_2972, n4685);
  not g7585 (n_2973, n4686);
  and g7586 (n4687, n_2972, n_2973);
  and g7587 (n4688, n_2894, n_2898);
  and g7588 (n4689, n4687, n4688);
  not g7589 (n_2974, n4687);
  not g7590 (n_2975, n4688);
  and g7591 (n4690, n_2974, n_2975);
  not g7592 (n_2976, n4689);
  not g7593 (n_2977, n4690);
  and g7594 (n4691, n_2976, n_2977);
  not g7606 (n_2978, n4702);
  and g7607 (n4703, n4691, n_2978);
  not g7608 (n_2979, n4691);
  and g7609 (n4704, n_2979, n4702);
  not g7610 (n_2980, n4703);
  not g7611 (n_2981, n4704);
  and g7612 (n4705, n_2980, n_2981);
  not g7613 (n_2982, n4618);
  and g7614 (n4706, n_2982, n4705);
  not g7615 (n_2983, n4705);
  and g7616 (n4707, n4618, n_2983);
  not g7617 (n_2984, n4706);
  not g7618 (n_2985, n4707);
  and g7619 (n4708, n_2984, n_2985);
  and g7620 (n4709, n4611, n4708);
  not g7621 (n_2986, n4708);
  and g7622 (n4710, n_2910, n_2986);
  not g7623 (n_2987, n4709);
  not g7624 (n_2988, n4710);
  and g7625 (n4711, n_2987, n_2988);
  and g7626 (n4712, n_2912, n4613);
  not g7627 (n_2989, n4712);
  and g7628 (n4713, n_2468, n_2989);
  not g7629 (n_2990, n4711);
  and g7630 (n4714, n_2990, n4713);
  not g7631 (n_2991, n4713);
  and g7632 (n4715, n4711, n_2991);
  or g7633 (\sin[7] , n4714, n4715);
  and g7634 (n4717, n_2980, n_2984);
  and g7655 (n4738, n_2970, n_2971);
  not g7656 (n_2992, n4738);
  and g7657 (n4739, n_2977, n_2992);
  and g7658 (n4740, n_2925, n_2967);
  and g7659 (n4741, n2808, n3750);
  and g7660 (n4742, n2810, n3896);
  not g7661 (n_2993, n4741);
  not g7662 (n_2994, n4742);
  and g7663 (n4743, n_2993, n_2994);
  and g7664 (n4744, n2817, n4056);
  not g7665 (n_2995, n4744);
  and g7666 (n4745, n4743, n_2995);
  not g7667 (n_2996, n4745);
  and g7668 (n4746, n_404, n_2996);
  not g7669 (n_2997, n4746);
  and g7670 (n4747, n_2996, n_2997);
  and g7671 (n4748, n_404, n_2997);
  not g7672 (n_2998, n4747);
  not g7673 (n_2999, n4748);
  and g7674 (n4749, n_2998, n_2999);
  and g7675 (n4750, n_2958, n_2963);
  and g7676 (n4751, n_2945, n_2946);
  not g7677 (n_3000, n4751);
  and g7678 (n4752, n_2942, n_3000);
  and g7679 (n4753, n_240, n2562);
  and g7680 (n4754, n_2935, n_2939);
  not g7681 (n_3001, n4753);
  not g7682 (n_3002, n4754);
  and g7683 (n4755, n_3001, n_3002);
  not g7684 (n_3003, n4755);
  and g7685 (n4756, n_3001, n_3003);
  and g7686 (n4757, n_3002, n_3003);
  not g7687 (n_3004, n4756);
  not g7688 (n_3005, n4757);
  and g7689 (n4758, n_3004, n_3005);
  and g7690 (n4759, n2668, n3277);
  and g7691 (n4760, n_1368, n2776);
  and g7692 (n4761, n_1359, n2666);
  not g7693 (n_3006, n4760);
  not g7694 (n_3007, n4761);
  and g7695 (n4762, n_3006, n_3007);
  not g7696 (n_3008, n4759);
  and g7697 (n4763, n_3008, n4762);
  and g7698 (n4764, n_1543, n4763);
  not g7699 (n_3009, n3332);
  and g7700 (n4765, n_3009, n4763);
  not g7701 (n_3010, n4764);
  not g7702 (n_3011, n4765);
  and g7703 (n4766, n_3010, n_3011);
  not g7704 (n_3012, n4766);
  and g7705 (n4767, n525, n_3012);
  and g7706 (n4768, n_240, n4766);
  not g7707 (n_3013, n4767);
  not g7708 (n_3014, n4768);
  and g7709 (n4769, n_3013, n_3014);
  not g7710 (n_3015, n4758);
  and g7711 (n4770, n_3015, n4769);
  not g7712 (n_3016, n4769);
  and g7713 (n4771, n4758, n_3016);
  not g7714 (n_3017, n4770);
  not g7715 (n_3018, n4771);
  and g7716 (n4772, n_3017, n_3018);
  not g7717 (n_3019, n4752);
  and g7718 (n4773, n_3019, n4772);
  not g7719 (n_3020, n4773);
  and g7720 (n4774, n_3019, n_3020);
  and g7721 (n4775, n4772, n_3020);
  not g7722 (n_3021, n4774);
  not g7723 (n_3022, n4775);
  and g7724 (n4776, n_3021, n_3022);
  and g7725 (n4777, n2699, n_2220);
  and g7726 (n4778, n2695, n_1931);
  and g7727 (n4779, n2697, n3272);
  and g7733 (n4782, n2690, n3641);
  not g7736 (n_3027, n4783);
  and g7737 (n4784, n_272, n_3027);
  and g7738 (n4785, n669, n4783);
  not g7739 (n_3028, n4784);
  not g7740 (n_3029, n4785);
  and g7741 (n4786, n_3028, n_3029);
  not g7742 (n_3030, n4776);
  and g7743 (n4787, n_3030, n4786);
  not g7744 (n_3031, n4786);
  and g7745 (n4788, n_3022, n_3031);
  and g7746 (n4789, n_3021, n4788);
  not g7747 (n_3032, n4787);
  not g7748 (n_3033, n4789);
  and g7749 (n4790, n_3032, n_3033);
  not g7750 (n_3034, n4750);
  and g7751 (n4791, n_3034, n4790);
  not g7752 (n_3035, n4790);
  and g7753 (n4792, n4750, n_3035);
  not g7754 (n_3036, n4791);
  not g7755 (n_3037, n4792);
  and g7756 (n4793, n_3036, n_3037);
  not g7757 (n_3038, n4749);
  and g7758 (n4794, n_3038, n4793);
  not g7759 (n_3039, n4793);
  and g7760 (n4795, n4749, n_3039);
  not g7761 (n_3040, n4794);
  not g7762 (n_3041, n4795);
  and g7763 (n4796, n_3040, n_3041);
  not g7764 (n_3042, n4740);
  and g7765 (n4797, n_3042, n4796);
  not g7766 (n_3043, n4796);
  and g7767 (n4798, n4740, n_3043);
  not g7768 (n_3044, n4797);
  not g7769 (n_3045, n4798);
  and g7770 (n4799, n_3044, n_3045);
  not g7771 (n_3046, n4739);
  and g7772 (n4800, n_3046, n4799);
  not g7773 (n_3047, n4799);
  and g7774 (n4801, n4739, n_3047);
  not g7775 (n_3048, n4800);
  not g7776 (n_3049, n4801);
  and g7777 (n4802, n_3048, n_3049);
  not g7778 (n_3050, n4802);
  and g7779 (n4803, n4737, n_3050);
  not g7780 (n_3051, n4737);
  and g7781 (n4804, n_3051, n4802);
  not g7782 (n_3052, n4803);
  not g7783 (n_3053, n4804);
  and g7784 (n4805, n_3052, n_3053);
  not g7785 (n_3054, n4717);
  and g7786 (n4806, n_3054, n4805);
  not g7787 (n_3055, n4805);
  and g7788 (n4807, n4717, n_3055);
  not g7789 (n_3056, n4806);
  not g7790 (n_3057, n4807);
  and g7791 (n4808, n_3056, n_3057);
  not g7792 (n_3058, n4808);
  and g7793 (n4809, n_2987, n_3058);
  and g7794 (n4810, n4709, n4808);
  not g7795 (n_3059, n4809);
  not g7796 (n_3060, n4810);
  and g7797 (n4811, n_3059, n_3060);
  and g7798 (n4812, n_2990, n4712);
  not g7799 (n_3061, n4812);
  and g7800 (n4813, n_2468, n_3061);
  not g7801 (n_3062, n4811);
  and g7802 (n4814, n_3062, n4813);
  not g7803 (n_3063, n4813);
  and g7804 (n4815, n4811, n_3063);
  or g7805 (\sin[8] , n4814, n4815);
  and g7806 (n4817, n_3053, n_3056);
  and g7819 (n4830, n_3036, n_3040);
  and g7820 (n4831, n_3003, n_3017);
  and g7821 (n4832, n2668, n_1931);
  and g7822 (n4833, n_1359, n2776);
  and g7823 (n4834, n2666, n3277);
  and g7829 (n4837, n2674, n3318);
  not g7832 (n_3068, n4838);
  and g7833 (n4839, n_240, n_3068);
  not g7834 (n_3069, n4839);
  and g7835 (n4840, n_3068, n_3069);
  and g7836 (n4841, n_240, n_3069);
  not g7837 (n_3070, n4840);
  not g7838 (n_3071, n4841);
  and g7839 (n4842, n_3070, n_3071);
  and g7840 (n4843, n_240, n2644);
  not g7841 (n_3072, n4842);
  not g7842 (n_3073, n4843);
  and g7843 (n4844, n_3072, n_3073);
  not g7844 (n_3074, n4844);
  and g7845 (n4845, n_3072, n_3074);
  and g7846 (n4846, n_3073, n_3074);
  not g7847 (n_3075, n4845);
  not g7848 (n_3076, n4846);
  and g7849 (n4847, n_3075, n_3076);
  not g7850 (n_3077, n4831);
  and g7851 (n4848, n_3077, n4847);
  not g7852 (n_3078, n4847);
  and g7853 (n4849, n4831, n_3078);
  not g7854 (n_3079, n4848);
  not g7855 (n_3080, n4849);
  and g7856 (n4850, n_3079, n_3080);
  and g7857 (n4851, n2699, n3750);
  and g7858 (n4852, n2695, n3272);
  and g7859 (n4853, n2697, n_2220);
  and g7865 (n4856, n2690, n3762);
  not g7868 (n_3085, n4857);
  and g7869 (n4858, n_272, n_3085);
  and g7870 (n4859, n669, n4857);
  not g7871 (n_3086, n4858);
  not g7872 (n_3087, n4859);
  and g7873 (n4860, n_3086, n_3087);
  not g7874 (n_3088, n4850);
  and g7875 (n4861, n_3088, n4860);
  not g7876 (n_3089, n4861);
  and g7877 (n4862, n_3088, n_3089);
  and g7878 (n4863, n4860, n_3089);
  not g7879 (n_3090, n4862);
  not g7880 (n_3091, n4863);
  and g7881 (n4864, n_3090, n_3091);
  and g7882 (n4865, n_3020, n_3032);
  and g7883 (n4866, n2808, n3896);
  and g7884 (n4867, n2817, n4054);
  not g7885 (n_3092, n4866);
  not g7886 (n_3093, n4867);
  and g7887 (n4868, n_3092, n_3093);
  and g7888 (n4869, n_404, n4868);
  not g7889 (n_3094, n4868);
  and g7890 (n4870, n1021, n_3094);
  not g7891 (n_3095, n4869);
  not g7892 (n_3096, n4870);
  and g7893 (n4871, n_3095, n_3096);
  not g7894 (n_3097, n4865);
  not g7895 (n_3098, n4871);
  and g7896 (n4872, n_3097, n_3098);
  and g7897 (n4873, n4865, n4871);
  not g7898 (n_3099, n4872);
  not g7899 (n_3100, n4873);
  and g7900 (n4874, n_3099, n_3100);
  not g7901 (n_3101, n4864);
  and g7902 (n4875, n_3101, n4874);
  not g7903 (n_3102, n4875);
  and g7904 (n4876, n_3101, n_3102);
  and g7905 (n4877, n4874, n_3102);
  not g7906 (n_3103, n4876);
  not g7907 (n_3104, n4877);
  and g7908 (n4878, n_3103, n_3104);
  not g7909 (n_3105, n4830);
  and g7910 (n4879, n_3105, n4878);
  not g7911 (n_3106, n4878);
  and g7912 (n4880, n4830, n_3106);
  not g7913 (n_3107, n4879);
  not g7914 (n_3108, n4880);
  and g7915 (n4881, n_3107, n_3108);
  and g7916 (n4882, n_3044, n_3048);
  and g7917 (n4883, n4881, n4882);
  not g7918 (n_3109, n4881);
  not g7919 (n_3110, n4882);
  and g7920 (n4884, n_3109, n_3110);
  not g7921 (n_3111, n4883);
  not g7922 (n_3112, n4884);
  and g7923 (n4885, n_3111, n_3112);
  not g7924 (n_3113, n4885);
  and g7925 (n4886, n4829, n_3113);
  not g7926 (n_3114, n4829);
  and g7927 (n4887, n_3114, n4885);
  not g7928 (n_3115, n4886);
  not g7929 (n_3116, n4887);
  and g7930 (n4888, n_3115, n_3116);
  not g7931 (n_3117, n4817);
  and g7932 (n4889, n_3117, n4888);
  not g7933 (n_3118, n4888);
  and g7934 (n4890, n4817, n_3118);
  not g7935 (n_3119, n4889);
  not g7936 (n_3120, n4890);
  and g7937 (n4891, n_3119, n_3120);
  not g7938 (n_3121, n4891);
  and g7939 (n4892, n_3060, n_3121);
  and g7940 (n4893, n4810, n4891);
  not g7941 (n_3122, n4892);
  not g7942 (n_3123, n4893);
  and g7943 (n4894, n_3122, n_3123);
  and g7944 (n4895, n_3062, n4812);
  not g7945 (n_3124, n4895);
  and g7946 (n4896, n_2468, n_3124);
  not g7947 (n_3125, n4894);
  and g7948 (n4897, n_3125, n4896);
  not g7949 (n_3126, n4896);
  and g7950 (n4898, n4894, n_3126);
  or g7951 (\sin[9] , n4897, n4898);
  and g7952 (n4900, n_3116, n_3119);
  and g7964 (n4912, n_3105, n_3106);
  not g7965 (n_3127, n4912);
  and g7966 (n4913, n_3112, n_3127);
  and g7967 (n4914, n_3099, n_3102);
  and g7968 (n4915, n_1368, n_3001);
  and g7969 (n4916, n_240, n4915);
  not g7970 (n_3128, n4916);
  and g7971 (n4917, n_3074, n_3128);
  and g7972 (n4918, n_240, n_1359);
  not g7973 (n_3129, n4918);
  and g7974 (n4919, n_404, n_3129);
  and g7975 (n4920, n1021, n4918);
  not g7976 (n_3130, n4920);
  and g7977 (n4921, n4753, n_3130);
  not g7978 (n_3131, n4919);
  and g7979 (n4922, n_3131, n4921);
  not g7980 (n_3132, n4922);
  and g7981 (n4923, n4753, n_3132);
  and g7982 (n4924, n_3130, n_3132);
  and g7983 (n4925, n_3131, n4924);
  not g7984 (n_3133, n4923);
  not g7985 (n_3134, n4925);
  and g7986 (n4926, n_3133, n_3134);
  not g7987 (n_3135, n4917);
  not g7988 (n_3136, n4926);
  and g7989 (n4927, n_3135, n_3136);
  not g7990 (n_3137, n4927);
  and g7991 (n4928, n_3135, n_3137);
  and g7992 (n4929, n_3136, n_3137);
  not g7993 (n_3138, n4928);
  not g7994 (n_3139, n4929);
  and g7995 (n4930, n_3138, n_3139);
  and g7996 (n4931, n2668, n3272);
  and g7997 (n4932, n2776, n3277);
  and g7998 (n4933, n2666, n_1931);
  and g8004 (n4936, n2674, n3302);
  not g8007 (n_3144, n4937);
  and g8008 (n4938, n_240, n_3144);
  not g8009 (n_3145, n4938);
  and g8010 (n4939, n_240, n_3145);
  and g8011 (n4940, n_3144, n_3145);
  not g8012 (n_3146, n4939);
  not g8013 (n_3147, n4940);
  and g8014 (n4941, n_3146, n_3147);
  not g8015 (n_3148, n4930);
  not g8016 (n_3149, n4941);
  and g8017 (n4942, n_3148, n_3149);
  not g8018 (n_3150, n4942);
  and g8019 (n4943, n_3148, n_3150);
  and g8020 (n4944, n_3149, n_3150);
  not g8021 (n_3151, n4943);
  not g8022 (n_3152, n4944);
  and g8023 (n4945, n_3151, n_3152);
  and g8024 (n4946, n_3077, n_3078);
  not g8025 (n_3153, n4946);
  and g8026 (n4947, n_3089, n_3153);
  and g8027 (n4948, n2699, n3896);
  and g8028 (n4949, n2695, n_2220);
  and g8029 (n4950, n2697, n3750);
  not g8030 (n_3154, n4949);
  not g8031 (n_3155, n4950);
  and g8032 (n4951, n_3154, n_3155);
  not g8033 (n_3156, n4948);
  and g8034 (n4952, n_3156, n4951);
  and g8035 (n4953, n_1484, n4952);
  and g8036 (n4954, n_2917, n4952);
  not g8037 (n_3157, n4953);
  not g8038 (n_3158, n4954);
  and g8039 (n4955, n_3157, n_3158);
  not g8040 (n_3159, n4955);
  and g8041 (n4956, n669, n_3159);
  and g8042 (n4957, n_272, n4955);
  not g8043 (n_3160, n4956);
  not g8044 (n_3161, n4957);
  and g8045 (n4958, n_3160, n_3161);
  not g8046 (n_3162, n4947);
  and g8047 (n4959, n_3162, n4958);
  not g8048 (n_3163, n4959);
  and g8049 (n4960, n_3162, n_3163);
  and g8050 (n4961, n4958, n_3163);
  not g8051 (n_3164, n4960);
  not g8052 (n_3165, n4961);
  and g8053 (n4962, n_3164, n_3165);
  not g8054 (n_3166, n4945);
  not g8055 (n_3167, n4962);
  and g8056 (n4963, n_3166, n_3167);
  and g8057 (n4964, n4945, n_3165);
  and g8058 (n4965, n_3164, n4964);
  not g8059 (n_3168, n4963);
  not g8060 (n_3169, n4965);
  and g8061 (n4966, n_3168, n_3169);
  not g8062 (n_3170, n4914);
  and g8063 (n4967, n_3170, n4966);
  not g8064 (n_3171, n4966);
  and g8065 (n4968, n4914, n_3171);
  not g8066 (n_3172, n4967);
  not g8067 (n_3173, n4968);
  and g8068 (n4969, n_3172, n_3173);
  not g8069 (n_3174, n4913);
  and g8070 (n4970, n_3174, n4969);
  not g8071 (n_3175, n4969);
  and g8072 (n4971, n4913, n_3175);
  not g8073 (n_3176, n4970);
  not g8074 (n_3177, n4971);
  and g8075 (n4972, n_3176, n_3177);
  not g8076 (n_3178, n4972);
  and g8077 (n4973, n4911, n_3178);
  not g8078 (n_3179, n4911);
  and g8079 (n4974, n_3179, n4972);
  not g8080 (n_3180, n4973);
  not g8081 (n_3181, n4974);
  and g8082 (n4975, n_3180, n_3181);
  not g8083 (n_3182, n4900);
  and g8084 (n4976, n_3182, n4975);
  not g8085 (n_3183, n4975);
  and g8086 (n4977, n4900, n_3183);
  not g8087 (n_3184, n4976);
  not g8088 (n_3185, n4977);
  and g8089 (n4978, n_3184, n_3185);
  not g8090 (n_3186, n4978);
  and g8091 (n4979, n_3123, n_3186);
  and g8092 (n4980, n4893, n4978);
  not g8093 (n_3187, n4979);
  not g8094 (n_3188, n4980);
  and g8095 (n4981, n_3187, n_3188);
  and g8096 (n4982, n_3125, n4895);
  not g8097 (n_3189, n4982);
  and g8098 (n4983, n_2468, n_3189);
  not g8099 (n_3190, n4981);
  and g8100 (n4984, n_3190, n4983);
  not g8101 (n_3191, n4983);
  and g8102 (n4985, n4981, n_3191);
  or g8103 (\sin[10] , n4984, n4985);
  and g8104 (n4987, n_3181, n_3184);
  and g8111 (n4994, n_3172, n_3176);
  and g8112 (n4995, n_3163, n_3168);
  and g8113 (n4996, n_3137, n_3150);
  and g8114 (n4997, n_240, n3277);
  not g8115 (n_3192, n4924);
  and g8116 (n4998, n_3192, n4997);
  not g8117 (n_3193, n4997);
  and g8118 (n4999, n4924, n_3193);
  not g8119 (n_3194, n4998);
  not g8120 (n_3195, n4999);
  and g8121 (n5000, n_3194, n_3195);
  and g8122 (n5001, n2668, n_2220);
  and g8123 (n5002, n2776, n_1931);
  and g8124 (n5003, n2666, n3272);
  not g8125 (n_3196, n5002);
  not g8126 (n_3197, n5003);
  and g8127 (n5004, n_3196, n_3197);
  not g8128 (n_3198, n5001);
  and g8129 (n5005, n_3198, n5004);
  and g8130 (n5006, n_1543, n5005);
  and g8131 (n5007, n_2230, n5005);
  not g8132 (n_3199, n5006);
  not g8133 (n_3200, n5007);
  and g8134 (n5008, n_3199, n_3200);
  not g8135 (n_3201, n5008);
  and g8136 (n5009, n525, n_3201);
  and g8137 (n5010, n_240, n5008);
  not g8138 (n_3202, n5009);
  not g8139 (n_3203, n5010);
  and g8140 (n5011, n_3202, n_3203);
  not g8141 (n_3204, n5000);
  and g8142 (n5012, n_3204, n5011);
  not g8143 (n_3205, n5011);
  and g8144 (n5013, n5000, n_3205);
  not g8145 (n_3206, n5012);
  not g8146 (n_3207, n5013);
  and g8147 (n5014, n_3206, n_3207);
  not g8148 (n_3208, n4996);
  and g8149 (n5015, n_3208, n5014);
  not g8150 (n_3209, n5015);
  and g8151 (n5016, n_3208, n_3209);
  and g8152 (n5017, n5014, n_3209);
  not g8153 (n_3210, n5016);
  not g8154 (n_3211, n5017);
  and g8155 (n5018, n_3210, n_3211);
  and g8156 (n5019, n2695, n3750);
  and g8157 (n5020, n2697, n3896);
  not g8158 (n_3212, n5019);
  not g8159 (n_3213, n5020);
  and g8160 (n5021, n_3212, n_3213);
  and g8161 (n5022, n2690, n4056);
  not g8162 (n_3214, n5022);
  and g8163 (n5023, n5021, n_3214);
  not g8164 (n_3215, n5023);
  and g8165 (n5024, n_272, n_3215);
  and g8166 (n5025, n669, n5023);
  not g8167 (n_3216, n5024);
  not g8168 (n_3217, n5025);
  and g8169 (n5026, n_3216, n_3217);
  not g8170 (n_3218, n5018);
  and g8171 (n5027, n_3218, n5026);
  not g8172 (n_3219, n5026);
  and g8173 (n5028, n_3211, n_3219);
  and g8174 (n5029, n_3210, n5028);
  not g8175 (n_3220, n5027);
  not g8176 (n_3221, n5029);
  and g8177 (n5030, n_3220, n_3221);
  not g8178 (n_3222, n4995);
  and g8179 (n5031, n_3222, n5030);
  not g8180 (n_3223, n5030);
  and g8181 (n5032, n4995, n_3223);
  not g8182 (n_3224, n5031);
  not g8183 (n_3225, n5032);
  and g8184 (n5033, n_3224, n_3225);
  not g8185 (n_3226, n4994);
  and g8186 (n5034, n_3226, n5033);
  not g8187 (n_3227, n5033);
  and g8188 (n5035, n4994, n_3227);
  not g8189 (n_3228, n5034);
  not g8190 (n_3229, n5035);
  and g8191 (n5036, n_3228, n_3229);
  not g8192 (n_3230, n5036);
  and g8193 (n5037, n4993, n_3230);
  not g8194 (n_3231, n4993);
  and g8195 (n5038, n_3231, n5036);
  not g8196 (n_3232, n5037);
  not g8197 (n_3233, n5038);
  and g8198 (n5039, n_3232, n_3233);
  not g8199 (n_3234, n4987);
  and g8200 (n5040, n_3234, n5039);
  not g8201 (n_3235, n5039);
  and g8202 (n5041, n4987, n_3235);
  not g8203 (n_3236, n5040);
  not g8204 (n_3237, n5041);
  and g8205 (n5042, n_3236, n_3237);
  not g8206 (n_3238, n5042);
  and g8207 (n5043, n_3188, n_3238);
  and g8208 (n5044, n4980, n5042);
  not g8209 (n_3239, n5043);
  not g8210 (n_3240, n5044);
  and g8211 (n5045, n_3239, n_3240);
  and g8212 (n5046, n_3190, n4982);
  not g8213 (n_3241, n5046);
  and g8214 (n5047, n_2468, n_3241);
  not g8215 (n_3242, n5045);
  and g8216 (n5048, n_3242, n5047);
  not g8217 (n_3243, n5047);
  and g8218 (n5049, n5045, n_3243);
  or g8219 (\sin[11] , n5048, n5049);
  and g8220 (n5051, n_3233, n_3236);
  and g8233 (n5064, n_3224, n_3228);
  and g8234 (n5065, n_3209, n_3220);
  and g8235 (n5066, n2695, n3896);
  and g8236 (n5067, n2690, n4054);
  not g8237 (n_3244, n5066);
  not g8238 (n_3245, n5067);
  and g8239 (n5068, n_3244, n_3245);
  not g8240 (n_3246, n5068);
  and g8241 (n5069, n_272, n_3246);
  and g8242 (n5070, n669, n5068);
  not g8243 (n_3247, n5069);
  not g8244 (n_3248, n5070);
  and g8245 (n5071, n_3247, n_3248);
  and g8246 (n5072, n2668, n3750);
  and g8247 (n5073, n2776, n3272);
  and g8248 (n5074, n2666, n_2220);
  and g8254 (n5077, n2674, n3762);
  not g8257 (n_3253, n5078);
  and g8258 (n5079, n_240, n_3253);
  not g8259 (n_3254, n5079);
  and g8260 (n5080, n_240, n_3254);
  and g8261 (n5081, n_3253, n_3254);
  not g8262 (n_3255, n5080);
  not g8263 (n_3256, n5081);
  and g8264 (n5082, n_3255, n_3256);
  not g8265 (n_3257, n5082);
  and g8266 (n5083, n5071, n_3257);
  not g8267 (n_3258, n5083);
  and g8268 (n5084, n5071, n_3258);
  and g8269 (n5085, n_3257, n_3258);
  not g8270 (n_3259, n5084);
  not g8271 (n_3260, n5085);
  and g8272 (n5086, n_3259, n_3260);
  and g8273 (n5087, n_3192, n_3193);
  not g8274 (n_3261, n5087);
  and g8275 (n5088, n_3206, n_3261);
  and g8276 (n5089, n_240, n_1931);
  and g8277 (n5090, n_3193, n5089);
  not g8278 (n_3262, n5089);
  and g8279 (n5091, n4997, n_3262);
  not g8280 (n_3263, n5088);
  not g8281 (n_3264, n5091);
  and g8282 (n5092, n_3263, n_3264);
  not g8283 (n_3265, n5090);
  and g8284 (n5093, n_3265, n5092);
  not g8285 (n_3266, n5093);
  and g8286 (n5094, n_3263, n_3266);
  and g8287 (n5095, n_3264, n_3266);
  and g8288 (n5096, n_3265, n5095);
  not g8289 (n_3267, n5094);
  not g8290 (n_3268, n5096);
  and g8291 (n5097, n_3267, n_3268);
  not g8292 (n_3269, n5086);
  and g8293 (n5098, n_3269, n5097);
  not g8294 (n_3270, n5097);
  and g8295 (n5099, n5086, n_3270);
  not g8296 (n_3271, n5098);
  not g8297 (n_3272, n5099);
  and g8298 (n5100, n_3271, n_3272);
  not g8299 (n_3273, n5065);
  not g8300 (n_3274, n5100);
  and g8301 (n5101, n_3273, n_3274);
  and g8302 (n5102, n5065, n5100);
  not g8303 (n_3275, n5101);
  not g8304 (n_3276, n5102);
  and g8305 (n5103, n_3275, n_3276);
  not g8306 (n_3277, n5064);
  and g8307 (n5104, n_3277, n5103);
  not g8308 (n_3278, n5103);
  and g8309 (n5105, n5064, n_3278);
  not g8310 (n_3279, n5104);
  not g8311 (n_3280, n5105);
  and g8312 (n5106, n_3279, n_3280);
  not g8313 (n_3281, n5106);
  and g8314 (n5107, n5063, n_3281);
  not g8315 (n_3282, n5063);
  and g8316 (n5108, n_3282, n5106);
  not g8317 (n_3283, n5107);
  not g8318 (n_3284, n5108);
  and g8319 (n5109, n_3283, n_3284);
  not g8320 (n_3285, n5051);
  and g8321 (n5110, n_3285, n5109);
  not g8322 (n_3286, n5109);
  and g8323 (n5111, n5051, n_3286);
  not g8324 (n_3287, n5110);
  not g8325 (n_3288, n5111);
  and g8326 (n5112, n_3287, n_3288);
  not g8327 (n_3289, n5112);
  and g8328 (n5113, n_3240, n_3289);
  and g8329 (n5114, n5044, n5112);
  not g8330 (n_3290, n5113);
  not g8331 (n_3291, n5114);
  and g8332 (n5115, n_3290, n_3291);
  and g8333 (n5116, n_3242, n5046);
  not g8334 (n_3292, n5116);
  and g8335 (n5117, n_2468, n_3292);
  not g8336 (n_3293, n5115);
  and g8337 (n5118, n_3293, n5117);
  not g8338 (n_3294, n5117);
  and g8339 (n5119, n5115, n_3294);
  or g8340 (\sin[12] , n5118, n5119);
  and g8341 (n5121, n_3284, n_3287);
  and g8359 (n5139, n_3275, n_3279);
  and g8360 (n5140, n2668, n3896);
  and g8361 (n5141, n2776, n_2220);
  and g8362 (n5142, n2666, n3750);
  and g8368 (n5145, n2674, n3908);
  not g8371 (n_3299, n5146);
  and g8372 (n5147, n_240, n_3299);
  not g8373 (n_3300, n5147);
  and g8374 (n5148, n_3299, n_3300);
  and g8375 (n5149, n_240, n_3300);
  not g8376 (n_3301, n5148);
  not g8377 (n_3302, n5149);
  and g8378 (n5150, n_3301, n_3302);
  and g8379 (n5151, n669, n5089);
  and g8380 (n5152, n_272, n_3262);
  not g8381 (n_3303, n5151);
  not g8382 (n_3304, n5152);
  and g8383 (n5153, n_3303, n_3304);
  and g8384 (n5154, n_240, n3272);
  and g8385 (n5155, n5153, n5154);
  not g8386 (n_3305, n5153);
  not g8387 (n_3306, n5154);
  and g8388 (n5156, n_3305, n_3306);
  not g8389 (n_3307, n5155);
  not g8390 (n_3308, n5156);
  and g8391 (n5157, n_3307, n_3308);
  not g8392 (n_3309, n5150);
  and g8393 (n5158, n_3309, n5157);
  not g8394 (n_3310, n5158);
  and g8395 (n5159, n_3309, n_3310);
  and g8396 (n5160, n5157, n_3310);
  not g8397 (n_3311, n5159);
  not g8398 (n_3312, n5160);
  and g8399 (n5161, n_3311, n_3312);
  not g8400 (n_3313, n5095);
  and g8401 (n5162, n_3313, n5161);
  not g8402 (n_3314, n5161);
  and g8403 (n5163, n5095, n_3314);
  not g8404 (n_3315, n5162);
  not g8405 (n_3316, n5163);
  and g8406 (n5164, n_3315, n_3316);
  and g8407 (n5165, n_3269, n_3270);
  not g8408 (n_3317, n5165);
  and g8409 (n5166, n_3258, n_3317);
  not g8410 (n_3318, n5164);
  not g8411 (n_3319, n5166);
  and g8412 (n5167, n_3318, n_3319);
  and g8413 (n5168, n5164, n5166);
  not g8414 (n_3320, n5167);
  not g8415 (n_3321, n5168);
  and g8416 (n5169, n_3320, n_3321);
  not g8417 (n_3322, n5139);
  and g8418 (n5170, n_3322, n5169);
  not g8419 (n_3323, n5169);
  and g8420 (n5171, n5139, n_3323);
  not g8421 (n_3324, n5170);
  not g8422 (n_3325, n5171);
  and g8423 (n5172, n_3324, n_3325);
  not g8424 (n_3326, n5138);
  and g8425 (n5173, n_3326, n5172);
  not g8426 (n_3327, n5172);
  and g8427 (n5174, n5138, n_3327);
  not g8428 (n_3328, n5121);
  not g8429 (n_3329, n5174);
  and g8430 (n5175, n_3328, n_3329);
  not g8431 (n_3330, n5173);
  and g8432 (n5176, n_3330, n5175);
  not g8433 (n_3331, n5176);
  and g8434 (n5177, n_3328, n_3331);
  and g8435 (n5178, n_3330, n_3331);
  and g8436 (n5179, n_3329, n5178);
  not g8437 (n_3332, n5177);
  not g8438 (n_3333, n5179);
  and g8439 (n5180, n_3332, n_3333);
  and g8440 (n5181, n_3291, n5180);
  not g8441 (n_3334, n5180);
  and g8442 (n5182, n5114, n_3334);
  not g8443 (n_3335, n5181);
  not g8444 (n_3336, n5182);
  and g8445 (n5183, n_3335, n_3336);
  and g8446 (n5184, n_3293, n5116);
  not g8447 (n_3337, n5184);
  and g8448 (n5185, n_2468, n_3337);
  not g8449 (n_3338, n5183);
  and g8450 (n5186, n_3338, n5185);
  not g8451 (n_3339, n5185);
  and g8452 (n5187, n5183, n_3339);
  or g8453 (\sin[13] , n5186, n5187);
  and g8468 (n5203, n_3320, n_3324);
  and g8469 (n5204, n_3313, n_3314);
  not g8470 (n_3340, n5204);
  and g8471 (n5205, n_3310, n_3340);
  and g8472 (n5206, n_240, n_2220);
  and g8473 (n5207, n_3303, n_3307);
  not g8474 (n_3341, n5206);
  not g8475 (n_3342, n5207);
  and g8476 (n5208, n_3341, n_3342);
  not g8477 (n_3343, n5208);
  and g8478 (n5209, n_3341, n_3343);
  and g8479 (n5210, n_3342, n_3343);
  not g8480 (n_3344, n5209);
  not g8481 (n_3345, n5210);
  and g8482 (n5211, n_3344, n_3345);
  and g8483 (n5212, n2776, n3750);
  and g8484 (n5213, n2666, n3896);
  not g8485 (n_3346, n5212);
  not g8486 (n_3347, n5213);
  and g8487 (n5214, n_3346, n_3347);
  and g8488 (n5215, n_1543, n5214);
  not g8489 (n_3348, n4056);
  and g8490 (n5216, n_3348, n5214);
  not g8491 (n_3349, n5215);
  not g8492 (n_3350, n5216);
  and g8493 (n5217, n_3349, n_3350);
  not g8494 (n_3351, n5217);
  and g8495 (n5218, n525, n_3351);
  and g8496 (n5219, n_240, n5217);
  not g8497 (n_3352, n5218);
  not g8498 (n_3353, n5219);
  and g8499 (n5220, n_3352, n_3353);
  not g8500 (n_3354, n5211);
  and g8501 (n5221, n_3354, n5220);
  not g8502 (n_3355, n5220);
  and g8503 (n5222, n5211, n_3355);
  not g8504 (n_3356, n5221);
  not g8505 (n_3357, n5222);
  and g8506 (n5223, n_3356, n_3357);
  not g8507 (n_3358, n5205);
  and g8508 (n5224, n_3358, n5223);
  not g8509 (n_3359, n5223);
  and g8510 (n5225, n5205, n_3359);
  not g8511 (n_3360, n5224);
  not g8512 (n_3361, n5225);
  and g8513 (n5226, n_3360, n_3361);
  not g8514 (n_3362, n5203);
  and g8515 (n5227, n_3362, n5226);
  not g8516 (n_3363, n5226);
  and g8517 (n5228, n5203, n_3363);
  not g8518 (n_3364, n5227);
  not g8519 (n_3365, n5228);
  and g8520 (n5229, n_3364, n_3365);
  not g8521 (n_3366, n5229);
  and g8522 (n5230, n5202, n_3366);
  not g8523 (n_3367, n5202);
  and g8524 (n5231, n_3367, n5229);
  not g8525 (n_3368, n5230);
  not g8526 (n_3369, n5231);
  and g8527 (n5232, n_3368, n_3369);
  not g8528 (n_3370, n5178);
  and g8529 (n5233, n_3370, n5232);
  not g8530 (n_3371, n5232);
  and g8531 (n5234, n5178, n_3371);
  not g8532 (n_3372, n5233);
  not g8533 (n_3373, n5234);
  and g8534 (n5235, n_3372, n_3373);
  not g8535 (n_3374, n5235);
  and g8536 (n5236, n_3336, n_3374);
  and g8537 (n5237, n5182, n5235);
  not g8538 (n_3375, n5236);
  not g8539 (n_3376, n5237);
  and g8540 (n5238, n_3375, n_3376);
  and g8541 (n5239, n_3338, n5184);
  not g8542 (n_3377, n5239);
  and g8543 (n5240, n_2468, n_3377);
  not g8544 (n_3378, n5238);
  and g8545 (n5241, n_3378, n5240);
  not g8546 (n_3379, n5240);
  and g8547 (n5242, n5238, n_3379);
  or g8548 (\sin[14] , n5241, n5242);
  and g8549 (n5244, n_3369, n_3372);
  and g8564 (n5259, n2776, n3896);
  and g8565 (n5260, n2674, n4054);
  not g8566 (n_3380, n5259);
  not g8567 (n_3381, n5260);
  and g8568 (n5261, n_3380, n_3381);
  not g8569 (n_3382, n5261);
  and g8570 (n5262, n_240, n_3382);
  not g8571 (n_3383, n5262);
  and g8572 (n5263, n_3382, n_3383);
  and g8573 (n5264, n_240, n_3383);
  not g8574 (n_3384, n5263);
  not g8575 (n_3385, n5264);
  and g8576 (n5265, n_3384, n_3385);
  and g8577 (n5266, n_240, n3759);
  not g8578 (n_3386, n5265);
  not g8579 (n_3387, n5266);
  and g8580 (n5267, n_3386, n_3387);
  not g8581 (n_3388, n5267);
  and g8582 (n5268, n_3386, n_3388);
  and g8583 (n5269, n_3387, n_3388);
  not g8584 (n_3389, n5268);
  not g8585 (n_3390, n5269);
  and g8586 (n5270, n_3389, n_3390);
  and g8587 (n5271, n_3343, n_3356);
  and g8588 (n5272, n5270, n5271);
  not g8589 (n_3391, n5270);
  not g8590 (n_3392, n5271);
  and g8591 (n5273, n_3391, n_3392);
  not g8592 (n_3393, n5272);
  not g8593 (n_3394, n5273);
  and g8594 (n5274, n_3393, n_3394);
  and g8595 (n5275, n_3360, n_3364);
  not g8596 (n_3395, n5274);
  and g8597 (n5276, n_3395, n5275);
  not g8598 (n_3396, n5275);
  and g8599 (n5277, n5274, n_3396);
  not g8600 (n_3397, n5276);
  not g8601 (n_3398, n5277);
  and g8602 (n5278, n_3397, n_3398);
  not g8603 (n_3399, n5258);
  and g8604 (n5279, n_3399, n5278);
  not g8605 (n_3400, n5278);
  and g8606 (n5280, n5258, n_3400);
  not g8607 (n_3401, n5244);
  not g8608 (n_3402, n5280);
  and g8609 (n5281, n_3401, n_3402);
  not g8610 (n_3403, n5279);
  and g8611 (n5282, n_3403, n5281);
  not g8612 (n_3404, n5282);
  and g8613 (n5283, n_3401, n_3404);
  and g8614 (n5284, n_3403, n_3404);
  and g8615 (n5285, n_3402, n5284);
  not g8616 (n_3405, n5283);
  not g8617 (n_3406, n5285);
  and g8618 (n5286, n_3405, n_3406);
  and g8619 (n5287, n_3376, n5286);
  not g8620 (n_3407, n5286);
  and g8621 (n5288, n5237, n_3407);
  not g8622 (n_3408, n5287);
  not g8623 (n_3409, n5288);
  and g8624 (n5289, n_3408, n_3409);
  and g8625 (n5290, n_3378, n5239);
  not g8626 (n_3410, n5290);
  and g8627 (n5291, n_2468, n_3410);
  not g8628 (n_3411, n5289);
  and g8629 (n5292, n_3411, n5291);
  not g8630 (n_3412, n5291);
  and g8631 (n5293, n5289, n_3412);
  or g8632 (\sin[15] , n5292, n5293);
  and g8642 (n5304, n_3394, n_3398);
  and g8643 (n5305, n3750, n_3341);
  and g8644 (n5306, n_240, n5305);
  not g8645 (n_3413, n5306);
  and g8646 (n5307, n_3388, n_3413);
  not g8647 (n_3414, n5304);
  and g8648 (n5308, n_3414, n5307);
  not g8649 (n_3415, n5307);
  and g8650 (n5309, n5304, n_3415);
  not g8651 (n_3416, n5308);
  not g8652 (n_3417, n5309);
  and g8653 (n5310, n_3416, n_3417);
  and g8654 (n5311, n3896, n_3341);
  and g8655 (n5312, n_2368, n5206);
  not g8656 (n_3418, n5311);
  not g8657 (n_3419, n5312);
  and g8658 (n5313, n_3418, n_3419);
  and g8659 (n5314, n_240, n5313);
  not g8660 (n_3420, n5314);
  and g8661 (n5315, n5310, n_3420);
  not g8662 (n_3421, n5310);
  and g8663 (n5316, n_3421, n5314);
  not g8664 (n_3422, n5315);
  not g8665 (n_3423, n5316);
  and g8666 (n5317, n_3422, n_3423);
  not g8667 (n_3424, n5303);
  not g8668 (n_3425, n5317);
  and g8669 (n5318, n_3424, n_3425);
  and g8670 (n5319, n5303, n5317);
  not g8671 (n_3426, n5284);
  not g8672 (n_3427, n5319);
  and g8673 (n5320, n_3426, n_3427);
  not g8674 (n_3428, n5318);
  and g8675 (n5321, n_3428, n5320);
  not g8676 (n_3429, n5321);
  and g8677 (n5322, n_3426, n_3429);
  and g8678 (n5323, n_3428, n_3429);
  and g8679 (n5324, n_3427, n5323);
  not g8680 (n_3430, n5322);
  not g8681 (n_3431, n5324);
  and g8682 (n5325, n_3430, n_3431);
  and g8683 (n5326, n_3409, n5325);
  not g8684 (n_3432, n5325);
  and g8685 (n5327, n5288, n_3432);
  not g8686 (n_3433, n5326);
  not g8687 (n_3434, n5327);
  and g8688 (n5328, n_3433, n_3434);
  and g8689 (n5329, n_3411, n5290);
  not g8690 (n_3435, n5329);
  and g8691 (n5330, n_2468, n_3435);
  not g8692 (n_3436, n5328);
  and g8693 (n5331, n_3436, n5330);
  not g8694 (n_3437, n5330);
  and g8695 (n5332, n5328, n_3437);
  or g8696 (\sin[16] , n5331, n5332);
  not g8708 (n_3438, n5323);
  not g8709 (n_3439, n5344);
  and g8710 (n5345, n_3438, n_3439);
  and g8711 (n5346, n5323, n5344);
  not g8712 (n_3440, n5345);
  not g8713 (n_3441, n5346);
  and g8714 (n5347, n_3440, n_3441);
  and g8715 (n5348, n_3434, n5347);
  not g8716 (n_3442, n5347);
  and g8717 (n5349, n5327, n_3442);
  not g8718 (n_3443, n5348);
  not g8719 (n_3444, n5349);
  and g8720 (n5350, n_3443, n_3444);
  and g8721 (n5351, n_3436, n5329);
  not g8722 (n_3445, n5351);
  and g8723 (n5352, n_2468, n_3445);
  not g8724 (n_3446, n5350);
  and g8725 (n5353, n_3446, n5352);
  not g8726 (n_3447, n5352);
  and g8727 (n5354, n5350, n_3447);
  not g8728 (n_3448, n5353);
  not g8729 (n_3449, n5354);
  and g8730 (\sin[17] , n_3448, n_3449);
  and g8731 (n5356, n5327, n5347);
  not g8743 (n_3450, n5367);
  and g8744 (n5368, n5345, n_3450);
  and g8745 (n5369, n_3440, n5367);
  not g8746 (n_3451, n5368);
  not g8747 (n_3452, n5369);
  and g8748 (n5370, n_3451, n_3452);
  not g8749 (n_3453, n5356);
  not g8750 (n_3454, n5370);
  and g8751 (n5371, n_3453, n_3454);
  and g8752 (n5372, n5356, n_3452);
  not g8753 (n_3455, n5371);
  not g8754 (n_3456, n5372);
  and g8755 (n5373, n_3455, n_3456);
  and g8756 (n5374, n5350, n5351);
  not g8757 (n_3457, n5374);
  and g8758 (n5375, n_2468, n_3457);
  not g8759 (n_3458, n5373);
  and g8760 (n5376, n_3458, n5375);
  not g8761 (n_3459, n5375);
  and g8762 (n5377, n5373, n_3459);
  or g8763 (\sin[18] , n5376, n5377);
  and g8775 (n5390, n_3451, n5389);
  not g8776 (n_3460, n5389);
  and g8777 (n5391, n5368, n_3460);
  not g8778 (n_3461, n5390);
  not g8779 (n_3462, n5391);
  and g8780 (n5392, n_3461, n_3462);
  not g8781 (n_3463, n5392);
  and g8782 (n5393, n_3456, n_3463);
  and g8783 (n5394, n5372, n5392);
  not g8784 (n_3464, n5393);
  not g8785 (n_3465, n5394);
  and g8786 (n5395, n_3464, n_3465);
  and g8787 (n5396, n_3458, n5374);
  not g8788 (n_3466, n5396);
  and g8789 (n5397, n_2468, n_3466);
  not g8790 (n_3467, n5395);
  and g8791 (n5398, n_3467, n5397);
  not g8792 (n_3468, n5397);
  and g8793 (n5399, n5395, n_3468);
  or g8794 (\sin[19] , n5398, n5399);
  not g8807 (n_3469, n5412);
  and g8808 (n5413, n5391, n_3469);
  and g8809 (n5414, n_3462, n5412);
  not g8810 (n_3470, n5413);
  not g8811 (n_3471, n5414);
  and g8812 (n5415, n_3470, n_3471);
  not g8813 (n_3472, n5415);
  and g8814 (n5416, n_3465, n_3472);
  and g8815 (n5417, n5394, n_3471);
  not g8816 (n_3473, n5416);
  not g8817 (n_3474, n5417);
  and g8818 (n5418, n_3473, n_3474);
  and g8819 (n5419, n_3467, n5396);
  not g8820 (n_3475, n5419);
  and g8821 (n5420, n_2468, n_3475);
  not g8822 (n_3476, n5418);
  and g8823 (n5421, n_3476, n5420);
  not g8824 (n_3477, n5420);
  and g8825 (n5422, n5418, n_3477);
  or g8826 (\sin[20] , n5421, n5422);
  and g8831 (n5428, n_3470, n5427);
  not g8832 (n_3478, n5427);
  and g8833 (n5429, n5413, n_3478);
  not g8834 (n_3479, n5428);
  not g8835 (n_3480, n5429);
  and g8836 (n5430, n_3479, n_3480);
  not g8837 (n_3481, n5430);
  and g8838 (n5431, n_3474, n_3481);
  and g8839 (n5432, n5417, n5430);
  not g8840 (n_3482, n5431);
  not g8841 (n_3483, n5432);
  and g8842 (n5433, n_3482, n_3483);
  and g8843 (n5434, n_3476, n5419);
  not g8844 (n_3484, n5434);
  and g8845 (n5435, n_2468, n_3484);
  not g8846 (n_3485, n5433);
  and g8847 (n5436, n_3485, n5435);
  not g8848 (n_3486, n5435);
  and g8849 (n5437, n5433, n_3486);
  or g8850 (\sin[21] , n5436, n5437);
  and g8851 (n5439, n444, n517);
  not g8852 (n_3487, n5439);
  and g8853 (n5440, n5429, n_3487);
  and g8854 (n5441, n_3480, n5439);
  not g8855 (n_3488, n5440);
  not g8856 (n_3489, n5441);
  and g8857 (n5442, n_3488, n_3489);
  not g8858 (n_3490, n5442);
  and g8859 (n5443, n_3483, n_3490);
  and g8860 (n5444, n5432, n_3489);
  not g8861 (n_3491, n5443);
  not g8862 (n_3492, n5444);
  and g8863 (n5445, n_3491, n_3492);
  and g8864 (n5446, n_3485, n5434);
  not g8865 (n_3493, n5446);
  and g8866 (n5447, n_2468, n_3493);
  not g8867 (n_3494, n5445);
  and g8868 (n5448, n_3494, n5447);
  not g8869 (n_3495, n5447);
  and g8870 (n5449, n5445, n_3495);
  or g8871 (\sin[22] , n5448, n5449);
  and g8872 (n5451, n_49, n71);
  and g8873 (n5452, n_3488, n_3492);
  and g8874 (n5453, n5440, n5444);
  not g8875 (n_3496, n5452);
  not g8876 (n_3497, n5453);
  and g8877 (n5454, n_3496, n_3497);
  and g8878 (n5455, n_3494, n5446);
  not g8879 (n_3498, n5455);
  and g8880 (n5456, n_2468, n_3498);
  not g8881 (n_3499, n5456);
  and g8882 (n5457, n5454, n_3499);
  not g8883 (n_3500, n5454);
  and g8884 (n5458, n_3500, n5456);
  not g8885 (n_3501, n5457);
  not g8886 (n_3502, n5458);
  and g8887 (n5459, n_3501, n_3502);
  not g8888 (n_3503, n5459);
  or g8889 (\sin[23] , n5451, n_3503);
  and g8890 (n5461, n_3496, n5455);
  and g8891 (n5462, n_3497, n_3498);
  not g8892 (n_3504, n5461);
  not g8893 (n_3505, n5462);
  and g8894 (n5463, n_3504, n_3505);
  not g8895 (n_3506, n5451);
  and g8896 (n5464, n_3506, n5463);
  not g8897 (n_3507, n5464);
  and g8898 (\sin[24] , n_2468, n_3507);
  and g8899 (n_3532, n_196, n_88, n_141);
  and g8900 (n_3533, n210, n623, n643);
  and g8901 (n_3534, n2311, n1459, n806);
  and g8902 (n_3535, n239, n1093);
  and g8903 (n3861, n_3532, n_3533, n_3534, n_3535);
  and g8904 (n_3536, n_190, n_204, n_133);
  and g8905 (n_3537, n_144, n_107, n_210);
  and g8906 (n_3538, n614, n505);
  and g8907 (n_3539, n153, n432);
  and g8908 (n623, n_3536, n_3537, n_3538, n_3539);
  and g8909 (n_3540, n_177, n_176);
  and g8910 (n_3541, n_101, n_109);
  and g8911 (n643, n637, n638, n_3540, n_3541);
  and g8912 (n_3542, n_197, n_215, n_217);
  and g8913 (n_3543, n_191, n369);
  and g8914 (n_3544, n644, n944);
  and g8915 (n_3545, n141, n1116);
  and g8916 (n2311, n_3542, n_3543, n_3544, n_3545);
  and g8917 (n_3546, n_150, n_149, n_148, n_147);
  and g8918 (n_3547, n_146, n_145, n_144);
  and g8919 (n_3548, n165, n204, n210);
  and g8920 (n_3549, n253, n256, n259);
  and g8921 (n271, n_3546, n_3547, n_3548, n_3549);
  and g8922 (n_3550, n_91, n_188);
  and g8923 (n_3551, n_198, n_118);
  and g8924 (n614, n474, n609, n_3550, n_3551);
  and g8925 (n_3552, n_194, n_321);
  and g8926 (n_3553, n_96, n_110);
  and g8927 (n_3554, n_132, n_98);
  and g8928 (n944, n_136, n_3552, n_3553, n_3554);
  and g8929 (n_3555, n_194, n_222, n_193, n_180);
  and g8930 (n_3556, n_87, n_218, n_189);
  and g8931 (n_3557, n_140, n_94, n980);
  and g8932 (n_3558, n3666, n2454, n3678);
  and g8933 (n3690, n_3555, n_3556, n_3557, n_3558);
  and g8934 (n_3559, n_97, n_96);
  and g8935 (n_3560, n_95, n_94);
  and g8936 (n_3561, n_93, n141);
  and g8937 (n_3562, n145, n158);
  and g8938 (n165, n_3559, n_3560, n_3561, n_3562);
  and g8939 (n_3563, n_114, n_113);
  and g8940 (n204, n185, n189, n200, n_3563);
  and g8941 (n_3564, n_139, n_138);
  and g8942 (n253, n_137, n_136, n249, n_3564);
  and g8943 (n_3565, n_150, n_85, n_202);
  and g8944 (n_3566, n_96, n_182, n_106);
  and g8945 (n_3567, n_89, n_83);
  and g8946 (n_3568, n806, n3657);
  and g8947 (n3666, n_3565, n_3566, n_3567, n_3568);
  and g8948 (n_3569, n_260, n_197);
  and g8949 (n2454, n_118, n_90, n1117, n_3569);
  and g8950 (n3678, n_179, n_213, n789, n3675);
  and g8951 (n_3570, n_177, n_132, n_102, n_131);
  and g8952 (n_3571, n_184, n_89, n_212, n2364);
  and g8953 (n_3572, n3699, n3702, n344);
  and g8954 (n_3573, n2433, n460, n2422);
  and g8955 (n3715, n_3570, n_3571, n_3572, n_3573);
  and g8956 (n_3574, n_105, n_104);
  and g8957 (n_3575, n_103, n_102);
  and g8958 (n_3576, n_101, n_100);
  and g8959 (n185, n179, n_3574, n_3575, n_3576);
  and g8960 (n_3577, n_112, n_111);
  and g8961 (n200, n_110, n_108, n_109, n_3577);
  and g8962 (n_3578, n_135, n_134, n_133);
  and g8963 (n_3579, n_132, n_131, n_130);
  and g8964 (n_3580, n_129, n_128, n233);
  and g8965 (n_3581, n236, n239);
  and g8966 (n249, n_3578, n_3579, n_3580, n_3581);
  and g8967 (n_3582, n_91, n_181);
  and g8968 (n3657, n_321, n_148, n_228, n_3582);
  and g8969 (n_3583, n_135, n_221, n_225);
  and g8970 (n_3584, n_261, n_226, n_141);
  and g8971 (n_3585, n_133, n1134);
  and g8972 (n_3586, n372, n505);
  and g8973 (n3675, n_3583, n_3584, n_3585, n_3586);
  and g8974 (n_3587, n_125, n_261);
  and g8975 (n_3588, n_122, n_182);
  and g8976 (n_3589, n_213, n141);
  and g8977 (n2364, n_185, n_3587, n_3588, n_3589);
  and g8978 (n_3590, n_219, n_205);
  and g8979 (n_3591, n_229, n_86);
  and g8980 (n_3592, n2303, n397);
  and g8981 (n3699, n2278, n_3590, n_3591, n_3592);
  and g8982 (n3702, n_92, n_94, n341, n813);
  and g8983 (n_3593, n_123, n_122);
  and g8984 (n_3594, n_121, n_120);
  and g8985 (n233, n_118, n_119, n_3593, n_3594);
  and g8986 (n_3595, n_214, n_130);
  and g8987 (n1134, n807, n459, n1116, n_3595);
  and g8988 (n_3596, n_105, n_134);
  and g8989 (n_3597, n_204, n_124);
  and g8990 (n_3598, n_103, n_146);
  and g8991 (n_3599, n_93, n_118);
  and g8992 (n2303, n_3596, n_3597, n_3598, n_3599);
  and g8993 (n_3600, n_193, n_192);
  and g8994 (n341, n_101, n_107, n_191, n_3600);
  and g8995 (n_3601, n_206, n_143);
  and g8996 (n813, n149, n301, n809, n_3601);
  nor g8997 (n3764, n3751, n3752, n3753, n3763);
  nor g8998 (n3334, n3326, n3327, n3328, n3333);
  nor g8999 (n3522, n3516, n3517, n3518, n3521);
  nor g9000 (n3551, n3545, n3546, n3547, n3550);
  nor g9001 (n3506, n3500, n3501, n3502, n3505);
  nor g9002 (n3494, n3344, n3347, n3349, n3491);
  nor g9003 (n2654, n2555, n2563, n2568, n2653);
  and g9004 (n_3602, n_123, n_97, n_139, n_260);
  and g9005 (n_3603, n_132, n_98, n_184, n_128);
  and g9006 (n_3604, n2418, n3734, n1162);
  and g9007 (n_3605, n334, n353, n_224);
  and g9008 (n3747, n_3602, n_3603, n_3604, n_3605);
  and g9009 (n_3606, n_84, n3259, n453);
  and g9010 (n_3607, n502, n485, n314);
  and g9011 (n_3608, n437, n397, n1165);
  and g9012 (n_3609, n349, n423);
  and g9013 (n3269, n_3606, n_3607, n_3608, n_3609);
  nor g9014 (n3024, n3016, n3017, n3018, n3023);
  and g9015 (n_3610, n_223, n_225);
  and g9016 (n_3611, n_115, n_182);
  and g9017 (n_3612, n_146, n_209);
  and g9018 (n_3613, n239, n590);
  and g9019 (n3734, n_3610, n_3611, n_3612, n_3613);
  and g9020 (n_3614, n_135, n_91, n_196);
  and g9021 (n_3615, n_143, n_192, n_113);
  and g9022 (n_3616, n475, n1152, n_186);
  and g9023 (n_3617, n560, n969);
  and g9024 (n1162, n_3614, n_3615, n_3616, n_3617);
  and g9025 (n334, n_190, n_105, n_189, n331);
  and g9026 (n_3618, n_122, n_131);
  and g9027 (n_3619, n_107, n404);
  and g9028 (n_3620, n414, n485);
  and g9029 (n_3621, n514, n3617);
  and g9030 (n3624, n_3618, n_3619, n_3620, n_3621);
  and g9031 (n502, n_202, n_117, n_124, n499);
  and g9032 (n_3622, n_221, n_220);
  and g9033 (n_3623, n_208, n_150);
  and g9034 (n_3624, n473, n474);
  and g9035 (n_3625, n476, n478);
  and g9036 (n485, n_3622, n_3623, n_3624, n_3625);
  and g9037 (n_3626, n_96, n_120);
  and g9038 (n_3627, n_185, n_101);
  and g9039 (n437, n_99, n_118, n_3626, n_3627);
  and g9040 (n1165, n_149, n_85, n_116, n_210);
  and g9041 (n_3628, n_126, n_143, n_138, n_180);
  and g9042 (n_3629, n_227, n976, n2418);
  and g9043 (n_3630, n2333, n2244, n431);
  and g9044 (n_3631, n485, n_186, n809);
  and g9045 (n3229, n_3628, n_3629, n_3630, n_3631);
  and g9046 (n_3632, n_219, n_201, n_218, n_106);
  and g9047 (n_3633, n_118, n_130, n_100, n_89);
  and g9048 (n_3634, n210, n3243, n768);
  and g9049 (n_3635, n156, n744, n2366);
  and g9050 (n3256, n_3632, n_3633, n_3634, n_3635);
  nor g9051 (n3486, n3355, n3358, n3359, n3483);
  and g9052 (n_3636, n_321, n_263);
  and g9053 (n_3637, n_178, n_198);
  and g9054 (n_3638, n_136, n_108);
  and g9055 (n_3639, n637, n911);
  and g9056 (n1152, n_3636, n_3637, n_3638, n_3639);
  and g9057 (n_3640, n_113, n395);
  and g9058 (n_3641, n_119, n_116);
  and g9059 (n_3642, n141, n314);
  and g9060 (n_3643, n396, n397);
  and g9061 (n404, n_3640, n_3641, n_3642, n_3643);
  and g9062 (n414, n_146, n_211, n407, n411);
  and g9063 (n_3644, n_229, n_148);
  and g9064 (n_3645, n_104, n_179);
  and g9065 (n_3646, n_177, n505);
  and g9066 (n514, n508, n_3644, n_3645, n_3646);
  and g9067 (n499, n_183, n_203, n_226, n496);
  and g9068 (n_3647, n_121, n_131);
  and g9069 (n421, n_145, n153, n189, n_3647);
  and g9070 (n2333, n_196, n_321, n_137, n508);
  and g9071 (n_3648, n_127, n_149);
  and g9072 (n_3649, n_88, n_215);
  and g9073 (n2244, n_140, n906, n_3648, n_3649);
  and g9074 (n_3650, n_95, n_136, n_100);
  and g9075 (n_3651, n_144, n_86);
  and g9076 (n_3652, n_128, n414);
  and g9077 (n_3653, n416, n423);
  and g9078 (n431, n_3650, n_3651, n_3652, n_3653);
  and g9079 (n_3654, n_194, n_150, n_203, n_148);
  and g9080 (n_3655, n_193, n_215, n_207);
  and g9081 (n_3656, n_137, n_120, n_212);
  and g9082 (n_3657, n2166, n200, n3231);
  and g9083 (n3243, n_3654, n_3655, n_3656, n_3657);
  and g9084 (n_3658, n_225, n_263, n_85);
  and g9085 (n_3659, n_142, n_107);
  and g9086 (n_3660, n753, n757);
  and g9087 (n_3661, n759, n760);
  and g9088 (n768, n_3658, n_3659, n_3660, n_3661);
  and g9089 (n_3662, n_125, n_199);
  and g9090 (n_3663, n_228, n_229);
  and g9091 (n744, n_191, n_226, n_3662, n_3663);
  and g9092 (n_3664, n_123, n_260, n_263);
  and g9093 (n_3665, n945, n_178, n149);
  and g9094 (n_3666, n653, n2540, n1468);
  and g9095 (n_3667, n2339, n478, n1091);
  and g9096 (n2551, n_3664, n_3665, n_3666, n_3667);
  and g9097 (n411, n_178, n_130, n_93, n_210);
  and g9098 (n_3668, n_88, n_132);
  and g9099 (n757, n_209, n_198, n645, n_3668);
  and g9100 (n_3669, n_97, n_221);
  and g9101 (n_3670, n_129, n_86);
  and g9102 (n653, n256, n648, n_3669, n_3670);
  and g9103 (n_3671, n_206, n_102);
  and g9104 (n_3672, n_118, n_107);
  and g9105 (n2540, n_210, n796, n_3671, n_3672);
  and g9106 (n_3673, n_208, n_124, n_213);
  and g9107 (n_3674, n_136, n_191, n644);
  and g9108 (n_3675, n968, n1459);
  and g9109 (n_3676, n432, n584);
  and g9110 (n1468, n_3673, n_3674, n_3675, n_3676);
  and g9111 (n_3677, n_223, n_190);
  and g9112 (n_3678, n_148, n_104);
  and g9113 (n_3679, n931, n303);
  and g9114 (n2339, n759, n_3677, n_3678, n_3679);
  and g9115 (n_3680, n_135, n_208, n_227, n_98);
  and g9116 (n_3681, n_119, n_187, n2166, n2178);
  and g9117 (n_3682, n2190, n2196, n773);
  and g9118 (n_3683, n397, n153, n808);
  and g9119 (n2209, n_3680, n_3681, n_3682, n_3683);
  nor g9120 (n3477, n3365, n3368, n3369, n3474);
  and g9121 (n584, n_216, n_188, n_132, n_195);
  and g9122 (n_3684, n_95, n_116, n311);
  and g9123 (n_3685, n323, n325, n334);
  and g9124 (n_3686, n341, n344, n259);
  and g9125 (n_3687, n346, n349, n382);
  and g9126 (n393, n_3684, n_3685, n_3686, n_3687);
  and g9127 (n_3688, n_126, n_105, n_203, n_180);
  and g9128 (n_3689, n_217, n1104, n606, n967);
  and g9129 (n_3690, n739, n637, n474);
  and g9130 (n_3691, n319, n145, n794);
  and g9131 (n2225, n_3688, n_3689, n_3690, n_3691);
  and g9132 (n_3692, n_321, n_262, n_112);
  and g9133 (n_3693, n_117, n_113);
  and g9134 (n_3694, n_132, n_120);
  and g9135 (n_3695, n760, n2170);
  and g9136 (n2178, n_3692, n_3693, n_3694, n_3695);
  and g9137 (n_3696, n_91, n753);
  and g9138 (n_3697, n986, n2181);
  and g9139 (n_3698, n1091, n476);
  and g9140 (n_3699, n555, n2183);
  and g9141 (n2190, n_3696, n_3697, n_3698, n_3699);
  and g9142 (n_3700, n_261, n_88);
  and g9143 (n_3701, n_204, n_217);
  and g9144 (n_3702, n_178, n_84);
  and g9145 (n2196, n792, n_3700, n_3701, n_3702);
  and g9146 (n_3703, n_221, n_105);
  and g9147 (n_3704, n_183, n_215);
  and g9148 (n773, n_94, n_182, n_3703, n_3704);
  nor g9149 (n2832, n2824, n2825, n2826, n2831);
  and g9150 (n_3705, n_181, n_180, n_179);
  and g9151 (n_3706, n_111, n_178);
  and g9152 (n_3707, n_94, n301);
  and g9153 (n_3708, n179, n303);
  and g9154 (n311, n_3705, n_3706, n_3707, n_3708);
  and g9155 (n_3709, n_138, n_185);
  and g9156 (n323, n314, n316, n319, n_3709);
  and g9157 (n_3710, n_223, n_138, n_189);
  and g9158 (n_3711, n_109, n149);
  and g9159 (n_3712, n983, n1091);
  and g9160 (n_3713, n1093, n1096);
  and g9161 (n1104, n_3710, n_3711, n_3712, n_3713);
  and g9162 (n_3714, n_260, n_228);
  and g9163 (n_3715, n_179, n_103);
  and g9164 (n_3716, n_95, n_130);
  and g9165 (n_3717, n141, n373);
  and g9166 (n606, n_3714, n_3715, n_3716, n_3717);
  and g9167 (n_3718, n_204, n_202);
  and g9168 (n_3719, n_124, n_132);
  and g9169 (n_3720, n_209, n_92);
  and g9170 (n967, n961, n_3718, n_3719, n_3720);
  and g9171 (n739, n_321, n_134, n_146, n_113);
  and g9172 (n_3721, n_194, n_190);
  and g9173 (n2170, n_203, n_140, n_188, n_3721);
  and g9174 (n986, n_216, n_109, n_144, n_99);
  and g9175 (n2181, n_205, n_180, n_212, n626);
  and g9176 (n792, n_123, n_197, n_104, n_106);
  nor g9177 (n3085, n3079, n3080, n3081, n3084);
  nor g9178 (n3776, n3770, n3771, n3772, n3775);
  and g9179 (n_3722, n_123, n_87);
  and g9180 (n_3723, n_96, n_102);
  and g9181 (n_3724, n355, n366);
  and g9182 (n_3725, n372, n373);
  and g9183 (n380, n_3722, n_3723, n_3724, n_3725);
  and g9184 (n983, n_213, n_119, n_214, n980);
  and g9185 (n1096, n_220, n_229, n_101, n_195);
  nor g9186 (n3563, n3557, n3558, n3559, n3562);
  nor g9187 (n2752, n2743, n2744, n2745, n2751);
  and g9188 (n_3726, n_260, n_192, n_184);
  and g9189 (n_3727, n2239, n2250, n644);
  and g9190 (n_3728, n577, n156, n2252);
  and g9191 (n_3729, n478, n2254);
  and g9192 (n2264, n_3726, n_3727, n_3728, n_3729);
  and g9193 (n_3730, n_205, n_204);
  and g9194 (n366, n_203, n_202, n362, n_3730);
  nor g9195 (n3453, n3376, n3379, n3380, n3450);
  nor g9196 (n2956, n2950, n2951, n2952, n2955);
  and g9197 (n_3731, n_182, n_200, n_113);
  and g9198 (n_3732, n_195, n_100, n980);
  and g9199 (n_3733, n2276, n2196, n325);
  and g9200 (n_3734, n2278, n1459, n2281);
  and g9201 (n2292, n_3731, n_3732, n_3733, n_3734);
  and g9202 (n_3735, n_117, n_121, n_214);
  and g9203 (n_3736, n_129, n355, n2166);
  and g9204 (n_3737, n637, n301, n236);
  and g9205 (n_3738, n331, n2183);
  and g9206 (n2239, n_3735, n_3736, n_3737, n_3738);
  and g9207 (n_3739, n_321, n_146);
  and g9208 (n_3740, n_213, n_118);
  and g9209 (n_3741, n2244, n581);
  and g9210 (n2250, n628, n_3739, n_3740, n_3741);
  and g9211 (n_3742, n_222, n_138);
  and g9212 (n577, n_200, n_191, n573, n_3742);
  and g9213 (n_3743, n_214, n_184);
  and g9214 (n_3744, n_109, n_187);
  and g9215 (n_3745, n404, n431);
  and g9216 (n_3746, n432, n437);
  and g9217 (n444, n_3743, n_3744, n_3745, n_3746);
  nor g9218 (n2770, n2762, n2763, n2764, n2769);
  nor g9219 (n2863, n2857, n2858, n2859, n2862);
  and g9220 (n_3747, n_264, n_208, n_193);
  and g9221 (n_3748, n_202, n_144, n_107);
  and g9222 (n_3749, n_83, n451);
  and g9223 (n_3750, n396, n2252);
  and g9224 (n2276, n_3747, n_3748, n_3749, n_3750);
  and g9225 (n2281, n_135, n_181, n_90, n2239);
  and g9226 (n581, n_223, n_229, n_148, n578);
  nor g9227 (n3462, n3456, n3457, n3458, n3461);
  and g9228 (n_3751, n_264, n_112, n_203);
  and g9229 (n_3752, n_110, n_213, n2190);
  and g9230 (n_3753, n739, n2395, n373);
  and g9231 (n_3754, n914, n777, n1096);
  and g9232 (n2495, n_3751, n_3752, n_3753, n_3754);
  and g9233 (n_3755, n_123, n_225);
  and g9234 (n_3756, n_206, n467);
  and g9235 (n494, n_224, n489, n_3755, n_3756);
  nor g9236 (n692, n685, n686, n688, n689);
  nor g9237 (n3113, n3107, n3108, n3109, n3112);
  and g9238 (n_3757, n_123, n_190);
  and g9239 (n_3758, n_148, n_200);
  and g9240 (n_3759, n411, n906);
  and g9241 (n_3760, n564, n2254);
  and g9242 (n2395, n_3757, n_3758, n_3759, n_3760);
  and g9243 (n914, n_196, n_209, n_128, n911);
  and g9244 (n_3761, n_149, n_218);
  and g9245 (n_3762, n_137, n453);
  and g9246 (n_3763, n457, n459);
  and g9247 (n_3764, n349, n460);
  and g9248 (n467, n_3761, n_3762, n_3763, n_3764);
  and g9249 (n_3765, n_223, n_181);
  and g9250 (n489, n_105, n_222, n485, n_3765);
  and g9251 (n517, n473, n475, n467, n514);
  nor g9252 (n3428, n3387, n3390, n3391, n3425);
  nor g9253 (n3574, n3568, n3569, n3570, n3573);
  nor g9254 (n3790, n3784, n3785, n3786, n3789);
  and g9255 (n_3766, n_225, n450, n_179);
  and g9256 (n_3767, n_131, n_108, n_210);
  and g9257 (n_3768, n_187, n2303, n2311);
  and g9258 (n_3769, n2313, n2317);
  and g9259 (n2327, n_3766, n_3767, n_3768, n_3769);
  and g9260 (n_3770, n_226, n_133, n_90, n2333);
  and g9261 (n_3771, n930, n995, n2339);
  and g9262 (n_3772, n314, n344, n1106);
  and g9263 (n_3773, n2340, n432, n2342);
  and g9264 (n2354, n_3770, n_3771, n_3772, n_3773);
  and g9265 (n_3774, n_220, n_197, n_113);
  and g9266 (n_3775, n_214, n_129, n_109);
  and g9267 (n_3776, n2364, n753, n2375);
  and g9268 (n_3777, n382, n448);
  and g9269 (n2385, n_3774, n_3775, n_3776, n_3777);
  and g9270 (n_3778, n_85, n_138);
  and g9271 (n457, n_122, n_140, n_195, n_3778);
  nor g9272 (n3167, n3161, n3162, n3163, n3166);
  nor g9273 (n2919, n2913, n2914, n2915, n2918);
  nor g9274 (n2966, n2960, n2961, n2962, n2965);
  and g9275 (n_3779, n_223, n_139);
  and g9276 (n2317, n_87, n_133, n_119, n_3779);
  and g9277 (n_3780, n_208, n_262);
  and g9278 (n930, n_134, n_145, n407, n_3780);
  and g9279 (n_3781, n_123, n787, n_103);
  and g9280 (n_3782, n_130, n_100, n_187);
  and g9281 (n_3783, n926, n983);
  and g9282 (n_3784, n256, n986);
  and g9283 (n995, n_3781, n_3782, n_3783, n_3784);
  and g9284 (n_3785, n_181, n_194, n_260, n_143);
  and g9285 (n_3786, n_124, n_192, n_120, n_131);
  and g9286 (n_3787, n_119, n149, n986, n752);
  and g9287 (n_3788, n2395, n590, n2400);
  and g9288 (n2414, n_3785, n_3786, n_3787, n_3788);
  and g9289 (n_3789, n_229, n_111, n_188);
  and g9290 (n_3790, n_198, n_189);
  and g9291 (n_3791, n_107, n910);
  and g9292 (n_3792, n2366, n2367);
  and g9293 (n2375, n_3789, n_3790, n_3791, n_3792);
  nor g9294 (n711, n705, n706, n707, n708);
  nor g9295 (n3437, n3431, n3432, n3433, n3436);
  and g9296 (n_3793, n_91, n_226, n_227);
  and g9297 (n_3794, n_106, n_109, n_90);
  and g9298 (n_3795, n910, n323);
  and g9299 (n_3796, n303, n914);
  and g9300 (n923, n_3793, n_3794, n_3795, n_3796);
  and g9301 (n926, n_225, n_197, n_207, n_224);
  and g9302 (n_3797, n_127, n_200, n_142, n_136);
  and g9303 (n_3798, n_187, n165, n2432, n983);
  and g9304 (n_3799, n323, n325, n2400);
  and g9305 (n_3800, n2433, n396, n806);
  and g9306 (n2446, n_3797, n_3798, n_3799, n_3800);
  and g9307 (n_3801, n_127, n_150, n_117);
  and g9308 (n_3802, n_180, n_227);
  and g9309 (n_3803, n_83, n739);
  and g9310 (n_3804, n476, n744);
  and g9311 (n752, n_3801, n_3802, n_3803, n_3804);
  and g9312 (n_3805, n_208, n_122);
  and g9313 (n_3806, n_147, n_179);
  and g9314 (n2400, n416, n473, n_3805, n_3806);
  and g9315 (n_3807, n_225, n_204, n_122, n_146);
  and g9316 (n_3808, n_110, n_95, n_116, n_191);
  and g9317 (n_3809, n789, n2464, n2339);
  and g9318 (n_3810, n474, n256, n2422);
  and g9319 (n2477, n_3807, n_3808, n_3809, n_3810);
  and g9320 (n_3811, n_181, n_127);
  and g9321 (n910, n_263, n145, n906, n_3811);
  nor g9322 (n_3812, n3392, n3393);
  nor g9323 (n_3813, n3399, n3400);
  nor g9324 (n_3814, n3401, n3402);
  and g9325 (n3408, n_171, n_3812, n_3813, n_3814);
  and g9326 (n_3815, n_123, n_220, n_203);
  and g9327 (n_3816, n_202, n926, n2333);
  and g9328 (n_3817, n373, n2278, n2421);
  and g9329 (n_3818, n970, n2422);
  and g9330 (n2432, n_3815, n_3816, n_3817, n_3818);
  and g9331 (n_3819, n_91, n_263);
  and g9332 (n_3820, n_202, n_217);
  and g9333 (n_3821, n_195, n2454);
  and g9334 (n2464, n2458, n_3819, n_3820, n_3821);
  nor g9335 (n905, n899, n900, n901, n902);
  nor g9336 (n852, n845, n846, n848, n849);
  nor g9337 (n859, n853, n854, n855, n856);
  nor g9338 (n3416, n3410, n3411, n3412, n3415);
  and g9339 (n2421, n_219, n_149, n_193, n2418);
  and g9340 (n_3822, n_97, n_201);
  and g9341 (n2458, n_207, n_100, n_185, n_3822);
  nor g9342 (n879, n873, n874, n875, n876);
  and g9343 (n_3823, n_263, n355, n571);
  and g9344 (n_3824, n577, n581);
  and g9345 (n_3825, n584, n586);
  and g9346 (n_3826, n588, n590);
  and g9347 (n598, n_3823, n_3824, n_3825, n_3826);
  and g9348 (n_3827, n_208, n_263, n362);
  and g9349 (n_3828, n636, n643);
  and g9350 (n_3829, n644, n646);
  and g9351 (n_3830, n179, n655);
  and g9352 (n663, n_3827, n_3828, n_3829, n_3830);
  nor g9353 (n1041, n1034, n1035, n1037, n1038);
  nor g9354 (n1048, n1042, n1043, n1044, n1045);
  and g9355 (n_3831, n_261, n_198);
  and g9356 (n_3832, n_144, n185);
  and g9357 (n_3833, n558, n560);
  and g9358 (n_3834, n562, n564);
  and g9359 (n571, n_3831, n_3832, n_3833, n_3834);
  and g9360 (n_3835, n_139, n_264, n_218);
  and g9361 (n_3836, n_111, n606);
  and g9362 (n_3837, n608, n344);
  and g9363 (n_3838, n625, n628);
  and g9364 (n636, n_3835, n_3836, n_3837, n_3838);
  nor g9365 (n1032, n1026, n1027, n1028, n1029);
  and g9366 (n_3839, n_126, n_96, n_120);
  and g9367 (n_3840, n_210, n735, n752);
  and g9368 (n_3841, n768, n773);
  and g9369 (n_3842, n775, n777);
  and g9370 (n786, n_3839, n_3840, n_3841, n_3842);
  and g9371 (n_3843, n_181, n_321, n_203);
  and g9372 (n_3844, n578, n_103, n789);
  and g9373 (n_3845, n805, n806, n807);
  and g9374 (n_3846, n808, n625, n815);
  and g9375 (n826, n_3843, n_3844, n_3845, n_3846);
  and g9376 (n558, n_208, n_129, n_116, n555);
  and g9377 (n_3847, n_196, n_206);
  and g9378 (n_3848, n_222, n_114);
  and g9379 (n_3849, n_202, n_131);
  and g9380 (n_3850, n_128, n_212);
  and g9381 (n735, n_3847, n_3848, n_3849, n_3850);
  and g9382 (n_3851, n_150, n_183, n_96);
  and g9383 (n_3852, n_213, n_209, n_131);
  and g9384 (n_3853, n792, n648);
  and g9385 (n_3854, n794, n796);
  and g9386 (n805, n_3851, n_3852, n_3853, n_3854);
  nor g9387 (n1577, n1571, n1572, n1573, n1574);
  nor g9388 (n1835, n1829, n1830, n1831, n1832);
  nor g9389 (n1708, n1702, n1703, n1704, n1705);
  nor g9390 (n1633, n1627, n1628, n1629, n1630);
  nor g9391 (n1640, n1634, n1635, n1636, n1637);
  nor g9392 (n1526, n1520, n1521, n1522, n1523);
  nor g9393 (n1862, n1856, n1857, n1858, n1859);
  nor g9394 (n1757, n1751, n1752, n1753, n1754);
  nor g9395 (n1497, n1491, n1492, n1493, n1494);
  nor g9396 (n1584, n1578, n1579, n1580, n1581);
  nor g9397 (n1591, n1585, n1586, n1587, n1588);
  nor g9398 (n1569, n1563, n1564, n1565, n1566);
  nor g9399 (n1081, n1075, n1076, n1077, n1078);
  nor g9400 (n1088, n1082, n1083, n1084, n1085);
  nor g9401 (n1210, n1204, n1205, n1206, n1207);
  nor g9402 (n1302, n1296, n1297, n1298, n1299);
  and g9403 (n1680, n_3855, n_3856, n_3857, n665);
  not g9404 (n_3855, n1676);
  not g9405 (n_3856, n847);
  not g9406 (n_3857, n1677);
  nor g9407 (n1764, n1758, n1759, n1760, n1761);
  nor g9408 (n1771, n1765, n1766, n1767, n1768);
  and g9409 (n_3858, n_139, n_264, n_143);
  and g9410 (n_3859, n_201, n_147, n_116);
  and g9411 (n_3860, n_99, n1457, n421);
  and g9412 (n_3861, n1468, n373, n1476);
  and g9413 (n1487, n_3858, n_3859, n_3860, n_3861);
  and g9414 (n_3862, n_261, n_143, n_141);
  and g9415 (n_3863, n_176, n923, n938);
  and g9416 (n_3864, n944, n325, n946);
  and g9417 (n_3865, n948, n496, n573);
  and g9418 (n959, n_3862, n_3863, n_3864, n_3865);
  and g9419 (n_3866, n_208, n_229, n_178);
  and g9420 (n_3867, n614, n967);
  and g9421 (n_3868, n975, n141);
  and g9422 (n_3869, n979, n999);
  and g9423 (n1007, n_3866, n_3867, n_3868, n_3869);
  nor g9424 (n1688, n1682, n1683, n1684, n1685);
  nor g9425 (n1695, n1689, n1690, n1691, n1692);
  nor g9426 (n1721, n1715, n1716, n1717, n1718);
  nor g9427 (n1815, n1809, n1810, n1811, n1812);
  nor g9428 (n1823, n1817, n1818, n1819, n1820);
  and g9429 (n_3870, n_263, n_114, n_117, n_96);
  and g9430 (n_3871, n_107, n1104, n311, n1108);
  and g9431 (n_3872, n1115, n325, n558);
  and g9432 (n_3873, n609, n1116, n1117);
  and g9433 (n1130, n_3870, n_3871, n_3872, n_3873);
  and g9434 (n_3874, n_261, n_263, n_197);
  and g9435 (n_3875, n_138, n_146);
  and g9436 (n_3876, n_176, n_102);
  and g9437 (n_3877, n_129, n809);
  and g9438 (n1457, n_3874, n_3875, n_3876, n_3877);
  and g9439 (n_3878, n_91, n_194, n_134);
  and g9440 (n_3879, n_205, n_229);
  and g9441 (n_3880, n_103, n_218);
  and g9442 (n_3881, n_186, n_200);
  and g9443 (n1476, n_3878, n_3879, n_3880, n_3881);
  nor g9444 (n1511, n1505, n1506, n1507, n1508);
  nor g9445 (n1518, n1512, n1513, n1514, n1515);
  nor g9446 (n1364, n1358, n1359, n1360, n1361);
  nor g9447 (n1389, n1383, n1384, n1385, n1386);
  nor g9448 (n1396, n1390, n1391, n1392, n1393);
  nor g9449 (n1404, n1398, n1399, n1400, n1401);
  nor g9450 (n1256, n1250, n1251, n1252, n1253);
  nor g9451 (n1263, n1257, n1258, n1259, n1260);
  and g9452 (n_3882, n_88, n_178);
  and g9453 (n_3883, n_131, n926);
  and g9454 (n_3884, n930, n931);
  and g9455 (n_3885, n562, n638);
  and g9456 (n938, n_3882, n_3883, n_3884, n_3885);
  and g9457 (n_3886, n_183, n_218);
  and g9458 (n_3887, n_189, n_86);
  and g9459 (n975, n969, n970, n_3886, n_3887);
  and g9460 (n_3888, n_199, n_263);
  and g9461 (n999, n_101, n_191, n995, n_3888);
  nor g9462 (n1334, n1328, n1329, n1330, n1331);
  nor g9463 (n1341, n1335, n1336, n1337, n1338);
  nor g9464 (n1249, n1242, n1243, n1245, n1246);
  nor g9465 (n1904, n1898, n1899, n1900, n1901);
  nor g9466 (n1911, n1905, n1906, n1907, n1908);
  and g9467 (n_3889, n_196, n_203);
  and g9468 (n_3890, n_227, n_132);
  and g9469 (n_3891, n_136, n_100);
  and g9470 (n_3892, n460, n_224);
  and g9471 (n1115, n_3889, n_3890, n_3891, n_3892);
  nor g9472 (n1448, n1442, n1443, n1444, n1445);
  nor g9473 (n1376, n1369, n1370, n1372, n1373);
  nor g9474 (n1349, n1343, n1344, n1345, n1346);
  nor g9475 (n1897, n1891, n1892, n1893, n1894);
  nor g9476 (n1976, n1970, n1971, n1972, n1973);
  nor g9477 (n1983, n1977, n1978, n1979, n1980);
  and g9478 (n_3893, n_193, n_131, n_90);
  and g9479 (n_3894, n1145, n1162, n141);
  and g9480 (n_3895, n366, n505, n451);
  and g9481 (n_3896, n760, n1165);
  and g9482 (n1175, n_3893, n_3894, n_3895, n_3896);
  and g9483 (n1939, n_3897, n_3898, n_3899, n1009);
  not g9484 (n_3897, n1935);
  not g9485 (n_3898, n1244);
  not g9486 (n_3899, n1936);
  and g9487 (n_3900, n_190, n_183, n_104);
  and g9488 (n_3901, n_137, n_89, n_109);
  and g9489 (n_3902, n_144, n1134, n1108);
  and g9490 (n_3903, n314, n646, n948);
  and g9491 (n1145, n_3900, n_3901, n_3902, n_3903);
  nor g9492 (n2007, n2001, n2002, n2003, n2004);
  nor g9493 (n1949, n1943, n1944, n1945, n1946);
  nor g9494 (n1956, n1950, n1951, n1952, n1953);
  nor g9495 (n_3907, n2025, n2026);
  and g9496 (n2051, n_3904, n_3905, n_3906, n_3907);
  not g9497 (n_3904, n2027);
  not g9498 (n_3905, n2046);
  not g9499 (n_3906, n2047);
  and g9500 (n_3908, n_225, n_147, n_111, n_189);
  and g9501 (n_3909, n_92, n_101, n3231, n210);
  and g9502 (n_3910, n4002, n753, n249);
  and g9503 (n_3911, n2276, n637, n2340);
  and g9504 (n4015, n_3908, n_3909, n_3910, n_3911);
  and g9505 (n4002, n_143, n_201, n_84, n_211);
  nor g9506 (n3910, n3897, n3898, n3899, n3909);
  and g9507 (n_3912, n_190, n_208, n_222);
  and g9508 (n_3913, n_226, n976, n2432);
  and g9509 (n_3914, n3883, n1476, n815);
  and g9510 (n_3915, n316, n555);
  and g9511 (n3893, n_3912, n_3913, n_3914, n_3915);
  and g9512 (n_3916, n_105, n_114);
  and g9513 (n_3917, n_147, n_104);
  and g9514 (n_3918, n753, n457);
  and g9515 (n_3919, n236, n2433);
  and g9516 (n3883, n_3916, n_3917, n_3918, n_3919);
  nor g9517 (n3922, n3916, n3917, n3918, n3921);
  nor g9518 (n3937, n3931, n3932, n3933, n3936);
  and g9519 (n_3920, n_190, n_228, n_87);
  and g9520 (n_3921, n_179, n_227, n_217);
  and g9521 (n_3922, n_182, n3699, n4037);
  and g9522 (n_3923, n805, n416, n608);
  and g9523 (n4048, n_3920, n_3921, n_3922, n_3923);
  and g9524 (n_3924, n_97, n_85);
  and g9525 (n_3925, n_119, n_144);
  and g9526 (n4037, n346, n_210, n_3924, n_3925);
  nor g9527 (n4070, n4064, n4065, n4066, n4069);
  nor g9528 (n4085, n4079, n4080, n4081, n4084);
  and g9529 (n_3926, n_127, n_143, n_149, n_207);
  and g9530 (n_3927, n_101, n_184, n355, n735);
  and g9531 (n_3928, n1468, n2196, n946);
  and g9532 (n_3929, n397, n2340, n3657);
  and g9533 (n4175, n_3926, n_3927, n_3928, n_3929);
  nor g9534 (n4192, n4186, n4187, n4188, n4191);
  nor g9535 (n4207, n4201, n4202, n4203, n4206);
  and g9536 (n_3930, n_262, n_108, n_99);
  and g9537 (n_3931, n2418, n644, n752);
  and g9538 (n_3932, n975, n2464, n301);
  and g9539 (n_3933, n346, n496);
  and g9540 (n4291, n_3930, n_3931, n_3932, n_3933);
  nor g9541 (n4363, n4357, n4358, n4359, n4362);
  nor g9542 (n4346, n4340, n4341, n4342, n4345);
  nor g9543 (n4329, n4323, n4324, n4325, n4328);
  nor g9544 (n4302, n4296, n4297, n4298, n4301);
  and g9545 (n_3934, n_126, n_178, n_213, n_99);
  and g9546 (n_3935, n369, n4002, n3243);
  and g9547 (n_3936, n3883, n314, n2317);
  and g9548 (n_3937, n4392, n189, n807);
  and g9549 (n4404, n_3934, n_3935, n_3936, n_3937);
  nor g9550 (n4415, n4409, n4410, n4411, n4414);
  nor g9551 (n4453, n4447, n4448, n4449, n4452);
  and g9552 (n_3938, n_88, n_215, n_104);
  and g9553 (n_3939, n_103, n_89, n_191);
  and g9554 (n_3940, n4513, n3259, n2458);
  and g9555 (n_3941, n253, n970);
  and g9556 (n4523, n_3938, n_3939, n_3940, n_3941);
  and g9557 (n_3942, n_204, n976, n369);
  and g9558 (n_3943, n156, n2340);
  and g9559 (n_3944, n2421, n586);
  and g9560 (n_3945, n316, n1117);
  and g9561 (n4513, n_3942, n_3943, n_3944, n_3945);
  nor g9562 (n4542, n4536, n4537, n4538, n4541);
  nor g9563 (n4579, n4573, n4574, n4575, n4578);
  and g9564 (n_3946, n_225, n_105, n1090);
  and g9565 (n_3947, n_132, n_94, n_108);
  and g9566 (n_3948, n_144, n4513, n809);
  and g9567 (n_3949, n4392, n931, n2281);
  and g9568 (n4702, n_3946, n_3947, n_3948, n_3949);
  nor g9569 (n4643, n4637, n4638, n4639, n4642);
  and g9570 (n_3950, n_223, n_190, n_122);
  and g9571 (n_3951, n_201, n_115, n_142);
  and g9572 (n_3952, n_210, n4726, n3678);
  and g9573 (n_3953, n979, n961, n2342);
  and g9574 (n4737, n_3950, n_3951, n_3952, n_3953);
  and g9575 (n_3954, n_139, n_149, n_218);
  and g9576 (n_3955, n_121, n_113, n_131);
  and g9577 (n_3956, n_129, n165);
  and g9578 (n_3957, n609, n2181);
  and g9579 (n4726, n_3954, n_3955, n_3956, n_3957);
  nor g9580 (n4783, n4777, n4778, n4779, n4782);
  and g9581 (n_3958, n_134, n_205, n_124, n_96);
  and g9582 (n_3959, n_121, n_189, n_191);
  and g9583 (n_3960, n3259, n2432, n3231);
  and g9584 (n_3961, n204, n757, n809);
  and g9585 (n4829, n_3958, n_3959, n_3960, n_3961);
  nor g9586 (n4857, n4851, n4852, n4853, n4856);
  nor g9587 (n4838, n4832, n4833, n4834, n4837);
  and g9588 (n_3962, n_183, n_110, n_185);
  and g9589 (n_3963, n977, n3259, n1104);
  and g9590 (n_3964, n3666, n210, n505);
  and g9591 (n_3965, n476, n259, n655);
  and g9592 (n4911, n_3962, n_3963, n_3964, n_3965);
  nor g9593 (n4937, n4931, n4932, n4933, n4936);
  and g9594 (n_3966, n_192, n453);
  and g9595 (n_3967, n636, n3734);
  and g9596 (n_3968, n499, n911);
  and g9597 (n4993, n969, n_3966, n_3967, n_3968);
  and g9598 (n_3969, n_139, n_95, n_83);
  and g9599 (n_3970, n380, n2250);
  and g9600 (n_3971, n4037, n946);
  and g9601 (n_3972, n2367, n5055);
  and g9602 (n5063, n_3969, n_3970, n_3971, n_3972);
  and g9603 (n_3973, n_193, n_124);
  and g9604 (n5055, n_115, n_98, n_106, n_3973);
  nor g9605 (n5078, n5072, n5073, n5074, n5077);
  and g9606 (n_3974, n_199, n_222, n_85, n_104);
  and g9607 (n_3975, n_142, n_195, n_109, n3699);
  and g9608 (n_3976, n980, n2178, n311);
  and g9609 (n_3977, n4002, n156, n5125);
  and g9610 (n5138, n_3974, n_3975, n_3976, n_3977);
  and g9611 (n_3978, n_147, n_200);
  and g9612 (n5125, n_141, n_108, n_214, n_3978);
  nor g9613 (n5146, n5140, n5141, n5142, n5145);
  and g9614 (n_3979, n_228, n_192, n_207, n_195);
  and g9615 (n_3980, n_145, n_100, n_93, n3259);
  and g9616 (n_3981, n983, n1457, n2190, n967);
  and g9617 (n_3982, n473, n2367, n2433);
  and g9618 (n5202, n_3979, n_3980, n_3981, n_3982);
  and g9619 (n_3983, n_321, n_228, n_205);
  and g9620 (n_3984, n_133, n_120, n_145);
  and g9621 (n_3985, n1115, n2375, n5055);
  and g9622 (n_3986, n344, n970, n5247);
  and g9623 (n5258, n_3983, n_3984, n_3985, n_3986);
  and g9624 (n5247, n_140, n_187, n_191, n1145);
  and g9625 (n_3987, n_219, n_215, n_116);
  and g9626 (n_3988, n3702, n475, n233);
  and g9627 (n_3989, n5125, n2252);
  and g9628 (n_3990, n638, n2313);
  and g9629 (n5303, n_3987, n_3988, n_3989, n_3990);
  and g9630 (n_3991, n_135, n_206, n_180);
  and g9631 (n_3992, n_115, n_83, n980);
  and g9632 (n_3993, n571, n3243, n259);
  and g9633 (n_3994, n906, n158, n775);
  and g9634 (n5344, n_3991, n_3992, n_3993, n_3994);
  and g9635 (n_3995, n_127, n_204, n_115);
  and g9636 (n_3996, n_118, n_100, n3675);
  and g9637 (n_3997, n986, n1108, n1152);
  and g9638 (n_3998, n608, n588, n2170);
  and g9639 (n5367, n_3995, n_3996, n_3997, n_3998);
  and g9640 (n_3999, n_117, n_179, n_218);
  and g9641 (n_4000, n_84, n_116, n_90);
  and g9642 (n_4001, n_86, n938, n2540);
  and g9643 (n_4002, n373, n4392, n5247);
  and g9644 (n5389, n_3999, n_4000, n_4001, n_4002);
  and g9645 (n_4003, n_260, n_138, n_137, n_132);
  and g9646 (n_4004, n_185, n_118, n_108);
  and g9647 (n_4005, n369, n4726, n502);
  and g9648 (n_4006, n999, n189, n459);
  and g9649 (n5412, n_4003, n_4004, n_4005, n_4006);
  and g9650 (n_4007, n_200, n_195);
  and g9651 (n5427, n444, n489, n3617, n_4007);
endmodule

