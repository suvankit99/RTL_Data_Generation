
module int2float(\B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6]
     , \B[7] , \B[8] , \B[9] , \B[10] , \M[0] , \M[1] , \M[2] , \M[3] ,
     \E[0] , \E[1] , \E[2] );
  input \B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] ,
       \B[8] , \B[9] , \B[10] ;
  output \M[0] , \M[1] , \M[2] , \M[3] , \E[0] , \E[1] , \E[2] ;
  wire \B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] ,
       \B[8] , \B[9] , \B[10] ;
  wire \M[0] , \M[1] , \M[2] , \M[3] , \E[0] , \E[1] , \E[2] ;
  wire n19, n20, n21, n22, n23, n24, n25, n26;
  wire n27, n28, n29, n30, n31, n32, n33, n34;
  wire n35, n36, n37, n38, n39, n40, n41, n42;
  wire n43, n44, n45, n46, n47, n48, n49, n50;
  wire n51, n52, n53, n54, n55, n56, n57, n58;
  wire n59, n60, n61, n62, n63, n64, n65, n66;
  wire n67, n68, n69, n70, n71, n72, n73, n74;
  wire n75, n76, n77, n79, n80, n81, n82, n83;
  wire n84, n85, n86, n87, n88, n89, n90, n91;
  wire n92, n93, n96, n97, n98, n99, n100, n101;
  wire n102, n103, n104, n105, n106, n107, n108, n109;
  wire n110, n111, n112, n113, n114, n115, n116, n117;
  wire n118, n119, n120, n121, n122, n123, n124, n125;
  wire n126, n127, n128, n129, n130, n131, n132, n133;
  wire n134, n135, n138, n139, n140, n141, n144, n145;
  wire n149, n150, n151, n152, n153, n154, n155, n156;
  wire n157, n158, n159, n160, n161, n162, n163, n164;
  wire n165, n166, n167, n168, n169, n170, n171, n172;
  wire n173, n174, n175, n176, n177, n178, n179, n180;
  wire n181, n182, n183, n184, n185, n186, n187, n188;
  wire n189, n190, n191, n192, n193, n194, n195, n196;
  wire n197, n198, n199, n200, n201, n202, n203, n204;
  wire n205, n206, n207, n208, n213, n214, n215, n216;
  wire n220, n221, n222, n223, n224, n225, n226, n227;
  wire n228, n229, n230, n231, n232, n233, n238, n239;
  wire n240, n241, n246, n247, n248, n249, n250, n252;
  wire n253, n258, n259, n260, n263, n264, n265, n266;
  wire n267, n268, n269, n270, n274, n275, n_2, n_5;
  wire n_6, n_7, n_8, n_10, n_11, n_12, n_13, n_15;
  wire n_16, n_18, n_19, n_20, n_22, n_23, n_25, n_26;
  wire n_27, n_29, n_30, n_31, n_32, n_33, n_34, n_35;
  wire n_36, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_50, n_51, n_52, n_53;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93;
  wire n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_173, n_174, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_202, n_203, n_204;
  wire n_207, n_208, n_209, n_211, n_212, n_213, n_217, n_218;
  not g1 (n_2, \B[1] );
  and g2 (n19, n_2, \B[4] );
  not g3 (n_5, \B[4] );
  not g4 (n_6, \B[8] );
  and g5 (n20, n_5, n_6);
  not g6 (n_7, n19);
  not g7 (n_8, n20);
  and g8 (n21, n_7, n_8);
  not g9 (n_10, n21);
  and g10 (n22, \B[0] , n_10);
  and g11 (n23, \B[1] , \B[4] );
  not g12 (n_11, \B[0] );
  and g13 (n24, n_11, n23);
  not g14 (n_12, n22);
  not g15 (n_13, n24);
  and g16 (n25, n_12, n_13);
  not g17 (n_15, \B[6] );
  not g18 (n_16, n25);
  and g19 (n26, n_15, n_16);
  not g20 (n_18, \B[7] );
  and g21 (n27, n_18, n26);
  and g22 (n28, \B[4] , \B[8] );
  not g23 (n_19, n27);
  not g24 (n_20, n28);
  and g25 (n29, n_19, n_20);
  not g26 (n_22, \B[5] );
  not g27 (n_23, n29);
  and g28 (n30, n_22, n_23);
  and g29 (n31, n_5, \B[7] );
  not g30 (n_25, \B[2] );
  and g31 (n32, \B[1] , n_25);
  and g32 (n33, \B[5] , n_18);
  and g33 (n34, n32, n33);
  not g34 (n_26, n31);
  not g35 (n_27, n34);
  and g36 (n35, n_26, n_27);
  not g37 (n_29, n35);
  and g38 (n36, \B[3] , n_29);
  and g39 (n37, \B[4] , \B[7] );
  not g40 (n_30, \B[3] );
  and g41 (n38, n_30, n37);
  not g42 (n_31, n36);
  not g43 (n_32, n38);
  and g44 (n39, n_31, n_32);
  not g45 (n_33, n39);
  and g46 (n40, n_6, n_33);
  and g47 (n41, \B[5] , \B[8] );
  and g48 (n42, n_5, n41);
  not g49 (n_34, n40);
  not g50 (n_35, n42);
  and g51 (n43, n_34, n_35);
  not g52 (n_36, n30);
  and g53 (n44, n_36, n43);
  not g54 (n_38, \B[9] );
  not g55 (n_39, n44);
  and g56 (n45, n_38, n_39);
  and g57 (n46, \B[4] , n_6);
  and g58 (n47, n_30, n46);
  and g59 (n48, n_5, n_18);
  not g60 (n_40, n47);
  not g61 (n_41, n48);
  and g62 (n49, n_40, n_41);
  not g63 (n_42, n49);
  and g64 (n50, n_25, n_42);
  and g65 (n51, \B[1] , n50);
  and g66 (n52, n_2, \B[2] );
  and g67 (n53, n_18, n_6);
  and g68 (n54, n52, n53);
  not g69 (n_43, n54);
  and g70 (n55, n_38, n_43);
  not g71 (n_44, n51);
  and g72 (n56, n_44, n55);
  not g73 (n_45, n56);
  and g74 (n57, n_15, n_45);
  and g75 (n58, \B[5] , n57);
  and g76 (n59, \B[6] , \B[9] );
  and g77 (n60, n_22, n59);
  not g78 (n_46, n58);
  not g79 (n_47, n60);
  and g80 (n61, n_46, n_47);
  not g81 (n_48, n45);
  and g82 (n62, n_48, n61);
  not g83 (n_50, \B[10] );
  not g84 (n_51, n62);
  and g85 (n63, n_50, n_51);
  and g86 (n64, n_25, \B[3] );
  and g87 (n65, \B[2] , n_30);
  not g88 (n_52, n64);
  not g89 (n_53, n65);
  and g90 (n66, n_52, n_53);
  not g91 (n_54, n66);
  and g92 (n67, n_38, n_54);
  and g93 (n68, n_6, n67);
  not g94 (n_55, n68);
  and g95 (n69, n_50, n_55);
  not g96 (n_56, n69);
  and g97 (n70, n_18, n_56);
  and g98 (n71, \B[9] , \B[10] );
  and g99 (n72, \B[8] , n71);
  not g100 (n_57, n70);
  not g101 (n_58, n72);
  and g102 (n73, n_57, n_58);
  not g103 (n_59, n73);
  and g104 (n74, \B[6] , n_59);
  and g105 (n75, n_15, \B[10] );
  and g106 (n76, \B[7] , n75);
  not g107 (n_60, n74);
  not g108 (n_61, n76);
  and g109 (n77, n_60, n_61);
  not g110 (n_62, n77);
  or g111 (\M[0] , n63, n_62);
  and g112 (n79, n_5, n_38);
  and g113 (n80, n_25, n_18);
  not g114 (n_63, n79);
  not g115 (n_64, n80);
  and g116 (n81, n_63, n_64);
  not g117 (n_65, n81);
  and g118 (n82, n_2, n_65);
  and g119 (n83, \B[1] , \B[2] );
  and g120 (n84, \B[0] , n83);
  and g121 (n85, n_11, n_25);
  not g122 (n_66, n84);
  not g123 (n_67, n85);
  and g124 (n86, n_66, n_67);
  not g125 (n_68, n86);
  and g126 (n87, n_18, n_68);
  and g127 (n88, \B[4] , n87);
  and g128 (n89, \B[8] , n_38);
  not g129 (n_69, n88);
  not g130 (n_70, n89);
  and g131 (n90, n_69, n_70);
  not g132 (n_71, n82);
  and g133 (n91, n_71, n90);
  not g134 (n_72, n91);
  and g135 (n92, n_15, n_72);
  and g136 (n93, \B[3] , \B[4] );
  not g137 (n_73, n93);
  and g141 (n97, n_18, \B[9] );
  not g142 (n_74, n96);
  not g143 (n_75, n97);
  and g144 (n98, n_74, n_75);
  not g145 (n_76, n92);
  and g146 (n99, n_76, n98);
  not g147 (n_77, n99);
  and g148 (n100, n_22, n_77);
  and g149 (n101, n_6, n_38);
  and g150 (n102, \B[4] , n101);
  and g151 (n103, n_15, n_18);
  and g152 (n104, n_5, n103);
  not g153 (n_78, n102);
  not g154 (n_79, n104);
  and g155 (n105, n_78, n_79);
  not g156 (n_80, n105);
  and g157 (n106, \B[2] , n_80);
  and g158 (n107, \B[1] , n106);
  and g159 (n108, \B[7] , n_38);
  and g160 (n109, n46, n108);
  not g161 (n_81, n107);
  not g162 (n_82, n109);
  and g163 (n110, n_81, n_82);
  not g164 (n_83, n110);
  and g165 (n111, \B[3] , n_83);
  and g166 (n112, \B[4] , n89);
  and g167 (n113, \B[7] , \B[9] );
  not g168 (n_84, n112);
  not g169 (n_85, n113);
  and g170 (n114, n_84, n_85);
  not g171 (n_86, n114);
  and g172 (n115, \B[6] , n_86);
  not g173 (n_87, n111);
  not g174 (n_88, n115);
  and g175 (n116, n_87, n_88);
  not g176 (n_89, n116);
  and g177 (n117, \B[5] , n_89);
  and g178 (n118, n_5, n89);
  not g179 (n_90, n118);
  and g180 (n119, n_75, n_90);
  not g181 (n_91, n119);
  and g182 (n120, n_15, n_91);
  not g183 (n_92, n117);
  not g184 (n_93, n120);
  and g185 (n121, n_92, n_93);
  not g186 (n_94, n100);
  and g187 (n122, n_94, n121);
  not g188 (n_95, n122);
  and g189 (n123, n_50, n_95);
  and g190 (n124, \B[6] , n_38);
  and g191 (n125, n_5, n124);
  and g192 (n126, \B[5] , n_15);
  and g193 (n127, n_30, n126);
  not g194 (n_96, n125);
  not g195 (n_97, n127);
  and g196 (n128, n_96, n_97);
  not g197 (n_98, n128);
  and g198 (n129, n_25, n_98);
  and g199 (n130, n_2, n126);
  not g200 (n_99, n130);
  and g201 (n131, n_96, n_99);
  not g202 (n_100, n131);
  and g203 (n132, n_30, n_100);
  and g204 (n133, \B[2] , \B[3] );
  and g205 (n134, \B[4] , n124);
  and g206 (n135, n133, n134);
  not g213 (n_104, n138);
  and g214 (n139, n_18, n_104);
  not g215 (n_105, n75);
  not g216 (n_106, n139);
  and g217 (n140, n_105, n_106);
  not g218 (n_107, n140);
  and g219 (n141, n_6, n_107);
  not g223 (n_108, n141);
  not g224 (n_109, n144);
  and g225 (n145, n_108, n_109);
  not g226 (n_110, n123);
  and g227 (\M[1] , n_110, n145);
  and g231 (n150, n_5, \B[5] );
  and g232 (n151, \B[3] , n150);
  not g233 (n_111, n149);
  not g234 (n_112, n151);
  and g235 (n152, n_111, n_112);
  not g236 (n_113, n152);
  and g237 (n153, \B[1] , n_113);
  and g238 (n154, n_5, n_15);
  and g239 (n155, \B[0] , \B[1] );
  not g240 (n_114, n155);
  and g241 (n156, \B[4] , n_114);
  and g242 (n157, \B[3] , n156);
  not g243 (n_115, n154);
  not g244 (n_116, n157);
  and g245 (n158, n_115, n_116);
  not g246 (n_117, n158);
  and g247 (n159, n_22, n_117);
  not g248 (n_118, n153);
  not g249 (n_119, n159);
  and g250 (n160, n_118, n_119);
  not g251 (n_120, n160);
  and g252 (n161, \B[2] , n_120);
  and g253 (n162, \B[3] , n_15);
  and g254 (n163, n_25, n162);
  and g255 (n164, n_30, \B[5] );
  not g256 (n_121, n163);
  not g257 (n_122, n164);
  and g258 (n165, n_121, n_122);
  not g259 (n_123, n165);
  and g260 (n166, \B[4] , n_123);
  not g261 (n_124, n161);
  not g262 (n_125, n166);
  and g263 (n167, n_124, n_125);
  not g264 (n_126, n167);
  and g265 (n168, n_18, n_126);
  and g266 (n169, n_22, \B[6] );
  and g267 (n170, \B[2] , n169);
  not g268 (n_127, n170);
  and g269 (n171, n_99, n_127);
  not g270 (n_128, n171);
  and g271 (n172, \B[4] , n_128);
  and g272 (n173, \B[3] , n172);
  and g273 (n174, \B[5] , n_73);
  and g274 (n175, \B[6] , n174);
  not g275 (n_129, n173);
  not g276 (n_130, n175);
  and g277 (n176, n_129, n_130);
  not g278 (n_131, n168);
  and g279 (n177, n_131, n176);
  not g280 (n_132, n177);
  and g281 (n178, n_6, n_132);
  and g282 (n179, n_15, \B[7] );
  and g283 (n180, \B[3] , n179);
  and g284 (n181, \B[6] , n_18);
  and g285 (n182, n_25, n181);
  not g286 (n_133, n180);
  not g287 (n_134, n182);
  and g288 (n183, n_133, n_134);
  not g289 (n_135, n183);
  and g290 (n184, \B[5] , n_135);
  and g291 (n185, \B[4] , n184);
  and g292 (n186, \B[4] , \B[5] );
  not g293 (n_136, n186);
  and g294 (n187, \B[7] , n_136);
  and g295 (n188, \B[6] , n187);
  not g296 (n_137, n185);
  not g297 (n_138, n188);
  and g298 (n189, n_137, n_138);
  not g299 (n_139, n178);
  and g300 (n190, n_139, n189);
  not g301 (n_140, n190);
  and g302 (n191, n_38, n_140);
  and g303 (n192, \B[4] , \B[6] );
  and g304 (n193, n33, n192);
  not g305 (n_141, n179);
  not g306 (n_142, n193);
  and g307 (n194, n_141, n_142);
  not g308 (n_143, n194);
  and g309 (n195, \B[8] , n_143);
  not g310 (n_144, n191);
  not g311 (n_145, n195);
  and g312 (n196, n_144, n_145);
  not g313 (n_146, n196);
  and g314 (n197, n_50, n_146);
  and g315 (n198, \B[8] , \B[10] );
  and g316 (n199, n_6, \B[9] );
  and g317 (n200, \B[5] , n199);
  not g318 (n_147, n198);
  not g319 (n_148, n200);
  and g320 (n201, n_147, n_148);
  not g321 (n_149, n201);
  and g322 (n202, \B[7] , n_149);
  and g323 (n203, \B[6] , n202);
  and g324 (n204, \B[5] , \B[7] );
  not g325 (n_150, n204);
  and g326 (n205, \B[8] , n_150);
  not g327 (n_151, n205);
  and g328 (n206, n_50, n_151);
  not g329 (n_152, n206);
  and g330 (n207, \B[9] , n_152);
  not g331 (n_153, n203);
  not g332 (n_154, n207);
  and g333 (n208, n_153, n_154);
  not g334 (n_155, n208);
  or g335 (\M[2] , n197, n_155);
  and g340 (n214, n_22, n20);
  and g341 (n215, n103, n214);
  not g342 (n_156, n213);
  not g343 (n_157, n215);
  and g344 (n216, n_156, n_157);
  and g350 (n220, \B[5] , \B[6] );
  and g351 (n221, \B[4] , n_18);
  and g352 (n222, n220, n221);
  and g353 (n223, n_22, n_15);
  and g354 (n224, n155, n223);
  not g355 (n_160, n222);
  not g356 (n_161, n224);
  and g357 (n225, n_160, n_161);
  not g358 (n_162, n225);
  and g359 (n226, \B[3] , n_162);
  and g360 (n227, \B[2] , n226);
  not g361 (n_163, n181);
  and g362 (n228, n_5, n_163);
  not g363 (n_164, n126);
  and g364 (n229, n_18, n_164);
  not g365 (n_165, n229);
  and g366 (n230, n_30, n_165);
  not g367 (n_166, n220);
  and g368 (n231, \B[7] , n_166);
  not g369 (n_167, n83);
  and g370 (n232, n_15, n_167);
  and g371 (n233, \B[5] , n232);
  not g382 (n_173, n238);
  and g383 (n239, n_6, n_173);
  and g384 (n240, \B[3] , \B[8] );
  not g385 (n_174, n240);
  and g386 (n241, n_53, n_174);
  and g393 (n247, \B[7] , n220);
  not g394 (n_176, n247);
  and g395 (n248, \B[9] , n_176);
  not g396 (n_177, n246);
  not g397 (n_178, n248);
  and g398 (n249, n_177, n_178);
  not g399 (n_179, n239);
  and g400 (n250, n_179, n249);
  or g401 (\E[0] , \B[10] , n250);
  and g402 (n252, \B[6] , \B[8] );
  and g403 (n253, n204, n252);
  not g409 (n_180, n253);
  not g410 (n_181, n258);
  and g411 (n259, n_180, n_181);
  not g412 (n_182, n259);
  and g413 (n260, \B[2] , n_182);
  not g417 (n_183, n260);
  not g418 (n_184, n263);
  and g419 (n264, n_183, n_184);
  not g420 (n_185, n264);
  and g421 (n265, \B[4] , n_185);
  and g422 (n266, n133, n192);
  not g423 (n_186, n266);
  and g424 (n267, \B[5] , n_186);
  not g425 (n_187, n169);
  not g426 (n_188, n267);
  and g427 (n268, n_187, n_188);
  not g428 (n_189, n268);
  and g429 (n269, n_18, n_189);
  and g430 (n270, n_6, n269);
  and g436 (n274, \B[2] , n93);
  and g437 (n275, n220, n274);
  and g444 (n144, n89, \B[7] , \B[6] , \B[10] );
  and g445 (n138, n_202, n_203, n_204, n_50);
  not g446 (n_202, n129);
  not g447 (n_203, n132);
  not g448 (n_204, n135);
  and g449 (n96, n_6, n_38, \B[7] , n_73);
  and g450 (n149, \B[4] , n_15, \B[0] , n_30);
  or g451 (\M[3] , \B[10] , \B[9] , \B[3] , n216);
  and g454 (n_207, n_25, \B[6] );
  and g455 (n213, \B[7] , \B[5] , n28, n_207);
  and g456 (n_209, n_208, \B[4] );
  not g457 (n_208, n241);
  and g459 (n246, \B[5] , \B[6] , n_209, n108);
  nor g460 (n_212, n227, n228);
  nor g461 (n_213, n230, n231);
  and g462 (n238, n_211, n_38, n_212, n_213);
  not g463 (n_211, n233);
  or g464 (\E[1] , \B[9] , \B[10] , n265, n270);
  and g467 (n263, \B[8] , n204, \B[3] , \B[6] );
  and g469 (n_217, \B[3] , n_6);
  and g470 (n258, n_22, n_18, n155, n_217);
  or g471 (\E[2] , n_218, \B[10] , \B[9] , n275);
  not g472 (n_218, n53);
endmodule

