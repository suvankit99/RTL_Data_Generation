
module log2(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] ,
     \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14]
     , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
     \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
     \a[29] , \a[30] , \a[31] , \result[0] , \result[1] , \result[2] ,
     \result[3] , \result[4] , \result[5] , \result[6] , \result[7] ,
     \result[8] , \result[9] , \result[10] , \result[11] , \result[12]
     , \result[13] , \result[14] , \result[15] , \result[16] ,
     \result[17] , \result[18] , \result[19] , \result[20] ,
     \result[21] , \result[22] , \result[23] , \result[24] ,
     \result[25] , \result[26] , \result[27] , \result[28] ,
     \result[29] , \result[30] , \result[31] );
  input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4]
       , \result[5] , \result[6] , \result[7] , \result[8] , \result[9]
       , \result[10] , \result[11] , \result[12] , \result[13] ,
       \result[14] , \result[15] , \result[16] , \result[17] ,
       \result[18] , \result[19] , \result[20] , \result[21] ,
       \result[22] , \result[23] , \result[24] , \result[25] ,
       \result[26] , \result[27] , \result[28] , \result[29] ,
       \result[30] , \result[31] ;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] ;
  wire \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
       \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
       \result[10] , \result[11] , \result[12] , \result[13] ,
       \result[14] , \result[15] , \result[16] , \result[17] ,
       \result[18] , \result[19] , \result[20] , \result[21] ,
       \result[22] , \result[23] , \result[24] , \result[25] ,
       \result[26] , \result[27] , \result[28] , \result[29] ,
       \result[30] , \result[31] ;
  wire n65, n66, n67, n68, n69, n70, n71, n72;
  wire n73, n74, n75, n76, n77, n78, n79, n80;
  wire n81, n82, n83, n84, n85, n86, n87, n88;
  wire n89, n90, n91, n92, n93, n94, n95, n96;
  wire n97, n98, n99, n100, n101, n102, n103, n104;
  wire n105, n106, n107, n108, n109, n110, n111, n112;
  wire n113, n114, n115, n116, n117, n118, n119, n120;
  wire n121, n122, n123, n124, n125, n126, n127, n128;
  wire n129, n130, n131, n132, n133, n134, n135, n136;
  wire n137, n141, n142, n143, n144, n145, n146, n147;
  wire n148, n149, n150, n151, n152, n153, n154, n155;
  wire n156, n157, n158, n159, n160, n161, n162, n163;
  wire n164, n165, n166, n167, n168, n169, n170, n171;
  wire n172, n173, n174, n175, n176, n177, n178, n179;
  wire n187, n188, n189, n190, n191, n192, n193, n194;
  wire n198, n199, n200, n201, n202, n203, n204, n205;
  wire n206, n207, n221, n222, n223, n224, n225, n226;
  wire n227, n228, n229, n230, n231, n232, n233, n234;
  wire n235, n236, n237, n238, n239, n240, n241, n242;
  wire n243, n244, n245, n246, n247, n248, n249, n250;
  wire n251, n252, n253, n254, n255, n256, n268, n269;
  wire n270, n271, n272, n273, n274, n275, n276, n277;
  wire n278, n279, n280, n281, n282, n283, n284, n285;
  wire n286, n287, n288, n289, n290, n291, n292, n293;
  wire n294, n295, n296, n297, n298, n299, n300, n301;
  wire n302, n303, n304, n305, n306, n307, n308, n324;
  wire n325, n326, n327, n328, n329, n330, n331, n332;
  wire n333, n334, n335, n336, n337, n338, n339, n340;
  wire n341, n342, n343, n351, n352, n353, n354, n355;
  wire n356, n357, n358, n359, n362, n363, n364, n365;
  wire n366, n367, n368, n369, n370, n371, n372, n373;
  wire n374, n375, n376, n392, n393, n394, n395, n396;
  wire n397, n398, n399, n400, n401, n402, n403, n404;
  wire n405, n415, n416, n417, n418, n419, n420, n421;
  wire n422, n423, n424, n425, n426, n427, n428, n429;
  wire n430, n431, n434, n435, n436, n437, n438, n439;
  wire n448, n449, n450, n451, n452, n453, n454, n459;
  wire n460, n461, n462, n465, n466, n467, n468, n469;
  wire n470, n471, n472, n473, n474, n475, n488, n489;
  wire n490, n491, n492, n493, n494, n495, n496, n497;
  wire n503, n504, n505, n506, n507, n508, n509, n510;
  wire n511, n512, n513, n514, n515, n516, n517, n518;
  wire n519, n520, n524, n525, n526, n527, n528, n529;
  wire n530, n531, n532, n533, n534, n535, n536, n537;
  wire n538, n539, n540, n541, n556, n557, n558, n561;
  wire n562, n563, n564, n565, n566, n567, n568, n569;
  wire n570, n571, n572, n573, n587, n588, n589, n590;
  wire n591, n592, n593, n594, n595, n600, n601, n602;
  wire n603, n604, n614, n615, n616, n617, n618, n619;
  wire n620, n621, n622, n623, n624, n631, n632, n633;
  wire n634, n635, n636, n637, n638, n639, n640, n641;
  wire n642, n653, n654, n655, n656, n657, n658, n664;
  wire n665, n666, n667, n671, n672, n673, n674, n675;
  wire n688, n689, n690, n691, n692, n693, n694, n710;
  wire n711, n712, n713, n714, n715, n716, n719, n720;
  wire n721, n722, n723, n730, n731, n732, n733, n734;
  wire n735, n745, n746, n747, n751, n752, n753, n754;
  wire n757, n770, n771, n772, n773, n774, n775, n776;
  wire n777, n778, n787, n788, n789, n790, n791, n792;
  wire n793, n802, n803, n804, n805, n808, n809, n810;
  wire n811, n812, n813, n814, n815, n816, n824, n825;
  wire n826, n827, n830, n831, n832, n844, n845, n846;
  wire n847, n848, n849, n850, n851, n867, n868, n869;
  wire n872, n873, n874, n875, n876, n877, n882, n883;
  wire n884, n885, n886, n887, n888, n889, n895, n896;
  wire n897, n898, n899, n916, n917, n918, n921, n931;
  wire n932, n933, n936, n937, n940, n941, n958, n959;
  wire n960, n961, n962, n967, n968, n976, n977, n978;
  wire n979, n980, n981, n982, n988, n989, n990, n991;
  wire n992, n1008, n1009, n1010, n1011, n1012, n1020, n1021;
  wire n1024, n1025, n1029, n1039, n1040, n1044, n1045, n1046;
  wire n1047, n1060, n1061, n1062, n1063, n1064, n1065, n1069;
  wire n1070, n1071, n1072, n1073, n1080, n1084, n1085, n1100;
  wire n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108;
  wire n1109, n1119, n1120, n1121, n1126, n1127, n1128, n1129;
  wire n1130, n1131, n1132, n1135, n1138, n1139, n1140, n1141;
  wire n1142, n1143, n1154, n1155, n1158, n1159, n1160, n1161;
  wire n1162, n1163, n1178, n1179, n1180, n1181, n1182, n1183;
  wire n1184, n1185, n1202, n1203, n1204, n1205, n1206, n1211;
  wire n1216, n1219, n1220, n1221, n1235, n1236, n1237, n1240;
  wire n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252;
  wire n1253, n1254, n1255, n1264, n1268, n1269, n1270, n1271;
  wire n1272, n1273, n1274, n1291, n1292, n1293, n1294, n1305;
  wire n1306, n1307, n1308, n1313, n1314, n1315, n1323, n1324;
  wire n1328, n1329, n1330, n1331, n1332, n1333, n1345, n1346;
  wire n1347, n1364, n1365, n1366, n1367, n1368, n1369, n1372;
  wire n1378, n1379, n1380, n1384, n1387, n1388, n1389, n1390;
  wire n1391, n1392, n1393, n1394, n1407, n1408, n1409, n1419;
  wire n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1435;
  wire n1436, n1437, n1438, n1439, n1440, n1454, n1455, n1456;
  wire n1457, n1458, n1472, n1473, n1474, n1475, n1476, n1477;
  wire n1478, n1479, n1480, n1488, n1489, n1490, n1496, n1497;
  wire n1498, n1499, n1511, n1521, n1522, n1523, n1524, n1527;
  wire n1528, n1529, n1530, n1531, n1532, n1533, n1549, n1550;
  wire n1555, n1556, n1557, n1572, n1573, n1574, n1575, n1576;
  wire n1577, n1578, n1585, n1586, n1587, n1588, n1600, n1601;
  wire n1602, n1603, n1604, n1610, n1611, n1615, n1616, n1617;
  wire n1621, n1635, n1636, n1640, n1643, n1644, n1645, n1646;
  wire n1665, n1666, n1667, n1668, n1669, n1679, n1680, n1681;
  wire n1687, n1691, n1692, n1693, n1694, n1695, n1696, n1697;
  wire n1708, n1709, n1719, n1720, n1721, n1725, n1726, n1727;
  wire n1731, n1732, n1735, n1736, n1737, n1738, n1739, n1740;
  wire n1754, n1755, n1759, n1760, n1761, n1762, n1763, n1779;
  wire n1780, n1781, n1782, n1783, n1784, n1785, n1794, n1795;
  wire n1798, n1799, n1800, n1814, n1819, n1823, n1824, n1825;
  wire n1826, n1827, n1828, n1838, n1839, n1844, n1857, n1858;
  wire n1859, n1860, n1861, n1877, n1878, n1879, n1884, n1887;
  wire n1890, n1893, n1894, n1895, n1896, n1897, n1898, n1913;
  wire n1914, n1915, n1916, n1917, n1925, n1928, n1931, n1940;
  wire n1941, n1942, n1943, n1944, n1958, n1959, n1960, n1969;
  wire n1970, n1971, n1972, n1973, n1992, n1993, n1994, n1995;
  wire n1996, n2006, n2007, n2010, n2011, n2012, n2013, n2014;
  wire n2017, n2020, n2021, n2022, n2025, n2026, n2040, n2057;
  wire n2058, n2059, n2068, n2072, n2073, n2074, n2075, n2088;
  wire n2089, n2090, n2091, n2092, n2093, n2104, n2105, n2112;
  wire n2113, n2114, n2115, n2127, n2132, n2133, n2152, n2153;
  wire n2154, n2167, n2168, n2169, n2170, n2171, n2172, n2173;
  wire n2174, n2175, n2176, n2189, n2190, n2191, n2192, n2202;
  wire n2208, n2209, n2210, n2217, n2218, n2219, n2220, n2229;
  wire n2230, n2237, n2240, n2241, n2258, n2262, n2263, n2264;
  wire n2265, n2266, n2267, n2273, n2274, n2275, n2276, n2277;
  wire n2278, n2291, n2292, n2293, n2296, n2297, n2301, n2302;
  wire n2303, n2317, n2325, n2330, n2331, n2332, n2333, n2334;
  wire n2345, n2346, n2347, n2348, n2349, n2360, n2361, n2362;
  wire n2363, n2370, n2371, n2388, n2389, n2390, n2405, n2406;
  wire n2409, n2410, n2417, n2422, n2423, n2424, n2425, n2426;
  wire n2427, n2439, n2440, n2441, n2442, n2443, n2444, n2445;
  wire n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2483;
  wire n2484, n2487, n2500, n2506, n2507, n2508, n2512, n2515;
  wire n2533, n2534, n2537, n2543, n2544, n2545, n2546, n2555;
  wire n2556, n2571, n2572, n2573, n2581, n2582, n2583, n2584;
  wire n2591, n2592, n2593, n2594, n2595, n2605, n2606, n2607;
  wire n2608, n2623, n2624, n2625, n2626, n2627, n2632, n2633;
  wire n2634, n2635, n2636, n2637, n2650, n2651, n2652, n2653;
  wire n2656, n2674, n2675, n2678, n2682, n2683, n2684, n2697;
  wire n2698, n2703, n2704, n2705, n2716, n2719, n2720, n2721;
  wire n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2751;
  wire n2752, n2753, n2758, n2759, n2760, n2772, n2778, n2782;
  wire n2783, n2784, n2796, n2806, n2807, n2808, n2809, n2810;
  wire n2811, n2829, n2830, n2831, n2832, n2833, n2834, n2835;
  wire n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843;
  wire n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851;
  wire n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859;
  wire n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867;
  wire n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875;
  wire n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883;
  wire n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891;
  wire n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899;
  wire n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907;
  wire n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915;
  wire n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923;
  wire n2924, n2925, n2926, n2927, n2928, n2931, n2940, n2943;
  wire n2958, n2961, n2962, n2963, n2979, n2987, n2990, n2991;
  wire n2992, n2993, n2994, n2995, n3012, n3013, n3014, n3015;
  wire n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023;
  wire n3024, n3025, n3026, n3027, n3028, n3029, n3032, n3039;
  wire n3040, n3041, n3042, n3043, n3044, n3045, n3057, n3058;
  wire n3059, n3065, n3068, n3083, n3084, n3085, n3094, n3108;
  wire n3113, n3114, n3115, n3127, n3128, n3146, n3147, n3148;
  wire n3155, n3159, n3160, n3161, n3162, n3163, n3164, n3165;
  wire n3180, n3191, n3192, n3193, n3194, n3205, n3206, n3219;
  wire n3225, n3226, n3239, n3240, n3241, n3242, n3243, n3244;
  wire n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252;
  wire n3259, n3260, n3261, n3264, n3265, n3266, n3267, n3268;
  wire n3282, n3290, n3296, n3297, n3298, n3299, n3300, n3312;
  wire n3313, n3314, n3327, n3328, n3329, n3330, n3331, n3332;
  wire n3333, n3334, n3335, n3338, n3339, n3340, n3341, n3342;
  wire n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350;
  wire n3351, n3354, n3355, n3356, n3357, n3358, n3359, n3360;
  wire n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368;
  wire n3369, n3370, n3378, n3379, n3380, n3386, n3389, n3390;
  wire n3391, n3392, n3393, n3405, n3408, n3409, n3415, n3416;
  wire n3432, n3435, n3436, n3437, n3438, n3456, n3457, n3458;
  wire n3459, n3464, n3470, n3471, n3472, n3473, n3474, n3489;
  wire n3490, n3497, n3510, n3511, n3512, n3513, n3514, n3521;
  wire n3522, n3523, n3524, n3539, n3540, n3541, n3542, n3543;
  wire n3544, n3548, n3549, n3559, n3565, n3569, n3570, n3580;
  wire n3581, n3582, n3583, n3587, n3605, n3606, n3607, n3608;
  wire n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616;
  wire n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624;
  wire n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632;
  wire n3633, n3634, n3635, n3636, n3644, n3645, n3651, n3663;
  wire n3675, n3681, n3685, n3686, n3687, n3702, n3703, n3704;
  wire n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712;
  wire n3713, n3714, n3715, n3716, n3719, n3720, n3721, n3722;
  wire n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3733;
  wire n3739, n3743, n3757, n3764, n3768, n3771, n3782, n3790;
  wire n3791, n3792, n3805, n3806, n3807, n3808, n3809, n3810;
  wire n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818;
  wire n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826;
  wire n3827, n3831, n3832, n3839, n3848, n3852, n3856, n3857;
  wire n3858, n3866, n3869, n3873, n3874, n3877, n3878, n3879;
  wire n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3901;
  wire n3905, n3906, n3912, n3913, n3914, n3929, n3930, n3931;
  wire n3939, n3947, n3948, n3949, n3964, n3965, n3966, n3967;
  wire n3968, n3972, n3978, n3984, n3985, n3986, n3987, n3990;
  wire n3997, n4003, n4009, n4010, n4011, n4017, n4030, n4034;
  wire n4040, n4045, n4046, n4047, n4050, n4051, n4052, n4053;
  wire n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061;
  wire n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069;
  wire n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077;
  wire n4078, n4079, n4080, n4083, n4084, n4085, n4086, n4087;
  wire n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095;
  wire n4096, n4097, n4098, n4099, n4100, n4101, n4104, n4121;
  wire n4127, n4130, n4131, n4132, n4148, n4151, n4152, n4153;
  wire n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178;
  wire n4179, n4180, n4181, n4182, n4183, n4186, n4187, n4188;
  wire n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196;
  wire n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204;
  wire n4205, n4208, n4209, n4215, n4216, n4217, n4218, n4232;
  wire n4233, n4234, n4247, n4266, n4267, n4268, n4269, n4274;
  wire n4279, n4293, n4294, n4295, n4298, n4311, n4312, n4313;
  wire n4325, n4326, n4327, n4332, n4333, n4334, n4335, n4351;
  wire n4356, n4357, n4366, n4367, n4375, n4388, n4405, n4421;
  wire n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429;
  wire n4430, n4431, n4432, n4433, n4436, n4437, n4438, n4439;
  wire n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447;
  wire n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455;
  wire n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463;
  wire n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471;
  wire n4472, n4473, n4476, n4477, n4478, n4479, n4480, n4481;
  wire n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4493;
  wire n4502, n4511, n4514, n4515, n4516, n4517, n4518, n4519;
  wire n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527;
  wire n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535;
  wire n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543;
  wire n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551;
  wire n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559;
  wire n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567;
  wire n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577;
  wire n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585;
  wire n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593;
  wire n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601;
  wire n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609;
  wire n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617;
  wire n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625;
  wire n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633;
  wire n4634, n4637, n4638, n4639, n4640, n4641, n4644, n4645;
  wire n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653;
  wire n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4663;
  wire n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671;
  wire n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679;
  wire n4680, n4683, n4684, n4685, n4686, n4687, n4688, n4689;
  wire n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697;
  wire n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707;
  wire n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715;
  wire n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723;
  wire n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731;
  wire n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739;
  wire n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747;
  wire n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755;
  wire n4756, n4757, n4758, n4759, n4760, n4761, n4767, n4768;
  wire n4769, n4770, n4771, n4785, n4786, n4787, n4788, n4794;
  wire n4797, n4798, n4799, n4815, n4819, n4827, n4828, n4844;
  wire n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852;
  wire n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862;
  wire n4863, n4864, n4865, n4868, n4869, n4870, n4871, n4872;
  wire n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880;
  wire n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888;
  wire n4889, n4890, n4891, n4892, n4893, n4894, n4897, n4898;
  wire n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906;
  wire n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914;
  wire n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924;
  wire n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932;
  wire n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940;
  wire n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948;
  wire n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956;
  wire n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4966;
  wire n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974;
  wire n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982;
  wire n4983, n4986, n4987, n4988, n4989, n4990, n4991, n4992;
  wire n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000;
  wire n5001, n5002, n5013, n5019, n5020, n5021, n5034, n5035;
  wire n5036, n5037, n5038, n5039, n5040, n5053, n5056, n5063;
  wire n5064, n5065, n5066, n5082, n5085, n5106, n5107, n5108;
  wire n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116;
  wire n5117, n5118, n5121, n5122, n5123, n5124, n5125, n5126;
  wire n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134;
  wire n5135, n5136, n5137, n5138, n5139, n5140, n5143, n5144;
  wire n5148, n5149, n5150, n5151, n5152, n5168, n5169, n5170;
  wire n5171, n5172, n5173, n5188, n5189, n5190, n5193, n5199;
  wire n5200, n5201, n5209, n5224, n5233, n5239, n5254, n5264;
  wire n5269, n5270, n5271, n5286, n5296, n5304, n5320, n5321;
  wire n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329;
  wire n5330, n5331, n5332, n5335, n5336, n5337, n5338, n5339;
  wire n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347;
  wire n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355;
  wire n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363;
  wire n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371;
  wire n5372, n5373, n5374, n5377, n5378, n5379, n5380, n5381;
  wire n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389;
  wire n5390, n5393, n5394, n5395, n5396, n5397, n5398, n5399;
  wire n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407;
  wire n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415;
  wire n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423;
  wire n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431;
  wire n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439;
  wire n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5449;
  wire n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457;
  wire n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465;
  wire n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473;
  wire n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481;
  wire n5482, n5485, n5486, n5487, n5488, n5489, n5490, n5491;
  wire n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499;
  wire n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509;
  wire n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517;
  wire n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525;
  wire n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533;
  wire n5534, n5535, n5536, n5539, n5540, n5541, n5542, n5543;
  wire n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551;
  wire n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559;
  wire n5560, n5561, n5562, n5565, n5566, n5567, n5568, n5569;
  wire n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579;
  wire n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587;
  wire n5588, n5591, n5592, n5593, n5594, n5595, n5596, n5597;
  wire n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605;
  wire n5606, n5607, n5608, n5611, n5612, n5613, n5614, n5615;
  wire n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623;
  wire n5624, n5627, n5628, n5629, n5630, n5631, n5632, n5633;
  wire n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641;
  wire n5642, n5645, n5646, n5647, n5648, n5649, n5650, n5651;
  wire n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659;
  wire n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667;
  wire n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675;
  wire n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683;
  wire n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691;
  wire n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699;
  wire n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707;
  wire n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715;
  wire n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723;
  wire n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731;
  wire n5732, n5733, n5734, n5746, n5747, n5748, n5765, n5766;
  wire n5767, n5773, n5774, n5775, n5776, n5777, n5785, n5786;
  wire n5787, n5791, n5792, n5793, n5806, n5807, n5808, n5825;
  wire n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833;
  wire n5834, n5835, n5836, n5837, n5838, n5841, n5842, n5843;
  wire n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851;
  wire n5852, n5853, n5854, n5855, n5858, n5859, n5860, n5861;
  wire n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869;
  wire n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877;
  wire n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5887;
  wire n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895;
  wire n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903;
  wire n5904, n5907, n5908, n5909, n5910, n5911, n5912, n5913;
  wire n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5923;
  wire n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931;
  wire n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939;
  wire n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947;
  wire n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955;
  wire n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963;
  wire n5964, n5967, n5968, n5969, n5970, n5971, n5972, n5973;
  wire n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981;
  wire n5982, n5983, n5984, n5987, n5988, n5989, n5990, n5991;
  wire n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999;
  wire n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007;
  wire n6008, n6011, n6012, n6013, n6014, n6015, n6020, n6026;
  wire n6041, n6042, n6043, n6054, n6055, n6056, n6074, n6075;
  wire n6076, n6083, n6084, n6097, n6102, n6103, n6104, n6118;
  wire n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126;
  wire n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136;
  wire n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144;
  wire n6145, n6146, n6147, n6150, n6151, n6152, n6153, n6154;
  wire n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162;
  wire n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170;
  wire n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178;
  wire n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6188;
  wire n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196;
  wire n6197, n6198, n6199, n6200, n6201, n6204, n6205, n6206;
  wire n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214;
  wire n6215, n6216, n6217, n6218, n6219, n6222, n6223, n6224;
  wire n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232;
  wire n6233, n6234, n6235, n6236, n6239, n6240, n6241, n6242;
  wire n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250;
  wire n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258;
  wire n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266;
  wire n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274;
  wire n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282;
  wire n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290;
  wire n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298;
  wire n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306;
  wire n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314;
  wire n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322;
  wire n6323, n6324, n6327, n6328, n6329, n6330, n6331, n6332;
  wire n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340;
  wire n6341, n6342, n6343, n6344, n6347, n6348, n6349, n6350;
  wire n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358;
  wire n6359, n6360, n6363, n6364, n6365, n6366, n6367, n6368;
  wire n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376;
  wire n6377, n6378, n6379, n6380, n6383, n6384, n6385, n6386;
  wire n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394;
  wire n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402;
  wire n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410;
  wire n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418;
  wire n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426;
  wire n6427, n6428, n6431, n6432, n6433, n6434, n6435, n6436;
  wire n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444;
  wire n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6454;
  wire n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462;
  wire n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470;
  wire n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478;
  wire n6479, n6480, n6483, n6484, n6485, n6486, n6487, n6488;
  wire n6489, n6490, n6491, n6492, n6493, n6496, n6497, n6498;
  wire n6499, n6500, n6514, n6517, n6520, n6536, n6537, n6538;
  wire n6539, n6540, n6541, n6542, n6545, n6546, n6547, n6548;
  wire n6561, n6565, n6566, n6567, n6586, n6587, n6588, n6589;
  wire n6590, n6591, n6592, n6595, n6596, n6604, n6607, n6610;
  wire n6625, n6628, n6641, n6642, n6643, n6644, n6645, n6646;
  wire n6647, n6650, n6651, n6662, n6663, n6664, n6667, n6670;
  wire n6671, n6672, n6690, n6691, n6692, n6693, n6694, n6695;
  wire n6696, n6699, n6700, n6705, n6706, n6707, n6714, n6715;
  wire n6716, n6717, n6732, n6733, n6734, n6748, n6755, n6769;
  wire n6770, n6771, n6791, n6792, n6793, n6794, n6795, n6796;
  wire n6797, n6798, n6799, n6802, n6803, n6804, n6805, n6806;
  wire n6807, n6808, n6809, n6810, n6813, n6814, n6815, n6816;
  wire n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824;
  wire n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832;
  wire n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840;
  wire n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848;
  wire n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856;
  wire n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864;
  wire n6865, n6866, n6867, n6868, n6869, n6872, n6873, n6874;
  wire n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882;
  wire n6883, n6884, n6885, n6886, n6887, n6890, n6891, n6892;
  wire n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900;
  wire n6901, n6902, n6903, n6906, n6907, n6908, n6909, n6910;
  wire n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918;
  wire n6919, n6920, n6921, n6924, n6925, n6926, n6927, n6928;
  wire n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936;
  wire n6937, n6940, n6941, n6942, n6943, n6944, n6945, n6946;
  wire n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954;
  wire n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962;
  wire n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970;
  wire n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978;
  wire n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986;
  wire n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994;
  wire n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002;
  wire n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010;
  wire n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018;
  wire n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026;
  wire n7027, n7028, n7029, n7030, n7031, n7034, n7035, n7036;
  wire n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044;
  wire n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7054;
  wire n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062;
  wire n7063, n7064, n7065, n7066, n7067, n7070, n7071, n7072;
  wire n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080;
  wire n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7090;
  wire n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098;
  wire n7099, n7100, n7101, n7102, n7103, n7104, n7107, n7108;
  wire n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116;
  wire n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124;
  wire n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132;
  wire n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140;
  wire n7141, n7142, n7145, n7146, n7147, n7148, n7149, n7150;
  wire n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158;
  wire n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7168;
  wire n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176;
  wire n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184;
  wire n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192;
  wire n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200;
  wire n7201, n7202, n7205, n7206, n7207, n7208, n7209, n7210;
  wire n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218;
  wire n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228;
  wire n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236;
  wire n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246;
  wire n7247, n7248, n7249, n7250, n7251, n7252, n7255, n7256;
  wire n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264;
  wire n7265, n7266, n7267, n7268, n7269, n7270, n7273, n7274;
  wire n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282;
  wire n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290;
  wire n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298;
  wire n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306;
  wire n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314;
  wire n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322;
  wire n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330;
  wire n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338;
  wire n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346;
  wire n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354;
  wire n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362;
  wire n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370;
  wire n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378;
  wire n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386;
  wire n7387, n7390, n7391, n7392, n7393, n7394, n7395, n7396;
  wire n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404;
  wire n7405, n7408, n7409, n7410, n7411, n7412, n7413, n7414;
  wire n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422;
  wire n7423, n7426, n7427, n7428, n7429, n7430, n7431, n7432;
  wire n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440;
  wire n7441, n7444, n7445, n7446, n7447, n7448, n7449, n7450;
  wire n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458;
  wire n7459, n7462, n7463, n7464, n7465, n7466, n7467, n7468;
  wire n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476;
  wire n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484;
  wire n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492;
  wire n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500;
  wire n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508;
  wire n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518;
  wire n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526;
  wire n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534;
  wire n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542;
  wire n7543, n7544, n7545, n7548, n7549, n7550, n7551, n7552;
  wire n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560;
  wire n7561, n7562, n7563, n7566, n7567, n7568, n7569, n7570;
  wire n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578;
  wire n7579, n7582, n7583, n7584, n7585, n7586, n7587, n7588;
  wire n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596;
  wire n7597, n7598, n7599, n7602, n7603, n7604, n7605, n7606;
  wire n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614;
  wire n7615, n7618, n7619, n7620, n7621, n7622, n7623, n7624;
  wire n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632;
  wire n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640;
  wire n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648;
  wire n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656;
  wire n7657, n7658, n7659, n7660, n7663, n7664, n7665, n7666;
  wire n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674;
  wire n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682;
  wire n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690;
  wire n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698;
  wire n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706;
  wire n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714;
  wire n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722;
  wire n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730;
  wire n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738;
  wire n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746;
  wire n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754;
  wire n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762;
  wire n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770;
  wire n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778;
  wire n7779, n7780, n7781, n7782, n7785, n7786, n7787, n7788;
  wire n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796;
  wire n7797, n7798, n7799, n7802, n7803, n7804, n7805, n7806;
  wire n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814;
  wire n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822;
  wire n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830;
  wire n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838;
  wire n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846;
  wire n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854;
  wire n7855, n7856, n7857, n7858, n7861, n7862, n7863, n7864;
  wire n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872;
  wire n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880;
  wire n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888;
  wire n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896;
  wire n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904;
  wire n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912;
  wire n7913, n7914, n7915, n7916, n7917, n7920, n7921, n7922;
  wire n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930;
  wire n7931, n7932, n7933, n7934, n7935, n7938, n7939, n7940;
  wire n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948;
  wire n7949, n7950, n7951, n7954, n7955, n7956, n7957, n7958;
  wire n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966;
  wire n7967, n7968, n7969, n7972, n7973, n7974, n7975, n7976;
  wire n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984;
  wire n7985, n7986, n7989, n7990, n7991, n7992, n7993, n7994;
  wire n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002;
  wire n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010;
  wire n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018;
  wire n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026;
  wire n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034;
  wire n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042;
  wire n8043, n8044, n8045, n8046, n8047, n8050, n8051, n8052;
  wire n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060;
  wire n8061, n8062, n8063, n8064, n8065, n8068, n8069, n8070;
  wire n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078;
  wire n8079, n8080, n8081, n8082, n8083, n8086, n8087, n8088;
  wire n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096;
  wire n8097, n8098, n8099, n8100, n8101, n8104, n8105, n8106;
  wire n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114;
  wire n8115, n8116, n8117, n8118, n8119, n8122, n8123, n8124;
  wire n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132;
  wire n8133, n8134, n8135, n8136, n8137, n8140, n8141, n8142;
  wire n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150;
  wire n8151, n8152, n8153, n8154, n8155, n8158, n8159, n8160;
  wire n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168;
  wire n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176;
  wire n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184;
  wire n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192;
  wire n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200;
  wire n8201, n8204, n8205, n8206, n8207, n8208, n8209, n8210;
  wire n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218;
  wire n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226;
  wire n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8236;
  wire n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244;
  wire n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252;
  wire n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260;
  wire n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268;
  wire n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276;
  wire n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284;
  wire n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292;
  wire n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302;
  wire n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310;
  wire n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318;
  wire n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326;
  wire n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334;
  wire n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342;
  wire n8343, n8346, n8347, n8348, n8349, n8350, n8351, n8352;
  wire n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360;
  wire n8361, n8364, n8365, n8366, n8367, n8368, n8369, n8370;
  wire n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8380;
  wire n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388;
  wire n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396;
  wire n8397, n8400, n8401, n8402, n8403, n8404, n8405, n8406;
  wire n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414;
  wire n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422;
  wire n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430;
  wire n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438;
  wire n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446;
  wire n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454;
  wire n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462;
  wire n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470;
  wire n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478;
  wire n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486;
  wire n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494;
  wire n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502;
  wire n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510;
  wire n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518;
  wire n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526;
  wire n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534;
  wire n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542;
  wire n8543, n8544, n8545, n8546, n8547, n8550, n8551, n8552;
  wire n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560;
  wire n8561, n8562, n8563, n8564, n8567, n8568, n8569, n8570;
  wire n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578;
  wire n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586;
  wire n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594;
  wire n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602;
  wire n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610;
  wire n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618;
  wire n8619, n8620, n8621, n8622, n8623, n8624, n8627, n8628;
  wire n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636;
  wire n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644;
  wire n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652;
  wire n8653, n8654, n8655, n8656, n8659, n8660, n8661, n8662;
  wire n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670;
  wire n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678;
  wire n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686;
  wire n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694;
  wire n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702;
  wire n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710;
  wire n8711, n8712, n8713, n8714, n8715, n8718, n8719, n8720;
  wire n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728;
  wire n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736;
  wire n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744;
  wire n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752;
  wire n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760;
  wire n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768;
  wire n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776;
  wire n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784;
  wire n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792;
  wire n8793, n8794, n8795, n8796, n8799, n8800, n8801, n8802;
  wire n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810;
  wire n8811, n8812, n8813, n8814, n8817, n8818, n8819, n8820;
  wire n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828;
  wire n8829, n8830, n8833, n8834, n8835, n8836, n8837, n8838;
  wire n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846;
  wire n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854;
  wire n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862;
  wire n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870;
  wire n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878;
  wire n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886;
  wire n8887, n8888, n8891, n8892, n8893, n8894, n8895, n8896;
  wire n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904;
  wire n8905, n8906, n8909, n8910, n8911, n8912, n8913, n8914;
  wire n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922;
  wire n8923, n8924, n8927, n8928, n8929, n8930, n8931, n8932;
  wire n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940;
  wire n8941, n8942, n8945, n8946, n8947, n8948, n8949, n8950;
  wire n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958;
  wire n8959, n8960, n8963, n8964, n8965, n8966, n8967, n8968;
  wire n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976;
  wire n8977, n8978, n8981, n8982, n8983, n8984, n8985, n8986;
  wire n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994;
  wire n8995, n8996, n8999, n9000, n9001, n9002, n9003, n9004;
  wire n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012;
  wire n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020;
  wire n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028;
  wire n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036;
  wire n9037, n9038, n9039, n9040, n9041, n9042, n9045, n9046;
  wire n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054;
  wire n9055, n9056, n9057, n9058, n9059, n9062, n9063, n9064;
  wire n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072;
  wire n9073, n9074, n9075, n9076, n9077, n9080, n9081, n9082;
  wire n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090;
  wire n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098;
  wire n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106;
  wire n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114;
  wire n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122;
  wire n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130;
  wire n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9140;
  wire n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148;
  wire n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156;
  wire n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164;
  wire n9165, n9166, n9167, n9168, n9169, n9172, n9173, n9174;
  wire n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182;
  wire n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190;
  wire n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198;
  wire n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206;
  wire n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214;
  wire n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222;
  wire n9223, n9224, n9225, n9226, n9227, n9228, n9231, n9232;
  wire n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240;
  wire n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248;
  wire n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256;
  wire n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264;
  wire n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272;
  wire n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280;
  wire n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288;
  wire n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296;
  wire n9297, n9298, n9299, n9302, n9303, n9304, n9305, n9306;
  wire n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314;
  wire n9315, n9316, n9317, n9320, n9321, n9322, n9323, n9324;
  wire n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332;
  wire n9333, n9334, n9337, n9338, n9339, n9340, n9341, n9342;
  wire n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350;
  wire n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358;
  wire n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366;
  wire n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374;
  wire n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382;
  wire n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390;
  wire n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398;
  wire n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406;
  wire n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414;
  wire n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422;
  wire n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430;
  wire n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438;
  wire n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446;
  wire n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454;
  wire n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462;
  wire n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470;
  wire n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480;
  wire n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9490;
  wire n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498;
  wire n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506;
  wire n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514;
  wire n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522;
  wire n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530;
  wire n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538;
  wire n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546;
  wire n9547, n9550, n9551, n9552, n9553, n9554, n9555, n9556;
  wire n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564;
  wire n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574;
  wire n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582;
  wire n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592;
  wire n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600;
  wire n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608;
  wire n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616;
  wire n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624;
  wire n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632;
  wire n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640;
  wire n9641, n9642, n9645, n9646, n9647, n9648, n9649, n9650;
  wire n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658;
  wire n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666;
  wire n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674;
  wire n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684;
  wire n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692;
  wire n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700;
  wire n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708;
  wire n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716;
  wire n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724;
  wire n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732;
  wire n9733, n9736, n9737, n9738, n9739, n9740, n9741, n9742;
  wire n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750;
  wire n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758;
  wire n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766;
  wire n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774;
  wire n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782;
  wire n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790;
  wire n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798;
  wire n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806;
  wire n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814;
  wire n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822;
  wire n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830;
  wire n9831, n9832, n9833, n9834, n9837, n9838, n9839, n9840;
  wire n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848;
  wire n9849, n9850, n9851, n9852, n9855, n9856, n9857, n9858;
  wire n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866;
  wire n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874;
  wire n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882;
  wire n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890;
  wire n9891, n9892, n9893, n9896, n9897, n9898, n9899, n9900;
  wire n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908;
  wire n9909, n9910, n9911, n9914, n9915, n9916, n9917, n9918;
  wire n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926;
  wire n9927, n9928, n9929, n9932, n9933, n9934, n9935, n9936;
  wire n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944;
  wire n9945, n9946, n9947, n9950, n9951, n9952, n9953, n9954;
  wire n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962;
  wire n9963, n9964, n9965, n9968, n9969, n9970, n9971, n9972;
  wire n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980;
  wire n9981, n9982, n9983, n9986, n9987, n9988, n9989, n9990;
  wire n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998;
  wire n9999, n10000, n10001, n10004, n10005, n10006, n10007, n10008;
  wire n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016;
  wire n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024;
  wire n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032;
  wire n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040;
  wire n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10050;
  wire n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058;
  wire n10059, n10060, n10061, n10062, n10063, n10064, n10067, n10068;
  wire n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076;
  wire n10077, n10078, n10079, n10080, n10081, n10082, n10085, n10086;
  wire n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094;
  wire n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102;
  wire n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110;
  wire n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118;
  wire n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126;
  wire n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134;
  wire n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142;
  wire n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152;
  wire n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10162;
  wire n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170;
  wire n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10180;
  wire n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188;
  wire n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196;
  wire n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204;
  wire n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212;
  wire n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220;
  wire n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228;
  wire n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236;
  wire n10237, n10240, n10241, n10242, n10243, n10244, n10245, n10246;
  wire n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254;
  wire n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262;
  wire n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10272;
  wire n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280;
  wire n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288;
  wire n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296;
  wire n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304;
  wire n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312;
  wire n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320;
  wire n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328;
  wire n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338;
  wire n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346;
  wire n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354;
  wire n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362;
  wire n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370;
  wire n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378;
  wire n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386;
  wire n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394;
  wire n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402;
  wire n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410;
  wire n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418;
  wire n10419, n10422, n10423, n10424, n10425, n10426, n10427, n10428;
  wire n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436;
  wire n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444;
  wire n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452;
  wire n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460;
  wire n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468;
  wire n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476;
  wire n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484;
  wire n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492;
  wire n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500;
  wire n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508;
  wire n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516;
  wire n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524;
  wire n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532;
  wire n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540;
  wire n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548;
  wire n10549, n10550, n10551, n10552, n10553, n10554, n10557, n10558;
  wire n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566;
  wire n10567, n10568, n10569, n10570, n10571, n10574, n10575, n10576;
  wire n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584;
  wire n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592;
  wire n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600;
  wire n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608;
  wire n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616;
  wire n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624;
  wire n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10634;
  wire n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642;
  wire n10643, n10644, n10645, n10646, n10647, n10648, n10651, n10652;
  wire n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660;
  wire n10661, n10662, n10663, n10664, n10665, n10666, n10669, n10670;
  wire n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678;
  wire n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686;
  wire n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694;
  wire n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702;
  wire n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710;
  wire n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718;
  wire n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726;
  wire n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736;
  wire n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10746;
  wire n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754;
  wire n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10764;
  wire n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772;
  wire n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780;
  wire n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788;
  wire n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796;
  wire n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804;
  wire n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812;
  wire n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820;
  wire n10821, n10824, n10825, n10826, n10827, n10828, n10829, n10830;
  wire n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838;
  wire n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846;
  wire n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10856;
  wire n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864;
  wire n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872;
  wire n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880;
  wire n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888;
  wire n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896;
  wire n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904;
  wire n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912;
  wire n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922;
  wire n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930;
  wire n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938;
  wire n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946;
  wire n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954;
  wire n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962;
  wire n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970;
  wire n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978;
  wire n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986;
  wire n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994;
  wire n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002;
  wire n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010;
  wire n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018;
  wire n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026;
  wire n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034;
  wire n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044;
  wire n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052;
  wire n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060;
  wire n11061, n11062, n11063, n11064, n11065, n11066, n11069, n11070;
  wire n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078;
  wire n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086;
  wire n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11096;
  wire n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104;
  wire n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11114;
  wire n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122;
  wire n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11132;
  wire n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140;
  wire n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11150;
  wire n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158;
  wire n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11168;
  wire n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176;
  wire n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11186;
  wire n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194;
  wire n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202;
  wire n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210;
  wire n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218;
  wire n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226;
  wire n11227, n11228, n11229, n11232, n11233, n11234, n11235, n11236;
  wire n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244;
  wire n11245, n11246, n11249, n11250, n11251, n11252, n11253, n11254;
  wire n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262;
  wire n11263, n11264, n11267, n11268, n11269, n11270, n11271, n11272;
  wire n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280;
  wire n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288;
  wire n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296;
  wire n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304;
  wire n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312;
  wire n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320;
  wire n11321, n11322, n11323, n11324, n11327, n11328, n11329, n11330;
  wire n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338;
  wire n11339, n11340, n11341, n11344, n11345, n11346, n11347, n11348;
  wire n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356;
  wire n11357, n11358, n11359, n11362, n11363, n11364, n11365, n11366;
  wire n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374;
  wire n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382;
  wire n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390;
  wire n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398;
  wire n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406;
  wire n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414;
  wire n11415, n11416, n11417, n11418, n11419, n11422, n11423, n11424;
  wire n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432;
  wire n11433, n11434, n11435, n11436, n11439, n11440, n11441, n11442;
  wire n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450;
  wire n11451, n11452, n11453, n11454, n11457, n11458, n11459, n11460;
  wire n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468;
  wire n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476;
  wire n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484;
  wire n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492;
  wire n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500;
  wire n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508;
  wire n11509, n11510, n11511, n11512, n11513, n11514, n11517, n11518;
  wire n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526;
  wire n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534;
  wire n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542;
  wire n11543, n11544, n11545, n11546, n11549, n11550, n11551, n11552;
  wire n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560;
  wire n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568;
  wire n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576;
  wire n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584;
  wire n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592;
  wire n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600;
  wire n11601, n11602, n11603, n11604, n11605, n11608, n11609, n11610;
  wire n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618;
  wire n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626;
  wire n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634;
  wire n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642;
  wire n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650;
  wire n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658;
  wire n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666;
  wire n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674;
  wire n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682;
  wire n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690;
  wire n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698;
  wire n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706;
  wire n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714;
  wire n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722;
  wire n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730;
  wire n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738;
  wire n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746;
  wire n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754;
  wire n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762;
  wire n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770;
  wire n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778;
  wire n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786;
  wire n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794;
  wire n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802;
  wire n11803, n11804, n11805, n11806, n11807, n11808, n11814, n11815;
  wire n11816, n11817, n11818, n11819, n11822, n11823, n11824, n11825;
  wire n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833;
  wire n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841;
  wire n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849;
  wire n11850, n11853, n11854, n11855, n11856, n11857, n11858, n11859;
  wire n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867;
  wire n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875;
  wire n11876, n11877, n11878, n11879, n11880, n11881, n11884, n11885;
  wire n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893;
  wire n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901;
  wire n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909;
  wire n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917;
  wire n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925;
  wire n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933;
  wire n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941;
  wire n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949;
  wire n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959;
  wire n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11969;
  wire n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977;
  wire n11978, n11979, n11980, n11983, n11984, n11985, n11986, n11987;
  wire n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995;
  wire n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003;
  wire n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011;
  wire n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019;
  wire n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027;
  wire n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035;
  wire n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043;
  wire n12044, n12045, n12046, n12047, n12048, n12051, n12052, n12053;
  wire n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061;
  wire n12062, n12063, n12064, n12065, n12068, n12069, n12070, n12071;
  wire n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079;
  wire n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089;
  wire n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097;
  wire n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105;
  wire n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113;
  wire n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121;
  wire n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129;
  wire n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137;
  wire n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145;
  wire n12146, n12147, n12150, n12151, n12152, n12153, n12154, n12155;
  wire n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163;
  wire n12164, n12167, n12168, n12169, n12170, n12171, n12172, n12173;
  wire n12174, n12175, n12176, n12177, n12178, n12181, n12182, n12183;
  wire n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191;
  wire n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199;
  wire n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207;
  wire n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215;
  wire n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223;
  wire n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231;
  wire n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239;
  wire n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12249;
  wire n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257;
  wire n12258, n12259, n12260, n12263, n12264, n12265, n12266, n12267;
  wire n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275;
  wire n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283;
  wire n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291;
  wire n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299;
  wire n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307;
  wire n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315;
  wire n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323;
  wire n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331;
  wire n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339;
  wire n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347;
  wire n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355;
  wire n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363;
  wire n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371;
  wire n12372, n12373, n12374, n12375, n12378, n12379, n12380, n12381;
  wire n12382, n12383, n12384, n12387, n12390, n12396, n12397, n12404;
  wire n12409, n12412, n12428, n12431, n12448, n12449, n12450, n12451;
  wire n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459;
  wire n12460, n12463, n12464, n12465, n12466, n12467, n12468, n12469;
  wire n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477;
  wire n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485;
  wire n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493;
  wire n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501;
  wire n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509;
  wire n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517;
  wire n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525;
  wire n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533;
  wire n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541;
  wire n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549;
  wire n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557;
  wire n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565;
  wire n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573;
  wire n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581;
  wire n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589;
  wire n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597;
  wire n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605;
  wire n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613;
  wire n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621;
  wire n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629;
  wire n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637;
  wire n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645;
  wire n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653;
  wire n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661;
  wire n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669;
  wire n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677;
  wire n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685;
  wire n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693;
  wire n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12703;
  wire n12710, n12711, n12712, n12730, n12731, n12732, n12733, n12734;
  wire n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742;
  wire n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750;
  wire n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758;
  wire n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766;
  wire n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774;
  wire n12775, n12776, n12777, n12778, n12779, n12780, n12783, n12784;
  wire n12785, n12795, n12805, n12810, n12811, n12812, n12828, n12829;
  wire n12830, n12842, n12843, n12844, n12845, n12846, n12847, n12848;
  wire n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856;
  wire n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864;
  wire n12865, n12866, n12867, n12868, n12871, n12872, n12873, n12874;
  wire n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882;
  wire n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890;
  wire n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898;
  wire n12899, n12902, n12909, n12910, n12911, n12919, n12924, n12932;
  wire n12939, n12940, n12941, n12944, n12958, n12973, n12977, n12995;
  wire n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003;
  wire n13006, n13007, n13008, n13009, n13012, n13013, n13014, n13015;
  wire n13016, n13031, n13041, n13056, n13059, n13063, n13074, n13075;
  wire n13081, n13082, n13083, n13087, n13095, n13096, n13097, n13098;
  wire n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106;
  wire n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114;
  wire n13123, n13135, n13138, n13158, n13161, n13172, n13173, n13174;
  wire n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182;
  wire n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190;
  wire n13191, n13192, n13193, n13194, n13195, n13196, n13210, n13221;
  wire n13238, n13239, n13240, n13247, n13248, n13249, n13265, n13268;
  wire n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290;
  wire n13291, n13292, n13293, n13296, n13297, n13298, n13299, n13300;
  wire n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308;
  wire n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318;
  wire n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326;
  wire n13327, n13328, n13329, n13332, n13333, n13334, n13335, n13336;
  wire n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344;
  wire n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352;
  wire n13353, n13354, n13355, n13358, n13359, n13360, n13361, n13362;
  wire n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370;
  wire n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378;
  wire n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386;
  wire n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394;
  wire n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404;
  wire n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412;
  wire n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420;
  wire n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428;
  wire n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436;
  wire n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444;
  wire n13445, n13458, n13474, n13475, n13476, n13477, n13478, n13479;
  wire n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487;
  wire n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495;
  wire n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503;
  wire n13504, n13507, n13508, n13509, n13510, n13511, n13512, n13513;
  wire n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521;
  wire n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529;
  wire n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537;
  wire n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545;
  wire n13546, n13547, n13548, n13549, n13560, n13574, n13575, n13576;
  wire n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584;
  wire n13585, n13586, n13587, n13588, n13591, n13592, n13593, n13594;
  wire n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602;
  wire n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610;
  wire n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618;
  wire n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626;
  wire n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634;
  wire n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644;
  wire n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652;
  wire n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660;
  wire n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668;
  wire n13669, n13670, n13671, n13677, n13695, n13698, n13699, n13700;
  wire n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722;
  wire n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730;
  wire n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13740;
  wire n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748;
  wire n13749, n13750, n13751, n13752, n13755, n13756, n13757, n13758;
  wire n13768, n13773, n13774, n13787, n13788, n13789, n13805, n13806;
  wire n13807, n13808, n13821, n13826, n13827, n13843, n13844, n13845;
  wire n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853;
  wire n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861;
  wire n13862, n13863, n13864, n13867, n13868, n13869, n13870, n13871;
  wire n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879;
  wire n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887;
  wire n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895;
  wire n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903;
  wire n13904, n13907, n13908, n13909, n13910, n13911, n13912, n13913;
  wire n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921;
  wire n13922, n13923, n13924, n13925, n13928, n13929, n13930, n13931;
  wire n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939;
  wire n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947;
  wire n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955;
  wire n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963;
  wire n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971;
  wire n13972, n13975, n13976, n13977, n13978, n13979, n13980, n13981;
  wire n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989;
  wire n13990, n13991, n13994, n13995, n13996, n13997, n13998, n13999;
  wire n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14009;
  wire n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017;
  wire n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14027;
  wire n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035;
  wire n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043;
  wire n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051;
  wire n14052, n14053, n14054, n14055, n14058, n14059, n14060, n14061;
  wire n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069;
  wire n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077;
  wire n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085;
  wire n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095;
  wire n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103;
  wire n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113;
  wire n14114, n14115, n14116, n14117, n14118, n14119, n14122, n14123;
  wire n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131;
  wire n14132, n14135, n14136, n14137, n14138, n14139, n14140, n14141;
  wire n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149;
  wire n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157;
  wire n14158, n14159, n14160, n14161, n14162, n14163, n14166, n14167;
  wire n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175;
  wire n14176, n14177, n14178, n14179, n14180, n14181, n14184, n14189;
  wire n14202, n14210, n14228, n14229, n14230, n14231, n14232, n14233;
  wire n14234, n14235, n14236, n14237, n14240, n14241, n14242, n14243;
  wire n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251;
  wire n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259;
  wire n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267;
  wire n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275;
  wire n14276, n14279, n14280, n14281, n14282, n14283, n14284, n14285;
  wire n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293;
  wire n14294, n14297, n14298, n14299, n14300, n14301, n14302, n14303;
  wire n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311;
  wire n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319;
  wire n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327;
  wire n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335;
  wire n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345;
  wire n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353;
  wire n14354, n14355, n14356, n14359, n14360, n14361, n14362, n14363;
  wire n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371;
  wire n14381, n14386, n14403, n14407, n14422, n14423, n14424, n14425;
  wire n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433;
  wire n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441;
  wire n14442, n14443, n14444, n14447, n14448, n14449, n14450, n14451;
  wire n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14461;
  wire n14462, n14463, n14464, n14465, n14466, n14467, n14476, n14479;
  wire n14482, n14498, n14514, n14515, n14516, n14517, n14518, n14525;
  wire n14534, n14544, n14559, n14560, n14561, n14565, n14572, n14588;
  wire n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596;
  wire n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604;
  wire n14605, n14606, n14607, n14608, n14609, n14612, n14613, n14614;
  wire n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622;
  wire n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630;
  wire n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638;
  wire n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646;
  wire n14647, n14648, n14649, n14652, n14653, n14654, n14655, n14656;
  wire n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664;
  wire n14665, n14668, n14669, n14670, n14671, n14672, n14673, n14674;
  wire n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682;
  wire n14683, n14686, n14687, n14688, n14689, n14690, n14691, n14692;
  wire n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700;
  wire n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708;
  wire n14709, n14710, n14713, n14714, n14715, n14716, n14717, n14718;
  wire n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726;
  wire n14727, n14730, n14731, n14732, n14733, n14734, n14735, n14736;
  wire n14737, n14738, n14739, n14740, n14741, n14742, n14745, n14746;
  wire n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754;
  wire n14755, n14756, n14757, n14758, n14759, n14760, n14763, n14764;
  wire n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772;
  wire n14773, n14774, n14775, n14776, n14779, n14780, n14781, n14782;
  wire n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14792;
  wire n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800;
  wire n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808;
  wire n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816;
  wire n14817, n14820, n14821, n14822, n14823, n14824, n14825, n14826;
  wire n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834;
  wire n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14844;
  wire n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852;
  wire n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860;
  wire n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868;
  wire n14869, n14870, n14871, n14874, n14875, n14876, n14877, n14878;
  wire n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886;
  wire n14887, n14888, n14889, n14892, n14893, n14894, n14895, n14896;
  wire n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904;
  wire n14905, n14908, n14909, n14910, n14911, n14912, n14913, n14914;
  wire n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922;
  wire n14923, n14926, n14927, n14928, n14929, n14930, n14931, n14932;
  wire n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940;
  wire n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948;
  wire n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956;
  wire n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964;
  wire n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974;
  wire n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982;
  wire n14983, n14984, n14985, n14986, n14987, n14988, n14991, n14992;
  wire n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000;
  wire n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15010;
  wire n15011, n15012, n15028, n15029, n15030, n15031, n15032, n15033;
  wire n15034, n15035, n15047, n15050, n15061, n15074, n15075, n15076;
  wire n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084;
  wire n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092;
  wire n15093, n15094, n15095, n15096, n15097, n15100, n15101, n15102;
  wire n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110;
  wire n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118;
  wire n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126;
  wire n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134;
  wire n15135, n15136, n15137, n15138, n15141, n15142, n15143, n15144;
  wire n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152;
  wire n15153, n15154, n15155, n15156, n15159, n15160, n15161, n15162;
  wire n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170;
  wire n15171, n15172, n15175, n15176, n15177, n15178, n15179, n15180;
  wire n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188;
  wire n15189, n15190, n15193, n15194, n15195, n15196, n15197, n15198;
  wire n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206;
  wire n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214;
  wire n15215, n15216, n15217, n15220, n15221, n15222, n15223, n15224;
  wire n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232;
  wire n15233, n15234, n15235, n15236, n15237, n15238, n15241, n15242;
  wire n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250;
  wire n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258;
  wire n15259, n15262, n15263, n15264, n15265, n15266, n15283, n15284;
  wire n15285, n15286, n15305, n15306, n15312, n15324, n15330, n15337;
  wire n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359;
  wire n15360, n15363, n15364, n15365, n15366, n15367, n15368, n15369;
  wire n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377;
  wire n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385;
  wire n15386, n15387, n15388, n15389, n15392, n15393, n15394, n15395;
  wire n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403;
  wire n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411;
  wire n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419;
  wire n15420, n15421, n15422, n15423, n15424, n15425, n15428, n15429;
  wire n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437;
  wire n15438, n15439, n15440, n15441, n15444, n15445, n15446, n15447;
  wire n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455;
  wire n15456, n15457, n15458, n15459, n15462, n15463, n15464, n15465;
  wire n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473;
  wire n15474, n15475, n15478, n15479, n15480, n15481, n15482, n15483;
  wire n15484, n15485, n15486, n15487, n15488, n15491, n15492, n15493;
  wire n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501;
  wire n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509;
  wire n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15519;
  wire n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527;
  wire n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535;
  wire n15536, n15537, n15538, n15539, n15542, n15543, n15544, n15545;
  wire n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553;
  wire n15554, n15555, n15556, n15559, n15560, n15561, n15562, n15563;
  wire n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571;
  wire n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581;
  wire n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589;
  wire n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599;
  wire n15600, n15601, n15602, n15603, n15604, n15605, n15608, n15609;
  wire n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617;
  wire n15618, n15619, n15620, n15621, n15622, n15623, n15626, n15627;
  wire n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635;
  wire n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643;
  wire n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651;
  wire n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659;
  wire n15660, n15661, n15662, n15663, n15664, n15667, n15668, n15669;
  wire n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677;
  wire n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685;
  wire n15686, n15687, n15690, n15691, n15692, n15693, n15694, n15695;
  wire n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703;
  wire n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711;
  wire n15712, n15715, n15716, n15717, n15718, n15719, n15720, n15721;
  wire n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15731;
  wire n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15743;
  wire n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15768;
  wire n15769, n15785, n15786, n15787, n15788, n15789, n15790, n15791;
  wire n15792, n15795, n15796, n15810, n15811, n15812, n15813, n15814;
  wire n15815, n15816, n15817, n15820, n15821, n15826, n15842, n15843;
  wire n15844, n15845, n15846, n15847, n15848, n15851, n15852, n15853;
  wire n15854, n15867, n15880, n15881, n15882, n15899, n15900, n15901;
  wire n15902, n15903, n15904, n15905, n15906, n15909, n15910, n15924;
  wire n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945;
  wire n15948, n15949, n15953, n15956, n15970, n15984, n15985, n15986;
  wire n15987, n15988, n15989, n15990, n15993, n15994, n16008, n16009;
  wire n16010, n16011, n16012, n16013, n16014, n16017, n16018, n16019;
  wire n16020, n16031, n16049, n16055, n16067, n16081, n16082, n16083;
  wire n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091;
  wire n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16101;
  wire n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109;
  wire n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117;
  wire n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125;
  wire n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133;
  wire n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141;
  wire n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149;
  wire n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157;
  wire n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165;
  wire n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173;
  wire n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183;
  wire n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191;
  wire n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201;
  wire n16202, n16203, n16204, n16205, n16206, n16207, n16210, n16211;
  wire n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219;
  wire n16220, n16221, n16222, n16223, n16224, n16225, n16228, n16229;
  wire n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237;
  wire n16238, n16239, n16240, n16241, n16244, n16245, n16246, n16247;
  wire n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255;
  wire n16256, n16257, n16258, n16259, n16262, n16263, n16264, n16265;
  wire n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273;
  wire n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281;
  wire n16282, n16283, n16284, n16285, n16286, n16289, n16290, n16291;
  wire n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299;
  wire n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307;
  wire n16308, n16309, n16310, n16313, n16314, n16315, n16316, n16317;
  wire n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325;
  wire n16326, n16327, n16330, n16331, n16332, n16333, n16334, n16335;
  wire n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16345;
  wire n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353;
  wire n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16363;
  wire n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371;
  wire n16372, n16373, n16374, n16375, n16376, n16379, n16380, n16381;
  wire n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389;
  wire n16390, n16391, n16392, n16393, n16394, n16397, n16398, n16399;
  wire n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407;
  wire n16408, n16409, n16410, n16413, n16414, n16415, n16416, n16417;
  wire n16418, n16419, n16420, n16421, n16422, n16423, n16426, n16427;
  wire n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435;
  wire n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443;
  wire n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451;
  wire n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461;
  wire n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469;
  wire n16470, n16471, n16472, n16473, n16474, n16477, n16478, n16479;
  wire n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487;
  wire n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16497;
  wire n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505;
  wire n16506, n16507, n16508, n16509, n16512, n16513, n16514, n16515;
  wire n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523;
  wire n16524, n16525, n16528, n16529, n16530, n16531, n16532, n16533;
  wire n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541;
  wire n16542, n16543, n16546, n16547, n16548, n16549, n16550, n16551;
  wire n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559;
  wire n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569;
  wire n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577;
  wire n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587;
  wire n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595;
  wire n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603;
  wire n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611;
  wire n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16621;
  wire n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629;
  wire n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637;
  wire n16638, n16639, n16640, n16641, n16644, n16645, n16646, n16647;
  wire n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655;
  wire n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663;
  wire n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671;
  wire n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679;
  wire n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687;
  wire n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695;
  wire n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703;
  wire n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711;
  wire n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719;
  wire n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727;
  wire n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735;
  wire n16736, n16737, n16740, n16741, n16742, n16743, n16744, n16745;
  wire n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753;
  wire n16754, n16755, n16758, n16759, n16760, n16761, n16762, n16763;
  wire n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771;
  wire n16772, n16773, n16776, n16777, n16778, n16779, n16780, n16781;
  wire n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789;
  wire n16790, n16791, n16794, n16795, n16796, n16797, n16798, n16799;
  wire n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807;
  wire n16808, n16809, n16812, n16813, n16814, n16815, n16816, n16817;
  wire n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825;
  wire n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833;
  wire n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841;
  wire n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849;
  wire n16850, n16851, n16852, n16853, n16856, n16857, n16858, n16859;
  wire n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867;
  wire n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875;
  wire n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883;
  wire n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891;
  wire n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899;
  wire n16900, n16901, n16902, n16903, n16904, n16907, n16908, n16909;
  wire n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917;
  wire n16918, n16919, n16920, n16923, n16924, n16925, n16926, n16927;
  wire n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935;
  wire n16936, n16939, n16940, n16941, n16942, n16943, n16944, n16945;
  wire n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953;
  wire n16954, n16957, n16958, n16959, n16960, n16961, n16962, n16963;
  wire n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16973;
  wire n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981;
  wire n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16991;
  wire n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999;
  wire n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007;
  wire n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015;
  wire n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025;
  wire n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033;
  wire n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041;
  wire n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049;
  wire n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057;
  wire n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065;
  wire n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073;
  wire n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081;
  wire n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089;
  wire n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097;
  wire n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105;
  wire n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113;
  wire n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121;
  wire n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129;
  wire n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137;
  wire n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145;
  wire n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153;
  wire n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161;
  wire n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169;
  wire n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177;
  wire n17178, n17179, n17180, n17183, n17184, n17185, n17186, n17187;
  wire n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195;
  wire n17196, n17197, n17200, n17201, n17202, n17203, n17204, n17205;
  wire n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213;
  wire n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221;
  wire n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229;
  wire n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237;
  wire n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245;
  wire n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253;
  wire n17254, n17255, n17256, n17259, n17260, n17261, n17262, n17263;
  wire n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271;
  wire n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279;
  wire n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287;
  wire n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295;
  wire n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303;
  wire n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311;
  wire n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319;
  wire n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327;
  wire n17328, n17329, n17332, n17333, n17334, n17335, n17336, n17337;
  wire n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345;
  wire n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355;
  wire n17356, n17357, n17358, n17359, n17360, n17361, n17364, n17365;
  wire n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373;
  wire n17374, n17375, n17376, n17377, n17378, n17379, n17382, n17383;
  wire n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391;
  wire n17392, n17393, n17394, n17395, n17398, n17399, n17400, n17401;
  wire n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17411;
  wire n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419;
  wire n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427;
  wire n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435;
  wire n17436, n17439, n17440, n17441, n17442, n17443, n17444, n17445;
  wire n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453;
  wire n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17463;
  wire n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471;
  wire n17472, n17473, n17474, n17475, n17476, n17477, n17480, n17481;
  wire n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489;
  wire n17490, n17491, n17492, n17493, n17494, n17495, n17498, n17499;
  wire n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507;
  wire n17508, n17509, n17510, n17511, n17512, n17513, n17516, n17517;
  wire n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525;
  wire n17526, n17527, n17528, n17529, n17530, n17531, n17534, n17535;
  wire n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543;
  wire n17544, n17545, n17546, n17547, n17548, n17549, n17552, n17553;
  wire n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561;
  wire n17562, n17563, n17564, n17565, n17566, n17567, n17570, n17571;
  wire n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579;
  wire n17580, n17581, n17582, n17583, n17584, n17585, n17588, n17589;
  wire n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597;
  wire n17598, n17599, n17600, n17601, n17602, n17603, n17606, n17607;
  wire n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615;
  wire n17616, n17617, n17618, n17619, n17620, n17621, n17624, n17625;
  wire n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633;
  wire n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641;
  wire n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649;
  wire n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657;
  wire n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665;
  wire n17666, n17667, n17670, n17671, n17672, n17673, n17674, n17675;
  wire n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683;
  wire n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691;
  wire n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699;
  wire n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709;
  wire n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717;
  wire n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725;
  wire n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733;
  wire n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741;
  wire n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749;
  wire n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757;
  wire n17758, n17761, n17762, n17763, n17764, n17765, n17766, n17767;
  wire n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775;
  wire n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783;
  wire n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791;
  wire n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799;
  wire n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807;
  wire n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815;
  wire n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825;
  wire n17826, n17827, n17828, n17829, n17830, n17831, n17834, n17835;
  wire n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843;
  wire n17844, n17845, n17846, n17847, n17850, n17851, n17852, n17853;
  wire n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861;
  wire n17862, n17863, n17864, n17865, n17868, n17869, n17870, n17871;
  wire n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879;
  wire n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887;
  wire n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895;
  wire n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903;
  wire n17904, n17905, n17906, n17909, n17910, n17911, n17912, n17913;
  wire n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921;
  wire n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929;
  wire n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937;
  wire n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945;
  wire n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953;
  wire n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961;
  wire n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969;
  wire n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977;
  wire n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985;
  wire n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993;
  wire n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001;
  wire n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009;
  wire n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017;
  wire n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025;
  wire n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033;
  wire n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041;
  wire n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049;
  wire n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057;
  wire n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065;
  wire n18066, n18067, n18068, n18069, n18070, n18073, n18074, n18075;
  wire n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083;
  wire n18084, n18085, n18086, n18087, n18090, n18091, n18092, n18093;
  wire n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101;
  wire n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109;
  wire n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117;
  wire n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125;
  wire n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133;
  wire n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141;
  wire n18142, n18143, n18144, n18145, n18146, n18147, n18150, n18151;
  wire n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159;
  wire n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167;
  wire n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175;
  wire n18176, n18177, n18178, n18179, n18182, n18183, n18184, n18185;
  wire n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193;
  wire n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201;
  wire n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209;
  wire n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217;
  wire n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225;
  wire n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233;
  wire n18234, n18235, n18236, n18237, n18238, n18241, n18242, n18243;
  wire n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251;
  wire n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259;
  wire n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267;
  wire n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275;
  wire n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283;
  wire n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291;
  wire n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299;
  wire n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307;
  wire n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315;
  wire n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323;
  wire n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331;
  wire n18332, n18333, n18336, n18337, n18338, n18339, n18340, n18341;
  wire n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349;
  wire n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359;
  wire n18360, n18361, n18362, n18363, n18364, n18365, n18368, n18369;
  wire n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377;
  wire n18378, n18379, n18380, n18381, n18382, n18383, n18386, n18387;
  wire n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395;
  wire n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403;
  wire n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411;
  wire n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421;
  wire n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18431;
  wire n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439;
  wire n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18449;
  wire n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457;
  wire n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18467;
  wire n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475;
  wire n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18485;
  wire n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493;
  wire n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18503;
  wire n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511;
  wire n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18521;
  wire n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529;
  wire n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18539;
  wire n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547;
  wire n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18557;
  wire n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565;
  wire n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18575;
  wire n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583;
  wire n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591;
  wire n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599;
  wire n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607;
  wire n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615;
  wire n18616, n18617, n18618, n18621, n18622, n18623, n18624, n18625;
  wire n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633;
  wire n18634, n18635, n18638, n18639, n18640, n18641, n18642, n18643;
  wire n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651;
  wire n18652, n18653, n18656, n18657, n18658, n18659, n18660, n18661;
  wire n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669;
  wire n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677;
  wire n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685;
  wire n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693;
  wire n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701;
  wire n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709;
  wire n18710, n18711, n18712, n18713, n18716, n18717, n18718, n18719;
  wire n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727;
  wire n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735;
  wire n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743;
  wire n18744, n18745, n18748, n18749, n18750, n18751, n18752, n18753;
  wire n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761;
  wire n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769;
  wire n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777;
  wire n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785;
  wire n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793;
  wire n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801;
  wire n18802, n18803, n18804, n18807, n18808, n18809, n18810, n18811;
  wire n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819;
  wire n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827;
  wire n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835;
  wire n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843;
  wire n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851;
  wire n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859;
  wire n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867;
  wire n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875;
  wire n18876, n18877, n18878, n18879, n18880, n18881, n18884, n18885;
  wire n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893;
  wire n18894, n18895, n18896, n18897, n18900, n18901, n18902, n18903;
  wire n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911;
  wire n18912, n18913, n18916, n18917, n18918, n18919, n18920, n18921;
  wire n18922, n18923, n18924, n18925, n18926, n18929, n18930, n18931;
  wire n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939;
  wire n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947;
  wire n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955;
  wire n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963;
  wire n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971;
  wire n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979;
  wire n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987;
  wire n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995;
  wire n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003;
  wire n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011;
  wire n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019;
  wire n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027;
  wire n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035;
  wire n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043;
  wire n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051;
  wire n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059;
  wire n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067;
  wire n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075;
  wire n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083;
  wire n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091;
  wire n19092, n19093, n19094, n19095, n19098, n19099, n19100, n19101;
  wire n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109;
  wire n19110, n19111, n19112, n19115, n19116, n19117, n19118, n19119;
  wire n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127;
  wire n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135;
  wire n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143;
  wire n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151;
  wire n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159;
  wire n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167;
  wire n19168, n19169, n19170, n19171, n19172, n19175, n19176, n19177;
  wire n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185;
  wire n19186, n19187, n19188, n19189, n19192, n19193, n19194, n19195;
  wire n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203;
  wire n19204, n19205, n19206, n19207, n19210, n19211, n19212, n19213;
  wire n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221;
  wire n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229;
  wire n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237;
  wire n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245;
  wire n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253;
  wire n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261;
  wire n19262, n19263, n19264, n19265, n19266, n19267, n19270, n19271;
  wire n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279;
  wire n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287;
  wire n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295;
  wire n19296, n19297, n19298, n19299, n19302, n19303, n19304, n19305;
  wire n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313;
  wire n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321;
  wire n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329;
  wire n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337;
  wire n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345;
  wire n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353;
  wire n19354, n19355, n19356, n19357, n19358, n19361, n19362, n19363;
  wire n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371;
  wire n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379;
  wire n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387;
  wire n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395;
  wire n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403;
  wire n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411;
  wire n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419;
  wire n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427;
  wire n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435;
  wire n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443;
  wire n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451;
  wire n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459;
  wire n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467;
  wire n19468, n19469, n19470, n19471, n19472, n19473, n19476, n19477;
  wire n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485;
  wire n19486, n19487, n19488, n19489, n19492, n19493, n19494, n19495;
  wire n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503;
  wire n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511;
  wire n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519;
  wire n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527;
  wire n19528, n19529, n19530, n19531, n19534, n19535, n19536, n19537;
  wire n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545;
  wire n19546, n19547, n19548, n19551, n19552, n19553, n19554, n19555;
  wire n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563;
  wire n19564, n19565, n19566, n19569, n19570, n19571, n19572, n19573;
  wire n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581;
  wire n19582, n19583, n19584, n19587, n19588, n19589, n19590, n19591;
  wire n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599;
  wire n19600, n19601, n19602, n19605, n19606, n19607, n19608, n19609;
  wire n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617;
  wire n19618, n19619, n19620, n19623, n19624, n19625, n19626, n19627;
  wire n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635;
  wire n19636, n19637, n19638, n19641, n19642, n19643, n19644, n19645;
  wire n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653;
  wire n19654, n19655, n19656, n19659, n19660, n19661, n19662, n19663;
  wire n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671;
  wire n19672, n19673, n19674, n19677, n19678, n19679, n19680, n19681;
  wire n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689;
  wire n19690, n19691, n19692, n19695, n19696, n19697, n19698, n19699;
  wire n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707;
  wire n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715;
  wire n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723;
  wire n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731;
  wire n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19741;
  wire n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749;
  wire n19750, n19751, n19752, n19753, n19754, n19755, n19758, n19759;
  wire n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767;
  wire n19768, n19769, n19770, n19771, n19772, n19773, n19776, n19777;
  wire n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785;
  wire n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793;
  wire n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801;
  wire n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809;
  wire n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817;
  wire n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825;
  wire n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833;
  wire n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843;
  wire n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19853;
  wire n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861;
  wire n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19871;
  wire n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879;
  wire n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887;
  wire n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895;
  wire n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903;
  wire n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911;
  wire n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919;
  wire n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927;
  wire n19928, n19931, n19932, n19933, n19934, n19935, n19936, n19937;
  wire n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945;
  wire n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953;
  wire n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19963;
  wire n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971;
  wire n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979;
  wire n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987;
  wire n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995;
  wire n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003;
  wire n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011;
  wire n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019;
  wire n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029;
  wire n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037;
  wire n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045;
  wire n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053;
  wire n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061;
  wire n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069;
  wire n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077;
  wire n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085;
  wire n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093;
  wire n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101;
  wire n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109;
  wire n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20119;
  wire n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127;
  wire n20128, n20129, n20130, n20131, n20132, n20135, n20136, n20137;
  wire n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145;
  wire n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153;
  wire n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161;
  wire n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169;
  wire n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177;
  wire n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185;
  wire n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193;
  wire n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201;
  wire n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209;
  wire n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217;
  wire n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225;
  wire n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233;
  wire n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241;
  wire n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249;
  wire n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257;
  wire n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265;
  wire n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273;
  wire n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281;
  wire n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289;
  wire n20290, n20291, n20292, n20293, n20294, n20297, n20298, n20299;
  wire n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307;
  wire n20308, n20309, n20310, n20311, n20314, n20315, n20316, n20317;
  wire n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325;
  wire n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333;
  wire n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341;
  wire n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349;
  wire n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357;
  wire n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365;
  wire n20366, n20367, n20368, n20369, n20370, n20371, n20374, n20375;
  wire n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383;
  wire n20384, n20385, n20386, n20387, n20388, n20391, n20392, n20393;
  wire n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401;
  wire n20402, n20403, n20404, n20405, n20406, n20409, n20410, n20411;
  wire n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419;
  wire n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427;
  wire n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435;
  wire n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443;
  wire n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451;
  wire n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459;
  wire n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20469;
  wire n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477;
  wire n20478, n20479, n20480, n20481, n20482, n20483, n20486, n20487;
  wire n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495;
  wire n20496, n20497, n20498, n20499, n20500, n20501, n20504, n20505;
  wire n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513;
  wire n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521;
  wire n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529;
  wire n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537;
  wire n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545;
  wire n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553;
  wire n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561;
  wire n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571;
  wire n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579;
  wire n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587;
  wire n20588, n20589, n20590, n20591, n20592, n20593, n20596, n20597;
  wire n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605;
  wire n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613;
  wire n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621;
  wire n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629;
  wire n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637;
  wire n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645;
  wire n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20655;
  wire n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663;
  wire n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671;
  wire n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679;
  wire n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687;
  wire n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695;
  wire n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703;
  wire n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711;
  wire n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719;
  wire n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727;
  wire n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735;
  wire n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743;
  wire n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751;
  wire n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759;
  wire n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767;
  wire n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775;
  wire n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783;
  wire n20784, n20785, n20786, n20787, n20790, n20791, n20792, n20793;
  wire n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801;
  wire n20802, n20803, n20804, n20805, n20806, n20809, n20810, n20811;
  wire n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819;
  wire n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827;
  wire n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835;
  wire n20836, n20837, n20838, n20839, n20840, n20841, n20844, n20845;
  wire n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853;
  wire n20854, n20855, n20856, n20857, n20858, n20859, n20862, n20863;
  wire n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871;
  wire n20872, n20873, n20874, n20875, n20876, n20877, n20880, n20881;
  wire n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889;
  wire n20890, n20891, n20892, n20893, n20894, n20895, n20898, n20899;
  wire n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907;
  wire n20908, n20909, n20910, n20911, n20912, n20913, n20916, n20917;
  wire n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925;
  wire n20926, n20927, n20928, n20929, n20930, n20931, n20934, n20935;
  wire n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943;
  wire n20944, n20945, n20946, n20947, n20948, n20949, n20952, n20953;
  wire n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961;
  wire n20962, n20963, n20964, n20965, n20966, n20967, n20970, n20971;
  wire n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979;
  wire n20980, n20981, n20982, n20983, n20984, n20985, n20988, n20989;
  wire n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997;
  wire n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005;
  wire n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013;
  wire n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021;
  wire n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029;
  wire n21030, n21031, n21034, n21035, n21036, n21037, n21038, n21039;
  wire n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047;
  wire n21048, n21051, n21052, n21053, n21054, n21055, n21056, n21057;
  wire n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065;
  wire n21066, n21069, n21070, n21071, n21072, n21073, n21074, n21075;
  wire n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083;
  wire n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091;
  wire n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099;
  wire n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107;
  wire n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115;
  wire n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123;
  wire n21124, n21125, n21126, n21129, n21130, n21131, n21132, n21133;
  wire n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141;
  wire n21142, n21143, n21146, n21147, n21148, n21149, n21150, n21151;
  wire n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159;
  wire n21160, n21161, n21164, n21165, n21166, n21167, n21168, n21169;
  wire n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177;
  wire n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185;
  wire n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193;
  wire n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201;
  wire n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209;
  wire n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217;
  wire n21218, n21219, n21220, n21221, n21224, n21225, n21226, n21227;
  wire n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235;
  wire n21236, n21237, n21238, n21241, n21242, n21243, n21244, n21245;
  wire n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253;
  wire n21254, n21255, n21256, n21259, n21260, n21261, n21262, n21263;
  wire n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271;
  wire n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279;
  wire n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287;
  wire n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295;
  wire n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303;
  wire n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311;
  wire n21312, n21313, n21314, n21315, n21316, n21319, n21320, n21321;
  wire n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329;
  wire n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337;
  wire n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345;
  wire n21346, n21347, n21348, n21351, n21352, n21353, n21354, n21355;
  wire n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363;
  wire n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371;
  wire n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379;
  wire n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387;
  wire n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395;
  wire n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403;
  wire n21404, n21405, n21406, n21407, n21410, n21411, n21412, n21413;
  wire n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421;
  wire n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429;
  wire n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437;
  wire n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445;
  wire n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453;
  wire n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461;
  wire n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469;
  wire n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477;
  wire n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485;
  wire n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493;
  wire n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501;
  wire n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509;
  wire n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517;
  wire n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525;
  wire n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533;
  wire n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541;
  wire n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549;
  wire n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557;
  wire n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565;
  wire n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573;
  wire n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581;
  wire n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589;
  wire n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597;
  wire n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605;
  wire n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613;
  wire n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621;
  wire n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629;
  wire n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637;
  wire n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645;
  wire n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653;
  wire n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661;
  wire n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21674;
  wire n21675, n21676, n21677, n21678, n21679, n21682, n21683, n21684;
  wire n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692;
  wire n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700;
  wire n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708;
  wire n21709, n21710, n21713, n21714, n21715, n21716, n21717, n21718;
  wire n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726;
  wire n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734;
  wire n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21744;
  wire n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752;
  wire n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760;
  wire n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768;
  wire n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776;
  wire n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784;
  wire n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792;
  wire n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800;
  wire n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808;
  wire n21809, n21812, n21813, n21814, n21815, n21816, n21817, n21818;
  wire n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826;
  wire n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836;
  wire n21837, n21838, n21839, n21840, n21843, n21844, n21845, n21846;
  wire n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854;
  wire n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862;
  wire n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870;
  wire n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878;
  wire n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886;
  wire n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894;
  wire n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902;
  wire n21903, n21904, n21905, n21906, n21907, n21908, n21911, n21912;
  wire n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920;
  wire n21921, n21922, n21923, n21924, n21925, n21928, n21929, n21930;
  wire n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938;
  wire n21939, n21942, n21943, n21944, n21945, n21946, n21947, n21948;
  wire n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956;
  wire n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964;
  wire n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972;
  wire n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980;
  wire n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988;
  wire n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996;
  wire n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004;
  wire n22005, n22006, n22007, n22010, n22011, n22012, n22013, n22014;
  wire n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022;
  wire n22023, n22024, n22027, n22028, n22029, n22030, n22031, n22032;
  wire n22033, n22034, n22035, n22036, n22037, n22038, n22041, n22042;
  wire n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050;
  wire n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058;
  wire n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066;
  wire n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074;
  wire n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082;
  wire n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090;
  wire n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098;
  wire n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106;
  wire n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116;
  wire n22117, n22118, n22119, n22120, n22123, n22124, n22125, n22126;
  wire n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134;
  wire n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142;
  wire n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150;
  wire n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158;
  wire n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166;
  wire n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174;
  wire n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182;
  wire n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190;
  wire n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198;
  wire n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206;
  wire n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214;
  wire n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222;
  wire n22223, n22224, n22225, n22226, n22227, n22230, n22231, n22232;
  wire n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240;
  wire n22241, n22242, n22243, n22246, n22247, n22248, n22249, n22250;
  wire n22251, n22252, n22268, n22269, n22270, n22271, n22272, n22273;
  wire n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281;
  wire n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22291;
  wire n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299;
  wire n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307;
  wire n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315;
  wire n22316, n22319, n22320, n22321, n22322, n22323, n22324, n22325;
  wire n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333;
  wire n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341;
  wire n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349;
  wire n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357;
  wire n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365;
  wire n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373;
  wire n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381;
  wire n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389;
  wire n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397;
  wire n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405;
  wire n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413;
  wire n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421;
  wire n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429;
  wire n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437;
  wire n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445;
  wire n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453;
  wire n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461;
  wire n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469;
  wire n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477;
  wire n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485;
  wire n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493;
  wire n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501;
  wire n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509;
  wire n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517;
  wire n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525;
  wire n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533;
  wire n22534, n22535, n22536, n22537, n22538, n22541, n22542, n22543;
  wire n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551;
  wire n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561;
  wire n22562, n22563, n22564, n22565, n22568, n22569, n22570, n22571;
  wire n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22581;
  wire n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589;
  wire n22590, n22591, n22594, n22595, n22596, n22597, n22598, n22599;
  wire n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607;
  wire n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615;
  wire n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623;
  wire n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631;
  wire n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639;
  wire n22640, n22641, n22642, n22643, n22644, n22645, n22648, n22649;
  wire n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657;
  wire n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665;
  wire n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673;
  wire n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681;
  wire n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689;
  wire n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697;
  wire n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705;
  wire n22706, n22707, n22708, n22711, n22712, n22713, n22714, n22715;
  wire n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723;
  wire n22724, n22725, n22726, n22727, n22728, n22729, n22732, n22733;
  wire n22734, n22735, n22736, n22737, n22748, n22762, n22779, n22780;
  wire n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788;
  wire n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796;
  wire n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804;
  wire n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812;
  wire n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820;
  wire n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828;
  wire n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836;
  wire n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844;
  wire n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852;
  wire n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22862;
  wire n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870;
  wire n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878;
  wire n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886;
  wire n22887, n22888, n22889, n22890, n22891, n22894, n22895, n22896;
  wire n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904;
  wire n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912;
  wire n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920;
  wire n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928;
  wire n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936;
  wire n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944;
  wire n22945, n22946, n22947, n22948, n22949, n22950, n22953, n22954;
  wire n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962;
  wire n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970;
  wire n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978;
  wire n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986;
  wire n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994;
  wire n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002;
  wire n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012;
  wire n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020;
  wire n23021, n23024, n23025, n23026, n23027, n23028, n23029, n23030;
  wire n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038;
  wire n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046;
  wire n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054;
  wire n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062;
  wire n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070;
  wire n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078;
  wire n23079, n23080, n23081, n23082, n23083, n23086, n23087, n23088;
  wire n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096;
  wire n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104;
  wire n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112;
  wire n23113, n23114, n23115, n23118, n23119, n23120, n23121, n23122;
  wire n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130;
  wire n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138;
  wire n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146;
  wire n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154;
  wire n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162;
  wire n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170;
  wire n23171, n23172, n23173, n23174, n23177, n23178, n23179, n23180;
  wire n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188;
  wire n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196;
  wire n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204;
  wire n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212;
  wire n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220;
  wire n23221, n23222, n23225, n23226, n23227, n23228, n23229, n23230;
  wire n23231, n23232, n23233, n23234, n23237, n23238, n23239, n23240;
  wire n23241, n23242, n23243, n23244, n23245, n23246, n23249, n23250;
  wire n23251, n23269, n23270, n23271, n23272, n23273, n23274, n23275;
  wire n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283;
  wire n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291;
  wire n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299;
  wire n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307;
  wire n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315;
  wire n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323;
  wire n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331;
  wire n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339;
  wire n23340, n23343, n23344, n23345, n23346, n23347, n23348, n23349;
  wire n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357;
  wire n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365;
  wire n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373;
  wire n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381;
  wire n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389;
  wire n23390, n23391, n23394, n23395, n23396, n23397, n23398, n23399;
  wire n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407;
  wire n23408, n23411, n23412, n23413, n23414, n23415, n23416, n23417;
  wire n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425;
  wire n23426, n23429, n23430, n23431, n23432, n23433, n23434, n23435;
  wire n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443;
  wire n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451;
  wire n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459;
  wire n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467;
  wire n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475;
  wire n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483;
  wire n23484, n23485, n23486, n23489, n23490, n23491, n23492, n23493;
  wire n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501;
  wire n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509;
  wire n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517;
  wire n23518, n23521, n23522, n23523, n23524, n23525, n23526, n23527;
  wire n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535;
  wire n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543;
  wire n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551;
  wire n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559;
  wire n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567;
  wire n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575;
  wire n23576, n23577, n23580, n23581, n23582, n23583, n23584, n23585;
  wire n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593;
  wire n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601;
  wire n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609;
  wire n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617;
  wire n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625;
  wire n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633;
  wire n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641;
  wire n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649;
  wire n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657;
  wire n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665;
  wire n23666, n23667, n23668, n23671, n23672, n23673, n23674, n23675;
  wire n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683;
  wire n23684, n23685, n23686, n23687, n23690, n23691, n23692, n23693;
  wire n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701;
  wire n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709;
  wire n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717;
  wire n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725;
  wire n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733;
  wire n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741;
  wire n23742, n23743, n23744, n23745, n23746, n23747, n23750, n23751;
  wire n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759;
  wire n23760, n23761, n23762, n23763, n23764, n23767, n23768, n23769;
  wire n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777;
  wire n23778, n23779, n23780, n23781, n23782, n23785, n23786, n23787;
  wire n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795;
  wire n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803;
  wire n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811;
  wire n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819;
  wire n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827;
  wire n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835;
  wire n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23845;
  wire n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853;
  wire n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861;
  wire n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869;
  wire n23870, n23871, n23872, n23873, n23874, n23877, n23878, n23879;
  wire n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887;
  wire n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895;
  wire n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903;
  wire n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911;
  wire n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919;
  wire n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927;
  wire n23928, n23929, n23930, n23931, n23932, n23933, n23936, n23937;
  wire n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945;
  wire n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953;
  wire n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961;
  wire n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969;
  wire n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977;
  wire n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985;
  wire n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993;
  wire n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001;
  wire n24002, n24003, n24004, n24005, n24006, n24009, n24010, n24011;
  wire n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24021;
  wire n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029;
  wire n24030, n24033, n24034, n24035, n24036, n24037, n24038, n24039;
  wire n24040, n24041, n24057, n24058, n24059, n24060, n24061, n24064;
  wire n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072;
  wire n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080;
  wire n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088;
  wire n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096;
  wire n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104;
  wire n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112;
  wire n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120;
  wire n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128;
  wire n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136;
  wire n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144;
  wire n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152;
  wire n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160;
  wire n24161, n24162, n24165, n24166, n24167, n24168, n24169, n24170;
  wire n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178;
  wire n24179, n24180, n24181, n24182, n24183, n24186, n24187, n24188;
  wire n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196;
  wire n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204;
  wire n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212;
  wire n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220;
  wire n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228;
  wire n24229, n24230, n24231, n24232, n24235, n24236, n24237, n24238;
  wire n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246;
  wire n24247, n24248, n24249, n24252, n24253, n24254, n24255, n24256;
  wire n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264;
  wire n24265, n24266, n24267, n24270, n24271, n24272, n24273, n24274;
  wire n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282;
  wire n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290;
  wire n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298;
  wire n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306;
  wire n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314;
  wire n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322;
  wire n24323, n24324, n24325, n24326, n24327, n24330, n24331, n24332;
  wire n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340;
  wire n24341, n24342, n24343, n24344, n24347, n24348, n24349, n24350;
  wire n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358;
  wire n24359, n24360, n24361, n24362, n24365, n24366, n24367, n24368;
  wire n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376;
  wire n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384;
  wire n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392;
  wire n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400;
  wire n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408;
  wire n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416;
  wire n24417, n24418, n24419, n24420, n24421, n24422, n24425, n24426;
  wire n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434;
  wire n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442;
  wire n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450;
  wire n24451, n24452, n24453, n24454, n24457, n24458, n24459, n24460;
  wire n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468;
  wire n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476;
  wire n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484;
  wire n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492;
  wire n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500;
  wire n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508;
  wire n24509, n24510, n24511, n24512, n24513, n24516, n24517, n24518;
  wire n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526;
  wire n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534;
  wire n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542;
  wire n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550;
  wire n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558;
  wire n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566;
  wire n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574;
  wire n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582;
  wire n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590;
  wire n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598;
  wire n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606;
  wire n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614;
  wire n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622;
  wire n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630;
  wire n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638;
  wire n24639, n24640, n24641, n24642, n24645, n24646, n24647, n24648;
  wire n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656;
  wire n24657, n24658, n24659, n24662, n24663, n24664, n24665, n24666;
  wire n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674;
  wire n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682;
  wire n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690;
  wire n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698;
  wire n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706;
  wire n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714;
  wire n24715, n24716, n24717, n24718, n24719, n24722, n24723, n24724;
  wire n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732;
  wire n24733, n24734, n24735, n24736, n24739, n24740, n24741, n24742;
  wire n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750;
  wire n24751, n24752, n24753, n24754, n24757, n24758, n24759, n24760;
  wire n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768;
  wire n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776;
  wire n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784;
  wire n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792;
  wire n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800;
  wire n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808;
  wire n24809, n24810, n24811, n24812, n24813, n24814, n24817, n24818;
  wire n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826;
  wire n24827, n24828, n24829, n24830, n24831, n24834, n24835, n24836;
  wire n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844;
  wire n24845, n24846, n24847, n24848, n24849, n24852, n24853, n24854;
  wire n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862;
  wire n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870;
  wire n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878;
  wire n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886;
  wire n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894;
  wire n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902;
  wire n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24912;
  wire n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920;
  wire n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928;
  wire n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936;
  wire n24937, n24938, n24939, n24940, n24941, n24944, n24945, n24946;
  wire n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954;
  wire n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962;
  wire n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970;
  wire n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978;
  wire n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986;
  wire n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994;
  wire n24995, n24996, n24997, n24998, n24999, n25000, n25003, n25004;
  wire n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012;
  wire n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020;
  wire n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028;
  wire n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036;
  wire n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044;
  wire n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052;
  wire n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060;
  wire n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068;
  wire n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076;
  wire n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084;
  wire n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092;
  wire n25093, n25094, n25095, n25096, n25097, n25098, n25101, n25102;
  wire n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110;
  wire n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120;
  wire n25121, n25122, n25125, n25126, n25127, n25128, n25129, n25130;
  wire n25131, n25132, n25133, n25134, n25137, n25138, n25139, n25140;
  wire n25141, n25142, n25143, n25157, n25158, n25159, n25160, n25161;
  wire n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171;
  wire n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179;
  wire n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187;
  wire n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195;
  wire n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203;
  wire n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211;
  wire n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219;
  wire n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227;
  wire n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235;
  wire n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243;
  wire n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251;
  wire n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259;
  wire n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267;
  wire n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275;
  wire n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283;
  wire n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25293;
  wire n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301;
  wire n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309;
  wire n25310, n25313, n25314, n25315, n25316, n25317, n25318, n25319;
  wire n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327;
  wire n25328, n25329, n25330, n25331, n25334, n25335, n25336, n25337;
  wire n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345;
  wire n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353;
  wire n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361;
  wire n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369;
  wire n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377;
  wire n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387;
  wire n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25397;
  wire n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405;
  wire n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25415;
  wire n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423;
  wire n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431;
  wire n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439;
  wire n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447;
  wire n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455;
  wire n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463;
  wire n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471;
  wire n25472, n25475, n25476, n25477, n25478, n25479, n25480, n25481;
  wire n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489;
  wire n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499;
  wire n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507;
  wire n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517;
  wire n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525;
  wire n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533;
  wire n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541;
  wire n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549;
  wire n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557;
  wire n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565;
  wire n25566, n25567, n25570, n25571, n25572, n25573, n25574, n25575;
  wire n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583;
  wire n25584, n25587, n25588, n25589, n25590, n25591, n25592, n25593;
  wire n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601;
  wire n25602, n25605, n25606, n25607, n25608, n25609, n25610, n25611;
  wire n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619;
  wire n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627;
  wire n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635;
  wire n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643;
  wire n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651;
  wire n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659;
  wire n25660, n25661, n25662, n25665, n25666, n25667, n25668, n25669;
  wire n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677;
  wire n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685;
  wire n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693;
  wire n25694, n25697, n25698, n25699, n25700, n25701, n25702, n25703;
  wire n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711;
  wire n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719;
  wire n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727;
  wire n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735;
  wire n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743;
  wire n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751;
  wire n25752, n25753, n25756, n25757, n25758, n25759, n25760, n25761;
  wire n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769;
  wire n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777;
  wire n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785;
  wire n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793;
  wire n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801;
  wire n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809;
  wire n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817;
  wire n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825;
  wire n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833;
  wire n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841;
  wire n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849;
  wire n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25863;
  wire n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881;
  wire n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891;
  wire n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899;
  wire n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907;
  wire n25908, n25909, n25910, n25913, n25914, n25915, n25916, n25917;
  wire n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25927;
  wire n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947;
  wire n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955;
  wire n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963;
  wire n25964, n25965, n25966, n25967, n25968, n25969, n25972, n25973;
  wire n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981;
  wire n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989;
  wire n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997;
  wire n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005;
  wire n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015;
  wire n26016, n26021, n26022, n26023, n26024, n26025, n26026, n26027;
  wire n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035;
  wire n26036, n26037, n26040, n26041, n26042, n26043, n26044, n26045;
  wire n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053;
  wire n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061;
  wire n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069;
  wire n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077;
  wire n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085;
  wire n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093;
  wire n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101;
  wire n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109;
  wire n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117;
  wire n26123, n26124, n26125, n26126, n26127, n26128, n26131, n26132;
  wire n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140;
  wire n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148;
  wire n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156;
  wire n26157, n26158, n26159, n26162, n26163, n26164, n26165, n26166;
  wire n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174;
  wire n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182;
  wire n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190;
  wire n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200;
  wire n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208;
  wire n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216;
  wire n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224;
  wire n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232;
  wire n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240;
  wire n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248;
  wire n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256;
  wire n26257, n26258, n26261, n26262, n26263, n26264, n26265, n26266;
  wire n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274;
  wire n26275, n26278, n26279, n26280, n26281, n26282, n26283, n26284;
  wire n26285, n26286, n26287, n26288, n26289, n26292, n26293, n26294;
  wire n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302;
  wire n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310;
  wire n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318;
  wire n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326;
  wire n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334;
  wire n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342;
  wire n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350;
  wire n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26360;
  wire n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368;
  wire n26369, n26370, n26371, n26372, n26373, n26374, n26377, n26378;
  wire n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386;
  wire n26387, n26388, n26391, n26392, n26393, n26394, n26395, n26396;
  wire n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404;
  wire n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412;
  wire n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420;
  wire n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428;
  wire n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436;
  wire n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444;
  wire n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452;
  wire n26453, n26454, n26455, n26456, n26459, n26460, n26461, n26462;
  wire n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470;
  wire n26471, n26472, n26473, n26476, n26477, n26478, n26479, n26480;
  wire n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26490;
  wire n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498;
  wire n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506;
  wire n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514;
  wire n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522;
  wire n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530;
  wire n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538;
  wire n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546;
  wire n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554;
  wire n26555, n26558, n26559, n26560, n26561, n26562, n26563, n26564;
  wire n26565, n26566, n26567, n26568, n26569, n26572, n26573, n26574;
  wire n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582;
  wire n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590;
  wire n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598;
  wire n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606;
  wire n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614;
  wire n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622;
  wire n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630;
  wire n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638;
  wire n26639, n26640, n26641, n26642, n26643, n26646, n26647, n26648;
  wire n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26658;
  wire n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666;
  wire n26667, n26670, n26671, n26672, n26673, n26674, n26675, n26676;
  wire n26677, n26678, n26679, n26682, n26683, n26684, n26685, n26686;
  wire n26687, n26688, n26689, n26690, n26691, n26694, n26695, n26696;
  wire n26697, n26698, n26699, n26700, n26715, n26716, n26717, n26718;
  wire n26719, n26722, n26723, n26724, n26725, n26726, n26727, n26728;
  wire n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736;
  wire n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744;
  wire n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752;
  wire n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760;
  wire n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768;
  wire n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776;
  wire n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784;
  wire n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792;
  wire n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800;
  wire n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808;
  wire n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816;
  wire n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824;
  wire n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832;
  wire n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840;
  wire n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848;
  wire n26849, n26850, n26851, n26852, n26855, n26856, n26859, n26860;
  wire n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868;
  wire n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876;
  wire n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884;
  wire n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892;
  wire n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900;
  wire n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908;
  wire n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916;
  wire n26917, n26918, n26919, n26920, n26922, n26923, n26924, n26925;
  wire n26926, n26929, n26930, n26931, n26932, n26933, n26934, n26935;
  wire n26936, n26937, n26938, n26941, n26942, n26943, n26944, n26945;
  wire n26946, n26947, n26948, n26949, n26950, n26953, n26954, n26955;
  wire n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26965;
  wire n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973;
  wire n26991, n26992, n26993, n26994, n26995, n26998, n26999, n27000;
  wire n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008;
  wire n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016;
  wire n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024;
  wire n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032;
  wire n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040;
  wire n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048;
  wire n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056;
  wire n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064;
  wire n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072;
  wire n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080;
  wire n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088;
  wire n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096;
  wire n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104;
  wire n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112;
  wire n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120;
  wire n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128;
  wire n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136;
  wire n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144;
  wire n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152;
  wire n27153, n27154, n27155, n27156, n27157, n27160, n27161, n27162;
  wire n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170;
  wire n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178;
  wire n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186;
  wire n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194;
  wire n27195, n27196, n27197, n27198, n27200, n27201, n27202, n27203;
  wire n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213;
  wire n27214, n27215, n27218, n27219, n27220, n27221, n27222, n27223;
  wire n27224, n27225, n27226, n27227, n27230, n27231, n27232, n27233;
  wire n27234, n27235, n27236, n27237, n27238, n27239, n27242, n27243;
  wire n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27267;
  wire n27268, n27269, n27270, n27271, n27274, n27275, n27276, n27277;
  wire n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285;
  wire n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293;
  wire n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301;
  wire n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309;
  wire n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317;
  wire n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325;
  wire n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333;
  wire n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341;
  wire n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349;
  wire n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357;
  wire n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365;
  wire n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373;
  wire n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381;
  wire n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389;
  wire n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397;
  wire n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405;
  wire n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413;
  wire n27414, n27417, n27418, n27419, n27420, n27421, n27422, n27423;
  wire n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431;
  wire n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439;
  wire n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447;
  wire n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455;
  wire n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463;
  wire n27464, n27465, n27466, n27467, n27468, n27470, n27471, n27472;
  wire n27473, n27476, n27477, n27478, n27479, n27480, n27481, n27482;
  wire n27483, n27484, n27485, n27488, n27489, n27490, n27491, n27492;
  wire n27493, n27494, n27495, n27496, n27497, n27500, n27501, n27502;
  wire n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27512;
  wire n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520;
  wire n27521, n27522, n27535, n27536, n27537, n27538, n27539, n27542;
  wire n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550;
  wire n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558;
  wire n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566;
  wire n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574;
  wire n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582;
  wire n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590;
  wire n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598;
  wire n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606;
  wire n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614;
  wire n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622;
  wire n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630;
  wire n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638;
  wire n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646;
  wire n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654;
  wire n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662;
  wire n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670;
  wire n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678;
  wire n27679, n27682, n27683, n27684, n27685, n27686, n27687, n27688;
  wire n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696;
  wire n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704;
  wire n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712;
  wire n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720;
  wire n27721, n27722, n27723, n27724, n27725, n27726, n27728, n27729;
  wire n27730, n27731, n27734, n27735, n27736, n27737, n27738, n27739;
  wire n27740, n27741, n27742, n27743, n27746, n27747, n27748, n27749;
  wire n27750, n27751, n27752, n27753, n27754, n27755, n27758, n27759;
  wire n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767;
  wire n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777;
  wire n27778, n27789, n27807, n27808, n27809, n27810, n27811, n27814;
  wire n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822;
  wire n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830;
  wire n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838;
  wire n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846;
  wire n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854;
  wire n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862;
  wire n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870;
  wire n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878;
  wire n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886;
  wire n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894;
  wire n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902;
  wire n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910;
  wire n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918;
  wire n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926;
  wire n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934;
  wire n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942;
  wire n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950;
  wire n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958;
  wire n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966;
  wire n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974;
  wire n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982;
  wire n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27991;
  wire n27992, n27993, n27994, n27997, n27998, n27999, n28000, n28001;
  wire n28002, n28003, n28004, n28005, n28006, n28009, n28010, n28011;
  wire n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28021;
  wire n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029;
  wire n28030, n28033, n28034, n28035, n28036, n28037, n28038, n28039;
  wire n28040, n28041, n28059, n28060, n28061, n28062, n28063, n28066;
  wire n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074;
  wire n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082;
  wire n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090;
  wire n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098;
  wire n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106;
  wire n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114;
  wire n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122;
  wire n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130;
  wire n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138;
  wire n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146;
  wire n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154;
  wire n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162;
  wire n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170;
  wire n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178;
  wire n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186;
  wire n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194;
  wire n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202;
  wire n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210;
  wire n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218;
  wire n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226;
  wire n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234;
  wire n28235, n28236, n28238, n28239, n28240, n28243, n28244, n28245;
  wire n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28255;
  wire n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263;
  wire n28264, n28267, n28268, n28269, n28270, n28271, n28272, n28273;
  wire n28274, n28275, n28276, n28279, n28280, n28281, n28282, n28283;
  wire n28284, n28285, n28286, n28287, n28294, n28314, n28315, n28316;
  wire n28317, n28318, n28321, n28322, n28323, n28324, n28325, n28326;
  wire n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334;
  wire n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342;
  wire n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350;
  wire n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358;
  wire n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366;
  wire n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374;
  wire n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382;
  wire n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390;
  wire n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398;
  wire n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406;
  wire n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414;
  wire n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422;
  wire n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430;
  wire n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438;
  wire n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446;
  wire n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454;
  wire n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462;
  wire n28463, n28464, n28465, n28467, n28468, n28469, n28470, n28471;
  wire n28474, n28492, n28493, n28494, n28495, n28496, n28497, n28498;
  wire n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506;
  wire n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514;
  wire n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522;
  wire n28523, n28524, n28525, n28526, n28527, n28528, n28531, n28532;
  wire n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540;
  wire n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28550;
  wire n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558;
  wire n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566;
  wire n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576;
  wire n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584;
  wire n28585, n28588, n28589, n28590, n28591, n28592, n28593, n28594;
  wire n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602;
  wire n28603, n28604, n28607, n28608, n28609, n28610, n28611, n28612;
  wire n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620;
  wire n28621, n28622, n28623, n28626, n28627, n28628, n28629, n28630;
  wire n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638;
  wire n28639, n28640, n28641, n28642, n28645, n28646, n28647, n28648;
  wire n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656;
  wire n28657, n28658, n28659, n28660, n28661, n28664, n28665, n28666;
  wire n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674;
  wire n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682;
  wire n28683, n28688, n28706, n28707, n28708, n28709, n28710, n28711;
  wire n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28721;
  wire n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729;
  wire n28730, n28731, n28732, n28735, n28736, n28737, n28738, n28739;
  wire n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747;
  wire n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757;
  wire n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765;
  wire n28766, n28769, n28770, n28771, n28772, n28773, n28774, n28775;
  wire n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783;
  wire n28784, n28785, n28788, n28789, n28790, n28791, n28792, n28793;
  wire n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801;
  wire n28802, n28803, n28804, n28807, n28808, n28809, n28810, n28811;
  wire n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819;
  wire n28820, n28821, n28822, n28823, n28826, n28827, n28828, n28829;
  wire n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837;
  wire n28838, n28839, n28840, n28841, n28842, n28845, n28846, n28847;
  wire n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855;
  wire n28856, n28857, n28858, n28859, n28860, n28861, n28864, n28865;
  wire n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873;
  wire n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28883;
  wire n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891;
  wire n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899;
  wire n28900, n28901, n28902, n28919, n28920, n28921, n28922, n28923;
  wire n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931;
  wire n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941;
  wire n28942, n28943, n28944, n28945, n28948, n28949, n28950, n28951;
  wire n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959;
  wire n28960, n28963, n28964, n28965, n28966, n28967, n28968, n28969;
  wire n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977;
  wire n28978, n28979, n28982, n28983, n28984, n28985, n28986, n28987;
  wire n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995;
  wire n28996, n28997, n28998, n29001, n29002, n29003, n29004, n29005;
  wire n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013;
  wire n29014, n29015, n29016, n29017, n29020, n29021, n29022, n29023;
  wire n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031;
  wire n29032, n29033, n29034, n29035, n29036, n29039, n29040, n29041;
  wire n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049;
  wire n29050, n29051, n29052, n29053, n29054, n29055, n29058, n29059;
  wire n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067;
  wire n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29077;
  wire n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085;
  wire n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093;
  wire n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101;
  wire n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109;
  wire n29110, n29111, n29112, n29113, n29115, n29116, n29117, n29132;
  wire n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140;
  wire n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148;
  wire n29149, n29150, n29151, n29154, n29155, n29156, n29157, n29158;
  wire n29159, n29160, n29161, n29162, n29163, n29166, n29167, n29168;
  wire n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176;
  wire n29177, n29178, n29181, n29182, n29183, n29184, n29185, n29186;
  wire n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194;
  wire n29195, n29196, n29197, n29200, n29201, n29202, n29203, n29204;
  wire n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212;
  wire n29213, n29214, n29215, n29216, n29219, n29220, n29221, n29222;
  wire n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230;
  wire n29231, n29232, n29233, n29234, n29235, n29238, n29239, n29240;
  wire n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248;
  wire n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29258;
  wire n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266;
  wire n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29276;
  wire n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284;
  wire n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292;
  wire n29293, n29296, n29297, n29298, n29299, n29300, n29301, n29302;
  wire n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310;
  wire n29311, n29312, n29313, n29314, n29315, n29316, n29318, n29319;
  wire n29320, n29321, n29322, n29325, n29337, n29355, n29356, n29357;
  wire n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365;
  wire n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373;
  wire n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381;
  wire n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389;
  wire n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399;
  wire n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407;
  wire n29408, n29411, n29412, n29413, n29414, n29415, n29416, n29417;
  wire n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425;
  wire n29426, n29427, n29430, n29431, n29432, n29433, n29434, n29435;
  wire n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443;
  wire n29444, n29445, n29446, n29449, n29450, n29451, n29452, n29453;
  wire n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461;
  wire n29462, n29463, n29464, n29465, n29468, n29469, n29470, n29471;
  wire n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479;
  wire n29480, n29481, n29482, n29483, n29484, n29485, n29488, n29489;
  wire n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497;
  wire n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29507;
  wire n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515;
  wire n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523;
  wire n29524, n29525, n29526, n29527, n29529, n29530, n29538, n29550;
  wire n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571;
  wire n29572, n29573, n29574, n29575, n29576, n29579, n29580, n29581;
  wire n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589;
  wire n29590, n29593, n29594, n29595, n29596, n29597, n29598, n29599;
  wire n29600, n29601, n29602, n29603, n29604, n29605, n29608, n29609;
  wire n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617;
  wire n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29627;
  wire n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635;
  wire n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643;
  wire n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653;
  wire n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661;
  wire n29662, n29665, n29666, n29667, n29668, n29669, n29670, n29671;
  wire n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679;
  wire n29680, n29681, n29684, n29685, n29686, n29687, n29688, n29689;
  wire n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697;
  wire n29698, n29699, n29700, n29703, n29704, n29705, n29706, n29707;
  wire n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715;
  wire n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723;
  wire n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731;
  wire n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739;
  wire n29741, n29742, n29743, n29744, n29745, n29746, n29749, n29750;
  wire n29751, n29752, n29753, n29767, n29768, n29769, n29770, n29771;
  wire n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779;
  wire n29780, n29781, n29782, n29783, n29786, n29787, n29788, n29789;
  wire n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797;
  wire n29798, n29799, n29800, n29801, n29802, n29805, n29806, n29807;
  wire n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815;
  wire n29816, n29817, n29818, n29819, n29820, n29821, n29824, n29825;
  wire n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833;
  wire n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29843;
  wire n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851;
  wire n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859;
  wire n29860, n29863, n29864, n29865, n29866, n29867, n29868, n29869;
  wire n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877;
  wire n29878, n29881, n29882, n29883, n29884, n29885, n29886, n29887;
  wire n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895;
  wire n29896, n29897, n29898, n29901, n29902, n29903, n29904, n29905;
  wire n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913;
  wire n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921;
  wire n29923, n29924, n29925, n29926, n29927, n29930, n29931, n29946;
  wire n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954;
  wire n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962;
  wire n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970;
  wire n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29980;
  wire n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988;
  wire n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996;
  wire n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006;
  wire n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014;
  wire n30015, n30018, n30019, n30020, n30021, n30022, n30023, n30024;
  wire n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032;
  wire n30033, n30034, n30037, n30038, n30039, n30040, n30041, n30042;
  wire n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050;
  wire n30051, n30052, n30053, n30054, n30057, n30058, n30059, n30060;
  wire n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068;
  wire n30069, n30070, n30071, n30072, n30073, n30076, n30077, n30078;
  wire n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086;
  wire n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094;
  wire n30095, n30096, n30098, n30099, n30117, n30118, n30119, n30120;
  wire n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128;
  wire n30129, n30132, n30133, n30134, n30135, n30136, n30137, n30138;
  wire n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146;
  wire n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154;
  wire n30155, n30156, n30159, n30160, n30161, n30162, n30163, n30164;
  wire n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172;
  wire n30173, n30174, n30175, n30178, n30179, n30180, n30181, n30182;
  wire n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190;
  wire n30191, n30192, n30193, n30194, n30197, n30198, n30199, n30200;
  wire n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208;
  wire n30209, n30210, n30211, n30212, n30213, n30216, n30217, n30218;
  wire n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226;
  wire n30227, n30228, n30229, n30230, n30231, n30232, n30235, n30236;
  wire n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244;
  wire n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252;
  wire n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260;
  wire n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268;
  wire n30269, n30270, n30271, n30272, n30274, n30275, n30276, n30277;
  wire n30278, n30279, n30280, n30283, n30284, n30285, n30286, n30287;
  wire n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310;
  wire n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318;
  wire n30319, n30320, n30321, n30322, n30323, n30324, n30327, n30328;
  wire n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336;
  wire n30337, n30338, n30339, n30342, n30343, n30344, n30345, n30346;
  wire n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354;
  wire n30355, n30356, n30357, n30358, n30361, n30362, n30363, n30364;
  wire n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372;
  wire n30373, n30374, n30375, n30376, n30377, n30378, n30381, n30382;
  wire n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390;
  wire n30391, n30392, n30393, n30394, n30395, n30396, n30399, n30400;
  wire n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408;
  wire n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416;
  wire n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426;
  wire n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434;
  wire n30435, n30436, n30437, n30438, n30439, n30441, n30442, n30443;
  wire n30444, n30445, n30448, n30449, n30464, n30465, n30466, n30467;
  wire n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475;
  wire n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483;
  wire n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491;
  wire n30492, n30493, n30494, n30495, n30498, n30499, n30500, n30501;
  wire n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509;
  wire n30510, n30511, n30512, n30513, n30514, n30517, n30518, n30519;
  wire n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527;
  wire n30528, n30529, n30530, n30531, n30532, n30533, n30536, n30537;
  wire n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545;
  wire n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553;
  wire n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563;
  wire n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571;
  wire n30572, n30575, n30576, n30577, n30578, n30579, n30580, n30581;
  wire n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589;
  wire n30590, n30591, n30592, n30593, n30594, n30595, n30597, n30598;
  wire n30599, n30600, n30601, n30604, n30621, n30622, n30623, n30624;
  wire n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632;
  wire n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640;
  wire n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650;
  wire n30651, n30652, n30653, n30654, n30655, n30658, n30659, n30660;
  wire n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668;
  wire n30669, n30670, n30671, n30672, n30673, n30674, n30677, n30678;
  wire n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686;
  wire n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30696;
  wire n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704;
  wire n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712;
  wire n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722;
  wire n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730;
  wire n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738;
  wire n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746;
  wire n30747, n30748, n30749, n30750, n30751, n30753, n30754, n30755;
  wire n30756, n30757, n30758, n30761, n30762, n30763, n30764, n30765;
  wire n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784;
  wire n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792;
  wire n30793, n30796, n30797, n30798, n30799, n30800, n30801, n30802;
  wire n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810;
  wire n30811, n30812, n30815, n30816, n30817, n30818, n30819, n30820;
  wire n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828;
  wire n30829, n30830, n30831, n30832, n30835, n30836, n30837, n30838;
  wire n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846;
  wire n30847, n30848, n30849, n30850, n30853, n30854, n30855, n30856;
  wire n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864;
  wire n30865, n30866, n30867, n30868, n30869, n30870, n30873, n30874;
  wire n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882;
  wire n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890;
  wire n30891, n30892, n30893, n30895, n30896, n30897, n30898, n30899;
  wire n30902, n30903, n30919, n30920, n30921, n30922, n30923, n30924;
  wire n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932;
  wire n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940;
  wire n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948;
  wire n30949, n30950, n30953, n30954, n30955, n30956, n30957, n30958;
  wire n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966;
  wire n30967, n30968, n30969, n30972, n30973, n30974, n30975, n30976;
  wire n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984;
  wire n30985, n30986, n30987, n30988, n30989, n30992, n30993, n30994;
  wire n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002;
  wire n31003, n31004, n31005, n31006, n31007, n31008, n31011, n31012;
  wire n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020;
  wire n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028;
  wire n31029, n31030, n31031, n31033, n31034, n31035, n31036, n31052;
  wire n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060;
  wire n31061, n31062, n31063, n31064, n31067, n31068, n31069, n31070;
  wire n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078;
  wire n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086;
  wire n31087, n31088, n31089, n31090, n31091, n31094, n31095, n31096;
  wire n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104;
  wire n31105, n31106, n31107, n31108, n31109, n31110, n31113, n31114;
  wire n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122;
  wire n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31132;
  wire n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140;
  wire n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148;
  wire n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156;
  wire n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164;
  wire n31165, n31166, n31167, n31168, n31169, n31171, n31172, n31173;
  wire n31174, n31175, n31176, n31177, n31180, n31181, n31182, n31183;
  wire n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191;
  wire n31192, n31193, n31194, n31197, n31198, n31199, n31200, n31201;
  wire n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221;
  wire n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229;
  wire n31230, n31231, n31232, n31233, n31234, n31235, n31238, n31239;
  wire n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247;
  wire n31248, n31249, n31250, n31251, n31252, n31253, n31256, n31257;
  wire n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265;
  wire n31266, n31267, n31268, n31269, n31270, n31271, n31274, n31275;
  wire n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283;
  wire n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291;
  wire n31292, n31293, n31294, n31296, n31297, n31298, n31299, n31300;
  wire n31303, n31304, n31319, n31320, n31321, n31322, n31323, n31324;
  wire n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332;
  wire n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340;
  wire n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348;
  wire n31349, n31350, n31353, n31354, n31355, n31356, n31357, n31358;
  wire n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366;
  wire n31367, n31368, n31369, n31370, n31371, n31374, n31375, n31376;
  wire n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384;
  wire n31385, n31386, n31387, n31388, n31389, n31390, n31393, n31394;
  wire n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402;
  wire n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410;
  wire n31411, n31412, n31413, n31415, n31416, n31417, n31418, n31419;
  wire n31422, n31435, n31436, n31437, n31438, n31439, n31440, n31441;
  wire n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449;
  wire n31450, n31451, n31452, n31453, n31454, n31457, n31458, n31459;
  wire n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467;
  wire n31468, n31469, n31472, n31473, n31474, n31475, n31476, n31477;
  wire n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485;
  wire n31486, n31487, n31488, n31491, n31492, n31493, n31494, n31495;
  wire n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503;
  wire n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511;
  wire n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519;
  wire n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527;
  wire n31529, n31530, n31531, n31532, n31533, n31534, n31537, n31538;
  wire n31539, n31540, n31541, n31558, n31559, n31560, n31561, n31562;
  wire n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570;
  wire n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578;
  wire n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588;
  wire n31589, n31590, n31591, n31592, n31593, n31596, n31597, n31598;
  wire n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606;
  wire n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31616;
  wire n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624;
  wire n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632;
  wire n31633, n31634, n31635, n31636, n31638, n31639, n31640, n31641;
  wire n31642, n31645, n31646, n31661, n31662, n31663, n31664, n31665;
  wire n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673;
  wire n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681;
  wire n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689;
  wire n31690, n31691, n31692, n31695, n31696, n31697, n31698, n31699;
  wire n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707;
  wire n31708, n31709, n31710, n31711, n31714, n31715, n31716, n31717;
  wire n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725;
  wire n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733;
  wire n31734, n31736, n31751, n31752, n31753, n31754, n31755, n31756;
  wire n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31766;
  wire n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774;
  wire n31775, n31776, n31777, n31780, n31781, n31782, n31783, n31784;
  wire n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792;
  wire n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802;
  wire n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810;
  wire n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818;
  wire n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826;
  wire n31827, n31828, n31829, n31830, n31831, n31832, n31834, n31835;
  wire n31836, n31837, n31838, n31839, n31842, n31843, n31844, n31845;
  wire n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853;
  wire n31854, n31855, n31858, n31859, n31860, n31861, n31862, n31876;
  wire n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884;
  wire n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892;
  wire n31893, n31894, n31895, n31896, n31899, n31900, n31901, n31902;
  wire n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910;
  wire n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918;
  wire n31919, n31921, n31922, n31923, n31924, n31925, n31928, n31929;
  wire n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952;
  wire n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960;
  wire n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968;
  wire n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976;
  wire n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986;
  wire n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994;
  wire n31995, n31996, n31997, n31998, n31999, n32000, n32002, n32003;
  wire n32004, n32005, n32012, n32013, n32014, n32015, n32016, n32017;
  wire n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32027;
  wire n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035;
  wire n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043;
  wire n32044, n32045, n32046, n32047, n32050, n32051, n32052, n32053;
  wire n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061;
  wire n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069;
  wire n32070, n32072, n32073, n32074, n32075, n32078, n32079, n32080;
  wire n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088;
  wire n32089, n32090, n32093, n32094, n32095, n32096, n32097, n32098;
  wire n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106;
  wire n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114;
  wire n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122;
  wire n32123, n_3, n_4, n_5, n_6, n_9, n_10, n_11;
  wire n_12, n_13, n_15, n_17, n_18, n_19, n_21, n_24;
  wire n_25, n_27, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
  wire n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340;
  wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
  wire n_349, n_350, n_351, n_352, n_353, n_354, n_355, n_356;
  wire n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364;
  wire n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_373, n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  wire n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_430, n_431, n_432;
  wire n_433, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_452, n_453;
  wire n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
  wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_596;
  wire n_597, n_599, n_600, n_601, n_602, n_603, n_604, n_605;
  wire n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613;
  wire n_614, n_615, n_617, n_618, n_619, n_620, n_621, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_652, n_653, n_654, n_655;
  wire n_656, n_661, n_662, n_663, n_664, n_665, n_666, n_667;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_692, n_693, n_694, n_695, n_699, n_700, n_702, n_703;
  wire n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711;
  wire n_712, n_713, n_714, n_715, n_716, n_717, n_719, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_764, n_765;
  wire n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781;
  wire n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789;
  wire n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813;
  wire n_814, n_815, n_816, n_821, n_822, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837;
  wire n_838, n_839, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_863, n_864, n_865, n_866, n_867, n_868, n_869;
  wire n_870, n_871, n_872, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929;
  wire n_930, n_935, n_936, n_937, n_938, n_939, n_940, n_941;
  wire n_942, n_947, n_948, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969;
  wire n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981;
  wire n_982, n_983, n_984, n_985, n_986, n_987, n_992, n_993;
  wire n_994, n_995, n_996, n_997, n_999, n_1001, n_1002, n_1003;
  wire n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011;
  wire n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019;
  wire n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1037, n_1038, n_1039;
  wire n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047;
  wire n_1048, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059;
  wire n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067;
  wire n_1068, n_1069, n_1071, n_1072, n_1073, n_1074, n_1075, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088;
  wire n_1089, n_1090, n_1091, n_1092, n_1093, n_1098, n_1099, n_1100;
  wire n_1101, n_1102, n_1103, n_1104, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121;
  wire n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129;
  wire n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137;
  wire n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1157;
  wire n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165;
  wire n_1166, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177;
  wire n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185;
  wire n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193;
  wire n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201;
  wire n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209;
  wire n_1210, n_1211, n_1212, n_1213, n_1214, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1253, n_1254, n_1255, n_1256, n_1257;
  wire n_1258, n_1259, n_1260, n_1261, n_1262, n_1267, n_1268, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1297;
  wire n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305;
  wire n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1317;
  wire n_1318, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329;
  wire n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1359, n_1360, n_1361;
  wire n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1390, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1397, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411;
  wire n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419;
  wire n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427;
  wire n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435;
  wire n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443;
  wire n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467;
  wire n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487;
  wire n_1488, n_1489, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1539;
  wire n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567;
  wire n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575;
  wire n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583;
  wire n_1584, n_1585, n_1586, n_1587, n_1592, n_1593, n_1594, n_1595;
  wire n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603;
  wire n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1627;
  wire n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635;
  wire n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647;
  wire n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683;
  wire n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691;
  wire n_1692, n_1693, n_1694, n_1699, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1705, n_1706, n_1707, n_1708, n_1713, n_1714, n_1715;
  wire n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723;
  wire n_1724, n_1725, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1744, n_1745, n_1746, n_1747;
  wire n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755;
  wire n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763;
  wire n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771;
  wire n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779;
  wire n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787;
  wire n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795;
  wire n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803;
  wire n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1834, n_1835;
  wire n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843;
  wire n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855;
  wire n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1867;
  wire n_1868, n_1869, n_1870, n_1871, n_1872, n_1874, n_1875, n_1876;
  wire n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885;
  wire n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893;
  wire n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901;
  wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1913;
  wire n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921;
  wire n_1922, n_1923, n_1924, n_1925, n_1926, n_1931, n_1932, n_1933;
  wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1953;
  wire n_1954, n_1955, n_1956, n_1957, n_1958, n_1963, n_1964, n_1965;
  wire n_1966, n_1967, n_1968, n_1973, n_1974, n_1975, n_1976, n_1981;
  wire n_1982, n_1983, n_1984, n_1989, n_1990, n_1991, n_1992, n_1997;
  wire n_1998, n_1999, n_2000, n_2001, n_2006, n_2007, n_2008, n_2009;
  wire n_2010, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021;
  wire n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029;
  wire n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037;
  wire n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045;
  wire n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053;
  wire n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061;
  wire n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069;
  wire n_2070, n_2071, n_2072, n_2073, n_2074, n_2079, n_2080, n_2081;
  wire n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089;
  wire n_2090, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101;
  wire n_2102, n_2103, n_2104, n_2109, n_2110, n_2111, n_2112, n_2113;
  wire n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121;
  wire n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133;
  wire n_2134, n_2135, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145;
  wire n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153;
  wire n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161;
  wire n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177;
  wire n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185;
  wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
  wire n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201;
  wire n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209;
  wire n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2220, n_2221;
  wire n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229;
  wire n_2230, n_2231, n_2232, n_2233, n_2238, n_2239, n_2240, n_2241;
  wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2252, n_2253;
  wire n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261;
  wire n_2262, n_2263, n_2264, n_2265, n_2266, n_2271, n_2272, n_2273;
  wire n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2285;
  wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
  wire n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301;
  wire n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309;
  wire n_2310, n_2311, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321;
  wire n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329;
  wire n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341;
  wire n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349;
  wire n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357;
  wire n_2358, n_2359, n_2360, n_2365, n_2366, n_2367, n_2368, n_2369;
  wire n_2370, n_2371, n_2372, n_2373, n_2374, n_2379, n_2380, n_2381;
  wire n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389;
  wire n_2390, n_2391, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401;
  wire n_2402, n_2403, n_2404, n_2405, n_2410, n_2411, n_2412, n_2413;
  wire n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421;
  wire n_2422, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2434;
  wire n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443;
  wire n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451;
  wire n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459;
  wire n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467;
  wire n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475;
  wire n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483;
  wire n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491;
  wire n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499;
  wire n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507;
  wire n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515;
  wire n_2516, n_2517, n_2518, n_2523, n_2524, n_2525, n_2526, n_2527;
  wire n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2538, n_2539;
  wire n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547;
  wire n_2548, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559;
  wire n_2560, n_2561, n_2562, n_2563, n_2568, n_2569, n_2570, n_2571;
  wire n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2583;
  wire n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591;
  wire n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599;
  wire n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607;
  wire n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615;
  wire n_2616, n_2617, n_2618, n_2623, n_2624, n_2625, n_2626, n_2627;
  wire n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635;
  wire n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643;
  wire n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
  wire n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659;
  wire n_2660, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671;
  wire n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2682, n_2683;
  wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
  wire n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703;
  wire n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2715;
  wire n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723;
  wire n_2724, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735;
  wire n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743;
  wire n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751;
  wire n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759;
  wire n_2760, n_2761, n_2762, n_2763, n_2764, n_2769, n_2770, n_2771;
  wire n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779;
  wire n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787;
  wire n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795;
  wire n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803;
  wire n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811;
  wire n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819;
  wire n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827;
  wire n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835;
  wire n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843;
  wire n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851;
  wire n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2863;
  wire n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871;
  wire n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883;
  wire n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891;
  wire n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899;
  wire n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907;
  wire n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915;
  wire n_2916, n_2917, n_2918, n_2923, n_2924, n_2925, n_2926, n_2927;
  wire n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935;
  wire n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943;
  wire n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951;
  wire n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959;
  wire n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967;
  wire n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975;
  wire n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983;
  wire n_2984, n_2985, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995;
  wire n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3007;
  wire n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015;
  wire n_3016, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027;
  wire n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3038, n_3039;
  wire n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047;
  wire n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059;
  wire n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067;
  wire n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075;
  wire n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083;
  wire n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091;
  wire n_3092, n_3093, n_3094, n_3099, n_3100, n_3101, n_3102, n_3103;
  wire n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3114, n_3115;
  wire n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123;
  wire n_3124, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135;
  wire n_3136, n_3137, n_3138, n_3139, n_3144, n_3145, n_3146, n_3147;
  wire n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, n_3159;
  wire n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167;
  wire n_3168, n_3169, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179;
  wire n_3180, n_3181, n_3182, n_3183, n_3184, n_3189, n_3190, n_3191;
  wire n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199;
  wire n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207;
  wire n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215;
  wire n_3216, n_3217, n_3218, n_3219, n_3224, n_3225, n_3226, n_3227;
  wire n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235;
  wire n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243;
  wire n_3244, n_3245, n_3246, n_3251, n_3252, n_3253, n_3254, n_3255;
  wire n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263;
  wire n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271;
  wire n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279;
  wire n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287;
  wire n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3298, n_3299;
  wire n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307;
  wire n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315;
  wire n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323;
  wire n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330, n_3331;
  wire n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, n_3339;
  wire n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347;
  wire n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3359;
  wire n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367;
  wire n_3368, n_3369, n_3370, n_3371, n_3376, n_3377, n_3378, n_3379;
  wire n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3390, n_3391;
  wire n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399;
  wire n_3400, n_3401, n_3402, n_3403, n_3404, n_3409, n_3410, n_3411;
  wire n_3412, n_3413, n_3414, n_3416, n_3418, n_3419, n_3420, n_3421;
  wire n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429;
  wire n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437;
  wire n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445;
  wire n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453;
  wire n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461;
  wire n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469;
  wire n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477;
  wire n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485;
  wire n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493;
  wire n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501;
  wire n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509;
  wire n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517;
  wire n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3528, n_3529;
  wire n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537;
  wire n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549;
  wire n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557;
  wire n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565;
  wire n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573;
  wire n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581;
  wire n_3582, n_3583, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593;
  wire n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609;
  wire n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621;
  wire n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629;
  wire n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637;
  wire n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645;
  wire n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653;
  wire n_3654, n_3655, n_3656, n_3661, n_3662, n_3663, n_3664, n_3665;
  wire n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673;
  wire n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681;
  wire n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689;
  wire n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697;
  wire n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705;
  wire n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713;
  wire n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721;
  wire n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729;
  wire n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737;
  wire n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745;
  wire n_3746, n_3747, n_3748, n_3749, n_3750, n_3755, n_3756, n_3757;
  wire n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765;
  wire n_3766, n_3767, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777;
  wire n_3778, n_3779, n_3780, n_3781, n_3786, n_3787, n_3788, n_3789;
  wire n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797;
  wire n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805;
  wire n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813;
  wire n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3821;
  wire n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829;
  wire n_3830, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841;
  wire n_3842, n_3843, n_3844, n_3845, n_3850, n_3851, n_3852, n_3853;
  wire n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3865;
  wire n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873;
  wire n_3874, n_3875, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885;
  wire n_3886, n_3887, n_3888, n_3889, n_3890, n_3895, n_3896, n_3897;
  wire n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905;
  wire n_3910, n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917;
  wire n_3918, n_3919, n_3920, n_3925, n_3926, n_3927, n_3928, n_3929;
  wire n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937;
  wire n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945;
  wire n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953;
  wire n_3954, n_3955, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965;
  wire n_3966, n_3967, n_3968, n_3969, n_3974, n_3975, n_3976, n_3977;
  wire n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3989;
  wire n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997;
  wire n_3998, n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005;
  wire n_4006, n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013;
  wire n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021;
  wire n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029;
  wire n_4030, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041;
  wire n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049;
  wire n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4061;
  wire n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069;
  wire n_4070, n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077;
  wire n_4078, n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085;
  wire n_4086, n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093;
  wire n_4094, n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101;
  wire n_4102, n_4103, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113;
  wire n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121;
  wire n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129;
  wire n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137;
  wire n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145;
  wire n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153;
  wire n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161;
  wire n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169;
  wire n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177;
  wire n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185;
  wire n_4186, n_4187, n_4188, n_4189, n_4190, n_4195, n_4196, n_4197;
  wire n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205;
  wire n_4206, n_4207, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217;
  wire n_4218, n_4219, n_4220, n_4221, n_4226, n_4227, n_4228, n_4229;
  wire n_4230, n_4231, n_4232, n_4233, n_4234, n_4235, n_4236, n_4237;
  wire n_4238, n_4239, n_4240, n_4241, n_4242, n_4243, n_4244, n_4245;
  wire n_4246, n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253;
  wire n_4254, n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261;
  wire n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4268, n_4269;
  wire n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277;
  wire n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284, n_4285;
  wire n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293;
  wire n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301;
  wire n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309;
  wire n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317;
  wire n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325;
  wire n_4330, n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337;
  wire n_4338, n_4339, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349;
  wire n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357;
  wire n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365;
  wire n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373;
  wire n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381;
  wire n_4382, n_4383, n_4384, n_4389, n_4390, n_4391, n_4392, n_4393;
  wire n_4394, n_4395, n_4396, n_4397, n_4398, n_4403, n_4404, n_4405;
  wire n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413;
  wire n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425;
  wire n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433;
  wire n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440, n_4441;
  wire n_4442, n_4443, n_4444, n_4445, n_4446, n_4447, n_4448, n_4449;
  wire n_4450, n_4451, n_4452, n_4453, n_4454, n_4455, n_4456, n_4457;
  wire n_4458, n_4459, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469;
  wire n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477;
  wire n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485;
  wire n_4490, n_4491, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497;
  wire n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505;
  wire n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513;
  wire n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521;
  wire n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529;
  wire n_4530, n_4531, n_4532, n_4537, n_4538, n_4539, n_4540, n_4541;
  wire n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549;
  wire n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557;
  wire n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565;
  wire n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573;
  wire n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581;
  wire n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589;
  wire n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597;
  wire n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605;
  wire n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613;
  wire n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621;
  wire n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629;
  wire n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637;
  wire n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645;
  wire n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4657;
  wire n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665;
  wire n_4666, n_4667, n_4668, n_4669, n_4674, n_4675, n_4676, n_4677;
  wire n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685;
  wire n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693;
  wire n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701;
  wire n_4702, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713;
  wire n_4714, n_4715, n_4716, n_4717, n_4722, n_4723, n_4724, n_4725;
  wire n_4726, n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4737;
  wire n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745;
  wire n_4746, n_4747, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757;
  wire n_4758, n_4759, n_4760, n_4761, n_4762, n_4767, n_4768, n_4769;
  wire n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4776, n_4777;
  wire n_4782, n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789;
  wire n_4790, n_4791, n_4792, n_4797, n_4798, n_4799, n_4800, n_4801;
  wire n_4802, n_4803, n_4804, n_4805, n_4806, n_4807, n_4808, n_4809;
  wire n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4816, n_4817;
  wire n_4818, n_4819, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825;
  wire n_4826, n_4827, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837;
  wire n_4838, n_4839, n_4840, n_4841, n_4846, n_4847, n_4848, n_4849;
  wire n_4850, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4861;
  wire n_4862, n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869;
  wire n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877;
  wire n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885;
  wire n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893;
  wire n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901;
  wire n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913;
  wire n_4914, n_4915, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925;
  wire n_4926, n_4927, n_4928, n_4929, n_4930, n_4935, n_4936, n_4937;
  wire n_4938, n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945;
  wire n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953;
  wire n_4954, n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961;
  wire n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969;
  wire n_4970, n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4981;
  wire n_4982, n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989;
  wire n_4990, n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997;
  wire n_4998, n_4999, n_5000, n_5001, n_5002, n_5007, n_5008, n_5009;
  wire n_5010, n_5011, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017;
  wire n_5018, n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025;
  wire n_5026, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032, n_5033;
  wire n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040, n_5041;
  wire n_5042, n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049;
  wire n_5054, n_5055, n_5056, n_5057, n_5058, n_5059, n_5060, n_5061;
  wire n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068, n_5069;
  wire n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076, n_5077;
  wire n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084, n_5085;
  wire n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092, n_5093;
  wire n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100, n_5101;
  wire n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108, n_5109;
  wire n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116, n_5117;
  wire n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124, n_5125;
  wire n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132, n_5133;
  wire n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140, n_5141;
  wire n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148, n_5149;
  wire n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156, n_5157;
  wire n_5158, n_5159, n_5160, n_5161, n_5162, n_5167, n_5168, n_5169;
  wire n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176, n_5177;
  wire n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185;
  wire n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193;
  wire n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5201;
  wire n_5202, n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5209;
  wire n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5216, n_5217;
  wire n_5218, n_5219, n_5220, n_5221, n_5222, n_5223, n_5224, n_5225;
  wire n_5226, n_5227, n_5228, n_5229, n_5230, n_5231, n_5232, n_5233;
  wire n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240, n_5241;
  wire n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248, n_5249;
  wire n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256, n_5257;
  wire n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264, n_5265;
  wire n_5266, n_5271, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277;
  wire n_5278, n_5279, n_5280, n_5285, n_5286, n_5287, n_5288, n_5289;
  wire n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296, n_5297;
  wire n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304, n_5305;
  wire n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313;
  wire n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320, n_5321;
  wire n_5322, n_5323, n_5324, n_5325, n_5330, n_5331, n_5332, n_5333;
  wire n_5334, n_5335, n_5336, n_5337, n_5338, n_5339, n_5344, n_5345;
  wire n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353;
  wire n_5354, n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365;
  wire n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373;
  wire n_5374, n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381;
  wire n_5382, n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389;
  wire n_5390, n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397;
  wire n_5398, n_5399, n_5404, n_5405, n_5406, n_5407, n_5408, n_5409;
  wire n_5410, n_5411, n_5412, n_5413, n_5418, n_5419, n_5420, n_5421;
  wire n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5433;
  wire n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440, n_5441;
  wire n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448, n_5449;
  wire n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456, n_5457;
  wire n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464, n_5465;
  wire n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472, n_5473;
  wire n_5474, n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485;
  wire n_5486, n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493;
  wire n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5505;
  wire n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512, n_5513;
  wire n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520, n_5521;
  wire n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528, n_5529;
  wire n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537;
  wire n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544, n_5545;
  wire n_5546, n_5547, n_5552, n_5553, n_5554, n_5555, n_5556, n_5557;
  wire n_5558, n_5559, n_5560, n_5561, n_5562, n_5563, n_5564, n_5565;
  wire n_5566, n_5567, n_5568, n_5569, n_5570, n_5571, n_5572, n_5573;
  wire n_5574, n_5575, n_5576, n_5577, n_5578, n_5579, n_5580, n_5581;
  wire n_5582, n_5583, n_5584, n_5585, n_5586, n_5587, n_5588, n_5589;
  wire n_5590, n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597;
  wire n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605;
  wire n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613;
  wire n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621;
  wire n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629;
  wire n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637;
  wire n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645;
  wire n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653;
  wire n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661;
  wire n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669;
  wire n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677;
  wire n_5678, n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685;
  wire n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5697;
  wire n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704, n_5705;
  wire n_5706, n_5707, n_5708, n_5709, n_5711, n_5712, n_5713, n_5715;
  wire n_5716, n_5717, n_5718, n_5719, n_5720, n_5721, n_5722, n_5727;
  wire n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735;
  wire n_5736, n_5737, n_5738, n_5739, n_5740, n_5741, n_5742, n_5743;
  wire n_5744, n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755;
  wire n_5756, n_5757, n_5758, n_5759, n_5764, n_5765, n_5766, n_5767;
  wire n_5768, n_5769, n_5770, n_5771, n_5772, n_5773, n_5774, n_5779;
  wire n_5780, n_5781, n_5782, n_5783, n_5784, n_5785, n_5786, n_5787;
  wire n_5788, n_5789, n_5794, n_5795, n_5796, n_5797, n_5798, n_5799;
  wire n_5800, n_5801, n_5802, n_5803, n_5804, n_5809, n_5810, n_5811;
  wire n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819;
  wire n_5824, n_5825, n_5826, n_5827, n_5828, n_5829, n_5830, n_5831;
  wire n_5832, n_5833, n_5834, n_5835, n_5836, n_5837, n_5838, n_5839;
  wire n_5840, n_5841, n_5842, n_5843, n_5844, n_5845, n_5846, n_5847;
  wire n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854, n_5859;
  wire n_5860, n_5861, n_5862, n_5863, n_5864, n_5865, n_5866, n_5867;
  wire n_5868, n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879;
  wire n_5880, n_5881, n_5882, n_5883, n_5888, n_5889, n_5890, n_5891;
  wire n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898, n_5899;
  wire n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907;
  wire n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915;
  wire n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923;
  wire n_5924, n_5925, n_5926, n_5927, n_5928, n_5933, n_5934, n_5935;
  wire n_5936, n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5947;
  wire n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955;
  wire n_5956, n_5957, n_5962, n_5963, n_5964, n_5965, n_5966, n_5967;
  wire n_5968, n_5969, n_5970, n_5971, n_5972, n_5973, n_5974, n_5975;
  wire n_5976, n_5977, n_5978, n_5979, n_5980, n_5981, n_5982, n_5983;
  wire n_5984, n_5985, n_5986, n_5987, n_5988, n_5989, n_5990, n_5991;
  wire n_5992, n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999;
  wire n_6000, n_6001, n_6002, n_6007, n_6008, n_6009, n_6010, n_6011;
  wire n_6012, n_6013, n_6014, n_6015, n_6016, n_6021, n_6022, n_6023;
  wire n_6024, n_6025, n_6026, n_6027, n_6028, n_6029, n_6030, n_6031;
  wire n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043;
  wire n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051;
  wire n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059;
  wire n_6060, n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067;
  wire n_6068, n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075;
  wire n_6076, n_6077, n_6082, n_6083, n_6084, n_6085, n_6086, n_6087;
  wire n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094, n_6095;
  wire n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103;
  wire n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115;
  wire n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123;
  wire n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131;
  wire n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139;
  wire n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147;
  wire n_6148, n_6149, n_6150, n_6155, n_6156, n_6157, n_6158, n_6159;
  wire n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166, n_6167;
  wire n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6174, n_6175;
  wire n_6176, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183;
  wire n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191;
  wire n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199;
  wire n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207;
  wire n_6208, n_6209, n_6210, n_6211, n_6212, n_6213, n_6214, n_6215;
  wire n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223;
  wire n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231;
  wire n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239;
  wire n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247;
  wire n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255;
  wire n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263;
  wire n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271;
  wire n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279;
  wire n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287;
  wire n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295;
  wire n_6296, n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303;
  wire n_6304, n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311;
  wire n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319;
  wire n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327;
  wire n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335;
  wire n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343;
  wire n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351;
  wire n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6365;
  wire n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376, n_6377;
  wire n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384, n_6385;
  wire n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392, n_6393;
  wire n_6398, n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405;
  wire n_6406, n_6407, n_6408, n_6409, n_6410, n_6411, n_6412, n_6413;
  wire n_6414, n_6415, n_6416, n_6417, n_6418, n_6419, n_6420, n_6425;
  wire n_6426, n_6427, n_6428, n_6429, n_6430, n_6431, n_6432, n_6433;
  wire n_6434, n_6435, n_6436, n_6437, n_6438, n_6439, n_6440, n_6441;
  wire n_6442, n_6443, n_6444, n_6445, n_6446, n_6447, n_6448, n_6449;
  wire n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457;
  wire n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, n_6465;
  wire n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472, n_6473;
  wire n_6474, n_6475, n_6476, n_6477, n_6482, n_6483, n_6484, n_6485;
  wire n_6486, n_6487, n_6488, n_6489, n_6490, n_6491, n_6496, n_6497;
  wire n_6498, n_6499, n_6500, n_6501, n_6502, n_6503, n_6504, n_6509;
  wire n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516, n_6517;
  wire n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524, n_6525;
  wire n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532, n_6533;
  wire n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540, n_6541;
  wire n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548, n_6549;
  wire n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556, n_6557;
  wire n_6558, n_6559, n_6560, n_6565, n_6566, n_6567, n_6568, n_6569;
  wire n_6570, n_6571, n_6572, n_6573, n_6574, n_6579, n_6580, n_6581;
  wire n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6592, n_6593;
  wire n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601;
  wire n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608, n_6609;
  wire n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617;
  wire n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6625;
  wire n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633;
  wire n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641;
  wire n_6642, n_6643, n_6648, n_6649, n_6650, n_6651, n_6652, n_6653;
  wire n_6654, n_6655, n_6656, n_6657, n_6662, n_6663, n_6664, n_6665;
  wire n_6666, n_6667, n_6668, n_6669, n_6670, n_6675, n_6676, n_6677;
  wire n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684, n_6685;
  wire n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692, n_6693;
  wire n_6694, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700, n_6701;
  wire n_6702, n_6703, n_6704, n_6705, n_6706, n_6707, n_6708, n_6709;
  wire n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716, n_6717;
  wire n_6718, n_6719, n_6720, n_6721, n_6722, n_6723, n_6724, n_6725;
  wire n_6726, n_6731, n_6732, n_6733, n_6734, n_6735, n_6736, n_6737;
  wire n_6738, n_6739, n_6744, n_6745, n_6746, n_6747, n_6748, n_6749;
  wire n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757;
  wire n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764, n_6765;
  wire n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772, n_6773;
  wire n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780, n_6781;
  wire n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788, n_6789;
  wire n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796, n_6797;
  wire n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804, n_6805;
  wire n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812, n_6813;
  wire n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820, n_6821;
  wire n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828, n_6829;
  wire n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836, n_6837;
  wire n_6838, n_6839, n_6840, n_6841, n_6842, n_6843, n_6844, n_6845;
  wire n_6846, n_6847, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853;
  wire n_6854, n_6855, n_6856, n_6857, n_6858, n_6859, n_6860, n_6861;
  wire n_6862, n_6863, n_6868, n_6869, n_6870, n_6871, n_6872, n_6873;
  wire n_6874, n_6875, n_6876, n_6877, n_6882, n_6883, n_6884, n_6885;
  wire n_6886, n_6887, n_6888, n_6889, n_6890, n_6891, n_6892, n_6893;
  wire n_6894, n_6895, n_6896, n_6897, n_6898, n_6899, n_6900, n_6901;
  wire n_6902, n_6903, n_6904, n_6905, n_6906, n_6907, n_6908, n_6909;
  wire n_6910, n_6911, n_6912, n_6913, n_6914, n_6915, n_6916, n_6917;
  wire n_6918, n_6919, n_6920, n_6921, n_6922, n_6923, n_6924, n_6925;
  wire n_6926, n_6927, n_6928, n_6929, n_6930, n_6931, n_6932, n_6933;
  wire n_6934, n_6935, n_6936, n_6937, n_6938, n_6939, n_6940, n_6941;
  wire n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948, n_6949;
  wire n_6950, n_6951, n_6952, n_6953, n_6954, n_6955, n_6956, n_6957;
  wire n_6958, n_6959, n_6960, n_6961, n_6962, n_6963, n_6964, n_6965;
  wire n_6966, n_6967, n_6968, n_6969, n_6970, n_6971, n_6972, n_6973;
  wire n_6974, n_6975, n_6976, n_6977, n_6978, n_6979, n_6980, n_6981;
  wire n_6982, n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6989;
  wire n_6990, n_6991, n_6992, n_6993, n_6994, n_6995, n_6996, n_6997;
  wire n_6998, n_6999, n_7000, n_7001, n_7002, n_7003, n_7004, n_7005;
  wire n_7006, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012, n_7013;
  wire n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020, n_7021;
  wire n_7022, n_7023, n_7024, n_7025, n_7026, n_7027, n_7028, n_7029;
  wire n_7030, n_7031, n_7032, n_7033, n_7034, n_7035, n_7036, n_7037;
  wire n_7038, n_7039, n_7040, n_7041, n_7042, n_7043, n_7044, n_7045;
  wire n_7046, n_7047, n_7048, n_7049, n_7050, n_7051, n_7052, n_7053;
  wire n_7054, n_7055, n_7056, n_7057, n_7058, n_7059, n_7060, n_7061;
  wire n_7062, n_7063, n_7064, n_7065, n_7066, n_7067, n_7068, n_7069;
  wire n_7070, n_7071, n_7072, n_7073, n_7074, n_7075, n_7076, n_7077;
  wire n_7078, n_7079, n_7080, n_7081, n_7082, n_7083, n_7084, n_7085;
  wire n_7086, n_7087, n_7088, n_7089, n_7090, n_7091, n_7092, n_7093;
  wire n_7094, n_7095, n_7096, n_7097, n_7098, n_7099, n_7100, n_7101;
  wire n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108, n_7109;
  wire n_7110, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120, n_7121;
  wire n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129;
  wire n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136, n_7137;
  wire n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145;
  wire n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153;
  wire n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7164, n_7165;
  wire n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172, n_7173;
  wire n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181;
  wire n_7182, n_7183, n_7184, n_7189, n_7190, n_7191, n_7192, n_7193;
  wire n_7194, n_7195, n_7196, n_7197, n_7198, n_7199, n_7200, n_7201;
  wire n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208, n_7209;
  wire n_7210, n_7211, n_7212, n_7213, n_7214, n_7215, n_7216, n_7221;
  wire n_7222, n_7223, n_7224, n_7229, n_7230, n_7231, n_7232, n_7233;
  wire n_7234, n_7235, n_7236, n_7237, n_7238, n_7239, n_7240, n_7241;
  wire n_7242, n_7243, n_7244, n_7245, n_7246, n_7247, n_7248, n_7249;
  wire n_7250, n_7251, n_7252, n_7253, n_7254, n_7255, n_7256, n_7257;
  wire n_7258, n_7259, n_7260, n_7261, n_7262, n_7263, n_7264, n_7265;
  wire n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273;
  wire n_7274, n_7275, n_7276, n_7277, n_7278, n_7283, n_7284, n_7285;
  wire n_7286, n_7287, n_7288, n_7289, n_7290, n_7291, n_7292, n_7297;
  wire n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304, n_7305;
  wire n_7306, n_7307, n_7308, n_7309, n_7310, n_7315, n_7316, n_7317;
  wire n_7318, n_7319, n_7320, n_7321, n_7322, n_7323, n_7324, n_7325;
  wire n_7326, n_7327, n_7328, n_7329, n_7330, n_7331, n_7332, n_7333;
  wire n_7338, n_7339, n_7340, n_7341, n_7342, n_7343, n_7344, n_7345;
  wire n_7346, n_7347, n_7348, n_7349, n_7350, n_7351, n_7352, n_7353;
  wire n_7354, n_7355, n_7356, n_7357, n_7358, n_7359, n_7360, n_7361;
  wire n_7362, n_7363, n_7364, n_7365, n_7366, n_7367, n_7372, n_7373;
  wire n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, n_7380, n_7381;
  wire n_7382, n_7383, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389;
  wire n_7390, n_7391, n_7392, n_7393, n_7394, n_7395, n_7396, n_7397;
  wire n_7398, n_7399, n_7400, n_7401, n_7402, n_7403, n_7404, n_7405;
  wire n_7406, n_7407, n_7408, n_7409, n_7410, n_7411, n_7412, n_7413;
  wire n_7414, n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7421;
  wire n_7422, n_7423, n_7424, n_7425, n_7426, n_7427, n_7428, n_7429;
  wire n_7430, n_7431, n_7432, n_7433, n_7434, n_7435, n_7436, n_7437;
  wire n_7438, n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445;
  wire n_7446, n_7447, n_7452, n_7453, n_7454, n_7455, n_7456, n_7457;
  wire n_7458, n_7459, n_7460, n_7461, n_7462, n_7463, n_7464, n_7465;
  wire n_7466, n_7467, n_7468, n_7469, n_7470, n_7471, n_7472, n_7473;
  wire n_7474, n_7475, n_7476, n_7477, n_7478, n_7479, n_7480, n_7481;
  wire n_7482, n_7483, n_7484, n_7485, n_7486, n_7487, n_7488, n_7489;
  wire n_7490, n_7491, n_7492, n_7493, n_7494, n_7495, n_7496, n_7497;
  wire n_7498, n_7499, n_7500, n_7501, n_7502, n_7507, n_7508, n_7509;
  wire n_7510, n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517;
  wire n_7518, n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525;
  wire n_7526, n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533;
  wire n_7534, n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541;
  wire n_7542, n_7543, n_7547, n_7548, n_7549, n_7550, n_7551, n_7552;
  wire n_7553, n_7554, n_7555, n_7556, n_7557, n_7558, n_7559, n_7560;
  wire n_7561, n_7562, n_7563, n_7565, n_7566, n_7567, n_7568, n_7569;
  wire n_7570, n_7571, n_7572, n_7573, n_7574, n_7575, n_7576, n_7577;
  wire n_7578, n_7579, n_7580, n_7581, n_7582, n_7583, n_7584, n_7585;
  wire n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7592, n_7593;
  wire n_7594, n_7599, n_7600, n_7601, n_7602, n_7603, n_7604, n_7605;
  wire n_7606, n_7607, n_7612, n_7613, n_7614, n_7615, n_7616, n_7617;
  wire n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625;
  wire n_7626, n_7627, n_7628, n_7629, n_7630, n_7631, n_7632, n_7633;
  wire n_7638, n_7639, n_7640, n_7641, n_7642, n_7643, n_7644, n_7645;
  wire n_7646, n_7647, n_7648, n_7649, n_7650, n_7651, n_7652, n_7653;
  wire n_7654, n_7655, n_7656, n_7657, n_7658, n_7659, n_7660, n_7661;
  wire n_7662, n_7663, n_7664, n_7665, n_7666, n_7667, n_7668, n_7669;
  wire n_7670, n_7671, n_7675, n_7676, n_7677, n_7679, n_7680, n_7681;
  wire n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688, n_7689;
  wire n_7690, n_7694, n_7695, n_7697, n_7698, n_7699, n_7700, n_7701;
  wire n_7702, n_7703, n_7704, n_7705, n_7706, n_7707, n_7708, n_7709;
  wire n_7710, n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717;
  wire n_7718, n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725;
  wire n_7726, n_7727, n_7728, n_7729, n_7730, n_7731, n_7732, n_7736;
  wire n_7737, n_7739, n_7740, n_7741, n_7742, n_7743, n_7744, n_7745;
  wire n_7746, n_7747, n_7748, n_7749, n_7754, n_7755, n_7756, n_7757;
  wire n_7758, n_7759, n_7760, n_7761, n_7765, n_7767, n_7768, n_7769;
  wire n_7770, n_7771, n_7772, n_7773, n_7774, n_7775, n_7776, n_7777;
  wire n_7778, n_7779, n_7780, n_7784, n_7786, n_7787, n_7788, n_7789;
  wire n_7790, n_7791, n_7792, n_7793, n_7794, n_7795, n_7796, n_7797;
  wire n_7798, n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7809;
  wire n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816, n_7817;
  wire n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824, n_7825;
  wire n_7826, n_7827, n_7828, n_7829, n_7830, n_7831, n_7832, n_7837;
  wire n_7838, n_7839, n_7840, n_7841, n_7842, n_7843, n_7844, n_7845;
  wire n_7846, n_7847, n_7848, n_7849, n_7854, n_7855, n_7856, n_7857;
  wire n_7858, n_7859, n_7860, n_7861, n_7862, n_7863, n_7868, n_7869;
  wire n_7870, n_7871, n_7872, n_7873, n_7877, n_7878, n_7880, n_7881;
  wire n_7882, n_7883, n_7884, n_7885, n_7886, n_7887, n_7888, n_7889;
  wire n_7890, n_7891, n_7892, n_7893, n_7894, n_7895, n_7896, n_7897;
  wire n_7898, n_7899, n_7900, n_7905, n_7906, n_7907, n_7908, n_7909;
  wire n_7910, n_7911, n_7912, n_7913, n_7914, n_7915, n_7920, n_7921;
  wire n_7922, n_7923, n_7928, n_7929, n_7930, n_7931, n_7932, n_7933;
  wire n_7934, n_7935, n_7936, n_7937, n_7938, n_7939, n_7940, n_7941;
  wire n_7942, n_7943, n_7944, n_7945, n_7946, n_7947, n_7948, n_7949;
  wire n_7950, n_7951, n_7952, n_7953, n_7954, n_7955, n_7956, n_7957;
  wire n_7958, n_7959, n_7960, n_7961, n_7966, n_7967, n_7968, n_7969;
  wire n_7970, n_7971, n_7972, n_7973, n_7974, n_7975, n_7976, n_7977;
  wire n_7978, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988, n_7989;
  wire n_7990, n_7991, n_7992, n_7993, n_7994, n_7995, n_7996, n_7997;
  wire n_7998, n_7999, n_8000, n_8001, n_8002, n_8003, n_8004, n_8005;
  wire n_8006, n_8007, n_8008, n_8009, n_8010, n_8011, n_8012, n_8017;
  wire n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025;
  wire n_8026, n_8027, n_8028, n_8033, n_8034, n_8035, n_8036, n_8037;
  wire n_8038, n_8039, n_8040, n_8041, n_8042, n_8043, n_8044, n_8045;
  wire n_8046, n_8047, n_8048, n_8049, n_8050, n_8051, n_8052, n_8053;
  wire n_8054, n_8055, n_8056, n_8057, n_8058, n_8059, n_8060, n_8061;
  wire n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072, n_8073;
  wire n_8078, n_8079, n_8080, n_8081, n_8082, n_8083, n_8084, n_8085;
  wire n_8086, n_8087, n_8088, n_8089, n_8090, n_8091, n_8092, n_8093;
  wire n_8094, n_8095, n_8096, n_8097, n_8098, n_8099, n_8100, n_8101;
  wire n_8102, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112, n_8113;
  wire n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120, n_8121;
  wire n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128, n_8129;
  wire n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136, n_8137;
  wire n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8148, n_8149;
  wire n_8150, n_8151, n_8152, n_8153, n_8154, n_8155, n_8156, n_8157;
  wire n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168, n_8169;
  wire n_8170, n_8171, n_8172, n_8173, n_8174, n_8179, n_8180, n_8181;
  wire n_8182, n_8183, n_8184, n_8185, n_8186, n_8187, n_8188, n_8189;
  wire n_8190, n_8191, n_8192, n_8193, n_8194, n_8195, n_8200, n_8201;
  wire n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208, n_8209;
  wire n_8214, n_8215, n_8216, n_8217, n_8218, n_8219, n_8220, n_8221;
  wire n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232, n_8233;
  wire n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8244, n_8245;
  wire n_8246, n_8247, n_8248, n_8249, n_8250, n_8251, n_8252, n_8253;
  wire n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8268, n_8269;
  wire n_8270, n_8271, n_8272, n_8273, n_8274, n_8275, n_8276, n_8277;
  wire n_8278, n_8279, n_8280, n_8281, n_8282, n_8283, n_8284, n_8285;
  wire n_8286, n_8287, n_8292, n_8293, n_8294, n_8295, n_8296, n_8297;
  wire n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304, n_8305;
  wire n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316, n_8317;
  wire n_8318, n_8319, n_8320, n_8321, n_8322, n_8323, n_8324, n_8325;
  wire n_8326, n_8327, n_8328, n_8329, n_8330, n_8331, n_8332, n_8337;
  wire n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345;
  wire n_8346, n_8347, n_8348, n_8349, n_8354, n_8355, n_8356, n_8357;
  wire n_8358, n_8359, n_8360, n_8361, n_8362, n_8363, n_8368, n_8369;
  wire n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376, n_8377;
  wire n_8378, n_8379, n_8380, n_8385, n_8386, n_8387, n_8388, n_8389;
  wire n_8390, n_8391, n_8392, n_8393, n_8394, n_8395, n_8396, n_8397;
  wire n_8398, n_8399, n_8400, n_8401, n_8402, n_8403, n_8404, n_8405;
  wire n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412, n_8413;
  wire n_8414, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424, n_8425;
  wire n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432, n_8437;
  wire n_8438, n_8439, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445;
  wire n_8446, n_8447, n_8448, n_8453, n_8454, n_8455, n_8456, n_8457;
  wire n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464, n_8465;
  wire n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472, n_8473;
  wire n_8474, n_8475, n_8476, n_8477, n_8482, n_8483, n_8484, n_8485;
  wire n_8486, n_8487, n_8488, n_8489, n_8490, n_8491, n_8492, n_8493;
  wire n_8494, n_8495, n_8496, n_8497, n_8498, n_8499, n_8500, n_8501;
  wire n_8502, n_8503, n_8504, n_8505, n_8506, n_8507, n_8508, n_8509;
  wire n_8510, n_8511, n_8512, n_8513, n_8514, n_8515, n_8516, n_8517;
  wire n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528, n_8529;
  wire n_8530, n_8531, n_8532, n_8533, n_8534, n_8539, n_8540, n_8541;
  wire n_8542, n_8543, n_8544, n_8545, n_8546, n_8547, n_8548, n_8553;
  wire n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560, n_8561;
  wire n_8562, n_8563, n_8564, n_8565, n_8570, n_8571, n_8572, n_8573;
  wire n_8574, n_8575, n_8576, n_8577, n_8578, n_8579, n_8580, n_8581;
  wire n_8582, n_8583, n_8584, n_8585, n_8586, n_8591, n_8592, n_8593;
  wire n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600, n_8601;
  wire n_8602, n_8607, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613;
  wire n_8614, n_8615, n_8616, n_8617, n_8618, n_8619, n_8624, n_8625;
  wire n_8626, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632, n_8633;
  wire n_8634, n_8639, n_8640, n_8641, n_8642, n_8643, n_8644, n_8645;
  wire n_8646, n_8647, n_8648, n_8649, n_8650, n_8651, n_8652, n_8653;
  wire n_8654, n_8655, n_8656, n_8657, n_8658, n_8659, n_8664, n_8665;
  wire n_8666, n_8667, n_8668, n_8669, n_8670, n_8671, n_8672, n_8673;
  wire n_8674, n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681;
  wire n_8682, n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689;
  wire n_8690, n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8701;
  wire n_8702, n_8703, n_8704, n_8705, n_8706, n_8707, n_8708, n_8709;
  wire n_8710, n_8715, n_8716, n_8717, n_8718, n_8719, n_8720, n_8721;
  wire n_8722, n_8723, n_8724, n_8725, n_8726, n_8727, n_8732, n_8733;
  wire n_8734, n_8735, n_8736, n_8737, n_8738, n_8739, n_8740, n_8741;
  wire n_8746, n_8747, n_8748, n_8749, n_8750, n_8751, n_8756, n_8757;
  wire n_8758, n_8759, n_8760, n_8761, n_8762, n_8763, n_8764, n_8765;
  wire n_8766, n_8767, n_8768, n_8769, n_8770, n_8771, n_8772, n_8773;
  wire n_8774, n_8775, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785;
  wire n_8786, n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8797;
  wire n_8798, n_8799, n_8800, n_8801, n_8802, n_8803, n_8804, n_8805;
  wire n_8810, n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817;
  wire n_8822, n_8823, n_8824, n_8825, n_8826, n_8827, n_8828, n_8829;
  wire n_8830, n_8831, n_8832, n_8833, n_8834, n_8835, n_8840, n_8841;
  wire n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8848, n_8849;
  wire n_8854, n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861;
  wire n_8862, n_8863, n_8864, n_8865, n_8866, n_8871, n_8872, n_8873;
  wire n_8874, n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881;
  wire n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889;
  wire n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897;
  wire n_8898, n_8899, n_8900, n_8905, n_8906, n_8907, n_8908, n_8909;
  wire n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916, n_8917;
  wire n_8922, n_8923, n_8924, n_8925, n_8926, n_8927, n_8928, n_8929;
  wire n_8930, n_8931, n_8932, n_8933, n_8934, n_8935, n_8936, n_8941;
  wire n_8942, n_8943, n_8944, n_8945, n_8946, n_8947, n_8948, n_8949;
  wire n_8954, n_8955, n_8956, n_8957, n_8958, n_8959, n_8960, n_8961;
  wire n_8962, n_8967, n_8968, n_8969, n_8970, n_8971, n_8976, n_8977;
  wire n_8978, n_8979, n_8980, n_8985, n_8986, n_8987, n_8988, n_8993;
  wire n_8994, n_8995, n_8996, n_8997, n_9002, n_9003, n_9004, n_9005;
  wire n_9006, n_9011, n_9012, n_9013, n_9014, n_9019, n_9020, n_9021;
  wire n_9022, n_9027, n_9028, n_9029, n_9030, n_9031, n_9032, n_9033;
  wire n_9034, n_9035, n_9036, n_9037, n_9038, n_9039, n_9040, n_9041;
  wire n_9046, n_9047, n_9048, n_9049, n_9050, n_9051, n_9052, n_9053;
  wire n_9054, n_9055, n_9056, n_9057, n_9058, n_9059, n_9060, n_9061;
  wire n_9062, n_9063, n_9064, n_9065, n_9066, n_9067, n_9068, n_9069;
  wire n_9070, n_9071, n_9072, n_9073, n_9074, n_9075, n_9076, n_9077;
  wire n_9078, n_9079, n_9080, n_9081, n_9082, n_9083, n_9084, n_9085;
  wire n_9086, n_9087, n_9088, n_9089, n_9090, n_9091, n_9092, n_9093;
  wire n_9094, n_9095, n_9096, n_9097, n_9098, n_9099, n_9100, n_9101;
  wire n_9102, n_9103, n_9104, n_9105, n_9106, n_9107, n_9108, n_9109;
  wire n_9110, n_9111, n_9112, n_9113, n_9114, n_9115, n_9116, n_9117;
  wire n_9118, n_9119, n_9120, n_9121, n_9122, n_9123, n_9128, n_9129;
  wire n_9130, n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137;
  wire n_9138, n_9139, n_9144, n_9145, n_9146, n_9147, n_9148, n_9149;
  wire n_9150, n_9151, n_9152, n_9153, n_9158, n_9159, n_9160, n_9161;
  wire n_9162, n_9163, n_9164, n_9165, n_9166, n_9167, n_9168, n_9169;
  wire n_9170, n_9175, n_9176, n_9177, n_9178, n_9179, n_9180, n_9181;
  wire n_9182, n_9183, n_9184, n_9189, n_9190, n_9191, n_9192, n_9193;
  wire n_9194, n_9195, n_9196, n_9197, n_9198, n_9199, n_9200, n_9201;
  wire n_9206, n_9207, n_9208, n_9209, n_9210, n_9211, n_9212, n_9213;
  wire n_9214, n_9215, n_9216, n_9217, n_9218, n_9219, n_9220, n_9221;
  wire n_9222, n_9227, n_9228, n_9229, n_9230, n_9231, n_9232, n_9233;
  wire n_9234, n_9235, n_9236, n_9237, n_9238, n_9239, n_9240, n_9245;
  wire n_9246, n_9247, n_9248, n_9249, n_9250, n_9251, n_9252, n_9253;
  wire n_9254, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265;
  wire n_9266, n_9271, n_9272, n_9273, n_9274, n_9275, n_9276, n_9277;
  wire n_9278, n_9279, n_9280, n_9281, n_9282, n_9283, n_9284, n_9289;
  wire n_9290, n_9291, n_9292, n_9293, n_9294, n_9295, n_9296, n_9297;
  wire n_9298, n_9303, n_9304, n_9305, n_9306, n_9307, n_9308, n_9309;
  wire n_9310, n_9311, n_9312, n_9313, n_9314, n_9315, n_9320, n_9321;
  wire n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9328, n_9329;
  wire n_9334, n_9335, n_9336, n_9337, n_9338, n_9339, n_9344, n_9345;
  wire n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353;
  wire n_9354, n_9355, n_9356, n_9357, n_9358, n_9359, n_9360, n_9361;
  wire n_9362, n_9363, n_9368, n_9369, n_9370, n_9371, n_9372, n_9373;
  wire n_9374, n_9375, n_9376, n_9377, n_9378, n_9379, n_9380, n_9385;
  wire n_9386, n_9387, n_9388, n_9389, n_9390, n_9391, n_9392, n_9393;
  wire n_9394, n_9395, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405;
  wire n_9406, n_9407, n_9412, n_9413, n_9414, n_9415, n_9416, n_9417;
  wire n_9418, n_9419, n_9420, n_9421, n_9422, n_9427, n_9428, n_9429;
  wire n_9430, n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437;
  wire n_9438, n_9439, n_9444, n_9445, n_9446, n_9447, n_9448, n_9449;
  wire n_9450, n_9451, n_9452, n_9453, n_9458, n_9459, n_9460, n_9461;
  wire n_9462, n_9463, n_9464, n_9465, n_9466, n_9467, n_9468, n_9469;
  wire n_9470, n_9475, n_9476, n_9477, n_9478, n_9479, n_9480, n_9481;
  wire n_9482, n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489;
  wire n_9490, n_9491, n_9492, n_9493, n_9494, n_9495, n_9496, n_9497;
  wire n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9504, n_9509;
  wire n_9510, n_9511, n_9512, n_9513, n_9514, n_9515, n_9516, n_9517;
  wire n_9518, n_9519, n_9520, n_9521, n_9526, n_9527, n_9528, n_9529;
  wire n_9530, n_9531, n_9532, n_9533, n_9534, n_9535, n_9536, n_9537;
  wire n_9538, n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545;
  wire n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552, n_9553;
  wire n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9560, n_9561;
  wire n_9562, n_9563, n_9564, n_9565, n_9566, n_9567, n_9568, n_9569;
  wire n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576, n_9577;
  wire n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584, n_9585;
  wire n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592, n_9593;
  wire n_9594, n_9595, n_9596, n_9597, n_9598, n_9599, n_9604, n_9605;
  wire n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612, n_9613;
  wire n_9614, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624, n_9625;
  wire n_9626, n_9627, n_9628, n_9629, n_9634, n_9635, n_9636, n_9637;
  wire n_9638, n_9639, n_9640, n_9641, n_9642, n_9643, n_9644, n_9649;
  wire n_9650, n_9651, n_9652, n_9653, n_9654, n_9655, n_9656, n_9657;
  wire n_9658, n_9659, n_9664, n_9665, n_9666, n_9667, n_9668, n_9669;
  wire n_9670, n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677;
  wire n_9678, n_9679, n_9680, n_9681, n_9682, n_9683, n_9684, n_9685;
  wire n_9686, n_9687, n_9688, n_9689, n_9690, n_9691, n_9692, n_9697;
  wire n_9698, n_9699, n_9700, n_9701, n_9702, n_9703, n_9704, n_9705;
  wire n_9706, n_9707, n_9708, n_9709, n_9710, n_9711, n_9712, n_9713;
  wire n_9714, n_9715, n_9716, n_9717, n_9718, n_9719, n_9720, n_9721;
  wire n_9722, n_9723, n_9724, n_9725, n_9726, n_9727, n_9728, n_9729;
  wire n_9730, n_9731, n_9732, n_9733, n_9734, n_9735, n_9736, n_9737;
  wire n_9738, n_9739, n_9740, n_9741, n_9742, n_9743, n_9744, n_9745;
  wire n_9746, n_9747, n_9748, n_9749, n_9754, n_9755, n_9756, n_9757;
  wire n_9758, n_9759, n_9760, n_9761, n_9762, n_9763, n_9768, n_9769;
  wire n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776, n_9777;
  wire n_9782, n_9783, n_9784, n_9785, n_9786, n_9787, n_9788, n_9789;
  wire n_9790, n_9791, n_9792, n_9793, n_9794, n_9799, n_9800, n_9801;
  wire n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808, n_9813;
  wire n_9814, n_9815, n_9816, n_9817, n_9818, n_9819, n_9820, n_9821;
  wire n_9822, n_9823, n_9824, n_9825, n_9830, n_9831, n_9832, n_9833;
  wire n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841;
  wire n_9842, n_9843, n_9844, n_9845, n_9846, n_9851, n_9852, n_9853;
  wire n_9854, n_9855, n_9856, n_9857, n_9858, n_9859, n_9860, n_9861;
  wire n_9862, n_9863, n_9864, n_9865, n_9866, n_9867, n_9868, n_9869;
  wire n_9870, n_9871, n_9872, n_9873, n_9874, n_9875, n_9876, n_9877;
  wire n_9878, n_9879, n_9880, n_9881, n_9882, n_9883, n_9884, n_9885;
  wire n_9886, n_9887, n_9888, n_9889, n_9890, n_9891, n_9892, n_9893;
  wire n_9894, n_9895, n_9896, n_9897, n_9898, n_9899, n_9900, n_9901;
  wire n_9902, n_9903, n_9904, n_9905, n_9906, n_9907, n_9908, n_9909;
  wire n_9910, n_9911, n_9912, n_9913, n_9914, n_9915, n_9916, n_9917;
  wire n_9918, n_9919, n_9920, n_9921, n_9922, n_9923, n_9924, n_9925;
  wire n_9926, n_9927, n_9928, n_9929, n_9930, n_9931, n_9932, n_9933;
  wire n_9934, n_9935, n_9936, n_9937, n_9938, n_9939, n_9940, n_9941;
  wire n_9942, n_9943, n_9944, n_9945, n_9946, n_9947, n_9948, n_9949;
  wire n_9950, n_9951, n_9952, n_9953, n_9954, n_9955, n_9956, n_9957;
  wire n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964, n_9965;
  wire n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972, n_9973;
  wire n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984, n_9985;
  wire n_9986, n_9991, n_9992, n_9993, n_9994, n_9995, n_9996, n_9997;
  wire n_9998, n_9999, n_10000, n_10001, n_10002, n_10003, n_10004,
       n_10005;
  wire n_10006, n_10007, n_10008, n_10009, n_10010, n_10011, n_10012,
       n_10013;
  wire n_10014, n_10015, n_10016, n_10017, n_10018, n_10019, n_10020,
       n_10021;
  wire n_10022, n_10023, n_10024, n_10025, n_10026, n_10027, n_10028,
       n_10029;
  wire n_10030, n_10031, n_10032, n_10033, n_10038, n_10039, n_10040,
       n_10041;
  wire n_10042, n_10043, n_10044, n_10045, n_10046, n_10047, n_10048,
       n_10049;
  wire n_10050, n_10051, n_10052, n_10053, n_10054, n_10055, n_10056,
       n_10057;
  wire n_10058, n_10059, n_10060, n_10061, n_10062, n_10063, n_10064,
       n_10065;
  wire n_10066, n_10067, n_10068, n_10069, n_10070, n_10071, n_10072,
       n_10073;
  wire n_10074, n_10075, n_10076, n_10077, n_10078, n_10079, n_10080,
       n_10081;
  wire n_10082, n_10083, n_10084, n_10085, n_10086, n_10087, n_10088,
       n_10089;
  wire n_10090, n_10091, n_10092, n_10093, n_10094, n_10095, n_10096,
       n_10097;
  wire n_10098, n_10099, n_10100, n_10101, n_10102, n_10103, n_10104,
       n_10105;
  wire n_10106, n_10107, n_10108, n_10109, n_10110, n_10111, n_10112,
       n_10113;
  wire n_10114, n_10115, n_10116, n_10117, n_10118, n_10123, n_10124,
       n_10125;
  wire n_10126, n_10127, n_10128, n_10129, n_10130, n_10131, n_10132,
       n_10137;
  wire n_10138, n_10139, n_10140, n_10141, n_10142, n_10143, n_10144,
       n_10145;
  wire n_10146, n_10151, n_10152, n_10153, n_10154, n_10155, n_10156,
       n_10157;
  wire n_10158, n_10159, n_10160, n_10161, n_10162, n_10163, n_10168,
       n_10169;
  wire n_10170, n_10171, n_10172, n_10173, n_10174, n_10175, n_10176,
       n_10177;
  wire n_10182, n_10183, n_10184, n_10185, n_10186, n_10187, n_10192,
       n_10193;
  wire n_10194, n_10195, n_10196, n_10197, n_10198, n_10199, n_10200,
       n_10201;
  wire n_10202, n_10203, n_10204, n_10205, n_10206, n_10207, n_10208,
       n_10209;
  wire n_10210, n_10211, n_10216, n_10217, n_10218, n_10219, n_10220,
       n_10221;
  wire n_10222, n_10223, n_10224, n_10225, n_10226, n_10227, n_10228,
       n_10229;
  wire n_10234, n_10235, n_10236, n_10237, n_10238, n_10239, n_10240,
       n_10241;
  wire n_10242, n_10243, n_10248, n_10249, n_10250, n_10251, n_10252,
       n_10253;
  wire n_10254, n_10255, n_10256, n_10257, n_10258, n_10263, n_10264,
       n_10265;
  wire n_10266, n_10267, n_10268, n_10269, n_10270, n_10271, n_10272,
       n_10273;
  wire n_10278, n_10279, n_10280, n_10281, n_10282, n_10283, n_10284,
       n_10285;
  wire n_10286, n_10287, n_10288, n_10293, n_10294, n_10295, n_10296,
       n_10297;
  wire n_10298, n_10299, n_10300, n_10301, n_10302, n_10303, n_10308,
       n_10309;
  wire n_10310, n_10311, n_10312, n_10313, n_10314, n_10315, n_10316,
       n_10317;
  wire n_10318, n_10323, n_10324, n_10325, n_10326, n_10327, n_10328,
       n_10329;
  wire n_10330, n_10331, n_10332, n_10333, n_10338, n_10339, n_10340,
       n_10341;
  wire n_10342, n_10343, n_10344, n_10345, n_10346, n_10347, n_10348,
       n_10353;
  wire n_10354, n_10355, n_10356, n_10357, n_10358, n_10359, n_10360,
       n_10361;
  wire n_10362, n_10363, n_10368, n_10369, n_10370, n_10371, n_10372,
       n_10373;
  wire n_10374, n_10375, n_10376, n_10377, n_10378, n_10379, n_10380,
       n_10381;
  wire n_10382, n_10383, n_10384, n_10385, n_10386, n_10387, n_10388,
       n_10389;
  wire n_10390, n_10391, n_10392, n_10393, n_10394, n_10395, n_10396,
       n_10397;
  wire n_10398, n_10403, n_10404, n_10405, n_10406, n_10407, n_10408,
       n_10409;
  wire n_10410, n_10411, n_10412, n_10413, n_10414, n_10415, n_10416,
       n_10417;
  wire n_10418, n_10419, n_10420, n_10421, n_10422, n_10423, n_10424,
       n_10429;
  wire n_10430, n_10431, n_10432, n_10433, n_10434, n_10435, n_10436,
       n_10437;
  wire n_10438, n_10439, n_10440, n_10441, n_10442, n_10443, n_10444,
       n_10445;
  wire n_10446, n_10447, n_10448, n_10449, n_10450, n_10451, n_10452,
       n_10453;
  wire n_10454, n_10455, n_10456, n_10457, n_10458, n_10459, n_10460,
       n_10461;
  wire n_10462, n_10463, n_10464, n_10465, n_10466, n_10467, n_10468,
       n_10469;
  wire n_10470, n_10471, n_10476, n_10477, n_10478, n_10479, n_10480,
       n_10481;
  wire n_10482, n_10483, n_10484, n_10485, n_10486, n_10487, n_10488,
       n_10489;
  wire n_10490, n_10491, n_10492, n_10493, n_10494, n_10495, n_10496,
       n_10497;
  wire n_10498, n_10499, n_10500, n_10501, n_10502, n_10503, n_10504,
       n_10505;
  wire n_10506, n_10507, n_10508, n_10509, n_10510, n_10511, n_10512,
       n_10513;
  wire n_10514, n_10515, n_10516, n_10517, n_10518, n_10519, n_10520,
       n_10521;
  wire n_10522, n_10523, n_10524, n_10525, n_10526, n_10527, n_10528,
       n_10529;
  wire n_10530, n_10531, n_10532, n_10533, n_10534, n_10535, n_10536,
       n_10537;
  wire n_10538, n_10539, n_10540, n_10541, n_10542, n_10547, n_10548,
       n_10549;
  wire n_10550, n_10551, n_10552, n_10553, n_10554, n_10555, n_10556,
       n_10561;
  wire n_10562, n_10563, n_10564, n_10565, n_10566, n_10567, n_10568,
       n_10569;
  wire n_10570, n_10575, n_10576, n_10577, n_10578, n_10579, n_10580,
       n_10581;
  wire n_10582, n_10583, n_10584, n_10585, n_10586, n_10587, n_10592,
       n_10593;
  wire n_10594, n_10595, n_10596, n_10597, n_10598, n_10599, n_10600,
       n_10601;
  wire n_10602, n_10603, n_10604, n_10605, n_10606, n_10607, n_10608,
       n_10609;
  wire n_10610, n_10611, n_10612, n_10613, n_10614, n_10615, n_10616,
       n_10617;
  wire n_10618, n_10619, n_10620, n_10621, n_10626, n_10627, n_10628,
       n_10629;
  wire n_10630, n_10631, n_10632, n_10633, n_10634, n_10635, n_10636,
       n_10637;
  wire n_10638, n_10639, n_10640, n_10641, n_10642, n_10643, n_10644,
       n_10645;
  wire n_10646, n_10647, n_10648, n_10649, n_10650, n_10651, n_10652,
       n_10653;
  wire n_10654, n_10655, n_10656, n_10657, n_10658, n_10659, n_10660,
       n_10661;
  wire n_10662, n_10663, n_10664, n_10665, n_10666, n_10667, n_10668,
       n_10669;
  wire n_10670, n_10671, n_10672, n_10673, n_10674, n_10675, n_10676,
       n_10677;
  wire n_10678, n_10679, n_10680, n_10681, n_10682, n_10683, n_10684,
       n_10685;
  wire n_10686, n_10687, n_10688, n_10689, n_10690, n_10691, n_10692,
       n_10693;
  wire n_10694, n_10695, n_10696, n_10697, n_10698, n_10699, n_10700,
       n_10701;
  wire n_10702, n_10703, n_10704, n_10705, n_10706, n_10707, n_10708,
       n_10709;
  wire n_10710, n_10711, n_10712, n_10713, n_10714, n_10715, n_10716,
       n_10717;
  wire n_10718, n_10719, n_10720, n_10721, n_10722, n_10723, n_10724,
       n_10725;
  wire n_10726, n_10727, n_10728, n_10729, n_10730, n_10731, n_10732,
       n_10733;
  wire n_10734, n_10735, n_10736, n_10737, n_10738, n_10739, n_10740,
       n_10741;
  wire n_10746, n_10747, n_10748, n_10749, n_10750, n_10751, n_10752,
       n_10753;
  wire n_10754, n_10755, n_10760, n_10761, n_10762, n_10763, n_10764,
       n_10765;
  wire n_10766, n_10767, n_10768, n_10769, n_10770, n_10771, n_10772,
       n_10773;
  wire n_10774, n_10775, n_10776, n_10777, n_10778, n_10779, n_10780,
       n_10781;
  wire n_10782, n_10783, n_10784, n_10785, n_10786, n_10787, n_10788,
       n_10789;
  wire n_10790, n_10791, n_10792, n_10793, n_10794, n_10795, n_10796,
       n_10797;
  wire n_10798, n_10799, n_10800, n_10801, n_10806, n_10807, n_10808,
       n_10809;
  wire n_10810, n_10811, n_10812, n_10813, n_10814, n_10815, n_10816,
       n_10817;
  wire n_10818, n_10819, n_10820, n_10821, n_10822, n_10823, n_10824,
       n_10825;
  wire n_10826, n_10827, n_10832, n_10833, n_10834, n_10835, n_10836,
       n_10837;
  wire n_10838, n_10839, n_10840, n_10841, n_10842, n_10843, n_10844,
       n_10845;
  wire n_10846, n_10847, n_10848, n_10849, n_10850, n_10851, n_10852,
       n_10853;
  wire n_10854, n_10855, n_10856, n_10857, n_10858, n_10859, n_10860,
       n_10861;
  wire n_10862, n_10863, n_10864, n_10865, n_10866, n_10867, n_10868,
       n_10869;
  wire n_10870, n_10871, n_10872, n_10873, n_10874, n_10879, n_10880,
       n_10881;
  wire n_10882, n_10883, n_10884, n_10885, n_10886, n_10887, n_10888,
       n_10889;
  wire n_10890, n_10891, n_10892, n_10893, n_10894, n_10895, n_10896,
       n_10897;
  wire n_10898, n_10899, n_10900, n_10901, n_10902, n_10903, n_10904,
       n_10905;
  wire n_10906, n_10907, n_10908, n_10909, n_10910, n_10911, n_10912,
       n_10913;
  wire n_10914, n_10915, n_10916, n_10917, n_10918, n_10919, n_10920,
       n_10921;
  wire n_10922, n_10923, n_10924, n_10925, n_10926, n_10927, n_10928,
       n_10929;
  wire n_10930, n_10931, n_10932, n_10933, n_10934, n_10935, n_10936,
       n_10937;
  wire n_10938, n_10939, n_10940, n_10941, n_10942, n_10943, n_10944,
       n_10945;
  wire n_10946, n_10947, n_10948, n_10949, n_10950, n_10951, n_10952,
       n_10953;
  wire n_10954, n_10955, n_10956, n_10957, n_10958, n_10959, n_10960,
       n_10961;
  wire n_10962, n_10963, n_10964, n_10965, n_10966, n_10967, n_10968,
       n_10969;
  wire n_10970, n_10971, n_10972, n_10973, n_10974, n_10975, n_10976,
       n_10977;
  wire n_10978, n_10979, n_10980, n_10981, n_10982, n_10983, n_10984,
       n_10985;
  wire n_10986, n_10991, n_10992, n_10993, n_10994, n_10995, n_10996,
       n_10997;
  wire n_10998, n_10999, n_11000, n_11005, n_11006, n_11007, n_11008,
       n_11009;
  wire n_11010, n_11011, n_11012, n_11013, n_11014, n_11019, n_11020,
       n_11021;
  wire n_11022, n_11023, n_11024, n_11025, n_11026, n_11027, n_11028,
       n_11029;
  wire n_11030, n_11031, n_11036, n_11037, n_11038, n_11039, n_11040,
       n_11041;
  wire n_11042, n_11043, n_11044, n_11045, n_11046, n_11047, n_11048,
       n_11049;
  wire n_11050, n_11051, n_11052, n_11053, n_11058, n_11059, n_11060,
       n_11061;
  wire n_11062, n_11063, n_11064, n_11065, n_11066, n_11067, n_11072,
       n_11073;
  wire n_11074, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080,
       n_11081;
  wire n_11082, n_11087, n_11088, n_11089, n_11090, n_11091, n_11092,
       n_11093;
  wire n_11094, n_11095, n_11096, n_11097, n_11102, n_11103, n_11104,
       n_11105;
  wire n_11106, n_11107, n_11108, n_11109, n_11110, n_11111, n_11112,
       n_11117;
  wire n_11118, n_11119, n_11120, n_11121, n_11122, n_11123, n_11124,
       n_11125;
  wire n_11126, n_11127, n_11132, n_11133, n_11134, n_11135, n_11136,
       n_11137;
  wire n_11138, n_11139, n_11140, n_11141, n_11142, n_11147, n_11148,
       n_11149;
  wire n_11150, n_11151, n_11152, n_11153, n_11154, n_11155, n_11156,
       n_11157;
  wire n_11162, n_11163, n_11164, n_11165, n_11166, n_11167, n_11168,
       n_11169;
  wire n_11170, n_11171, n_11172, n_11177, n_11178, n_11179, n_11180,
       n_11181;
  wire n_11182, n_11183, n_11184, n_11185, n_11186, n_11187, n_11192,
       n_11193;
  wire n_11194, n_11195, n_11196, n_11197, n_11198, n_11199, n_11200,
       n_11201;
  wire n_11202, n_11203, n_11204, n_11205, n_11206, n_11207, n_11208,
       n_11209;
  wire n_11210, n_11211, n_11212, n_11213, n_11214, n_11215, n_11216,
       n_11217;
  wire n_11218, n_11219, n_11220, n_11221, n_11222, n_11227, n_11228,
       n_11229;
  wire n_11230, n_11231, n_11232, n_11233, n_11234, n_11235, n_11236,
       n_11241;
  wire n_11242, n_11243, n_11244, n_11245, n_11246, n_11247, n_11248,
       n_11249;
  wire n_11250, n_11251, n_11256, n_11257, n_11258, n_11259, n_11260,
       n_11261;
  wire n_11262, n_11263, n_11264, n_11265, n_11266, n_11267, n_11268,
       n_11269;
  wire n_11270, n_11271, n_11272, n_11273, n_11274, n_11275, n_11276,
       n_11277;
  wire n_11278, n_11279, n_11280, n_11281, n_11282, n_11283, n_11284,
       n_11285;
  wire n_11286, n_11287, n_11288, n_11289, n_11290, n_11291, n_11292,
       n_11293;
  wire n_11294, n_11295, n_11296, n_11297, n_11302, n_11303, n_11304,
       n_11305;
  wire n_11306, n_11307, n_11308, n_11309, n_11310, n_11311, n_11312,
       n_11313;
  wire n_11314, n_11315, n_11316, n_11317, n_11318, n_11319, n_11320,
       n_11321;
  wire n_11322, n_11323, n_11328, n_11329, n_11330, n_11331, n_11332,
       n_11333;
  wire n_11334, n_11335, n_11336, n_11337, n_11338, n_11339, n_11340,
       n_11341;
  wire n_11342, n_11343, n_11344, n_11345, n_11346, n_11347, n_11348,
       n_11349;
  wire n_11350, n_11351, n_11352, n_11353, n_11354, n_11355, n_11356,
       n_11357;
  wire n_11358, n_11359, n_11360, n_11361, n_11362, n_11363, n_11364,
       n_11365;
  wire n_11366, n_11367, n_11368, n_11369, n_11370, n_11375, n_11376,
       n_11377;
  wire n_11378, n_11379, n_11380, n_11381, n_11382, n_11383, n_11384,
       n_11385;
  wire n_11386, n_11387, n_11388, n_11389, n_11390, n_11391, n_11392,
       n_11393;
  wire n_11394, n_11395, n_11396, n_11397, n_11398, n_11399, n_11400,
       n_11401;
  wire n_11402, n_11403, n_11404, n_11405, n_11406, n_11407, n_11408,
       n_11409;
  wire n_11410, n_11411, n_11412, n_11413, n_11414, n_11415, n_11416,
       n_11417;
  wire n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424,
       n_11425;
  wire n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432,
       n_11433;
  wire n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440,
       n_11441;
  wire n_11442, n_11443, n_11444, n_11445, n_11446, n_11447, n_11448,
       n_11449;
  wire n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11456,
       n_11457;
  wire n_11458, n_11459, n_11460, n_11461, n_11462, n_11463, n_11464,
       n_11465;
  wire n_11466, n_11467, n_11472, n_11473, n_11474, n_11475, n_11476,
       n_11477;
  wire n_11478, n_11479, n_11480, n_11481, n_11486, n_11487, n_11488,
       n_11489;
  wire n_11490, n_11491, n_11492, n_11493, n_11494, n_11495, n_11500,
       n_11501;
  wire n_11502, n_11503, n_11504, n_11505, n_11510, n_11511, n_11512,
       n_11513;
  wire n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520,
       n_11521;
  wire n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528,
       n_11529;
  wire n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536,
       n_11537;
  wire n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544,
       n_11545;
  wire n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552,
       n_11553;
  wire n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560,
       n_11561;
  wire n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568,
       n_11569;
  wire n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576,
       n_11577;
  wire n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584,
       n_11585;
  wire n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592,
       n_11593;
  wire n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600,
       n_11601;
  wire n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11608,
       n_11609;
  wire n_11610, n_11611, n_11612, n_11613, n_11614, n_11615, n_11616,
       n_11617;
  wire n_11618, n_11619, n_11620, n_11621, n_11622, n_11623, n_11624,
       n_11625;
  wire n_11626, n_11627, n_11628, n_11629, n_11630, n_11631, n_11636,
       n_11637;
  wire n_11638, n_11639, n_11640, n_11641, n_11642, n_11643, n_11644,
       n_11645;
  wire n_11650, n_11651, n_11652, n_11653, n_11654, n_11655, n_11656,
       n_11657;
  wire n_11658, n_11659, n_11660, n_11661, n_11662, n_11663, n_11664,
       n_11665;
  wire n_11666, n_11667, n_11668, n_11669, n_11670, n_11671, n_11672,
       n_11673;
  wire n_11674, n_11675, n_11676, n_11677, n_11678, n_11679, n_11680,
       n_11681;
  wire n_11682, n_11683, n_11684, n_11685, n_11686, n_11687, n_11688,
       n_11689;
  wire n_11690, n_11695, n_11696, n_11697, n_11698, n_11699, n_11700,
       n_11701;
  wire n_11702, n_11703, n_11704, n_11709, n_11710, n_11711, n_11712,
       n_11713;
  wire n_11714, n_11715, n_11716, n_11717, n_11718, n_11719, n_11724,
       n_11725;
  wire n_11726, n_11727, n_11728, n_11729, n_11730, n_11731, n_11732,
       n_11733;
  wire n_11734, n_11735, n_11736, n_11737, n_11738, n_11739, n_11740,
       n_11741;
  wire n_11742, n_11743, n_11744, n_11745, n_11746, n_11747, n_11748,
       n_11749;
  wire n_11750, n_11751, n_11752, n_11753, n_11754, n_11755, n_11756,
       n_11757;
  wire n_11758, n_11759, n_11760, n_11761, n_11762, n_11763, n_11764,
       n_11765;
  wire n_11770, n_11771, n_11772, n_11773, n_11774, n_11775, n_11776,
       n_11777;
  wire n_11778, n_11779, n_11780, n_11781, n_11782, n_11783, n_11784,
       n_11785;
  wire n_11786, n_11787, n_11788, n_11789, n_11790, n_11791, n_11796,
       n_11797;
  wire n_11798, n_11799, n_11800, n_11801, n_11802, n_11803, n_11804,
       n_11805;
  wire n_11806, n_11807, n_11808, n_11809, n_11810, n_11811, n_11812,
       n_11813;
  wire n_11814, n_11815, n_11816, n_11817, n_11818, n_11819, n_11820,
       n_11821;
  wire n_11822, n_11823, n_11824, n_11825, n_11826, n_11827, n_11828,
       n_11829;
  wire n_11830, n_11831, n_11832, n_11833, n_11834, n_11835, n_11836,
       n_11837;
  wire n_11838, n_11843, n_11844, n_11845, n_11846, n_11847, n_11848,
       n_11849;
  wire n_11850, n_11851, n_11852, n_11853, n_11854, n_11855, n_11856,
       n_11857;
  wire n_11858, n_11859, n_11860, n_11861, n_11862, n_11863, n_11864,
       n_11865;
  wire n_11866, n_11867, n_11868, n_11869, n_11870, n_11871, n_11872,
       n_11873;
  wire n_11874, n_11875, n_11876, n_11877, n_11878, n_11879, n_11880,
       n_11881;
  wire n_11882, n_11883, n_11884, n_11885, n_11886, n_11887, n_11888,
       n_11889;
  wire n_11890, n_11891, n_11892, n_11893, n_11894, n_11895, n_11896,
       n_11897;
  wire n_11898, n_11899, n_11900, n_11901, n_11902, n_11903, n_11904,
       n_11905;
  wire n_11906, n_11907, n_11908, n_11909, n_11910, n_11911, n_11912,
       n_11913;
  wire n_11914, n_11915, n_11916, n_11917, n_11918, n_11919, n_11920,
       n_11921;
  wire n_11922, n_11923, n_11924, n_11925, n_11926, n_11927, n_11928,
       n_11929;
  wire n_11930, n_11931, n_11932, n_11933, n_11934, n_11935, n_11936,
       n_11937;
  wire n_11938, n_11939, n_11940, n_11941, n_11942, n_11943, n_11944,
       n_11945;
  wire n_11946, n_11947, n_11948, n_11949, n_11950, n_11951, n_11952,
       n_11953;
  wire n_11954, n_11955, n_11956, n_11957, n_11958, n_11959, n_11960,
       n_11961;
  wire n_11962, n_11963, n_11964, n_11965, n_11966, n_11967, n_11968,
       n_11969;
  wire n_11970, n_11971, n_11972, n_11973, n_11974, n_11975, n_11976,
       n_11981;
  wire n_11982, n_11983, n_11984, n_11985, n_11986, n_11987, n_11988,
       n_11989;
  wire n_11990, n_11995, n_11996, n_11997, n_11998, n_11999, n_12000,
       n_12001;
  wire n_12002, n_12003, n_12004, n_12005, n_12006, n_12007, n_12008,
       n_12009;
  wire n_12010, n_12011, n_12012, n_12013, n_12014, n_12015, n_12016,
       n_12017;
  wire n_12018, n_12019, n_12020, n_12021, n_12022, n_12023, n_12024,
       n_12025;
  wire n_12030, n_12031, n_12032, n_12033, n_12034, n_12035, n_12036,
       n_12037;
  wire n_12038, n_12039, n_12044, n_12045, n_12046, n_12047, n_12048,
       n_12049;
  wire n_12050, n_12051, n_12052, n_12053, n_12054, n_12059, n_12060,
       n_12061;
  wire n_12062, n_12063, n_12064, n_12065, n_12066, n_12067, n_12068,
       n_12069;
  wire n_12074, n_12075, n_12076, n_12077, n_12078, n_12079, n_12080,
       n_12081;
  wire n_12082, n_12083, n_12084, n_12089, n_12090, n_12091, n_12092,
       n_12093;
  wire n_12094, n_12095, n_12096, n_12097, n_12098, n_12099, n_12104,
       n_12105;
  wire n_12106, n_12107, n_12108, n_12109, n_12110, n_12111, n_12112,
       n_12113;
  wire n_12114, n_12119, n_12120, n_12121, n_12122, n_12123, n_12124,
       n_12125;
  wire n_12126, n_12127, n_12128, n_12129, n_12134, n_12135, n_12136,
       n_12137;
  wire n_12138, n_12139, n_12140, n_12141, n_12142, n_12143, n_12144,
       n_12149;
  wire n_12150, n_12151, n_12152, n_12153, n_12154, n_12155, n_12156,
       n_12157;
  wire n_12158, n_12159, n_12164, n_12165, n_12166, n_12167, n_12168,
       n_12169;
  wire n_12170, n_12171, n_12172, n_12173, n_12174, n_12175, n_12176,
       n_12177;
  wire n_12178, n_12179, n_12180, n_12181, n_12182, n_12183, n_12184,
       n_12185;
  wire n_12186, n_12187, n_12188, n_12189, n_12190, n_12191, n_12192,
       n_12193;
  wire n_12194, n_12199, n_12200, n_12201, n_12202, n_12203, n_12204,
       n_12205;
  wire n_12206, n_12207, n_12208, n_12213, n_12214, n_12215, n_12216,
       n_12217;
  wire n_12218, n_12219, n_12220, n_12221, n_12222, n_12223, n_12228,
       n_12229;
  wire n_12230, n_12231, n_12232, n_12233, n_12234, n_12235, n_12236,
       n_12237;
  wire n_12238, n_12239, n_12240, n_12241, n_12242, n_12243, n_12244,
       n_12245;
  wire n_12246, n_12247, n_12248, n_12249, n_12250, n_12251, n_12252,
       n_12253;
  wire n_12254, n_12255, n_12256, n_12257, n_12258, n_12259, n_12260,
       n_12261;
  wire n_12262, n_12263, n_12264, n_12265, n_12266, n_12267, n_12268,
       n_12273;
  wire n_12274, n_12275, n_12276, n_12277, n_12278, n_12279, n_12280,
       n_12281;
  wire n_12282, n_12287, n_12288, n_12289, n_12290, n_12291, n_12292,
       n_12293;
  wire n_12294, n_12295, n_12296, n_12297, n_12302, n_12303, n_12304,
       n_12305;
  wire n_12306, n_12307, n_12308, n_12309, n_12310, n_12311, n_12312,
       n_12313;
  wire n_12314, n_12315, n_12316, n_12317, n_12318, n_12319, n_12320,
       n_12321;
  wire n_12322, n_12323, n_12324, n_12325, n_12326, n_12327, n_12328,
       n_12329;
  wire n_12330, n_12331, n_12332, n_12333, n_12334, n_12335, n_12336,
       n_12337;
  wire n_12338, n_12339, n_12340, n_12341, n_12342, n_12343, n_12348,
       n_12349;
  wire n_12350, n_12351, n_12352, n_12353, n_12354, n_12355, n_12356,
       n_12357;
  wire n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364,
       n_12365;
  wire n_12366, n_12367, n_12368, n_12369, n_12374, n_12375, n_12376,
       n_12377;
  wire n_12378, n_12379, n_12380, n_12381, n_12382, n_12383, n_12384,
       n_12385;
  wire n_12386, n_12387, n_12388, n_12389, n_12390, n_12391, n_12392,
       n_12393;
  wire n_12394, n_12395, n_12396, n_12397, n_12398, n_12399, n_12400,
       n_12401;
  wire n_12402, n_12403, n_12404, n_12405, n_12406, n_12407, n_12408,
       n_12409;
  wire n_12410, n_12411, n_12412, n_12413, n_12414, n_12415, n_12416,
       n_12421;
  wire n_12422, n_12423, n_12424, n_12425, n_12426, n_12427, n_12428,
       n_12429;
  wire n_12430, n_12431, n_12432, n_12433, n_12434, n_12435, n_12436,
       n_12437;
  wire n_12438, n_12439, n_12440, n_12441, n_12442, n_12443, n_12444,
       n_12445;
  wire n_12446, n_12447, n_12448, n_12449, n_12450, n_12451, n_12452,
       n_12453;
  wire n_12454, n_12455, n_12456, n_12457, n_12458, n_12459, n_12460,
       n_12461;
  wire n_12462, n_12463, n_12464, n_12465, n_12466, n_12467, n_12468,
       n_12469;
  wire n_12470, n_12471, n_12472, n_12473, n_12474, n_12475, n_12476,
       n_12477;
  wire n_12478, n_12479, n_12480, n_12481, n_12482, n_12483, n_12484,
       n_12485;
  wire n_12486, n_12487, n_12488, n_12489, n_12490, n_12491, n_12492,
       n_12493;
  wire n_12494, n_12495, n_12496, n_12497, n_12498, n_12499, n_12500,
       n_12501;
  wire n_12502, n_12503, n_12504, n_12505, n_12506, n_12507, n_12508,
       n_12509;
  wire n_12510, n_12511, n_12512, n_12513, n_12514, n_12515, n_12516,
       n_12517;
  wire n_12518, n_12519, n_12520, n_12521, n_12522, n_12523, n_12524,
       n_12525;
  wire n_12526, n_12527, n_12528, n_12529, n_12530, n_12531, n_12532,
       n_12533;
  wire n_12534, n_12535, n_12536, n_12537, n_12538, n_12539, n_12544,
       n_12545;
  wire n_12546, n_12547, n_12548, n_12549, n_12550, n_12551, n_12552,
       n_12553;
  wire n_12558, n_12559, n_12560, n_12561, n_12562, n_12563, n_12564,
       n_12565;
  wire n_12566, n_12567, n_12568, n_12569, n_12570, n_12571, n_12572,
       n_12573;
  wire n_12574, n_12575, n_12576, n_12577, n_12578, n_12579, n_12580,
       n_12581;
  wire n_12582, n_12583, n_12584, n_12585, n_12586, n_12587, n_12588,
       n_12589;
  wire n_12590, n_12591, n_12592, n_12593, n_12594, n_12595, n_12596,
       n_12597;
  wire n_12598, n_12599, n_12600, n_12601, n_12602, n_12603, n_12604,
       n_12605;
  wire n_12606, n_12607, n_12608, n_12609, n_12610, n_12611, n_12612,
       n_12613;
  wire n_12614, n_12615, n_12616, n_12617, n_12618, n_12619, n_12620,
       n_12621;
  wire n_12622, n_12623, n_12624, n_12625, n_12626, n_12627, n_12628,
       n_12629;
  wire n_12630, n_12631, n_12632, n_12633, n_12634, n_12635, n_12636,
       n_12637;
  wire n_12638, n_12639, n_12640, n_12641, n_12642, n_12643, n_12644,
       n_12645;
  wire n_12646, n_12647, n_12648, n_12649, n_12650, n_12651, n_12652,
       n_12653;
  wire n_12654, n_12655, n_12656, n_12657, n_12658, n_12659, n_12660,
       n_12661;
  wire n_12662, n_12663, n_12664, n_12665, n_12666, n_12667, n_12668,
       n_12669;
  wire n_12670, n_12671, n_12672, n_12673, n_12678, n_12679, n_12680,
       n_12681;
  wire n_12682, n_12683, n_12684, n_12685, n_12686, n_12687, n_12692,
       n_12693;
  wire n_12694, n_12695, n_12696, n_12697, n_12698, n_12699, n_12700,
       n_12701;
  wire n_12702, n_12703, n_12704, n_12705, n_12706, n_12707, n_12708,
       n_12709;
  wire n_12710, n_12711, n_12712, n_12713, n_12714, n_12715, n_12716,
       n_12717;
  wire n_12718, n_12719, n_12720, n_12721, n_12722, n_12723, n_12724,
       n_12725;
  wire n_12726, n_12727, n_12728, n_12729, n_12730, n_12731, n_12732,
       n_12737;
  wire n_12738, n_12739, n_12740, n_12741, n_12742, n_12743, n_12744,
       n_12745;
  wire n_12746, n_12751, n_12752, n_12753, n_12754, n_12755, n_12756,
       n_12757;
  wire n_12758, n_12759, n_12760, n_12761, n_12766, n_12767, n_12768,
       n_12769;
  wire n_12770, n_12771, n_12772, n_12773, n_12774, n_12775, n_12776,
       n_12777;
  wire n_12778, n_12779, n_12780, n_12781, n_12782, n_12783, n_12784,
       n_12785;
  wire n_12786, n_12787, n_12788, n_12789, n_12790, n_12791, n_12792,
       n_12793;
  wire n_12794, n_12795, n_12796, n_12797, n_12798, n_12799, n_12800,
       n_12801;
  wire n_12802, n_12803, n_12804, n_12805, n_12806, n_12811, n_12812,
       n_12813;
  wire n_12814, n_12815, n_12816, n_12817, n_12818, n_12819, n_12820,
       n_12825;
  wire n_12826, n_12827, n_12828, n_12829, n_12830, n_12831, n_12832,
       n_12833;
  wire n_12834, n_12835, n_12840, n_12841, n_12842, n_12843, n_12844,
       n_12845;
  wire n_12846, n_12847, n_12848, n_12849, n_12850, n_12851, n_12852,
       n_12853;
  wire n_12854, n_12855, n_12856, n_12857, n_12858, n_12859, n_12860,
       n_12861;
  wire n_12862, n_12863, n_12864, n_12865, n_12866, n_12867, n_12868,
       n_12869;
  wire n_12870, n_12871, n_12872, n_12873, n_12874, n_12875, n_12876,
       n_12877;
  wire n_12878, n_12879, n_12880, n_12881, n_12886, n_12887, n_12888,
       n_12889;
  wire n_12890, n_12891, n_12892, n_12893, n_12894, n_12895, n_12896,
       n_12897;
  wire n_12898, n_12899, n_12900, n_12901, n_12902, n_12903, n_12904,
       n_12905;
  wire n_12906, n_12907, n_12912, n_12913, n_12914, n_12915, n_12916,
       n_12917;
  wire n_12918, n_12919, n_12920, n_12921, n_12922, n_12923, n_12924,
       n_12925;
  wire n_12926, n_12927, n_12928, n_12929, n_12930, n_12931, n_12932,
       n_12933;
  wire n_12934, n_12935, n_12936, n_12937, n_12938, n_12939, n_12940,
       n_12941;
  wire n_12942, n_12943, n_12944, n_12945, n_12946, n_12947, n_12948,
       n_12949;
  wire n_12950, n_12951, n_12952, n_12953, n_12954, n_12959, n_12960,
       n_12961;
  wire n_12962, n_12963, n_12964, n_12965, n_12966, n_12967, n_12968,
       n_12969;
  wire n_12970, n_12971, n_12972, n_12973, n_12974, n_12975, n_12976,
       n_12977;
  wire n_12978, n_12979, n_12980, n_12981, n_12982, n_12983, n_12984,
       n_12985;
  wire n_12986, n_12987, n_12988, n_12989, n_12990, n_12991, n_12992,
       n_12993;
  wire n_12994, n_12995, n_12996, n_12997, n_12998, n_12999, n_13000,
       n_13001;
  wire n_13002, n_13003, n_13004, n_13005, n_13006, n_13007, n_13008,
       n_13009;
  wire n_13010, n_13011, n_13012, n_13013, n_13014, n_13015, n_13016,
       n_13017;
  wire n_13018, n_13019, n_13020, n_13021, n_13022, n_13023, n_13024,
       n_13025;
  wire n_13026, n_13027, n_13028, n_13029, n_13030, n_13031, n_13032,
       n_13033;
  wire n_13034, n_13035, n_13036, n_13037, n_13038, n_13039, n_13040,
       n_13041;
  wire n_13042, n_13043, n_13044, n_13045, n_13046, n_13047, n_13048,
       n_13049;
  wire n_13050, n_13051, n_13052, n_13053, n_13054, n_13055, n_13056,
       n_13057;
  wire n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064,
       n_13065;
  wire n_13066, n_13067, n_13068, n_13069, n_13070, n_13071, n_13072,
       n_13073;
  wire n_13074, n_13075, n_13076, n_13077, n_13078, n_13079, n_13080,
       n_13081;
  wire n_13082, n_13083, n_13084, n_13085, n_13086, n_13087, n_13088,
       n_13089;
  wire n_13090, n_13091, n_13092, n_13093, n_13094, n_13095, n_13096,
       n_13097;
  wire n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104,
       n_13105;
  wire n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13112,
       n_13113;
  wire n_13114, n_13115, n_13116, n_13117, n_13118, n_13123, n_13124,
       n_13125;
  wire n_13126, n_13127, n_13128, n_13129, n_13130, n_13131, n_13132,
       n_13133;
  wire n_13134, n_13139, n_13140, n_13141, n_13142, n_13143, n_13144,
       n_13145;
  wire n_13146, n_13147, n_13148, n_13149, n_13150, n_13151, n_13152,
       n_13153;
  wire n_13154, n_13155, n_13156, n_13157, n_13158, n_13159, n_13160,
       n_13161;
  wire n_13162, n_13163, n_13164, n_13165, n_13166, n_13167, n_13172,
       n_13173;
  wire n_13174, n_13175, n_13176, n_13177, n_13178, n_13179, n_13180,
       n_13181;
  wire n_13182, n_13187, n_13188, n_13189, n_13190, n_13191, n_13192,
       n_13193;
  wire n_13194, n_13195, n_13196, n_13197, n_13202, n_13203, n_13204,
       n_13205;
  wire n_13206, n_13207, n_13208, n_13209, n_13210, n_13211, n_13212,
       n_13217;
  wire n_13218, n_13219, n_13220, n_13221, n_13222, n_13223, n_13224,
       n_13225;
  wire n_13226, n_13227, n_13232, n_13233, n_13234, n_13235, n_13236,
       n_13237;
  wire n_13238, n_13239, n_13240, n_13241, n_13242, n_13247, n_13248,
       n_13249;
  wire n_13250, n_13251, n_13252, n_13253, n_13254, n_13255, n_13256,
       n_13257;
  wire n_13262, n_13263, n_13264, n_13265, n_13266, n_13267, n_13268,
       n_13269;
  wire n_13270, n_13271, n_13272, n_13277, n_13278, n_13279, n_13280,
       n_13281;
  wire n_13282, n_13283, n_13284, n_13285, n_13286, n_13287, n_13292,
       n_13293;
  wire n_13294, n_13295, n_13296, n_13297, n_13298, n_13299, n_13300,
       n_13301;
  wire n_13302, n_13303, n_13304, n_13305, n_13306, n_13307, n_13308,
       n_13309;
  wire n_13310, n_13311, n_13312, n_13313, n_13314, n_13315, n_13316,
       n_13317;
  wire n_13318, n_13319, n_13320, n_13321, n_13322, n_13327, n_13328,
       n_13329;
  wire n_13330, n_13331, n_13332, n_13333, n_13334, n_13335, n_13336,
       n_13341;
  wire n_13342, n_13343, n_13344, n_13345, n_13346, n_13347, n_13348,
       n_13349;
  wire n_13350, n_13351, n_13356, n_13357, n_13358, n_13359, n_13360,
       n_13361;
  wire n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368,
       n_13369;
  wire n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376,
       n_13377;
  wire n_13378, n_13379, n_13380, n_13381, n_13382, n_13383, n_13384,
       n_13385;
  wire n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392,
       n_13393;
  wire n_13394, n_13395, n_13396, n_13401, n_13402, n_13403, n_13404,
       n_13405;
  wire n_13406, n_13407, n_13408, n_13409, n_13410, n_13415, n_13416,
       n_13417;
  wire n_13418, n_13419, n_13420, n_13421, n_13422, n_13423, n_13424,
       n_13425;
  wire n_13430, n_13431, n_13432, n_13433, n_13434, n_13435, n_13436,
       n_13437;
  wire n_13438, n_13439, n_13440, n_13441, n_13442, n_13443, n_13444,
       n_13445;
  wire n_13446, n_13447, n_13448, n_13449, n_13450, n_13451, n_13452,
       n_13453;
  wire n_13454, n_13455, n_13456, n_13457, n_13458, n_13459, n_13460,
       n_13461;
  wire n_13462, n_13463, n_13464, n_13465, n_13466, n_13467, n_13468,
       n_13469;
  wire n_13470, n_13475, n_13476, n_13477, n_13478, n_13479, n_13480,
       n_13481;
  wire n_13482, n_13483, n_13484, n_13489, n_13490, n_13491, n_13492,
       n_13493;
  wire n_13494, n_13495, n_13496, n_13497, n_13498, n_13499, n_13504,
       n_13505;
  wire n_13506, n_13507, n_13508, n_13509, n_13510, n_13511, n_13512,
       n_13513;
  wire n_13514, n_13515, n_13516, n_13517, n_13518, n_13519, n_13520,
       n_13521;
  wire n_13522, n_13523, n_13524, n_13525, n_13526, n_13527, n_13528,
       n_13529;
  wire n_13530, n_13531, n_13532, n_13533, n_13534, n_13535, n_13536,
       n_13537;
  wire n_13538, n_13539, n_13540, n_13541, n_13542, n_13543, n_13544,
       n_13545;
  wire n_13550, n_13551, n_13552, n_13553, n_13554, n_13555, n_13556,
       n_13557;
  wire n_13558, n_13559, n_13560, n_13561, n_13562, n_13563, n_13564,
       n_13565;
  wire n_13566, n_13567, n_13568, n_13569, n_13570, n_13571, n_13576,
       n_13577;
  wire n_13578, n_13579, n_13580, n_13581, n_13582, n_13583, n_13584,
       n_13585;
  wire n_13586, n_13587, n_13588, n_13589, n_13590, n_13591, n_13592,
       n_13593;
  wire n_13594, n_13595, n_13596, n_13597, n_13598, n_13599, n_13600,
       n_13601;
  wire n_13602, n_13603, n_13604, n_13605, n_13606, n_13607, n_13608,
       n_13609;
  wire n_13610, n_13611, n_13612, n_13613, n_13614, n_13615, n_13616,
       n_13617;
  wire n_13618, n_13623, n_13624, n_13625, n_13626, n_13627, n_13628,
       n_13629;
  wire n_13630, n_13631, n_13632, n_13633, n_13634, n_13635, n_13636,
       n_13637;
  wire n_13638, n_13639, n_13640, n_13641, n_13642, n_13643, n_13644,
       n_13645;
  wire n_13646, n_13647, n_13648, n_13649, n_13650, n_13651, n_13652,
       n_13653;
  wire n_13654, n_13655, n_13656, n_13657, n_13658, n_13659, n_13660,
       n_13661;
  wire n_13662, n_13663, n_13664, n_13665, n_13666, n_13667, n_13668,
       n_13669;
  wire n_13670, n_13671, n_13672, n_13673, n_13674, n_13675, n_13676,
       n_13677;
  wire n_13678, n_13679, n_13680, n_13681, n_13682, n_13683, n_13684,
       n_13685;
  wire n_13686, n_13687, n_13688, n_13689, n_13690, n_13691, n_13692,
       n_13693;
  wire n_13694, n_13695, n_13696, n_13697, n_13698, n_13699, n_13700,
       n_13701;
  wire n_13702, n_13703, n_13704, n_13705, n_13706, n_13707, n_13708,
       n_13709;
  wire n_13710, n_13711, n_13712, n_13713, n_13714, n_13715, n_13716,
       n_13717;
  wire n_13718, n_13719, n_13720, n_13721, n_13722, n_13723, n_13724,
       n_13725;
  wire n_13726, n_13727, n_13728, n_13729, n_13730, n_13731, n_13732,
       n_13733;
  wire n_13734, n_13735, n_13736, n_13737, n_13738, n_13739, n_13740,
       n_13741;
  wire n_13742, n_13743, n_13744, n_13745, n_13746, n_13747, n_13748,
       n_13749;
  wire n_13750, n_13751, n_13752, n_13753, n_13754, n_13755, n_13756,
       n_13757;
  wire n_13758, n_13759, n_13760, n_13761, n_13762, n_13763, n_13764,
       n_13765;
  wire n_13766, n_13767, n_13768, n_13769, n_13770, n_13771, n_13772,
       n_13773;
  wire n_13774, n_13775, n_13776, n_13777, n_13778, n_13779, n_13780,
       n_13781;
  wire n_13782, n_13783, n_13784, n_13785, n_13786, n_13787, n_13788,
       n_13789;
  wire n_13790, n_13791, n_13792, n_13793, n_13794, n_13795, n_13796,
       n_13797;
  wire n_13798, n_13799, n_13800, n_13801, n_13802, n_13803, n_13804,
       n_13805;
  wire n_13806, n_13807, n_13808, n_13809, n_13810, n_13811, n_13812,
       n_13813;
  wire n_13814, n_13815, n_13816, n_13817, n_13818, n_13819, n_13820,
       n_13821;
  wire n_13822, n_13823, n_13824, n_13825, n_13826, n_13827, n_13828,
       n_13829;
  wire n_13830, n_13831, n_13832, n_13833, n_13834, n_13835, n_13836,
       n_13837;
  wire n_13838, n_13839, n_13840, n_13841, n_13842, n_13843, n_13844,
       n_13845;
  wire n_13846, n_13847, n_13848, n_13849, n_13850, n_13851, n_13852,
       n_13853;
  wire n_13854, n_13855, n_13856, n_13857, n_13858, n_13859, n_13860,
       n_13861;
  wire n_13862, n_13863, n_13864, n_13865, n_13866, n_13867, n_13868,
       n_13869;
  wire n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13882,
       n_13887;
  wire n_13888, n_13889, n_13890, n_13891, n_13892, n_13893, n_13894,
       n_13895;
  wire n_13896, n_13897, n_13898, n_13899, n_13900, n_13901, n_13902,
       n_13903;
  wire n_13904, n_13905, n_13906, n_13907, n_13908, n_13909, n_13910,
       n_13915;
  wire n_13916, n_13917, n_13918, n_13919, n_13920, n_13921, n_13922,
       n_13923;
  wire n_13924, n_13925, n_13926, n_13927, n_13928, n_13929, n_13930,
       n_13931;
  wire n_13932, n_13933, n_13934, n_13935, n_13936, n_13937, n_13942,
       n_13943;
  wire n_13944, n_13945, n_13946, n_13947, n_13948, n_13949, n_13950,
       n_13951;
  wire n_13952, n_13953, n_13954, n_13955, n_13956, n_13957, n_13958,
       n_13959;
  wire n_13960, n_13961, n_13962, n_13963, n_13964, n_13965, n_13966,
       n_13967;
  wire n_13968, n_13969, n_13970, n_13971, n_13972, n_13973, n_13974,
       n_13975;
  wire n_13976, n_13977, n_13978, n_13979, n_13980, n_13981, n_13982,
       n_13983;
  wire n_13984, n_13985, n_13986, n_13987, n_13988, n_13989, n_13990,
       n_13991;
  wire n_13992, n_13993, n_13994, n_13999, n_14000, n_14001, n_14002,
       n_14003;
  wire n_14004, n_14005, n_14006, n_14007, n_14008, n_14013, n_14014,
       n_14015;
  wire n_14016, n_14017, n_14018, n_14019, n_14020, n_14021, n_14026,
       n_14027;
  wire n_14028, n_14029, n_14030, n_14031, n_14032, n_14033, n_14034,
       n_14035;
  wire n_14036, n_14037, n_14038, n_14039, n_14040, n_14041, n_14042,
       n_14043;
  wire n_14044, n_14045, n_14046, n_14047, n_14048, n_14049, n_14050,
       n_14051;
  wire n_14052, n_14053, n_14054, n_14055, n_14056, n_14057, n_14058,
       n_14059;
  wire n_14060, n_14061, n_14062, n_14063, n_14064, n_14065, n_14066,
       n_14067;
  wire n_14068, n_14069, n_14070, n_14071, n_14072, n_14073, n_14074,
       n_14075;
  wire n_14076, n_14077, n_14082, n_14083, n_14084, n_14085, n_14086,
       n_14087;
  wire n_14088, n_14089, n_14090, n_14091, n_14096, n_14097, n_14098,
       n_14099;
  wire n_14100, n_14101, n_14102, n_14103, n_14104, n_14109, n_14110,
       n_14111;
  wire n_14112, n_14113, n_14114, n_14115, n_14116, n_14117, n_14118,
       n_14119;
  wire n_14120, n_14121, n_14122, n_14123, n_14124, n_14125, n_14126,
       n_14127;
  wire n_14128, n_14129, n_14130, n_14131, n_14132, n_14133, n_14134,
       n_14135;
  wire n_14136, n_14137, n_14138, n_14139, n_14140, n_14141, n_14142,
       n_14143;
  wire n_14144, n_14145, n_14146, n_14147, n_14148, n_14149, n_14150,
       n_14151;
  wire n_14152, n_14153, n_14154, n_14155, n_14156, n_14157, n_14158,
       n_14159;
  wire n_14160, n_14165, n_14166, n_14167, n_14168, n_14169, n_14170,
       n_14171;
  wire n_14172, n_14173, n_14174, n_14179, n_14180, n_14181, n_14182,
       n_14183;
  wire n_14184, n_14185, n_14186, n_14187, n_14192, n_14193, n_14194,
       n_14195;
  wire n_14196, n_14197, n_14198, n_14199, n_14200, n_14201, n_14202,
       n_14203;
  wire n_14204, n_14205, n_14206, n_14207, n_14208, n_14209, n_14210,
       n_14211;
  wire n_14212, n_14213, n_14214, n_14215, n_14216, n_14217, n_14218,
       n_14219;
  wire n_14220, n_14221, n_14222, n_14223, n_14224, n_14225, n_14226,
       n_14227;
  wire n_14228, n_14229, n_14230, n_14231, n_14232, n_14233, n_14234,
       n_14235;
  wire n_14236, n_14237, n_14238, n_14239, n_14240, n_14241, n_14242,
       n_14243;
  wire n_14248, n_14249, n_14250, n_14251, n_14252, n_14253, n_14254,
       n_14255;
  wire n_14256, n_14261, n_14262, n_14263, n_14264, n_14265, n_14266,
       n_14267;
  wire n_14268, n_14269, n_14270, n_14271, n_14272, n_14273, n_14274,
       n_14275;
  wire n_14276, n_14277, n_14278, n_14279, n_14280, n_14281, n_14282,
       n_14283;
  wire n_14284, n_14285, n_14286, n_14287, n_14288, n_14289, n_14290,
       n_14291;
  wire n_14292, n_14293, n_14294, n_14295, n_14296, n_14297, n_14298,
       n_14299;
  wire n_14300, n_14301, n_14302, n_14303, n_14304, n_14305, n_14306,
       n_14307;
  wire n_14308, n_14309, n_14310, n_14311, n_14312, n_14313, n_14314,
       n_14315;
  wire n_14316, n_14317, n_14318, n_14319, n_14320, n_14321, n_14322,
       n_14323;
  wire n_14324, n_14325, n_14326, n_14327, n_14328, n_14329, n_14330,
       n_14331;
  wire n_14332, n_14333, n_14334, n_14335, n_14336, n_14337, n_14338,
       n_14339;
  wire n_14340, n_14341, n_14342, n_14343, n_14344, n_14345, n_14346,
       n_14347;
  wire n_14348, n_14349, n_14350, n_14351, n_14352, n_14353, n_14354,
       n_14355;
  wire n_14356, n_14357, n_14358, n_14359, n_14360, n_14361, n_14362,
       n_14363;
  wire n_14364, n_14365, n_14366, n_14367, n_14368, n_14369, n_14370,
       n_14371;
  wire n_14372, n_14373, n_14374, n_14375, n_14376, n_14377, n_14378,
       n_14379;
  wire n_14380, n_14381, n_14386, n_14387, n_14388, n_14389, n_14390,
       n_14391;
  wire n_14392, n_14393, n_14394, n_14399, n_14400, n_14401, n_14402,
       n_14403;
  wire n_14404, n_14405, n_14406, n_14407, n_14408, n_14409, n_14410,
       n_14411;
  wire n_14412, n_14413, n_14414, n_14415, n_14416, n_14417, n_14418,
       n_14419;
  wire n_14420, n_14421, n_14422, n_14427, n_14428, n_14429, n_14430,
       n_14431;
  wire n_14432, n_14433, n_14434, n_14435, n_14436, n_14437, n_14438,
       n_14439;
  wire n_14440, n_14441, n_14442, n_14443, n_14444, n_14445, n_14446,
       n_14447;
  wire n_14448, n_14449, n_14453, n_14454, n_14455, n_14456, n_14457,
       n_14458;
  wire n_14459, n_14460, n_14461, n_14462, n_14463, n_14464, n_14465,
       n_14466;
  wire n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, n_14473,
       n_14474;
  wire n_14475, n_14476, n_14477, n_14478, n_14479, n_14480, n_14481,
       n_14482;
  wire n_14483, n_14484, n_14485, n_14486, n_14487, n_14488, n_14489,
       n_14490;
  wire n_14491, n_14492, n_14493, n_14494, n_14495, n_14496, n_14497,
       n_14498;
  wire n_14499, n_14500, n_14501, n_14502, n_14503, n_14504, n_14505,
       n_14506;
  wire n_14507, n_14508, n_14509, n_14510, n_14511, n_14512, n_14513,
       n_14514;
  wire n_14515, n_14516, n_14517, n_14518, n_14519, n_14520, n_14521,
       n_14522;
  wire n_14523, n_14524, n_14525, n_14526, n_14527, n_14528, n_14529,
       n_14530;
  wire n_14531, n_14532, n_14533, n_14534, n_14535, n_14536, n_14537,
       n_14538;
  wire n_14539, n_14540, n_14541, n_14542, n_14543, n_14544, n_14545,
       n_14546;
  wire n_14547, n_14548, n_14549, n_14550, n_14551, n_14552, n_14553,
       n_14554;
  wire n_14555, n_14556, n_14557, n_14558, n_14559, n_14560, n_14561,
       n_14562;
  wire n_14563, n_14564, n_14565, n_14566, n_14567, n_14568, n_14569,
       n_14570;
  wire n_14571, n_14572, n_14573, n_14574, n_14575, n_14576, n_14577,
       n_14578;
  wire n_14579, n_14580, n_14581, n_14582, n_14583, n_14584, n_14585,
       n_14586;
  wire n_14587, n_14588, n_14589, n_14590, n_14591, n_14592, n_14593,
       n_14594;
  wire n_14595, n_14596, n_14597, n_14598, n_14599, n_14600, n_14601,
       n_14602;
  wire n_14603, n_14604, n_14605, n_14606, n_14607, n_14608, n_14609,
       n_14610;
  wire n_14611, n_14612, n_14613, n_14614, n_14615, n_14616, n_14617,
       n_14618;
  wire n_14619, n_14620, n_14621, n_14622, n_14623, n_14624, n_14625,
       n_14626;
  wire n_14627, n_14628, n_14629, n_14630, n_14631, n_14632, n_14633,
       n_14634;
  wire n_14635, n_14636, n_14637, n_14638, n_14639, n_14640, n_14641,
       n_14642;
  wire n_14643, n_14644, n_14645, n_14646, n_14647, n_14648, n_14649,
       n_14650;
  wire n_14651, n_14652, n_14653, n_14654, n_14655, n_14656, n_14657,
       n_14659;
  wire n_14660, n_14661, n_14662, n_14666, n_14667, n_14669, n_14670,
       n_14671;
  wire n_14672, n_14676, n_14677, n_14678, n_14680, n_14681, n_14682,
       n_14683;
  wire n_14687, n_14688, n_14690, n_14691, n_14692, n_14693, n_14697,
       n_14698;
  wire n_14700, n_14701, n_14702, n_14703, n_14707, n_14708, n_14710,
       n_14711;
  wire n_14712, n_14713, n_14714, n_14715, n_14716, n_14717, n_14718,
       n_14719;
  wire n_14720, n_14721, n_14722, n_14723, n_14724, n_14725, n_14726,
       n_14727;
  wire n_14728, n_14729, n_14730, n_14731, n_14732, n_14733, n_14734,
       n_14735;
  wire n_14736, n_14737, n_14738, n_14739, n_14740, n_14741, n_14742,
       n_14743;
  wire n_14744, n_14745, n_14746, n_14747, n_14748, n_14749, n_14753,
       n_14754;
  wire n_14756, n_14757, n_14758, n_14759, n_14760, n_14761, n_14762,
       n_14763;
  wire n_14764, n_14765, n_14766, n_14767, n_14768, n_14769, n_14770,
       n_14771;
  wire n_14772, n_14773, n_14774, n_14775, n_14776, n_14777, n_14778,
       n_14779;
  wire n_14780, n_14781, n_14782, n_14783, n_14784, n_14785, n_14786,
       n_14787;
  wire n_14788, n_14789, n_14790, n_14791, n_14792, n_14793, n_14794,
       n_14795;
  wire n_14796, n_14797, n_14798, n_14799, n_14800, n_14805, n_14806,
       n_14807;
  wire n_14808, n_14809, n_14810, n_14811, n_14812, n_14813, n_14814,
       n_14815;
  wire n_14816, n_14817, n_14818, n_14819, n_14820, n_14821, n_14822,
       n_14827;
  wire n_14828, n_14829, n_14830, n_14831, n_14832, n_14833, n_14834,
       n_14835;
  wire n_14836, n_14837, n_14838, n_14839, n_14840, n_14841, n_14842,
       n_14843;
  wire n_14844, n_14845, n_14846, n_14847, n_14848, n_14849, n_14850,
       n_14851;
  wire n_14852, n_14853, n_14854, n_14855, n_14856, n_14857, n_14858,
       n_14859;
  wire n_14860, n_14861, n_14862, n_14863, n_14864, n_14865, n_14866,
       n_14867;
  wire n_14868, n_14869, n_14870, n_14871, n_14872, n_14873, n_14874,
       n_14875;
  wire n_14876, n_14877, n_14878, n_14879, n_14880, n_14881, n_14882,
       n_14883;
  wire n_14884, n_14885, n_14886, n_14887, n_14888, n_14889, n_14890,
       n_14891;
  wire n_14892, n_14893, n_14894, n_14895, n_14896, n_14897, n_14898,
       n_14899;
  wire n_14900, n_14905, n_14906, n_14907, n_14908, n_14909, n_14910,
       n_14911;
  wire n_14912, n_14913, n_14914, n_14915, n_14916, n_14917, n_14918,
       n_14919;
  wire n_14920, n_14921, n_14922, n_14923, n_14924, n_14925, n_14926,
       n_14927;
  wire n_14932, n_14933, n_14934, n_14935, n_14936, n_14937, n_14938,
       n_14939;
  wire n_14940, n_14941, n_14942, n_14943, n_14944, n_14945, n_14946,
       n_14947;
  wire n_14948, n_14949, n_14950, n_14951, n_14952, n_14953, n_14954,
       n_14955;
  wire n_14956, n_14957, n_14958, n_14959, n_14960, n_14961, n_14962,
       n_14963;
  wire n_14964, n_14965, n_14966, n_14967, n_14968, n_14969, n_14970,
       n_14971;
  wire n_14972, n_14973, n_14974, n_14979, n_14980, n_14981, n_14982,
       n_14983;
  wire n_14984, n_14985, n_14986, n_14987, n_14988, n_14989, n_14990,
       n_14991;
  wire n_14992, n_14993, n_14994, n_14995, n_14996, n_14997, n_14998,
       n_14999;
  wire n_15000, n_15001, n_15002, n_15003, n_15004, n_15005, n_15006,
       n_15007;
  wire n_15008, n_15009, n_15010, n_15011, n_15012, n_15013, n_15014,
       n_15015;
  wire n_15016, n_15017, n_15018, n_15019, n_15020, n_15021, n_15022,
       n_15023;
  wire n_15024, n_15025, n_15026, n_15030, n_15031, n_15033, n_15034,
       n_15035;
  wire n_15036, n_15037, n_15038, n_15039, n_15040, n_15041, n_15042,
       n_15046;
  wire n_15047, n_15049, n_15050, n_15051, n_15052, n_15053, n_15054,
       n_15055;
  wire n_15056, n_15057, n_15058, n_15059, n_15060, n_15061, n_15062,
       n_15063;
  wire n_15064, n_15065, n_15066, n_15067, n_15068, n_15069, n_15070,
       n_15071;
  wire n_15072, n_15073, n_15074, n_15075, n_15076, n_15077, n_15078,
       n_15079;
  wire n_15080, n_15081, n_15082, n_15083, n_15084, n_15085, n_15086,
       n_15087;
  wire n_15088, n_15089, n_15090, n_15091, n_15096, n_15097, n_15098,
       n_15099;
  wire n_15100, n_15101, n_15102, n_15103, n_15104, n_15105, n_15106,
       n_15107;
  wire n_15108, n_15109, n_15110, n_15111, n_15112, n_15113, n_15114,
       n_15115;
  wire n_15116, n_15117, n_15122, n_15123, n_15124, n_15125, n_15126,
       n_15127;
  wire n_15128, n_15129, n_15130, n_15131, n_15132, n_15133, n_15134,
       n_15135;
  wire n_15136, n_15137, n_15138, n_15139, n_15140, n_15141, n_15142,
       n_15143;
  wire n_15144, n_15145, n_15146, n_15147, n_15148, n_15149, n_15150,
       n_15151;
  wire n_15152, n_15153, n_15154, n_15155, n_15156, n_15157, n_15158,
       n_15159;
  wire n_15160, n_15161, n_15162, n_15163, n_15164, n_15169, n_15170,
       n_15171;
  wire n_15172, n_15173, n_15174, n_15175, n_15176, n_15177, n_15178,
       n_15179;
  wire n_15180, n_15181, n_15182, n_15183, n_15184, n_15185, n_15186,
       n_15187;
  wire n_15188, n_15189, n_15190, n_15191, n_15192, n_15193, n_15194,
       n_15195;
  wire n_15196, n_15197, n_15198, n_15199, n_15200, n_15201, n_15202,
       n_15203;
  wire n_15204, n_15205, n_15206, n_15207, n_15208, n_15209, n_15210,
       n_15211;
  wire n_15212, n_15213, n_15214, n_15215, n_15216, n_15217, n_15218,
       n_15219;
  wire n_15224, n_15225, n_15226, n_15227, n_15232, n_15233, n_15234,
       n_15235;
  wire n_15236, n_15241, n_15242, n_15243, n_15244, n_15245, n_15246,
       n_15247;
  wire n_15248, n_15249, n_15250, n_15251, n_15252, n_15253, n_15254,
       n_15255;
  wire n_15256, n_15257, n_15258, n_15259, n_15260, n_15261, n_15262,
       n_15263;
  wire n_15264, n_15265, n_15266, n_15267, n_15268, n_15269, n_15270,
       n_15271;
  wire n_15272, n_15273, n_15274, n_15275, n_15276, n_15277, n_15278,
       n_15279;
  wire n_15280, n_15281, n_15282, n_15283, n_15284, n_15285, n_15286,
       n_15287;
  wire n_15288, n_15289, n_15290, n_15291, n_15292, n_15293, n_15294,
       n_15295;
  wire n_15296, n_15297, n_15298, n_15299, n_15300, n_15301, n_15302,
       n_15303;
  wire n_15304, n_15305, n_15306, n_15310, n_15311, n_15312, n_15314,
       n_15315;
  wire n_15316, n_15317, n_15318, n_15319, n_15320, n_15321, n_15322,
       n_15323;
  wire n_15324, n_15325, n_15326, n_15327, n_15328, n_15329, n_15330,
       n_15331;
  wire n_15332, n_15333, n_15334, n_15335, n_15336, n_15337, n_15338,
       n_15339;
  wire n_15340, n_15341, n_15342, n_15343, n_15344, n_15345, n_15346,
       n_15347;
  wire n_15351, n_15353, n_15354, n_15355, n_15356, n_15357, n_15358,
       n_15359;
  wire n_15360, n_15361, n_15362, n_15367, n_15368, n_15369, n_15370,
       n_15371;
  wire n_15372, n_15373, n_15374, n_15375, n_15376, n_15377, n_15382,
       n_15383;
  wire n_15384, n_15385, n_15386, n_15387, n_15388, n_15389, n_15390,
       n_15391;
  wire n_15392, n_15393, n_15394, n_15395, n_15396, n_15397, n_15398,
       n_15399;
  wire n_15400, n_15401, n_15402, n_15403, n_15404, n_15405, n_15406,
       n_15407;
  wire n_15408, n_15409, n_15410, n_15411, n_15412, n_15413, n_15414,
       n_15415;
  wire n_15416, n_15417, n_15418, n_15419, n_15420, n_15421, n_15422,
       n_15423;
  wire n_15428, n_15429, n_15430, n_15431, n_15432, n_15433, n_15434,
       n_15435;
  wire n_15436, n_15437, n_15438, n_15439, n_15440, n_15441, n_15442,
       n_15443;
  wire n_15444, n_15445, n_15446, n_15447, n_15448, n_15449, n_15454,
       n_15455;
  wire n_15456, n_15457, n_15458, n_15459, n_15460, n_15461, n_15462,
       n_15463;
  wire n_15464, n_15465, n_15466, n_15467, n_15468, n_15469, n_15470,
       n_15471;
  wire n_15472, n_15473, n_15474, n_15475, n_15476, n_15477, n_15478,
       n_15479;
  wire n_15480, n_15481, n_15482, n_15483, n_15484, n_15485, n_15486,
       n_15487;
  wire n_15488, n_15489, n_15490, n_15491, n_15492, n_15493, n_15494,
       n_15495;
  wire n_15496, n_15501, n_15502, n_15503, n_15504, n_15505, n_15506,
       n_15507;
  wire n_15508, n_15509, n_15510, n_15511, n_15512, n_15513, n_15514,
       n_15515;
  wire n_15516, n_15517, n_15518, n_15519, n_15520, n_15521, n_15522,
       n_15523;
  wire n_15524, n_15525, n_15526, n_15527, n_15528, n_15529, n_15530,
       n_15531;
  wire n_15532, n_15533, n_15534, n_15535, n_15536, n_15537, n_15538,
       n_15539;
  wire n_15540, n_15541, n_15542, n_15543, n_15544, n_15545, n_15546,
       n_15547;
  wire n_15548, n_15549, n_15550, n_15551, n_15552, n_15553, n_15554,
       n_15555;
  wire n_15556, n_15557, n_15558, n_15559, n_15560, n_15561, n_15562,
       n_15563;
  wire n_15564, n_15565, n_15566, n_15567, n_15568, n_15569, n_15570,
       n_15571;
  wire n_15572, n_15573, n_15574, n_15575, n_15576, n_15577, n_15578,
       n_15579;
  wire n_15580, n_15581, n_15582, n_15583, n_15584, n_15585, n_15586,
       n_15587;
  wire n_15588, n_15589, n_15593, n_15594, n_15596, n_15597, n_15598,
       n_15599;
  wire n_15600, n_15601, n_15602, n_15603, n_15604, n_15605, n_15610,
       n_15611;
  wire n_15612, n_15613, n_15614, n_15615, n_15616, n_15617, n_15618,
       n_15619;
  wire n_15620, n_15621, n_15622, n_15623, n_15624, n_15625, n_15626,
       n_15627;
  wire n_15628, n_15629, n_15630, n_15631, n_15632, n_15633, n_15634,
       n_15635;
  wire n_15636, n_15637, n_15638, n_15639, n_15640, n_15641, n_15642,
       n_15643;
  wire n_15644, n_15645, n_15646, n_15647, n_15648, n_15649, n_15650,
       n_15655;
  wire n_15656, n_15657, n_15658, n_15659, n_15660, n_15661, n_15662,
       n_15663;
  wire n_15664, n_15669, n_15670, n_15671, n_15672, n_15673, n_15674,
       n_15675;
  wire n_15676, n_15677, n_15678, n_15679, n_15684, n_15685, n_15686,
       n_15687;
  wire n_15688, n_15689, n_15690, n_15691, n_15692, n_15693, n_15694,
       n_15695;
  wire n_15696, n_15697, n_15698, n_15699, n_15700, n_15701, n_15702,
       n_15703;
  wire n_15704, n_15705, n_15706, n_15707, n_15708, n_15709, n_15710,
       n_15711;
  wire n_15712, n_15713, n_15714, n_15715, n_15716, n_15717, n_15718,
       n_15719;
  wire n_15720, n_15721, n_15722, n_15723, n_15724, n_15725, n_15730,
       n_15731;
  wire n_15732, n_15733, n_15734, n_15735, n_15736, n_15737, n_15738,
       n_15739;
  wire n_15740, n_15741, n_15742, n_15743, n_15744, n_15745, n_15746,
       n_15747;
  wire n_15748, n_15749, n_15750, n_15751, n_15756, n_15757, n_15758,
       n_15759;
  wire n_15760, n_15761, n_15762, n_15763, n_15764, n_15765, n_15766,
       n_15767;
  wire n_15768, n_15769, n_15770, n_15771, n_15772, n_15773, n_15774,
       n_15775;
  wire n_15776, n_15777, n_15778, n_15779, n_15780, n_15781, n_15782,
       n_15783;
  wire n_15784, n_15785, n_15786, n_15787, n_15788, n_15789, n_15790,
       n_15791;
  wire n_15792, n_15793, n_15794, n_15795, n_15796, n_15797, n_15798,
       n_15803;
  wire n_15804, n_15805, n_15806, n_15807, n_15808, n_15809, n_15810,
       n_15811;
  wire n_15812, n_15813, n_15814, n_15815, n_15816, n_15817, n_15818,
       n_15819;
  wire n_15820, n_15821, n_15822, n_15823, n_15824, n_15825, n_15826,
       n_15827;
  wire n_15828, n_15829, n_15830, n_15831, n_15832, n_15833, n_15834,
       n_15835;
  wire n_15836, n_15837, n_15838, n_15839, n_15840, n_15841, n_15842,
       n_15843;
  wire n_15844, n_15845, n_15846, n_15847, n_15848, n_15849, n_15850,
       n_15851;
  wire n_15852, n_15853, n_15854, n_15855, n_15856, n_15857, n_15858,
       n_15859;
  wire n_15860, n_15861, n_15862, n_15863, n_15864, n_15865, n_15866,
       n_15867;
  wire n_15868, n_15869, n_15870, n_15871, n_15872, n_15873, n_15874,
       n_15875;
  wire n_15876, n_15877, n_15878, n_15879, n_15880, n_15881, n_15882,
       n_15883;
  wire n_15884, n_15885, n_15890, n_15891, n_15892, n_15893, n_15898,
       n_15899;
  wire n_15900, n_15901, n_15906, n_15907, n_15908, n_15909, n_15914,
       n_15915;
  wire n_15916, n_15917, n_15918, n_15919, n_15920, n_15921, n_15922,
       n_15923;
  wire n_15924, n_15925, n_15926, n_15927, n_15928, n_15929, n_15930,
       n_15931;
  wire n_15932, n_15933, n_15934, n_15935, n_15936, n_15937, n_15938,
       n_15939;
  wire n_15940, n_15941, n_15942, n_15943, n_15944, n_15945, n_15946,
       n_15947;
  wire n_15948, n_15949, n_15950, n_15951, n_15952, n_15953, n_15954,
       n_15955;
  wire n_15956, n_15957, n_15958, n_15959, n_15960, n_15961, n_15962,
       n_15963;
  wire n_15964, n_15965, n_15966, n_15967, n_15968, n_15969, n_15970,
       n_15971;
  wire n_15972, n_15973, n_15974, n_15975, n_15976, n_15977, n_15978,
       n_15979;
  wire n_15980, n_15981, n_15982, n_15983, n_15984, n_15985, n_15986,
       n_15987;
  wire n_15988, n_15989, n_15990, n_15991, n_15992, n_15993, n_15994,
       n_15995;
  wire n_15996, n_15997, n_15998, n_15999, n_16000, n_16001, n_16002,
       n_16003;
  wire n_16004, n_16005, n_16006, n_16007, n_16008, n_16009, n_16013,
       n_16014;
  wire n_16015, n_16017, n_16018, n_16019, n_16020, n_16021, n_16022,
       n_16023;
  wire n_16024, n_16025, n_16026, n_16027, n_16031, n_16032, n_16033,
       n_16035;
  wire n_16036, n_16037, n_16038, n_16039, n_16040, n_16041, n_16042,
       n_16043;
  wire n_16044, n_16045, n_16046, n_16047, n_16048, n_16049, n_16050,
       n_16051;
  wire n_16052, n_16053, n_16054, n_16055, n_16056, n_16057, n_16058,
       n_16059;
  wire n_16060, n_16061, n_16062, n_16063, n_16064, n_16065, n_16069,
       n_16071;
  wire n_16072, n_16073, n_16074, n_16075, n_16076, n_16077, n_16078,
       n_16079;
  wire n_16080, n_16085, n_16086, n_16087, n_16088, n_16089, n_16090,
       n_16091;
  wire n_16092, n_16093, n_16094, n_16095, n_16100, n_16101, n_16102,
       n_16103;
  wire n_16104, n_16105, n_16106, n_16107, n_16108, n_16109, n_16110,
       n_16111;
  wire n_16112, n_16113, n_16114, n_16115, n_16116, n_16117, n_16118,
       n_16119;
  wire n_16120, n_16121, n_16122, n_16123, n_16124, n_16125, n_16126,
       n_16127;
  wire n_16128, n_16129, n_16130, n_16131, n_16132, n_16133, n_16134,
       n_16135;
  wire n_16136, n_16137, n_16138, n_16139, n_16140, n_16145, n_16146,
       n_16147;
  wire n_16148, n_16149, n_16150, n_16151, n_16152, n_16153, n_16154,
       n_16159;
  wire n_16160, n_16161, n_16162, n_16163, n_16164, n_16165, n_16166,
       n_16167;
  wire n_16168, n_16169, n_16174, n_16175, n_16176, n_16177, n_16178,
       n_16179;
  wire n_16180, n_16181, n_16182, n_16183, n_16184, n_16185, n_16186,
       n_16187;
  wire n_16188, n_16189, n_16190, n_16191, n_16192, n_16193, n_16194,
       n_16195;
  wire n_16196, n_16197, n_16198, n_16199, n_16200, n_16201, n_16202,
       n_16203;
  wire n_16204, n_16205, n_16206, n_16207, n_16208, n_16209, n_16210,
       n_16211;
  wire n_16212, n_16213, n_16214, n_16215, n_16220, n_16221, n_16222,
       n_16223;
  wire n_16224, n_16225, n_16226, n_16227, n_16228, n_16229, n_16230,
       n_16231;
  wire n_16232, n_16233, n_16234, n_16235, n_16236, n_16237, n_16238,
       n_16239;
  wire n_16240, n_16241, n_16246, n_16247, n_16248, n_16249, n_16250,
       n_16251;
  wire n_16252, n_16253, n_16254, n_16255, n_16256, n_16257, n_16258,
       n_16259;
  wire n_16260, n_16261, n_16262, n_16263, n_16264, n_16265, n_16266,
       n_16267;
  wire n_16268, n_16269, n_16270, n_16271, n_16272, n_16273, n_16274,
       n_16275;
  wire n_16276, n_16277, n_16278, n_16279, n_16280, n_16281, n_16282,
       n_16283;
  wire n_16284, n_16285, n_16286, n_16287, n_16288, n_16293, n_16294,
       n_16295;
  wire n_16296, n_16297, n_16298, n_16299, n_16300, n_16301, n_16302,
       n_16303;
  wire n_16304, n_16305, n_16306, n_16307, n_16308, n_16309, n_16310,
       n_16311;
  wire n_16312, n_16313, n_16314, n_16315, n_16316, n_16317, n_16318,
       n_16319;
  wire n_16320, n_16321, n_16322, n_16323, n_16324, n_16325, n_16326,
       n_16327;
  wire n_16328, n_16329, n_16330, n_16331, n_16332, n_16333, n_16334,
       n_16335;
  wire n_16336, n_16337, n_16338, n_16339, n_16340, n_16341, n_16342,
       n_16343;
  wire n_16344, n_16345, n_16346, n_16347, n_16348, n_16349, n_16350,
       n_16351;
  wire n_16352, n_16353, n_16354, n_16355, n_16356, n_16357, n_16358,
       n_16359;
  wire n_16360, n_16361, n_16362, n_16363, n_16364, n_16365, n_16366,
       n_16367;
  wire n_16368, n_16369, n_16370, n_16371, n_16372, n_16373, n_16374,
       n_16375;
  wire n_16376, n_16377, n_16378, n_16379, n_16380, n_16381, n_16382,
       n_16383;
  wire n_16384, n_16385, n_16386, n_16387, n_16388, n_16389, n_16390,
       n_16391;
  wire n_16392, n_16393, n_16394, n_16395, n_16396, n_16397, n_16398,
       n_16399;
  wire n_16400, n_16401, n_16402, n_16403, n_16404, n_16405, n_16406,
       n_16407;
  wire n_16408, n_16409, n_16410, n_16411, n_16412, n_16413, n_16414,
       n_16415;
  wire n_16416, n_16417, n_16418, n_16419, n_16420, n_16421, n_16422,
       n_16423;
  wire n_16428, n_16429, n_16430, n_16431, n_16432, n_16433, n_16434,
       n_16435;
  wire n_16436, n_16437, n_16442, n_16443, n_16444, n_16445, n_16446,
       n_16447;
  wire n_16448, n_16449, n_16450, n_16451, n_16452, n_16453, n_16454,
       n_16455;
  wire n_16456, n_16457, n_16458, n_16459, n_16460, n_16461, n_16462,
       n_16463;
  wire n_16464, n_16465, n_16466, n_16467, n_16468, n_16469, n_16470,
       n_16471;
  wire n_16472, n_16473, n_16474, n_16475, n_16476, n_16477, n_16478,
       n_16479;
  wire n_16480, n_16481, n_16482, n_16487, n_16488, n_16489, n_16490,
       n_16491;
  wire n_16492, n_16493, n_16494, n_16495, n_16496, n_16501, n_16502,
       n_16503;
  wire n_16504, n_16505, n_16506, n_16507, n_16508, n_16509, n_16510,
       n_16511;
  wire n_16516, n_16517, n_16518, n_16519, n_16520, n_16521, n_16522,
       n_16523;
  wire n_16524, n_16525, n_16526, n_16527, n_16528, n_16529, n_16530,
       n_16531;
  wire n_16532, n_16533, n_16534, n_16535, n_16536, n_16537, n_16538,
       n_16539;
  wire n_16540, n_16541, n_16542, n_16543, n_16544, n_16545, n_16546,
       n_16547;
  wire n_16548, n_16549, n_16550, n_16551, n_16552, n_16553, n_16554,
       n_16555;
  wire n_16556, n_16561, n_16562, n_16563, n_16564, n_16565, n_16566,
       n_16567;
  wire n_16568, n_16569, n_16570, n_16575, n_16576, n_16577, n_16578,
       n_16579;
  wire n_16580, n_16581, n_16582, n_16583, n_16584, n_16585, n_16590,
       n_16591;
  wire n_16592, n_16593, n_16594, n_16595, n_16596, n_16597, n_16598,
       n_16599;
  wire n_16600, n_16601, n_16602, n_16603, n_16604, n_16605, n_16606,
       n_16607;
  wire n_16608, n_16609, n_16610, n_16611, n_16612, n_16613, n_16614,
       n_16615;
  wire n_16616, n_16617, n_16618, n_16619, n_16620, n_16621, n_16622,
       n_16623;
  wire n_16624, n_16625, n_16626, n_16627, n_16628, n_16629, n_16630,
       n_16631;
  wire n_16636, n_16637, n_16638, n_16639, n_16640, n_16641, n_16642,
       n_16643;
  wire n_16644, n_16645, n_16646, n_16647, n_16648, n_16649, n_16650,
       n_16651;
  wire n_16652, n_16653, n_16654, n_16655, n_16656, n_16657, n_16662,
       n_16663;
  wire n_16664, n_16665, n_16666, n_16667, n_16668, n_16669, n_16670,
       n_16671;
  wire n_16672, n_16673, n_16674, n_16675, n_16676, n_16677, n_16678,
       n_16679;
  wire n_16680, n_16681, n_16682, n_16683, n_16684, n_16685, n_16686,
       n_16687;
  wire n_16688, n_16689, n_16690, n_16691, n_16692, n_16693, n_16694,
       n_16695;
  wire n_16696, n_16697, n_16698, n_16699, n_16700, n_16701, n_16702,
       n_16703;
  wire n_16704, n_16709, n_16710, n_16711, n_16712, n_16713, n_16714,
       n_16715;
  wire n_16716, n_16717, n_16718, n_16719, n_16720, n_16721, n_16722,
       n_16723;
  wire n_16724, n_16725, n_16726, n_16727, n_16728, n_16729, n_16730,
       n_16731;
  wire n_16732, n_16733, n_16734, n_16735, n_16736, n_16737, n_16738,
       n_16739;
  wire n_16740, n_16741, n_16742, n_16743, n_16744, n_16745, n_16746,
       n_16747;
  wire n_16748, n_16749, n_16750, n_16751, n_16752, n_16753, n_16754,
       n_16755;
  wire n_16756, n_16757, n_16758, n_16759, n_16760, n_16761, n_16762,
       n_16763;
  wire n_16764, n_16765, n_16766, n_16767, n_16768, n_16769, n_16770,
       n_16771;
  wire n_16772, n_16773, n_16774, n_16775, n_16776, n_16777, n_16778,
       n_16779;
  wire n_16780, n_16781, n_16782, n_16783, n_16784, n_16785, n_16786,
       n_16787;
  wire n_16788, n_16789, n_16790, n_16791, n_16792, n_16793, n_16794,
       n_16795;
  wire n_16796, n_16797, n_16798, n_16799, n_16800, n_16801, n_16802,
       n_16803;
  wire n_16804, n_16805, n_16806, n_16807, n_16808, n_16809, n_16810,
       n_16811;
  wire n_16812, n_16813, n_16814, n_16815, n_16816, n_16817, n_16818,
       n_16819;
  wire n_16820, n_16821, n_16822, n_16823, n_16827, n_16829, n_16830,
       n_16831;
  wire n_16832, n_16837, n_16838, n_16839, n_16840, n_16845, n_16846,
       n_16847;
  wire n_16848, n_16853, n_16854, n_16855, n_16856, n_16861, n_16862,
       n_16863;
  wire n_16864, n_16865, n_16866, n_16867, n_16868, n_16869, n_16870,
       n_16871;
  wire n_16872, n_16873, n_16874, n_16875, n_16876, n_16877, n_16878,
       n_16879;
  wire n_16880, n_16881, n_16882, n_16883, n_16884, n_16885, n_16886,
       n_16887;
  wire n_16888, n_16889, n_16890, n_16891, n_16892, n_16893, n_16894,
       n_16895;
  wire n_16896, n_16897, n_16898, n_16899, n_16900, n_16901, n_16902,
       n_16903;
  wire n_16904, n_16905, n_16906, n_16907, n_16908, n_16909, n_16910,
       n_16911;
  wire n_16912, n_16913, n_16914, n_16915, n_16916, n_16917, n_16918,
       n_16919;
  wire n_16920, n_16921, n_16922, n_16923, n_16924, n_16925, n_16926,
       n_16927;
  wire n_16928, n_16929, n_16930, n_16931, n_16932, n_16933, n_16934,
       n_16935;
  wire n_16936, n_16937, n_16938, n_16939, n_16940, n_16941, n_16942,
       n_16943;
  wire n_16944, n_16945, n_16946, n_16947, n_16948, n_16949, n_16950,
       n_16951;
  wire n_16952, n_16953, n_16954, n_16955, n_16956, n_16957, n_16958,
       n_16959;
  wire n_16960, n_16961, n_16962, n_16963, n_16964, n_16965, n_16966,
       n_16967;
  wire n_16968, n_16969, n_16970, n_16971, n_16972, n_16973, n_16974,
       n_16975;
  wire n_16976, n_16977, n_16978, n_16979, n_16980, n_16981, n_16985,
       n_16986;
  wire n_16988, n_16989, n_16990, n_16991, n_16992, n_16993, n_16994,
       n_16995;
  wire n_16996, n_16997, n_16998, n_17002, n_17003, n_17004, n_17006,
       n_17007;
  wire n_17008, n_17009, n_17010, n_17011, n_17012, n_17013, n_17014,
       n_17015;
  wire n_17016, n_17020, n_17022, n_17023, n_17024, n_17025, n_17026,
       n_17027;
  wire n_17028, n_17029, n_17030, n_17031, n_17032, n_17033, n_17034,
       n_17035;
  wire n_17036, n_17037, n_17038, n_17039, n_17040, n_17041, n_17042,
       n_17043;
  wire n_17044, n_17045, n_17046, n_17047, n_17048, n_17049, n_17050,
       n_17051;
  wire n_17052, n_17057, n_17058, n_17059, n_17060, n_17061, n_17062,
       n_17063;
  wire n_17064, n_17065, n_17066, n_17071, n_17072, n_17073, n_17074,
       n_17075;
  wire n_17076, n_17077, n_17078, n_17079, n_17080, n_17081, n_17086,
       n_17087;
  wire n_17088, n_17089, n_17090, n_17091, n_17092, n_17093, n_17094,
       n_17095;
  wire n_17096, n_17097, n_17098, n_17099, n_17100, n_17101, n_17102,
       n_17103;
  wire n_17104, n_17105, n_17106, n_17107, n_17108, n_17109, n_17110,
       n_17111;
  wire n_17112, n_17113, n_17114, n_17115, n_17116, n_17117, n_17118,
       n_17119;
  wire n_17120, n_17121, n_17122, n_17123, n_17124, n_17125, n_17126,
       n_17131;
  wire n_17132, n_17133, n_17134, n_17135, n_17136, n_17137, n_17138,
       n_17139;
  wire n_17140, n_17145, n_17146, n_17147, n_17148, n_17149, n_17150,
       n_17151;
  wire n_17152, n_17153, n_17154, n_17155, n_17160, n_17161, n_17162,
       n_17163;
  wire n_17164, n_17165, n_17166, n_17167, n_17168, n_17169, n_17170,
       n_17171;
  wire n_17172, n_17173, n_17174, n_17175, n_17176, n_17177, n_17178,
       n_17179;
  wire n_17180, n_17181, n_17182, n_17183, n_17184, n_17185, n_17186,
       n_17187;
  wire n_17188, n_17189, n_17190, n_17191, n_17192, n_17193, n_17194,
       n_17195;
  wire n_17196, n_17197, n_17198, n_17199, n_17200, n_17205, n_17206,
       n_17207;
  wire n_17208, n_17209, n_17210, n_17211, n_17212, n_17213, n_17214,
       n_17219;
  wire n_17220, n_17221, n_17222, n_17223, n_17224, n_17225, n_17226,
       n_17227;
  wire n_17228, n_17229, n_17234, n_17235, n_17236, n_17237, n_17238,
       n_17239;
  wire n_17240, n_17241, n_17242, n_17243, n_17244, n_17245, n_17246,
       n_17247;
  wire n_17248, n_17249, n_17250, n_17251, n_17252, n_17253, n_17254,
       n_17255;
  wire n_17256, n_17257, n_17258, n_17259, n_17260, n_17261, n_17262,
       n_17263;
  wire n_17264, n_17265, n_17266, n_17267, n_17268, n_17269, n_17270,
       n_17271;
  wire n_17272, n_17273, n_17274, n_17275, n_17280, n_17281, n_17282,
       n_17283;
  wire n_17284, n_17285, n_17286, n_17287, n_17288, n_17289, n_17290,
       n_17291;
  wire n_17292, n_17293, n_17294, n_17295, n_17296, n_17297, n_17298,
       n_17299;
  wire n_17300, n_17301, n_17306, n_17307, n_17308, n_17309, n_17310,
       n_17311;
  wire n_17312, n_17313, n_17314, n_17315, n_17316, n_17317, n_17318,
       n_17319;
  wire n_17320, n_17321, n_17322, n_17323, n_17324, n_17325, n_17326,
       n_17327;
  wire n_17328, n_17329, n_17330, n_17331, n_17332, n_17333, n_17334,
       n_17335;
  wire n_17336, n_17337, n_17338, n_17339, n_17340, n_17341, n_17342,
       n_17343;
  wire n_17344, n_17345, n_17346, n_17347, n_17348, n_17353, n_17354,
       n_17355;
  wire n_17356, n_17357, n_17358, n_17359, n_17360, n_17361, n_17362,
       n_17363;
  wire n_17364, n_17365, n_17366, n_17367, n_17368, n_17369, n_17370,
       n_17371;
  wire n_17372, n_17373, n_17374, n_17375, n_17376, n_17377, n_17378,
       n_17379;
  wire n_17380, n_17381, n_17382, n_17383, n_17384, n_17385, n_17386,
       n_17387;
  wire n_17388, n_17389, n_17390, n_17391, n_17392, n_17393, n_17394,
       n_17395;
  wire n_17396, n_17397, n_17398, n_17399, n_17400, n_17401, n_17402,
       n_17403;
  wire n_17404, n_17405, n_17406, n_17407, n_17408, n_17409, n_17410,
       n_17411;
  wire n_17412, n_17413, n_17414, n_17415, n_17416, n_17417, n_17418,
       n_17419;
  wire n_17420, n_17421, n_17422, n_17423, n_17424, n_17425, n_17426,
       n_17427;
  wire n_17428, n_17429, n_17430, n_17431, n_17432, n_17433, n_17434,
       n_17435;
  wire n_17436, n_17437, n_17438, n_17439, n_17440, n_17441, n_17442,
       n_17443;
  wire n_17444, n_17445, n_17446, n_17447, n_17448, n_17449, n_17450,
       n_17451;
  wire n_17452, n_17453, n_17454, n_17455, n_17456, n_17457, n_17458,
       n_17459;
  wire n_17460, n_17461, n_17462, n_17463, n_17464, n_17465, n_17466,
       n_17467;
  wire n_17468, n_17469, n_17470, n_17471, n_17472, n_17473, n_17474,
       n_17475;
  wire n_17476, n_17477, n_17478, n_17479, n_17480, n_17485, n_17486,
       n_17487;
  wire n_17488, n_17489, n_17490, n_17491, n_17492, n_17493, n_17494,
       n_17495;
  wire n_17496, n_17497, n_17498, n_17499, n_17500, n_17501, n_17502,
       n_17503;
  wire n_17504, n_17505, n_17506, n_17507, n_17508, n_17513, n_17514,
       n_17515;
  wire n_17516, n_17517, n_17518, n_17523, n_17524, n_17525, n_17526,
       n_17527;
  wire n_17528, n_17529, n_17530, n_17531, n_17532, n_17533, n_17534,
       n_17535;
  wire n_17536, n_17537, n_17538, n_17539, n_17540, n_17541, n_17542,
       n_17543;
  wire n_17544, n_17545, n_17546, n_17547, n_17552, n_17553, n_17554,
       n_17555;
  wire n_17556, n_17557, n_17558, n_17559, n_17560, n_17561, n_17562,
       n_17563;
  wire n_17564, n_17565, n_17566, n_17567, n_17568, n_17569, n_17570,
       n_17571;
  wire n_17572, n_17573, n_17574, n_17575, n_17576, n_17577, n_17578,
       n_17579;
  wire n_17580, n_17581, n_17586, n_17587, n_17588, n_17589, n_17590,
       n_17591;
  wire n_17592, n_17593, n_17594, n_17595, n_17596, n_17597, n_17598,
       n_17599;
  wire n_17600, n_17601, n_17602, n_17603, n_17604, n_17605, n_17610,
       n_17611;
  wire n_17612, n_17613, n_17614, n_17615, n_17616, n_17617, n_17618,
       n_17619;
  wire n_17620, n_17621, n_17622, n_17623, n_17624, n_17625, n_17626,
       n_17627;
  wire n_17628, n_17629, n_17630, n_17631, n_17632, n_17633, n_17634,
       n_17635;
  wire n_17636, n_17637, n_17638, n_17639, n_17640, n_17641, n_17642,
       n_17643;
  wire n_17644, n_17645, n_17646, n_17647, n_17648, n_17649, n_17650,
       n_17651;
  wire n_17652, n_17653, n_17654, n_17655, n_17656, n_17657, n_17658,
       n_17659;
  wire n_17660, n_17661, n_17662, n_17663, n_17664, n_17665, n_17666,
       n_17667;
  wire n_17668, n_17669, n_17670, n_17671, n_17672, n_17673, n_17674,
       n_17675;
  wire n_17676, n_17683, n_17688, n_17689, n_17690, n_17691, n_17692,
       n_17693;
  wire n_17694, n_17695, n_17696, n_17697, n_17698, n_17699, n_17700,
       n_17701;
  wire n_17702, n_17703, n_17704, n_17705, n_17706, n_17707, n_17708,
       n_17709;
  wire n_17710, n_17711, n_17716, n_17717, n_17718, n_17719, n_17720,
       n_17721;
  wire n_17722, n_17723, n_17724, n_17725, n_17726, n_17727, n_17728,
       n_17729;
  wire n_17730, n_17731, n_17732, n_17733, n_17734, n_17735, n_17736,
       n_17737;
  wire n_17738, n_17743, n_17744, n_17745, n_17746, n_17747, n_17748,
       n_17749;
  wire n_17750, n_17751, n_17752, n_17753, n_17754, n_17755, n_17756,
       n_17757;
  wire n_17758, n_17759, n_17760, n_17761, n_17762, n_17763, n_17764,
       n_17765;
  wire n_17766, n_17767, n_17768, n_17769, n_17770, n_17771, n_17772,
       n_17773;
  wire n_17774, n_17775, n_17776, n_17777, n_17778, n_17779, n_17780,
       n_17781;
  wire n_17782, n_17783, n_17784, n_17785, n_17786, n_17787, n_17788,
       n_17789;
  wire n_17790, n_17791, n_17792, n_17793, n_17794, n_17795, n_17800,
       n_17801;
  wire n_17802, n_17803, n_17804, n_17805, n_17806, n_17807, n_17808,
       n_17809;
  wire n_17814, n_17815, n_17816, n_17817, n_17818, n_17819, n_17820,
       n_17821;
  wire n_17822, n_17827, n_17828, n_17829, n_17830, n_17831, n_17832,
       n_17833;
  wire n_17834, n_17835, n_17836, n_17837, n_17838, n_17839, n_17840,
       n_17841;
  wire n_17842, n_17843, n_17844, n_17845, n_17846, n_17847, n_17848,
       n_17849;
  wire n_17850, n_17851, n_17852, n_17853, n_17854, n_17855, n_17856,
       n_17857;
  wire n_17858, n_17859, n_17860, n_17861, n_17862, n_17863, n_17864,
       n_17865;
  wire n_17866, n_17867, n_17868, n_17869, n_17870, n_17871, n_17872,
       n_17873;
  wire n_17874, n_17875, n_17876, n_17877, n_17878, n_17883, n_17884,
       n_17885;
  wire n_17886, n_17887, n_17888, n_17889, n_17890, n_17891, n_17892,
       n_17897;
  wire n_17898, n_17899, n_17900, n_17901, n_17902, n_17903, n_17904,
       n_17905;
  wire n_17910, n_17911, n_17912, n_17913, n_17914, n_17915, n_17916,
       n_17917;
  wire n_17918, n_17919, n_17920, n_17921, n_17922, n_17923, n_17924,
       n_17925;
  wire n_17926, n_17927, n_17928, n_17929, n_17930, n_17931, n_17932,
       n_17933;
  wire n_17934, n_17935, n_17936, n_17937, n_17938, n_17939, n_17940,
       n_17941;
  wire n_17942, n_17943, n_17944, n_17945, n_17946, n_17947, n_17948,
       n_17949;
  wire n_17950, n_17951, n_17952, n_17953, n_17954, n_17955, n_17956,
       n_17957;
  wire n_17958, n_17959, n_17960, n_17961, n_17966, n_17967, n_17968,
       n_17969;
  wire n_17970, n_17971, n_17972, n_17973, n_17974, n_17975, n_17980,
       n_17981;
  wire n_17982, n_17983, n_17984, n_17985, n_17986, n_17987, n_17988,
       n_17993;
  wire n_17994, n_17995, n_17996, n_17997, n_17998, n_17999, n_18000,
       n_18001;
  wire n_18002, n_18003, n_18004, n_18005, n_18006, n_18007, n_18008,
       n_18009;
  wire n_18010, n_18011, n_18012, n_18013, n_18014, n_18015, n_18016,
       n_18017;
  wire n_18018, n_18019, n_18020, n_18021, n_18022, n_18023, n_18024,
       n_18025;
  wire n_18026, n_18027, n_18028, n_18029, n_18030, n_18031, n_18032,
       n_18033;
  wire n_18034, n_18035, n_18036, n_18037, n_18038, n_18039, n_18040,
       n_18041;
  wire n_18042, n_18043, n_18044, n_18049, n_18050, n_18051, n_18052,
       n_18053;
  wire n_18054, n_18055, n_18056, n_18057, n_18062, n_18063, n_18064,
       n_18065;
  wire n_18066, n_18067, n_18068, n_18069, n_18070, n_18071, n_18072,
       n_18073;
  wire n_18074, n_18075, n_18076, n_18077, n_18078, n_18079, n_18080,
       n_18081;
  wire n_18082, n_18083, n_18084, n_18085, n_18086, n_18087, n_18088,
       n_18089;
  wire n_18090, n_18091, n_18092, n_18093, n_18094, n_18095, n_18096,
       n_18097;
  wire n_18098, n_18099, n_18100, n_18101, n_18102, n_18103, n_18104,
       n_18105;
  wire n_18106, n_18107, n_18108, n_18109, n_18110, n_18111, n_18112,
       n_18113;
  wire n_18114, n_18115, n_18116, n_18117, n_18118, n_18119, n_18120,
       n_18124;
  wire n_18126, n_18127, n_18128, n_18129, n_18133, n_18135, n_18136,
       n_18137;
  wire n_18138, n_18142, n_18144, n_18145, n_18146, n_18147, n_18151,
       n_18153;
  wire n_18154, n_18155, n_18156, n_18161, n_18162, n_18163, n_18164,
       n_18169;
  wire n_18170, n_18171, n_18172, n_18173, n_18174, n_18175, n_18176,
       n_18177;
  wire n_18178, n_18179, n_18180, n_18181, n_18182, n_18183, n_18184,
       n_18185;
  wire n_18186, n_18187, n_18188, n_18189, n_18190, n_18191, n_18192,
       n_18193;
  wire n_18194, n_18195, n_18196, n_18197, n_18198, n_18199, n_18200,
       n_18201;
  wire n_18202, n_18203, n_18204, n_18205, n_18206, n_18207, n_18208,
       n_18209;
  wire n_18210, n_18211, n_18212, n_18213, n_18214, n_18215, n_18216,
       n_18217;
  wire n_18218, n_18219, n_18220, n_18221, n_18222, n_18223, n_18224,
       n_18225;
  wire n_18226, n_18227, n_18228, n_18229, n_18230, n_18231, n_18232,
       n_18233;
  wire n_18234, n_18235, n_18236, n_18237, n_18238, n_18239, n_18240,
       n_18241;
  wire n_18242, n_18243, n_18244, n_18245, n_18246, n_18247, n_18248,
       n_18249;
  wire n_18250, n_18251, n_18252, n_18253, n_18254, n_18255, n_18256,
       n_18257;
  wire n_18258, n_18259, n_18260, n_18261, n_18262, n_18263, n_18264,
       n_18265;
  wire n_18266, n_18267, n_18268, n_18269, n_18270, n_18271, n_18272,
       n_18273;
  wire n_18274, n_18275, n_18276, n_18277, n_18278, n_18279, n_18280,
       n_18281;
  wire n_18282, n_18283, n_18284, n_18285, n_18286, n_18287, n_18288,
       n_18289;
  wire n_18290, n_18291, n_18292, n_18297, n_18298, n_18299, n_18300,
       n_18301;
  wire n_18302, n_18303, n_18304, n_18305, n_18306, n_18307, n_18308,
       n_18309;
  wire n_18310, n_18311, n_18312, n_18313, n_18314, n_18315, n_18316,
       n_18317;
  wire n_18318, n_18319, n_18320, n_18321, n_18322, n_18323, n_18324,
       n_18325;
  wire n_18326, n_18327, n_18328, n_18329, n_18330, n_18331, n_18332,
       n_18333;
  wire n_18334, n_18335, n_18336, n_18337, n_18338, n_18339, n_18340,
       n_18341;
  wire n_18342, n_18343, n_18344, n_18345, n_18346, n_18347, n_18348,
       n_18349;
  wire n_18350, n_18351, n_18352, n_18353, n_18354, n_18355, n_18359,
       n_18361;
  wire n_18362, n_18363, n_18364, n_18369, n_18370, n_18371, n_18372,
       n_18377;
  wire n_18378, n_18379, n_18380, n_18385, n_18386, n_18387, n_18388,
       n_18393;
  wire n_18394, n_18395, n_18396, n_18397, n_18398, n_18399, n_18400,
       n_18401;
  wire n_18402, n_18403, n_18404, n_18405, n_18406, n_18407, n_18408,
       n_18409;
  wire n_18410, n_18411, n_18412, n_18413, n_18414, n_18415, n_18416,
       n_18417;
  wire n_18418, n_18419, n_18420, n_18421, n_18422, n_18423, n_18424,
       n_18425;
  wire n_18426, n_18427, n_18428, n_18429, n_18430, n_18431, n_18432,
       n_18433;
  wire n_18434, n_18435, n_18436, n_18437, n_18438, n_18439, n_18440,
       n_18441;
  wire n_18442, n_18443, n_18444, n_18445, n_18446, n_18447, n_18448,
       n_18449;
  wire n_18450, n_18451, n_18452, n_18453, n_18454, n_18455, n_18456,
       n_18457;
  wire n_18458, n_18459, n_18460, n_18461, n_18462, n_18463, n_18464,
       n_18465;
  wire n_18466, n_18467, n_18468, n_18469, n_18470, n_18471, n_18472,
       n_18473;
  wire n_18474, n_18475, n_18476, n_18477, n_18478, n_18479, n_18480,
       n_18481;
  wire n_18482, n_18483, n_18484, n_18485, n_18486, n_18487, n_18488,
       n_18489;
  wire n_18490, n_18491, n_18492, n_18493, n_18494, n_18495, n_18496,
       n_18497;
  wire n_18498, n_18499, n_18500, n_18501, n_18502, n_18503, n_18504,
       n_18505;
  wire n_18506, n_18507, n_18508, n_18509, n_18510, n_18511, n_18512,
       n_18513;
  wire n_18514, n_18515, n_18516, n_18517, n_18518, n_18519, n_18520,
       n_18521;
  wire n_18522, n_18523, n_18524, n_18525, n_18526, n_18527, n_18528,
       n_18529;
  wire n_18530, n_18531, n_18532, n_18533, n_18534, n_18535, n_18536,
       n_18537;
  wire n_18538, n_18539, n_18540, n_18541, n_18542, n_18543, n_18548,
       n_18549;
  wire n_18550, n_18551, n_18552, n_18553, n_18554, n_18555, n_18556,
       n_18557;
  wire n_18558, n_18559, n_18560, n_18561, n_18562, n_18563, n_18564,
       n_18565;
  wire n_18566, n_18567, n_18568, n_18569, n_18570, n_18571, n_18572,
       n_18573;
  wire n_18574, n_18575, n_18576, n_18577, n_18578, n_18579, n_18580,
       n_18581;
  wire n_18582, n_18583, n_18584, n_18585, n_18586, n_18587, n_18588,
       n_18589;
  wire n_18590, n_18591, n_18592, n_18596, n_18598, n_18599, n_18600,
       n_18601;
  wire n_18606, n_18607, n_18608, n_18609, n_18614, n_18615, n_18616,
       n_18617;
  wire n_18622, n_18623, n_18624, n_18625, n_18630, n_18631, n_18632,
       n_18633;
  wire n_18634, n_18635, n_18636, n_18637, n_18638, n_18639, n_18640,
       n_18641;
  wire n_18642, n_18643, n_18644, n_18645, n_18646, n_18647, n_18648,
       n_18649;
  wire n_18650, n_18651, n_18652, n_18653, n_18654, n_18655, n_18656,
       n_18657;
  wire n_18658, n_18659, n_18660, n_18661, n_18662, n_18663, n_18664,
       n_18665;
  wire n_18666, n_18667, n_18668, n_18669, n_18670, n_18671, n_18672,
       n_18673;
  wire n_18674, n_18675, n_18676, n_18677, n_18678, n_18679, n_18680,
       n_18681;
  wire n_18682, n_18683, n_18684, n_18685, n_18686, n_18687, n_18688,
       n_18689;
  wire n_18690, n_18691, n_18692, n_18693, n_18694, n_18695, n_18696,
       n_18697;
  wire n_18698, n_18699, n_18700, n_18701, n_18702, n_18703, n_18704,
       n_18705;
  wire n_18706, n_18707, n_18708, n_18709, n_18710, n_18711, n_18712,
       n_18713;
  wire n_18714, n_18715, n_18716, n_18717, n_18718, n_18719, n_18720,
       n_18721;
  wire n_18722, n_18723, n_18724, n_18725, n_18726, n_18727, n_18728,
       n_18729;
  wire n_18730, n_18731, n_18732, n_18733, n_18734, n_18735, n_18736,
       n_18737;
  wire n_18738, n_18739, n_18740, n_18741, n_18742, n_18743, n_18744,
       n_18745;
  wire n_18746, n_18747, n_18748, n_18749, n_18750, n_18751, n_18752,
       n_18753;
  wire n_18754, n_18755, n_18756, n_18757, n_18758, n_18759, n_18760,
       n_18765;
  wire n_18766, n_18767, n_18768, n_18769, n_18770, n_18771, n_18772,
       n_18773;
  wire n_18774, n_18775, n_18776, n_18777, n_18778, n_18779, n_18780,
       n_18781;
  wire n_18782, n_18783, n_18784, n_18785, n_18786, n_18787, n_18788,
       n_18789;
  wire n_18790, n_18791, n_18792, n_18793, n_18794, n_18795, n_18796,
       n_18797;
  wire n_18798, n_18799, n_18800, n_18801, n_18802, n_18803, n_18804,
       n_18805;
  wire n_18806, n_18807, n_18808, n_18809, n_18810, n_18811, n_18812,
       n_18813;
  wire n_18814, n_18815, n_18816, n_18817, n_18818, n_18819, n_18823,
       n_18825;
  wire n_18826, n_18827, n_18828, n_18833, n_18834, n_18835, n_18836,
       n_18841;
  wire n_18842, n_18843, n_18844, n_18849, n_18850, n_18851, n_18852,
       n_18857;
  wire n_18858, n_18859, n_18860, n_18861, n_18862, n_18863, n_18864,
       n_18865;
  wire n_18866, n_18867, n_18868, n_18869, n_18870, n_18871, n_18872,
       n_18873;
  wire n_18874, n_18875, n_18876, n_18877, n_18878, n_18879, n_18880,
       n_18881;
  wire n_18882, n_18883, n_18884, n_18885, n_18886, n_18887, n_18888,
       n_18889;
  wire n_18890, n_18891, n_18892, n_18893, n_18894, n_18895, n_18896,
       n_18897;
  wire n_18898, n_18899, n_18900, n_18901, n_18902, n_18903, n_18904,
       n_18905;
  wire n_18906, n_18907, n_18908, n_18909, n_18910, n_18911, n_18912,
       n_18913;
  wire n_18914, n_18915, n_18916, n_18917, n_18918, n_18919, n_18920,
       n_18921;
  wire n_18922, n_18923, n_18924, n_18925, n_18926, n_18927, n_18928,
       n_18929;
  wire n_18930, n_18931, n_18932, n_18933, n_18934, n_18935, n_18936,
       n_18937;
  wire n_18938, n_18939, n_18940, n_18941, n_18942, n_18943, n_18944,
       n_18945;
  wire n_18946, n_18947, n_18948, n_18949, n_18950, n_18951, n_18952,
       n_18953;
  wire n_18954, n_18955, n_18956, n_18957, n_18958, n_18959, n_18960,
       n_18961;
  wire n_18962, n_18963, n_18964, n_18965, n_18966, n_18967, n_18968,
       n_18969;
  wire n_18970, n_18971, n_18972, n_18973, n_18974, n_18975, n_18976,
       n_18977;
  wire n_18978, n_18979, n_18980, n_18981, n_18982, n_18983, n_18984,
       n_18985;
  wire n_18986, n_18991, n_18992, n_18993, n_18994, n_18995, n_18996,
       n_18997;
  wire n_18998, n_18999, n_19000, n_19001, n_19002, n_19003, n_19004,
       n_19005;
  wire n_19006, n_19007, n_19008, n_19009, n_19010, n_19011, n_19012,
       n_19013;
  wire n_19014, n_19015, n_19016, n_19017, n_19018, n_19019, n_19020,
       n_19021;
  wire n_19022, n_19023, n_19024, n_19025, n_19026, n_19027, n_19028,
       n_19029;
  wire n_19030, n_19031, n_19032, n_19037, n_19038, n_19039, n_19040,
       n_19045;
  wire n_19046, n_19047, n_19048, n_19053, n_19054, n_19055, n_19056,
       n_19061;
  wire n_19062, n_19063, n_19064, n_19065, n_19070, n_19071, n_19072,
       n_19073;
  wire n_19074, n_19075, n_19076, n_19077, n_19078, n_19079, n_19080,
       n_19081;
  wire n_19082, n_19083, n_19084, n_19085, n_19086, n_19087, n_19088,
       n_19089;
  wire n_19090, n_19091, n_19092, n_19093, n_19094, n_19095, n_19096,
       n_19097;
  wire n_19098, n_19099, n_19100, n_19101, n_19102, n_19103, n_19104,
       n_19105;
  wire n_19106, n_19107, n_19108, n_19109, n_19110, n_19111, n_19112,
       n_19113;
  wire n_19114, n_19115, n_19116, n_19117, n_19118, n_19119, n_19120,
       n_19121;
  wire n_19122, n_19123, n_19124, n_19125, n_19126, n_19127, n_19128,
       n_19129;
  wire n_19130, n_19131, n_19132, n_19133, n_19134, n_19135, n_19136,
       n_19137;
  wire n_19138, n_19139, n_19140, n_19141, n_19142, n_19143, n_19144,
       n_19145;
  wire n_19146, n_19147, n_19148, n_19149, n_19150, n_19151, n_19152,
       n_19153;
  wire n_19154, n_19155, n_19156, n_19157, n_19158, n_19159, n_19160,
       n_19161;
  wire n_19162, n_19163, n_19164, n_19165, n_19166, n_19167, n_19168,
       n_19169;
  wire n_19170, n_19171, n_19172, n_19173, n_19174, n_19175, n_19176,
       n_19177;
  wire n_19178, n_19179, n_19180, n_19181, n_19182, n_19183, n_19184,
       n_19185;
  wire n_19186, n_19187, n_19188, n_19189, n_19190, n_19191, n_19192,
       n_19193;
  wire n_19194, n_19195, n_19196, n_19197, n_19198, n_19199, n_19200,
       n_19201;
  wire n_19202, n_19203, n_19204, n_19205, n_19206, n_19207, n_19208,
       n_19209;
  wire n_19210, n_19211, n_19212, n_19213, n_19214, n_19215, n_19216,
       n_19217;
  wire n_19218, n_19219, n_19220, n_19221, n_19222, n_19223, n_19224,
       n_19225;
  wire n_19226, n_19227, n_19228, n_19229, n_19230, n_19231, n_19232,
       n_19233;
  wire n_19234, n_19235, n_19236, n_19237, n_19238, n_19239, n_19240,
       n_19241;
  wire n_19242, n_19247, n_19248, n_19249, n_19250, n_19255, n_19256,
       n_19257;
  wire n_19258, n_19263, n_19264, n_19265, n_19266, n_19271, n_19272,
       n_19273;
  wire n_19274, n_19279, n_19280, n_19281, n_19282, n_19283, n_19284,
       n_19285;
  wire n_19286, n_19287, n_19288, n_19289, n_19290, n_19291, n_19292,
       n_19293;
  wire n_19294, n_19295, n_19296, n_19297, n_19298, n_19299, n_19300,
       n_19301;
  wire n_19302, n_19303, n_19304, n_19305, n_19306, n_19307, n_19308,
       n_19309;
  wire n_19310, n_19311, n_19312, n_19313, n_19314, n_19315, n_19316,
       n_19317;
  wire n_19318, n_19319, n_19320, n_19321, n_19322, n_19323, n_19324,
       n_19325;
  wire n_19326, n_19327, n_19328, n_19329, n_19330, n_19331, n_19332,
       n_19333;
  wire n_19334, n_19335, n_19336, n_19337, n_19338, n_19339, n_19340,
       n_19341;
  wire n_19342, n_19343, n_19344, n_19345, n_19346, n_19347, n_19348,
       n_19349;
  wire n_19350, n_19351, n_19352, n_19353, n_19354, n_19355, n_19356,
       n_19357;
  wire n_19358, n_19359, n_19360, n_19361, n_19362, n_19363, n_19364,
       n_19365;
  wire n_19366, n_19367, n_19368, n_19369, n_19370, n_19371, n_19372,
       n_19373;
  wire n_19374, n_19375, n_19376, n_19377, n_19378, n_19379, n_19380,
       n_19381;
  wire n_19382, n_19383, n_19384, n_19385, n_19386, n_19387, n_19388,
       n_19389;
  wire n_19390, n_19391, n_19392, n_19393, n_19394, n_19395, n_19396,
       n_19397;
  wire n_19398, n_19399, n_19400, n_19401, n_19402, n_19403, n_19404,
       n_19405;
  wire n_19406, n_19407, n_19408, n_19409, n_19410, n_19411, n_19412,
       n_19413;
  wire n_19414, n_19415, n_19416, n_19417, n_19418, n_19419, n_19420,
       n_19421;
  wire n_19422, n_19423, n_19424, n_19425, n_19426, n_19427, n_19428,
       n_19429;
  wire n_19430, n_19431, n_19432, n_19433, n_19434, n_19435, n_19436,
       n_19437;
  wire n_19438, n_19439, n_19440, n_19441, n_19442, n_19446, n_19448,
       n_19449;
  wire n_19450, n_19451, n_19456, n_19457, n_19458, n_19459, n_19464,
       n_19465;
  wire n_19466, n_19467, n_19472, n_19473, n_19474, n_19475, n_19480,
       n_19481;
  wire n_19482, n_19483, n_19484, n_19485, n_19486, n_19487, n_19488,
       n_19489;
  wire n_19490, n_19491, n_19492, n_19493, n_19494, n_19495, n_19496,
       n_19497;
  wire n_19498, n_19499, n_19500, n_19501, n_19502, n_19503, n_19504,
       n_19505;
  wire n_19506, n_19507, n_19508, n_19509, n_19510, n_19511, n_19512,
       n_19513;
  wire n_19514, n_19515, n_19516, n_19517, n_19518, n_19519, n_19520,
       n_19521;
  wire n_19522, n_19523, n_19524, n_19525, n_19526, n_19527, n_19528,
       n_19529;
  wire n_19530, n_19531, n_19532, n_19533, n_19534, n_19535, n_19536,
       n_19537;
  wire n_19538, n_19539, n_19540, n_19541, n_19542, n_19543, n_19544,
       n_19545;
  wire n_19546, n_19547, n_19548, n_19549, n_19550, n_19551, n_19552,
       n_19553;
  wire n_19554, n_19555, n_19556, n_19557, n_19558, n_19559, n_19560,
       n_19561;
  wire n_19562, n_19563, n_19564, n_19565, n_19566, n_19567, n_19568,
       n_19569;
  wire n_19570, n_19571, n_19572, n_19573, n_19574, n_19575, n_19576,
       n_19577;
  wire n_19578, n_19579, n_19580, n_19581, n_19582, n_19583, n_19584,
       n_19585;
  wire n_19586, n_19587, n_19588, n_19589, n_19590, n_19591, n_19592,
       n_19593;
  wire n_19594, n_19595, n_19596, n_19597, n_19598, n_19599, n_19600,
       n_19601;
  wire n_19602, n_19603, n_19604, n_19605, n_19606, n_19607, n_19608,
       n_19609;
  wire n_19610, n_19611, n_19612, n_19613, n_19614, n_19615, n_19616,
       n_19617;
  wire n_19618, n_19619, n_19620, n_19621, n_19626, n_19627, n_19628,
       n_19629;
  wire n_19630, n_19631, n_19632, n_19633, n_19634, n_19635, n_19636,
       n_19637;
  wire n_19638, n_19639, n_19640, n_19641, n_19642, n_19643, n_19644,
       n_19645;
  wire n_19646, n_19647, n_19648, n_19649, n_19650, n_19651, n_19652,
       n_19653;
  wire n_19654, n_19655, n_19656, n_19661, n_19662, n_19663, n_19664,
       n_19665;
  wire n_19666, n_19667, n_19668, n_19669, n_19670, n_19671, n_19672,
       n_19677;
  wire n_19678, n_19679, n_19680, n_19681, n_19682, n_19683, n_19684,
       n_19685;
  wire n_19686, n_19687, n_19688, n_19693, n_19694, n_19695, n_19696,
       n_19697;
  wire n_19698, n_19699, n_19700, n_19701, n_19702, n_19703, n_19704,
       n_19709;
  wire n_19710, n_19711, n_19712, n_19713, n_19714, n_19715, n_19716,
       n_19717;
  wire n_19718, n_19719, n_19720, n_19725, n_19726, n_19727, n_19728,
       n_19729;
  wire n_19730, n_19731, n_19732, n_19733, n_19734, n_19735, n_19736,
       n_19741;
  wire n_19742, n_19743, n_19744, n_19745, n_19746, n_19747, n_19748,
       n_19749;
  wire n_19750, n_19751, n_19752, n_19757, n_19758, n_19759, n_19760,
       n_19761;
  wire n_19762, n_19763, n_19764, n_19765, n_19766, n_19767, n_19768,
       n_19773;
  wire n_19774, n_19775, n_19776, n_19777, n_19778, n_19779, n_19780,
       n_19781;
  wire n_19782, n_19783, n_19784, n_19785, n_19786, n_19787, n_19788,
       n_19789;
  wire n_19790, n_19791, n_19792, n_19793, n_19794, n_19795, n_19796,
       n_19797;
  wire n_19798, n_19803, n_19804, n_19805, n_19806, n_19807, n_19808,
       n_19809;
  wire n_19810, n_19811, n_19816, n_19817, n_19818, n_19819, n_19820,
       n_19821;
  wire n_19822, n_19823, n_19828, n_19829, n_19830, n_19831, n_19832,
       n_19833;
  wire n_19834, n_19835, n_19836, n_19837, n_19838, n_19839, n_19840,
       n_19845;
  wire n_19846, n_19847, n_19848, n_19849, n_19850, n_19851, n_19852,
       n_19853;
  wire n_19854, n_19855, n_19856, n_19861, n_19862, n_19863, n_19864,
       n_19865;
  wire n_19866, n_19867, n_19868, n_19869, n_19870, n_19871, n_19872,
       n_19877;
  wire n_19878, n_19879, n_19880, n_19881, n_19882, n_19883, n_19884,
       n_19885;
  wire n_19886, n_19887, n_19888, n_19893, n_19894, n_19895, n_19896,
       n_19897;
  wire n_19898, n_19899, n_19900, n_19901, n_19902, n_19903, n_19904,
       n_19909;
  wire n_19910, n_19911, n_19912, n_19913, n_19914, n_19915, n_19916,
       n_19917;
  wire n_19918, n_19919, n_19920, n_19925, n_19926, n_19927, n_19928,
       n_19929;
  wire n_19930, n_19931, n_19932, n_19933, n_19934, n_19935, n_19936,
       n_19940;
  wire n_19942, n_19943, n_19944, n_19945, n_19946, n_19947, n_19948,
       n_19949;
  wire n_19950, n_19951, n_19952, n_19953, n_19954, n_19955, n_19956,
       n_19957;
  wire n_19958, n_19959, n_19960, n_19961, n_19962, n_19963, n_19964,
       n_19965;
  wire n_19966, n_19967, n_19972, n_19973, n_19974, n_19975, n_19976,
       n_19977;
  wire n_19978, n_19979, n_19980, n_19985, n_19986, n_19987, n_19988,
       n_19989;
  wire n_19990, n_19991, n_19992, n_19997, n_19998, n_19999, n_20000,
       n_20001;
  wire n_20002, n_20003, n_20004, n_20005, n_20006, n_20007, n_20008,
       n_20009;
  wire n_20014, n_20015, n_20016, n_20017, n_20018, n_20019, n_20020,
       n_20021;
  wire n_20022, n_20023, n_20024, n_20025, n_20030, n_20031, n_20032,
       n_20033;
  wire n_20034, n_20035, n_20036, n_20037, n_20038, n_20039, n_20040,
       n_20041;
  wire n_20046, n_20047, n_20048, n_20049, n_20050, n_20051, n_20052,
       n_20053;
  wire n_20054, n_20055, n_20056, n_20057, n_20062, n_20063, n_20064,
       n_20065;
  wire n_20066, n_20067, n_20068, n_20069, n_20070, n_20071, n_20072,
       n_20073;
  wire n_20078, n_20079, n_20080, n_20081, n_20082, n_20083, n_20084,
       n_20085;
  wire n_20086, n_20087, n_20088, n_20089, n_20094, n_20095, n_20096,
       n_20097;
  wire n_20098, n_20099, n_20100, n_20101, n_20102, n_20103, n_20104,
       n_20105;
  wire n_20106, n_20107, n_20108, n_20109, n_20110, n_20111, n_20112,
       n_20113;
  wire n_20114, n_20115, n_20116, n_20117, n_20118, n_20119, n_20120,
       n_20121;
  wire n_20122, n_20123, n_20124, n_20125, n_20126, n_20127, n_20128,
       n_20129;
  wire n_20130, n_20131, n_20132, n_20133, n_20134, n_20135, n_20136,
       n_20137;
  wire n_20138, n_20139, n_20140, n_20141, n_20146, n_20147, n_20148,
       n_20149;
  wire n_20150, n_20151, n_20152, n_20153, n_20158, n_20159, n_20160,
       n_20161;
  wire n_20162, n_20163, n_20164, n_20165, n_20170, n_20171, n_20172,
       n_20173;
  wire n_20174, n_20175, n_20176, n_20177, n_20178, n_20179, n_20180,
       n_20181;
  wire n_20182, n_20187, n_20188, n_20189, n_20190, n_20191, n_20192,
       n_20193;
  wire n_20194, n_20195, n_20196, n_20197, n_20198, n_20203, n_20204,
       n_20205;
  wire n_20206, n_20207, n_20208, n_20209, n_20210, n_20211, n_20212,
       n_20213;
  wire n_20214, n_20219, n_20220, n_20221, n_20222, n_20223, n_20224,
       n_20225;
  wire n_20226, n_20227, n_20228, n_20229, n_20230, n_20235, n_20236,
       n_20237;
  wire n_20238, n_20239, n_20240, n_20241, n_20242, n_20243, n_20244,
       n_20245;
  wire n_20246, n_20247, n_20252, n_20253, n_20254, n_20255, n_20256,
       n_20257;
  wire n_20258, n_20259, n_20260, n_20261, n_20262, n_20263, n_20268,
       n_20269;
  wire n_20270, n_20271, n_20272, n_20273, n_20274, n_20275, n_20276,
       n_20277;
  wire n_20278, n_20279, n_20280, n_20281, n_20282, n_20283, n_20284,
       n_20285;
  wire n_20286, n_20287, n_20288, n_20289, n_20290, n_20291, n_20296,
       n_20297;
  wire n_20298, n_20299, n_20300, n_20301, n_20302, n_20303, n_20304,
       n_20305;
  wire n_20306, n_20307, n_20308, n_20309, n_20310, n_20311, n_20312,
       n_20313;
  wire n_20314, n_20315, n_20316, n_20317, n_20318, n_20319, n_20320,
       n_20321;
  wire n_20322, n_20323, n_20324, n_20325, n_20330, n_20331, n_20332,
       n_20333;
  wire n_20334, n_20335, n_20336, n_20337, n_20338, n_20339, n_20340,
       n_20341;
  wire n_20346, n_20347, n_20348, n_20349, n_20350, n_20351, n_20352,
       n_20353;
  wire n_20354, n_20355, n_20356, n_20357, n_20362, n_20363, n_20364,
       n_20365;
  wire n_20366, n_20367, n_20368, n_20369, n_20370, n_20371, n_20372,
       n_20373;
  wire n_20378, n_20379, n_20380, n_20381, n_20382, n_20383, n_20384,
       n_20385;
  wire n_20386, n_20387, n_20388, n_20389, n_20394, n_20395, n_20396,
       n_20397;
  wire n_20398, n_20399, n_20400, n_20401, n_20402, n_20403, n_20404,
       n_20405;
  wire n_20406, n_20411, n_20412, n_20413, n_20414, n_20415, n_20416,
       n_20417;
  wire n_20418, n_20419, n_20420, n_20421, n_20422, n_20423, n_20428,
       n_20429;
  wire n_20430, n_20431, n_20432, n_20433, n_20434, n_20435, n_20436,
       n_20437;
  wire n_20438, n_20439, n_20440, n_20441, n_20442, n_20443, n_20444,
       n_20445;
  wire n_20446, n_20447, n_20448, n_20449, n_20450, n_20451, n_20452,
       n_20457;
  wire n_20458, n_20459, n_20460, n_20461, n_20462, n_20463, n_20464,
       n_20465;
  wire n_20470, n_20471, n_20472, n_20473, n_20474, n_20475, n_20476,
       n_20477;
  wire n_20482, n_20483, n_20484, n_20485, n_20486, n_20487, n_20488,
       n_20489;
  wire n_20490, n_20491, n_20492, n_20493, n_20494, n_20499, n_20500,
       n_20501;
  wire n_20502, n_20503, n_20504, n_20505, n_20506, n_20507, n_20508,
       n_20509;
  wire n_20510, n_20515, n_20516, n_20517, n_20518, n_20519, n_20520,
       n_20521;
  wire n_20522, n_20523, n_20524, n_20525, n_20526, n_20531, n_20532,
       n_20533;
  wire n_20534, n_20535, n_20536, n_20537, n_20538, n_20539, n_20540,
       n_20541;
  wire n_20542, n_20547, n_20548, n_20549, n_20550, n_20551, n_20552,
       n_20553;
  wire n_20554, n_20555, n_20556, n_20557, n_20558, n_20563, n_20564,
       n_20565;
  wire n_20566, n_20567, n_20568, n_20569, n_20570, n_20571, n_20572,
       n_20573;
  wire n_20574, n_20575, n_20576, n_20577, n_20578, n_20579, n_20580,
       n_20581;
  wire n_20582, n_20583, n_20584, n_20585, n_20586, n_20587, n_20588,
       n_20589;
  wire n_20590, n_20591, n_20592, n_20593, n_20594, n_20595, n_20596,
       n_20597;
  wire n_20602, n_20603, n_20604, n_20605, n_20606, n_20607, n_20608,
       n_20609;
  wire n_20610, n_20611, n_20612, n_20613, n_20614, n_20615, n_20616,
       n_20617;
  wire n_20618, n_20619, n_20624, n_20625, n_20626, n_20627, n_20628,
       n_20629;
  wire n_20630, n_20631, n_20632, n_20633, n_20634, n_20635, n_20636,
       n_20641;
  wire n_20642, n_20643, n_20644, n_20645, n_20646, n_20647, n_20648,
       n_20649;
  wire n_20650, n_20651, n_20652, n_20657, n_20658, n_20659, n_20660,
       n_20661;
  wire n_20662, n_20663, n_20664, n_20665, n_20666, n_20667, n_20668,
       n_20673;
  wire n_20674, n_20675, n_20676, n_20677, n_20678, n_20679, n_20680,
       n_20681;
  wire n_20682, n_20683, n_20684, n_20689, n_20690, n_20691, n_20692,
       n_20693;
  wire n_20694, n_20695, n_20696, n_20697, n_20698, n_20699, n_20700,
       n_20701;
  wire n_20706, n_20707, n_20708, n_20709, n_20710, n_20711, n_20712,
       n_20713;
  wire n_20714, n_20715, n_20716, n_20717, n_20722, n_20723, n_20724,
       n_20725;
  wire n_20726, n_20727, n_20728, n_20729, n_20730, n_20731, n_20732,
       n_20733;
  wire n_20734, n_20735, n_20736, n_20737, n_20738, n_20739, n_20740,
       n_20741;
  wire n_20742, n_20743, n_20744, n_20745, n_20750, n_20751, n_20752,
       n_20753;
  wire n_20754, n_20755, n_20756, n_20757, n_20758, n_20759, n_20760,
       n_20761;
  wire n_20762, n_20763, n_20764, n_20765, n_20766, n_20767, n_20768,
       n_20769;
  wire n_20770, n_20771, n_20772, n_20773, n_20774, n_20775, n_20776,
       n_20777;
  wire n_20782, n_20783, n_20784, n_20785, n_20786, n_20787, n_20788,
       n_20789;
  wire n_20790, n_20791, n_20792, n_20793, n_20798, n_20799, n_20800,
       n_20801;
  wire n_20802, n_20803, n_20804, n_20805, n_20806, n_20807, n_20808,
       n_20809;
  wire n_20814, n_20815, n_20816, n_20817, n_20818, n_20819, n_20820,
       n_20821;
  wire n_20822, n_20823, n_20824, n_20825, n_20830, n_20831, n_20832,
       n_20833;
  wire n_20834, n_20835, n_20836, n_20837, n_20838, n_20839, n_20840,
       n_20841;
  wire n_20842, n_20847, n_20848, n_20849, n_20850, n_20851, n_20852,
       n_20853;
  wire n_20854, n_20855, n_20856, n_20857, n_20858, n_20859, n_20864,
       n_20865;
  wire n_20866, n_20867, n_20868, n_20869, n_20870, n_20871, n_20872,
       n_20873;
  wire n_20874, n_20875, n_20876, n_20877, n_20878, n_20879, n_20880,
       n_20881;
  wire n_20882, n_20883, n_20884, n_20885, n_20886, n_20887, n_20888,
       n_20893;
  wire n_20894, n_20895, n_20896, n_20897, n_20898, n_20899, n_20900,
       n_20901;
  wire n_20902, n_20903, n_20904, n_20905, n_20906, n_20907, n_20908,
       n_20909;
  wire n_20910, n_20911, n_20912, n_20913, n_20918, n_20919, n_20920,
       n_20921;
  wire n_20922, n_20923, n_20924, n_20925, n_20926, n_20927, n_20928,
       n_20929;
  wire n_20934, n_20935, n_20936, n_20937, n_20938, n_20939, n_20940,
       n_20941;
  wire n_20942, n_20943, n_20944, n_20945, n_20950, n_20951, n_20952,
       n_20953;
  wire n_20954, n_20955, n_20956, n_20957, n_20958, n_20959, n_20960,
       n_20961;
  wire n_20966, n_20967, n_20968, n_20969, n_20970, n_20971, n_20972,
       n_20973;
  wire n_20974, n_20975, n_20976, n_20977, n_20982, n_20983, n_20984,
       n_20985;
  wire n_20986, n_20987, n_20988, n_20989, n_20990, n_20991, n_20992,
       n_20993;
  wire n_20994, n_20995, n_20996, n_20997, n_20998, n_20999, n_21000,
       n_21001;
  wire n_21002, n_21003, n_21004, n_21005, n_21006, n_21007, n_21008,
       n_21009;
  wire n_21010, n_21011, n_21012, n_21013, n_21014, n_21015, n_21016,
       n_21021;
  wire n_21022, n_21023, n_21024, n_21025, n_21026, n_21027, n_21028,
       n_21029;
  wire n_21030, n_21031, n_21032, n_21033, n_21034, n_21035, n_21036,
       n_21037;
  wire n_21038, n_21039, n_21040, n_21041, n_21042, n_21043, n_21044,
       n_21049;
  wire n_21050, n_21051, n_21052, n_21053, n_21054, n_21055, n_21056,
       n_21057;
  wire n_21062, n_21063, n_21064, n_21065, n_21066, n_21067, n_21068,
       n_21069;
  wire n_21070, n_21071, n_21072, n_21073, n_21074, n_21079, n_21080,
       n_21081;
  wire n_21082, n_21083, n_21084, n_21085, n_21086, n_21087, n_21088,
       n_21089;
  wire n_21090, n_21095, n_21096, n_21097, n_21098, n_21099, n_21100,
       n_21101;
  wire n_21102, n_21103, n_21104, n_21105, n_21106, n_21107, n_21112,
       n_21113;
  wire n_21114, n_21115, n_21116, n_21117, n_21118, n_21119, n_21120,
       n_21121;
  wire n_21122, n_21123, n_21128, n_21129, n_21130, n_21131, n_21132,
       n_21133;
  wire n_21134, n_21135, n_21136, n_21137, n_21138, n_21139, n_21140,
       n_21141;
  wire n_21142, n_21143, n_21144, n_21145, n_21146, n_21147, n_21148,
       n_21149;
  wire n_21150, n_21151, n_21156, n_21157, n_21158, n_21159, n_21160,
       n_21161;
  wire n_21162, n_21163, n_21164, n_21165, n_21166, n_21167, n_21168,
       n_21169;
  wire n_21170, n_21171, n_21172, n_21173, n_21174, n_21175, n_21176,
       n_21177;
  wire n_21178, n_21179, n_21180, n_21181, n_21182, n_21183, n_21188,
       n_21189;
  wire n_21190, n_21191, n_21192, n_21193, n_21194, n_21195, n_21196,
       n_21197;
  wire n_21198, n_21199, n_21204, n_21205, n_21206, n_21207, n_21208,
       n_21209;
  wire n_21210, n_21211, n_21212, n_21213, n_21214, n_21215, n_21220,
       n_21221;
  wire n_21222, n_21223, n_21224, n_21225, n_21226, n_21227, n_21228,
       n_21229;
  wire n_21230, n_21231, n_21232, n_21237, n_21238, n_21239, n_21240,
       n_21241;
  wire n_21242, n_21243, n_21244, n_21245, n_21246, n_21247, n_21248,
       n_21249;
  wire n_21254, n_21255, n_21256, n_21257, n_21258, n_21259, n_21260,
       n_21261;
  wire n_21262, n_21263, n_21264, n_21265, n_21266, n_21267, n_21268,
       n_21269;
  wire n_21270, n_21271, n_21276, n_21277, n_21278, n_21279, n_21280,
       n_21281;
  wire n_21282, n_21283, n_21284, n_21285, n_21286, n_21287, n_21288,
       n_21289;
  wire n_21290, n_21295, n_21296, n_21297, n_21298, n_21299, n_21300,
       n_21301;
  wire n_21302, n_21307, n_21308, n_21309, n_21310, n_21311, n_21312,
       n_21313;
  wire n_21314, n_21315, n_21316, n_21317, n_21318, n_21319, n_21324,
       n_21325;
  wire n_21326, n_21327, n_21328, n_21329, n_21330, n_21331, n_21332,
       n_21333;
  wire n_21334, n_21335, n_21340, n_21341, n_21342, n_21343, n_21344,
       n_21345;
  wire n_21346, n_21347, n_21348, n_21349, n_21350, n_21351, n_21356,
       n_21357;
  wire n_21358, n_21359, n_21360, n_21361, n_21362, n_21363, n_21364,
       n_21365;
  wire n_21366, n_21367, n_21368, n_21369, n_21370, n_21371, n_21372,
       n_21373;
  wire n_21374, n_21375, n_21376, n_21377, n_21378, n_21379, n_21380,
       n_21381;
  wire n_21382, n_21383, n_21384, n_21385, n_21386, n_21387, n_21388,
       n_21389;
  wire n_21390, n_21395, n_21396, n_21397, n_21398, n_21399, n_21400,
       n_21401;
  wire n_21402, n_21403, n_21404, n_21405, n_21406, n_21407, n_21408,
       n_21409;
  wire n_21410, n_21411, n_21412, n_21417, n_21418, n_21419, n_21420,
       n_21421;
  wire n_21422, n_21423, n_21424, n_21425, n_21426, n_21427, n_21428,
       n_21429;
  wire n_21434, n_21435, n_21436, n_21437, n_21438, n_21439, n_21440,
       n_21441;
  wire n_21442, n_21443, n_21444, n_21445, n_21450, n_21451, n_21452,
       n_21453;
  wire n_21454, n_21455, n_21456, n_21457, n_21458, n_21459, n_21460,
       n_21461;
  wire n_21462, n_21467, n_21468, n_21469, n_21470, n_21471, n_21472,
       n_21473;
  wire n_21474, n_21475, n_21476, n_21477, n_21478, n_21483, n_21484,
       n_21485;
  wire n_21486, n_21487, n_21488, n_21489, n_21490, n_21491, n_21492,
       n_21493;
  wire n_21494, n_21495, n_21496, n_21497, n_21498, n_21499, n_21500,
       n_21501;
  wire n_21502, n_21503, n_21504, n_21505, n_21506, n_21511, n_21512,
       n_21513;
  wire n_21514, n_21515, n_21516, n_21517, n_21518, n_21519, n_21520,
       n_21521;
  wire n_21522, n_21523, n_21524, n_21525, n_21526, n_21527, n_21528,
       n_21529;
  wire n_21530, n_21531, n_21532, n_21533, n_21534, n_21535, n_21536,
       n_21537;
  wire n_21538, n_21543, n_21544, n_21545, n_21546, n_21547, n_21548,
       n_21549;
  wire n_21550, n_21551, n_21552, n_21553, n_21554, n_21559, n_21560,
       n_21561;
  wire n_21562, n_21563, n_21564, n_21565, n_21566, n_21567, n_21568,
       n_21569;
  wire n_21570, n_21571, n_21576, n_21577, n_21578, n_21579, n_21580,
       n_21581;
  wire n_21582, n_21583, n_21584, n_21585, n_21586, n_21587, n_21588,
       n_21593;
  wire n_21594, n_21595, n_21596, n_21597, n_21598, n_21599, n_21600,
       n_21601;
  wire n_21602, n_21603, n_21604, n_21605, n_21606, n_21607, n_21608,
       n_21609;
  wire n_21610, n_21611, n_21612, n_21613, n_21614, n_21615, n_21616,
       n_21617;
  wire n_21622, n_21623, n_21624, n_21625, n_21626, n_21627, n_21628,
       n_21629;
  wire n_21630, n_21631, n_21632, n_21633, n_21634, n_21635, n_21636,
       n_21637;
  wire n_21638, n_21639, n_21640, n_21641, n_21642, n_21647, n_21648,
       n_21649;
  wire n_21650, n_21651, n_21652, n_21653, n_21654, n_21655, n_21656,
       n_21657;
  wire n_21658, n_21663, n_21664, n_21665, n_21666, n_21667, n_21668,
       n_21669;
  wire n_21670, n_21671, n_21672, n_21673, n_21674, n_21679, n_21680,
       n_21681;
  wire n_21682, n_21683, n_21684, n_21685, n_21686, n_21687, n_21688,
       n_21689;
  wire n_21690, n_21691, n_21692, n_21693, n_21694, n_21695, n_21696,
       n_21697;
  wire n_21698, n_21699, n_21700, n_21701, n_21702, n_21703, n_21704,
       n_21705;
  wire n_21706, n_21707, n_21708, n_21709, n_21710, n_21711, n_21712,
       n_21713;
  wire n_21718, n_21719, n_21720, n_21721, n_21722, n_21723, n_21724,
       n_21725;
  wire n_21726, n_21731, n_21732, n_21733, n_21734, n_21735, n_21736,
       n_21737;
  wire n_21738, n_21739, n_21740, n_21741, n_21742, n_21743, n_21744,
       n_21745;
  wire n_21746, n_21747, n_21748, n_21749, n_21750, n_21751, n_21752,
       n_21753;
  wire n_21754, n_21759, n_21760, n_21761, n_21762, n_21763, n_21764,
       n_21765;
  wire n_21766, n_21767, n_21768, n_21769, n_21770, n_21771, n_21776,
       n_21777;
  wire n_21778, n_21779, n_21780, n_21781, n_21782, n_21783, n_21784,
       n_21785;
  wire n_21786, n_21787, n_21792, n_21793, n_21794, n_21795, n_21796,
       n_21797;
  wire n_21798, n_21799, n_21800, n_21801, n_21802, n_21803, n_21804,
       n_21805;
  wire n_21806, n_21807, n_21808, n_21809, n_21810, n_21811, n_21812,
       n_21813;
  wire n_21814, n_21815, n_21820, n_21821, n_21822, n_21823, n_21824,
       n_21825;
  wire n_21826, n_21827, n_21828, n_21829, n_21830, n_21831, n_21832,
       n_21833;
  wire n_21834, n_21835, n_21836, n_21837, n_21838, n_21839, n_21840,
       n_21841;
  wire n_21842, n_21843, n_21844, n_21845, n_21846, n_21847, n_21852,
       n_21853;
  wire n_21854, n_21855, n_21856, n_21857, n_21858, n_21859, n_21860,
       n_21861;
  wire n_21862, n_21863, n_21864, n_21865, n_21870, n_21871, n_21872,
       n_21873;
  wire n_21874, n_21875, n_21876, n_21877, n_21878, n_21879, n_21880,
       n_21881;
  wire n_21882, n_21887, n_21888, n_21889, n_21890, n_21891, n_21892,
       n_21893;
  wire n_21894, n_21895, n_21896, n_21897, n_21898, n_21899, n_21900,
       n_21901;
  wire n_21902, n_21903, n_21904, n_21909, n_21910, n_21911, n_21912,
       n_21913;
  wire n_21914, n_21915, n_21916, n_21917, n_21918, n_21919, n_21920,
       n_21921;
  wire n_21922, n_21923, n_21928, n_21929, n_21930, n_21931, n_21932,
       n_21933;
  wire n_21934, n_21935, n_21940, n_21941, n_21942, n_21943, n_21944,
       n_21945;
  wire n_21946, n_21947, n_21948, n_21949, n_21950, n_21951, n_21952,
       n_21957;
  wire n_21958, n_21959, n_21960, n_21961, n_21962, n_21963, n_21964,
       n_21965;
  wire n_21966, n_21967, n_21968, n_21969, n_21970, n_21971, n_21972,
       n_21973;
  wire n_21974, n_21975, n_21976, n_21977, n_21978, n_21979, n_21980,
       n_21981;
  wire n_21982, n_21983, n_21984, n_21985, n_21986, n_21987, n_21988,
       n_21989;
  wire n_21990, n_21991, n_21996, n_21997, n_21998, n_21999, n_22000,
       n_22001;
  wire n_22002, n_22003, n_22004, n_22005, n_22006, n_22007, n_22008,
       n_22009;
  wire n_22010, n_22011, n_22012, n_22013, n_22014, n_22015, n_22016,
       n_22017;
  wire n_22022, n_22023, n_22024, n_22025, n_22026, n_22027, n_22028,
       n_22029;
  wire n_22034, n_22035, n_22036, n_22037, n_22038, n_22039, n_22040,
       n_22041;
  wire n_22042, n_22043, n_22044, n_22045, n_22046, n_22051, n_22052,
       n_22053;
  wire n_22054, n_22055, n_22056, n_22057, n_22058, n_22059, n_22060,
       n_22061;
  wire n_22062, n_22063, n_22064, n_22065, n_22066, n_22067, n_22068,
       n_22069;
  wire n_22070, n_22071, n_22072, n_22073, n_22074, n_22079, n_22080,
       n_22081;
  wire n_22082, n_22083, n_22084, n_22085, n_22086, n_22087, n_22088,
       n_22089;
  wire n_22090, n_22091, n_22092, n_22093, n_22094, n_22095, n_22096,
       n_22097;
  wire n_22098, n_22099, n_22100, n_22101, n_22102, n_22103, n_22104,
       n_22105;
  wire n_22106, n_22111, n_22112, n_22113, n_22114, n_22115, n_22116,
       n_22117;
  wire n_22118, n_22119, n_22120, n_22121, n_22122, n_22127, n_22128,
       n_22129;
  wire n_22130, n_22131, n_22132, n_22133, n_22134, n_22135, n_22136,
       n_22137;
  wire n_22138, n_22139, n_22140, n_22141, n_22142, n_22143, n_22144,
       n_22145;
  wire n_22146, n_22147, n_22148, n_22149, n_22150, n_22151, n_22156,
       n_22157;
  wire n_22158, n_22159, n_22160, n_22161, n_22162, n_22163, n_22164,
       n_22169;
  wire n_22170, n_22171, n_22172, n_22173, n_22174, n_22175, n_22176,
       n_22181;
  wire n_22182, n_22183, n_22184, n_22185, n_22186, n_22187, n_22188,
       n_22189;
  wire n_22190, n_22191, n_22192, n_22193, n_22194, n_22195, n_22196,
       n_22197;
  wire n_22198, n_22199, n_22200, n_22201, n_22202, n_22203, n_22204,
       n_22205;
  wire n_22206, n_22207, n_22208, n_22209, n_22210, n_22211, n_22212,
       n_22213;
  wire n_22214, n_22215, n_22216, n_22221, n_22222, n_22223, n_22224,
       n_22225;
  wire n_22226, n_22227, n_22228, n_22229, n_22234, n_22235, n_22236,
       n_22237;
  wire n_22238, n_22239, n_22240, n_22241, n_22242, n_22243, n_22244,
       n_22245;
  wire n_22246, n_22247, n_22248, n_22249, n_22250, n_22251, n_22252,
       n_22253;
  wire n_22254, n_22255, n_22260, n_22261, n_22262, n_22263, n_22264,
       n_22265;
  wire n_22266, n_22267, n_22268, n_22269, n_22270, n_22271, n_22272,
       n_22273;
  wire n_22274, n_22275, n_22276, n_22277, n_22278, n_22279, n_22280,
       n_22281;
  wire n_22282, n_22287, n_22288, n_22289, n_22290, n_22291, n_22292,
       n_22293;
  wire n_22294, n_22295, n_22296, n_22297, n_22298, n_22299, n_22300,
       n_22301;
  wire n_22302, n_22303, n_22304, n_22305, n_22306, n_22307, n_22308,
       n_22309;
  wire n_22310, n_22311, n_22312, n_22313, n_22314, n_22319, n_22320,
       n_22321;
  wire n_22322, n_22323, n_22324, n_22325, n_22326, n_22327, n_22328,
       n_22329;
  wire n_22330, n_22331, n_22332, n_22333, n_22334, n_22335, n_22336,
       n_22337;
  wire n_22338, n_22339, n_22340, n_22341, n_22342, n_22343, n_22344,
       n_22349;
  wire n_22350, n_22351, n_22352, n_22353, n_22354, n_22355, n_22356,
       n_22357;
  wire n_22358, n_22359, n_22360, n_22361, n_22362, n_22363, n_22364,
       n_22369;
  wire n_22370, n_22371, n_22372, n_22373, n_22374, n_22375, n_22376,
       n_22377;
  wire n_22378, n_22379, n_22380, n_22381, n_22382, n_22383, n_22384,
       n_22385;
  wire n_22386, n_22387, n_22388, n_22389, n_22390, n_22391, n_22392,
       n_22393;
  wire n_22398, n_22399, n_22400, n_22401, n_22402, n_22403, n_22404,
       n_22409;
  wire n_22410, n_22411, n_22412, n_22413, n_22414, n_22415, n_22416,
       n_22417;
  wire n_22418, n_22419, n_22420, n_22421, n_22422, n_22423, n_22424,
       n_22425;
  wire n_22426, n_22427, n_22428, n_22429, n_22430, n_22431, n_22432,
       n_22433;
  wire n_22434, n_22435, n_22436, n_22437, n_22438, n_22439, n_22472,
       n_22473;
  wire n_22474, n_22475, n_22476, n_22477, n_22478, n_22479, n_22480,
       n_22481;
  wire n_22482, n_22483, n_22484, n_22485, n_22486, n_22487, n_22488,
       n_22489;
  wire n_22490, n_22491, n_22492, n_22493, n_22494, n_22495, n_22496,
       n_22497;
  wire n_22498, n_22499, n_22500, n_22501, n_22502, n_22503, n_22504,
       n_22505;
  wire n_22506, n_22507, n_22508, n_22509, n_22510, n_22511, n_22512,
       n_22513;
  wire n_22514, n_22515, n_22516, n_22517, n_22518, n_22519, n_22520,
       n_22521;
  wire n_22522, n_22523, n_22524, n_22525, n_22526, n_22527, n_22528,
       n_22529;
  wire n_22530, n_22531, n_22532, n_22533, n_22534, n_22535, n_22536,
       n_22537;
  wire n_22538, n_22539, n_22540, n_22541, n_22542, n_22543, n_22544,
       n_22545;
  wire n_22546, n_22547, n_22548, n_22549, n_22550, n_22551, n_22552,
       n_22553;
  wire n_22554, n_22555, n_22556, n_22557, n_22558, n_22559, n_22560,
       n_22561;
  wire n_22562, n_22563, n_22564, n_22565, n_22566, n_22567, n_22568,
       n_22569;
  wire n_22570, n_22571, n_22572, n_22573, n_22574, n_22575, n_22576,
       n_22577;
  wire n_22578, n_22579, n_22580, n_22581, n_22582, n_22583, n_22584,
       n_22585;
  wire n_22586, n_22587, n_22588, n_22589, n_22590, n_22591, n_22592,
       n_22593;
  wire n_22594, n_22595, n_22596, n_22597, n_22598, n_22599, n_22600,
       n_22601;
  wire n_22602, n_22603, n_22604, n_22605, n_22606, n_22607, n_22608,
       n_22609;
  wire n_22610, n_22611, n_22612, n_22613, n_22614, n_22615, n_22616,
       n_22617;
  wire n_22618, n_22619, n_22620, n_22621, n_22622, n_22623, n_22624,
       n_22625;
  wire n_22626, n_22627, n_22628, n_22629, n_22630, n_22631, n_22632,
       n_22633;
  wire n_22634, n_22635, n_22636, n_22637, n_22638, n_22639, n_22640,
       n_22641;
  wire n_22642, n_22643, n_22644, n_22645, n_22646, n_22647, n_22648,
       n_22650;
  wire n_22651, n_22652, n_22653, n_22654, n_22655, n_22656, n_22657,
       n_22658;
  wire n_22659, n_22660, n_22661, n_22662, n_22663, n_22664, n_22665,
       n_22666;
  wire n_22667, n_22668, n_22669, n_22670, n_22671, n_22672, n_22673,
       n_22674;
  wire n_22675, n_22676, n_22677, n_22678, n_22679, n_22680, n_22681,
       n_22682;
  wire n_22683, n_22684, n_22685, n_22686, n_22687, n_22688, n_22689,
       n_22690;
  wire n_22691, n_22692, n_22693, n_22694, n_22695, n_22696, n_22697,
       n_22698;
  wire n_22699, n_22700, n_22701, n_22702, n_22703, n_22704, n_22705,
       n_22706;
  wire n_22707, n_22708, n_22709, n_22710, n_22711, n_22712, n_22713,
       n_22714;
  wire n_22715, n_22716, n_22717, n_22718, n_22719, n_22720, n_22721,
       n_22722;
  wire n_22723, n_22724, n_22725, n_22726, n_22727, n_22728, n_22729,
       n_22730;
  wire n_22731, n_22732, n_22733, n_22734, n_22735, n_22736, n_22737,
       n_22738;
  wire n_22739, n_22740, n_22741, n_22742, n_22743, n_22744, n_22745,
       n_22746;
  wire n_22747, n_22748, n_22749, n_22750, n_22751, n_22752, n_22753,
       n_22754;
  wire n_22755, n_22756, n_22757, n_22758, n_22759, n_22760, n_22761,
       n_22762;
  wire n_22763, n_22764, n_22765, n_22766, n_22767, n_22768, n_22769,
       n_22770;
  wire n_22771, n_22772, n_22773, n_22774, n_22775, n_22776, n_22777,
       n_22778;
  wire n_22779, n_22780, n_22781, n_22782, n_22783, n_22784, n_22785,
       n_22786;
  wire n_22787, n_22788, n_22789, n_22790, n_22791, n_22792, n_22793,
       n_22794;
  wire n_22795, n_22796, n_22797, n_22798, n_22799, n_22800, n_22801,
       n_22802;
  wire n_22803, n_22804, n_22805, n_22806, n_22807, n_22808, n_22809,
       n_22810;
  wire n_22811, n_22812, n_22813, n_22814, n_22815, n_22816, n_22817,
       n_22818;
  wire n_22819, n_22820, n_22821, n_22822, n_22823, n_22824, n_22825,
       n_22826;
  wire n_22827, n_22828, n_22829, n_22830, n_22831, n_22832, n_22833,
       n_22834;
  wire n_22835, n_22836, n_22837, n_22838, n_22839, n_22840, n_22841,
       n_22842;
  wire n_22843, n_22844, n_22845, n_22846, n_22847, n_22848, n_22849,
       n_22850;
  wire n_22851, n_22852, n_22853, n_22854, n_22855, n_22856, n_22857,
       n_22858;
  wire n_22859, n_22860, n_22861, n_22862, n_22863, n_22864, n_22865,
       n_22866;
  wire n_22867, n_22868, n_22869, n_22870, n_22871, n_22872, n_22873,
       n_22874;
  wire n_22875, n_22876, n_22877, n_22878, n_22879, n_22880, n_22881,
       n_22882;
  wire n_22883, n_22884, n_22885, n_22886, n_22887, n_22888, n_22889,
       n_22890;
  wire n_22891, n_22892, n_22893, n_22894, n_22895, n_22896, n_22897,
       n_22898;
  wire n_22899, n_22900, n_22901, n_22902, n_22903, n_22904, n_22905,
       n_22906;
  wire n_22907, n_22908, n_22909, n_22910, n_22911, n_22912, n_22913,
       n_22914;
  wire n_22915, n_22916, n_22917, n_22918, n_22919, n_22920, n_22921,
       n_22922;
  wire n_22923, n_22924, n_22925, n_22926, n_22927, n_22928, n_22929,
       n_22930;
  wire n_22931, n_22932, n_22933, n_22934, n_22935, n_22936, n_22937,
       n_22938;
  wire n_22939, n_22940, n_22941, n_22942, n_22943, n_22944, n_22945,
       n_22946;
  wire n_22947, n_22948, n_22949, n_22950, n_22951, n_22952, n_22953,
       n_22954;
  wire n_22955, n_22956, n_22957, n_22958, n_22959, n_22960, n_22961,
       n_22962;
  wire n_22963, n_22964, n_22965, n_22966, n_22967, n_22968, n_22969,
       n_22970;
  wire n_22971, n_22972, n_22973, n_22974, n_22975, n_22976, n_22977,
       n_22978;
  wire n_22979, n_22980, n_22981, n_22982, n_22983, n_22984, n_22985,
       n_22986;
  wire n_22987, n_22988, n_22989, n_22990, n_22991, n_22992, n_22993,
       n_22994;
  wire n_22995, n_22996, n_22997, n_22998, n_22999, n_23000, n_23001,
       n_23002;
  wire n_23003, n_23004, n_23005, n_23006, n_23007, n_23008, n_23009,
       n_23010;
  wire n_23011, n_23012, n_23013, n_23014, n_23015, n_23016, n_23017,
       n_23018;
  wire n_23019, n_23020, n_23021, n_23022, n_23023, n_23024, n_23025,
       n_23026;
  wire n_23027, n_23028, n_23029, n_23030, n_23031, n_23032, n_23033,
       n_23034;
  wire n_23035, n_23036, n_23037, n_23038, n_23039, n_23040, n_23041,
       n_23042;
  wire n_23043, n_23044, n_23045, n_23046, n_23047, n_23048, n_23049,
       n_23050;
  wire n_23051, n_23052, n_23053, n_23054, n_23055, n_23056, n_23057,
       n_23058;
  wire n_23059, n_23060, n_23061, n_23062, n_23063, n_23064, n_23065,
       n_23066;
  wire n_23067, n_23068, n_23069, n_23070, n_23071, n_23072, n_23073,
       n_23074;
  wire n_23075, n_23076, n_23077, n_23078, n_23080, n_23081, n_23082,
       n_23083;
  wire n_23084, n_23085, n_23086, n_23087, n_23088, n_23089, n_23090,
       n_23091;
  wire n_23092, n_23093, n_23094, n_23095, n_23096, n_23097, n_23098,
       n_23099;
  wire n_23100, n_23101, n_23102, n_23103, n_23104, n_23105, n_23106,
       n_23107;
  wire n_23108, n_23109, n_23110, n_23111, n_23112, n_23113, n_23114,
       n_23115;
  wire n_23116, n_23117, n_23118, n_23119, n_23120, n_23121, n_23122,
       n_23123;
  wire n_23124, n_23125, n_23126, n_23127, n_23128, n_23129, n_23130,
       n_23131;
  wire n_23132, n_23133, n_23134, n_23135, n_23136, n_23137, n_23138,
       n_23139;
  wire n_23140, n_23141, n_23142, n_23143, n_23144, n_23145, n_23146,
       n_23147;
  wire n_23148, n_23149, n_23150, n_23151, n_23152, n_23153, n_23154,
       n_23155;
  wire n_23156, n_23157, n_23158, n_23159, n_23160, n_23161, n_23162,
       n_23163;
  wire n_23164, n_23165, n_23166, n_23167, n_23168, n_23169, n_23170,
       n_23171;
  wire n_23172, n_23173, n_23174, n_23175, n_23176, n_23177, n_23178,
       n_23179;
  wire n_23180, n_23181, n_23182, n_23183, n_23184, n_23185, n_23186,
       n_23187;
  wire n_23188, n_23189, n_23190, n_23191, n_23192, n_23193, n_23194,
       n_23195;
  wire n_23196, n_23197, n_23198, n_23199, n_23200, n_23201, n_23202,
       n_23203;
  wire n_23204, n_23205, n_23206, n_23207, n_23208, n_23209, n_23210,
       n_23211;
  wire n_23212, n_23213, n_23214, n_23215, n_23216, n_23217, n_23218,
       n_23219;
  wire n_23220, n_23221, n_23222, n_23223, n_23224, n_23225, n_23226,
       n_23227;
  wire n_23228, n_23229, n_23230, n_23231, n_23232, n_23233, n_23234,
       n_23235;
  wire n_23236, n_23237, n_23238, n_23239, n_23240, n_23241, n_23242,
       n_23243;
  wire n_23244, n_23245, n_23246, n_23247, n_23248, n_23249, n_23250,
       n_23251;
  wire n_23252, n_23253, n_23254, n_23255, n_23256, n_23257, n_23258,
       n_23259;
  wire n_23260, n_23261, n_23262, n_23263, n_23264, n_23265, n_23267,
       n_23268;
  wire n_23269, n_23270, n_23271, n_23272, n_23273, n_23274, n_23275,
       n_23276;
  wire n_23277, n_23278, n_23279, n_23280, n_23281, n_23282, n_23283,
       n_23284;
  wire n_23285, n_23286, n_23287, n_23288, n_23289, n_23290, n_23291,
       n_23292;
  wire n_23293, n_23294, n_23295, n_23296, n_23297, n_23298, n_23299,
       n_23300;
  wire n_23301, n_23302, n_23303, n_23304, n_23305, n_23306, n_23307,
       n_23308;
  wire n_23309, n_23310, n_23311, n_23312, n_23313, n_23314, n_23315,
       n_23316;
  wire n_23317, n_23318, n_23319, n_23320, n_23321, n_23322, n_23323,
       n_23324;
  wire n_23325, n_23326, n_23327, n_23328, n_23329, n_23330, n_23331,
       n_23332;
  wire n_23333, n_23334, n_23335, n_23336, n_23337, n_23338, n_23339,
       n_23340;
  wire n_23341, n_23342, n_23343, n_23344, n_23345, n_23346, n_23347,
       n_23348;
  wire n_23349, n_23350, n_23351, n_23352, n_23353, n_23354, n_23355,
       n_23356;
  wire n_23357, n_23358, n_23359, n_23360, n_23361, n_23362, n_23363,
       n_23364;
  wire n_23365, n_23366, n_23367, n_23368, n_23369, n_23370, n_23371,
       n_23372;
  wire n_23373, n_23374, n_23375, n_23376, n_23377, n_23378, n_23379,
       n_23380;
  wire n_23381, n_23382, n_23383, n_23384, n_23385, n_23386, n_23387,
       n_23388;
  wire n_23389, n_23390, n_23391, n_23392, n_23393, n_23394, n_23395,
       n_23396;
  wire n_23397, n_23398, n_23399, n_23400, n_23401, n_23402, n_23403,
       n_23404;
  wire n_23405, n_23406, n_23407, n_23408, n_23409, n_23410, n_23411,
       n_23412;
  wire n_23413, n_23414, n_23415, n_23416, n_23417, n_23418, n_23419,
       n_23420;
  wire n_23421, n_23422, n_23423, n_23424, n_23425, n_23426, n_23427,
       n_23428;
  wire n_23429, n_23430, n_23431, n_23432, n_23433, n_23434, n_23435,
       n_23436;
  wire n_23437, n_23438, n_23439, n_23440, n_23441, n_23442, n_23443,
       n_23444;
  wire n_23445, n_23446, n_23447, n_23448, n_23449, n_23450, n_23451,
       n_23452;
  wire n_23453, n_23454, n_23455, n_23456, n_23457, n_23458, n_23459,
       n_23460;
  wire n_23461, n_23462, n_23463, n_23464, n_23465, n_23466, n_23467,
       n_23468;
  wire n_23469, n_23470, n_23471, n_23472, n_23473, n_23474, n_23475,
       n_23476;
  wire n_23477, n_23478, n_23479, n_23480, n_23481, n_23482, n_23483,
       n_23484;
  wire n_23485, n_23486, n_23487, n_23488, n_23489, n_23490, n_23491,
       n_23492;
  wire n_23493, n_23494, n_23495, n_23496, n_23497, n_23498, n_23499,
       n_23500;
  wire n_23501, n_23502, n_23503, n_23504, n_23505, n_23506, n_23507,
       n_23508;
  wire n_23509, n_23510, n_23511, n_23512, n_23513, n_23514, n_23515,
       n_23516;
  wire n_23517, n_23518, n_23519, n_23520, n_23521, n_23522, n_23523,
       n_23524;
  wire n_23525, n_23526, n_23527, n_23528, n_23529, n_23530, n_23531,
       n_23532;
  wire n_23533, n_23534, n_23535, n_23536, n_23537, n_23538, n_23539,
       n_23540;
  wire n_23541, n_23542, n_23543, n_23544, n_23545, n_23546, n_23547,
       n_23548;
  wire n_23549, n_23550, n_23551, n_23552, n_23553, n_23554, n_23555,
       n_23556;
  wire n_23557, n_23558, n_23559, n_23560, n_23561, n_23562, n_23563,
       n_23564;
  wire n_23565, n_23566, n_23567, n_23568, n_23569, n_23570, n_23571,
       n_23572;
  wire n_23573, n_23574, n_23575, n_23576, n_23577, n_23578, n_23579,
       n_23580;
  wire n_23581, n_23582, n_23583, n_23584, n_23585, n_23586, n_23587,
       n_23588;
  wire n_23589, n_23590, n_23591, n_23592, n_23593, n_23594, n_23595,
       n_23596;
  wire n_23597, n_23598, n_23599, n_23600, n_23601, n_23602, n_23603,
       n_23604;
  wire n_23605, n_23606, n_23607, n_23608, n_23609, n_23610, n_23611,
       n_23612;
  wire n_23613, n_23614, n_23615, n_23616, n_23617, n_23618, n_23619,
       n_23620;
  wire n_23621, n_23622, n_23623, n_23624, n_23625, n_23626, n_23627,
       n_23628;
  wire n_23629, n_23630, n_23631, n_23632, n_23633, n_23634, n_23635,
       n_23636;
  wire n_23637, n_23638, n_23639, n_23640, n_23641, n_23642, n_23643,
       n_23644;
  wire n_23645, n_23646, n_23647, n_23648, n_23649, n_23650, n_23651,
       n_23652;
  wire n_23653, n_23654, n_23655, n_23656, n_23657, n_23658, n_23659,
       n_23660;
  wire n_23661, n_23662, n_23663, n_23664, n_23665, n_23666, n_23667,
       n_23668;
  wire n_23669, n_23670, n_23671, n_23672, n_23673, n_23674, n_23675,
       n_23676;
  wire n_23677, n_23678, n_23679, n_23680, n_23681, n_23682, n_23683,
       n_23684;
  wire n_23685, n_23686, n_23687, n_23688, n_23689, n_23690, n_23691,
       n_23692;
  wire n_23693, n_23694, n_23695, n_23696, n_23697, n_23698, n_23699,
       n_23700;
  wire n_23701, n_23702, n_23703, n_23704, n_23705, n_23706, n_23707,
       n_23708;
  wire n_23709, n_23710, n_23711, n_23712, n_23713, n_23714, n_23715,
       n_23716;
  wire n_23717, n_23718, n_23719, n_23720, n_23721, n_23722, n_23723,
       n_23724;
  wire n_23725, n_23726, n_23727, n_23728, n_23729, n_23730, n_23731,
       n_23732;
  wire n_23733, n_23734, n_23735, n_23736, n_23737, n_23738, n_23739,
       n_23740;
  wire n_23741, n_23742, n_23743, n_23744, n_23745, n_23746, n_23747,
       n_23748;
  wire n_23749, n_23750, n_23751, n_23752, n_23753, n_23754, n_23755,
       n_23756;
  wire n_23757, n_23758, n_23759, n_23760, n_23761, n_23762, n_23763,
       n_23764;
  wire n_23765, n_23766, n_23767, n_23768, n_23769, n_23770, n_23771,
       n_23772;
  wire n_23773, n_23774, n_23775, n_23776, n_23777, n_23778, n_23779,
       n_23780;
  wire n_23781, n_23782, n_23783, n_23784, n_23785, n_23786, n_23787,
       n_23788;
  wire n_23789, n_23790, n_23791, n_23792, n_23793, n_23794, n_23795,
       n_23796;
  wire n_23797, n_23798, n_23799, n_23800, n_23801, n_23802, n_23803,
       n_23804;
  wire n_23805, n_23806, n_23807, n_23808, n_23809, n_23810, n_23811,
       n_23812;
  wire n_23813, n_23814, n_23815, n_23816, n_23817, n_23818, n_23819,
       n_23820;
  wire n_23821, n_23822, n_23823, n_23824, n_23825, n_23826, n_23827,
       n_23828;
  wire n_23829, n_23830, n_23831, n_23832, n_23833, n_23834, n_23835,
       n_23836;
  wire n_23837, n_23839, n_23840, n_23841, n_23842, n_23843, n_23844,
       n_23845;
  wire n_23846, n_23847, n_23848, n_23849, n_23850, n_23851, n_23852,
       n_23853;
  wire n_23854, n_23855, n_23856, n_23857, n_23858, n_23859, n_23860,
       n_23863;
  wire n_23864, n_23865, n_23866, n_23867, n_23869, n_23870, n_23871,
       n_23872;
  wire n_23873, n_23874, n_23875, n_23876, n_23877, n_23878, n_23879,
       n_23880;
  wire n_23881, n_23882, n_23883, n_23884, n_23885, n_23886, n_23887,
       n_23888;
  wire n_23889, n_23890, n_23891, n_23892, n_23893, n_23894, n_23895,
       n_23896;
  wire n_23897, n_23898, n_23899, n_23900, n_23901, n_23902, n_23903,
       n_23904;
  wire n_23905, n_23906, n_23907, n_23908, n_23909, n_23910, n_23911,
       n_23912;
  wire n_23913, n_23914, n_23915, n_23916, n_23917, n_23918, n_23919,
       n_23920;
  wire n_23921, n_23922, n_23923, n_23924, n_23925, n_23926, n_23927,
       n_23928;
  wire n_23929, n_23930, n_23931, n_23932, n_23933, n_23934, n_23935,
       n_23936;
  wire n_23937, n_23938, n_23939, n_23940, n_23941, n_23942, n_23943,
       n_23944;
  wire n_23945, n_23946, n_23947, n_23948, n_23949, n_23950, n_23951,
       n_23952;
  wire n_23953, n_23954, n_23955, n_23956, n_23957, n_23958, n_23959,
       n_23960;
  wire n_23961, n_23962, n_23963, n_23964, n_23965, n_23966, n_23967,
       n_23968;
  wire n_23969, n_23970, n_23971, n_23972, n_23973, n_23974, n_23975,
       n_23976;
  wire n_23977, n_23978, n_23979, n_23980, n_23981, n_23982, n_23983,
       n_23984;
  wire n_23985, n_23986, n_23987, n_23988, n_23989, n_23990, n_23991,
       n_23992;
  wire n_23993, n_23994, n_23995, n_23996, n_23997, n_23998, n_23999,
       n_24000;
  wire n_24001, n_24002, n_24003, n_24004, n_24005, n_24006, n_24007,
       n_24008;
  wire n_24009, n_24010, n_24011, n_24012, n_24013, n_24014, n_24015,
       n_24016;
  wire n_24017, n_24018, n_24019, n_24020, n_24021, n_24022, n_24023,
       n_24024;
  wire n_24025, n_24026, n_24027, n_24028, n_24029, n_24030, n_24031,
       n_24032;
  wire n_24033, n_24034, n_24035, n_24036, n_24037, n_24038, n_24039,
       n_24040;
  wire n_24041, n_24042, n_24043, n_24044, n_24045, n_24046, n_24047,
       n_24048;
  wire n_24049, n_24050, n_24051, n_24052, n_24053, n_24054, n_24055,
       n_24056;
  wire n_24057, n_24058, n_24059, n_24060, n_24061, n_24062, n_24063,
       n_24064;
  wire n_24065, n_24066, n_24067, n_24068, n_24069, n_24070, n_24071,
       n_24072;
  wire n_24073, n_24074, n_24075, n_24076, n_24077, n_24078, n_24079,
       n_24080;
  wire n_24081, n_24082, n_24083, n_24084, n_24085, n_24086, n_24087,
       n_24088;
  wire n_24089, n_24090, n_24091, n_24092, n_24093, n_24094, n_24095,
       n_24096;
  wire n_24097, n_24098, n_24099, n_24100, n_24101, n_24102, n_24103,
       n_24104;
  wire n_24105, n_24106, n_24107, n_24108, n_24109, n_24110, n_24111,
       n_24112;
  wire n_24113, n_24114, n_24115, n_24116, n_24117, n_24118, n_24119,
       n_24120;
  wire n_24121, n_24122, n_24123, n_24124, n_24125, n_24126, n_24127,
       n_24129;
  wire n_24130, n_24131, n_24132, n_24133, n_24134, n_24135, n_24136,
       n_24137;
  wire n_24138, n_24139, n_24140, n_24141, n_24142, n_24143, n_24144,
       n_24145;
  wire n_24146, n_24147, n_24148, n_24149, n_24150, n_24151, n_24152,
       n_24153;
  wire n_24154, n_24155, n_24156, n_24157, n_24158, n_24159, n_24160,
       n_24161;
  wire n_24162, n_24163, n_24164, n_24165, n_24166, n_24167, n_24169,
       n_24170;
  wire n_24171, n_24172, n_24173, n_24174, n_24175, n_24176, n_24177,
       n_24178;
  wire n_24179, n_24180, n_24181, n_24182, n_24183, n_24184, n_24185,
       n_24186;
  wire n_24187, n_24188, n_24189, n_24190, n_24191, n_24192, n_24193,
       n_24194;
  wire n_24195, n_24196, n_24197, n_24198, n_24199, n_24200, n_24201,
       n_24202;
  wire n_24203, n_24204, n_24205, n_24206, n_24207, n_24208, n_24209,
       n_24210;
  wire n_24211, n_24212, n_24213, n_24214, n_24215, n_24216, n_24217,
       n_24218;
  wire n_24219, n_24220, n_24221, n_24222, n_24223, n_24224, n_24225,
       n_24226;
  wire n_24227, n_24228, n_24229, n_24230, n_24231, n_24232, n_24233,
       n_24234;
  wire n_24235, n_24236, n_24237, n_24238, n_24239, n_24240, n_24241,
       n_24242;
  wire n_24243, n_24244, n_24245, n_24246, n_24247, n_24248, n_24249,
       n_24250;
  wire n_24251, n_24252, n_24253, n_24254, n_24255, n_24256, n_24257,
       n_24258;
  wire n_24259, n_24260, n_24261, n_24262, n_24263, n_24264, n_24265,
       n_24266;
  wire n_24267, n_24268, n_24269, n_24270, n_24271, n_24272, n_24273,
       n_24274;
  wire n_24275, n_24276, n_24277, n_24278, n_24279, n_24281, n_24282,
       n_24283;
  wire n_24284, n_24285, n_24286, n_24287, n_24288, n_24289, n_24290,
       n_24291;
  wire n_24292, n_24293, n_24294, n_24295, n_24296, n_24297, n_24298,
       n_24299;
  wire n_24300, n_24301, n_24302, n_24303, n_24304, n_24305, n_24306,
       n_24307;
  wire n_24308, n_24309, n_24310, n_24311, n_24312, n_24313, n_24314,
       n_24315;
  wire n_24316, n_24317, n_24318, n_24319, n_24320, n_24321, n_24322,
       n_24323;
  wire n_24324, n_24325, n_24326, n_24327, n_24328, n_24329, n_24330,
       n_24331;
  wire n_24332, n_24333, n_24334, n_24335, n_24336, n_24337, n_24338,
       n_24339;
  wire n_24340, n_24341, n_24342, n_24343, n_24344, n_24345, n_24346,
       n_24347;
  wire n_24348, n_24349, n_24350, n_24351, n_24352, n_24353, n_24354,
       n_24355;
  wire n_24356, n_24357, n_24358, n_24359, n_24360, n_24361, n_24362,
       n_24363;
  wire n_24364, n_24365, n_24366, n_24367, n_24368, n_24369, n_24370,
       n_24371;
  wire n_24372, n_24373, n_24374, n_24375, n_24376, n_24377, n_24378,
       n_24379;
  wire n_24380, n_24381, n_24382, n_24383, n_24384, n_24385, n_24386,
       n_24387;
  wire n_24388, n_24389, n_24390, n_24391, n_24392, n_24393, n_24394,
       n_24395;
  wire n_24396, n_24397, n_24398, n_24399, n_24400, n_24401, n_24402,
       n_24403;
  wire n_24404, n_24405, n_24406, n_24407, n_24408, n_24409, n_24410,
       n_24411;
  wire n_24412, n_24413;
  not g1 (n_3, \a[5] );
  and g2 (n65, \a[4] , n_3);
  not g3 (n_4, \a[4] );
  and g4 (n66, n_4, \a[5] );
  not g5 (n_5, n65);
  not g6 (n_6, n66);
  and g7 (n67, n_5, n_6);
  not g8 (n_9, \a[3] );
  and g9 (n68, \a[2] , n_9);
  not g10 (n_10, \a[2] );
  and g11 (n69, n_10, \a[3] );
  not g12 (n_11, n68);
  not g13 (n_12, n69);
  and g14 (n70, n_11, n_12);
  not g15 (n_13, n70);
  and g16 (n71, n67, n_13);
  not g17 (n_15, \a[29] );
  and g18 (n72, n_15, \a[30] );
  not g19 (n_17, \a[30] );
  and g20 (n73, \a[29] , n_17);
  not g21 (n_18, n72);
  not g22 (n_19, n73);
  and g23 (n74, n_18, n_19);
  not g24 (n_21, n74);
  and g25 (n75, \a[31] , n_21);
  not g26 (n_24, \a[24] );
  not g27 (n_25, \a[25] );
  and g28 (n76, n_24, n_25);
  not g29 (n_27, \a[23] );
  and g30 (n77, n_27, \a[26] );
  and g31 (n78, n76, n77);
  and g32 (n79, \a[27] , \a[28] );
  and g33 (n80, n73, n79);
  and g34 (n81, n78, n80);
  not g35 (n_31, \a[27] );
  not g36 (n_32, \a[28] );
  and g37 (n82, n_31, n_32);
  and g38 (n83, n73, n82);
  and g39 (n84, \a[24] , \a[25] );
  and g40 (n85, n77, n84);
  and g41 (n86, n83, n85);
  not g42 (n_33, \a[26] );
  and g43 (n87, n_27, n_33);
  and g44 (n88, n76, n87);
  and g45 (n89, \a[29] , \a[30] );
  and g46 (n90, n79, n89);
  and g47 (n91, n88, n90);
  and g48 (n92, \a[23] , n_33);
  and g49 (n93, n_24, \a[25] );
  and g50 (n94, n92, n93);
  and g51 (n95, n83, n94);
  and g52 (n96, n84, n92);
  and g53 (n97, n_15, n_17);
  and g54 (n98, n82, n97);
  and g55 (n99, n96, n98);
  not g56 (n_34, n95);
  not g57 (n_35, n99);
  and g58 (n100, n_34, n_35);
  and g59 (n101, n87, n93);
  and g60 (n102, n90, n101);
  and g61 (n103, \a[27] , n_32);
  and g62 (n104, n89, n103);
  and g63 (n105, \a[23] , \a[26] );
  and g64 (n106, n93, n105);
  and g65 (n107, n104, n106);
  not g66 (n_36, n102);
  not g67 (n_37, n107);
  and g68 (n108, n_36, n_37);
  and g69 (n109, n_31, \a[28] );
  and g70 (n110, n72, n109);
  and g71 (n111, n96, n110);
  and g72 (n112, \a[24] , n_25);
  and g73 (n113, n92, n112);
  and g74 (n114, n72, n103);
  and g75 (n115, n113, n114);
  not g76 (n_38, n111);
  not g77 (n_39, n115);
  and g78 (n116, n_38, n_39);
  and g79 (n117, n82, n89);
  and g80 (n118, n94, n117);
  and g81 (n119, n83, n106);
  not g82 (n_40, n118);
  not g83 (n_41, n119);
  and g84 (n120, n_40, n_41);
  and g85 (n121, n88, n117);
  and g86 (n122, n87, n112);
  and g87 (n123, n110, n122);
  and g88 (n124, n77, n93);
  and g89 (n125, n83, n124);
  and g90 (n126, n105, n112);
  and g91 (n127, n83, n126);
  not g92 (n_42, n125);
  not g93 (n_43, n127);
  and g94 (n128, n_42, n_43);
  and g95 (n129, n97, n109);
  and g96 (n130, n113, n129);
  and g97 (n131, n76, n92);
  and g98 (n132, n129, n131);
  not g99 (n_44, n130);
  not g100 (n_45, n132);
  and g101 (n133, n_44, n_45);
  and g102 (n134, n72, n82);
  and g103 (n135, n113, n134);
  and g104 (n136, n110, n126);
  not g105 (n_46, n135);
  not g106 (n_47, n136);
  and g107 (n137, n_46, n_47);
  not g110 (n_48, n123);
  not g112 (n_49, n121);
  and g114 (n142, n98, n126);
  and g115 (n143, n79, n97);
  and g116 (n144, n122, n143);
  and g117 (n145, n78, n143);
  and g118 (n146, n104, n126);
  and g119 (n147, n78, n117);
  and g120 (n148, n77, n112);
  and g121 (n149, n117, n148);
  and g122 (n150, n114, n124);
  and g123 (n151, n114, n122);
  and g124 (n152, n101, n134);
  and g125 (n153, n72, n79);
  and g126 (n154, n126, n153);
  and g127 (n155, n117, n124);
  not g128 (n_50, n154);
  not g129 (n_51, n155);
  and g130 (n156, n_50, n_51);
  and g131 (n157, n94, n129);
  and g132 (n158, n83, n148);
  not g133 (n_52, n157);
  not g134 (n_53, n158);
  and g135 (n159, n_52, n_53);
  and g136 (n160, n73, n109);
  and g137 (n161, n94, n160);
  and g138 (n162, n84, n105);
  and g139 (n163, n129, n162);
  and g140 (n164, n85, n143);
  and g141 (n165, n124, n143);
  and g142 (n166, n97, n103);
  and g143 (n167, n124, n166);
  and g144 (n168, n114, n126);
  and g145 (n169, n85, n153);
  and g146 (n170, n129, n148);
  and g147 (n171, n114, n131);
  not g148 (n_54, n170);
  not g149 (n_55, n171);
  and g150 (n172, n_54, n_55);
  and g151 (n173, n88, n143);
  and g152 (n174, n89, n109);
  and g153 (n175, n106, n174);
  and g154 (n176, n84, n87);
  and g155 (n177, n117, n176);
  not g156 (n_56, n175);
  not g157 (n_57, n177);
  and g158 (n178, n_56, n_57);
  not g159 (n_58, n173);
  and g160 (n179, n_58, n178);
  not g162 (n_59, n169);
  not g164 (n_60, n168);
  not g166 (n_61, n167);
  not g168 (n_62, n165);
  not g170 (n_63, n164);
  not g172 (n_64, n163);
  not g174 (n_65, n161);
  and g176 (n188, n80, n124);
  and g177 (n189, n106, n114);
  and g178 (n190, n122, n153);
  and g179 (n191, n98, n162);
  and g180 (n192, n101, n166);
  not g181 (n_66, n191);
  not g182 (n_67, n192);
  and g183 (n193, n_66, n_67);
  and g184 (n194, n110, n113);
  not g185 (n_68, n194);
  not g187 (n_69, n190);
  not g189 (n_70, n189);
  not g191 (n_71, n188);
  and g193 (n199, n73, n103);
  and g194 (n200, n176, n199);
  and g195 (n201, n126, n199);
  not g196 (n_72, n200);
  not g197 (n_73, n201);
  and g198 (n202, n_72, n_73);
  and g199 (n203, n126, n174);
  not g200 (n_74, n203);
  and g201 (n204, n202, n_74);
  and g202 (n205, n94, n143);
  and g203 (n206, n90, n148);
  not g204 (n_75, n205);
  not g205 (n_76, n206);
  and g206 (n207, n_75, n_76);
  not g212 (n_77, n152);
  not g214 (n_78, n151);
  not g216 (n_79, n150);
  not g218 (n_80, n149);
  not g220 (n_81, n147);
  not g222 (n_82, n146);
  not g224 (n_83, n145);
  not g226 (n_84, n144);
  not g228 (n_85, n142);
  and g230 (n222, n80, n85);
  and g231 (n223, n117, n162);
  and g232 (n224, n85, n134);
  and g233 (n225, n88, n199);
  and g234 (n226, n94, n104);
  not g235 (n_86, n225);
  not g236 (n_87, n226);
  and g237 (n227, n_86, n_87);
  and g238 (n228, n90, n122);
  and g239 (n229, n78, n153);
  not g240 (n_88, n228);
  not g241 (n_89, n229);
  and g242 (n230, n_88, n_89);
  and g243 (n231, n80, n106);
  and g244 (n232, n126, n134);
  and g245 (n233, n78, n174);
  not g246 (n_90, n232);
  not g247 (n_91, n233);
  and g248 (n234, n_90, n_91);
  not g249 (n_92, n231);
  and g250 (n235, n_92, n234);
  and g251 (n236, n85, n110);
  and g252 (n237, n148, n199);
  not g253 (n_93, n236);
  not g254 (n_94, n237);
  and g255 (n238, n_93, n_94);
  and g256 (n239, n85, n117);
  and g257 (n240, n143, n148);
  not g258 (n_95, n239);
  not g259 (n_96, n240);
  and g260 (n241, n_95, n_96);
  and g261 (n242, n153, n176);
  and g262 (n243, n143, n176);
  not g263 (n_97, n242);
  not g264 (n_98, n243);
  and g265 (n244, n_97, n_98);
  and g266 (n245, n98, n124);
  and g267 (n246, n126, n166);
  not g268 (n_99, n245);
  not g269 (n_100, n246);
  and g270 (n247, n_99, n_100);
  and g271 (n248, n104, n162);
  and g272 (n249, n80, n131);
  not g273 (n_101, n248);
  not g274 (n_102, n249);
  and g275 (n250, n_101, n_102);
  and g276 (n251, n83, n131);
  and g277 (n252, n106, n199);
  not g278 (n_103, n251);
  not g279 (n_104, n252);
  and g280 (n253, n_103, n_104);
  and g281 (n254, n114, n176);
  and g282 (n255, n106, n134);
  not g283 (n_105, n254);
  not g284 (n_106, n255);
  and g285 (n256, n_105, n_106);
  not g295 (n_107, n224);
  not g297 (n_108, n223);
  not g299 (n_109, n222);
  and g301 (n269, n76, n105);
  and g302 (n270, n80, n269);
  and g303 (n271, n83, n88);
  and g304 (n272, n131, n199);
  and g305 (n273, n126, n129);
  and g306 (n274, n131, n143);
  and g307 (n275, n113, n117);
  and g308 (n276, n110, n131);
  and g309 (n277, n96, n160);
  and g310 (n278, n134, n162);
  not g311 (n_110, n277);
  not g312 (n_111, n278);
  and g313 (n279, n_110, n_111);
  and g314 (n280, n101, n114);
  and g315 (n281, n96, n134);
  not g316 (n_112, n280);
  not g317 (n_113, n281);
  and g318 (n282, n_112, n_113);
  and g319 (n283, n98, n131);
  and g320 (n284, n134, n148);
  not g321 (n_114, n283);
  not g322 (n_115, n284);
  and g323 (n285, n_114, n_115);
  and g324 (n286, n131, n166);
  and g325 (n287, n90, n94);
  not g326 (n_116, n286);
  not g327 (n_117, n287);
  and g328 (n288, n_116, n_117);
  and g329 (n289, n94, n134);
  and g330 (n290, n96, n104);
  not g331 (n_118, n289);
  not g332 (n_119, n290);
  and g333 (n291, n_118, n_119);
  and g334 (n292, n104, n131);
  and g335 (n293, n83, n162);
  not g336 (n_120, n292);
  not g337 (n_121, n293);
  and g338 (n294, n_120, n_121);
  and g339 (n295, n124, n160);
  and g340 (n296, n94, n166);
  not g341 (n_122, n295);
  not g342 (n_123, n296);
  and g343 (n297, n_122, n_123);
  and g344 (n298, n98, n176);
  and g345 (n299, n117, n131);
  not g346 (n_124, n298);
  not g347 (n_125, n299);
  and g348 (n300, n_124, n_125);
  and g349 (n301, n110, n176);
  and g350 (n302, n90, n124);
  not g351 (n_126, n301);
  not g352 (n_127, n302);
  and g353 (n303, n_126, n_127);
  and g354 (n304, n88, n160);
  and g355 (n305, n104, n269);
  and g356 (n306, n129, n269);
  not g357 (n_128, n305);
  not g358 (n_129, n306);
  and g359 (n307, n_128, n_129);
  not g360 (n_130, n304);
  and g361 (n308, n_130, n307);
  not g371 (n_131, n276);
  not g373 (n_132, n275);
  not g375 (n_133, n274);
  not g377 (n_134, n273);
  not g379 (n_135, n272);
  not g381 (n_136, n271);
  not g383 (n_137, n270);
  and g385 (n325, n83, n101);
  and g386 (n326, n90, n162);
  and g387 (n327, n162, n174);
  and g388 (n328, n88, n114);
  and g389 (n329, n78, n134);
  and g390 (n330, n94, n153);
  and g391 (n331, n162, n166);
  and g392 (n332, n160, n269);
  not g393 (n_138, n331);
  not g394 (n_139, n332);
  and g395 (n333, n_138, n_139);
  and g396 (n334, n174, n176);
  and g397 (n335, n94, n114);
  not g398 (n_140, n334);
  not g399 (n_141, n335);
  and g400 (n336, n_140, n_141);
  and g401 (n337, n80, n101);
  and g402 (n338, n85, n199);
  and g403 (n339, n101, n174);
  and g404 (n340, n113, n160);
  not g405 (n_142, n339);
  not g406 (n_143, n340);
  and g407 (n341, n_142, n_143);
  not g408 (n_144, n338);
  and g409 (n342, n_144, n341);
  not g410 (n_145, n337);
  and g411 (n343, n_145, n342);
  not g414 (n_146, n330);
  not g416 (n_147, n329);
  not g418 (n_148, n328);
  not g420 (n_149, n327);
  not g422 (n_150, n326);
  not g424 (n_151, n325);
  and g426 (n352, n122, n174);
  and g427 (n353, n134, n176);
  and g428 (n354, n124, n134);
  and g429 (n355, n134, n269);
  not g430 (n_152, n354);
  not g431 (n_153, n355);
  and g432 (n356, n_152, n_153);
  and g433 (n357, n90, n269);
  and g434 (n358, n83, n269);
  not g435 (n_154, n357);
  not g436 (n_155, n358);
  and g437 (n359, n_154, n_155);
  not g439 (n_156, n353);
  not g441 (n_157, n352);
  and g443 (n363, n80, n94);
  and g444 (n364, n110, n162);
  not g445 (n_158, n363);
  not g446 (n_159, n364);
  and g447 (n365, n_158, n_159);
  and g448 (n366, n96, n199);
  and g449 (n367, n104, n113);
  and g450 (n368, n98, n113);
  not g451 (n_160, n367);
  not g452 (n_161, n368);
  and g453 (n369, n_160, n_161);
  not g454 (n_162, n366);
  and g455 (n370, n_162, n369);
  and g456 (n371, n85, n160);
  and g457 (n372, n88, n98);
  not g458 (n_163, n371);
  not g459 (n_164, n372);
  and g460 (n373, n_163, n_164);
  and g461 (n374, n90, n96);
  and g462 (n375, n78, n129);
  not g463 (n_165, n374);
  not g464 (n_166, n375);
  and g465 (n376, n_165, n_166);
  not g479 (n_167, n91);
  not g481 (n_168, n86);
  not g483 (n_169, n81);
  and g485 (n393, n85, n129);
  and g486 (n394, n124, n129);
  and g487 (n395, n90, n113);
  and g488 (n396, n78, n104);
  and g489 (n397, n106, n110);
  and g490 (n398, n131, n153);
  not g491 (n_170, n398);
  and g492 (n399, n_149, n_170);
  and g493 (n400, n88, n104);
  not g494 (n_171, n400);
  and g495 (n401, n_141, n_171);
  and g496 (n402, n101, n104);
  and g497 (n403, n104, n148);
  not g498 (n_172, n402);
  not g499 (n_173, n403);
  and g500 (n404, n_172, n_173);
  and g501 (n405, n_166, n404);
  not g505 (n_174, n397);
  not g509 (n_175, n396);
  not g511 (n_176, n395);
  and g515 (n416, n78, n90);
  and g516 (n417, n117, n122);
  not g517 (n_177, n417);
  and g518 (n418, n_159, n_177);
  and g519 (n419, n96, n117);
  and g520 (n420, n106, n153);
  not g521 (n_178, n419);
  not g522 (n_179, n420);
  and g523 (n421, n_178, n_179);
  and g524 (n422, n98, n148);
  not g525 (n_180, n422);
  and g526 (n423, n_82, n_180);
  and g527 (n424, n101, n143);
  and g528 (n425, n166, n269);
  and g529 (n426, n114, n148);
  and g530 (n427, n110, n148);
  and g531 (n428, n80, n176);
  and g532 (n429, n80, n148);
  and g533 (n430, n148, n166);
  not g534 (n_181, n430);
  and g535 (n431, n_84, n_181);
  not g537 (n_182, n429);
  not g539 (n_183, n428);
  and g541 (n435, n117, n269);
  and g542 (n436, n160, n176);
  not g543 (n_184, n435);
  not g544 (n_185, n436);
  and g545 (n437, n_184, n_185);
  and g546 (n438, n88, n166);
  not g547 (n_186, n438);
  and g548 (n439, n_163, n_186);
  not g551 (n_187, n427);
  not g554 (n_188, n426);
  not g558 (n_189, n425);
  not g560 (n_190, n424);
  and g562 (n449, n80, n122);
  not g563 (n_191, n449);
  and g564 (n450, n_136, n_191);
  and g565 (n451, n199, n269);
  and g566 (n452, n85, n98);
  and g567 (n453, n98, n101);
  not g568 (n_192, n452);
  not g569 (n_193, n453);
  and g570 (n454, n_192, n_193);
  not g575 (n_194, n451);
  and g577 (n460, n104, n176);
  and g578 (n461, n85, n104);
  and g579 (n462, n148, n153);
  not g580 (n_195, n461);
  not g581 (n_196, n462);
  not g583 (n_197, n460);
  and g586 (n466, n96, n143);
  not g587 (n_198, n466);
  and g588 (n467, n_91, n_198);
  and g589 (n468, n106, n129);
  and g590 (n469, n94, n110);
  and g591 (n470, n94, n199);
  not g592 (n_199, n470);
  and g593 (n471, n_162, n_199);
  not g594 (n_200, n469);
  and g595 (n472, n_200, n471);
  not g596 (n_201, n468);
  and g597 (n473, n_201, n472);
  and g598 (n474, n101, n160);
  not g599 (n_202, n474);
  and g600 (n475, n_71, n_202);
  not g612 (n_203, n416);
  and g615 (n489, n83, n176);
  and g616 (n490, n90, n106);
  not g617 (n_204, n489);
  not g618 (n_205, n490);
  and g619 (n491, n_204, n_205);
  and g620 (n492, n166, n176);
  and g621 (n493, n129, n176);
  not g622 (n_206, n493);
  and g623 (n494, n_61, n_206);
  and g624 (n495, n85, n174);
  and g625 (n496, n78, n166);
  not g626 (n_207, n495);
  not g627 (n_208, n496);
  and g628 (n497, n_207, n_208);
  not g633 (n_209, n492);
  and g636 (n504, n143, n162);
  and g637 (n505, n96, n166);
  and g638 (n506, n96, n174);
  not g639 (n_210, n506);
  and g640 (n507, n_169, n_210);
  and g641 (n508, n_132, n_140);
  and g642 (n509, n101, n153);
  not g643 (n_211, n509);
  and g644 (n510, n_46, n_211);
  and g645 (n511, n114, n269);
  not g646 (n_212, n511);
  and g647 (n512, n_101, n_212);
  and g648 (n513, n104, n124);
  and g649 (n514, n174, n269);
  and g650 (n515, n_129, n_154);
  and g651 (n516, n_65, n515);
  and g652 (n517, n_139, n516);
  and g653 (n518, n96, n153);
  and g654 (n519, n122, n160);
  not g655 (n_213, n518);
  not g656 (n_214, n519);
  and g657 (n520, n_213, n_214);
  not g659 (n_215, n514);
  not g661 (n_216, n513);
  and g664 (n525, n160, n162);
  not g665 (n_217, n525);
  and g666 (n526, n_135, n_217);
  and g667 (n527, n104, n122);
  and g668 (n528, n_39, n_128);
  not g669 (n_218, n527);
  and g670 (n529, n_218, n528);
  and g671 (n530, n_43, n_108);
  and g672 (n531, n101, n199);
  and g673 (n532, n148, n160);
  not g674 (n_219, n532);
  and g675 (n533, n_143, n_219);
  not g676 (n_220, n531);
  and g677 (n534, n_220, n533);
  and g678 (n535, n_144, n534);
  and g679 (n536, n78, n98);
  and g680 (n537, n98, n122);
  not g681 (n_221, n537);
  and g682 (n538, n_161, n_221);
  not g683 (n_222, n536);
  and g684 (n539, n_222, n538);
  and g685 (n540, n_124, n539);
  and g686 (n541, n_155, n540);
  not g699 (n_223, n505);
  not g701 (n_224, n504);
  and g704 (n557, n88, n134);
  and g705 (n558, n88, n110);
  not g706 (n_225, n557);
  not g707 (n_226, n558);
  and g711 (n562, n80, n162);
  and g712 (n563, n85, n166);
  and g713 (n564, n78, n160);
  not g714 (n_227, n563);
  not g715 (n_228, n564);
  and g716 (n565, n_227, n_228);
  not g717 (n_229, n562);
  and g718 (n566, n_229, n565);
  and g719 (n567, n98, n269);
  and g720 (n568, n122, n166);
  and g721 (n569, n83, n122);
  not g722 (n_230, n568);
  not g723 (n_231, n569);
  and g724 (n570, n_230, n_231);
  and g725 (n571, n88, n174);
  not g726 (n_232, n571);
  and g727 (n572, n570, n_232);
  not g728 (n_233, n567);
  and g729 (n573, n_233, n572);
  not g741 (n_234, n394);
  not g743 (n_235, n393);
  not g746 (n_236, n392);
  not g747 (n_237, n587);
  and g748 (n588, n_236, n_237);
  and g749 (n589, n96, n129);
  and g750 (n590, n_71, n_109);
  and g751 (n591, n_68, n_205);
  and g752 (n592, n124, n199);
  not g753 (n_238, n592);
  and g754 (n593, n_88, n_238);
  and g755 (n594, n117, n126);
  not g756 (n_239, n594);
  and g757 (n595, n_75, n_239);
  and g763 (n601, n106, n143);
  and g764 (n602, n114, n162);
  and g765 (n603, n101, n129);
  not g766 (n_240, n603);
  and g767 (n604, n_206, n_240);
  not g769 (n_241, n602);
  not g774 (n_242, n601);
  and g780 (n615, n_78, n_149);
  and g781 (n616, n_89, n376);
  and g782 (n617, n110, n269);
  not g783 (n_243, n617);
  and g784 (n618, n_55, n_243);
  and g785 (n619, n124, n174);
  and g786 (n620, n131, n134);
  not g787 (n_244, n619);
  not g788 (n_245, n620);
  and g789 (n621, n_244, n_245);
  and g790 (n622, n_56, n_217);
  and g791 (n623, n162, n199);
  and g792 (n624, n_46, n_77);
  not g797 (n_246, n623);
  and g801 (n632, n_36, n_97);
  and g802 (n633, n80, n126);
  not g803 (n_247, n633);
  and g804 (n634, n_190, n_247);
  and g805 (n635, n_50, n634);
  and g806 (n636, n_171, n635);
  and g807 (n637, n101, n117);
  not g808 (n_248, n637);
  and g809 (n638, n_232, n_248);
  and g810 (n639, n90, n126);
  not g811 (n_249, n639);
  and g812 (n640, n_223, n_249);
  and g813 (n641, n78, n114);
  not g814 (n_250, n641);
  and g815 (n642, n_209, n_250);
  and g827 (n654, n_48, n_42);
  and g828 (n655, n80, n113);
  and g829 (n656, n94, n174);
  and g830 (n657, n113, n199);
  not g831 (n_251, n657);
  and g832 (n658, n_192, n_251);
  not g836 (n_252, n656);
  not g839 (n_253, n655);
  and g841 (n665, n_114, n_233);
  and g842 (n666, n83, n96);
  and g843 (n667, n153, n162);
  not g844 (n_254, n667);
  not g848 (n_255, n666);
  and g850 (n672, n106, n160);
  and g851 (n673, n143, n269);
  not g852 (n_256, n672);
  not g853 (n_257, n673);
  and g854 (n674, n_256, n_257);
  and g855 (n675, n_84, n_230);
  and g869 (n689, n113, n143);
  not g870 (n_258, n689);
  and g871 (n690, n_69, n_258);
  and g872 (n691, n_147, n_142);
  and g873 (n692, n_179, n_222);
  and g874 (n693, n_201, n692);
  and g875 (n694, n_83, n_105);
  not g891 (n_259, n589);
  not g893 (n_260, n710);
  and g894 (n711, n_237, n_260);
  and g895 (n712, n78, n199);
  and g896 (n713, n122, n134);
  and g897 (n714, n126, n143);
  and g898 (n715, n90, n131);
  and g899 (n716, n113, n166);
  not g902 (n_261, n716);
  and g904 (n720, n_63, n_103);
  and g905 (n721, n_51, n_200);
  and g906 (n722, n_165, n721);
  and g907 (n723, n_81, n_197);
  and g915 (n731, n_83, n_232);
  and g916 (n732, n_163, n_202);
  and g917 (n733, n_58, n_214);
  and g918 (n734, n_53, n733);
  and g919 (n735, n_222, n_252);
  and g930 (n746, n101, n110);
  and g931 (n747, n_76, n_127);
  not g932 (n_262, n746);
  and g937 (n752, n124, n153);
  not g938 (n_263, n752);
  and g939 (n753, n_50, n_263);
  and g940 (n754, n_227, n753);
  not g953 (n_264, n715);
  not g955 (n_265, n714);
  and g959 (n771, n80, n88);
  not g960 (n_266, n771);
  and g961 (n772, n_194, n_266);
  and g962 (n773, n_69, n_96);
  and g963 (n774, n_155, n_172);
  and g964 (n775, n_159, n_187);
  and g965 (n776, n_111, n_148);
  and g966 (n777, n85, n90);
  not g967 (n_267, n777);
  and g968 (n778, n_145, n_267);
  and g978 (n788, n_168, n_206);
  and g979 (n789, n_199, n_254);
  and g980 (n790, n_173, n_216);
  and g981 (n791, n98, n106);
  not g982 (n_268, n791);
  and g983 (n792, n_60, n_268);
  and g984 (n793, n_65, n_99);
  and g994 (n803, n96, n114);
  and g995 (n804, n_150, n_212);
  and g996 (n805, n_207, n_215);
  and g1000 (n809, n113, n174);
  not g1001 (n_269, n809);
  and g1002 (n810, n_181, n_269);
  and g1003 (n811, n_79, n_115);
  and g1004 (n812, n_80, n_177);
  and g1005 (n813, n_246, n_250);
  and g1006 (n814, n_255, n813);
  and g1007 (n815, n_59, n_245);
  and g1008 (n816, n_256, n815);
  and g1017 (n825, n90, n176);
  and g1018 (n826, n_100, n_179);
  and g1019 (n827, n_122, n_228);
  not g1022 (n_270, n825);
  and g1024 (n831, n_224, n_213);
  and g1025 (n832, n_137, n831);
  not g1035 (n_271, n803);
  and g1039 (n845, n120, n654);
  and g1040 (n846, n_70, n845);
  and g1041 (n847, n88, n153);
  not g1042 (n_272, n847);
  and g1043 (n848, n_226, n_272);
  and g1044 (n849, n_108, n848);
  and g1045 (n850, n_243, n849);
  and g1046 (n851, n_156, n850);
  not g1053 (n_273, n713);
  not g1061 (n_274, n712);
  not g1065 (n_275, n867);
  and g1066 (n868, n_260, n_275);
  and g1067 (n869, n_107, n_98);
  and g1071 (n873, n_84, n_273);
  and g1072 (n874, n_93, n_135);
  and g1073 (n875, n80, n96);
  and g1074 (n876, n_126, n_216);
  and g1075 (n877, n_146, n_264);
  not g1080 (n_276, n875);
  and g1082 (n883, n78, n83);
  and g1083 (n884, n106, n117);
  and g1084 (n885, n_168, n_123);
  and g1085 (n886, n83, n113);
  and g1086 (n887, n_188, n_229);
  and g1087 (n888, n_150, n_248);
  and g1088 (n889, n_208, n888);
  not g1093 (n_277, n886);
  and g1096 (n896, n_189, n_204);
  and g1097 (n897, n_144, n_187);
  and g1098 (n898, n_152, n719);
  and g1099 (n899, n_235, n898);
  not g1112 (n_278, n884);
  not g1116 (n_279, n883);
  and g1119 (n917, n_97, n_141);
  and g1120 (n918, n_266, n917);
  and g1134 (n932, n88, n129);
  not g1135 (n_280, n932);
  and g1136 (n933, n_185, n_280);
  and g1140 (n937, n_41, n_186);
  and g1144 (n941, n_81, n_122);
  not g1162 (n_281, n958);
  and g1163 (n959, n_275, n_281);
  and g1164 (n960, n_38, n_105);
  and g1165 (n961, n94, n98);
  not g1166 (n_282, n961);
  and g1167 (n962, n_174, n_282);
  and g1173 (n968, n_169, n_145);
  and g1182 (n977, n_234, n_182);
  and g1183 (n978, n_150, n_249);
  and g1184 (n979, n_156, n_245);
  and g1185 (n980, n106, n166);
  and g1186 (n981, n_74, n_116);
  and g1187 (n982, n_162, n981);
  not g1191 (n_283, n980);
  and g1195 (n989, n_185, n_259);
  and g1196 (n990, n_198, n_206);
  and g1197 (n991, n_80, n_243);
  and g1198 (n992, n_270, n991);
  and g1215 (n1009, n_79, n_104);
  and g1216 (n1010, n131, n160);
  and g1217 (n1011, n113, n153);
  and g1218 (n1012, n_171, n_256);
  not g1220 (n_284, n1011);
  not g1226 (n_285, n1010);
  and g1229 (n1021, n_69, n_107);
  and g1233 (n1025, n_50, n_134);
  and g1237 (n1029, n431, n_271);
  and g1248 (n1040, n_130, n_225);
  and g1253 (n1045, n_47, n282);
  and g1254 (n1046, n_61, n_100);
  and g1255 (n1047, n_64, n1046);
  not g1269 (n_286, n1060);
  and g1270 (n1061, n_281, n_286);
  and g1271 (n1062, n131, n174);
  and g1272 (n1063, n_57, n_203);
  and g1273 (n1064, n_178, n_284);
  and g1274 (n1065, n_145, n1064);
  and g1279 (n1070, n_104, n_211);
  and g1280 (n1071, n_62, n_94);
  and g1281 (n1072, n110, n124);
  not g1282 (n_287, n1072);
  and g1283 (n1073, n_51, n_287);
  and g1295 (n1085, n_133, n_220);
  not g1304 (n_288, n1062);
  and g1312 (n1101, n148, n174);
  and g1313 (n1102, n85, n114);
  not g1314 (n_289, n1102);
  and g1315 (n1103, n_198, n_289);
  and g1316 (n1104, n122, n199);
  not g1317 (n_290, n1104);
  and g1318 (n1105, n_214, n_290);
  and g1319 (n1106, n_240, n1105);
  and g1320 (n1107, n_266, n1106);
  and g1321 (n1108, n_55, n_263);
  and g1322 (n1109, n_274, n1108);
  not g1329 (n_291, n1101);
  and g1334 (n1120, n_95, n_100);
  and g1335 (n1121, n_134, n1120);
  and g1341 (n1127, n126, n160);
  not g1342 (n_292, n1127);
  and g1343 (n1128, n_279, n_292);
  and g1344 (n1129, n_183, n_200);
  and g1345 (n1130, n_78, n_225);
  and g1346 (n1131, n_210, n1130);
  and g1347 (n1132, n_190, n_271);
  and g1354 (n1139, n_75, n_120);
  and g1355 (n1140, n_228, n1139);
  and g1356 (n1141, n_137, n_144);
  and g1357 (n1142, n_132, n1141);
  and g1358 (n1143, n_64, n1142);
  and g1370 (n1155, n_130, n_285);
  and g1374 (n1159, n_35, n_128);
  and g1375 (n1160, n_121, n1159);
  and g1376 (n1161, n_66, n_201);
  and g1377 (n1162, n_113, n1161);
  and g1378 (n1163, n_265, n1162);
  not g1394 (n_293, n1178);
  and g1395 (n1179, n_286, n_293);
  and g1396 (n1180, n_46, n_251);
  and g1397 (n1181, n_77, n_223);
  and g1398 (n1182, n_169, n_147);
  and g1399 (n1183, n_178, n_184);
  and g1400 (n1184, n238, n937);
  and g1401 (n1185, n_68, n1184);
  and g1419 (n1203, n122, n129);
  and g1420 (n1204, n_231, n_283);
  and g1421 (n1205, n_143, n_218);
  and g1422 (n1206, n_276, n1205);
  not g1426 (n_294, n1203);
  and g1437 (n1220, n_180, n_252);
  and g1438 (n1221, n_109, n1220);
  not g1453 (n_295, n1235);
  and g1454 (n1236, n_293, n_295);
  and g1455 (n1237, n_107, n_174);
  and g1464 (n1246, n153, n269);
  and g1465 (n1247, n_133, n_200);
  and g1466 (n1248, n_157, n_291);
  and g1467 (n1249, n_67, n_103);
  and g1468 (n1250, n303, n1249);
  and g1469 (n1251, n_257, n1250);
  and g1470 (n1252, n_163, n_224);
  and g1471 (n1253, n_161, n_266);
  and g1472 (n1254, n_106, n_229);
  and g1473 (n1255, n_35, n_102);
  and g1487 (n1269, n_187, n_191);
  and g1488 (n1270, n_147, n1269);
  and g1489 (n1271, n_278, n1270);
  and g1490 (n1272, n_50, n_215);
  and g1491 (n1273, n533, n_243);
  and g1492 (n1274, n_170, n1273);
  not g1503 (n_296, n1246);
  and g1511 (n1292, n_226, n_271);
  and g1512 (n1293, n_166, n_249);
  and g1513 (n1294, n_134, n1293);
  and g1525 (n1306, n78, n110);
  and g1526 (n1307, n_176, n_258);
  and g1527 (n1308, n_193, n1307);
  not g1528 (n_297, n1306);
  and g1534 (n1314, n_234, n_175);
  and g1535 (n1315, n_194, n1314);
  and g1544 (n1324, n_213, n_230);
  and g1549 (n1329, n_80, n_241);
  and g1550 (n1330, n_272, n_277);
  and g1551 (n1331, n_94, n1330);
  and g1552 (n1332, n_72, n_125);
  and g1553 (n1333, n_65, n1332);
  and g1566 (n1346, n_40, n_152);
  and g1567 (n1347, n_160, n_171);
  not g1585 (n_298, n1364);
  and g1586 (n1365, n_295, n_298);
  and g1587 (n1366, n_86, n_242);
  and g1588 (n1367, n_54, n_134);
  and g1589 (n1368, n_66, n_157);
  and g1590 (n1369, n_135, n1368);
  and g1600 (n1379, n_220, n_297);
  and g1601 (n1380, n_147, n_202);
  and g1609 (n1388, n_138, n_280);
  and g1610 (n1389, n_74, n_195);
  and g1611 (n1390, n_245, n1389);
  and g1612 (n1391, n_214, n1390);
  and g1613 (n1392, n_132, n_166);
  and g1614 (n1393, n_173, n_289);
  and g1615 (n1394, n_72, n1393);
  and g1629 (n1408, n_37, n_264);
  and g1630 (n1409, n_247, n_282);
  and g1644 (n1423, n_167, n_63);
  and g1645 (n1424, n_62, n_207);
  and g1646 (n1425, n_244, n_266);
  and g1647 (n1426, n_131, n_238);
  and g1648 (n1427, n_258, n1426);
  and g1649 (n1428, n_182, n1427);
  and g1657 (n1436, n_176, n_232);
  and g1658 (n1437, n_270, n1436);
  and g1659 (n1438, n_118, n_288);
  and g1660 (n1439, n_241, n_250);
  and g1661 (n1440, n_79, n1439);
  and g1676 (n1455, n454, n1454);
  and g1677 (n1456, n_249, n1455);
  and g1678 (n1457, n_77, n_233);
  and g1679 (n1458, n_65, n1457);
  not g1694 (n_299, n1472);
  and g1695 (n1473, n_298, n_299);
  and g1696 (n1474, n_187, n_230);
  and g1697 (n1475, n_114, n1474);
  and g1698 (n1476, n_90, n_139);
  and g1699 (n1477, n_176, n_203);
  and g1700 (n1478, n_165, n1477);
  and g1701 (n1479, n_208, n_262);
  and g1702 (n1480, n_102, n_253);
  and g1711 (n1489, n_37, n_284);
  and g1712 (n1490, n_54, n1489);
  and g1719 (n1497, n_51, n_269);
  and g1720 (n1498, n_216, n_263);
  and g1721 (n1499, n_189, n1498);
  and g1744 (n1522, n_108, n_229);
  and g1745 (n1523, n_80, n_124);
  and g1746 (n1524, n_82, n_207);
  and g1750 (n1528, n_156, n_175);
  and g1751 (n1529, n_150, n1528);
  and g1752 (n1530, n_191, n1529);
  and g1753 (n1531, n_121, n_255);
  and g1754 (n1532, n1129, n1531);
  and g1755 (n1533, n_261, n1532);
  and g1772 (n1550, n_133, n_226);
  and g1778 (n1556, n_44, n_162);
  and g1779 (n1557, n_136, n_196);
  not g1795 (n_300, n1572);
  and g1796 (n1573, n_299, n_300);
  and g1797 (n1574, n_115, n_219);
  and g1798 (n1575, n_54, n_148);
  and g1799 (n1576, n_85, n_265);
  and g1800 (n1577, n_135, n_294);
  and g1801 (n1578, n_192, n772);
  and g1809 (n1586, n_249, n_251);
  and g1810 (n1587, n_133, n_224);
  and g1811 (n1588, n_73, n1587);
  and g1824 (n1601, n_57, n_93);
  and g1825 (n1602, n_65, n_152);
  and g1826 (n1603, n_69, n_112);
  and g1827 (n1604, n_240, n_284);
  and g1834 (n1611, n_209, n_285);
  and g1839 (n1616, n_38, n_242);
  and g1840 (n1617, n_256, n1616);
  and g1859 (n1636, n_190, n_297);
  and g1867 (n1644, n_88, n_267);
  and g1868 (n1645, n_108, n1254);
  and g1869 (n1646, n_138, n1645);
  not g1889 (n_301, n1665);
  and g1890 (n1666, n_300, n_301);
  and g1891 (n1667, n_45, n_102);
  and g1892 (n1668, n_167, n_196);
  and g1893 (n1669, n_183, n788);
  and g1904 (n1680, n_265, n_290);
  and g1905 (n1681, n_247, n1680);
  and g1916 (n1692, n_182, n_213);
  and g1917 (n1693, n_47, n_125);
  and g1918 (n1694, n_101, n1693);
  and g1919 (n1695, n_202, n1694);
  and g1920 (n1696, n_51, n_161);
  and g1921 (n1697, n_158, n1696);
  and g1933 (n1709, n_198, n_222);
  and g1944 (n1720, n_72, n_192);
  and g1945 (n1721, n_214, n1720);
  and g1950 (n1726, n_56, n_88);
  and g1951 (n1727, n_34, n_255);
  and g1956 (n1732, n_156, n_287);
  and g1960 (n1736, n_205, n1603);
  and g1961 (n1737, n_103, n1736);
  and g1962 (n1738, n_98, n_248);
  and g1963 (n1739, n_37, n_279);
  and g1964 (n1740, n_41, n_207);
  and g1979 (n1755, n_91, n_263);
  and g1984 (n1760, n_90, n_111);
  and g1985 (n1761, n_190, n_258);
  and g1986 (n1762, n_200, n1761);
  and g1987 (n1763, n_107, n1762);
  not g2004 (n_302, n1779);
  and g2005 (n1780, n_301, n_302);
  and g2006 (n1781, n_253, n_270);
  and g2007 (n1782, n_70, n_238);
  and g2008 (n1783, n_50, n_125);
  and g2009 (n1784, n_289, n1783);
  and g2010 (n1785, n_64, n_294);
  and g2020 (n1795, n_157, n_215);
  and g2024 (n1799, n_141, n_244);
  and g2025 (n1800, n_186, n1799);
  and g2049 (n1824, n_42, n_53);
  and g2050 (n1825, n_173, n_241);
  and g2051 (n1826, n_92, n_224);
  and g2052 (n1827, n_198, n_267);
  and g2053 (n1828, n_87, n_291);
  and g2064 (n1839, n_49, n_222);
  and g2083 (n1858, n_249, n1857);
  and g2084 (n1859, n_209, n1858);
  and g2085 (n1860, n_89, n_160);
  and g2086 (n1861, n_202, n1860);
  not g2103 (n_303, n1877);
  and g2104 (n1878, n_302, n_303);
  and g2105 (n1879, n_62, n_192);
  and g2120 (n1894, n_112, n_254);
  and g2121 (n1895, n618, n1894);
  and g2122 (n1896, n_81, n1895);
  and g2123 (n1897, n_53, n_212);
  and g2124 (n1898, n_121, n1897);
  not g2140 (n_304, n1913);
  and g2141 (n1914, n_303, n_304);
  and g2142 (n1915, n_107, n_220);
  and g2143 (n1916, n_95, n_218);
  and g2144 (n1917, n_232, n_246);
  and g2168 (n1941, n_126, n_278);
  and g2169 (n1942, n_165, n1941);
  and g2170 (n1943, n_44, n_125);
  and g2171 (n1944, n_290, n1943);
  and g2186 (n1959, n_200, n_249);
  and g2187 (n1960, n_41, n1959);
  and g2197 (n1970, n_49, n221);
  and g2198 (n1971, n_206, n1970);
  and g2199 (n1972, n418, n1248);
  and g2200 (n1973, n_34, n1972);
  not g2220 (n_305, n1992);
  and g2221 (n1993, n_304, n_305);
  and g2222 (n1994, n_127, n_289);
  and g2223 (n1995, n_60, n_174);
  and g2224 (n1996, n_259, n1995);
  and g2235 (n2007, n_209, n_221);
  and g2239 (n2011, n336, n979);
  and g2240 (n2012, n_164, n2011);
  and g2241 (n2013, n_143, n_284);
  and g2242 (n2014, n_62, n_96);
  and g2249 (n2021, n_64, n_261);
  and g2250 (n2022, n_34, n_262);
  and g2254 (n2026, n_109, n_186);
  not g2286 (n_306, n2057);
  and g2287 (n2058, n_305, n_306);
  and g2288 (n2059, n_77, n_69);
  and g2302 (n2073, n_59, n_248);
  and g2303 (n2074, n_101, n2073);
  and g2304 (n2075, n_290, n2074);
  and g2318 (n2089, n_159, n1129);
  and g2319 (n2090, n_85, n_250);
  and g2320 (n2091, n_158, n_226);
  and g2321 (n2092, n_61, n_210);
  and g2322 (n2093, n_35, n_108);
  and g2334 (n2105, n_215, n_273);
  and g2342 (n2113, n_87, n_211);
  and g2343 (n2114, n_287, n1128);
  and g2344 (n2115, n_82, n2114);
  and g2362 (n2133, n_216, n_288);
  not g2382 (n_307, n2152);
  and g2383 (n2153, n_306, n_307);
  and g2384 (n2154, n_40, n_287);
  and g2398 (n2168, n_209, n_215);
  and g2399 (n2169, n_217, n2168);
  and g2400 (n2170, n_235, n_283);
  and g2401 (n2171, n356, n2170);
  and g2402 (n2172, n_197, n2171);
  and g2403 (n2173, n156, n1893);
  and g2404 (n2174, n_56, n2173);
  and g2405 (n2175, n747, n773);
  and g2406 (n2176, n1141, n2175);
  not g2420 (n_308, n2189);
  and g2421 (n2190, n_307, n_308);
  and g2422 (n2191, n_52, n_131);
  and g2423 (n2192, n_84, n_291);
  and g2440 (n2209, n_265, n_282);
  and g2441 (n2210, n_81, n_67);
  and g2449 (n2218, n_68, n_244);
  and g2450 (n2219, n_270, n2218);
  and g2451 (n2220, n_134, n_210);
  and g2461 (n2230, n_93, n_197);
  and g2472 (n2241, n_37, n_227);
  and g2494 (n2263, n_262, n_269);
  and g2495 (n2264, n_65, n202);
  and g2496 (n2265, n_256, n2264);
  and g2497 (n2266, n526, n732);
  and g2498 (n2267, n_94, n2266);
  and g2505 (n2274, n_86, n2273);
  and g2506 (n2275, n_53, n2274);
  and g2507 (n2276, n_208, n_242);
  and g2508 (n2277, n_77, n2276);
  and g2509 (n2278, n_154, n2277);
  not g2523 (n_309, n2291);
  and g2524 (n2292, n_308, n_309);
  and g2525 (n2293, n_98, n_160);
  and g2529 (n2297, n_82, n_197);
  and g2534 (n2302, n1131, n1476);
  and g2535 (n2303, n_262, n2302);
  and g2563 (n2331, n_242, n_254);
  and g2564 (n2332, n_145, n2331);
  and g2565 (n2333, n_61, n_138);
  and g2566 (n2334, n_104, n2333);
  and g2578 (n2346, n_227, n_257);
  and g2579 (n2347, n_56, n2346);
  and g2580 (n2348, n_201, n_282);
  and g2581 (n2349, n_259, n_296);
  and g2593 (n2361, n_127, n_219);
  and g2594 (n2362, n_167, n_213);
  and g2595 (n2363, n_85, n2362);
  and g2603 (n2371, n_148, n_231);
  not g2621 (n_310, n2388);
  and g2622 (n2389, n_309, n_310);
  and g2623 (n2390, n_58, n_228);
  and g2639 (n2406, n_35, n_194);
  and g2643 (n2410, n_81, n_136);
  and g2656 (n2423, n_41, n_85);
  and g2657 (n2424, n_108, n_178);
  and g2658 (n2425, n_101, n_288);
  and g2659 (n2426, n_161, n2425);
  and g2660 (n2427, n156, n_280);
  and g2673 (n2440, n288, n2439);
  and g2674 (n2441, n_182, n2440);
  and g2675 (n2442, n_126, n_274);
  and g2676 (n2443, n_268, n2442);
  and g2677 (n2444, n_189, n2443);
  and g2678 (n2445, n_251, n2444);
  not g2698 (n_311, n2464);
  and g2699 (n2465, n_310, n_311);
  and g2700 (n2466, n_106, n_243);
  and g2701 (n2467, n_128, n_194);
  and g2702 (n2468, n_162, n_258);
  and g2703 (n2469, n202, n_207);
  and g2704 (n2470, n_104, n2469);
  and g2718 (n2484, n_61, n_181);
  and g2741 (n2507, n_64, n_296);
  and g2742 (n2508, n_179, n_224);
  not g2768 (n_312, n2533);
  and g2769 (n2534, n_311, n_312);
  and g2779 (n2544, n_170, n_239);
  and g2780 (n2545, n_97, n_223);
  and g2781 (n2546, n_52, n2545);
  and g2791 (n2556, n_95, n_247);
  not g2807 (n_313, n2571);
  and g2808 (n2572, n_312, n_313);
  and g2809 (n2573, n_151, n_279);
  and g2818 (n2582, n_158, n_276);
  and g2819 (n2583, n_211, n_246);
  and g2820 (n2584, n_170, n_201);
  and g2828 (n2592, n_96, n_99);
  and g2829 (n2593, n_294, n2592);
  and g2830 (n2594, n873, n1180);
  and g2831 (n2595, n_34, n2594);
  and g2842 (n2606, n_59, n_221);
  and g2843 (n2607, n_217, n2606);
  and g2844 (n2608, n_195, n_224);
  and g2860 (n2624, n_212, n616);
  and g2861 (n2625, n_44, n2624);
  and g2862 (n2626, n_68, n_226);
  and g2863 (n2627, n_265, n2626);
  and g2869 (n2633, n_48, n_235);
  and g2870 (n2634, n_57, n_73);
  and g2871 (n2635, n_104, n2634);
  and g2872 (n2636, n_76, n2635);
  and g2873 (n2637, n_155, n2636);
  and g2887 (n2651, n_167, n_223);
  and g2888 (n2652, n282, n2651);
  and g2889 (n2653, n_218, n2652);
  not g2911 (n_314, n2674);
  and g2912 (n2675, n_313, n_314);
  and g2920 (n2683, n_109, n_117);
  and g2921 (n2684, n_39, n2683);
  and g2935 (n2698, n_180, n_217);
  and g2941 (n2704, n_242, n_276);
  and g2942 (n2705, n_56, n_122);
  and g2957 (n2720, n_106, n_227);
  and g2958 (n2721, n_168, n2720);
  not g2974 (n_315, n2736);
  and g2975 (n2737, n_314, n_315);
  and g2976 (n2738, n_89, n_296);
  and g2977 (n2739, n_140, n_252);
  and g2978 (n2740, n_78, n_55);
  and g2979 (n2741, n_153, n804);
  and g2980 (n2742, n_276, n2741);
  and g2990 (n2752, n_185, n_233);
  and g2991 (n2753, n_171, n520);
  and g2996 (n2758, n_77, n_243);
  and g2997 (n2759, n_40, n2758);
  and g2998 (n2760, n1314, n2759);
  and g3021 (n2783, n418, n_209);
  and g3022 (n2784, n_99, n2783);
  and g3045 (n2807, n_45, n_151);
  and g3046 (n2808, n_68, n_277);
  and g3047 (n2809, n_121, n_164);
  and g3048 (n2810, n_63, n2073);
  and g3049 (n2811, n_110, n2810);
  and g3068 (n2830, n2674, n_315);
  not g3069 (n_316, n2829);
  and g3070 (n2831, n_316, n2830);
  not g3071 (n_317, n2737);
  not g3072 (n_318, n2831);
  and g3073 (n2832, n_317, n_318);
  and g3074 (n2833, n2571, n2674);
  not g3075 (n_319, n2675);
  not g3076 (n_320, n2833);
  and g3077 (n2834, n_319, n_320);
  not g3078 (n_321, n2832);
  and g3079 (n2835, n_321, n2834);
  not g3080 (n_322, n2835);
  and g3081 (n2836, n_319, n_322);
  and g3082 (n2837, n2533, n2571);
  not g3083 (n_323, n2572);
  not g3084 (n_324, n2837);
  and g3085 (n2838, n_323, n_324);
  not g3086 (n_325, n2836);
  and g3087 (n2839, n_325, n2838);
  not g3088 (n_326, n2839);
  and g3089 (n2840, n_323, n_326);
  and g3090 (n2841, n2464, n2533);
  not g3091 (n_327, n2534);
  not g3092 (n_328, n2841);
  and g3093 (n2842, n_327, n_328);
  not g3094 (n_329, n2840);
  and g3095 (n2843, n_329, n2842);
  not g3096 (n_330, n2843);
  and g3097 (n2844, n_327, n_330);
  and g3098 (n2845, n2388, n2464);
  not g3099 (n_331, n2465);
  not g3100 (n_332, n2845);
  and g3101 (n2846, n_331, n_332);
  not g3102 (n_333, n2844);
  and g3103 (n2847, n_333, n2846);
  not g3104 (n_334, n2847);
  and g3105 (n2848, n_331, n_334);
  and g3106 (n2849, n2291, n2388);
  not g3107 (n_335, n2389);
  not g3108 (n_336, n2849);
  and g3109 (n2850, n_335, n_336);
  not g3110 (n_337, n2848);
  and g3111 (n2851, n_337, n2850);
  not g3112 (n_338, n2851);
  and g3113 (n2852, n_335, n_338);
  and g3114 (n2853, n2189, n2291);
  not g3115 (n_339, n2292);
  not g3116 (n_340, n2853);
  and g3117 (n2854, n_339, n_340);
  not g3118 (n_341, n2852);
  and g3119 (n2855, n_341, n2854);
  not g3120 (n_342, n2855);
  and g3121 (n2856, n_339, n_342);
  and g3122 (n2857, n2152, n2189);
  not g3123 (n_343, n2190);
  not g3124 (n_344, n2857);
  and g3125 (n2858, n_343, n_344);
  not g3126 (n_345, n2856);
  and g3127 (n2859, n_345, n2858);
  not g3128 (n_346, n2859);
  and g3129 (n2860, n_343, n_346);
  and g3130 (n2861, n2057, n2152);
  not g3131 (n_347, n2153);
  not g3132 (n_348, n2861);
  and g3133 (n2862, n_347, n_348);
  not g3134 (n_349, n2860);
  and g3135 (n2863, n_349, n2862);
  not g3136 (n_350, n2863);
  and g3137 (n2864, n_347, n_350);
  and g3138 (n2865, n1992, n2057);
  not g3139 (n_351, n2058);
  not g3140 (n_352, n2865);
  and g3141 (n2866, n_351, n_352);
  not g3142 (n_353, n2864);
  and g3143 (n2867, n_353, n2866);
  not g3144 (n_354, n2867);
  and g3145 (n2868, n_351, n_354);
  and g3146 (n2869, n1913, n1992);
  not g3147 (n_355, n1993);
  not g3148 (n_356, n2869);
  and g3149 (n2870, n_355, n_356);
  not g3150 (n_357, n2868);
  and g3151 (n2871, n_357, n2870);
  not g3152 (n_358, n2871);
  and g3153 (n2872, n_355, n_358);
  and g3154 (n2873, n1877, n1913);
  not g3155 (n_359, n1914);
  not g3156 (n_360, n2873);
  and g3157 (n2874, n_359, n_360);
  not g3158 (n_361, n2872);
  and g3159 (n2875, n_361, n2874);
  not g3160 (n_362, n2875);
  and g3161 (n2876, n_359, n_362);
  and g3162 (n2877, n1779, n1877);
  not g3163 (n_363, n1878);
  not g3164 (n_364, n2877);
  and g3165 (n2878, n_363, n_364);
  not g3166 (n_365, n2876);
  and g3167 (n2879, n_365, n2878);
  not g3168 (n_366, n2879);
  and g3169 (n2880, n_363, n_366);
  and g3170 (n2881, n1665, n1779);
  not g3171 (n_367, n1780);
  not g3172 (n_368, n2881);
  and g3173 (n2882, n_367, n_368);
  not g3174 (n_369, n2880);
  and g3175 (n2883, n_369, n2882);
  not g3176 (n_370, n2883);
  and g3177 (n2884, n_367, n_370);
  and g3178 (n2885, n1572, n1665);
  not g3179 (n_371, n1666);
  not g3180 (n_372, n2885);
  and g3181 (n2886, n_371, n_372);
  not g3182 (n_373, n2884);
  and g3183 (n2887, n_373, n2886);
  not g3184 (n_374, n2887);
  and g3185 (n2888, n_371, n_374);
  and g3186 (n2889, n1472, n1572);
  not g3187 (n_375, n1573);
  not g3188 (n_376, n2889);
  and g3189 (n2890, n_375, n_376);
  not g3190 (n_377, n2888);
  and g3191 (n2891, n_377, n2890);
  not g3192 (n_378, n2891);
  and g3193 (n2892, n_375, n_378);
  and g3194 (n2893, n1364, n1472);
  not g3195 (n_379, n1473);
  not g3196 (n_380, n2893);
  and g3197 (n2894, n_379, n_380);
  not g3198 (n_381, n2892);
  and g3199 (n2895, n_381, n2894);
  not g3200 (n_382, n2895);
  and g3201 (n2896, n_379, n_382);
  and g3202 (n2897, n1235, n1364);
  not g3203 (n_383, n1365);
  not g3204 (n_384, n2897);
  and g3205 (n2898, n_383, n_384);
  not g3206 (n_385, n2896);
  and g3207 (n2899, n_385, n2898);
  not g3208 (n_386, n2899);
  and g3209 (n2900, n_383, n_386);
  and g3210 (n2901, n1178, n1235);
  not g3211 (n_387, n1236);
  not g3212 (n_388, n2901);
  and g3213 (n2902, n_387, n_388);
  not g3214 (n_389, n2900);
  and g3215 (n2903, n_389, n2902);
  not g3216 (n_390, n2903);
  and g3217 (n2904, n_387, n_390);
  and g3218 (n2905, n1060, n1178);
  not g3219 (n_391, n1179);
  not g3220 (n_392, n2905);
  and g3221 (n2906, n_391, n_392);
  not g3222 (n_393, n2904);
  and g3223 (n2907, n_393, n2906);
  not g3224 (n_394, n2907);
  and g3225 (n2908, n_391, n_394);
  and g3226 (n2909, n958, n1060);
  not g3227 (n_395, n1061);
  not g3228 (n_396, n2909);
  and g3229 (n2910, n_395, n_396);
  not g3230 (n_397, n2908);
  and g3231 (n2911, n_397, n2910);
  not g3232 (n_398, n2911);
  and g3233 (n2912, n_395, n_398);
  and g3234 (n2913, n867, n958);
  not g3235 (n_399, n959);
  not g3236 (n_400, n2913);
  and g3237 (n2914, n_399, n_400);
  not g3238 (n_401, n2912);
  and g3239 (n2915, n_401, n2914);
  not g3240 (n_402, n2915);
  and g3241 (n2916, n_399, n_402);
  and g3242 (n2917, n710, n867);
  not g3243 (n_403, n868);
  not g3244 (n_404, n2917);
  and g3245 (n2918, n_403, n_404);
  not g3246 (n_405, n2916);
  and g3247 (n2919, n_405, n2918);
  not g3248 (n_406, n2919);
  and g3249 (n2920, n_403, n_406);
  and g3250 (n2921, n587, n710);
  not g3251 (n_407, n711);
  not g3252 (n_408, n2921);
  and g3253 (n2922, n_407, n_408);
  not g3254 (n_409, n2920);
  and g3255 (n2923, n_409, n2922);
  not g3256 (n_410, n2923);
  and g3257 (n2924, n_407, n_410);
  and g3258 (n2925, n392, n587);
  not g3259 (n_411, n588);
  not g3260 (n_412, n2925);
  and g3261 (n2926, n_411, n_412);
  not g3262 (n_413, n2924);
  and g3263 (n2927, n_413, n2926);
  not g3264 (n_414, n2927);
  and g3265 (n2928, n_411, n_414);
  and g3299 (n2962, n_273, n1760);
  and g3300 (n2963, n_113, n2962);
  and g3328 (n2991, n_157, n421);
  and g3329 (n2992, n_144, n2991);
  and g3330 (n2993, n_49, n_57);
  and g3331 (n2994, n_170, n2993);
  and g3332 (n2995, n_39, n2994);
  not g3350 (n_415, n3012);
  and g3351 (n3013, n_236, n_415);
  and g3352 (n3014, n392, n3012);
  not g3353 (n_416, n3013);
  not g3354 (n_417, n3014);
  and g3355 (n3015, n_416, n_417);
  not g3356 (n_418, n2928);
  and g3357 (n3016, n_418, n3015);
  not g3358 (n_419, n3015);
  and g3359 (n3017, n2928, n_419);
  not g3360 (n_420, n3016);
  not g3361 (n_421, n3017);
  and g3362 (n3018, n_420, n_421);
  and g3363 (n3019, n75, n3018);
  not g3364 (n_422, \a[31] );
  and g3365 (n3020, n_422, n_21);
  and g3366 (n3021, n_415, n3020);
  and g3367 (n3022, \a[30] , n74);
  and g3368 (n3023, \a[31] , n3022);
  and g3369 (n3024, n_237, n3023);
  and g3370 (n3025, \a[30] , n_422);
  and g3371 (n3026, n_17, \a[31] );
  not g3372 (n_423, n3025);
  not g3373 (n_424, n3026);
  and g3374 (n3027, n_423, n_424);
  not g3375 (n_425, n3027);
  and g3376 (n3028, n74, n_425);
  and g3377 (n3029, n_236, n3028);
  and g3392 (n3040, n_116, n_193);
  and g3393 (n3041, n_151, n_292);
  and g3394 (n3042, n_71, n_252);
  and g3395 (n3043, n_69, n_218);
  and g3396 (n3044, n_171, n_273);
  and g3397 (n3045, n_66, n3044);
  and g3410 (n3058, n_250, n_263);
  and g3411 (n3059, n_248, n3058);
  and g3436 (n3084, n_74, n_268);
  and g3437 (n3085, n_219, n3084);
  and g3466 (n3114, n_132, n2347);
  and g3467 (n3115, n_60, n968);
  and g3480 (n3128, n618, n_272);
  and g3499 (n3147, n_140, n_196);
  and g3500 (n3148, n_220, n3147);
  and g3512 (n3160, n_151, n_271);
  and g3513 (n3161, n_274, n747);
  and g3514 (n3162, n_285, n3161);
  and g3515 (n3163, n_60, n_189);
  and g3516 (n3164, n_202, n3163);
  and g3517 (n3165, n_109, n3164);
  and g3544 (n3192, n507, n_284);
  and g3545 (n3193, n_131, n_146);
  and g3546 (n3194, n_77, n3193);
  and g3558 (n3206, n_107, n_147);
  and g3578 (n3226, n_91, n_176);
  not g3592 (n_430, n3146);
  not g3593 (n_431, n3239);
  and g3594 (n3240, n_430, n_431);
  and g3595 (n3241, n3146, n3239);
  not g3596 (n_432, n3240);
  not g3597 (n_433, n3241);
  and g3598 (n3242, n_432, n_433);
  not g3599 (n_435, \a[20] );
  and g3600 (n3243, n_435, n3242);
  not g3601 (n_436, n3243);
  and g3602 (n3244, n_432, n_436);
  not g3603 (n_437, n3244);
  and g3604 (n3245, n3083, n_437);
  not g3605 (n_438, n3083);
  and g3606 (n3246, n_438, n3244);
  not g3607 (n_439, n3245);
  not g3608 (n_440, n3246);
  and g3609 (n3247, n_439, n_440);
  not g3610 (n_441, n3032);
  and g3611 (n3248, n_441, n3247);
  not g3612 (n_442, n3248);
  and g3613 (n3249, n_441, n_442);
  and g3614 (n3250, n3247, n_442);
  not g3615 (n_443, n3249);
  not g3616 (n_444, n3250);
  and g3617 (n3251, n_443, n_444);
  and g3618 (n3252, n_58, n_87);
  and g3626 (n3260, n_106, n1394);
  and g3627 (n3261, n_134, n3260);
  and g3631 (n3265, n_136, n471);
  and g3632 (n3266, n_158, n3265);
  and g3633 (n3267, n1063, n1128);
  and g3634 (n3268, n_86, n3267);
  and g3663 (n3297, n_75, n2651);
  and g3664 (n3298, n_109, n3297);
  and g3665 (n3299, n_176, n_192);
  and g3666 (n3300, n_204, n3299);
  and g3679 (n3313, n_174, n_184);
  and g3680 (n3314, n_186, n3313);
  not g3694 (n_445, n3327);
  and g3695 (n3328, n3146, n_445);
  and g3696 (n3329, n_430, n3327);
  not g3697 (n_446, n2922);
  and g3698 (n3330, n2920, n_446);
  not g3699 (n_447, n3330);
  and g3700 (n3331, n_410, n_447);
  and g3701 (n3332, n75, n3331);
  and g3702 (n3333, n_237, n3020);
  and g3703 (n3334, n_275, n3023);
  and g3704 (n3335, n_260, n3028);
  not g3712 (n_452, n3328);
  not g3713 (n_453, n3338);
  and g3714 (n3339, n_452, n_453);
  not g3715 (n_454, n3329);
  and g3716 (n3340, n_454, n3339);
  not g3717 (n_455, n3340);
  and g3718 (n3341, n_452, n_455);
  and g3719 (n3342, n_435, n_436);
  and g3720 (n3343, n_433, n3244);
  not g3721 (n_456, n3342);
  not g3722 (n_457, n3343);
  and g3723 (n3344, n_456, n_457);
  not g3724 (n_458, n3341);
  not g3725 (n_459, n3344);
  and g3726 (n3345, n_458, n_459);
  not g3727 (n_460, n2926);
  and g3728 (n3346, n2924, n_460);
  not g3729 (n_461, n3346);
  and g3730 (n3347, n_414, n_461);
  and g3731 (n3348, n75, n3347);
  and g3732 (n3349, n_236, n3020);
  and g3733 (n3350, n_260, n3023);
  and g3734 (n3351, n_237, n3028);
  and g3742 (n3355, n3341, n3344);
  not g3743 (n_466, n3345);
  not g3744 (n_467, n3355);
  and g3745 (n3356, n_466, n_467);
  not g3746 (n_468, n3354);
  and g3747 (n3357, n_468, n3356);
  not g3748 (n_469, n3357);
  and g3749 (n3358, n_466, n_469);
  not g3750 (n_470, n3251);
  not g3751 (n_471, n3358);
  and g3752 (n3359, n_470, n_471);
  and g3753 (n3360, n3251, n3358);
  not g3754 (n_472, n3359);
  not g3755 (n_473, n3360);
  and g3756 (n3361, n_472, n_473);
  and g3757 (n3362, \a[28] , n_15);
  and g3758 (n3363, n_32, \a[29] );
  not g3759 (n_474, n3362);
  not g3760 (n_475, n3363);
  and g3761 (n3364, n_474, n_475);
  and g3762 (n3365, \a[26] , n_31);
  and g3763 (n3366, n_33, \a[27] );
  not g3764 (n_476, n3365);
  not g3765 (n_477, n3366);
  and g3766 (n3367, n_476, n_477);
  not g3767 (n_478, n3364);
  not g3768 (n_479, n3367);
  and g3769 (n3368, n_478, n_479);
  and g3770 (n3369, n_200, n_252);
  and g3771 (n3370, n_285, n3369);
  and g3780 (n3379, n_82, n_222);
  and g3781 (n3380, n_183, n3379);
  and g3791 (n3390, n_164, n_187);
  and g3792 (n3391, n_139, n3390);
  and g3793 (n3392, n937, n1181);
  and g3794 (n3393, n_250, n3392);
  and g3810 (n3409, n_105, n_141);
  and g3817 (n3416, n116, n515);
  and g3837 (n3436, n_230, n_261);
  and g3838 (n3437, n_85, n3436);
  and g3839 (n3438, n_168, n_96);
  and g3858 (n3457, n3364, n_479);
  not g3859 (n_480, n3456);
  and g3860 (n3458, n_480, n3457);
  and g3861 (n3459, n_41, n_136);
  and g3873 (n3471, n_138, n2105);
  and g3874 (n3472, n_193, n3471);
  and g3875 (n3473, n418, n_200);
  and g3876 (n3474, n_202, n3473);
  and g3892 (n3490, n_52, n_232);
  and g3913 (n3511, n_101, n_188);
  and g3914 (n3512, n_264, n3511);
  and g3915 (n3513, n968, n_288);
  and g3916 (n3514, n_189, n3513);
  and g3924 (n3522, n_49, n_83);
  and g3925 (n3523, n_144, n3522);
  and g3926 (n3524, n_116, n_139);
  not g3942 (n_481, n79);
  not g3943 (n_482, n82);
  and g3944 (n3540, n_481, n_482);
  and g3945 (n3541, n_478, n3367);
  not g3946 (n_483, n3540);
  and g3947 (n3542, n_483, n3541);
  not g3948 (n_484, n3539);
  and g3949 (n3543, n_484, n3542);
  and g3950 (n3544, n_91, n_278);
  and g3955 (n3549, n_87, n_292);
  and g3976 (n3570, n_183, n2582);
  and g3987 (n3581, n_153, n_188);
  and g3988 (n3582, n_175, n3581);
  and g3989 (n3583, n_199, n3582);
  and g4012 (n3606, n3367, n3540);
  not g4013 (n_485, n3605);
  and g4014 (n3607, n_485, n3606);
  not g4015 (n_486, n3543);
  not g4016 (n_487, n3607);
  and g4017 (n3608, n_486, n_487);
  not g4018 (n_488, n3458);
  and g4019 (n3609, n_488, n3608);
  not g4020 (n_489, n3368);
  and g4021 (n3610, n_489, n3609);
  and g4022 (n3611, n_484, n_485);
  and g4023 (n3612, n_415, n_484);
  and g4024 (n3613, n_416, n_420);
  and g4025 (n3614, n3012, n3539);
  not g4026 (n_490, n3612);
  not g4027 (n_491, n3614);
  and g4028 (n3615, n_490, n_491);
  not g4029 (n_492, n3613);
  and g4030 (n3616, n_492, n3615);
  not g4031 (n_493, n3616);
  and g4032 (n3617, n_490, n_493);
  and g4033 (n3618, n3539, n3605);
  not g4034 (n_494, n3611);
  not g4035 (n_495, n3618);
  and g4036 (n3619, n_494, n_495);
  not g4037 (n_496, n3617);
  and g4038 (n3620, n_496, n3619);
  not g4039 (n_497, n3620);
  and g4040 (n3621, n_494, n_497);
  and g4041 (n3622, n_480, n_485);
  and g4042 (n3623, n3456, n3605);
  not g4043 (n_498, n3622);
  not g4044 (n_499, n3623);
  and g4045 (n3624, n_498, n_499);
  not g4046 (n_500, n3621);
  and g4047 (n3625, n_500, n3624);
  not g4048 (n_501, n3624);
  and g4049 (n3626, n3621, n_501);
  not g4050 (n_502, n3625);
  not g4051 (n_503, n3626);
  and g4052 (n3627, n_502, n_503);
  not g4053 (n_504, n3627);
  and g4054 (n3628, n3609, n_504);
  not g4055 (n_505, n3610);
  not g4056 (n_506, n3628);
  and g4057 (n3629, n_505, n_506);
  not g4058 (n_507, n3629);
  and g4059 (n3630, \a[29] , n_507);
  and g4060 (n3631, n_15, n3629);
  not g4061 (n_508, n3630);
  not g4062 (n_509, n3631);
  and g4063 (n3632, n_508, n_509);
  not g4064 (n_510, n3632);
  and g4065 (n3633, n3361, n_510);
  not g4066 (n_511, n3633);
  and g4067 (n3634, n_472, n_511);
  and g4068 (n3635, n_439, n_442);
  and g4069 (n3636, n_244, n1531);
  and g4078 (n3645, n_45, n_64);
  and g4119 (n3686, n_206, n1380);
  and g4120 (n3687, n_285, n3686);
  not g4136 (n_512, n3702);
  and g4137 (n3703, n3083, n_512);
  and g4138 (n3704, n_438, n3702);
  not g4139 (n_513, n3635);
  not g4140 (n_514, n3704);
  and g4141 (n3705, n_513, n_514);
  not g4142 (n_515, n3703);
  and g4143 (n3706, n_515, n3705);
  not g4144 (n_516, n3706);
  and g4145 (n3707, n_513, n_516);
  and g4146 (n3708, n_514, n_516);
  and g4147 (n3709, n_515, n3708);
  not g4148 (n_517, n3707);
  not g4149 (n_518, n3709);
  and g4150 (n3710, n_517, n_518);
  and g4151 (n3711, n3020, n_484);
  and g4152 (n3712, n_415, n3028);
  and g4153 (n3713, n_236, n3023);
  not g4154 (n_519, n3615);
  and g4155 (n3714, n3613, n_519);
  not g4156 (n_520, n3714);
  and g4157 (n3715, n_493, n_520);
  and g4158 (n3716, n75, n3715);
  not g4166 (n_525, n3710);
  not g4167 (n_526, n3719);
  and g4168 (n3720, n_525, n_526);
  not g4169 (n_527, n3720);
  and g4170 (n3721, n_525, n_527);
  and g4171 (n3722, n_526, n_527);
  not g4172 (n_528, n3721);
  not g4173 (n_529, n3722);
  and g4174 (n3723, n_528, n_529);
  not g4175 (n_530, n3634);
  not g4176 (n_531, n3723);
  and g4177 (n3724, n_530, n_531);
  not g4178 (n_532, n3724);
  and g4179 (n3725, n_530, n_532);
  and g4180 (n3726, n_531, n_532);
  not g4181 (n_533, n3725);
  not g4182 (n_534, n3726);
  and g4183 (n3727, n_533, n_534);
  and g4184 (n3728, n_70, n_112);
  and g4185 (n3729, n_39, n3728);
  and g4247 (n3791, n_84, n_198);
  and g4248 (n3792, n_66, n3791);
  not g4262 (n_535, n3805);
  and g4263 (n3806, n3457, n_535);
  and g4264 (n3807, n3542, n_485);
  and g4265 (n3808, n_480, n3606);
  not g4266 (n_536, n3807);
  not g4267 (n_537, n3808);
  and g4268 (n3809, n_536, n_537);
  not g4269 (n_538, n3806);
  and g4270 (n3810, n_538, n3809);
  and g4271 (n3811, n_489, n3810);
  and g4272 (n3812, n_498, n_502);
  and g4273 (n3813, n_480, n_535);
  and g4274 (n3814, n3456, n3805);
  not g4275 (n_539, n3813);
  not g4276 (n_540, n3814);
  and g4277 (n3815, n_539, n_540);
  not g4278 (n_541, n3812);
  and g4279 (n3816, n_541, n3815);
  not g4280 (n_542, n3815);
  and g4281 (n3817, n3812, n_542);
  not g4282 (n_543, n3816);
  not g4283 (n_544, n3817);
  and g4284 (n3818, n_543, n_544);
  not g4285 (n_545, n3818);
  and g4286 (n3819, n3810, n_545);
  not g4287 (n_546, n3811);
  not g4288 (n_547, n3819);
  and g4289 (n3820, n_546, n_547);
  not g4290 (n_548, n3820);
  and g4291 (n3821, \a[29] , n_548);
  and g4292 (n3822, n_15, n3820);
  not g4293 (n_549, n3821);
  not g4294 (n_550, n3822);
  and g4295 (n3823, n_549, n_550);
  and g4296 (n3824, n3727, n3823);
  not g4297 (n_551, n3727);
  not g4298 (n_552, n3823);
  and g4299 (n3825, n_551, n_552);
  not g4300 (n_553, n3824);
  not g4301 (n_554, n3825);
  and g4302 (n3826, n_553, n_554);
  and g4303 (n3827, n_116, n_186);
  and g4308 (n3832, n_124, n_282);
  and g4333 (n3857, n_182, n590);
  and g4334 (n3858, n_92, n3857);
  and g4350 (n3874, n3856, n3873);
  and g4354 (n3878, \a[23] , n_24);
  and g4355 (n3879, n_27, \a[24] );
  not g4356 (n_555, n3878);
  not g4357 (n_556, n3879);
  and g4358 (n3880, n_555, n_556);
  and g4359 (n3881, \a[25] , n_33);
  and g4360 (n3882, n_25, \a[26] );
  not g4361 (n_557, n3881);
  not g4362 (n_558, n3882);
  and g4363 (n3883, n_557, n_558);
  not g4364 (n_559, n3880);
  and g4365 (n3884, n_559, n3883);
  not g4366 (n_560, n3877);
  and g4367 (n3885, n_560, n3884);
  and g4368 (n3886, n_43, n_110);
  and g4388 (n3906, n747, n978);
  and g4395 (n3913, n775, n3912);
  and g4396 (n3914, n_287, n3913);
  and g4412 (n3930, n_146, n2738);
  and g4413 (n3931, n_97, n3930);
  and g4430 (n3948, n_164, n1480);
  and g4431 (n3949, n_191, n3948);
  not g4447 (n_561, n76);
  not g4448 (n_562, n84);
  and g4449 (n3965, n_561, n_562);
  not g4450 (n_563, n3883);
  and g4451 (n3966, n3880, n_563);
  not g4452 (n_564, n3965);
  and g4453 (n3967, n_564, n3966);
  not g4454 (n_565, n3964);
  and g4455 (n3968, n_565, n3967);
  and g4472 (n3985, n_119, n_278);
  and g4473 (n3986, n_81, n3985);
  and g4474 (n3987, n_173, n3986);
  and g4497 (n4010, n_132, n2993);
  and g4498 (n4011, n_177, n4010);
  and g4533 (n4046, n3880, n3965);
  not g4534 (n_566, n4045);
  and g4535 (n4047, n_566, n4046);
  and g4541 (n4050, n_559, n_563);
  and g4542 (n4051, n_565, n_566);
  and g4543 (n4052, n_535, n_565);
  and g4544 (n4053, n_539, n_543);
  and g4545 (n4054, n3805, n3964);
  not g4546 (n_570, n4052);
  not g4547 (n_571, n4054);
  and g4548 (n4055, n_570, n_571);
  not g4549 (n_572, n4053);
  and g4550 (n4056, n_572, n4055);
  not g4551 (n_573, n4056);
  and g4552 (n4057, n_570, n_573);
  and g4553 (n4058, n3964, n4045);
  not g4554 (n_574, n4051);
  not g4555 (n_575, n4058);
  and g4556 (n4059, n_574, n_575);
  not g4557 (n_576, n4057);
  and g4558 (n4060, n_576, n4059);
  not g4559 (n_577, n4060);
  and g4560 (n4061, n_574, n_577);
  and g4561 (n4062, n_560, n_566);
  and g4562 (n4063, n3877, n4045);
  not g4563 (n_578, n4062);
  not g4564 (n_579, n4063);
  and g4565 (n4064, n_578, n_579);
  not g4566 (n_580, n4061);
  and g4567 (n4065, n_580, n4064);
  not g4568 (n_581, n4064);
  and g4569 (n4066, n4061, n_581);
  not g4570 (n_582, n4065);
  not g4571 (n_583, n4066);
  and g4572 (n4067, n_582, n_583);
  and g4573 (n4068, n4050, n4067);
  not g4576 (n_585, n4069);
  and g4577 (n4070, \a[26] , n_585);
  not g4578 (n_586, n4070);
  and g4579 (n4071, \a[26] , n_586);
  and g4580 (n4072, n_585, n_586);
  not g4581 (n_587, n4071);
  not g4582 (n_588, n4072);
  and g4583 (n4073, n_587, n_588);
  not g4584 (n_589, n4073);
  and g4585 (n4074, n3826, n_589);
  not g4586 (n_590, n4074);
  and g4587 (n4075, n3826, n_590);
  and g4588 (n4076, n_589, n_590);
  not g4589 (n_591, n4075);
  not g4590 (n_592, n4076);
  and g4591 (n4077, n_591, n_592);
  and g4592 (n4078, n3457, n_485);
  and g4593 (n4079, n_415, n3542);
  and g4594 (n4080, n_484, n3606);
  not g4600 (n_596, n3619);
  and g4601 (n4083, n3617, n_596);
  not g4602 (n_597, n4083);
  and g4603 (n4084, n_497, n_597);
  and g4604 (n4085, n3368, n4084);
  not g4607 (n_599, n4086);
  and g4608 (n4087, \a[29] , n_599);
  not g4609 (n_600, n4087);
  and g4610 (n4088, n_599, n_600);
  and g4611 (n4089, \a[29] , n_600);
  not g4612 (n_601, n4088);
  not g4613 (n_602, n4089);
  and g4614 (n4090, n_601, n_602);
  and g4615 (n4091, n_468, n_469);
  and g4616 (n4092, n3356, n_469);
  not g4617 (n_603, n4091);
  not g4618 (n_604, n4092);
  and g4619 (n4093, n_603, n_604);
  not g4620 (n_605, n4090);
  not g4621 (n_606, n4093);
  and g4622 (n4094, n_605, n_606);
  not g4623 (n_607, n4094);
  and g4624 (n4095, n_605, n_607);
  and g4625 (n4096, n_606, n_607);
  not g4626 (n_608, n4095);
  not g4627 (n_609, n4096);
  and g4628 (n4097, n_608, n_609);
  and g4629 (n4098, n_453, n_455);
  and g4630 (n4099, n_454, n3341);
  not g4631 (n_610, n4098);
  not g4632 (n_611, n4099);
  and g4633 (n4100, n_610, n_611);
  and g4634 (n4101, n_176, n_239);
  and g4664 (n4131, n_172, n1181);
  and g4665 (n4132, n_203, n4131);
  and g4685 (n4152, n279, n_259);
  and g4686 (n4153, n_234, n4152);
  not g4705 (n_612, n4121);
  not g4706 (n_613, n4171);
  and g4707 (n4172, n_612, n_613);
  and g4708 (n4173, n4121, n4171);
  not g4709 (n_614, n4172);
  not g4710 (n_615, n4173);
  and g4711 (n4174, n_614, n_615);
  not g4712 (n_617, \a[17] );
  and g4713 (n4175, n_617, n4174);
  not g4714 (n_618, n4175);
  and g4715 (n4176, n_614, n_618);
  not g4716 (n_619, n4176);
  and g4717 (n4177, n3146, n_619);
  not g4718 (n_620, n2918);
  and g4719 (n4178, n2916, n_620);
  not g4720 (n_621, n4178);
  and g4721 (n4179, n_406, n_621);
  and g4722 (n4180, n75, n4179);
  and g4723 (n4181, n_260, n3020);
  and g4724 (n4182, n_281, n3023);
  and g4725 (n4183, n_275, n3028);
  and g4733 (n4187, n_430, n4176);
  not g4734 (n_626, n4177);
  not g4735 (n_627, n4187);
  and g4736 (n4188, n_626, n_627);
  not g4737 (n_628, n4186);
  and g4738 (n4189, n_628, n4188);
  not g4739 (n_629, n4189);
  and g4740 (n4190, n_626, n_629);
  not g4741 (n_630, n4100);
  not g4742 (n_631, n4190);
  and g4743 (n4191, n_630, n_631);
  and g4744 (n4192, n4100, n4190);
  not g4745 (n_632, n4191);
  not g4746 (n_633, n4192);
  and g4747 (n4193, n_632, n_633);
  and g4748 (n4194, n_628, n_629);
  and g4749 (n4195, n4188, n_629);
  not g4750 (n_634, n4194);
  not g4751 (n_635, n4195);
  and g4752 (n4196, n_634, n_635);
  and g4753 (n4197, n_617, n_618);
  and g4754 (n4198, n_615, n4176);
  not g4755 (n_636, n4197);
  not g4756 (n_637, n4198);
  and g4757 (n4199, n_636, n_637);
  and g4758 (n4200, n_275, n3020);
  and g4759 (n4201, n_281, n3028);
  and g4760 (n4202, n_286, n3023);
  not g4761 (n_638, n2914);
  and g4762 (n4203, n2912, n_638);
  not g4763 (n_639, n4203);
  and g4764 (n4204, n_402, n_639);
  and g4765 (n4205, n75, n4204);
  not g4773 (n_644, n4199);
  not g4774 (n_645, n4208);
  and g4775 (n4209, n_644, n_645);
  and g4782 (n4216, n_175, n_181);
  and g4783 (n4217, n_93, n_292);
  and g4784 (n4218, n_276, n4217);
  and g4799 (n4233, n_208, n2468);
  and g4800 (n4234, n_279, n4233);
  not g4833 (n_646, n4266);
  and g4834 (n4267, n4121, n_646);
  and g4835 (n4268, n_612, n4266);
  and g4836 (n4269, n_79, n_51);
  and g4861 (n4294, n_142, n_165);
  and g4862 (n4295, n_144, n4294);
  and g4879 (n4312, n_46, n_192);
  and g4880 (n4313, n_114, n4312);
  and g4893 (n4326, n_133, n_188);
  and g4894 (n4327, n_247, n4326);
  and g4900 (n4333, n_67, n_211);
  and g4901 (n4334, n_143, n4333);
  and g4902 (n4335, n_91, n_264);
  and g4924 (n4357, n_257, n_297);
  and g4934 (n4367, n_36, n_121);
  not g4989 (n_647, n4351);
  not g4990 (n_648, n4421);
  and g4991 (n4422, n_647, n_648);
  and g4992 (n4423, n4351, n4421);
  not g4993 (n_649, n4422);
  not g4994 (n_650, n4423);
  and g4995 (n4424, n_649, n_650);
  not g4996 (n_652, \a[14] );
  and g4997 (n4425, n_652, n4424);
  not g4998 (n_653, n4425);
  and g4999 (n4426, n_649, n_653);
  not g5000 (n_654, n4426);
  and g5001 (n4427, n4266, n_654);
  not g5002 (n_655, n2906);
  and g5003 (n4428, n2904, n_655);
  not g5004 (n_656, n4428);
  and g5005 (n4429, n_394, n_656);
  and g5006 (n4430, n75, n4429);
  and g5007 (n4431, n_286, n3020);
  and g5008 (n4432, n_295, n3023);
  and g5009 (n4433, n_293, n3028);
  and g5017 (n4437, n_646, n4426);
  not g5018 (n_661, n4427);
  not g5019 (n_662, n4437);
  and g5020 (n4438, n_661, n_662);
  not g5021 (n_663, n4436);
  and g5022 (n4439, n_663, n4438);
  not g5023 (n_664, n4439);
  and g5024 (n4440, n_661, n_664);
  not g5025 (n_665, n4267);
  not g5026 (n_666, n4440);
  and g5027 (n4441, n_665, n_666);
  not g5028 (n_667, n4268);
  and g5029 (n4442, n_667, n4441);
  not g5030 (n_668, n4442);
  and g5031 (n4443, n_665, n_668);
  and g5032 (n4444, n4199, n4208);
  not g5033 (n_669, n4209);
  not g5034 (n_670, n4444);
  and g5035 (n4445, n_669, n_670);
  not g5036 (n_671, n4443);
  and g5037 (n4446, n_671, n4445);
  not g5038 (n_672, n4446);
  and g5039 (n4447, n_669, n_672);
  not g5040 (n_673, n4196);
  not g5041 (n_674, n4447);
  and g5042 (n4448, n_673, n_674);
  and g5043 (n4449, n4196, n4447);
  not g5044 (n_675, n4448);
  not g5045 (n_676, n4449);
  and g5046 (n4450, n_675, n_676);
  and g5047 (n4451, n_415, n3457);
  and g5048 (n4452, n_237, n3542);
  and g5049 (n4453, n_236, n3606);
  not g5050 (n_677, n4452);
  not g5051 (n_678, n4453);
  and g5052 (n4454, n_677, n_678);
  not g5053 (n_679, n4451);
  and g5054 (n4455, n_679, n4454);
  and g5055 (n4456, n_489, n4455);
  not g5056 (n_680, n3018);
  and g5057 (n4457, n_680, n4455);
  not g5058 (n_681, n4456);
  not g5059 (n_682, n4457);
  and g5060 (n4458, n_681, n_682);
  not g5061 (n_683, n4458);
  and g5062 (n4459, \a[29] , n_683);
  and g5063 (n4460, n_15, n4458);
  not g5064 (n_684, n4459);
  not g5065 (n_685, n4460);
  and g5066 (n4461, n_684, n_685);
  not g5067 (n_686, n4461);
  and g5068 (n4462, n4450, n_686);
  not g5069 (n_687, n4462);
  and g5070 (n4463, n_675, n_687);
  not g5071 (n_688, n4463);
  and g5072 (n4464, n4193, n_688);
  not g5073 (n_689, n4464);
  and g5074 (n4465, n_632, n_689);
  not g5075 (n_690, n4097);
  not g5076 (n_691, n4465);
  and g5077 (n4466, n_690, n_691);
  not g5078 (n_692, n4466);
  and g5079 (n4467, n_607, n_692);
  not g5080 (n_693, n3361);
  and g5081 (n4468, n_693, n3632);
  not g5082 (n_694, n4468);
  and g5083 (n4469, n_511, n_694);
  not g5084 (n_695, n4467);
  and g5085 (n4470, n_695, n4469);
  and g5086 (n4471, n3884, n_566);
  and g5087 (n4472, n_535, n3967);
  and g5088 (n4473, n_565, n4046);
  not g5094 (n_699, n4059);
  and g5095 (n4476, n4057, n_699);
  not g5096 (n_700, n4476);
  and g5097 (n4477, n_577, n_700);
  and g5098 (n4478, n4050, n4477);
  not g5101 (n_702, n4479);
  and g5102 (n4480, \a[26] , n_702);
  not g5103 (n_703, n4480);
  and g5104 (n4481, n_702, n_703);
  and g5105 (n4482, \a[26] , n_703);
  not g5106 (n_704, n4481);
  not g5107 (n_705, n4482);
  and g5108 (n4483, n_704, n_705);
  not g5109 (n_706, n4470);
  and g5110 (n4484, n_695, n_706);
  and g5111 (n4485, n4469, n_706);
  not g5112 (n_707, n4484);
  not g5113 (n_708, n4485);
  and g5114 (n4486, n_707, n_708);
  not g5115 (n_709, n4483);
  not g5116 (n_710, n4486);
  and g5117 (n4487, n_709, n_710);
  not g5118 (n_711, n4487);
  and g5119 (n4488, n_706, n_711);
  and g5146 (n4515, n3839, n4514);
  and g5147 (n4516, n_578, n_582);
  not g5148 (n_712, n4515);
  and g5149 (n4517, n_560, n_712);
  and g5150 (n4518, n3877, n4515);
  not g5151 (n_713, n4517);
  not g5152 (n_714, n4518);
  and g5153 (n4519, n_713, n_714);
  not g5154 (n_715, n4516);
  and g5155 (n4520, n_715, n4519);
  not g5156 (n_716, n4520);
  and g5157 (n4521, n3877, n_716);
  not g5158 (n_717, n4521);
  and g5159 (n4522, n_712, n_717);
  not g5160 (n_719, \a[21] );
  and g5161 (n4523, n_719, \a[22] );
  not g5162 (n_721, \a[22] );
  and g5163 (n4524, \a[21] , n_721);
  not g5164 (n_722, n4523);
  not g5165 (n_723, n4524);
  and g5166 (n4525, n_722, n_723);
  and g5167 (n4526, \a[20] , n_719);
  and g5168 (n4527, n_435, \a[21] );
  not g5169 (n_724, n4526);
  not g5170 (n_725, n4527);
  and g5171 (n4528, n_724, n_725);
  and g5172 (n4529, n_721, \a[23] );
  and g5173 (n4530, \a[22] , n_27);
  not g5174 (n_726, n4529);
  not g5175 (n_727, n4530);
  and g5176 (n4531, n_726, n_727);
  not g5177 (n_728, n4531);
  and g5178 (n4532, n4528, n_728);
  and g5179 (n4533, n4525, n4532);
  and g5180 (n4534, n_712, n4533);
  not g5181 (n_729, n4522);
  not g5182 (n_730, n4534);
  and g5183 (n4535, n_729, n_730);
  not g5184 (n_731, n4528);
  and g5185 (n4536, n_731, n_728);
  not g5186 (n_732, n4536);
  and g5187 (n4537, n_730, n_732);
  not g5188 (n_733, n4535);
  not g5189 (n_734, n4537);
  and g5190 (n4538, n_733, n_734);
  not g5191 (n_735, n4538);
  and g5192 (n4539, \a[23] , n_735);
  and g5193 (n4540, n_27, n4538);
  not g5194 (n_736, n4539);
  not g5195 (n_737, n4540);
  and g5196 (n4541, n_736, n_737);
  not g5197 (n_738, n4488);
  not g5198 (n_739, n4541);
  and g5199 (n4542, n_738, n_739);
  and g5200 (n4543, n4488, n4541);
  not g5201 (n_740, n4542);
  not g5202 (n_741, n4543);
  and g5203 (n4544, n_740, n_741);
  not g5204 (n_742, n4077);
  and g5205 (n4545, n_742, n4544);
  not g5206 (n_743, n4545);
  and g5207 (n4546, n_742, n_743);
  and g5208 (n4547, n4544, n_743);
  not g5209 (n_744, n4546);
  not g5210 (n_745, n4547);
  and g5211 (n4548, n_744, n_745);
  and g5212 (n4549, n4097, n4465);
  not g5213 (n_746, n4549);
  and g5214 (n4550, n_692, n_746);
  and g5215 (n4551, n3884, n_565);
  and g5216 (n4552, n_480, n3967);
  and g5217 (n4553, n_535, n4046);
  not g5218 (n_747, n4552);
  not g5219 (n_748, n4553);
  and g5220 (n4554, n_747, n_748);
  not g5221 (n_749, n4551);
  and g5222 (n4555, n_749, n4554);
  not g5223 (n_750, n4050);
  and g5224 (n4556, n_750, n4555);
  not g5225 (n_751, n4055);
  and g5226 (n4557, n4053, n_751);
  not g5227 (n_752, n4557);
  and g5228 (n4558, n_573, n_752);
  not g5229 (n_753, n4558);
  and g5230 (n4559, n4555, n_753);
  not g5231 (n_754, n4556);
  not g5232 (n_755, n4559);
  and g5233 (n4560, n_754, n_755);
  not g5234 (n_756, n4560);
  and g5235 (n4561, \a[26] , n_756);
  and g5236 (n4562, n_33, n4560);
  not g5237 (n_757, n4561);
  not g5238 (n_758, n4562);
  and g5239 (n4563, n_757, n_758);
  not g5240 (n_759, n4563);
  and g5241 (n4564, n4550, n_759);
  and g5242 (n4565, n_535, n3884);
  and g5243 (n4566, n_485, n3967);
  and g5244 (n4567, n_480, n4046);
  and g5250 (n4570, n3818, n4050);
  not g5253 (n_764, n4571);
  and g5254 (n4572, \a[26] , n_764);
  not g5255 (n_765, n4572);
  and g5256 (n4573, \a[26] , n_765);
  and g5257 (n4574, n_764, n_765);
  not g5258 (n_766, n4573);
  not g5259 (n_767, n4574);
  and g5260 (n4575, n_766, n_767);
  not g5261 (n_768, n4193);
  and g5262 (n4576, n_768, n4463);
  not g5263 (n_769, n4576);
  and g5264 (n4577, n_689, n_769);
  and g5265 (n4578, n3457, n_484);
  and g5266 (n4579, n_236, n3542);
  and g5267 (n4580, n_415, n3606);
  not g5268 (n_770, n4579);
  not g5269 (n_771, n4580);
  and g5270 (n4581, n_770, n_771);
  not g5271 (n_772, n4578);
  and g5272 (n4582, n_772, n4581);
  and g5273 (n4583, n_489, n4582);
  not g5274 (n_773, n3715);
  and g5275 (n4584, n_773, n4582);
  not g5276 (n_774, n4583);
  not g5277 (n_775, n4584);
  and g5278 (n4585, n_774, n_775);
  not g5279 (n_776, n4585);
  and g5280 (n4586, \a[29] , n_776);
  and g5281 (n4587, n_15, n4585);
  not g5282 (n_777, n4586);
  not g5283 (n_778, n4587);
  and g5284 (n4588, n_777, n_778);
  not g5285 (n_779, n4588);
  and g5286 (n4589, n4577, n_779);
  not g5287 (n_780, n4577);
  and g5288 (n4590, n_780, n4588);
  not g5289 (n_781, n4589);
  not g5290 (n_782, n4590);
  and g5291 (n4591, n_781, n_782);
  not g5292 (n_783, n4575);
  and g5293 (n4592, n_783, n4591);
  not g5294 (n_784, n4592);
  and g5295 (n4593, n_781, n_784);
  not g5296 (n_785, n4564);
  and g5297 (n4594, n4550, n_785);
  and g5298 (n4595, n_759, n_785);
  not g5299 (n_786, n4594);
  not g5300 (n_787, n4595);
  and g5301 (n4596, n_786, n_787);
  not g5302 (n_788, n4593);
  not g5303 (n_789, n4596);
  and g5304 (n4597, n_788, n_789);
  not g5305 (n_790, n4597);
  and g5306 (n4598, n_785, n_790);
  and g5307 (n4599, n4483, n_708);
  and g5308 (n4600, n_707, n4599);
  not g5309 (n_791, n4600);
  and g5310 (n4601, n_711, n_791);
  not g5311 (n_792, n4598);
  and g5312 (n4602, n_792, n4601);
  and g5313 (n4603, n_560, n4533);
  not g5314 (n_793, n4525);
  and g5315 (n4604, n_793, n4528);
  and g5316 (n4605, n_712, n4604);
  not g5317 (n_794, n4603);
  not g5318 (n_795, n4605);
  and g5319 (n4606, n_794, n_795);
  and g5320 (n4607, n_713, n_716);
  and g5321 (n4608, n4515, n4607);
  not g5322 (n_796, n4608);
  and g5323 (n4609, n_729, n_796);
  and g5324 (n4610, n4536, n4609);
  not g5325 (n_797, n4610);
  and g5326 (n4611, n4606, n_797);
  not g5327 (n_798, n4611);
  and g5328 (n4612, \a[23] , n_798);
  not g5329 (n_799, n4612);
  and g5330 (n4613, n_798, n_799);
  and g5331 (n4614, \a[23] , n_799);
  not g5332 (n_800, n4613);
  not g5333 (n_801, n4614);
  and g5334 (n4615, n_800, n_801);
  not g5335 (n_802, n4601);
  and g5336 (n4616, n4598, n_802);
  not g5337 (n_803, n4602);
  not g5338 (n_804, n4616);
  and g5339 (n4617, n_803, n_804);
  not g5340 (n_805, n4615);
  and g5341 (n4618, n_805, n4617);
  not g5342 (n_806, n4618);
  and g5343 (n4619, n_803, n_806);
  and g5344 (n4620, n4548, n4619);
  not g5345 (n_807, n4548);
  not g5346 (n_808, n4619);
  and g5347 (n4621, n_807, n_808);
  not g5348 (n_809, n4620);
  not g5349 (n_810, n4621);
  and g5350 (n4622, n_809, n_810);
  and g5351 (n4623, n4591, n_784);
  and g5352 (n4624, n_783, n_784);
  not g5353 (n_811, n4623);
  not g5354 (n_812, n4624);
  and g5355 (n4625, n_811, n_812);
  and g5356 (n4626, n_666, n_668);
  and g5357 (n4627, n_667, n4443);
  not g5358 (n_813, n4626);
  not g5359 (n_814, n4627);
  and g5360 (n4628, n_813, n_814);
  and g5361 (n4629, n_281, n3020);
  and g5362 (n4630, n_286, n3028);
  and g5363 (n4631, n_293, n3023);
  not g5364 (n_815, n2910);
  and g5365 (n4632, n2908, n_815);
  not g5366 (n_816, n4632);
  and g5367 (n4633, n_398, n_816);
  and g5368 (n4634, n75, n4633);
  not g5376 (n_821, n4628);
  not g5377 (n_822, n4637);
  and g5378 (n4638, n_821, n_822);
  and g5379 (n4639, n_237, n3457);
  and g5380 (n4640, n_275, n3542);
  and g5381 (n4641, n_260, n3606);
  and g5387 (n4644, n3331, n3368);
  not g5390 (n_827, n4645);
  and g5391 (n4646, \a[29] , n_827);
  not g5392 (n_828, n4646);
  and g5393 (n4647, n_827, n_828);
  and g5394 (n4648, \a[29] , n_828);
  not g5395 (n_829, n4647);
  not g5396 (n_830, n4648);
  and g5397 (n4649, n_829, n_830);
  not g5398 (n_831, n4638);
  and g5399 (n4650, n_821, n_831);
  and g5400 (n4651, n_822, n_831);
  not g5401 (n_832, n4650);
  not g5402 (n_833, n4651);
  and g5403 (n4652, n_832, n_833);
  not g5404 (n_834, n4649);
  not g5405 (n_835, n4652);
  and g5406 (n4653, n_834, n_835);
  not g5407 (n_836, n4653);
  and g5408 (n4654, n_831, n_836);
  not g5409 (n_837, n4445);
  and g5410 (n4655, n4443, n_837);
  not g5411 (n_838, n4655);
  and g5412 (n4656, n_672, n_838);
  not g5413 (n_839, n4654);
  and g5414 (n4657, n_839, n4656);
  and g5415 (n4658, n_236, n3457);
  and g5416 (n4659, n_260, n3542);
  and g5417 (n4660, n_237, n3606);
  and g5423 (n4663, n3347, n3368);
  not g5426 (n_844, n4664);
  and g5427 (n4665, \a[29] , n_844);
  not g5428 (n_845, n4665);
  and g5429 (n4666, \a[29] , n_845);
  and g5430 (n4667, n_844, n_845);
  not g5431 (n_846, n4666);
  not g5432 (n_847, n4667);
  and g5433 (n4668, n_846, n_847);
  not g5434 (n_848, n4656);
  and g5435 (n4669, n4654, n_848);
  not g5436 (n_849, n4657);
  not g5437 (n_850, n4669);
  and g5438 (n4670, n_849, n_850);
  not g5439 (n_851, n4668);
  and g5440 (n4671, n_851, n4670);
  not g5441 (n_852, n4671);
  and g5442 (n4672, n_849, n_852);
  not g5443 (n_853, n4450);
  and g5444 (n4673, n_853, n4461);
  not g5445 (n_854, n4673);
  and g5446 (n4674, n_687, n_854);
  not g5447 (n_855, n4672);
  and g5448 (n4675, n_855, n4674);
  not g5449 (n_856, n4674);
  and g5450 (n4676, n4672, n_856);
  not g5451 (n_857, n4675);
  not g5452 (n_858, n4676);
  and g5453 (n4677, n_857, n_858);
  and g5454 (n4678, n_480, n3884);
  and g5455 (n4679, n_484, n3967);
  and g5456 (n4680, n_485, n4046);
  and g5462 (n4683, n3627, n4050);
  not g5465 (n_863, n4684);
  and g5466 (n4685, \a[26] , n_863);
  not g5467 (n_864, n4685);
  and g5468 (n4686, \a[26] , n_864);
  and g5469 (n4687, n_863, n_864);
  not g5470 (n_865, n4686);
  not g5471 (n_866, n4687);
  and g5472 (n4688, n_865, n_866);
  not g5473 (n_867, n4688);
  and g5474 (n4689, n4677, n_867);
  not g5475 (n_868, n4689);
  and g5476 (n4690, n_857, n_868);
  not g5477 (n_869, n4625);
  not g5478 (n_870, n4690);
  and g5479 (n4691, n_869, n_870);
  and g5480 (n4692, n4625, n4690);
  not g5481 (n_871, n4691);
  not g5482 (n_872, n4692);
  and g5483 (n4693, n_871, n_872);
  and g5484 (n4694, n_731, n4531);
  and g5485 (n4695, n_560, n4694);
  and g5486 (n4696, n_565, n4533);
  and g5487 (n4697, n_566, n4604);
  and g5493 (n4700, n4067, n4536);
  not g5496 (n_877, n4701);
  and g5497 (n4702, \a[23] , n_877);
  not g5498 (n_878, n4702);
  and g5499 (n4703, \a[23] , n_878);
  and g5500 (n4704, n_877, n_878);
  not g5501 (n_879, n4703);
  not g5502 (n_880, n4704);
  and g5503 (n4705, n_879, n_880);
  not g5504 (n_881, n4705);
  and g5505 (n4706, n4693, n_881);
  not g5506 (n_882, n4706);
  and g5507 (n4707, n_871, n_882);
  and g5508 (n4708, n_712, n4694);
  and g5509 (n4709, n_566, n4533);
  and g5510 (n4710, n_560, n4604);
  not g5511 (n_883, n4709);
  not g5512 (n_884, n4710);
  and g5513 (n4711, n_883, n_884);
  not g5514 (n_885, n4708);
  and g5515 (n4712, n_885, n4711);
  and g5516 (n4713, n_732, n4712);
  not g5517 (n_886, n4519);
  and g5518 (n4714, n4516, n_886);
  not g5519 (n_887, n4714);
  and g5520 (n4715, n_716, n_887);
  not g5521 (n_888, n4715);
  and g5522 (n4716, n4712, n_888);
  not g5523 (n_889, n4713);
  not g5524 (n_890, n4716);
  and g5525 (n4717, n_889, n_890);
  not g5526 (n_891, n4717);
  and g5527 (n4718, \a[23] , n_891);
  and g5528 (n4719, n_27, n4717);
  not g5529 (n_892, n4718);
  not g5530 (n_893, n4719);
  and g5531 (n4720, n_892, n_893);
  not g5532 (n_894, n4707);
  not g5533 (n_895, n4720);
  and g5534 (n4721, n_894, n_895);
  and g5535 (n4722, n4707, n4720);
  not g5536 (n_896, n4721);
  not g5537 (n_897, n4722);
  and g5538 (n4723, n_896, n_897);
  and g5539 (n4724, n_788, n_790);
  and g5540 (n4725, n_789, n_790);
  not g5541 (n_898, n4724);
  not g5542 (n_899, n4725);
  and g5543 (n4726, n_898, n_899);
  not g5544 (n_900, n4726);
  and g5545 (n4727, n4723, n_900);
  not g5546 (n_901, n4727);
  and g5547 (n4728, n_896, n_901);
  not g5548 (n_902, n4617);
  and g5549 (n4729, n4615, n_902);
  not g5550 (n_903, n4729);
  and g5551 (n4730, n_806, n_903);
  not g5552 (n_904, n4728);
  and g5553 (n4731, n_904, n4730);
  and g5554 (n4732, n4723, n_901);
  and g5555 (n4733, n_900, n_901);
  not g5556 (n_905, n4732);
  not g5557 (n_906, n4733);
  and g5558 (n4734, n_905, n_906);
  and g5559 (n4735, n4677, n_868);
  and g5560 (n4736, n_867, n_868);
  not g5561 (n_907, n4735);
  not g5562 (n_908, n4736);
  and g5563 (n4737, n_907, n_908);
  and g5564 (n4738, n4670, n_852);
  and g5565 (n4739, n_851, n_852);
  not g5566 (n_909, n4738);
  not g5567 (n_910, n4739);
  and g5568 (n4740, n_909, n_910);
  and g5569 (n4741, n_485, n3884);
  and g5570 (n4742, n_415, n3967);
  and g5571 (n4743, n_484, n4046);
  not g5572 (n_911, n4742);
  not g5573 (n_912, n4743);
  and g5574 (n4744, n_911, n_912);
  not g5575 (n_913, n4741);
  and g5576 (n4745, n_913, n4744);
  and g5577 (n4746, n_750, n4745);
  not g5578 (n_914, n4084);
  and g5579 (n4747, n_914, n4745);
  not g5580 (n_915, n4746);
  not g5581 (n_916, n4747);
  and g5582 (n4748, n_915, n_916);
  not g5583 (n_917, n4748);
  and g5584 (n4749, \a[26] , n_917);
  and g5585 (n4750, n_33, n4748);
  not g5586 (n_918, n4749);
  not g5587 (n_919, n4750);
  and g5588 (n4751, n_918, n_919);
  not g5589 (n_920, n4740);
  not g5590 (n_921, n4751);
  and g5591 (n4752, n_920, n_921);
  and g5592 (n4753, n_834, n_836);
  and g5593 (n4754, n_835, n_836);
  not g5594 (n_922, n4753);
  not g5595 (n_923, n4754);
  and g5596 (n4755, n_922, n_923);
  and g5597 (n4756, n_663, n_664);
  and g5598 (n4757, n4438, n_664);
  not g5599 (n_924, n4756);
  not g5600 (n_925, n4757);
  and g5601 (n4758, n_924, n_925);
  and g5602 (n4759, n_652, n_653);
  and g5603 (n4760, n_650, n4426);
  not g5604 (n_926, n4759);
  not g5605 (n_927, n4760);
  and g5606 (n4761, n_926, n_927);
  and g5613 (n4768, n_228, n3490);
  and g5614 (n4769, n_277, n4768);
  and g5615 (n4770, n333, n1389);
  and g5616 (n4771, n_191, n4770);
  and g5631 (n4786, n_141, n_160);
  and g5632 (n4787, n_166, n_212);
  and g5633 (n4788, n_130, n4787);
  and g5643 (n4798, n1761, n4367);
  and g5644 (n4799, n_264, n4798);
  and g5673 (n4828, n_208, n_278);
  not g5690 (n_928, n4844);
  and g5691 (n4845, n4351, n_928);
  and g5692 (n4846, n_647, n4844);
  not g5693 (n_929, n2898);
  and g5694 (n4847, n2896, n_929);
  not g5695 (n_930, n4847);
  and g5696 (n4848, n_386, n_930);
  and g5697 (n4849, n75, n4848);
  and g5698 (n4850, n_295, n3020);
  and g5699 (n4851, n_299, n3023);
  and g5700 (n4852, n_298, n3028);
  not g5708 (n_935, n4845);
  not g5709 (n_936, n4855);
  and g5710 (n4856, n_935, n_936);
  not g5711 (n_937, n4846);
  and g5712 (n4857, n_937, n4856);
  not g5713 (n_938, n4857);
  and g5714 (n4858, n_935, n_938);
  not g5715 (n_939, n4761);
  not g5716 (n_940, n4858);
  and g5717 (n4859, n_939, n_940);
  not g5718 (n_941, n2902);
  and g5719 (n4860, n2900, n_941);
  not g5720 (n_942, n4860);
  and g5721 (n4861, n_390, n_942);
  and g5722 (n4862, n75, n4861);
  and g5723 (n4863, n_293, n3020);
  and g5724 (n4864, n_298, n3023);
  and g5725 (n4865, n_295, n3028);
  and g5733 (n4869, n4761, n4858);
  not g5734 (n_947, n4859);
  not g5735 (n_948, n4869);
  and g5736 (n4870, n_947, n_948);
  not g5737 (n_949, n4868);
  and g5738 (n4871, n_949, n4870);
  not g5739 (n_950, n4871);
  and g5740 (n4872, n_947, n_950);
  not g5741 (n_951, n4758);
  not g5742 (n_952, n4872);
  and g5743 (n4873, n_951, n_952);
  and g5744 (n4874, n4758, n4872);
  not g5745 (n_953, n4873);
  not g5746 (n_954, n4874);
  and g5747 (n4875, n_953, n_954);
  and g5748 (n4876, n_260, n3457);
  and g5749 (n4877, n_281, n3542);
  and g5750 (n4878, n_275, n3606);
  not g5751 (n_955, n4877);
  not g5752 (n_956, n4878);
  and g5753 (n4879, n_955, n_956);
  not g5754 (n_957, n4876);
  and g5755 (n4880, n_957, n4879);
  and g5756 (n4881, n_489, n4880);
  not g5757 (n_958, n4179);
  and g5758 (n4882, n_958, n4880);
  not g5759 (n_959, n4881);
  not g5760 (n_960, n4882);
  and g5761 (n4883, n_959, n_960);
  not g5762 (n_961, n4883);
  and g5763 (n4884, \a[29] , n_961);
  and g5764 (n4885, n_15, n4883);
  not g5765 (n_962, n4884);
  not g5766 (n_963, n4885);
  and g5767 (n4886, n_962, n_963);
  not g5768 (n_964, n4886);
  and g5769 (n4887, n4875, n_964);
  not g5770 (n_965, n4887);
  and g5771 (n4888, n_953, n_965);
  not g5772 (n_966, n4755);
  not g5773 (n_967, n4888);
  and g5774 (n4889, n_966, n_967);
  and g5775 (n4890, n4755, n4888);
  not g5776 (n_968, n4889);
  not g5777 (n_969, n4890);
  and g5778 (n4891, n_968, n_969);
  and g5779 (n4892, n_484, n3884);
  and g5780 (n4893, n_236, n3967);
  and g5781 (n4894, n_415, n4046);
  and g5787 (n4897, n3715, n4050);
  not g5790 (n_974, n4898);
  and g5791 (n4899, \a[26] , n_974);
  not g5792 (n_975, n4899);
  and g5793 (n4900, \a[26] , n_975);
  and g5794 (n4901, n_974, n_975);
  not g5795 (n_976, n4900);
  not g5796 (n_977, n4901);
  and g5797 (n4902, n_976, n_977);
  not g5798 (n_978, n4902);
  and g5799 (n4903, n4891, n_978);
  not g5800 (n_979, n4903);
  and g5801 (n4904, n_968, n_979);
  and g5802 (n4905, n4740, n4751);
  not g5803 (n_980, n4752);
  not g5804 (n_981, n4905);
  and g5805 (n4906, n_980, n_981);
  not g5806 (n_982, n4904);
  and g5807 (n4907, n_982, n4906);
  not g5808 (n_983, n4907);
  and g5809 (n4908, n_980, n_983);
  not g5810 (n_984, n4737);
  not g5811 (n_985, n4908);
  and g5812 (n4909, n_984, n_985);
  and g5813 (n4910, n4737, n4908);
  not g5814 (n_986, n4909);
  not g5815 (n_987, n4910);
  and g5816 (n4911, n_986, n_987);
  and g5817 (n4912, n_566, n4694);
  and g5818 (n4913, n_535, n4533);
  and g5819 (n4914, n_565, n4604);
  and g5825 (n4917, n4477, n4536);
  not g5828 (n_992, n4918);
  and g5829 (n4919, \a[23] , n_992);
  not g5830 (n_993, n4919);
  and g5831 (n4920, \a[23] , n_993);
  and g5832 (n4921, n_992, n_993);
  not g5833 (n_994, n4920);
  not g5834 (n_995, n4921);
  and g5835 (n4922, n_994, n_995);
  not g5836 (n_996, n4922);
  and g5837 (n4923, n4911, n_996);
  not g5838 (n_997, n4923);
  and g5839 (n4924, n_986, n_997);
  not g5840 (n_999, \a[18] );
  and g5841 (n4925, n_999, \a[19] );
  not g5842 (n_1001, \a[19] );
  and g5843 (n4926, \a[18] , n_1001);
  not g5844 (n_1002, n4925);
  not g5845 (n_1003, n4926);
  and g5846 (n4927, n_1002, n_1003);
  and g5847 (n4928, \a[19] , n_435);
  and g5848 (n4929, n_1001, \a[20] );
  not g5849 (n_1004, n4928);
  not g5850 (n_1005, n4929);
  and g5851 (n4930, n_1004, n_1005);
  and g5852 (n4931, \a[17] , n_999);
  and g5853 (n4932, n_617, \a[18] );
  not g5854 (n_1006, n4931);
  not g5855 (n_1007, n4932);
  and g5856 (n4933, n_1006, n_1007);
  not g5857 (n_1008, n4930);
  and g5858 (n4934, n_1008, n4933);
  and g5859 (n4935, n4927, n4934);
  and g5860 (n4936, n_712, n4935);
  not g5861 (n_1009, n4936);
  and g5862 (n4937, n_729, n_1009);
  not g5863 (n_1010, n4933);
  and g5864 (n4938, n_1008, n_1010);
  not g5865 (n_1011, n4938);
  and g5866 (n4939, n_1009, n_1011);
  not g5867 (n_1012, n4937);
  not g5868 (n_1013, n4939);
  and g5869 (n4940, n_1012, n_1013);
  not g5870 (n_1014, n4940);
  and g5871 (n4941, \a[20] , n_1014);
  and g5872 (n4942, n_435, n4940);
  not g5873 (n_1015, n4941);
  not g5874 (n_1016, n4942);
  and g5875 (n4943, n_1015, n_1016);
  not g5876 (n_1017, n4924);
  not g5877 (n_1018, n4943);
  and g5878 (n4944, n_1017, n_1018);
  and g5879 (n4945, n4693, n_882);
  and g5880 (n4946, n_881, n_882);
  not g5881 (n_1019, n4945);
  not g5882 (n_1020, n4946);
  and g5883 (n4947, n_1019, n_1020);
  and g5884 (n4948, n4924, n4943);
  not g5885 (n_1021, n4944);
  not g5886 (n_1022, n4948);
  and g5887 (n4949, n_1021, n_1022);
  not g5888 (n_1023, n4947);
  and g5889 (n4950, n_1023, n4949);
  not g5890 (n_1024, n4950);
  and g5891 (n4951, n_1021, n_1024);
  not g5892 (n_1025, n4734);
  not g5893 (n_1026, n4951);
  and g5894 (n4952, n_1025, n_1026);
  and g5895 (n4953, n4734, n4951);
  not g5896 (n_1027, n4952);
  not g5897 (n_1028, n4953);
  and g5898 (n4954, n_1027, n_1028);
  and g5899 (n4955, n_1023, n_1024);
  and g5900 (n4956, n4949, n_1024);
  not g5901 (n_1029, n4955);
  not g5902 (n_1030, n4956);
  and g5903 (n4957, n_1029, n_1030);
  and g5904 (n4958, n4911, n_997);
  and g5905 (n4959, n_996, n_997);
  not g5906 (n_1031, n4958);
  not g5907 (n_1032, n4959);
  and g5908 (n4960, n_1031, n_1032);
  and g5909 (n4961, n_565, n4694);
  and g5910 (n4962, n_480, n4533);
  and g5911 (n4963, n_535, n4604);
  and g5917 (n4966, n4536, n4558);
  not g5920 (n_1037, n4967);
  and g5921 (n4968, \a[23] , n_1037);
  not g5922 (n_1038, n4968);
  and g5923 (n4969, n_1037, n_1038);
  and g5924 (n4970, \a[23] , n_1038);
  not g5925 (n_1039, n4969);
  not g5926 (n_1040, n4970);
  and g5927 (n4971, n_1039, n_1040);
  not g5928 (n_1041, n4906);
  and g5929 (n4972, n4904, n_1041);
  not g5930 (n_1042, n4972);
  and g5931 (n4973, n_983, n_1042);
  not g5932 (n_1043, n4971);
  and g5933 (n4974, n_1043, n4973);
  not g5934 (n_1044, n4974);
  and g5935 (n4975, n_1043, n_1044);
  and g5936 (n4976, n4973, n_1044);
  not g5937 (n_1045, n4975);
  not g5938 (n_1046, n4976);
  and g5939 (n4977, n_1045, n_1046);
  and g5940 (n4978, n4891, n_979);
  and g5941 (n4979, n_978, n_979);
  not g5942 (n_1047, n4978);
  not g5943 (n_1048, n4979);
  and g5944 (n4980, n_1047, n_1048);
  and g5945 (n4981, n_275, n3457);
  and g5946 (n4982, n_286, n3542);
  and g5947 (n4983, n_281, n3606);
  and g5953 (n4986, n3368, n4204);
  not g5956 (n_1053, n4987);
  and g5957 (n4988, \a[29] , n_1053);
  not g5958 (n_1054, n4988);
  and g5959 (n4989, n_1053, n_1054);
  and g5960 (n4990, \a[29] , n_1054);
  not g5961 (n_1055, n4989);
  not g5962 (n_1056, n4990);
  and g5963 (n4991, n_1055, n_1056);
  and g5964 (n4992, n_949, n_950);
  and g5965 (n4993, n4870, n_950);
  not g5966 (n_1057, n4992);
  not g5967 (n_1058, n4993);
  and g5968 (n4994, n_1057, n_1058);
  not g5969 (n_1059, n4991);
  not g5970 (n_1060, n4994);
  and g5971 (n4995, n_1059, n_1060);
  not g5972 (n_1061, n4995);
  and g5973 (n4996, n_1059, n_1061);
  and g5974 (n4997, n_1060, n_1061);
  not g5975 (n_1062, n4996);
  not g5976 (n_1063, n4997);
  and g5977 (n4998, n_1062, n_1063);
  and g5978 (n4999, n_936, n_938);
  and g5979 (n5000, n_937, n4858);
  not g5980 (n_1064, n4999);
  not g5981 (n_1065, n5000);
  and g5982 (n5001, n_1064, n_1065);
  and g5983 (n5002, n_234, n_288);
  and g6001 (n5020, n_54, n_270);
  and g6002 (n5021, n_214, n5020);
  and g6016 (n5035, n_130, n_216);
  and g6017 (n5036, n_103, n5035);
  and g6018 (n5037, n_142, n_170);
  and g6019 (n5038, n_114, n5037);
  and g6020 (n5039, n979, n2406);
  and g6021 (n5040, n_287, n5039);
  and g6045 (n5064, n_86, n_261);
  and g6046 (n5065, n_112, n_272);
  and g6047 (n5066, n_172, n5065);
  not g6088 (n_1066, n5053);
  not g6089 (n_1067, n5106);
  and g6090 (n5107, n_1066, n_1067);
  and g6091 (n5108, n5053, n5106);
  not g6092 (n_1068, n5107);
  not g6093 (n_1069, n5108);
  and g6094 (n5109, n_1068, n_1069);
  not g6095 (n_1071, \a[11] );
  and g6096 (n5110, n_1071, n5109);
  not g6097 (n_1072, n5110);
  and g6098 (n5111, n_1068, n_1072);
  not g6099 (n_1073, n5111);
  and g6100 (n5112, n4351, n_1073);
  not g6101 (n_1074, n2894);
  and g6102 (n5113, n2892, n_1074);
  not g6103 (n_1075, n5113);
  and g6104 (n5114, n_382, n_1075);
  and g6105 (n5115, n75, n5114);
  and g6106 (n5116, n_298, n3020);
  and g6107 (n5117, n_300, n3023);
  and g6108 (n5118, n_299, n3028);
  and g6116 (n5122, n_647, n5111);
  not g6117 (n_1080, n5112);
  not g6118 (n_1081, n5122);
  and g6119 (n5123, n_1080, n_1081);
  not g6120 (n_1082, n5121);
  and g6121 (n5124, n_1082, n5123);
  not g6122 (n_1083, n5124);
  and g6123 (n5125, n_1080, n_1083);
  not g6124 (n_1084, n5001);
  not g6125 (n_1085, n5125);
  and g6126 (n5126, n_1084, n_1085);
  and g6127 (n5127, n5001, n5125);
  not g6128 (n_1086, n5126);
  not g6129 (n_1087, n5127);
  and g6130 (n5128, n_1086, n_1087);
  and g6131 (n5129, n_1082, n_1083);
  and g6132 (n5130, n5123, n_1083);
  not g6133 (n_1088, n5129);
  not g6134 (n_1089, n5130);
  and g6135 (n5131, n_1088, n_1089);
  and g6136 (n5132, n_1071, n_1072);
  and g6137 (n5133, n_1069, n5111);
  not g6138 (n_1090, n5132);
  not g6139 (n_1091, n5133);
  and g6140 (n5134, n_1090, n_1091);
  and g6141 (n5135, n_299, n3020);
  and g6142 (n5136, n_300, n3028);
  and g6143 (n5137, n_301, n3023);
  not g6144 (n_1092, n2890);
  and g6145 (n5138, n2888, n_1092);
  not g6146 (n_1093, n5138);
  and g6147 (n5139, n_378, n_1093);
  and g6148 (n5140, n75, n5139);
  not g6156 (n_1098, n5134);
  not g6157 (n_1099, n5143);
  and g6158 (n5144, n_1098, n_1099);
  and g6163 (n5149, n_183, n1523);
  and g6164 (n5150, n_137, n5149);
  and g6165 (n5151, n_60, n1330);
  and g6166 (n5152, n_104, n5151);
  not g6183 (n_1100, n5168);
  and g6184 (n5169, n5053, n_1100);
  and g6185 (n5170, n_1066, n5168);
  and g6186 (n5171, n_273, n_291);
  and g6187 (n5172, n_148, n1128);
  and g6188 (n5173, n_117, n5172);
  and g6204 (n5189, n_59, n_196);
  and g6205 (n5190, n_116, n5189);
  and g6215 (n5200, n_56, n_193);
  and g6216 (n5201, n_191, n5200);
  and g6285 (n5270, n202, n_216);
  and g6286 (n5271, n_183, n5270);
  not g6336 (n_1101, n5254);
  not g6337 (n_1102, n5320);
  and g6338 (n5321, n_1101, n_1102);
  and g6339 (n5322, n5254, n5320);
  not g6340 (n_1103, n5321);
  not g6341 (n_1104, n5322);
  and g6342 (n5323, n_1103, n_1104);
  not g6343 (n_1106, \a[8] );
  and g6344 (n5324, n_1106, n5323);
  not g6345 (n_1107, n5324);
  and g6346 (n5325, n_1103, n_1107);
  not g6347 (n_1108, n5325);
  and g6348 (n5326, n5053, n_1108);
  not g6349 (n_1109, n2882);
  and g6350 (n5327, n2880, n_1109);
  not g6351 (n_1110, n5327);
  and g6352 (n5328, n_370, n_1110);
  and g6353 (n5329, n75, n5328);
  and g6354 (n5330, n_301, n3020);
  and g6355 (n5331, n_303, n3023);
  and g6356 (n5332, n_302, n3028);
  and g6364 (n5336, n_1066, n5325);
  not g6365 (n_1115, n5326);
  not g6366 (n_1116, n5336);
  and g6367 (n5337, n_1115, n_1116);
  not g6368 (n_1117, n5335);
  and g6369 (n5338, n_1117, n5337);
  not g6370 (n_1118, n5338);
  and g6371 (n5339, n_1115, n_1118);
  not g6372 (n_1119, n5169);
  not g6373 (n_1120, n5339);
  and g6374 (n5340, n_1119, n_1120);
  not g6375 (n_1121, n5170);
  and g6376 (n5341, n_1121, n5340);
  not g6377 (n_1122, n5341);
  and g6378 (n5342, n_1119, n_1122);
  and g6379 (n5343, n5134, n5143);
  not g6380 (n_1123, n5144);
  not g6381 (n_1124, n5343);
  and g6382 (n5344, n_1123, n_1124);
  not g6383 (n_1125, n5342);
  and g6384 (n5345, n_1125, n5344);
  not g6385 (n_1126, n5345);
  and g6386 (n5346, n_1123, n_1126);
  not g6387 (n_1127, n5131);
  not g6388 (n_1128, n5346);
  and g6389 (n5347, n_1127, n_1128);
  and g6390 (n5348, n5131, n5346);
  not g6391 (n_1129, n5347);
  not g6392 (n_1130, n5348);
  and g6393 (n5349, n_1129, n_1130);
  and g6394 (n5350, n_286, n3457);
  and g6395 (n5351, n_295, n3542);
  and g6396 (n5352, n_293, n3606);
  not g6397 (n_1131, n5351);
  not g6398 (n_1132, n5352);
  and g6399 (n5353, n_1131, n_1132);
  not g6400 (n_1133, n5350);
  and g6401 (n5354, n_1133, n5353);
  and g6402 (n5355, n_489, n5354);
  not g6403 (n_1134, n4429);
  and g6404 (n5356, n_1134, n5354);
  not g6405 (n_1135, n5355);
  not g6406 (n_1136, n5356);
  and g6407 (n5357, n_1135, n_1136);
  not g6408 (n_1137, n5357);
  and g6409 (n5358, \a[29] , n_1137);
  and g6410 (n5359, n_15, n5357);
  not g6411 (n_1138, n5358);
  not g6412 (n_1139, n5359);
  and g6413 (n5360, n_1138, n_1139);
  not g6414 (n_1140, n5360);
  and g6415 (n5361, n5349, n_1140);
  not g6416 (n_1141, n5361);
  and g6417 (n5362, n_1129, n_1141);
  not g6418 (n_1142, n5362);
  and g6419 (n5363, n5128, n_1142);
  not g6420 (n_1143, n5363);
  and g6421 (n5364, n_1086, n_1143);
  not g6422 (n_1144, n4998);
  not g6423 (n_1145, n5364);
  and g6424 (n5365, n_1144, n_1145);
  not g6425 (n_1146, n5365);
  and g6426 (n5366, n_1061, n_1146);
  not g6427 (n_1147, n4875);
  and g6428 (n5367, n_1147, n4886);
  not g6429 (n_1148, n5367);
  and g6430 (n5368, n_965, n_1148);
  not g6431 (n_1149, n5366);
  and g6432 (n5369, n_1149, n5368);
  not g6433 (n_1150, n5368);
  and g6434 (n5370, n5366, n_1150);
  not g6435 (n_1151, n5369);
  not g6436 (n_1152, n5370);
  and g6437 (n5371, n_1151, n_1152);
  and g6438 (n5372, n_415, n3884);
  and g6439 (n5373, n_237, n3967);
  and g6440 (n5374, n_236, n4046);
  and g6446 (n5377, n3018, n4050);
  not g6449 (n_1157, n5378);
  and g6450 (n5379, \a[26] , n_1157);
  not g6451 (n_1158, n5379);
  and g6452 (n5380, \a[26] , n_1158);
  and g6453 (n5381, n_1157, n_1158);
  not g6454 (n_1159, n5380);
  not g6455 (n_1160, n5381);
  and g6456 (n5382, n_1159, n_1160);
  not g6457 (n_1161, n5382);
  and g6458 (n5383, n5371, n_1161);
  not g6459 (n_1162, n5383);
  and g6460 (n5384, n_1151, n_1162);
  not g6461 (n_1163, n4980);
  not g6462 (n_1164, n5384);
  and g6463 (n5385, n_1163, n_1164);
  and g6464 (n5386, n4980, n5384);
  not g6465 (n_1165, n5385);
  not g6466 (n_1166, n5386);
  and g6467 (n5387, n_1165, n_1166);
  and g6468 (n5388, n_535, n4694);
  and g6469 (n5389, n_485, n4533);
  and g6470 (n5390, n_480, n4604);
  and g6476 (n5393, n3818, n4536);
  not g6479 (n_1171, n5394);
  and g6480 (n5395, \a[23] , n_1171);
  not g6481 (n_1172, n5395);
  and g6482 (n5396, \a[23] , n_1172);
  and g6483 (n5397, n_1171, n_1172);
  not g6484 (n_1173, n5396);
  not g6485 (n_1174, n5397);
  and g6486 (n5398, n_1173, n_1174);
  not g6487 (n_1175, n5398);
  and g6488 (n5399, n5387, n_1175);
  not g6489 (n_1176, n5399);
  and g6490 (n5400, n_1165, n_1176);
  not g6491 (n_1177, n4977);
  not g6492 (n_1178, n5400);
  and g6493 (n5401, n_1177, n_1178);
  not g6494 (n_1179, n5401);
  and g6495 (n5402, n_1044, n_1179);
  not g6496 (n_1180, n4960);
  not g6497 (n_1181, n5402);
  and g6498 (n5403, n_1180, n_1181);
  and g6499 (n5404, n4960, n5402);
  not g6500 (n_1182, n5403);
  not g6501 (n_1183, n5404);
  and g6502 (n5405, n_1182, n_1183);
  and g6503 (n5406, n_560, n4935);
  not g6504 (n_1184, n4927);
  and g6505 (n5407, n_1184, n4933);
  and g6506 (n5408, n_712, n5407);
  not g6507 (n_1185, n5406);
  not g6508 (n_1186, n5408);
  and g6509 (n5409, n_1185, n_1186);
  and g6510 (n5410, n4609, n4938);
  not g6511 (n_1187, n5410);
  and g6512 (n5411, n5409, n_1187);
  not g6513 (n_1188, n5411);
  and g6514 (n5412, \a[20] , n_1188);
  not g6515 (n_1189, n5412);
  and g6516 (n5413, \a[20] , n_1189);
  and g6517 (n5414, n_1188, n_1189);
  not g6518 (n_1190, n5413);
  not g6519 (n_1191, n5414);
  and g6520 (n5415, n_1190, n_1191);
  not g6521 (n_1192, n5415);
  and g6522 (n5416, n5405, n_1192);
  not g6523 (n_1193, n5416);
  and g6524 (n5417, n_1182, n_1193);
  not g6525 (n_1194, n4957);
  not g6526 (n_1195, n5417);
  and g6527 (n5418, n_1194, n_1195);
  and g6528 (n5419, n4957, n5417);
  not g6529 (n_1196, n5418);
  not g6530 (n_1197, n5419);
  and g6531 (n5420, n_1196, n_1197);
  and g6532 (n5421, n5405, n_1193);
  and g6533 (n5422, n_1192, n_1193);
  not g6534 (n_1198, n5421);
  not g6535 (n_1199, n5422);
  and g6536 (n5423, n_1198, n_1199);
  and g6537 (n5424, n5387, n_1176);
  and g6538 (n5425, n_1175, n_1176);
  not g6539 (n_1200, n5424);
  not g6540 (n_1201, n5425);
  and g6541 (n5426, n_1200, n_1201);
  and g6542 (n5427, n5371, n_1162);
  and g6543 (n5428, n_1161, n_1162);
  not g6544 (n_1202, n5427);
  not g6545 (n_1203, n5428);
  and g6546 (n5429, n_1202, n_1203);
  and g6547 (n5430, n4998, n5364);
  not g6548 (n_1204, n5430);
  and g6549 (n5431, n_1146, n_1204);
  and g6550 (n5432, n_236, n3884);
  and g6551 (n5433, n_260, n3967);
  and g6552 (n5434, n_237, n4046);
  not g6553 (n_1205, n5433);
  not g6554 (n_1206, n5434);
  and g6555 (n5435, n_1205, n_1206);
  not g6556 (n_1207, n5432);
  and g6557 (n5436, n_1207, n5435);
  and g6558 (n5437, n_750, n5436);
  not g6559 (n_1208, n3347);
  and g6560 (n5438, n_1208, n5436);
  not g6561 (n_1209, n5437);
  not g6562 (n_1210, n5438);
  and g6563 (n5439, n_1209, n_1210);
  not g6564 (n_1211, n5439);
  and g6565 (n5440, \a[26] , n_1211);
  and g6566 (n5441, n_33, n5439);
  not g6567 (n_1212, n5440);
  not g6568 (n_1213, n5441);
  and g6569 (n5442, n_1212, n_1213);
  not g6570 (n_1214, n5442);
  and g6571 (n5443, n5431, n_1214);
  and g6572 (n5444, n_237, n3884);
  and g6573 (n5445, n_275, n3967);
  and g6574 (n5446, n_260, n4046);
  and g6580 (n5449, n3331, n4050);
  not g6583 (n_1219, n5450);
  and g6584 (n5451, \a[26] , n_1219);
  not g6585 (n_1220, n5451);
  and g6586 (n5452, \a[26] , n_1220);
  and g6587 (n5453, n_1219, n_1220);
  not g6588 (n_1221, n5452);
  not g6589 (n_1222, n5453);
  and g6590 (n5454, n_1221, n_1222);
  not g6591 (n_1223, n5128);
  and g6592 (n5455, n_1223, n5362);
  not g6593 (n_1224, n5455);
  and g6594 (n5456, n_1143, n_1224);
  and g6595 (n5457, n_281, n3457);
  and g6596 (n5458, n_293, n3542);
  and g6597 (n5459, n_286, n3606);
  not g6598 (n_1225, n5458);
  not g6599 (n_1226, n5459);
  and g6600 (n5460, n_1225, n_1226);
  not g6601 (n_1227, n5457);
  and g6602 (n5461, n_1227, n5460);
  and g6603 (n5462, n_489, n5461);
  not g6604 (n_1228, n4633);
  and g6605 (n5463, n_1228, n5461);
  not g6606 (n_1229, n5462);
  not g6607 (n_1230, n5463);
  and g6608 (n5464, n_1229, n_1230);
  not g6609 (n_1231, n5464);
  and g6610 (n5465, \a[29] , n_1231);
  and g6611 (n5466, n_15, n5464);
  not g6612 (n_1232, n5465);
  not g6613 (n_1233, n5466);
  and g6614 (n5467, n_1232, n_1233);
  not g6615 (n_1234, n5467);
  and g6616 (n5468, n5456, n_1234);
  not g6617 (n_1235, n5456);
  and g6618 (n5469, n_1235, n5467);
  not g6619 (n_1236, n5468);
  not g6620 (n_1237, n5469);
  and g6621 (n5470, n_1236, n_1237);
  not g6622 (n_1238, n5454);
  and g6623 (n5471, n_1238, n5470);
  not g6624 (n_1239, n5471);
  and g6625 (n5472, n_1236, n_1239);
  not g6626 (n_1240, n5431);
  and g6627 (n5473, n_1240, n5442);
  not g6628 (n_1241, n5443);
  not g6629 (n_1242, n5473);
  and g6630 (n5474, n_1241, n_1242);
  not g6631 (n_1243, n5472);
  and g6632 (n5475, n_1243, n5474);
  not g6633 (n_1244, n5475);
  and g6634 (n5476, n_1241, n_1244);
  not g6635 (n_1245, n5429);
  not g6636 (n_1246, n5476);
  and g6637 (n5477, n_1245, n_1246);
  and g6638 (n5478, n5429, n5476);
  not g6639 (n_1247, n5477);
  not g6640 (n_1248, n5478);
  and g6641 (n5479, n_1247, n_1248);
  and g6642 (n5480, n_480, n4694);
  and g6643 (n5481, n_484, n4533);
  and g6644 (n5482, n_485, n4604);
  and g6650 (n5485, n3627, n4536);
  not g6653 (n_1253, n5486);
  and g6654 (n5487, \a[23] , n_1253);
  not g6655 (n_1254, n5487);
  and g6656 (n5488, \a[23] , n_1254);
  and g6657 (n5489, n_1253, n_1254);
  not g6658 (n_1255, n5488);
  not g6659 (n_1256, n5489);
  and g6660 (n5490, n_1255, n_1256);
  not g6661 (n_1257, n5490);
  and g6662 (n5491, n5479, n_1257);
  not g6663 (n_1258, n5491);
  and g6664 (n5492, n_1247, n_1258);
  not g6665 (n_1259, n5426);
  not g6666 (n_1260, n5492);
  and g6667 (n5493, n_1259, n_1260);
  and g6668 (n5494, n5426, n5492);
  not g6669 (n_1261, n5493);
  not g6670 (n_1262, n5494);
  and g6671 (n5495, n_1261, n_1262);
  and g6672 (n5496, n4930, n_1010);
  and g6673 (n5497, n_560, n5496);
  and g6674 (n5498, n_565, n4935);
  and g6675 (n5499, n_566, n5407);
  and g6681 (n5502, n4067, n4938);
  not g6684 (n_1267, n5503);
  and g6685 (n5504, \a[20] , n_1267);
  not g6686 (n_1268, n5504);
  and g6687 (n5505, \a[20] , n_1268);
  and g6688 (n5506, n_1267, n_1268);
  not g6689 (n_1269, n5505);
  not g6690 (n_1270, n5506);
  and g6691 (n5507, n_1269, n_1270);
  not g6692 (n_1271, n5507);
  and g6693 (n5508, n5495, n_1271);
  not g6694 (n_1272, n5508);
  and g6695 (n5509, n_1261, n_1272);
  and g6696 (n5510, n_712, n5496);
  and g6697 (n5511, n_566, n4935);
  and g6698 (n5512, n_560, n5407);
  not g6699 (n_1273, n5511);
  not g6700 (n_1274, n5512);
  and g6701 (n5513, n_1273, n_1274);
  not g6702 (n_1275, n5510);
  and g6703 (n5514, n_1275, n5513);
  and g6704 (n5515, n_1011, n5514);
  and g6705 (n5516, n_888, n5514);
  not g6706 (n_1276, n5515);
  not g6707 (n_1277, n5516);
  and g6708 (n5517, n_1276, n_1277);
  not g6709 (n_1278, n5517);
  and g6710 (n5518, \a[20] , n_1278);
  and g6711 (n5519, n_435, n5517);
  not g6712 (n_1279, n5518);
  not g6713 (n_1280, n5519);
  and g6714 (n5520, n_1279, n_1280);
  not g6715 (n_1281, n5509);
  not g6716 (n_1282, n5520);
  and g6717 (n5521, n_1281, n_1282);
  and g6718 (n5522, n4977, n5400);
  not g6719 (n_1283, n5522);
  and g6720 (n5523, n_1179, n_1283);
  and g6721 (n5524, n5509, n5520);
  not g6722 (n_1284, n5521);
  not g6723 (n_1285, n5524);
  and g6724 (n5525, n_1284, n_1285);
  and g6725 (n5526, n5523, n5525);
  not g6726 (n_1286, n5526);
  and g6727 (n5527, n_1284, n_1286);
  not g6728 (n_1287, n5423);
  not g6729 (n_1288, n5527);
  and g6730 (n5528, n_1287, n_1288);
  and g6731 (n5529, n5423, n5527);
  not g6732 (n_1289, n5528);
  not g6733 (n_1290, n5529);
  and g6734 (n5530, n_1289, n_1290);
  and g6735 (n5531, n5479, n_1258);
  and g6736 (n5532, n_1257, n_1258);
  not g6737 (n_1291, n5531);
  not g6738 (n_1292, n5532);
  and g6739 (n5533, n_1291, n_1292);
  and g6740 (n5534, n_485, n4694);
  and g6741 (n5535, n_415, n4533);
  and g6742 (n5536, n_484, n4604);
  and g6748 (n5539, n4084, n4536);
  not g6751 (n_1297, n5540);
  and g6752 (n5541, \a[23] , n_1297);
  not g6753 (n_1298, n5541);
  and g6754 (n5542, n_1297, n_1298);
  and g6755 (n5543, \a[23] , n_1298);
  not g6756 (n_1299, n5542);
  not g6757 (n_1300, n5543);
  and g6758 (n5544, n_1299, n_1300);
  not g6759 (n_1301, n5474);
  and g6760 (n5545, n5472, n_1301);
  not g6761 (n_1302, n5545);
  and g6762 (n5546, n_1244, n_1302);
  not g6763 (n_1303, n5544);
  and g6764 (n5547, n_1303, n5546);
  not g6765 (n_1304, n5547);
  and g6766 (n5548, n_1303, n_1304);
  and g6767 (n5549, n5546, n_1304);
  not g6768 (n_1305, n5548);
  not g6769 (n_1306, n5549);
  and g6770 (n5550, n_1305, n_1306);
  and g6771 (n5551, n5470, n_1239);
  and g6772 (n5552, n_1238, n_1239);
  not g6773 (n_1307, n5551);
  not g6774 (n_1308, n5552);
  and g6775 (n5553, n_1307, n_1308);
  and g6776 (n5554, n_1120, n_1122);
  and g6777 (n5555, n_1121, n5342);
  not g6778 (n_1309, n5554);
  not g6779 (n_1310, n5555);
  and g6780 (n5556, n_1309, n_1310);
  and g6781 (n5557, n_300, n3020);
  and g6782 (n5558, n_301, n3028);
  and g6783 (n5559, n_302, n3023);
  not g6784 (n_1311, n2886);
  and g6785 (n5560, n2884, n_1311);
  not g6786 (n_1312, n5560);
  and g6787 (n5561, n_374, n_1312);
  and g6788 (n5562, n75, n5561);
  not g6796 (n_1317, n5556);
  not g6797 (n_1318, n5565);
  and g6798 (n5566, n_1317, n_1318);
  and g6799 (n5567, n_295, n3457);
  and g6800 (n5568, n_299, n3542);
  and g6801 (n5569, n_298, n3606);
  and g6807 (n5572, n3368, n4848);
  not g6810 (n_1323, n5573);
  and g6811 (n5574, \a[29] , n_1323);
  not g6812 (n_1324, n5574);
  and g6813 (n5575, n_1323, n_1324);
  and g6814 (n5576, \a[29] , n_1324);
  not g6815 (n_1325, n5575);
  not g6816 (n_1326, n5576);
  and g6817 (n5577, n_1325, n_1326);
  not g6818 (n_1327, n5566);
  and g6819 (n5578, n_1317, n_1327);
  and g6820 (n5579, n_1318, n_1327);
  not g6821 (n_1328, n5578);
  not g6822 (n_1329, n5579);
  and g6823 (n5580, n_1328, n_1329);
  not g6824 (n_1330, n5577);
  not g6825 (n_1331, n5580);
  and g6826 (n5581, n_1330, n_1331);
  not g6827 (n_1332, n5581);
  and g6828 (n5582, n_1327, n_1332);
  not g6829 (n_1333, n5344);
  and g6830 (n5583, n5342, n_1333);
  not g6831 (n_1334, n5583);
  and g6832 (n5584, n_1126, n_1334);
  not g6833 (n_1335, n5582);
  and g6834 (n5585, n_1335, n5584);
  and g6835 (n5586, n_293, n3457);
  and g6836 (n5587, n_298, n3542);
  and g6837 (n5588, n_295, n3606);
  and g6843 (n5591, n3368, n4861);
  not g6846 (n_1340, n5592);
  and g6847 (n5593, \a[29] , n_1340);
  not g6848 (n_1341, n5593);
  and g6849 (n5594, \a[29] , n_1341);
  and g6850 (n5595, n_1340, n_1341);
  not g6851 (n_1342, n5594);
  not g6852 (n_1343, n5595);
  and g6853 (n5596, n_1342, n_1343);
  not g6854 (n_1344, n5584);
  and g6855 (n5597, n5582, n_1344);
  not g6856 (n_1345, n5585);
  not g6857 (n_1346, n5597);
  and g6858 (n5598, n_1345, n_1346);
  not g6859 (n_1347, n5596);
  and g6860 (n5599, n_1347, n5598);
  not g6861 (n_1348, n5599);
  and g6862 (n5600, n_1345, n_1348);
  not g6863 (n_1349, n5349);
  and g6864 (n5601, n_1349, n5360);
  not g6865 (n_1350, n5601);
  and g6866 (n5602, n_1141, n_1350);
  not g6867 (n_1351, n5600);
  and g6868 (n5603, n_1351, n5602);
  not g6869 (n_1352, n5602);
  and g6870 (n5604, n5600, n_1352);
  not g6871 (n_1353, n5603);
  not g6872 (n_1354, n5604);
  and g6873 (n5605, n_1353, n_1354);
  and g6874 (n5606, n_260, n3884);
  and g6875 (n5607, n_281, n3967);
  and g6876 (n5608, n_275, n4046);
  and g6882 (n5611, n4050, n4179);
  not g6885 (n_1359, n5612);
  and g6886 (n5613, \a[26] , n_1359);
  not g6887 (n_1360, n5613);
  and g6888 (n5614, \a[26] , n_1360);
  and g6889 (n5615, n_1359, n_1360);
  not g6890 (n_1361, n5614);
  not g6891 (n_1362, n5615);
  and g6892 (n5616, n_1361, n_1362);
  not g6893 (n_1363, n5616);
  and g6894 (n5617, n5605, n_1363);
  not g6895 (n_1364, n5617);
  and g6896 (n5618, n_1353, n_1364);
  not g6897 (n_1365, n5553);
  not g6898 (n_1366, n5618);
  and g6899 (n5619, n_1365, n_1366);
  and g6900 (n5620, n5553, n5618);
  not g6901 (n_1367, n5619);
  not g6902 (n_1368, n5620);
  and g6903 (n5621, n_1367, n_1368);
  and g6904 (n5622, n_484, n4694);
  and g6905 (n5623, n_236, n4533);
  and g6906 (n5624, n_415, n4604);
  and g6912 (n5627, n3715, n4536);
  not g6915 (n_1373, n5628);
  and g6916 (n5629, \a[23] , n_1373);
  not g6917 (n_1374, n5629);
  and g6918 (n5630, \a[23] , n_1374);
  and g6919 (n5631, n_1373, n_1374);
  not g6920 (n_1375, n5630);
  not g6921 (n_1376, n5631);
  and g6922 (n5632, n_1375, n_1376);
  not g6923 (n_1377, n5632);
  and g6924 (n5633, n5621, n_1377);
  not g6925 (n_1378, n5633);
  and g6926 (n5634, n_1367, n_1378);
  not g6927 (n_1379, n5550);
  not g6928 (n_1380, n5634);
  and g6929 (n5635, n_1379, n_1380);
  not g6930 (n_1381, n5635);
  and g6931 (n5636, n_1304, n_1381);
  not g6932 (n_1382, n5533);
  not g6933 (n_1383, n5636);
  and g6934 (n5637, n_1382, n_1383);
  and g6935 (n5638, n5533, n5636);
  not g6936 (n_1384, n5637);
  not g6937 (n_1385, n5638);
  and g6938 (n5639, n_1384, n_1385);
  and g6939 (n5640, n_566, n5496);
  and g6940 (n5641, n_535, n4935);
  and g6941 (n5642, n_565, n5407);
  and g6947 (n5645, n4477, n4938);
  not g6950 (n_1390, n5646);
  and g6951 (n5647, \a[20] , n_1390);
  not g6952 (n_1391, n5647);
  and g6953 (n5648, \a[20] , n_1391);
  and g6954 (n5649, n_1390, n_1391);
  not g6955 (n_1392, n5648);
  not g6956 (n_1393, n5649);
  and g6957 (n5650, n_1392, n_1393);
  not g6958 (n_1394, n5650);
  and g6959 (n5651, n5639, n_1394);
  not g6960 (n_1395, n5651);
  and g6961 (n5652, n_1384, n_1395);
  not g6962 (n_1397, \a[15] );
  and g6963 (n5653, n_1397, \a[16] );
  not g6964 (n_1399, \a[16] );
  and g6965 (n5654, \a[15] , n_1399);
  not g6966 (n_1400, n5653);
  not g6967 (n_1401, n5654);
  and g6968 (n5655, n_1400, n_1401);
  and g6969 (n5656, \a[14] , n_1397);
  and g6970 (n5657, n_652, \a[15] );
  not g6971 (n_1402, n5656);
  not g6972 (n_1403, n5657);
  and g6973 (n5658, n_1402, n_1403);
  and g6974 (n5659, \a[16] , n_617);
  and g6975 (n5660, n_1399, \a[17] );
  not g6976 (n_1404, n5659);
  not g6977 (n_1405, n5660);
  and g6978 (n5661, n_1404, n_1405);
  not g6979 (n_1406, n5661);
  and g6980 (n5662, n5658, n_1406);
  and g6981 (n5663, n5655, n5662);
  and g6982 (n5664, n_712, n5663);
  not g6983 (n_1407, n5664);
  and g6984 (n5665, n_729, n_1407);
  not g6985 (n_1408, n5658);
  and g6986 (n5666, n_1408, n_1406);
  not g6987 (n_1409, n5666);
  and g6988 (n5667, n_1407, n_1409);
  not g6989 (n_1410, n5665);
  not g6990 (n_1411, n5667);
  and g6991 (n5668, n_1410, n_1411);
  not g6992 (n_1412, n5668);
  and g6993 (n5669, \a[17] , n_1412);
  and g6994 (n5670, n_617, n5668);
  not g6995 (n_1413, n5669);
  not g6996 (n_1414, n5670);
  and g6997 (n5671, n_1413, n_1414);
  not g6998 (n_1415, n5652);
  not g6999 (n_1416, n5671);
  and g7000 (n5672, n_1415, n_1416);
  and g7001 (n5673, n5495, n_1272);
  and g7002 (n5674, n_1271, n_1272);
  not g7003 (n_1417, n5673);
  not g7004 (n_1418, n5674);
  and g7005 (n5675, n_1417, n_1418);
  and g7006 (n5676, n5652, n5671);
  not g7007 (n_1419, n5672);
  not g7008 (n_1420, n5676);
  and g7009 (n5677, n_1419, n_1420);
  not g7010 (n_1421, n5675);
  and g7011 (n5678, n_1421, n5677);
  not g7012 (n_1422, n5678);
  and g7013 (n5679, n_1419, n_1422);
  not g7014 (n_1423, n5523);
  not g7015 (n_1424, n5525);
  and g7016 (n5680, n_1423, n_1424);
  not g7017 (n_1425, n5680);
  and g7018 (n5681, n_1286, n_1425);
  not g7019 (n_1426, n5679);
  and g7020 (n5682, n_1426, n5681);
  and g7021 (n5683, n_1421, n_1422);
  and g7022 (n5684, n5677, n_1422);
  not g7023 (n_1427, n5683);
  not g7024 (n_1428, n5684);
  and g7025 (n5685, n_1427, n_1428);
  and g7026 (n5686, n5639, n_1395);
  and g7027 (n5687, n_1394, n_1395);
  not g7028 (n_1429, n5686);
  not g7029 (n_1430, n5687);
  and g7030 (n5688, n_1429, n_1430);
  and g7031 (n5689, n5550, n5634);
  not g7032 (n_1431, n5689);
  and g7033 (n5690, n_1381, n_1431);
  and g7034 (n5691, n_565, n5496);
  and g7035 (n5692, n_480, n4935);
  and g7036 (n5693, n_535, n5407);
  not g7037 (n_1432, n5692);
  not g7038 (n_1433, n5693);
  and g7039 (n5694, n_1432, n_1433);
  not g7040 (n_1434, n5691);
  and g7041 (n5695, n_1434, n5694);
  and g7042 (n5696, n_1011, n5695);
  and g7043 (n5697, n_753, n5695);
  not g7044 (n_1435, n5696);
  not g7045 (n_1436, n5697);
  and g7046 (n5698, n_1435, n_1436);
  not g7047 (n_1437, n5698);
  and g7048 (n5699, \a[20] , n_1437);
  and g7049 (n5700, n_435, n5698);
  not g7050 (n_1438, n5699);
  not g7051 (n_1439, n5700);
  and g7052 (n5701, n_1438, n_1439);
  not g7053 (n_1440, n5701);
  and g7054 (n5702, n5690, n_1440);
  and g7055 (n5703, n5621, n_1378);
  and g7056 (n5704, n_1377, n_1378);
  not g7057 (n_1441, n5703);
  not g7058 (n_1442, n5704);
  and g7059 (n5705, n_1441, n_1442);
  and g7060 (n5706, n5605, n_1364);
  and g7061 (n5707, n_1363, n_1364);
  not g7062 (n_1443, n5706);
  not g7063 (n_1444, n5707);
  and g7064 (n5708, n_1443, n_1444);
  and g7065 (n5709, n5598, n_1348);
  and g7066 (n5710, n_1347, n_1348);
  not g7067 (n_1445, n5709);
  not g7068 (n_1446, n5710);
  and g7069 (n5711, n_1445, n_1446);
  and g7070 (n5712, n_275, n3884);
  and g7071 (n5713, n_286, n3967);
  and g7072 (n5714, n_281, n4046);
  not g7073 (n_1447, n5713);
  not g7074 (n_1448, n5714);
  and g7075 (n5715, n_1447, n_1448);
  not g7076 (n_1449, n5712);
  and g7077 (n5716, n_1449, n5715);
  and g7078 (n5717, n_750, n5716);
  not g7079 (n_1450, n4204);
  and g7080 (n5718, n_1450, n5716);
  not g7081 (n_1451, n5717);
  not g7082 (n_1452, n5718);
  and g7083 (n5719, n_1451, n_1452);
  not g7084 (n_1453, n5719);
  and g7085 (n5720, \a[26] , n_1453);
  and g7086 (n5721, n_33, n5719);
  not g7087 (n_1454, n5720);
  not g7088 (n_1455, n5721);
  and g7089 (n5722, n_1454, n_1455);
  not g7090 (n_1456, n5711);
  not g7091 (n_1457, n5722);
  and g7092 (n5723, n_1456, n_1457);
  and g7093 (n5724, n_1330, n_1332);
  and g7094 (n5725, n_1331, n_1332);
  not g7095 (n_1458, n5724);
  not g7096 (n_1459, n5725);
  and g7097 (n5726, n_1458, n_1459);
  and g7098 (n5727, n_1117, n_1118);
  and g7099 (n5728, n5337, n_1118);
  not g7100 (n_1460, n5727);
  not g7101 (n_1461, n5728);
  and g7102 (n5729, n_1460, n_1461);
  and g7103 (n5730, n_1106, n_1107);
  and g7104 (n5731, n_1104, n5325);
  not g7105 (n_1462, n5730);
  not g7106 (n_1463, n5731);
  and g7107 (n5732, n_1462, n_1463);
  and g7108 (n5733, n533, n591);
  and g7109 (n5734, n_123, n5733);
  and g7122 (n5747, n_118, n_159);
  and g7123 (n5748, n_117, n5747);
  not g7141 (n_1464, n5765);
  and g7142 (n5766, n5254, n_1464);
  and g7143 (n5767, n_1101, n5765);
  and g7150 (n5774, n_159, n_181);
  and g7151 (n5775, n_43, n5774);
  and g7152 (n5776, n_113, n_148);
  and g7153 (n5777, n_74, n5776);
  and g7162 (n5786, n_194, n_280);
  and g7163 (n5787, n_158, n5786);
  and g7168 (n5792, n_78, n_241);
  and g7169 (n5793, n_70, n5792);
  and g7183 (n5807, n_146, n_191);
  and g7184 (n5808, n_109, n5807);
  not g7202 (n_1465, n5825);
  and g7203 (n5826, n_10, n_1465);
  and g7204 (n5827, \a[2] , n_1465);
  and g7205 (n5828, n_10, n5825);
  not g7206 (n_1466, n5827);
  not g7207 (n_1467, n5828);
  and g7208 (n5829, n_1466, n_1467);
  not g7209 (n_1468, n5829);
  and g7210 (n5830, n_3, n_1468);
  not g7211 (n_1469, n5826);
  not g7212 (n_1470, n5830);
  and g7213 (n5831, n_1469, n_1470);
  not g7214 (n_1471, n5831);
  and g7215 (n5832, n5254, n_1471);
  not g7216 (n_1472, n2870);
  and g7217 (n5833, n2868, n_1472);
  not g7218 (n_1473, n5833);
  and g7219 (n5834, n_358, n_1473);
  and g7220 (n5835, n75, n5834);
  and g7221 (n5836, n_304, n3020);
  and g7222 (n5837, n_306, n3023);
  and g7223 (n5838, n_305, n3028);
  and g7231 (n5842, n_1101, n5831);
  not g7232 (n_1478, n5832);
  not g7233 (n_1479, n5842);
  and g7234 (n5843, n_1478, n_1479);
  not g7235 (n_1480, n5841);
  and g7236 (n5844, n_1480, n5843);
  not g7237 (n_1481, n5844);
  and g7238 (n5845, n_1478, n_1481);
  not g7239 (n_1482, n5766);
  not g7240 (n_1483, n5845);
  and g7241 (n5846, n_1482, n_1483);
  not g7242 (n_1484, n5767);
  and g7243 (n5847, n_1484, n5846);
  not g7244 (n_1485, n5847);
  and g7245 (n5848, n_1482, n_1485);
  not g7246 (n_1486, n5732);
  not g7247 (n_1487, n5848);
  and g7248 (n5849, n_1486, n_1487);
  not g7249 (n_1488, n2878);
  and g7250 (n5850, n2876, n_1488);
  not g7251 (n_1489, n5850);
  and g7252 (n5851, n_366, n_1489);
  and g7253 (n5852, n75, n5851);
  and g7254 (n5853, n_302, n3020);
  and g7255 (n5854, n_304, n3023);
  and g7256 (n5855, n_303, n3028);
  and g7264 (n5859, n5732, n5848);
  not g7265 (n_1494, n5849);
  not g7266 (n_1495, n5859);
  and g7267 (n5860, n_1494, n_1495);
  not g7268 (n_1496, n5858);
  and g7269 (n5861, n_1496, n5860);
  not g7270 (n_1497, n5861);
  and g7271 (n5862, n_1494, n_1497);
  not g7272 (n_1498, n5729);
  not g7273 (n_1499, n5862);
  and g7274 (n5863, n_1498, n_1499);
  and g7275 (n5864, n5729, n5862);
  not g7276 (n_1500, n5863);
  not g7277 (n_1501, n5864);
  and g7278 (n5865, n_1500, n_1501);
  and g7279 (n5866, n_298, n3457);
  and g7280 (n5867, n_300, n3542);
  and g7281 (n5868, n_299, n3606);
  not g7282 (n_1502, n5867);
  not g7283 (n_1503, n5868);
  and g7284 (n5869, n_1502, n_1503);
  not g7285 (n_1504, n5866);
  and g7286 (n5870, n_1504, n5869);
  and g7287 (n5871, n_489, n5870);
  not g7288 (n_1505, n5114);
  and g7289 (n5872, n_1505, n5870);
  not g7290 (n_1506, n5871);
  not g7291 (n_1507, n5872);
  and g7292 (n5873, n_1506, n_1507);
  not g7293 (n_1508, n5873);
  and g7294 (n5874, \a[29] , n_1508);
  and g7295 (n5875, n_15, n5873);
  not g7296 (n_1509, n5874);
  not g7297 (n_1510, n5875);
  and g7298 (n5876, n_1509, n_1510);
  not g7299 (n_1511, n5876);
  and g7300 (n5877, n5865, n_1511);
  not g7301 (n_1512, n5877);
  and g7302 (n5878, n_1500, n_1512);
  not g7303 (n_1513, n5726);
  not g7304 (n_1514, n5878);
  and g7305 (n5879, n_1513, n_1514);
  and g7306 (n5880, n5726, n5878);
  not g7307 (n_1515, n5879);
  not g7308 (n_1516, n5880);
  and g7309 (n5881, n_1515, n_1516);
  and g7310 (n5882, n_281, n3884);
  and g7311 (n5883, n_293, n3967);
  and g7312 (n5884, n_286, n4046);
  and g7318 (n5887, n4050, n4633);
  not g7321 (n_1521, n5888);
  and g7322 (n5889, \a[26] , n_1521);
  not g7323 (n_1522, n5889);
  and g7324 (n5890, \a[26] , n_1522);
  and g7325 (n5891, n_1521, n_1522);
  not g7326 (n_1523, n5890);
  not g7327 (n_1524, n5891);
  and g7328 (n5892, n_1523, n_1524);
  not g7329 (n_1525, n5892);
  and g7330 (n5893, n5881, n_1525);
  not g7331 (n_1526, n5893);
  and g7332 (n5894, n_1515, n_1526);
  and g7333 (n5895, n5711, n5722);
  not g7334 (n_1527, n5723);
  not g7335 (n_1528, n5895);
  and g7336 (n5896, n_1527, n_1528);
  not g7337 (n_1529, n5894);
  and g7338 (n5897, n_1529, n5896);
  not g7339 (n_1530, n5897);
  and g7340 (n5898, n_1527, n_1530);
  not g7341 (n_1531, n5708);
  not g7342 (n_1532, n5898);
  and g7343 (n5899, n_1531, n_1532);
  and g7344 (n5900, n5708, n5898);
  not g7345 (n_1533, n5899);
  not g7346 (n_1534, n5900);
  and g7347 (n5901, n_1533, n_1534);
  and g7348 (n5902, n_415, n4694);
  and g7349 (n5903, n_237, n4533);
  and g7350 (n5904, n_236, n4604);
  and g7356 (n5907, n3018, n4536);
  not g7359 (n_1539, n5908);
  and g7360 (n5909, \a[23] , n_1539);
  not g7361 (n_1540, n5909);
  and g7362 (n5910, \a[23] , n_1540);
  and g7363 (n5911, n_1539, n_1540);
  not g7364 (n_1541, n5910);
  not g7365 (n_1542, n5911);
  and g7366 (n5912, n_1541, n_1542);
  not g7367 (n_1543, n5912);
  and g7368 (n5913, n5901, n_1543);
  not g7369 (n_1544, n5913);
  and g7370 (n5914, n_1533, n_1544);
  not g7371 (n_1545, n5705);
  not g7372 (n_1546, n5914);
  and g7373 (n5915, n_1545, n_1546);
  and g7374 (n5916, n5705, n5914);
  not g7375 (n_1547, n5915);
  not g7376 (n_1548, n5916);
  and g7377 (n5917, n_1547, n_1548);
  and g7378 (n5918, n_535, n5496);
  and g7379 (n5919, n_485, n4935);
  and g7380 (n5920, n_480, n5407);
  and g7386 (n5923, n3818, n4938);
  not g7389 (n_1553, n5924);
  and g7390 (n5925, \a[20] , n_1553);
  not g7391 (n_1554, n5925);
  and g7392 (n5926, \a[20] , n_1554);
  and g7393 (n5927, n_1553, n_1554);
  not g7394 (n_1555, n5926);
  not g7395 (n_1556, n5927);
  and g7396 (n5928, n_1555, n_1556);
  not g7397 (n_1557, n5928);
  and g7398 (n5929, n5917, n_1557);
  not g7399 (n_1558, n5929);
  and g7400 (n5930, n_1547, n_1558);
  not g7401 (n_1559, n5690);
  and g7402 (n5931, n_1559, n5701);
  not g7403 (n_1560, n5702);
  not g7404 (n_1561, n5931);
  and g7405 (n5932, n_1560, n_1561);
  not g7406 (n_1562, n5930);
  and g7407 (n5933, n_1562, n5932);
  not g7408 (n_1563, n5933);
  and g7409 (n5934, n_1560, n_1563);
  not g7410 (n_1564, n5688);
  not g7411 (n_1565, n5934);
  and g7412 (n5935, n_1564, n_1565);
  and g7413 (n5936, n5688, n5934);
  not g7414 (n_1566, n5935);
  not g7415 (n_1567, n5936);
  and g7416 (n5937, n_1566, n_1567);
  and g7417 (n5938, n_560, n5663);
  not g7418 (n_1568, n5655);
  and g7419 (n5939, n_1568, n5658);
  and g7420 (n5940, n_712, n5939);
  not g7421 (n_1569, n5938);
  not g7422 (n_1570, n5940);
  and g7423 (n5941, n_1569, n_1570);
  and g7424 (n5942, n4609, n5666);
  not g7425 (n_1571, n5942);
  and g7426 (n5943, n5941, n_1571);
  not g7427 (n_1572, n5943);
  and g7428 (n5944, \a[17] , n_1572);
  not g7429 (n_1573, n5944);
  and g7430 (n5945, \a[17] , n_1573);
  and g7431 (n5946, n_1572, n_1573);
  not g7432 (n_1574, n5945);
  not g7433 (n_1575, n5946);
  and g7434 (n5947, n_1574, n_1575);
  not g7435 (n_1576, n5947);
  and g7436 (n5948, n5937, n_1576);
  not g7437 (n_1577, n5948);
  and g7438 (n5949, n_1566, n_1577);
  not g7439 (n_1578, n5685);
  not g7440 (n_1579, n5949);
  and g7441 (n5950, n_1578, n_1579);
  and g7442 (n5951, n5685, n5949);
  not g7443 (n_1580, n5950);
  not g7444 (n_1581, n5951);
  and g7445 (n5952, n_1580, n_1581);
  and g7446 (n5953, n5937, n_1577);
  and g7447 (n5954, n_1576, n_1577);
  not g7448 (n_1582, n5953);
  not g7449 (n_1583, n5954);
  and g7450 (n5955, n_1582, n_1583);
  and g7451 (n5956, n5917, n_1558);
  and g7452 (n5957, n_1557, n_1558);
  not g7453 (n_1584, n5956);
  not g7454 (n_1585, n5957);
  and g7455 (n5958, n_1584, n_1585);
  and g7456 (n5959, n5901, n_1544);
  and g7457 (n5960, n_1543, n_1544);
  not g7458 (n_1586, n5959);
  not g7459 (n_1587, n5960);
  and g7460 (n5961, n_1586, n_1587);
  and g7461 (n5962, n_236, n4694);
  and g7462 (n5963, n_260, n4533);
  and g7463 (n5964, n_237, n4604);
  and g7469 (n5967, n3347, n4536);
  not g7472 (n_1592, n5968);
  and g7473 (n5969, \a[23] , n_1592);
  not g7474 (n_1593, n5969);
  and g7475 (n5970, n_1592, n_1593);
  and g7476 (n5971, \a[23] , n_1593);
  not g7477 (n_1594, n5970);
  not g7478 (n_1595, n5971);
  and g7479 (n5972, n_1594, n_1595);
  not g7480 (n_1596, n5896);
  and g7481 (n5973, n5894, n_1596);
  not g7482 (n_1597, n5973);
  and g7483 (n5974, n_1530, n_1597);
  not g7484 (n_1598, n5972);
  and g7485 (n5975, n_1598, n5974);
  not g7486 (n_1599, n5975);
  and g7487 (n5976, n_1598, n_1599);
  and g7488 (n5977, n5974, n_1599);
  not g7489 (n_1600, n5976);
  not g7490 (n_1601, n5977);
  and g7491 (n5978, n_1600, n_1601);
  and g7492 (n5979, n5881, n_1526);
  and g7493 (n5980, n_1525, n_1526);
  not g7494 (n_1602, n5979);
  not g7495 (n_1603, n5980);
  and g7496 (n5981, n_1602, n_1603);
  and g7497 (n5982, n_299, n3457);
  and g7498 (n5983, n_301, n3542);
  and g7499 (n5984, n_300, n3606);
  and g7505 (n5987, n3368, n5139);
  not g7508 (n_1608, n5988);
  and g7509 (n5989, \a[29] , n_1608);
  not g7510 (n_1609, n5989);
  and g7511 (n5990, n_1608, n_1609);
  and g7512 (n5991, \a[29] , n_1609);
  not g7513 (n_1610, n5990);
  not g7514 (n_1611, n5991);
  and g7515 (n5992, n_1610, n_1611);
  and g7516 (n5993, n_1496, n_1497);
  and g7517 (n5994, n5860, n_1497);
  not g7518 (n_1612, n5993);
  not g7519 (n_1613, n5994);
  and g7520 (n5995, n_1612, n_1613);
  not g7521 (n_1614, n5992);
  not g7522 (n_1615, n5995);
  and g7523 (n5996, n_1614, n_1615);
  not g7524 (n_1616, n5996);
  and g7525 (n5997, n_1614, n_1616);
  and g7526 (n5998, n_1615, n_1616);
  not g7527 (n_1617, n5997);
  not g7528 (n_1618, n5998);
  and g7529 (n5999, n_1617, n_1618);
  and g7530 (n6000, n_1483, n_1485);
  and g7531 (n6001, n_1484, n5848);
  not g7532 (n_1619, n6000);
  not g7533 (n_1620, n6001);
  and g7534 (n6002, n_1619, n_1620);
  and g7535 (n6003, n_303, n3020);
  and g7536 (n6004, n_304, n3028);
  and g7537 (n6005, n_305, n3023);
  not g7538 (n_1621, n2874);
  and g7539 (n6006, n2872, n_1621);
  not g7540 (n_1622, n6006);
  and g7541 (n6007, n_362, n_1622);
  and g7542 (n6008, n75, n6007);
  not g7550 (n_1627, n6002);
  not g7551 (n_1628, n6011);
  and g7552 (n6012, n_1627, n_1628);
  and g7553 (n6013, n_1480, n_1481);
  and g7554 (n6014, n5843, n_1481);
  not g7555 (n_1629, n6013);
  not g7556 (n_1630, n6014);
  and g7557 (n6015, n_1629, n_1630);
  not g7584 (n_1631, n6041);
  and g7585 (n6042, \a[2] , n_1631);
  and g7586 (n6043, n_10, n6041);
  and g7598 (n6055, n690, n3252);
  and g7599 (n6056, n618, n6055);
  not g7618 (n_1632, n6074);
  and g7619 (n6075, \a[2] , n_1632);
  and g7620 (n6076, n_10, n6074);
  and g7628 (n6084, n_122, n_176);
  and g7647 (n6103, n_38, n4367);
  and g7648 (n6104, n_240, n6103);
  not g7663 (n_1633, n6118);
  and g7664 (n6119, \a[2] , n_1633);
  and g7665 (n6120, n_10, n6118);
  not g7666 (n_1634, n2854);
  and g7667 (n6121, n2852, n_1634);
  not g7668 (n_1635, n6121);
  and g7669 (n6122, n_342, n_1635);
  and g7670 (n6123, n75, n6122);
  and g7671 (n6124, n_308, n3020);
  and g7672 (n6125, n_310, n3023);
  and g7673 (n6126, n_309, n3028);
  not g7681 (n_1640, n6119);
  not g7682 (n_1641, n6129);
  and g7683 (n6130, n_1640, n_1641);
  not g7684 (n_1642, n6120);
  and g7685 (n6131, n_1642, n6130);
  not g7686 (n_1643, n6131);
  and g7687 (n6132, n_1640, n_1643);
  not g7688 (n_1644, n6075);
  not g7689 (n_1645, n6132);
  and g7690 (n6133, n_1644, n_1645);
  not g7691 (n_1646, n6076);
  and g7692 (n6134, n_1646, n6133);
  not g7693 (n_1647, n6134);
  and g7694 (n6135, n_1644, n_1647);
  not g7695 (n_1648, n6042);
  not g7696 (n_1649, n6135);
  and g7697 (n6136, n_1648, n_1649);
  not g7698 (n_1650, n6043);
  and g7699 (n6137, n_1650, n6136);
  not g7700 (n_1651, n6137);
  and g7701 (n6138, n_1648, n_1651);
  and g7702 (n6139, \a[5] , n5829);
  not g7703 (n_1652, n6139);
  and g7704 (n6140, n_1470, n_1652);
  not g7705 (n_1653, n6138);
  and g7706 (n6141, n_1653, n6140);
  not g7707 (n_1654, n2866);
  and g7708 (n6142, n2864, n_1654);
  not g7709 (n_1655, n6142);
  and g7710 (n6143, n_354, n_1655);
  and g7711 (n6144, n75, n6143);
  and g7712 (n6145, n_305, n3020);
  and g7713 (n6146, n_307, n3023);
  and g7714 (n6147, n_306, n3028);
  not g7722 (n_1660, n6140);
  and g7723 (n6151, n6138, n_1660);
  not g7724 (n_1661, n6141);
  not g7725 (n_1662, n6151);
  and g7726 (n6152, n_1661, n_1662);
  not g7727 (n_1663, n6150);
  and g7728 (n6153, n_1663, n6152);
  not g7729 (n_1664, n6153);
  and g7730 (n6154, n_1661, n_1664);
  not g7731 (n_1665, n6015);
  not g7732 (n_1666, n6154);
  and g7733 (n6155, n_1665, n_1666);
  and g7734 (n6156, n6015, n6154);
  not g7735 (n_1667, n6155);
  not g7736 (n_1668, n6156);
  and g7737 (n6157, n_1667, n_1668);
  and g7738 (n6158, n_301, n3457);
  and g7739 (n6159, n_303, n3542);
  and g7740 (n6160, n_302, n3606);
  not g7741 (n_1669, n6159);
  not g7742 (n_1670, n6160);
  and g7743 (n6161, n_1669, n_1670);
  not g7744 (n_1671, n6158);
  and g7745 (n6162, n_1671, n6161);
  and g7746 (n6163, n_489, n6162);
  not g7747 (n_1672, n5328);
  and g7748 (n6164, n_1672, n6162);
  not g7749 (n_1673, n6163);
  not g7750 (n_1674, n6164);
  and g7751 (n6165, n_1673, n_1674);
  not g7752 (n_1675, n6165);
  and g7753 (n6166, \a[29] , n_1675);
  and g7754 (n6167, n_15, n6165);
  not g7755 (n_1676, n6166);
  not g7756 (n_1677, n6167);
  and g7757 (n6168, n_1676, n_1677);
  not g7758 (n_1678, n6168);
  and g7759 (n6169, n6157, n_1678);
  not g7760 (n_1679, n6169);
  and g7761 (n6170, n_1667, n_1679);
  not g7762 (n_1680, n6012);
  and g7763 (n6171, n_1627, n_1680);
  and g7764 (n6172, n_1628, n_1680);
  not g7765 (n_1681, n6171);
  not g7766 (n_1682, n6172);
  and g7767 (n6173, n_1681, n_1682);
  not g7768 (n_1683, n6170);
  not g7769 (n_1684, n6173);
  and g7770 (n6174, n_1683, n_1684);
  not g7771 (n_1685, n6174);
  and g7772 (n6175, n_1680, n_1685);
  not g7773 (n_1686, n5999);
  not g7774 (n_1687, n6175);
  and g7775 (n6176, n_1686, n_1687);
  not g7776 (n_1688, n6176);
  and g7777 (n6177, n_1616, n_1688);
  not g7778 (n_1689, n5865);
  and g7779 (n6178, n_1689, n5876);
  not g7780 (n_1690, n6178);
  and g7781 (n6179, n_1512, n_1690);
  not g7782 (n_1691, n6177);
  and g7783 (n6180, n_1691, n6179);
  not g7784 (n_1692, n6179);
  and g7785 (n6181, n6177, n_1692);
  not g7786 (n_1693, n6180);
  not g7787 (n_1694, n6181);
  and g7788 (n6182, n_1693, n_1694);
  and g7789 (n6183, n_286, n3884);
  and g7790 (n6184, n_295, n3967);
  and g7791 (n6185, n_293, n4046);
  and g7797 (n6188, n4050, n4429);
  not g7800 (n_1699, n6189);
  and g7801 (n6190, \a[26] , n_1699);
  not g7802 (n_1700, n6190);
  and g7803 (n6191, \a[26] , n_1700);
  and g7804 (n6192, n_1699, n_1700);
  not g7805 (n_1701, n6191);
  not g7806 (n_1702, n6192);
  and g7807 (n6193, n_1701, n_1702);
  not g7808 (n_1703, n6193);
  and g7809 (n6194, n6182, n_1703);
  not g7810 (n_1704, n6194);
  and g7811 (n6195, n_1693, n_1704);
  not g7812 (n_1705, n5981);
  not g7813 (n_1706, n6195);
  and g7814 (n6196, n_1705, n_1706);
  and g7815 (n6197, n5981, n6195);
  not g7816 (n_1707, n6196);
  not g7817 (n_1708, n6197);
  and g7818 (n6198, n_1707, n_1708);
  and g7819 (n6199, n_237, n4694);
  and g7820 (n6200, n_275, n4533);
  and g7821 (n6201, n_260, n4604);
  and g7827 (n6204, n3331, n4536);
  not g7830 (n_1713, n6205);
  and g7831 (n6206, \a[23] , n_1713);
  not g7832 (n_1714, n6206);
  and g7833 (n6207, \a[23] , n_1714);
  and g7834 (n6208, n_1713, n_1714);
  not g7835 (n_1715, n6207);
  not g7836 (n_1716, n6208);
  and g7837 (n6209, n_1715, n_1716);
  not g7838 (n_1717, n6209);
  and g7839 (n6210, n6198, n_1717);
  not g7840 (n_1718, n6210);
  and g7841 (n6211, n_1707, n_1718);
  not g7842 (n_1719, n5978);
  not g7843 (n_1720, n6211);
  and g7844 (n6212, n_1719, n_1720);
  not g7845 (n_1721, n6212);
  and g7846 (n6213, n_1599, n_1721);
  not g7847 (n_1722, n5961);
  not g7848 (n_1723, n6213);
  and g7849 (n6214, n_1722, n_1723);
  and g7850 (n6215, n5961, n6213);
  not g7851 (n_1724, n6214);
  not g7852 (n_1725, n6215);
  and g7853 (n6216, n_1724, n_1725);
  and g7854 (n6217, n_480, n5496);
  and g7855 (n6218, n_484, n4935);
  and g7856 (n6219, n_485, n5407);
  and g7862 (n6222, n3627, n4938);
  not g7865 (n_1730, n6223);
  and g7866 (n6224, \a[20] , n_1730);
  not g7867 (n_1731, n6224);
  and g7868 (n6225, \a[20] , n_1731);
  and g7869 (n6226, n_1730, n_1731);
  not g7870 (n_1732, n6225);
  not g7871 (n_1733, n6226);
  and g7872 (n6227, n_1732, n_1733);
  not g7873 (n_1734, n6227);
  and g7874 (n6228, n6216, n_1734);
  not g7875 (n_1735, n6228);
  and g7876 (n6229, n_1724, n_1735);
  not g7877 (n_1736, n5958);
  not g7878 (n_1737, n6229);
  and g7879 (n6230, n_1736, n_1737);
  and g7880 (n6231, n5958, n6229);
  not g7881 (n_1738, n6230);
  not g7882 (n_1739, n6231);
  and g7883 (n6232, n_1738, n_1739);
  and g7884 (n6233, n_1408, n5661);
  and g7885 (n6234, n_560, n6233);
  and g7886 (n6235, n_565, n5663);
  and g7887 (n6236, n_566, n5939);
  and g7893 (n6239, n4067, n5666);
  not g7896 (n_1744, n6240);
  and g7897 (n6241, \a[17] , n_1744);
  not g7898 (n_1745, n6241);
  and g7899 (n6242, \a[17] , n_1745);
  and g7900 (n6243, n_1744, n_1745);
  not g7901 (n_1746, n6242);
  not g7902 (n_1747, n6243);
  and g7903 (n6244, n_1746, n_1747);
  not g7904 (n_1748, n6244);
  and g7905 (n6245, n6232, n_1748);
  not g7906 (n_1749, n6245);
  and g7907 (n6246, n_1738, n_1749);
  and g7908 (n6247, n_712, n6233);
  and g7909 (n6248, n_566, n5663);
  and g7910 (n6249, n_560, n5939);
  not g7911 (n_1750, n6248);
  not g7912 (n_1751, n6249);
  and g7913 (n6250, n_1750, n_1751);
  not g7914 (n_1752, n6247);
  and g7915 (n6251, n_1752, n6250);
  and g7916 (n6252, n_1409, n6251);
  and g7917 (n6253, n_888, n6251);
  not g7918 (n_1753, n6252);
  not g7919 (n_1754, n6253);
  and g7920 (n6254, n_1753, n_1754);
  not g7921 (n_1755, n6254);
  and g7922 (n6255, \a[17] , n_1755);
  and g7923 (n6256, n_617, n6254);
  not g7924 (n_1756, n6255);
  not g7925 (n_1757, n6256);
  and g7926 (n6257, n_1756, n_1757);
  not g7927 (n_1758, n6246);
  not g7928 (n_1759, n6257);
  and g7929 (n6258, n_1758, n_1759);
  and g7930 (n6259, n6246, n6257);
  not g7931 (n_1760, n6258);
  not g7932 (n_1761, n6259);
  and g7933 (n6260, n_1760, n_1761);
  not g7934 (n_1762, n5932);
  and g7935 (n6261, n5930, n_1762);
  not g7936 (n_1763, n6261);
  and g7937 (n6262, n_1563, n_1763);
  and g7938 (n6263, n6260, n6262);
  not g7939 (n_1764, n6263);
  and g7940 (n6264, n_1760, n_1764);
  not g7941 (n_1765, n5955);
  not g7942 (n_1766, n6264);
  and g7943 (n6265, n_1765, n_1766);
  and g7944 (n6266, n5955, n6264);
  not g7945 (n_1767, n6265);
  not g7946 (n_1768, n6266);
  and g7947 (n6267, n_1767, n_1768);
  and g7948 (n6268, n6216, n_1735);
  and g7949 (n6269, n_1734, n_1735);
  not g7950 (n_1769, n6268);
  not g7951 (n_1770, n6269);
  and g7952 (n6270, n_1769, n_1770);
  and g7953 (n6271, n5978, n6211);
  not g7954 (n_1771, n6271);
  and g7955 (n6272, n_1721, n_1771);
  and g7956 (n6273, n_485, n5496);
  and g7957 (n6274, n_415, n4935);
  and g7958 (n6275, n_484, n5407);
  not g7959 (n_1772, n6274);
  not g7960 (n_1773, n6275);
  and g7961 (n6276, n_1772, n_1773);
  not g7962 (n_1774, n6273);
  and g7963 (n6277, n_1774, n6276);
  and g7964 (n6278, n_1011, n6277);
  and g7965 (n6279, n_914, n6277);
  not g7966 (n_1775, n6278);
  not g7967 (n_1776, n6279);
  and g7968 (n6280, n_1775, n_1776);
  not g7969 (n_1777, n6280);
  and g7970 (n6281, \a[20] , n_1777);
  and g7971 (n6282, n_435, n6280);
  not g7972 (n_1778, n6281);
  not g7973 (n_1779, n6282);
  and g7974 (n6283, n_1778, n_1779);
  not g7975 (n_1780, n6283);
  and g7976 (n6284, n6272, n_1780);
  and g7977 (n6285, n6198, n_1718);
  and g7978 (n6286, n_1717, n_1718);
  not g7979 (n_1781, n6285);
  not g7980 (n_1782, n6286);
  and g7981 (n6287, n_1781, n_1782);
  and g7982 (n6288, n6182, n_1704);
  and g7983 (n6289, n_1703, n_1704);
  not g7984 (n_1783, n6288);
  not g7985 (n_1784, n6289);
  and g7986 (n6290, n_1783, n_1784);
  and g7987 (n6291, n5999, n6175);
  not g7988 (n_1785, n6291);
  and g7989 (n6292, n_1688, n_1785);
  and g7990 (n6293, n_293, n3884);
  and g7991 (n6294, n_298, n3967);
  and g7992 (n6295, n_295, n4046);
  not g7993 (n_1786, n6294);
  not g7994 (n_1787, n6295);
  and g7995 (n6296, n_1786, n_1787);
  not g7996 (n_1788, n6293);
  and g7997 (n6297, n_1788, n6296);
  and g7998 (n6298, n_750, n6297);
  not g7999 (n_1789, n4861);
  and g8000 (n6299, n_1789, n6297);
  not g8001 (n_1790, n6298);
  not g8002 (n_1791, n6299);
  and g8003 (n6300, n_1790, n_1791);
  not g8004 (n_1792, n6300);
  and g8005 (n6301, \a[26] , n_1792);
  and g8006 (n6302, n_33, n6300);
  not g8007 (n_1793, n6301);
  not g8008 (n_1794, n6302);
  and g8009 (n6303, n_1793, n_1794);
  not g8010 (n_1795, n6303);
  and g8011 (n6304, n6292, n_1795);
  and g8012 (n6305, n_1683, n_1685);
  and g8013 (n6306, n_1684, n_1685);
  not g8014 (n_1796, n6305);
  not g8015 (n_1797, n6306);
  and g8016 (n6307, n_1796, n_1797);
  and g8017 (n6308, n_300, n3457);
  and g8018 (n6309, n_302, n3542);
  and g8019 (n6310, n_301, n3606);
  not g8020 (n_1798, n6309);
  not g8021 (n_1799, n6310);
  and g8022 (n6311, n_1798, n_1799);
  not g8023 (n_1800, n6308);
  and g8024 (n6312, n_1800, n6311);
  and g8025 (n6313, n_489, n6312);
  not g8026 (n_1801, n5561);
  and g8027 (n6314, n_1801, n6312);
  not g8028 (n_1802, n6313);
  not g8029 (n_1803, n6314);
  and g8030 (n6315, n_1802, n_1803);
  not g8031 (n_1804, n6315);
  and g8032 (n6316, \a[29] , n_1804);
  and g8033 (n6317, n_15, n6315);
  not g8034 (n_1805, n6316);
  not g8035 (n_1806, n6317);
  and g8036 (n6318, n_1805, n_1806);
  not g8037 (n_1807, n6307);
  not g8038 (n_1808, n6318);
  and g8039 (n6319, n_1807, n_1808);
  and g8040 (n6320, n6307, n6318);
  not g8041 (n_1809, n6319);
  not g8042 (n_1810, n6320);
  and g8043 (n6321, n_1809, n_1810);
  and g8044 (n6322, n_295, n3884);
  and g8045 (n6323, n_299, n3967);
  and g8046 (n6324, n_298, n4046);
  and g8052 (n6327, n4050, n4848);
  not g8055 (n_1815, n6328);
  and g8056 (n6329, \a[26] , n_1815);
  not g8057 (n_1816, n6329);
  and g8058 (n6330, \a[26] , n_1816);
  and g8059 (n6331, n_1815, n_1816);
  not g8060 (n_1817, n6330);
  not g8061 (n_1818, n6331);
  and g8062 (n6332, n_1817, n_1818);
  not g8063 (n_1819, n6332);
  and g8064 (n6333, n6321, n_1819);
  not g8065 (n_1820, n6333);
  and g8066 (n6334, n_1809, n_1820);
  not g8067 (n_1821, n6292);
  and g8068 (n6335, n_1821, n6303);
  not g8069 (n_1822, n6304);
  not g8070 (n_1823, n6335);
  and g8071 (n6336, n_1822, n_1823);
  not g8072 (n_1824, n6334);
  and g8073 (n6337, n_1824, n6336);
  not g8074 (n_1825, n6337);
  and g8075 (n6338, n_1822, n_1825);
  not g8076 (n_1826, n6290);
  not g8077 (n_1827, n6338);
  and g8078 (n6339, n_1826, n_1827);
  and g8079 (n6340, n6290, n6338);
  not g8080 (n_1828, n6339);
  not g8081 (n_1829, n6340);
  and g8082 (n6341, n_1828, n_1829);
  and g8083 (n6342, n_260, n4694);
  and g8084 (n6343, n_281, n4533);
  and g8085 (n6344, n_275, n4604);
  and g8091 (n6347, n4179, n4536);
  not g8094 (n_1834, n6348);
  and g8095 (n6349, \a[23] , n_1834);
  not g8096 (n_1835, n6349);
  and g8097 (n6350, \a[23] , n_1835);
  and g8098 (n6351, n_1834, n_1835);
  not g8099 (n_1836, n6350);
  not g8100 (n_1837, n6351);
  and g8101 (n6352, n_1836, n_1837);
  not g8102 (n_1838, n6352);
  and g8103 (n6353, n6341, n_1838);
  not g8104 (n_1839, n6353);
  and g8105 (n6354, n_1828, n_1839);
  not g8106 (n_1840, n6287);
  not g8107 (n_1841, n6354);
  and g8108 (n6355, n_1840, n_1841);
  and g8109 (n6356, n6287, n6354);
  not g8110 (n_1842, n6355);
  not g8111 (n_1843, n6356);
  and g8112 (n6357, n_1842, n_1843);
  and g8113 (n6358, n_484, n5496);
  and g8114 (n6359, n_236, n4935);
  and g8115 (n6360, n_415, n5407);
  and g8121 (n6363, n3715, n4938);
  not g8124 (n_1848, n6364);
  and g8125 (n6365, \a[20] , n_1848);
  not g8126 (n_1849, n6365);
  and g8127 (n6366, \a[20] , n_1849);
  and g8128 (n6367, n_1848, n_1849);
  not g8129 (n_1850, n6366);
  not g8130 (n_1851, n6367);
  and g8131 (n6368, n_1850, n_1851);
  not g8132 (n_1852, n6368);
  and g8133 (n6369, n6357, n_1852);
  not g8134 (n_1853, n6369);
  and g8135 (n6370, n_1842, n_1853);
  not g8136 (n_1854, n6272);
  and g8137 (n6371, n_1854, n6283);
  not g8138 (n_1855, n6284);
  not g8139 (n_1856, n6371);
  and g8140 (n6372, n_1855, n_1856);
  not g8141 (n_1857, n6370);
  and g8142 (n6373, n_1857, n6372);
  not g8143 (n_1858, n6373);
  and g8144 (n6374, n_1855, n_1858);
  not g8145 (n_1859, n6270);
  not g8146 (n_1860, n6374);
  and g8147 (n6375, n_1859, n_1860);
  and g8148 (n6376, n6270, n6374);
  not g8149 (n_1861, n6375);
  not g8150 (n_1862, n6376);
  and g8151 (n6377, n_1861, n_1862);
  and g8152 (n6378, n_566, n6233);
  and g8153 (n6379, n_535, n5663);
  and g8154 (n6380, n_565, n5939);
  and g8160 (n6383, n4477, n5666);
  not g8163 (n_1867, n6384);
  and g8164 (n6385, \a[17] , n_1867);
  not g8165 (n_1868, n6385);
  and g8166 (n6386, \a[17] , n_1868);
  and g8167 (n6387, n_1867, n_1868);
  not g8168 (n_1869, n6386);
  not g8169 (n_1870, n6387);
  and g8170 (n6388, n_1869, n_1870);
  not g8171 (n_1871, n6388);
  and g8172 (n6389, n6377, n_1871);
  not g8173 (n_1872, n6389);
  and g8174 (n6390, n_1861, n_1872);
  not g8175 (n_1874, \a[12] );
  and g8176 (n6391, \a[11] , n_1874);
  and g8177 (n6392, n_1071, \a[12] );
  not g8178 (n_1875, n6391);
  not g8179 (n_1876, n6392);
  and g8180 (n6393, n_1875, n_1876);
  and g8181 (n6394, \a[13] , n_652);
  not g8182 (n_1878, \a[13] );
  and g8183 (n6395, n_1878, \a[14] );
  not g8184 (n_1879, n6394);
  not g8185 (n_1880, n6395);
  and g8186 (n6396, n_1879, n_1880);
  not g8187 (n_1881, n6393);
  not g8188 (n_1882, n6396);
  and g8189 (n6397, n_1881, n_1882);
  and g8190 (n6398, n_1874, \a[13] );
  and g8191 (n6399, \a[12] , n_1878);
  not g8192 (n_1883, n6398);
  not g8193 (n_1884, n6399);
  and g8194 (n6400, n_1883, n_1884);
  and g8195 (n6401, n6393, n_1882);
  and g8196 (n6402, n6400, n6401);
  and g8197 (n6403, n_712, n6402);
  not g8198 (n_1885, n6397);
  not g8199 (n_1886, n6403);
  and g8200 (n6404, n_1885, n_1886);
  and g8201 (n6405, n_729, n_1886);
  not g8202 (n_1887, n6404);
  not g8203 (n_1888, n6405);
  and g8204 (n6406, n_1887, n_1888);
  not g8205 (n_1889, n6406);
  and g8206 (n6407, \a[14] , n_1889);
  and g8207 (n6408, n_652, n6406);
  not g8208 (n_1890, n6407);
  not g8209 (n_1891, n6408);
  and g8210 (n6409, n_1890, n_1891);
  not g8211 (n_1892, n6390);
  not g8212 (n_1893, n6409);
  and g8213 (n6410, n_1892, n_1893);
  and g8214 (n6411, n6232, n_1749);
  and g8215 (n6412, n_1748, n_1749);
  not g8216 (n_1894, n6411);
  not g8217 (n_1895, n6412);
  and g8218 (n6413, n_1894, n_1895);
  and g8219 (n6414, n6390, n6409);
  not g8220 (n_1896, n6410);
  not g8221 (n_1897, n6414);
  and g8222 (n6415, n_1896, n_1897);
  not g8223 (n_1898, n6413);
  and g8224 (n6416, n_1898, n6415);
  not g8225 (n_1899, n6416);
  and g8226 (n6417, n_1896, n_1899);
  not g8227 (n_1900, n6260);
  not g8228 (n_1901, n6262);
  and g8229 (n6418, n_1900, n_1901);
  not g8230 (n_1902, n6418);
  and g8231 (n6419, n_1764, n_1902);
  not g8232 (n_1903, n6417);
  and g8233 (n6420, n_1903, n6419);
  not g8234 (n_1904, n6419);
  and g8235 (n6421, n6417, n_1904);
  not g8236 (n_1905, n6420);
  not g8237 (n_1906, n6421);
  and g8238 (n6422, n_1905, n_1906);
  and g8239 (n6423, n_1898, n_1899);
  and g8240 (n6424, n6415, n_1899);
  not g8241 (n_1907, n6423);
  not g8242 (n_1908, n6424);
  and g8243 (n6425, n_1907, n_1908);
  and g8244 (n6426, n_565, n6233);
  and g8245 (n6427, n_480, n5663);
  and g8246 (n6428, n_535, n5939);
  and g8252 (n6431, n4558, n5666);
  not g8255 (n_1913, n6432);
  and g8256 (n6433, \a[17] , n_1913);
  not g8257 (n_1914, n6433);
  and g8258 (n6434, n_1913, n_1914);
  and g8259 (n6435, \a[17] , n_1914);
  not g8260 (n_1915, n6434);
  not g8261 (n_1916, n6435);
  and g8262 (n6436, n_1915, n_1916);
  not g8263 (n_1917, n6372);
  and g8264 (n6437, n6370, n_1917);
  not g8265 (n_1918, n6437);
  and g8266 (n6438, n_1858, n_1918);
  not g8267 (n_1919, n6436);
  and g8268 (n6439, n_1919, n6438);
  not g8269 (n_1920, n6439);
  and g8270 (n6440, n_1919, n_1920);
  and g8271 (n6441, n6438, n_1920);
  not g8272 (n_1921, n6440);
  not g8273 (n_1922, n6441);
  and g8274 (n6442, n_1921, n_1922);
  and g8275 (n6443, n6357, n_1853);
  and g8276 (n6444, n_1852, n_1853);
  not g8277 (n_1923, n6443);
  not g8278 (n_1924, n6444);
  and g8279 (n6445, n_1923, n_1924);
  and g8280 (n6446, n6341, n_1839);
  and g8281 (n6447, n_1838, n_1839);
  not g8282 (n_1925, n6446);
  not g8283 (n_1926, n6447);
  and g8284 (n6448, n_1925, n_1926);
  and g8285 (n6449, n_275, n4694);
  and g8286 (n6450, n_286, n4533);
  and g8287 (n6451, n_281, n4604);
  and g8293 (n6454, n4204, n4536);
  not g8296 (n_1931, n6455);
  and g8297 (n6456, \a[23] , n_1931);
  not g8298 (n_1932, n6456);
  and g8299 (n6457, n_1931, n_1932);
  and g8300 (n6458, \a[23] , n_1932);
  not g8301 (n_1933, n6457);
  not g8302 (n_1934, n6458);
  and g8303 (n6459, n_1933, n_1934);
  not g8304 (n_1935, n6336);
  and g8305 (n6460, n6334, n_1935);
  not g8306 (n_1936, n6460);
  and g8307 (n6461, n_1825, n_1936);
  not g8308 (n_1937, n6459);
  and g8309 (n6462, n_1937, n6461);
  not g8310 (n_1938, n6462);
  and g8311 (n6463, n_1937, n_1938);
  and g8312 (n6464, n6461, n_1938);
  not g8313 (n_1939, n6463);
  not g8314 (n_1940, n6464);
  and g8315 (n6465, n_1939, n_1940);
  and g8316 (n6466, n6321, n_1820);
  and g8317 (n6467, n_1819, n_1820);
  not g8318 (n_1941, n6466);
  not g8319 (n_1942, n6467);
  and g8320 (n6468, n_1941, n_1942);
  and g8321 (n6469, n6152, n_1664);
  and g8322 (n6470, n_1663, n_1664);
  not g8323 (n_1943, n6469);
  not g8324 (n_1944, n6470);
  and g8325 (n6471, n_1943, n_1944);
  and g8326 (n6472, n_1649, n_1651);
  and g8327 (n6473, n_1650, n6138);
  not g8328 (n_1945, n6472);
  not g8329 (n_1946, n6473);
  and g8330 (n6474, n_1945, n_1946);
  and g8331 (n6475, n_306, n3020);
  and g8332 (n6476, n_307, n3028);
  and g8333 (n6477, n_308, n3023);
  not g8334 (n_1947, n2862);
  and g8335 (n6478, n2860, n_1947);
  not g8336 (n_1948, n6478);
  and g8337 (n6479, n_350, n_1948);
  and g8338 (n6480, n75, n6479);
  not g8346 (n_1953, n6474);
  not g8347 (n_1954, n6483);
  and g8348 (n6484, n_1953, n_1954);
  and g8349 (n6485, n_1645, n_1647);
  and g8350 (n6486, n_1646, n6135);
  not g8351 (n_1955, n6485);
  not g8352 (n_1956, n6486);
  and g8353 (n6487, n_1955, n_1956);
  and g8354 (n6488, n_307, n3020);
  and g8355 (n6489, n_308, n3028);
  and g8356 (n6490, n_309, n3023);
  not g8357 (n_1957, n2858);
  and g8358 (n6491, n2856, n_1957);
  not g8359 (n_1958, n6491);
  and g8360 (n6492, n_346, n_1958);
  and g8361 (n6493, n75, n6492);
  not g8369 (n_1963, n6487);
  not g8370 (n_1964, n6496);
  and g8371 (n6497, n_1963, n_1964);
  and g8372 (n6498, n_1641, n_1643);
  and g8373 (n6499, n_1642, n6132);
  not g8374 (n_1965, n6498);
  not g8375 (n_1966, n6499);
  and g8376 (n6500, n_1965, n_1966);
  and g8413 (n6537, n_309, n3020);
  and g8414 (n6538, n_310, n3028);
  and g8415 (n6539, n_311, n3023);
  not g8416 (n_1967, n2850);
  and g8417 (n6540, n2848, n_1967);
  not g8418 (n_1968, n6540);
  and g8419 (n6541, n_338, n_1968);
  and g8420 (n6542, n75, n6541);
  not g8428 (n_1973, n6536);
  not g8429 (n_1974, n6545);
  and g8430 (n6546, n_1973, n_1974);
  and g8431 (n6547, n_111, n_175);
  and g8432 (n6548, n_219, n6547);
  and g8450 (n6566, n_115, n1128);
  and g8451 (n6567, n_197, n6566);
  and g8471 (n6587, n_310, n3020);
  and g8472 (n6588, n_311, n3028);
  and g8473 (n6589, n_312, n3023);
  not g8474 (n_1975, n2846);
  and g8475 (n6590, n2844, n_1975);
  not g8476 (n_1976, n6590);
  and g8477 (n6591, n_334, n_1976);
  and g8478 (n6592, n75, n6591);
  not g8486 (n_1981, n6586);
  not g8487 (n_1982, n6595);
  and g8488 (n6596, n_1981, n_1982);
  and g8534 (n6642, n_311, n3020);
  and g8535 (n6643, n_312, n3028);
  and g8536 (n6644, n_313, n3023);
  not g8537 (n_1983, n2842);
  and g8538 (n6645, n2840, n_1983);
  not g8539 (n_1984, n6645);
  and g8540 (n6646, n_330, n_1984);
  and g8541 (n6647, n75, n6646);
  not g8549 (n_1989, n6641);
  not g8550 (n_1990, n6650);
  and g8551 (n6651, n_1989, n_1990);
  and g8563 (n6663, n_155, n_213);
  and g8564 (n6664, n_183, n6663);
  and g8571 (n6671, n_112, n604);
  and g8572 (n6672, n_139, n6671);
  and g8591 (n6691, n_312, n3020);
  and g8592 (n6692, n_313, n3028);
  and g8593 (n6693, n_314, n3023);
  not g8594 (n_1991, n2838);
  and g8595 (n6694, n2836, n_1991);
  not g8596 (n_1992, n6694);
  and g8597 (n6695, n_326, n_1992);
  and g8598 (n6696, n75, n6695);
  not g8606 (n_1997, n6690);
  not g8607 (n_1998, n6699);
  and g8608 (n6700, n_1997, n_1998);
  and g8614 (n6706, n_83, n_63);
  and g8615 (n6707, n_222, n6706);
  and g8623 (n6715, n_45, n3581);
  and g8624 (n6716, n_73, n6715);
  and g8625 (n6717, n_225, n2089);
  and g8641 (n6733, n_91, n885);
  and g8642 (n6734, n_84, n6733);
  and g8678 (n6770, n_292, n3636);
  and g8679 (n6771, n_247, n6770);
  and g8700 (n6792, n_314, n3020);
  and g8701 (n6793, n_315, n3028);
  and g8702 (n6794, n_316, n3023);
  and g8703 (n6795, n_315, n2829);
  not g8704 (n_1999, n6795);
  and g8705 (n6796, n2674, n_1999);
  and g8706 (n6797, n2737, n2829);
  not g8707 (n_2000, n6796);
  not g8708 (n_2001, n6797);
  and g8709 (n6798, n_2000, n_2001);
  and g8710 (n6799, n75, n6798);
  not g8718 (n_2006, n6791);
  not g8719 (n_2007, n6802);
  and g8720 (n6803, n_2006, n_2007);
  not g8721 (n_2008, n6748);
  and g8722 (n6804, n_2008, n6803);
  not g8723 (n_2009, n2834);
  and g8724 (n6805, n2832, n_2009);
  not g8725 (n_2010, n6805);
  and g8726 (n6806, n_322, n_2010);
  and g8727 (n6807, n75, n6806);
  and g8728 (n6808, n_313, n3020);
  and g8729 (n6809, n_315, n3023);
  and g8730 (n6810, n_314, n3028);
  not g8738 (n_2015, n6803);
  and g8739 (n6814, n6748, n_2015);
  not g8740 (n_2016, n6804);
  not g8741 (n_2017, n6814);
  and g8742 (n6815, n_2016, n_2017);
  not g8743 (n_2018, n6813);
  and g8744 (n6816, n_2018, n6815);
  not g8745 (n_2019, n6816);
  and g8746 (n6817, n_2016, n_2019);
  not g8747 (n_2020, n6700);
  and g8748 (n6818, n_1997, n_2020);
  and g8749 (n6819, n_1998, n_2020);
  not g8750 (n_2021, n6818);
  not g8751 (n_2022, n6819);
  and g8752 (n6820, n_2021, n_2022);
  not g8753 (n_2023, n6817);
  not g8754 (n_2024, n6820);
  and g8755 (n6821, n_2023, n_2024);
  not g8756 (n_2025, n6821);
  and g8757 (n6822, n_2020, n_2025);
  not g8758 (n_2026, n6651);
  and g8759 (n6823, n_1989, n_2026);
  and g8760 (n6824, n_1990, n_2026);
  not g8761 (n_2027, n6823);
  not g8762 (n_2028, n6824);
  and g8763 (n6825, n_2027, n_2028);
  not g8764 (n_2029, n6822);
  not g8765 (n_2030, n6825);
  and g8766 (n6826, n_2029, n_2030);
  not g8767 (n_2031, n6826);
  and g8768 (n6827, n_2026, n_2031);
  not g8769 (n_2032, n6596);
  and g8770 (n6828, n_1981, n_2032);
  and g8771 (n6829, n_1982, n_2032);
  not g8772 (n_2033, n6828);
  not g8773 (n_2034, n6829);
  and g8774 (n6830, n_2033, n_2034);
  not g8775 (n_2035, n6827);
  not g8776 (n_2036, n6830);
  and g8777 (n6831, n_2035, n_2036);
  not g8778 (n_2037, n6831);
  and g8779 (n6832, n_2032, n_2037);
  not g8780 (n_2038, n6546);
  and g8781 (n6833, n_1973, n_2038);
  and g8782 (n6834, n_1974, n_2038);
  not g8783 (n_2039, n6833);
  not g8784 (n_2040, n6834);
  and g8785 (n6835, n_2039, n_2040);
  not g8786 (n_2041, n6832);
  not g8787 (n_2042, n6835);
  and g8788 (n6836, n_2041, n_2042);
  not g8789 (n_2043, n6836);
  and g8790 (n6837, n_2038, n_2043);
  not g8791 (n_2044, n6500);
  not g8792 (n_2045, n6837);
  and g8793 (n6838, n_2044, n_2045);
  and g8794 (n6839, n6500, n6837);
  not g8795 (n_2046, n6838);
  not g8796 (n_2047, n6839);
  and g8797 (n6840, n_2046, n_2047);
  and g8798 (n6841, n_305, n3457);
  and g8799 (n6842, n_307, n3542);
  and g8800 (n6843, n_306, n3606);
  not g8801 (n_2048, n6842);
  not g8802 (n_2049, n6843);
  and g8803 (n6844, n_2048, n_2049);
  not g8804 (n_2050, n6841);
  and g8805 (n6845, n_2050, n6844);
  and g8806 (n6846, n_489, n6845);
  not g8807 (n_2051, n6143);
  and g8808 (n6847, n_2051, n6845);
  not g8809 (n_2052, n6846);
  not g8810 (n_2053, n6847);
  and g8811 (n6848, n_2052, n_2053);
  not g8812 (n_2054, n6848);
  and g8813 (n6849, \a[29] , n_2054);
  and g8814 (n6850, n_15, n6848);
  not g8815 (n_2055, n6849);
  not g8816 (n_2056, n6850);
  and g8817 (n6851, n_2055, n_2056);
  not g8818 (n_2057, n6851);
  and g8819 (n6852, n6840, n_2057);
  not g8820 (n_2058, n6852);
  and g8821 (n6853, n_2046, n_2058);
  not g8822 (n_2059, n6497);
  and g8823 (n6854, n_1963, n_2059);
  and g8824 (n6855, n_1964, n_2059);
  not g8825 (n_2060, n6854);
  not g8826 (n_2061, n6855);
  and g8827 (n6856, n_2060, n_2061);
  not g8828 (n_2062, n6853);
  not g8829 (n_2063, n6856);
  and g8830 (n6857, n_2062, n_2063);
  not g8831 (n_2064, n6857);
  and g8832 (n6858, n_2059, n_2064);
  not g8833 (n_2065, n6484);
  and g8834 (n6859, n_1953, n_2065);
  and g8835 (n6860, n_1954, n_2065);
  not g8836 (n_2066, n6859);
  not g8837 (n_2067, n6860);
  and g8838 (n6861, n_2066, n_2067);
  not g8839 (n_2068, n6858);
  not g8840 (n_2069, n6861);
  and g8841 (n6862, n_2068, n_2069);
  not g8842 (n_2070, n6862);
  and g8843 (n6863, n_2065, n_2070);
  not g8844 (n_2071, n6471);
  not g8845 (n_2072, n6863);
  and g8846 (n6864, n_2071, n_2072);
  and g8847 (n6865, n6471, n6863);
  not g8848 (n_2073, n6864);
  not g8849 (n_2074, n6865);
  and g8850 (n6866, n_2073, n_2074);
  and g8851 (n6867, n_302, n3457);
  and g8852 (n6868, n_304, n3542);
  and g8853 (n6869, n_303, n3606);
  and g8859 (n6872, n3368, n5851);
  not g8862 (n_2079, n6873);
  and g8863 (n6874, \a[29] , n_2079);
  not g8864 (n_2080, n6874);
  and g8865 (n6875, \a[29] , n_2080);
  and g8866 (n6876, n_2079, n_2080);
  not g8867 (n_2081, n6875);
  not g8868 (n_2082, n6876);
  and g8869 (n6877, n_2081, n_2082);
  not g8870 (n_2083, n6877);
  and g8871 (n6878, n6866, n_2083);
  not g8872 (n_2084, n6878);
  and g8873 (n6879, n_2073, n_2084);
  not g8874 (n_2085, n6157);
  and g8875 (n6880, n_2085, n6168);
  not g8876 (n_2086, n6880);
  and g8877 (n6881, n_1679, n_2086);
  not g8878 (n_2087, n6879);
  and g8879 (n6882, n_2087, n6881);
  not g8880 (n_2088, n6881);
  and g8881 (n6883, n6879, n_2088);
  not g8882 (n_2089, n6882);
  not g8883 (n_2090, n6883);
  and g8884 (n6884, n_2089, n_2090);
  and g8885 (n6885, n_298, n3884);
  and g8886 (n6886, n_300, n3967);
  and g8887 (n6887, n_299, n4046);
  and g8893 (n6890, n4050, n5114);
  not g8896 (n_2095, n6891);
  and g8897 (n6892, \a[26] , n_2095);
  not g8898 (n_2096, n6892);
  and g8899 (n6893, \a[26] , n_2096);
  and g8900 (n6894, n_2095, n_2096);
  not g8901 (n_2097, n6893);
  not g8902 (n_2098, n6894);
  and g8903 (n6895, n_2097, n_2098);
  not g8904 (n_2099, n6895);
  and g8905 (n6896, n6884, n_2099);
  not g8906 (n_2100, n6896);
  and g8907 (n6897, n_2089, n_2100);
  not g8908 (n_2101, n6468);
  not g8909 (n_2102, n6897);
  and g8910 (n6898, n_2101, n_2102);
  and g8911 (n6899, n6468, n6897);
  not g8912 (n_2103, n6898);
  not g8913 (n_2104, n6899);
  and g8914 (n6900, n_2103, n_2104);
  and g8915 (n6901, n_281, n4694);
  and g8916 (n6902, n_293, n4533);
  and g8917 (n6903, n_286, n4604);
  and g8923 (n6906, n4536, n4633);
  not g8926 (n_2109, n6907);
  and g8927 (n6908, \a[23] , n_2109);
  not g8928 (n_2110, n6908);
  and g8929 (n6909, \a[23] , n_2110);
  and g8930 (n6910, n_2109, n_2110);
  not g8931 (n_2111, n6909);
  not g8932 (n_2112, n6910);
  and g8933 (n6911, n_2111, n_2112);
  not g8934 (n_2113, n6911);
  and g8935 (n6912, n6900, n_2113);
  not g8936 (n_2114, n6912);
  and g8937 (n6913, n_2103, n_2114);
  not g8938 (n_2115, n6465);
  not g8939 (n_2116, n6913);
  and g8940 (n6914, n_2115, n_2116);
  not g8941 (n_2117, n6914);
  and g8942 (n6915, n_1938, n_2117);
  not g8943 (n_2118, n6448);
  not g8944 (n_2119, n6915);
  and g8945 (n6916, n_2118, n_2119);
  and g8946 (n6917, n6448, n6915);
  not g8947 (n_2120, n6916);
  not g8948 (n_2121, n6917);
  and g8949 (n6918, n_2120, n_2121);
  and g8950 (n6919, n_415, n5496);
  and g8951 (n6920, n_237, n4935);
  and g8952 (n6921, n_236, n5407);
  and g8958 (n6924, n3018, n4938);
  not g8961 (n_2126, n6925);
  and g8962 (n6926, \a[20] , n_2126);
  not g8963 (n_2127, n6926);
  and g8964 (n6927, \a[20] , n_2127);
  and g8965 (n6928, n_2126, n_2127);
  not g8966 (n_2128, n6927);
  not g8967 (n_2129, n6928);
  and g8968 (n6929, n_2128, n_2129);
  not g8969 (n_2130, n6929);
  and g8970 (n6930, n6918, n_2130);
  not g8971 (n_2131, n6930);
  and g8972 (n6931, n_2120, n_2131);
  not g8973 (n_2132, n6445);
  not g8974 (n_2133, n6931);
  and g8975 (n6932, n_2132, n_2133);
  and g8976 (n6933, n6445, n6931);
  not g8977 (n_2134, n6932);
  not g8978 (n_2135, n6933);
  and g8979 (n6934, n_2134, n_2135);
  and g8980 (n6935, n_535, n6233);
  and g8981 (n6936, n_485, n5663);
  and g8982 (n6937, n_480, n5939);
  and g8988 (n6940, n3818, n5666);
  not g8991 (n_2140, n6941);
  and g8992 (n6942, \a[17] , n_2140);
  not g8993 (n_2141, n6942);
  and g8994 (n6943, \a[17] , n_2141);
  and g8995 (n6944, n_2140, n_2141);
  not g8996 (n_2142, n6943);
  not g8997 (n_2143, n6944);
  and g8998 (n6945, n_2142, n_2143);
  not g8999 (n_2144, n6945);
  and g9000 (n6946, n6934, n_2144);
  not g9001 (n_2145, n6946);
  and g9002 (n6947, n_2134, n_2145);
  not g9003 (n_2146, n6442);
  not g9004 (n_2147, n6947);
  and g9005 (n6948, n_2146, n_2147);
  not g9006 (n_2148, n6948);
  and g9007 (n6949, n_1920, n_2148);
  and g9008 (n6950, n_560, n6402);
  not g9009 (n_2149, n6400);
  and g9010 (n6951, n6393, n_2149);
  and g9011 (n6952, n_712, n6951);
  not g9012 (n_2150, n6950);
  not g9013 (n_2151, n6952);
  and g9014 (n6953, n_2150, n_2151);
  and g9015 (n6954, n_1885, n6953);
  not g9016 (n_2152, n4609);
  and g9017 (n6955, n_2152, n6953);
  not g9018 (n_2153, n6954);
  not g9019 (n_2154, n6955);
  and g9020 (n6956, n_2153, n_2154);
  not g9021 (n_2155, n6956);
  and g9022 (n6957, \a[14] , n_2155);
  and g9023 (n6958, n_652, n6956);
  not g9024 (n_2156, n6957);
  not g9025 (n_2157, n6958);
  and g9026 (n6959, n_2156, n_2157);
  not g9027 (n_2158, n6949);
  not g9028 (n_2159, n6959);
  and g9029 (n6960, n_2158, n_2159);
  and g9030 (n6961, n6377, n_1872);
  and g9031 (n6962, n_1871, n_1872);
  not g9032 (n_2160, n6961);
  not g9033 (n_2161, n6962);
  and g9034 (n6963, n_2160, n_2161);
  and g9035 (n6964, n6949, n6959);
  not g9036 (n_2162, n6960);
  not g9037 (n_2163, n6964);
  and g9038 (n6965, n_2162, n_2163);
  not g9039 (n_2164, n6963);
  and g9040 (n6966, n_2164, n6965);
  not g9041 (n_2165, n6966);
  and g9042 (n6967, n_2162, n_2165);
  not g9043 (n_2166, n6425);
  not g9044 (n_2167, n6967);
  and g9045 (n6968, n_2166, n_2167);
  and g9046 (n6969, n6425, n6967);
  not g9047 (n_2168, n6968);
  not g9048 (n_2169, n6969);
  and g9049 (n6970, n_2168, n_2169);
  and g9050 (n6971, n6934, n_2145);
  and g9051 (n6972, n_2144, n_2145);
  not g9052 (n_2170, n6971);
  not g9053 (n_2171, n6972);
  and g9054 (n6973, n_2170, n_2171);
  and g9055 (n6974, n6918, n_2131);
  and g9056 (n6975, n_2130, n_2131);
  not g9057 (n_2172, n6974);
  not g9058 (n_2173, n6975);
  and g9059 (n6976, n_2172, n_2173);
  and g9060 (n6977, n6465, n6913);
  not g9061 (n_2174, n6977);
  and g9062 (n6978, n_2117, n_2174);
  and g9063 (n6979, n_236, n5496);
  and g9064 (n6980, n_260, n4935);
  and g9065 (n6981, n_237, n5407);
  not g9066 (n_2175, n6980);
  not g9067 (n_2176, n6981);
  and g9068 (n6982, n_2175, n_2176);
  not g9069 (n_2177, n6979);
  and g9070 (n6983, n_2177, n6982);
  and g9071 (n6984, n_1011, n6983);
  and g9072 (n6985, n_1208, n6983);
  not g9073 (n_2178, n6984);
  not g9074 (n_2179, n6985);
  and g9075 (n6986, n_2178, n_2179);
  not g9076 (n_2180, n6986);
  and g9077 (n6987, \a[20] , n_2180);
  and g9078 (n6988, n_435, n6986);
  not g9079 (n_2181, n6987);
  not g9080 (n_2182, n6988);
  and g9081 (n6989, n_2181, n_2182);
  not g9082 (n_2183, n6989);
  and g9083 (n6990, n6978, n_2183);
  and g9084 (n6991, n6900, n_2114);
  and g9085 (n6992, n_2113, n_2114);
  not g9086 (n_2184, n6991);
  not g9087 (n_2185, n6992);
  and g9088 (n6993, n_2184, n_2185);
  and g9089 (n6994, n6884, n_2100);
  and g9090 (n6995, n_2099, n_2100);
  not g9091 (n_2186, n6994);
  not g9092 (n_2187, n6995);
  and g9093 (n6996, n_2186, n_2187);
  and g9094 (n6997, n6866, n_2084);
  and g9095 (n6998, n_2083, n_2084);
  not g9096 (n_2188, n6997);
  not g9097 (n_2189, n6998);
  and g9098 (n6999, n_2188, n_2189);
  and g9099 (n7000, n_299, n3884);
  and g9100 (n7001, n_301, n3967);
  and g9101 (n7002, n_300, n4046);
  not g9102 (n_2190, n7001);
  not g9103 (n_2191, n7002);
  and g9104 (n7003, n_2190, n_2191);
  not g9105 (n_2192, n7000);
  and g9106 (n7004, n_2192, n7003);
  and g9107 (n7005, n_750, n7004);
  not g9108 (n_2193, n5139);
  and g9109 (n7006, n_2193, n7004);
  not g9110 (n_2194, n7005);
  not g9111 (n_2195, n7006);
  and g9112 (n7007, n_2194, n_2195);
  not g9113 (n_2196, n7007);
  and g9114 (n7008, \a[26] , n_2196);
  and g9115 (n7009, n_33, n7007);
  not g9116 (n_2197, n7008);
  not g9117 (n_2198, n7009);
  and g9118 (n7010, n_2197, n_2198);
  not g9119 (n_2199, n6999);
  not g9120 (n_2200, n7010);
  and g9121 (n7011, n_2199, n_2200);
  and g9122 (n7012, n_2068, n_2070);
  and g9123 (n7013, n_2069, n_2070);
  not g9124 (n_2201, n7012);
  not g9125 (n_2202, n7013);
  and g9126 (n7014, n_2201, n_2202);
  and g9127 (n7015, n_303, n3457);
  and g9128 (n7016, n_305, n3542);
  and g9129 (n7017, n_304, n3606);
  not g9130 (n_2203, n7016);
  not g9131 (n_2204, n7017);
  and g9132 (n7018, n_2203, n_2204);
  not g9133 (n_2205, n7015);
  and g9134 (n7019, n_2205, n7018);
  and g9135 (n7020, n_489, n7019);
  not g9136 (n_2206, n6007);
  and g9137 (n7021, n_2206, n7019);
  not g9138 (n_2207, n7020);
  not g9139 (n_2208, n7021);
  and g9140 (n7022, n_2207, n_2208);
  not g9141 (n_2209, n7022);
  and g9142 (n7023, \a[29] , n_2209);
  and g9143 (n7024, n_15, n7022);
  not g9144 (n_2210, n7023);
  not g9145 (n_2211, n7024);
  and g9146 (n7025, n_2210, n_2211);
  not g9147 (n_2212, n7014);
  not g9148 (n_2213, n7025);
  and g9149 (n7026, n_2212, n_2213);
  and g9150 (n7027, n7014, n7025);
  not g9151 (n_2214, n7026);
  not g9152 (n_2215, n7027);
  and g9153 (n7028, n_2214, n_2215);
  and g9154 (n7029, n_300, n3884);
  and g9155 (n7030, n_302, n3967);
  and g9156 (n7031, n_301, n4046);
  and g9162 (n7034, n4050, n5561);
  not g9165 (n_2220, n7035);
  and g9166 (n7036, \a[26] , n_2220);
  not g9167 (n_2221, n7036);
  and g9168 (n7037, \a[26] , n_2221);
  and g9169 (n7038, n_2220, n_2221);
  not g9170 (n_2222, n7037);
  not g9171 (n_2223, n7038);
  and g9172 (n7039, n_2222, n_2223);
  not g9173 (n_2224, n7039);
  and g9174 (n7040, n7028, n_2224);
  not g9175 (n_2225, n7040);
  and g9176 (n7041, n_2214, n_2225);
  and g9177 (n7042, n6999, n7010);
  not g9178 (n_2226, n7011);
  not g9179 (n_2227, n7042);
  and g9180 (n7043, n_2226, n_2227);
  not g9181 (n_2228, n7041);
  and g9182 (n7044, n_2228, n7043);
  not g9183 (n_2229, n7044);
  and g9184 (n7045, n_2226, n_2229);
  not g9185 (n_2230, n6996);
  not g9186 (n_2231, n7045);
  and g9187 (n7046, n_2230, n_2231);
  and g9188 (n7047, n6996, n7045);
  not g9189 (n_2232, n7046);
  not g9190 (n_2233, n7047);
  and g9191 (n7048, n_2232, n_2233);
  and g9192 (n7049, n_286, n4694);
  and g9193 (n7050, n_295, n4533);
  and g9194 (n7051, n_293, n4604);
  and g9200 (n7054, n4429, n4536);
  not g9203 (n_2238, n7055);
  and g9204 (n7056, \a[23] , n_2238);
  not g9205 (n_2239, n7056);
  and g9206 (n7057, \a[23] , n_2239);
  and g9207 (n7058, n_2238, n_2239);
  not g9208 (n_2240, n7057);
  not g9209 (n_2241, n7058);
  and g9210 (n7059, n_2240, n_2241);
  not g9211 (n_2242, n7059);
  and g9212 (n7060, n7048, n_2242);
  not g9213 (n_2243, n7060);
  and g9214 (n7061, n_2232, n_2243);
  not g9215 (n_2244, n6993);
  not g9216 (n_2245, n7061);
  and g9217 (n7062, n_2244, n_2245);
  and g9218 (n7063, n6993, n7061);
  not g9219 (n_2246, n7062);
  not g9220 (n_2247, n7063);
  and g9221 (n7064, n_2246, n_2247);
  and g9222 (n7065, n_237, n5496);
  and g9223 (n7066, n_275, n4935);
  and g9224 (n7067, n_260, n5407);
  and g9230 (n7070, n3331, n4938);
  not g9233 (n_2252, n7071);
  and g9234 (n7072, \a[20] , n_2252);
  not g9235 (n_2253, n7072);
  and g9236 (n7073, \a[20] , n_2253);
  and g9237 (n7074, n_2252, n_2253);
  not g9238 (n_2254, n7073);
  not g9239 (n_2255, n7074);
  and g9240 (n7075, n_2254, n_2255);
  not g9241 (n_2256, n7075);
  and g9242 (n7076, n7064, n_2256);
  not g9243 (n_2257, n7076);
  and g9244 (n7077, n_2246, n_2257);
  not g9245 (n_2258, n6978);
  and g9246 (n7078, n_2258, n6989);
  not g9247 (n_2259, n6990);
  not g9248 (n_2260, n7078);
  and g9249 (n7079, n_2259, n_2260);
  not g9250 (n_2261, n7077);
  and g9251 (n7080, n_2261, n7079);
  not g9252 (n_2262, n7080);
  and g9253 (n7081, n_2259, n_2262);
  not g9254 (n_2263, n6976);
  not g9255 (n_2264, n7081);
  and g9256 (n7082, n_2263, n_2264);
  and g9257 (n7083, n6976, n7081);
  not g9258 (n_2265, n7082);
  not g9259 (n_2266, n7083);
  and g9260 (n7084, n_2265, n_2266);
  and g9261 (n7085, n_480, n6233);
  and g9262 (n7086, n_484, n5663);
  and g9263 (n7087, n_485, n5939);
  and g9269 (n7090, n3627, n5666);
  not g9272 (n_2271, n7091);
  and g9273 (n7092, \a[17] , n_2271);
  not g9274 (n_2272, n7092);
  and g9275 (n7093, \a[17] , n_2272);
  and g9276 (n7094, n_2271, n_2272);
  not g9277 (n_2273, n7093);
  not g9278 (n_2274, n7094);
  and g9279 (n7095, n_2273, n_2274);
  not g9280 (n_2275, n7095);
  and g9281 (n7096, n7084, n_2275);
  not g9282 (n_2276, n7096);
  and g9283 (n7097, n_2265, n_2276);
  not g9284 (n_2277, n6973);
  not g9285 (n_2278, n7097);
  and g9286 (n7098, n_2277, n_2278);
  and g9287 (n7099, n6973, n7097);
  not g9288 (n_2279, n7098);
  not g9289 (n_2280, n7099);
  and g9290 (n7100, n_2279, n_2280);
  and g9291 (n7101, n_1881, n6396);
  and g9292 (n7102, n_560, n7101);
  and g9293 (n7103, n_565, n6402);
  and g9294 (n7104, n_566, n6951);
  and g9300 (n7107, n4067, n6397);
  not g9303 (n_2285, n7108);
  and g9304 (n7109, \a[14] , n_2285);
  not g9305 (n_2286, n7109);
  and g9306 (n7110, \a[14] , n_2286);
  and g9307 (n7111, n_2285, n_2286);
  not g9308 (n_2287, n7110);
  not g9309 (n_2288, n7111);
  and g9310 (n7112, n_2287, n_2288);
  not g9311 (n_2289, n7112);
  and g9312 (n7113, n7100, n_2289);
  not g9313 (n_2290, n7113);
  and g9314 (n7114, n_2279, n_2290);
  and g9315 (n7115, n_712, n7101);
  and g9316 (n7116, n_566, n6402);
  and g9317 (n7117, n_560, n6951);
  not g9318 (n_2291, n7116);
  not g9319 (n_2292, n7117);
  and g9320 (n7118, n_2291, n_2292);
  not g9321 (n_2293, n7115);
  and g9322 (n7119, n_2293, n7118);
  and g9323 (n7120, n_1885, n7119);
  and g9324 (n7121, n_888, n7119);
  not g9325 (n_2294, n7120);
  not g9326 (n_2295, n7121);
  and g9327 (n7122, n_2294, n_2295);
  not g9328 (n_2296, n7122);
  and g9329 (n7123, \a[14] , n_2296);
  and g9330 (n7124, n_652, n7122);
  not g9331 (n_2297, n7123);
  not g9332 (n_2298, n7124);
  and g9333 (n7125, n_2297, n_2298);
  not g9334 (n_2299, n7114);
  not g9335 (n_2300, n7125);
  and g9336 (n7126, n_2299, n_2300);
  and g9337 (n7127, n6442, n6947);
  not g9338 (n_2301, n7127);
  and g9339 (n7128, n_2148, n_2301);
  not g9340 (n_2302, n7126);
  and g9341 (n7129, n_2299, n_2302);
  and g9342 (n7130, n_2300, n_2302);
  not g9343 (n_2303, n7129);
  not g9344 (n_2304, n7130);
  and g9345 (n7131, n_2303, n_2304);
  not g9346 (n_2305, n7131);
  and g9347 (n7132, n7128, n_2305);
  not g9348 (n_2306, n7132);
  and g9349 (n7133, n_2302, n_2306);
  not g9350 (n_2307, n6965);
  and g9351 (n7134, n6963, n_2307);
  not g9352 (n_2308, n7134);
  and g9353 (n7135, n_2165, n_2308);
  not g9354 (n_2309, n7133);
  and g9355 (n7136, n_2309, n7135);
  and g9356 (n7137, n7084, n_2276);
  and g9357 (n7138, n_2275, n_2276);
  not g9358 (n_2310, n7137);
  not g9359 (n_2311, n7138);
  and g9360 (n7139, n_2310, n_2311);
  and g9361 (n7140, n_485, n6233);
  and g9362 (n7141, n_415, n5663);
  and g9363 (n7142, n_484, n5939);
  and g9369 (n7145, n4084, n5666);
  not g9372 (n_2316, n7146);
  and g9373 (n7147, \a[17] , n_2316);
  not g9374 (n_2317, n7147);
  and g9375 (n7148, n_2316, n_2317);
  and g9376 (n7149, \a[17] , n_2317);
  not g9377 (n_2318, n7148);
  not g9378 (n_2319, n7149);
  and g9379 (n7150, n_2318, n_2319);
  not g9380 (n_2320, n7079);
  and g9381 (n7151, n7077, n_2320);
  not g9382 (n_2321, n7151);
  and g9383 (n7152, n_2262, n_2321);
  not g9384 (n_2322, n7150);
  and g9385 (n7153, n_2322, n7152);
  not g9386 (n_2323, n7153);
  and g9387 (n7154, n_2322, n_2323);
  and g9388 (n7155, n7152, n_2323);
  not g9389 (n_2324, n7154);
  not g9390 (n_2325, n7155);
  and g9391 (n7156, n_2324, n_2325);
  and g9392 (n7157, n7064, n_2257);
  and g9393 (n7158, n_2256, n_2257);
  not g9394 (n_2326, n7157);
  not g9395 (n_2327, n7158);
  and g9396 (n7159, n_2326, n_2327);
  and g9397 (n7160, n7048, n_2243);
  and g9398 (n7161, n_2242, n_2243);
  not g9399 (n_2328, n7160);
  not g9400 (n_2329, n7161);
  and g9401 (n7162, n_2328, n_2329);
  and g9402 (n7163, n_293, n4694);
  and g9403 (n7164, n_298, n4533);
  and g9404 (n7165, n_295, n4604);
  and g9410 (n7168, n4536, n4861);
  not g9413 (n_2334, n7169);
  and g9414 (n7170, \a[23] , n_2334);
  not g9415 (n_2335, n7170);
  and g9416 (n7171, n_2334, n_2335);
  and g9417 (n7172, \a[23] , n_2335);
  not g9418 (n_2336, n7171);
  not g9419 (n_2337, n7172);
  and g9420 (n7173, n_2336, n_2337);
  not g9421 (n_2338, n7043);
  and g9422 (n7174, n7041, n_2338);
  not g9423 (n_2339, n7174);
  and g9424 (n7175, n_2229, n_2339);
  not g9425 (n_2340, n7173);
  and g9426 (n7176, n_2340, n7175);
  not g9427 (n_2341, n7176);
  and g9428 (n7177, n_2340, n_2341);
  and g9429 (n7178, n7175, n_2341);
  not g9430 (n_2342, n7177);
  not g9431 (n_2343, n7178);
  and g9432 (n7179, n_2342, n_2343);
  and g9433 (n7180, n7028, n_2225);
  and g9434 (n7181, n_2224, n_2225);
  not g9435 (n_2344, n7180);
  not g9436 (n_2345, n7181);
  and g9437 (n7182, n_2344, n_2345);
  and g9438 (n7183, n_2062, n_2064);
  and g9439 (n7184, n_2063, n_2064);
  not g9440 (n_2346, n7183);
  not g9441 (n_2347, n7184);
  and g9442 (n7185, n_2346, n_2347);
  and g9443 (n7186, n_304, n3457);
  and g9444 (n7187, n_306, n3542);
  and g9445 (n7188, n_305, n3606);
  not g9446 (n_2348, n7187);
  not g9447 (n_2349, n7188);
  and g9448 (n7189, n_2348, n_2349);
  not g9449 (n_2350, n7186);
  and g9450 (n7190, n_2350, n7189);
  and g9451 (n7191, n_489, n7190);
  not g9452 (n_2351, n5834);
  and g9453 (n7192, n_2351, n7190);
  not g9454 (n_2352, n7191);
  not g9455 (n_2353, n7192);
  and g9456 (n7193, n_2352, n_2353);
  not g9457 (n_2354, n7193);
  and g9458 (n7194, \a[29] , n_2354);
  and g9459 (n7195, n_15, n7193);
  not g9460 (n_2355, n7194);
  not g9461 (n_2356, n7195);
  and g9462 (n7196, n_2355, n_2356);
  not g9463 (n_2357, n7185);
  not g9464 (n_2358, n7196);
  and g9465 (n7197, n_2357, n_2358);
  and g9466 (n7198, n7185, n7196);
  not g9467 (n_2359, n7197);
  not g9468 (n_2360, n7198);
  and g9469 (n7199, n_2359, n_2360);
  and g9470 (n7200, n_301, n3884);
  and g9471 (n7201, n_303, n3967);
  and g9472 (n7202, n_302, n4046);
  and g9478 (n7205, n4050, n5328);
  not g9481 (n_2365, n7206);
  and g9482 (n7207, \a[26] , n_2365);
  not g9483 (n_2366, n7207);
  and g9484 (n7208, \a[26] , n_2366);
  and g9485 (n7209, n_2365, n_2366);
  not g9486 (n_2367, n7208);
  not g9487 (n_2368, n7209);
  and g9488 (n7210, n_2367, n_2368);
  not g9489 (n_2369, n7210);
  and g9490 (n7211, n7199, n_2369);
  not g9491 (n_2370, n7211);
  and g9492 (n7212, n_2359, n_2370);
  not g9493 (n_2371, n7182);
  not g9494 (n_2372, n7212);
  and g9495 (n7213, n_2371, n_2372);
  and g9496 (n7214, n7182, n7212);
  not g9497 (n_2373, n7213);
  not g9498 (n_2374, n7214);
  and g9499 (n7215, n_2373, n_2374);
  and g9500 (n7216, n_295, n4694);
  and g9501 (n7217, n_299, n4533);
  and g9502 (n7218, n_298, n4604);
  and g9508 (n7221, n4536, n4848);
  not g9511 (n_2379, n7222);
  and g9512 (n7223, \a[23] , n_2379);
  not g9513 (n_2380, n7223);
  and g9514 (n7224, \a[23] , n_2380);
  and g9515 (n7225, n_2379, n_2380);
  not g9516 (n_2381, n7224);
  not g9517 (n_2382, n7225);
  and g9518 (n7226, n_2381, n_2382);
  not g9519 (n_2383, n7226);
  and g9520 (n7227, n7215, n_2383);
  not g9521 (n_2384, n7227);
  and g9522 (n7228, n_2373, n_2384);
  not g9523 (n_2385, n7179);
  not g9524 (n_2386, n7228);
  and g9525 (n7229, n_2385, n_2386);
  not g9526 (n_2387, n7229);
  and g9527 (n7230, n_2341, n_2387);
  not g9528 (n_2388, n7162);
  not g9529 (n_2389, n7230);
  and g9530 (n7231, n_2388, n_2389);
  and g9531 (n7232, n7162, n7230);
  not g9532 (n_2390, n7231);
  not g9533 (n_2391, n7232);
  and g9534 (n7233, n_2390, n_2391);
  and g9535 (n7234, n_260, n5496);
  and g9536 (n7235, n_281, n4935);
  and g9537 (n7236, n_275, n5407);
  and g9543 (n7239, n4179, n4938);
  not g9546 (n_2396, n7240);
  and g9547 (n7241, \a[20] , n_2396);
  not g9548 (n_2397, n7241);
  and g9549 (n7242, \a[20] , n_2397);
  and g9550 (n7243, n_2396, n_2397);
  not g9551 (n_2398, n7242);
  not g9552 (n_2399, n7243);
  and g9553 (n7244, n_2398, n_2399);
  not g9554 (n_2400, n7244);
  and g9555 (n7245, n7233, n_2400);
  not g9556 (n_2401, n7245);
  and g9557 (n7246, n_2390, n_2401);
  not g9558 (n_2402, n7159);
  not g9559 (n_2403, n7246);
  and g9560 (n7247, n_2402, n_2403);
  and g9561 (n7248, n7159, n7246);
  not g9562 (n_2404, n7247);
  not g9563 (n_2405, n7248);
  and g9564 (n7249, n_2404, n_2405);
  and g9565 (n7250, n_484, n6233);
  and g9566 (n7251, n_236, n5663);
  and g9567 (n7252, n_415, n5939);
  and g9573 (n7255, n3715, n5666);
  not g9576 (n_2410, n7256);
  and g9577 (n7257, \a[17] , n_2410);
  not g9578 (n_2411, n7257);
  and g9579 (n7258, \a[17] , n_2411);
  and g9580 (n7259, n_2410, n_2411);
  not g9581 (n_2412, n7258);
  not g9582 (n_2413, n7259);
  and g9583 (n7260, n_2412, n_2413);
  not g9584 (n_2414, n7260);
  and g9585 (n7261, n7249, n_2414);
  not g9586 (n_2415, n7261);
  and g9587 (n7262, n_2404, n_2415);
  not g9588 (n_2416, n7156);
  not g9589 (n_2417, n7262);
  and g9590 (n7263, n_2416, n_2417);
  not g9591 (n_2418, n7263);
  and g9592 (n7264, n_2323, n_2418);
  not g9593 (n_2419, n7139);
  not g9594 (n_2420, n7264);
  and g9595 (n7265, n_2419, n_2420);
  and g9596 (n7266, n7139, n7264);
  not g9597 (n_2421, n7265);
  not g9598 (n_2422, n7266);
  and g9599 (n7267, n_2421, n_2422);
  and g9600 (n7268, n_566, n7101);
  and g9601 (n7269, n_535, n6402);
  and g9602 (n7270, n_565, n6951);
  and g9608 (n7273, n4477, n6397);
  not g9611 (n_2427, n7274);
  and g9612 (n7275, \a[14] , n_2427);
  not g9613 (n_2428, n7275);
  and g9614 (n7276, \a[14] , n_2428);
  and g9615 (n7277, n_2427, n_2428);
  not g9616 (n_2429, n7276);
  not g9617 (n_2430, n7277);
  and g9618 (n7278, n_2429, n_2430);
  not g9619 (n_2431, n7278);
  and g9620 (n7279, n7267, n_2431);
  not g9621 (n_2432, n7279);
  and g9622 (n7280, n_2421, n_2432);
  not g9623 (n_2434, \a[9] );
  and g9624 (n7281, n_2434, \a[10] );
  not g9625 (n_2436, \a[10] );
  and g9626 (n7282, \a[9] , n_2436);
  not g9627 (n_2437, n7281);
  not g9628 (n_2438, n7282);
  and g9629 (n7283, n_2437, n_2438);
  and g9630 (n7284, \a[10] , n_1071);
  and g9631 (n7285, n_2436, \a[11] );
  not g9632 (n_2439, n7284);
  not g9633 (n_2440, n7285);
  and g9634 (n7286, n_2439, n_2440);
  and g9635 (n7287, \a[8] , n_2434);
  and g9636 (n7288, n_1106, \a[9] );
  not g9637 (n_2441, n7287);
  not g9638 (n_2442, n7288);
  and g9639 (n7289, n_2441, n_2442);
  not g9640 (n_2443, n7286);
  and g9641 (n7290, n_2443, n7289);
  and g9642 (n7291, n7283, n7290);
  and g9643 (n7292, n_712, n7291);
  not g9644 (n_2444, n7292);
  and g9645 (n7293, n_729, n_2444);
  not g9646 (n_2445, n7289);
  and g9647 (n7294, n_2443, n_2445);
  not g9648 (n_2446, n7294);
  and g9649 (n7295, n_2444, n_2446);
  not g9650 (n_2447, n7293);
  not g9651 (n_2448, n7295);
  and g9652 (n7296, n_2447, n_2448);
  not g9653 (n_2449, n7296);
  and g9654 (n7297, \a[11] , n_2449);
  and g9655 (n7298, n_1071, n7296);
  not g9656 (n_2450, n7297);
  not g9657 (n_2451, n7298);
  and g9658 (n7299, n_2450, n_2451);
  not g9659 (n_2452, n7280);
  not g9660 (n_2453, n7299);
  and g9661 (n7300, n_2452, n_2453);
  and g9662 (n7301, n7100, n_2290);
  and g9663 (n7302, n_2289, n_2290);
  not g9664 (n_2454, n7301);
  not g9665 (n_2455, n7302);
  and g9666 (n7303, n_2454, n_2455);
  and g9667 (n7304, n7280, n7299);
  not g9668 (n_2456, n7300);
  not g9669 (n_2457, n7304);
  and g9670 (n7305, n_2456, n_2457);
  not g9671 (n_2458, n7303);
  and g9672 (n7306, n_2458, n7305);
  not g9673 (n_2459, n7306);
  and g9674 (n7307, n_2456, n_2459);
  not g9675 (n_2460, n7128);
  and g9676 (n7308, n_2460, n_2304);
  and g9677 (n7309, n_2303, n7308);
  not g9678 (n_2461, n7309);
  and g9679 (n7310, n_2306, n_2461);
  not g9680 (n_2462, n7307);
  and g9681 (n7311, n_2462, n7310);
  and g9682 (n7312, n_2458, n_2459);
  and g9683 (n7313, n7305, n_2459);
  not g9684 (n_2463, n7312);
  not g9685 (n_2464, n7313);
  and g9686 (n7314, n_2463, n_2464);
  and g9687 (n7315, n7156, n7262);
  not g9688 (n_2465, n7315);
  and g9689 (n7316, n_2418, n_2465);
  and g9690 (n7317, n_565, n7101);
  and g9691 (n7318, n_480, n6402);
  and g9692 (n7319, n_535, n6951);
  not g9693 (n_2466, n7318);
  not g9694 (n_2467, n7319);
  and g9695 (n7320, n_2466, n_2467);
  not g9696 (n_2468, n7317);
  and g9697 (n7321, n_2468, n7320);
  and g9698 (n7322, n_1885, n7321);
  and g9699 (n7323, n_753, n7321);
  not g9700 (n_2469, n7322);
  not g9701 (n_2470, n7323);
  and g9702 (n7324, n_2469, n_2470);
  not g9703 (n_2471, n7324);
  and g9704 (n7325, \a[14] , n_2471);
  and g9705 (n7326, n_652, n7324);
  not g9706 (n_2472, n7325);
  not g9707 (n_2473, n7326);
  and g9708 (n7327, n_2472, n_2473);
  not g9709 (n_2474, n7327);
  and g9710 (n7328, n7316, n_2474);
  and g9711 (n7329, n7249, n_2415);
  and g9712 (n7330, n_2414, n_2415);
  not g9713 (n_2475, n7329);
  not g9714 (n_2476, n7330);
  and g9715 (n7331, n_2475, n_2476);
  and g9716 (n7332, n7233, n_2401);
  and g9717 (n7333, n_2400, n_2401);
  not g9718 (n_2477, n7332);
  not g9719 (n_2478, n7333);
  and g9720 (n7334, n_2477, n_2478);
  and g9721 (n7335, n7179, n7228);
  not g9722 (n_2479, n7335);
  and g9723 (n7336, n_2387, n_2479);
  and g9724 (n7337, n_275, n5496);
  and g9725 (n7338, n_286, n4935);
  and g9726 (n7339, n_281, n5407);
  not g9727 (n_2480, n7338);
  not g9728 (n_2481, n7339);
  and g9729 (n7340, n_2480, n_2481);
  not g9730 (n_2482, n7337);
  and g9731 (n7341, n_2482, n7340);
  and g9732 (n7342, n_1011, n7341);
  and g9733 (n7343, n_1450, n7341);
  not g9734 (n_2483, n7342);
  not g9735 (n_2484, n7343);
  and g9736 (n7344, n_2483, n_2484);
  not g9737 (n_2485, n7344);
  and g9738 (n7345, \a[20] , n_2485);
  and g9739 (n7346, n_435, n7344);
  not g9740 (n_2486, n7345);
  not g9741 (n_2487, n7346);
  and g9742 (n7347, n_2486, n_2487);
  not g9743 (n_2488, n7347);
  and g9744 (n7348, n7336, n_2488);
  and g9745 (n7349, n7215, n_2384);
  and g9746 (n7350, n_2383, n_2384);
  not g9747 (n_2489, n7349);
  not g9748 (n_2490, n7350);
  and g9749 (n7351, n_2489, n_2490);
  and g9750 (n7352, n7199, n_2370);
  and g9751 (n7353, n_2369, n_2370);
  not g9752 (n_2491, n7352);
  not g9753 (n_2492, n7353);
  and g9754 (n7354, n_2491, n_2492);
  and g9755 (n7355, n_2041, n_2043);
  and g9756 (n7356, n_2042, n_2043);
  not g9757 (n_2493, n7355);
  not g9758 (n_2494, n7356);
  and g9759 (n7357, n_2493, n_2494);
  and g9760 (n7358, n_306, n3457);
  and g9761 (n7359, n_308, n3542);
  and g9762 (n7360, n_307, n3606);
  not g9763 (n_2495, n7359);
  not g9764 (n_2496, n7360);
  and g9765 (n7361, n_2495, n_2496);
  not g9766 (n_2497, n7358);
  and g9767 (n7362, n_2497, n7361);
  and g9768 (n7363, n_489, n7362);
  not g9769 (n_2498, n6479);
  and g9770 (n7364, n_2498, n7362);
  not g9771 (n_2499, n7363);
  not g9772 (n_2500, n7364);
  and g9773 (n7365, n_2499, n_2500);
  not g9774 (n_2501, n7365);
  and g9775 (n7366, \a[29] , n_2501);
  and g9776 (n7367, n_15, n7365);
  not g9777 (n_2502, n7366);
  not g9778 (n_2503, n7367);
  and g9779 (n7368, n_2502, n_2503);
  not g9780 (n_2504, n7357);
  not g9781 (n_2505, n7368);
  and g9782 (n7369, n_2504, n_2505);
  and g9783 (n7370, n_2035, n_2037);
  and g9784 (n7371, n_2036, n_2037);
  not g9785 (n_2506, n7370);
  not g9786 (n_2507, n7371);
  and g9787 (n7372, n_2506, n_2507);
  and g9788 (n7373, n_307, n3457);
  and g9789 (n7374, n_309, n3542);
  and g9790 (n7375, n_308, n3606);
  not g9791 (n_2508, n7374);
  not g9792 (n_2509, n7375);
  and g9793 (n7376, n_2508, n_2509);
  not g9794 (n_2510, n7373);
  and g9795 (n7377, n_2510, n7376);
  and g9796 (n7378, n_489, n7377);
  not g9797 (n_2511, n6492);
  and g9798 (n7379, n_2511, n7377);
  not g9799 (n_2512, n7378);
  not g9800 (n_2513, n7379);
  and g9801 (n7380, n_2512, n_2513);
  not g9802 (n_2514, n7380);
  and g9803 (n7381, \a[29] , n_2514);
  and g9804 (n7382, n_15, n7380);
  not g9805 (n_2515, n7381);
  not g9806 (n_2516, n7382);
  and g9807 (n7383, n_2515, n_2516);
  not g9808 (n_2517, n7372);
  not g9809 (n_2518, n7383);
  and g9810 (n7384, n_2517, n_2518);
  and g9811 (n7385, n_308, n3457);
  and g9812 (n7386, n_310, n3542);
  and g9813 (n7387, n_309, n3606);
  and g9819 (n7390, n3368, n6122);
  not g9822 (n_2523, n7391);
  and g9823 (n7392, \a[29] , n_2523);
  not g9824 (n_2524, n7392);
  and g9825 (n7393, n_2523, n_2524);
  and g9826 (n7394, \a[29] , n_2524);
  not g9827 (n_2525, n7393);
  not g9828 (n_2526, n7394);
  and g9829 (n7395, n_2525, n_2526);
  and g9830 (n7396, n_2029, n_2031);
  and g9831 (n7397, n_2030, n_2031);
  not g9832 (n_2527, n7396);
  not g9833 (n_2528, n7397);
  and g9834 (n7398, n_2527, n_2528);
  not g9835 (n_2529, n7395);
  not g9836 (n_2530, n7398);
  and g9837 (n7399, n_2529, n_2530);
  not g9838 (n_2531, n7399);
  and g9839 (n7400, n_2529, n_2531);
  and g9840 (n7401, n_2530, n_2531);
  not g9841 (n_2532, n7400);
  not g9842 (n_2533, n7401);
  and g9843 (n7402, n_2532, n_2533);
  and g9844 (n7403, n_309, n3457);
  and g9845 (n7404, n_311, n3542);
  and g9846 (n7405, n_310, n3606);
  and g9852 (n7408, n3368, n6541);
  not g9855 (n_2538, n7409);
  and g9856 (n7410, \a[29] , n_2538);
  not g9857 (n_2539, n7410);
  and g9858 (n7411, n_2538, n_2539);
  and g9859 (n7412, \a[29] , n_2539);
  not g9860 (n_2540, n7411);
  not g9861 (n_2541, n7412);
  and g9862 (n7413, n_2540, n_2541);
  and g9863 (n7414, n_2023, n_2025);
  and g9864 (n7415, n_2024, n_2025);
  not g9865 (n_2542, n7414);
  not g9866 (n_2543, n7415);
  and g9867 (n7416, n_2542, n_2543);
  not g9868 (n_2544, n7413);
  not g9869 (n_2545, n7416);
  and g9870 (n7417, n_2544, n_2545);
  not g9871 (n_2546, n7417);
  and g9872 (n7418, n_2544, n_2546);
  and g9873 (n7419, n_2545, n_2546);
  not g9874 (n_2547, n7418);
  not g9875 (n_2548, n7419);
  and g9876 (n7420, n_2547, n_2548);
  and g9877 (n7421, n_310, n3457);
  and g9878 (n7422, n_312, n3542);
  and g9879 (n7423, n_311, n3606);
  and g9885 (n7426, n3368, n6591);
  not g9888 (n_2553, n7427);
  and g9889 (n7428, \a[29] , n_2553);
  not g9890 (n_2554, n7428);
  and g9891 (n7429, n_2553, n_2554);
  and g9892 (n7430, \a[29] , n_2554);
  not g9893 (n_2555, n7429);
  not g9894 (n_2556, n7430);
  and g9895 (n7431, n_2555, n_2556);
  and g9896 (n7432, n_2018, n_2019);
  and g9897 (n7433, n6815, n_2019);
  not g9898 (n_2557, n7432);
  not g9899 (n_2558, n7433);
  and g9900 (n7434, n_2557, n_2558);
  not g9901 (n_2559, n7431);
  not g9902 (n_2560, n7434);
  and g9903 (n7435, n_2559, n_2560);
  not g9904 (n_2561, n7435);
  and g9905 (n7436, n_2559, n_2561);
  and g9906 (n7437, n_2560, n_2561);
  not g9907 (n_2562, n7436);
  not g9908 (n_2563, n7437);
  and g9909 (n7438, n_2562, n_2563);
  and g9910 (n7439, n_311, n3457);
  and g9911 (n7440, n_313, n3542);
  and g9912 (n7441, n_312, n3606);
  and g9918 (n7444, n3368, n6646);
  not g9921 (n_2568, n7445);
  and g9922 (n7446, \a[29] , n_2568);
  not g9923 (n_2569, n7446);
  and g9924 (n7447, n_2568, n_2569);
  and g9925 (n7448, \a[29] , n_2569);
  not g9926 (n_2570, n7447);
  not g9927 (n_2571, n7448);
  and g9928 (n7449, n_2570, n_2571);
  and g9929 (n7450, n_2006, n_2015);
  and g9930 (n7451, n_2007, n_2015);
  not g9931 (n_2572, n7450);
  not g9932 (n_2573, n7451);
  and g9933 (n7452, n_2572, n_2573);
  not g9934 (n_2574, n7449);
  not g9935 (n_2575, n7452);
  and g9936 (n7453, n_2574, n_2575);
  not g9937 (n_2576, n7453);
  and g9938 (n7454, n_2574, n_2576);
  and g9939 (n7455, n_2575, n_2576);
  not g9940 (n_2577, n7454);
  not g9941 (n_2578, n7455);
  and g9942 (n7456, n_2577, n_2578);
  and g9943 (n7457, n_312, n3457);
  and g9944 (n7458, n_314, n3542);
  and g9945 (n7459, n_313, n3606);
  and g9951 (n7462, n3368, n6695);
  not g9954 (n_2583, n7463);
  and g9955 (n7464, \a[29] , n_2583);
  not g9956 (n_2584, n7464);
  and g9957 (n7465, n_2583, n_2584);
  and g9958 (n7466, \a[29] , n_2584);
  not g9959 (n_2585, n7465);
  not g9960 (n_2586, n7466);
  and g9961 (n7467, n_2585, n_2586);
  and g9962 (n7468, n2736, n_316);
  not g9963 (n_2587, n7468);
  and g9964 (n7469, n_1999, n_2587);
  not g9965 (n_2588, n7469);
  and g9966 (n7470, n75, n_2588);
  and g9967 (n7471, n_316, n3028);
  and g9968 (n7472, n_315, n3020);
  not g9969 (n_2589, n7471);
  not g9970 (n_2590, n7472);
  and g9971 (n7473, n_2589, n_2590);
  not g9972 (n_2591, n7470);
  and g9973 (n7474, n_2591, n7473);
  not g9974 (n_2592, n7467);
  not g9975 (n_2593, n7474);
  and g9976 (n7475, n_2592, n_2593);
  not g9977 (n_2594, n7475);
  and g9978 (n7476, n_2592, n_2594);
  and g9979 (n7477, n_2593, n_2594);
  not g9980 (n_2595, n7476);
  not g9981 (n_2596, n7477);
  and g9982 (n7478, n_2595, n_2596);
  not g9983 (n_2597, n75);
  not g9984 (n_2598, n3020);
  and g9985 (n7479, n_2597, n_2598);
  not g9986 (n_2599, n7479);
  and g9987 (n7480, n_316, n_2599);
  and g9988 (n7481, n_316, n3606);
  and g9989 (n7482, n_315, n3457);
  not g9990 (n_2600, n7481);
  not g9991 (n_2601, n7482);
  and g9992 (n7483, n_2600, n_2601);
  and g9993 (n7484, n3368, n_2588);
  not g9994 (n_2602, n7484);
  and g9995 (n7485, n7483, n_2602);
  not g9996 (n_2603, n7485);
  and g9997 (n7486, \a[29] , n_2603);
  not g9998 (n_2604, n7486);
  and g9999 (n7487, \a[29] , n_2604);
  and g10000 (n7488, n_2603, n_2604);
  not g10001 (n_2605, n7487);
  not g10002 (n_2606, n7488);
  and g10003 (n7489, n_2605, n_2606);
  and g10004 (n7490, n_316, n_479);
  not g10005 (n_2607, n7490);
  and g10006 (n7491, \a[29] , n_2607);
  not g10007 (n_2608, n7489);
  and g10008 (n7492, n_2608, n7491);
  and g10009 (n7493, n_314, n3457);
  and g10010 (n7494, n_316, n3542);
  and g10011 (n7495, n_315, n3606);
  not g10012 (n_2609, n7494);
  not g10013 (n_2610, n7495);
  and g10014 (n7496, n_2609, n_2610);
  not g10015 (n_2611, n7493);
  and g10016 (n7497, n_2611, n7496);
  and g10017 (n7498, n_489, n7497);
  not g10018 (n_2612, n6798);
  and g10019 (n7499, n_2612, n7497);
  not g10020 (n_2613, n7498);
  not g10021 (n_2614, n7499);
  and g10022 (n7500, n_2613, n_2614);
  not g10023 (n_2615, n7500);
  and g10024 (n7501, \a[29] , n_2615);
  and g10025 (n7502, n_15, n7500);
  not g10026 (n_2616, n7501);
  not g10027 (n_2617, n7502);
  and g10028 (n7503, n_2616, n_2617);
  not g10029 (n_2618, n7503);
  and g10030 (n7504, n7492, n_2618);
  and g10031 (n7505, n7480, n7504);
  and g10032 (n7506, n_313, n3457);
  and g10033 (n7507, n_315, n3542);
  and g10034 (n7508, n_314, n3606);
  and g10040 (n7511, n3368, n6806);
  not g10043 (n_2623, n7512);
  and g10044 (n7513, \a[29] , n_2623);
  not g10045 (n_2624, n7513);
  and g10046 (n7514, n_2623, n_2624);
  and g10047 (n7515, \a[29] , n_2624);
  not g10048 (n_2625, n7514);
  not g10049 (n_2626, n7515);
  and g10050 (n7516, n_2625, n_2626);
  not g10051 (n_2627, n7480);
  and g10052 (n7517, n_2627, n7504);
  not g10053 (n_2628, n7504);
  and g10054 (n7518, n7480, n_2628);
  not g10055 (n_2629, n7517);
  not g10056 (n_2630, n7518);
  and g10057 (n7519, n_2629, n_2630);
  not g10058 (n_2631, n7516);
  not g10059 (n_2632, n7519);
  and g10060 (n7520, n_2631, n_2632);
  not g10061 (n_2633, n7505);
  not g10062 (n_2634, n7520);
  and g10063 (n7521, n_2633, n_2634);
  not g10064 (n_2635, n7478);
  not g10065 (n_2636, n7521);
  and g10066 (n7522, n_2635, n_2636);
  not g10067 (n_2637, n7522);
  and g10068 (n7523, n_2594, n_2637);
  not g10069 (n_2638, n7456);
  not g10070 (n_2639, n7523);
  and g10071 (n7524, n_2638, n_2639);
  not g10072 (n_2640, n7524);
  and g10073 (n7525, n_2576, n_2640);
  not g10074 (n_2641, n7438);
  not g10075 (n_2642, n7525);
  and g10076 (n7526, n_2641, n_2642);
  not g10077 (n_2643, n7526);
  and g10078 (n7527, n_2561, n_2643);
  not g10079 (n_2644, n7420);
  not g10080 (n_2645, n7527);
  and g10081 (n7528, n_2644, n_2645);
  not g10082 (n_2646, n7528);
  and g10083 (n7529, n_2546, n_2646);
  not g10084 (n_2647, n7402);
  not g10085 (n_2648, n7529);
  and g10086 (n7530, n_2647, n_2648);
  not g10087 (n_2649, n7530);
  and g10088 (n7531, n_2531, n_2649);
  and g10089 (n7532, n7372, n7383);
  not g10090 (n_2650, n7384);
  not g10091 (n_2651, n7532);
  and g10092 (n7533, n_2650, n_2651);
  not g10093 (n_2652, n7531);
  and g10094 (n7534, n_2652, n7533);
  not g10095 (n_2653, n7534);
  and g10096 (n7535, n_2650, n_2653);
  and g10097 (n7536, n7357, n7368);
  not g10098 (n_2654, n7369);
  not g10099 (n_2655, n7536);
  and g10100 (n7537, n_2654, n_2655);
  not g10101 (n_2656, n7535);
  and g10102 (n7538, n_2656, n7537);
  not g10103 (n_2657, n7538);
  and g10104 (n7539, n_2654, n_2657);
  not g10105 (n_2658, n6840);
  and g10106 (n7540, n_2658, n6851);
  not g10107 (n_2659, n7540);
  and g10108 (n7541, n_2058, n_2659);
  not g10109 (n_2660, n7539);
  and g10110 (n7542, n_2660, n7541);
  and g10111 (n7543, n_302, n3884);
  and g10112 (n7544, n_304, n3967);
  and g10113 (n7545, n_303, n4046);
  and g10119 (n7548, n4050, n5851);
  not g10122 (n_2665, n7549);
  and g10123 (n7550, \a[26] , n_2665);
  not g10124 (n_2666, n7550);
  and g10125 (n7551, n_2665, n_2666);
  and g10126 (n7552, \a[26] , n_2666);
  not g10127 (n_2667, n7551);
  not g10128 (n_2668, n7552);
  and g10129 (n7553, n_2667, n_2668);
  not g10130 (n_2669, n7541);
  and g10131 (n7554, n7539, n_2669);
  not g10132 (n_2670, n7542);
  not g10133 (n_2671, n7554);
  and g10134 (n7555, n_2670, n_2671);
  not g10135 (n_2672, n7553);
  and g10136 (n7556, n_2672, n7555);
  not g10137 (n_2673, n7556);
  and g10138 (n7557, n_2670, n_2673);
  not g10139 (n_2674, n7354);
  not g10140 (n_2675, n7557);
  and g10141 (n7558, n_2674, n_2675);
  and g10142 (n7559, n7354, n7557);
  not g10143 (n_2676, n7558);
  not g10144 (n_2677, n7559);
  and g10145 (n7560, n_2676, n_2677);
  and g10146 (n7561, n_298, n4694);
  and g10147 (n7562, n_300, n4533);
  and g10148 (n7563, n_299, n4604);
  and g10154 (n7566, n4536, n5114);
  not g10157 (n_2682, n7567);
  and g10158 (n7568, \a[23] , n_2682);
  not g10159 (n_2683, n7568);
  and g10160 (n7569, \a[23] , n_2683);
  and g10161 (n7570, n_2682, n_2683);
  not g10162 (n_2684, n7569);
  not g10163 (n_2685, n7570);
  and g10164 (n7571, n_2684, n_2685);
  not g10165 (n_2686, n7571);
  and g10166 (n7572, n7560, n_2686);
  not g10167 (n_2687, n7572);
  and g10168 (n7573, n_2676, n_2687);
  not g10169 (n_2688, n7351);
  not g10170 (n_2689, n7573);
  and g10171 (n7574, n_2688, n_2689);
  and g10172 (n7575, n7351, n7573);
  not g10173 (n_2690, n7574);
  not g10174 (n_2691, n7575);
  and g10175 (n7576, n_2690, n_2691);
  and g10176 (n7577, n_281, n5496);
  and g10177 (n7578, n_293, n4935);
  and g10178 (n7579, n_286, n5407);
  and g10184 (n7582, n4633, n4938);
  not g10187 (n_2696, n7583);
  and g10188 (n7584, \a[20] , n_2696);
  not g10189 (n_2697, n7584);
  and g10190 (n7585, \a[20] , n_2697);
  and g10191 (n7586, n_2696, n_2697);
  not g10192 (n_2698, n7585);
  not g10193 (n_2699, n7586);
  and g10194 (n7587, n_2698, n_2699);
  not g10195 (n_2700, n7587);
  and g10196 (n7588, n7576, n_2700);
  not g10197 (n_2701, n7588);
  and g10198 (n7589, n_2690, n_2701);
  not g10199 (n_2702, n7336);
  and g10200 (n7590, n_2702, n7347);
  not g10201 (n_2703, n7348);
  not g10202 (n_2704, n7590);
  and g10203 (n7591, n_2703, n_2704);
  not g10204 (n_2705, n7589);
  and g10205 (n7592, n_2705, n7591);
  not g10206 (n_2706, n7592);
  and g10207 (n7593, n_2703, n_2706);
  not g10208 (n_2707, n7334);
  not g10209 (n_2708, n7593);
  and g10210 (n7594, n_2707, n_2708);
  and g10211 (n7595, n7334, n7593);
  not g10212 (n_2709, n7594);
  not g10213 (n_2710, n7595);
  and g10214 (n7596, n_2709, n_2710);
  and g10215 (n7597, n_415, n6233);
  and g10216 (n7598, n_237, n5663);
  and g10217 (n7599, n_236, n5939);
  and g10223 (n7602, n3018, n5666);
  not g10226 (n_2715, n7603);
  and g10227 (n7604, \a[17] , n_2715);
  not g10228 (n_2716, n7604);
  and g10229 (n7605, \a[17] , n_2716);
  and g10230 (n7606, n_2715, n_2716);
  not g10231 (n_2717, n7605);
  not g10232 (n_2718, n7606);
  and g10233 (n7607, n_2717, n_2718);
  not g10234 (n_2719, n7607);
  and g10235 (n7608, n7596, n_2719);
  not g10236 (n_2720, n7608);
  and g10237 (n7609, n_2709, n_2720);
  not g10238 (n_2721, n7331);
  not g10239 (n_2722, n7609);
  and g10240 (n7610, n_2721, n_2722);
  and g10241 (n7611, n7331, n7609);
  not g10242 (n_2723, n7610);
  not g10243 (n_2724, n7611);
  and g10244 (n7612, n_2723, n_2724);
  and g10245 (n7613, n_535, n7101);
  and g10246 (n7614, n_485, n6402);
  and g10247 (n7615, n_480, n6951);
  and g10253 (n7618, n3818, n6397);
  not g10256 (n_2729, n7619);
  and g10257 (n7620, \a[14] , n_2729);
  not g10258 (n_2730, n7620);
  and g10259 (n7621, \a[14] , n_2730);
  and g10260 (n7622, n_2729, n_2730);
  not g10261 (n_2731, n7621);
  not g10262 (n_2732, n7622);
  and g10263 (n7623, n_2731, n_2732);
  not g10264 (n_2733, n7623);
  and g10265 (n7624, n7612, n_2733);
  not g10266 (n_2734, n7624);
  and g10267 (n7625, n_2723, n_2734);
  not g10268 (n_2735, n7328);
  and g10269 (n7626, n7316, n_2735);
  and g10270 (n7627, n_2474, n_2735);
  not g10271 (n_2736, n7626);
  not g10272 (n_2737, n7627);
  and g10273 (n7628, n_2736, n_2737);
  not g10274 (n_2738, n7625);
  not g10275 (n_2739, n7628);
  and g10276 (n7629, n_2738, n_2739);
  not g10277 (n_2740, n7629);
  and g10278 (n7630, n_2735, n_2740);
  and g10279 (n7631, n_560, n7291);
  not g10280 (n_2741, n7283);
  and g10281 (n7632, n_2741, n7289);
  and g10282 (n7633, n_712, n7632);
  not g10283 (n_2742, n7631);
  not g10284 (n_2743, n7633);
  and g10285 (n7634, n_2742, n_2743);
  and g10286 (n7635, n_2446, n7634);
  and g10287 (n7636, n_2152, n7634);
  not g10288 (n_2744, n7635);
  not g10289 (n_2745, n7636);
  and g10290 (n7637, n_2744, n_2745);
  not g10291 (n_2746, n7637);
  and g10292 (n7638, \a[11] , n_2746);
  and g10293 (n7639, n_1071, n7637);
  not g10294 (n_2747, n7638);
  not g10295 (n_2748, n7639);
  and g10296 (n7640, n_2747, n_2748);
  not g10297 (n_2749, n7630);
  not g10298 (n_2750, n7640);
  and g10299 (n7641, n_2749, n_2750);
  and g10300 (n7642, n7267, n_2432);
  and g10301 (n7643, n_2431, n_2432);
  not g10302 (n_2751, n7642);
  not g10303 (n_2752, n7643);
  and g10304 (n7644, n_2751, n_2752);
  and g10305 (n7645, n7630, n7640);
  not g10306 (n_2753, n7641);
  not g10307 (n_2754, n7645);
  and g10308 (n7646, n_2753, n_2754);
  not g10309 (n_2755, n7644);
  and g10310 (n7647, n_2755, n7646);
  not g10311 (n_2756, n7647);
  and g10312 (n7648, n_2753, n_2756);
  not g10313 (n_2757, n7314);
  not g10314 (n_2758, n7648);
  and g10315 (n7649, n_2757, n_2758);
  and g10316 (n7650, n7314, n7648);
  not g10317 (n_2759, n7649);
  not g10318 (n_2760, n7650);
  and g10319 (n7651, n_2759, n_2760);
  and g10320 (n7652, n7612, n_2734);
  and g10321 (n7653, n_2733, n_2734);
  not g10322 (n_2761, n7652);
  not g10323 (n_2762, n7653);
  and g10324 (n7654, n_2761, n_2762);
  and g10325 (n7655, n7596, n_2720);
  and g10326 (n7656, n_2719, n_2720);
  not g10327 (n_2763, n7655);
  not g10328 (n_2764, n7656);
  and g10329 (n7657, n_2763, n_2764);
  and g10330 (n7658, n_236, n6233);
  and g10331 (n7659, n_260, n5663);
  and g10332 (n7660, n_237, n5939);
  and g10338 (n7663, n3347, n5666);
  not g10341 (n_2769, n7664);
  and g10342 (n7665, \a[17] , n_2769);
  not g10343 (n_2770, n7665);
  and g10344 (n7666, n_2769, n_2770);
  and g10345 (n7667, \a[17] , n_2770);
  not g10346 (n_2771, n7666);
  not g10347 (n_2772, n7667);
  and g10348 (n7668, n_2771, n_2772);
  not g10349 (n_2773, n7591);
  and g10350 (n7669, n7589, n_2773);
  not g10351 (n_2774, n7669);
  and g10352 (n7670, n_2706, n_2774);
  not g10353 (n_2775, n7668);
  and g10354 (n7671, n_2775, n7670);
  not g10355 (n_2776, n7671);
  and g10356 (n7672, n_2775, n_2776);
  and g10357 (n7673, n7670, n_2776);
  not g10358 (n_2777, n7672);
  not g10359 (n_2778, n7673);
  and g10360 (n7674, n_2777, n_2778);
  and g10361 (n7675, n7576, n_2701);
  and g10362 (n7676, n_2700, n_2701);
  not g10363 (n_2779, n7675);
  not g10364 (n_2780, n7676);
  and g10365 (n7677, n_2779, n_2780);
  and g10366 (n7678, n7560, n_2687);
  and g10367 (n7679, n_2686, n_2687);
  not g10368 (n_2781, n7678);
  not g10369 (n_2782, n7679);
  and g10370 (n7680, n_2781, n_2782);
  not g10371 (n_2783, n7537);
  and g10372 (n7681, n7535, n_2783);
  not g10373 (n_2784, n7681);
  and g10374 (n7682, n_2657, n_2784);
  and g10375 (n7683, n_303, n3884);
  and g10376 (n7684, n_305, n3967);
  and g10377 (n7685, n_304, n4046);
  not g10378 (n_2785, n7684);
  not g10379 (n_2786, n7685);
  and g10380 (n7686, n_2785, n_2786);
  not g10381 (n_2787, n7683);
  and g10382 (n7687, n_2787, n7686);
  and g10383 (n7688, n_750, n7687);
  and g10384 (n7689, n_2206, n7687);
  not g10385 (n_2788, n7688);
  not g10386 (n_2789, n7689);
  and g10387 (n7690, n_2788, n_2789);
  not g10388 (n_2790, n7690);
  and g10389 (n7691, \a[26] , n_2790);
  and g10390 (n7692, n_33, n7690);
  not g10391 (n_2791, n7691);
  not g10392 (n_2792, n7692);
  and g10393 (n7693, n_2791, n_2792);
  not g10394 (n_2793, n7693);
  and g10395 (n7694, n7682, n_2793);
  not g10396 (n_2794, n7533);
  and g10397 (n7695, n7531, n_2794);
  not g10398 (n_2795, n7695);
  and g10399 (n7696, n_2653, n_2795);
  and g10400 (n7697, n_304, n3884);
  and g10401 (n7698, n_306, n3967);
  and g10402 (n7699, n_305, n4046);
  not g10403 (n_2796, n7698);
  not g10404 (n_2797, n7699);
  and g10405 (n7700, n_2796, n_2797);
  not g10406 (n_2798, n7697);
  and g10407 (n7701, n_2798, n7700);
  and g10408 (n7702, n_750, n7701);
  and g10409 (n7703, n_2351, n7701);
  not g10410 (n_2799, n7702);
  not g10411 (n_2800, n7703);
  and g10412 (n7704, n_2799, n_2800);
  not g10413 (n_2801, n7704);
  and g10414 (n7705, \a[26] , n_2801);
  and g10415 (n7706, n_33, n7704);
  not g10416 (n_2802, n7705);
  not g10417 (n_2803, n7706);
  and g10418 (n7707, n_2802, n_2803);
  not g10419 (n_2804, n7707);
  and g10420 (n7708, n7696, n_2804);
  and g10421 (n7709, n7402, n7529);
  not g10422 (n_2805, n7709);
  and g10423 (n7710, n_2649, n_2805);
  and g10424 (n7711, n_305, n3884);
  and g10425 (n7712, n_307, n3967);
  and g10426 (n7713, n_306, n4046);
  not g10427 (n_2806, n7712);
  not g10428 (n_2807, n7713);
  and g10429 (n7714, n_2806, n_2807);
  not g10430 (n_2808, n7711);
  and g10431 (n7715, n_2808, n7714);
  and g10432 (n7716, n_750, n7715);
  and g10433 (n7717, n_2051, n7715);
  not g10434 (n_2809, n7716);
  not g10435 (n_2810, n7717);
  and g10436 (n7718, n_2809, n_2810);
  not g10437 (n_2811, n7718);
  and g10438 (n7719, \a[26] , n_2811);
  and g10439 (n7720, n_33, n7718);
  not g10440 (n_2812, n7719);
  not g10441 (n_2813, n7720);
  and g10442 (n7721, n_2812, n_2813);
  not g10443 (n_2814, n7721);
  and g10444 (n7722, n7710, n_2814);
  and g10445 (n7723, n7420, n7527);
  not g10446 (n_2815, n7723);
  and g10447 (n7724, n_2646, n_2815);
  and g10448 (n7725, n_306, n3884);
  and g10449 (n7726, n_308, n3967);
  and g10450 (n7727, n_307, n4046);
  not g10451 (n_2816, n7726);
  not g10452 (n_2817, n7727);
  and g10453 (n7728, n_2816, n_2817);
  not g10454 (n_2818, n7725);
  and g10455 (n7729, n_2818, n7728);
  and g10456 (n7730, n_750, n7729);
  and g10457 (n7731, n_2498, n7729);
  not g10458 (n_2819, n7730);
  not g10459 (n_2820, n7731);
  and g10460 (n7732, n_2819, n_2820);
  not g10461 (n_2821, n7732);
  and g10462 (n7733, \a[26] , n_2821);
  and g10463 (n7734, n_33, n7732);
  not g10464 (n_2822, n7733);
  not g10465 (n_2823, n7734);
  and g10466 (n7735, n_2822, n_2823);
  not g10467 (n_2824, n7735);
  and g10468 (n7736, n7724, n_2824);
  and g10469 (n7737, n7438, n7525);
  not g10470 (n_2825, n7737);
  and g10471 (n7738, n_2643, n_2825);
  and g10472 (n7739, n_307, n3884);
  and g10473 (n7740, n_309, n3967);
  and g10474 (n7741, n_308, n4046);
  not g10475 (n_2826, n7740);
  not g10476 (n_2827, n7741);
  and g10477 (n7742, n_2826, n_2827);
  not g10478 (n_2828, n7739);
  and g10479 (n7743, n_2828, n7742);
  and g10480 (n7744, n_750, n7743);
  and g10481 (n7745, n_2511, n7743);
  not g10482 (n_2829, n7744);
  not g10483 (n_2830, n7745);
  and g10484 (n7746, n_2829, n_2830);
  not g10485 (n_2831, n7746);
  and g10486 (n7747, \a[26] , n_2831);
  and g10487 (n7748, n_33, n7746);
  not g10488 (n_2832, n7747);
  not g10489 (n_2833, n7748);
  and g10490 (n7749, n_2832, n_2833);
  not g10491 (n_2834, n7749);
  and g10492 (n7750, n7738, n_2834);
  and g10493 (n7751, n7456, n7523);
  not g10494 (n_2835, n7751);
  and g10495 (n7752, n_2640, n_2835);
  and g10496 (n7753, n_308, n3884);
  and g10497 (n7754, n_310, n3967);
  and g10498 (n7755, n_309, n4046);
  not g10499 (n_2836, n7754);
  not g10500 (n_2837, n7755);
  and g10501 (n7756, n_2836, n_2837);
  not g10502 (n_2838, n7753);
  and g10503 (n7757, n_2838, n7756);
  and g10504 (n7758, n_750, n7757);
  not g10505 (n_2839, n6122);
  and g10506 (n7759, n_2839, n7757);
  not g10507 (n_2840, n7758);
  not g10508 (n_2841, n7759);
  and g10509 (n7760, n_2840, n_2841);
  not g10510 (n_2842, n7760);
  and g10511 (n7761, \a[26] , n_2842);
  and g10512 (n7762, n_33, n7760);
  not g10513 (n_2843, n7761);
  not g10514 (n_2844, n7762);
  and g10515 (n7763, n_2843, n_2844);
  not g10516 (n_2845, n7763);
  and g10517 (n7764, n7752, n_2845);
  and g10518 (n7765, n_2635, n_2637);
  and g10519 (n7766, n_2636, n_2637);
  not g10520 (n_2846, n7765);
  not g10521 (n_2847, n7766);
  and g10522 (n7767, n_2846, n_2847);
  and g10523 (n7768, n_309, n3884);
  and g10524 (n7769, n_311, n3967);
  and g10525 (n7770, n_310, n4046);
  not g10526 (n_2848, n7769);
  not g10527 (n_2849, n7770);
  and g10528 (n7771, n_2848, n_2849);
  not g10529 (n_2850, n7768);
  and g10530 (n7772, n_2850, n7771);
  and g10531 (n7773, n_750, n7772);
  not g10532 (n_2851, n6541);
  and g10533 (n7774, n_2851, n7772);
  not g10534 (n_2852, n7773);
  not g10535 (n_2853, n7774);
  and g10536 (n7775, n_2852, n_2853);
  not g10537 (n_2854, n7775);
  and g10538 (n7776, \a[26] , n_2854);
  and g10539 (n7777, n_33, n7775);
  not g10540 (n_2855, n7776);
  not g10541 (n_2856, n7777);
  and g10542 (n7778, n_2855, n_2856);
  not g10543 (n_2857, n7767);
  not g10544 (n_2858, n7778);
  and g10545 (n7779, n_2857, n_2858);
  and g10546 (n7780, n_310, n3884);
  and g10547 (n7781, n_312, n3967);
  and g10548 (n7782, n_311, n4046);
  and g10554 (n7785, n4050, n6591);
  not g10557 (n_2863, n7786);
  and g10558 (n7787, \a[26] , n_2863);
  not g10559 (n_2864, n7787);
  and g10560 (n7788, n_2863, n_2864);
  and g10561 (n7789, \a[26] , n_2864);
  not g10562 (n_2865, n7788);
  not g10563 (n_2866, n7789);
  and g10564 (n7790, n_2865, n_2866);
  and g10565 (n7791, n7516, n7519);
  not g10566 (n_2867, n7791);
  and g10567 (n7792, n_2634, n_2867);
  not g10568 (n_2868, n7790);
  and g10569 (n7793, n_2868, n7792);
  not g10570 (n_2869, n7793);
  and g10571 (n7794, n_2868, n_2869);
  and g10572 (n7795, n7792, n_2869);
  not g10573 (n_2870, n7794);
  not g10574 (n_2871, n7795);
  and g10575 (n7796, n_2870, n_2871);
  and g10576 (n7797, n_311, n3884);
  and g10577 (n7798, n_313, n3967);
  and g10578 (n7799, n_312, n4046);
  and g10584 (n7802, n4050, n6646);
  not g10587 (n_2876, n7803);
  and g10588 (n7804, \a[26] , n_2876);
  not g10589 (n_2877, n7804);
  and g10590 (n7805, n_2876, n_2877);
  and g10591 (n7806, \a[26] , n_2877);
  not g10592 (n_2878, n7805);
  not g10593 (n_2879, n7806);
  and g10594 (n7807, n_2878, n_2879);
  not g10595 (n_2880, n7492);
  and g10596 (n7808, n_2880, n7503);
  not g10597 (n_2881, n7808);
  and g10598 (n7809, n_2628, n_2881);
  not g10599 (n_2882, n7807);
  and g10600 (n7810, n_2882, n7809);
  not g10601 (n_2883, n7810);
  and g10602 (n7811, n_2882, n_2883);
  and g10603 (n7812, n7809, n_2883);
  not g10604 (n_2884, n7811);
  not g10605 (n_2885, n7812);
  and g10606 (n7813, n_2884, n_2885);
  not g10607 (n_2886, n7491);
  and g10608 (n7814, n7489, n_2886);
  not g10609 (n_2887, n7814);
  and g10610 (n7815, n_2880, n_2887);
  and g10611 (n7816, n_312, n3884);
  and g10612 (n7817, n_314, n3967);
  and g10613 (n7818, n_313, n4046);
  not g10614 (n_2888, n7817);
  not g10615 (n_2889, n7818);
  and g10616 (n7819, n_2888, n_2889);
  not g10617 (n_2890, n7816);
  and g10618 (n7820, n_2890, n7819);
  and g10619 (n7821, n_750, n7820);
  not g10620 (n_2891, n6695);
  and g10621 (n7822, n_2891, n7820);
  not g10622 (n_2892, n7821);
  not g10623 (n_2893, n7822);
  and g10624 (n7823, n_2892, n_2893);
  not g10625 (n_2894, n7823);
  and g10626 (n7824, \a[26] , n_2894);
  and g10627 (n7825, n_33, n7823);
  not g10628 (n_2895, n7824);
  not g10629 (n_2896, n7825);
  and g10630 (n7826, n_2895, n_2896);
  not g10631 (n_2897, n7826);
  and g10632 (n7827, n7815, n_2897);
  and g10633 (n7828, n_316, n4046);
  and g10634 (n7829, n_315, n3884);
  not g10635 (n_2898, n7828);
  not g10636 (n_2899, n7829);
  and g10637 (n7830, n_2898, n_2899);
  and g10638 (n7831, n4050, n_2588);
  not g10639 (n_2900, n7831);
  and g10640 (n7832, n7830, n_2900);
  not g10641 (n_2901, n7832);
  and g10642 (n7833, \a[26] , n_2901);
  not g10643 (n_2902, n7833);
  and g10644 (n7834, \a[26] , n_2902);
  and g10645 (n7835, n_2901, n_2902);
  not g10646 (n_2903, n7834);
  not g10647 (n_2904, n7835);
  and g10648 (n7836, n_2903, n_2904);
  and g10649 (n7837, n_316, n_559);
  not g10650 (n_2905, n7837);
  and g10651 (n7838, \a[26] , n_2905);
  not g10652 (n_2906, n7836);
  and g10653 (n7839, n_2906, n7838);
  and g10654 (n7840, n_314, n3884);
  and g10655 (n7841, n_316, n3967);
  and g10656 (n7842, n_315, n4046);
  not g10657 (n_2907, n7841);
  not g10658 (n_2908, n7842);
  and g10659 (n7843, n_2907, n_2908);
  not g10660 (n_2909, n7840);
  and g10661 (n7844, n_2909, n7843);
  and g10662 (n7845, n_750, n7844);
  and g10663 (n7846, n_2612, n7844);
  not g10664 (n_2910, n7845);
  not g10665 (n_2911, n7846);
  and g10666 (n7847, n_2910, n_2911);
  not g10667 (n_2912, n7847);
  and g10668 (n7848, \a[26] , n_2912);
  and g10669 (n7849, n_33, n7847);
  not g10670 (n_2913, n7848);
  not g10671 (n_2914, n7849);
  and g10672 (n7850, n_2913, n_2914);
  not g10673 (n_2915, n7850);
  and g10674 (n7851, n7839, n_2915);
  and g10675 (n7852, n7490, n7851);
  not g10676 (n_2916, n7852);
  and g10677 (n7853, n7851, n_2916);
  and g10678 (n7854, n7490, n_2916);
  not g10679 (n_2917, n7853);
  not g10680 (n_2918, n7854);
  and g10681 (n7855, n_2917, n_2918);
  and g10682 (n7856, n_313, n3884);
  and g10683 (n7857, n_315, n3967);
  and g10684 (n7858, n_314, n4046);
  and g10690 (n7861, n4050, n6806);
  not g10693 (n_2923, n7862);
  and g10694 (n7863, \a[26] , n_2923);
  not g10695 (n_2924, n7863);
  and g10696 (n7864, \a[26] , n_2924);
  and g10697 (n7865, n_2923, n_2924);
  not g10698 (n_2925, n7864);
  not g10699 (n_2926, n7865);
  and g10700 (n7866, n_2925, n_2926);
  not g10701 (n_2927, n7855);
  not g10702 (n_2928, n7866);
  and g10703 (n7867, n_2927, n_2928);
  not g10704 (n_2929, n7867);
  and g10705 (n7868, n_2916, n_2929);
  not g10706 (n_2930, n7815);
  and g10707 (n7869, n_2930, n7826);
  not g10708 (n_2931, n7827);
  not g10709 (n_2932, n7869);
  and g10710 (n7870, n_2931, n_2932);
  not g10711 (n_2933, n7868);
  and g10712 (n7871, n_2933, n7870);
  not g10713 (n_2934, n7871);
  and g10714 (n7872, n_2931, n_2934);
  not g10715 (n_2935, n7813);
  not g10716 (n_2936, n7872);
  and g10717 (n7873, n_2935, n_2936);
  not g10718 (n_2937, n7873);
  and g10719 (n7874, n_2883, n_2937);
  not g10720 (n_2938, n7796);
  not g10721 (n_2939, n7874);
  and g10722 (n7875, n_2938, n_2939);
  not g10723 (n_2940, n7875);
  and g10724 (n7876, n_2869, n_2940);
  not g10725 (n_2941, n7779);
  and g10726 (n7877, n_2857, n_2941);
  and g10727 (n7878, n_2858, n_2941);
  not g10728 (n_2942, n7877);
  not g10729 (n_2943, n7878);
  and g10730 (n7879, n_2942, n_2943);
  not g10731 (n_2944, n7876);
  not g10732 (n_2945, n7879);
  and g10733 (n7880, n_2944, n_2945);
  not g10734 (n_2946, n7880);
  and g10735 (n7881, n_2941, n_2946);
  not g10736 (n_2947, n7764);
  and g10737 (n7882, n7752, n_2947);
  and g10738 (n7883, n_2845, n_2947);
  not g10739 (n_2948, n7882);
  not g10740 (n_2949, n7883);
  and g10741 (n7884, n_2948, n_2949);
  not g10742 (n_2950, n7881);
  not g10743 (n_2951, n7884);
  and g10744 (n7885, n_2950, n_2951);
  not g10745 (n_2952, n7885);
  and g10746 (n7886, n_2947, n_2952);
  not g10747 (n_2953, n7750);
  and g10748 (n7887, n7738, n_2953);
  and g10749 (n7888, n_2834, n_2953);
  not g10750 (n_2954, n7887);
  not g10751 (n_2955, n7888);
  and g10752 (n7889, n_2954, n_2955);
  not g10753 (n_2956, n7886);
  not g10754 (n_2957, n7889);
  and g10755 (n7890, n_2956, n_2957);
  not g10756 (n_2958, n7890);
  and g10757 (n7891, n_2953, n_2958);
  not g10758 (n_2959, n7736);
  and g10759 (n7892, n7724, n_2959);
  and g10760 (n7893, n_2824, n_2959);
  not g10761 (n_2960, n7892);
  not g10762 (n_2961, n7893);
  and g10763 (n7894, n_2960, n_2961);
  not g10764 (n_2962, n7891);
  not g10765 (n_2963, n7894);
  and g10766 (n7895, n_2962, n_2963);
  not g10767 (n_2964, n7895);
  and g10768 (n7896, n_2959, n_2964);
  not g10769 (n_2965, n7722);
  and g10770 (n7897, n7710, n_2965);
  and g10771 (n7898, n_2814, n_2965);
  not g10772 (n_2966, n7897);
  not g10773 (n_2967, n7898);
  and g10774 (n7899, n_2966, n_2967);
  not g10775 (n_2968, n7896);
  not g10776 (n_2969, n7899);
  and g10777 (n7900, n_2968, n_2969);
  not g10778 (n_2970, n7900);
  and g10779 (n7901, n_2965, n_2970);
  not g10780 (n_2971, n7708);
  and g10781 (n7902, n7696, n_2971);
  and g10782 (n7903, n_2804, n_2971);
  not g10783 (n_2972, n7902);
  not g10784 (n_2973, n7903);
  and g10785 (n7904, n_2972, n_2973);
  not g10786 (n_2974, n7901);
  not g10787 (n_2975, n7904);
  and g10788 (n7905, n_2974, n_2975);
  not g10789 (n_2976, n7905);
  and g10790 (n7906, n_2971, n_2976);
  not g10791 (n_2977, n7694);
  and g10792 (n7907, n7682, n_2977);
  and g10793 (n7908, n_2793, n_2977);
  not g10794 (n_2978, n7907);
  not g10795 (n_2979, n7908);
  and g10796 (n7909, n_2978, n_2979);
  not g10797 (n_2980, n7906);
  not g10798 (n_2981, n7909);
  and g10799 (n7910, n_2980, n_2981);
  not g10800 (n_2982, n7910);
  and g10801 (n7911, n_2977, n_2982);
  not g10802 (n_2983, n7555);
  and g10803 (n7912, n7553, n_2983);
  not g10804 (n_2984, n7912);
  and g10805 (n7913, n_2673, n_2984);
  not g10806 (n_2985, n7911);
  and g10807 (n7914, n_2985, n7913);
  and g10808 (n7915, n_299, n4694);
  and g10809 (n7916, n_301, n4533);
  and g10810 (n7917, n_300, n4604);
  and g10816 (n7920, n4536, n5139);
  not g10819 (n_2990, n7921);
  and g10820 (n7922, \a[23] , n_2990);
  not g10821 (n_2991, n7922);
  and g10822 (n7923, n_2990, n_2991);
  and g10823 (n7924, \a[23] , n_2991);
  not g10824 (n_2992, n7923);
  not g10825 (n_2993, n7924);
  and g10826 (n7925, n_2992, n_2993);
  not g10827 (n_2994, n7913);
  and g10828 (n7926, n7911, n_2994);
  not g10829 (n_2995, n7914);
  not g10830 (n_2996, n7926);
  and g10831 (n7927, n_2995, n_2996);
  not g10832 (n_2997, n7925);
  and g10833 (n7928, n_2997, n7927);
  not g10834 (n_2998, n7928);
  and g10835 (n7929, n_2995, n_2998);
  not g10836 (n_2999, n7680);
  not g10837 (n_3000, n7929);
  and g10838 (n7930, n_2999, n_3000);
  and g10839 (n7931, n7680, n7929);
  not g10840 (n_3001, n7930);
  not g10841 (n_3002, n7931);
  and g10842 (n7932, n_3001, n_3002);
  and g10843 (n7933, n_286, n5496);
  and g10844 (n7934, n_295, n4935);
  and g10845 (n7935, n_293, n5407);
  and g10851 (n7938, n4429, n4938);
  not g10854 (n_3007, n7939);
  and g10855 (n7940, \a[20] , n_3007);
  not g10856 (n_3008, n7940);
  and g10857 (n7941, \a[20] , n_3008);
  and g10858 (n7942, n_3007, n_3008);
  not g10859 (n_3009, n7941);
  not g10860 (n_3010, n7942);
  and g10861 (n7943, n_3009, n_3010);
  not g10862 (n_3011, n7943);
  and g10863 (n7944, n7932, n_3011);
  not g10864 (n_3012, n7944);
  and g10865 (n7945, n_3001, n_3012);
  not g10866 (n_3013, n7677);
  not g10867 (n_3014, n7945);
  and g10868 (n7946, n_3013, n_3014);
  and g10869 (n7947, n7677, n7945);
  not g10870 (n_3015, n7946);
  not g10871 (n_3016, n7947);
  and g10872 (n7948, n_3015, n_3016);
  and g10873 (n7949, n_237, n6233);
  and g10874 (n7950, n_275, n5663);
  and g10875 (n7951, n_260, n5939);
  and g10881 (n7954, n3331, n5666);
  not g10884 (n_3021, n7955);
  and g10885 (n7956, \a[17] , n_3021);
  not g10886 (n_3022, n7956);
  and g10887 (n7957, \a[17] , n_3022);
  and g10888 (n7958, n_3021, n_3022);
  not g10889 (n_3023, n7957);
  not g10890 (n_3024, n7958);
  and g10891 (n7959, n_3023, n_3024);
  not g10892 (n_3025, n7959);
  and g10893 (n7960, n7948, n_3025);
  not g10894 (n_3026, n7960);
  and g10895 (n7961, n_3015, n_3026);
  not g10896 (n_3027, n7674);
  not g10897 (n_3028, n7961);
  and g10898 (n7962, n_3027, n_3028);
  not g10899 (n_3029, n7962);
  and g10900 (n7963, n_2776, n_3029);
  not g10901 (n_3030, n7657);
  not g10902 (n_3031, n7963);
  and g10903 (n7964, n_3030, n_3031);
  and g10904 (n7965, n7657, n7963);
  not g10905 (n_3032, n7964);
  not g10906 (n_3033, n7965);
  and g10907 (n7966, n_3032, n_3033);
  and g10908 (n7967, n_480, n7101);
  and g10909 (n7968, n_484, n6402);
  and g10910 (n7969, n_485, n6951);
  and g10916 (n7972, n3627, n6397);
  not g10919 (n_3038, n7973);
  and g10920 (n7974, \a[14] , n_3038);
  not g10921 (n_3039, n7974);
  and g10922 (n7975, \a[14] , n_3039);
  and g10923 (n7976, n_3038, n_3039);
  not g10924 (n_3040, n7975);
  not g10925 (n_3041, n7976);
  and g10926 (n7977, n_3040, n_3041);
  not g10927 (n_3042, n7977);
  and g10928 (n7978, n7966, n_3042);
  not g10929 (n_3043, n7978);
  and g10930 (n7979, n_3032, n_3043);
  not g10931 (n_3044, n7654);
  not g10932 (n_3045, n7979);
  and g10933 (n7980, n_3044, n_3045);
  and g10934 (n7981, n7654, n7979);
  not g10935 (n_3046, n7980);
  not g10936 (n_3047, n7981);
  and g10937 (n7982, n_3046, n_3047);
  and g10938 (n7983, n7286, n_2445);
  and g10939 (n7984, n_560, n7983);
  and g10940 (n7985, n_565, n7291);
  and g10941 (n7986, n_566, n7632);
  and g10947 (n7989, n4067, n7294);
  not g10950 (n_3052, n7990);
  and g10951 (n7991, \a[11] , n_3052);
  not g10952 (n_3053, n7991);
  and g10953 (n7992, \a[11] , n_3053);
  and g10954 (n7993, n_3052, n_3053);
  not g10955 (n_3054, n7992);
  not g10956 (n_3055, n7993);
  and g10957 (n7994, n_3054, n_3055);
  not g10958 (n_3056, n7994);
  and g10959 (n7995, n7982, n_3056);
  not g10960 (n_3057, n7995);
  and g10961 (n7996, n_3046, n_3057);
  and g10962 (n7997, n_712, n7983);
  and g10963 (n7998, n_566, n7291);
  and g10964 (n7999, n_560, n7632);
  not g10965 (n_3058, n7998);
  not g10966 (n_3059, n7999);
  and g10967 (n8000, n_3058, n_3059);
  not g10968 (n_3060, n7997);
  and g10969 (n8001, n_3060, n8000);
  and g10970 (n8002, n_2446, n8001);
  and g10971 (n8003, n_888, n8001);
  not g10972 (n_3061, n8002);
  not g10973 (n_3062, n8003);
  and g10974 (n8004, n_3061, n_3062);
  not g10975 (n_3063, n8004);
  and g10976 (n8005, \a[11] , n_3063);
  and g10977 (n8006, n_1071, n8004);
  not g10978 (n_3064, n8005);
  not g10979 (n_3065, n8006);
  and g10980 (n8007, n_3064, n_3065);
  not g10981 (n_3066, n7996);
  not g10982 (n_3067, n8007);
  and g10983 (n8008, n_3066, n_3067);
  and g10984 (n8009, n7996, n8007);
  not g10985 (n_3068, n8008);
  not g10986 (n_3069, n8009);
  and g10987 (n8010, n_3068, n_3069);
  and g10988 (n8011, n_2738, n_2740);
  and g10989 (n8012, n_2739, n_2740);
  not g10990 (n_3070, n8011);
  not g10991 (n_3071, n8012);
  and g10992 (n8013, n_3070, n_3071);
  not g10993 (n_3072, n8013);
  and g10994 (n8014, n8010, n_3072);
  not g10995 (n_3073, n8014);
  and g10996 (n8015, n_3068, n_3073);
  not g10997 (n_3074, n7646);
  and g10998 (n8016, n7644, n_3074);
  not g10999 (n_3075, n8016);
  and g11000 (n8017, n_2756, n_3075);
  not g11001 (n_3076, n8015);
  and g11002 (n8018, n_3076, n8017);
  and g11003 (n8019, n8010, n_3073);
  and g11004 (n8020, n_3072, n_3073);
  not g11005 (n_3077, n8019);
  not g11006 (n_3078, n8020);
  and g11007 (n8021, n_3077, n_3078);
  and g11008 (n8022, n7966, n_3043);
  and g11009 (n8023, n_3042, n_3043);
  not g11010 (n_3079, n8022);
  not g11011 (n_3080, n8023);
  and g11012 (n8024, n_3079, n_3080);
  and g11013 (n8025, n7674, n7961);
  not g11014 (n_3081, n8025);
  and g11015 (n8026, n_3029, n_3081);
  and g11016 (n8027, n_485, n7101);
  and g11017 (n8028, n_415, n6402);
  and g11018 (n8029, n_484, n6951);
  not g11019 (n_3082, n8028);
  not g11020 (n_3083, n8029);
  and g11021 (n8030, n_3082, n_3083);
  not g11022 (n_3084, n8027);
  and g11023 (n8031, n_3084, n8030);
  and g11024 (n8032, n_1885, n8031);
  and g11025 (n8033, n_914, n8031);
  not g11026 (n_3085, n8032);
  not g11027 (n_3086, n8033);
  and g11028 (n8034, n_3085, n_3086);
  not g11029 (n_3087, n8034);
  and g11030 (n8035, \a[14] , n_3087);
  and g11031 (n8036, n_652, n8034);
  not g11032 (n_3088, n8035);
  not g11033 (n_3089, n8036);
  and g11034 (n8037, n_3088, n_3089);
  not g11035 (n_3090, n8037);
  and g11036 (n8038, n8026, n_3090);
  and g11037 (n8039, n7948, n_3026);
  and g11038 (n8040, n_3025, n_3026);
  not g11039 (n_3091, n8039);
  not g11040 (n_3092, n8040);
  and g11041 (n8041, n_3091, n_3092);
  and g11042 (n8042, n7932, n_3012);
  and g11043 (n8043, n_3011, n_3012);
  not g11044 (n_3093, n8042);
  not g11045 (n_3094, n8043);
  and g11046 (n8044, n_3093, n_3094);
  and g11047 (n8045, n_300, n4694);
  and g11048 (n8046, n_302, n4533);
  and g11049 (n8047, n_301, n4604);
  and g11055 (n8050, n4536, n5561);
  not g11058 (n_3099, n8051);
  and g11059 (n8052, \a[23] , n_3099);
  not g11060 (n_3100, n8052);
  and g11061 (n8053, n_3099, n_3100);
  and g11062 (n8054, \a[23] , n_3100);
  not g11063 (n_3101, n8053);
  not g11064 (n_3102, n8054);
  and g11065 (n8055, n_3101, n_3102);
  and g11066 (n8056, n_2980, n_2982);
  and g11067 (n8057, n_2981, n_2982);
  not g11068 (n_3103, n8056);
  not g11069 (n_3104, n8057);
  and g11070 (n8058, n_3103, n_3104);
  not g11071 (n_3105, n8055);
  not g11072 (n_3106, n8058);
  and g11073 (n8059, n_3105, n_3106);
  not g11074 (n_3107, n8059);
  and g11075 (n8060, n_3105, n_3107);
  and g11076 (n8061, n_3106, n_3107);
  not g11077 (n_3108, n8060);
  not g11078 (n_3109, n8061);
  and g11079 (n8062, n_3108, n_3109);
  and g11080 (n8063, n_301, n4694);
  and g11081 (n8064, n_303, n4533);
  and g11082 (n8065, n_302, n4604);
  and g11088 (n8068, n4536, n5328);
  not g11091 (n_3114, n8069);
  and g11092 (n8070, \a[23] , n_3114);
  not g11093 (n_3115, n8070);
  and g11094 (n8071, n_3114, n_3115);
  and g11095 (n8072, \a[23] , n_3115);
  not g11096 (n_3116, n8071);
  not g11097 (n_3117, n8072);
  and g11098 (n8073, n_3116, n_3117);
  and g11099 (n8074, n_2974, n_2976);
  and g11100 (n8075, n_2975, n_2976);
  not g11101 (n_3118, n8074);
  not g11102 (n_3119, n8075);
  and g11103 (n8076, n_3118, n_3119);
  not g11104 (n_3120, n8073);
  not g11105 (n_3121, n8076);
  and g11106 (n8077, n_3120, n_3121);
  not g11107 (n_3122, n8077);
  and g11108 (n8078, n_3120, n_3122);
  and g11109 (n8079, n_3121, n_3122);
  not g11110 (n_3123, n8078);
  not g11111 (n_3124, n8079);
  and g11112 (n8080, n_3123, n_3124);
  and g11113 (n8081, n_302, n4694);
  and g11114 (n8082, n_304, n4533);
  and g11115 (n8083, n_303, n4604);
  and g11121 (n8086, n4536, n5851);
  not g11124 (n_3129, n8087);
  and g11125 (n8088, \a[23] , n_3129);
  not g11126 (n_3130, n8088);
  and g11127 (n8089, n_3129, n_3130);
  and g11128 (n8090, \a[23] , n_3130);
  not g11129 (n_3131, n8089);
  not g11130 (n_3132, n8090);
  and g11131 (n8091, n_3131, n_3132);
  and g11132 (n8092, n_2968, n_2970);
  and g11133 (n8093, n_2969, n_2970);
  not g11134 (n_3133, n8092);
  not g11135 (n_3134, n8093);
  and g11136 (n8094, n_3133, n_3134);
  not g11137 (n_3135, n8091);
  not g11138 (n_3136, n8094);
  and g11139 (n8095, n_3135, n_3136);
  not g11140 (n_3137, n8095);
  and g11141 (n8096, n_3135, n_3137);
  and g11142 (n8097, n_3136, n_3137);
  not g11143 (n_3138, n8096);
  not g11144 (n_3139, n8097);
  and g11145 (n8098, n_3138, n_3139);
  and g11146 (n8099, n_303, n4694);
  and g11147 (n8100, n_305, n4533);
  and g11148 (n8101, n_304, n4604);
  and g11154 (n8104, n4536, n6007);
  not g11157 (n_3144, n8105);
  and g11158 (n8106, \a[23] , n_3144);
  not g11159 (n_3145, n8106);
  and g11160 (n8107, n_3144, n_3145);
  and g11161 (n8108, \a[23] , n_3145);
  not g11162 (n_3146, n8107);
  not g11163 (n_3147, n8108);
  and g11164 (n8109, n_3146, n_3147);
  and g11165 (n8110, n_2962, n_2964);
  and g11166 (n8111, n_2963, n_2964);
  not g11167 (n_3148, n8110);
  not g11168 (n_3149, n8111);
  and g11169 (n8112, n_3148, n_3149);
  not g11170 (n_3150, n8109);
  not g11171 (n_3151, n8112);
  and g11172 (n8113, n_3150, n_3151);
  not g11173 (n_3152, n8113);
  and g11174 (n8114, n_3150, n_3152);
  and g11175 (n8115, n_3151, n_3152);
  not g11176 (n_3153, n8114);
  not g11177 (n_3154, n8115);
  and g11178 (n8116, n_3153, n_3154);
  and g11179 (n8117, n_304, n4694);
  and g11180 (n8118, n_306, n4533);
  and g11181 (n8119, n_305, n4604);
  and g11187 (n8122, n4536, n5834);
  not g11190 (n_3159, n8123);
  and g11191 (n8124, \a[23] , n_3159);
  not g11192 (n_3160, n8124);
  and g11193 (n8125, n_3159, n_3160);
  and g11194 (n8126, \a[23] , n_3160);
  not g11195 (n_3161, n8125);
  not g11196 (n_3162, n8126);
  and g11197 (n8127, n_3161, n_3162);
  and g11198 (n8128, n_2956, n_2958);
  and g11199 (n8129, n_2957, n_2958);
  not g11200 (n_3163, n8128);
  not g11201 (n_3164, n8129);
  and g11202 (n8130, n_3163, n_3164);
  not g11203 (n_3165, n8127);
  not g11204 (n_3166, n8130);
  and g11205 (n8131, n_3165, n_3166);
  not g11206 (n_3167, n8131);
  and g11207 (n8132, n_3165, n_3167);
  and g11208 (n8133, n_3166, n_3167);
  not g11209 (n_3168, n8132);
  not g11210 (n_3169, n8133);
  and g11211 (n8134, n_3168, n_3169);
  and g11212 (n8135, n_305, n4694);
  and g11213 (n8136, n_307, n4533);
  and g11214 (n8137, n_306, n4604);
  and g11220 (n8140, n4536, n6143);
  not g11223 (n_3174, n8141);
  and g11224 (n8142, \a[23] , n_3174);
  not g11225 (n_3175, n8142);
  and g11226 (n8143, n_3174, n_3175);
  and g11227 (n8144, \a[23] , n_3175);
  not g11228 (n_3176, n8143);
  not g11229 (n_3177, n8144);
  and g11230 (n8145, n_3176, n_3177);
  and g11231 (n8146, n_2950, n_2952);
  and g11232 (n8147, n_2951, n_2952);
  not g11233 (n_3178, n8146);
  not g11234 (n_3179, n8147);
  and g11235 (n8148, n_3178, n_3179);
  not g11236 (n_3180, n8145);
  not g11237 (n_3181, n8148);
  and g11238 (n8149, n_3180, n_3181);
  not g11239 (n_3182, n8149);
  and g11240 (n8150, n_3180, n_3182);
  and g11241 (n8151, n_3181, n_3182);
  not g11242 (n_3183, n8150);
  not g11243 (n_3184, n8151);
  and g11244 (n8152, n_3183, n_3184);
  and g11245 (n8153, n_306, n4694);
  and g11246 (n8154, n_308, n4533);
  and g11247 (n8155, n_307, n4604);
  and g11253 (n8158, n4536, n6479);
  not g11256 (n_3189, n8159);
  and g11257 (n8160, \a[23] , n_3189);
  not g11258 (n_3190, n8160);
  and g11259 (n8161, n_3189, n_3190);
  and g11260 (n8162, \a[23] , n_3190);
  not g11261 (n_3191, n8161);
  not g11262 (n_3192, n8162);
  and g11263 (n8163, n_3191, n_3192);
  and g11264 (n8164, n_2944, n_2946);
  and g11265 (n8165, n_2945, n_2946);
  not g11266 (n_3193, n8164);
  not g11267 (n_3194, n8165);
  and g11268 (n8166, n_3193, n_3194);
  not g11269 (n_3195, n8163);
  not g11270 (n_3196, n8166);
  and g11271 (n8167, n_3195, n_3196);
  not g11272 (n_3197, n8167);
  and g11273 (n8168, n_3195, n_3197);
  and g11274 (n8169, n_3196, n_3197);
  not g11275 (n_3198, n8168);
  not g11276 (n_3199, n8169);
  and g11277 (n8170, n_3198, n_3199);
  and g11278 (n8171, n7796, n7874);
  not g11279 (n_3200, n8171);
  and g11280 (n8172, n_2940, n_3200);
  and g11281 (n8173, n_307, n4694);
  and g11282 (n8174, n_309, n4533);
  and g11283 (n8175, n_308, n4604);
  not g11284 (n_3201, n8174);
  not g11285 (n_3202, n8175);
  and g11286 (n8176, n_3201, n_3202);
  not g11287 (n_3203, n8173);
  and g11288 (n8177, n_3203, n8176);
  and g11289 (n8178, n_732, n8177);
  and g11290 (n8179, n_2511, n8177);
  not g11291 (n_3204, n8178);
  not g11292 (n_3205, n8179);
  and g11293 (n8180, n_3204, n_3205);
  not g11294 (n_3206, n8180);
  and g11295 (n8181, \a[23] , n_3206);
  and g11296 (n8182, n_27, n8180);
  not g11297 (n_3207, n8181);
  not g11298 (n_3208, n8182);
  and g11299 (n8183, n_3207, n_3208);
  not g11300 (n_3209, n8183);
  and g11301 (n8184, n8172, n_3209);
  and g11302 (n8185, n7813, n7872);
  not g11303 (n_3210, n8185);
  and g11304 (n8186, n_2937, n_3210);
  and g11305 (n8187, n_308, n4694);
  and g11306 (n8188, n_310, n4533);
  and g11307 (n8189, n_309, n4604);
  not g11308 (n_3211, n8188);
  not g11309 (n_3212, n8189);
  and g11310 (n8190, n_3211, n_3212);
  not g11311 (n_3213, n8187);
  and g11312 (n8191, n_3213, n8190);
  and g11313 (n8192, n_732, n8191);
  and g11314 (n8193, n_2839, n8191);
  not g11315 (n_3214, n8192);
  not g11316 (n_3215, n8193);
  and g11317 (n8194, n_3214, n_3215);
  not g11318 (n_3216, n8194);
  and g11319 (n8195, \a[23] , n_3216);
  and g11320 (n8196, n_27, n8194);
  not g11321 (n_3217, n8195);
  not g11322 (n_3218, n8196);
  and g11323 (n8197, n_3217, n_3218);
  not g11324 (n_3219, n8197);
  and g11325 (n8198, n8186, n_3219);
  and g11326 (n8199, n_309, n4694);
  and g11327 (n8200, n_311, n4533);
  and g11328 (n8201, n_310, n4604);
  and g11334 (n8204, n4536, n6541);
  not g11337 (n_3224, n8205);
  and g11338 (n8206, \a[23] , n_3224);
  not g11339 (n_3225, n8206);
  and g11340 (n8207, n_3224, n_3225);
  and g11341 (n8208, \a[23] , n_3225);
  not g11342 (n_3226, n8207);
  not g11343 (n_3227, n8208);
  and g11344 (n8209, n_3226, n_3227);
  not g11345 (n_3228, n7870);
  and g11346 (n8210, n7868, n_3228);
  not g11347 (n_3229, n8210);
  and g11348 (n8211, n_2934, n_3229);
  not g11349 (n_3230, n8209);
  and g11350 (n8212, n_3230, n8211);
  not g11351 (n_3231, n8212);
  and g11352 (n8213, n_3230, n_3231);
  and g11353 (n8214, n8211, n_3231);
  not g11354 (n_3232, n8213);
  not g11355 (n_3233, n8214);
  and g11356 (n8215, n_3232, n_3233);
  and g11357 (n8216, n_2927, n_2929);
  and g11358 (n8217, n_2928, n_2929);
  not g11359 (n_3234, n8216);
  not g11360 (n_3235, n8217);
  and g11361 (n8218, n_3234, n_3235);
  and g11362 (n8219, n_310, n4694);
  and g11363 (n8220, n_312, n4533);
  and g11364 (n8221, n_311, n4604);
  not g11365 (n_3236, n8220);
  not g11366 (n_3237, n8221);
  and g11367 (n8222, n_3236, n_3237);
  not g11368 (n_3238, n8219);
  and g11369 (n8223, n_3238, n8222);
  and g11370 (n8224, n_732, n8223);
  not g11371 (n_3239, n6591);
  and g11372 (n8225, n_3239, n8223);
  not g11373 (n_3240, n8224);
  not g11374 (n_3241, n8225);
  and g11375 (n8226, n_3240, n_3241);
  not g11376 (n_3242, n8226);
  and g11377 (n8227, \a[23] , n_3242);
  and g11378 (n8228, n_27, n8226);
  not g11379 (n_3243, n8227);
  not g11380 (n_3244, n8228);
  and g11381 (n8229, n_3243, n_3244);
  not g11382 (n_3245, n8218);
  not g11383 (n_3246, n8229);
  and g11384 (n8230, n_3245, n_3246);
  and g11385 (n8231, n_311, n4694);
  and g11386 (n8232, n_313, n4533);
  and g11387 (n8233, n_312, n4604);
  and g11393 (n8236, n4536, n6646);
  not g11396 (n_3251, n8237);
  and g11397 (n8238, \a[23] , n_3251);
  not g11398 (n_3252, n8238);
  and g11399 (n8239, n_3251, n_3252);
  and g11400 (n8240, \a[23] , n_3252);
  not g11401 (n_3253, n8239);
  not g11402 (n_3254, n8240);
  and g11403 (n8241, n_3253, n_3254);
  not g11404 (n_3255, n7839);
  and g11405 (n8242, n_3255, n7850);
  not g11406 (n_3256, n7851);
  not g11407 (n_3257, n8242);
  and g11408 (n8243, n_3256, n_3257);
  not g11409 (n_3258, n8241);
  and g11410 (n8244, n_3258, n8243);
  not g11411 (n_3259, n8244);
  and g11412 (n8245, n_3258, n_3259);
  and g11413 (n8246, n8243, n_3259);
  not g11414 (n_3260, n8245);
  not g11415 (n_3261, n8246);
  and g11416 (n8247, n_3260, n_3261);
  not g11417 (n_3262, n7838);
  and g11418 (n8248, n7836, n_3262);
  not g11419 (n_3263, n8248);
  and g11420 (n8249, n_3255, n_3263);
  and g11421 (n8250, n_312, n4694);
  and g11422 (n8251, n_314, n4533);
  and g11423 (n8252, n_313, n4604);
  not g11424 (n_3264, n8251);
  not g11425 (n_3265, n8252);
  and g11426 (n8253, n_3264, n_3265);
  not g11427 (n_3266, n8250);
  and g11428 (n8254, n_3266, n8253);
  and g11429 (n8255, n_732, n8254);
  and g11430 (n8256, n_2891, n8254);
  not g11431 (n_3267, n8255);
  not g11432 (n_3268, n8256);
  and g11433 (n8257, n_3267, n_3268);
  not g11434 (n_3269, n8257);
  and g11435 (n8258, \a[23] , n_3269);
  and g11436 (n8259, n_27, n8257);
  not g11437 (n_3270, n8258);
  not g11438 (n_3271, n8259);
  and g11439 (n8260, n_3270, n_3271);
  not g11440 (n_3272, n8260);
  and g11441 (n8261, n8249, n_3272);
  and g11442 (n8262, n_316, n4604);
  and g11443 (n8263, n_315, n4694);
  not g11444 (n_3273, n8262);
  not g11445 (n_3274, n8263);
  and g11446 (n8264, n_3273, n_3274);
  and g11447 (n8265, n4536, n_2588);
  not g11448 (n_3275, n8265);
  and g11449 (n8266, n8264, n_3275);
  not g11450 (n_3276, n8266);
  and g11451 (n8267, \a[23] , n_3276);
  not g11452 (n_3277, n8267);
  and g11453 (n8268, \a[23] , n_3277);
  and g11454 (n8269, n_3276, n_3277);
  not g11455 (n_3278, n8268);
  not g11456 (n_3279, n8269);
  and g11457 (n8270, n_3278, n_3279);
  and g11458 (n8271, n_316, n_731);
  not g11459 (n_3280, n8271);
  and g11460 (n8272, \a[23] , n_3280);
  not g11461 (n_3281, n8270);
  and g11462 (n8273, n_3281, n8272);
  and g11463 (n8274, n_314, n4694);
  and g11464 (n8275, n_316, n4533);
  and g11465 (n8276, n_315, n4604);
  not g11466 (n_3282, n8275);
  not g11467 (n_3283, n8276);
  and g11468 (n8277, n_3282, n_3283);
  not g11469 (n_3284, n8274);
  and g11470 (n8278, n_3284, n8277);
  and g11471 (n8279, n_732, n8278);
  and g11472 (n8280, n_2612, n8278);
  not g11473 (n_3285, n8279);
  not g11474 (n_3286, n8280);
  and g11475 (n8281, n_3285, n_3286);
  not g11476 (n_3287, n8281);
  and g11477 (n8282, \a[23] , n_3287);
  and g11478 (n8283, n_27, n8281);
  not g11479 (n_3288, n8282);
  not g11480 (n_3289, n8283);
  and g11481 (n8284, n_3288, n_3289);
  not g11482 (n_3290, n8284);
  and g11483 (n8285, n8273, n_3290);
  and g11484 (n8286, n7837, n8285);
  not g11485 (n_3291, n8286);
  and g11486 (n8287, n8285, n_3291);
  and g11487 (n8288, n7837, n_3291);
  not g11488 (n_3292, n8287);
  not g11489 (n_3293, n8288);
  and g11490 (n8289, n_3292, n_3293);
  and g11491 (n8290, n_313, n4694);
  and g11492 (n8291, n_315, n4533);
  and g11493 (n8292, n_314, n4604);
  and g11499 (n8295, n4536, n6806);
  not g11502 (n_3298, n8296);
  and g11503 (n8297, \a[23] , n_3298);
  not g11504 (n_3299, n8297);
  and g11505 (n8298, \a[23] , n_3299);
  and g11506 (n8299, n_3298, n_3299);
  not g11507 (n_3300, n8298);
  not g11508 (n_3301, n8299);
  and g11509 (n8300, n_3300, n_3301);
  not g11510 (n_3302, n8289);
  not g11511 (n_3303, n8300);
  and g11512 (n8301, n_3302, n_3303);
  not g11513 (n_3304, n8301);
  and g11514 (n8302, n_3291, n_3304);
  not g11515 (n_3305, n8249);
  and g11516 (n8303, n_3305, n8260);
  not g11517 (n_3306, n8261);
  not g11518 (n_3307, n8303);
  and g11519 (n8304, n_3306, n_3307);
  not g11520 (n_3308, n8302);
  and g11521 (n8305, n_3308, n8304);
  not g11522 (n_3309, n8305);
  and g11523 (n8306, n_3306, n_3309);
  not g11524 (n_3310, n8247);
  not g11525 (n_3311, n8306);
  and g11526 (n8307, n_3310, n_3311);
  not g11527 (n_3312, n8307);
  and g11528 (n8308, n_3259, n_3312);
  and g11529 (n8309, n8218, n8229);
  not g11530 (n_3313, n8230);
  not g11531 (n_3314, n8309);
  and g11532 (n8310, n_3313, n_3314);
  not g11533 (n_3315, n8308);
  and g11534 (n8311, n_3315, n8310);
  not g11535 (n_3316, n8311);
  and g11536 (n8312, n_3313, n_3316);
  not g11537 (n_3317, n8215);
  not g11538 (n_3318, n8312);
  and g11539 (n8313, n_3317, n_3318);
  not g11540 (n_3319, n8313);
  and g11541 (n8314, n_3231, n_3319);
  not g11542 (n_3320, n8198);
  and g11543 (n8315, n8186, n_3320);
  and g11544 (n8316, n_3219, n_3320);
  not g11545 (n_3321, n8315);
  not g11546 (n_3322, n8316);
  and g11547 (n8317, n_3321, n_3322);
  not g11548 (n_3323, n8314);
  not g11549 (n_3324, n8317);
  and g11550 (n8318, n_3323, n_3324);
  not g11551 (n_3325, n8318);
  and g11552 (n8319, n_3320, n_3325);
  not g11553 (n_3326, n8172);
  and g11554 (n8320, n_3326, n8183);
  not g11555 (n_3327, n8184);
  not g11556 (n_3328, n8320);
  and g11557 (n8321, n_3327, n_3328);
  not g11558 (n_3329, n8319);
  and g11559 (n8322, n_3329, n8321);
  not g11560 (n_3330, n8322);
  and g11561 (n8323, n_3327, n_3330);
  not g11562 (n_3331, n8170);
  not g11563 (n_3332, n8323);
  and g11564 (n8324, n_3331, n_3332);
  not g11565 (n_3333, n8324);
  and g11566 (n8325, n_3197, n_3333);
  not g11567 (n_3334, n8152);
  not g11568 (n_3335, n8325);
  and g11569 (n8326, n_3334, n_3335);
  not g11570 (n_3336, n8326);
  and g11571 (n8327, n_3182, n_3336);
  not g11572 (n_3337, n8134);
  not g11573 (n_3338, n8327);
  and g11574 (n8328, n_3337, n_3338);
  not g11575 (n_3339, n8328);
  and g11576 (n8329, n_3167, n_3339);
  not g11577 (n_3340, n8116);
  not g11578 (n_3341, n8329);
  and g11579 (n8330, n_3340, n_3341);
  not g11580 (n_3342, n8330);
  and g11581 (n8331, n_3152, n_3342);
  not g11582 (n_3343, n8098);
  not g11583 (n_3344, n8331);
  and g11584 (n8332, n_3343, n_3344);
  not g11585 (n_3345, n8332);
  and g11586 (n8333, n_3137, n_3345);
  not g11587 (n_3346, n8080);
  not g11588 (n_3347, n8333);
  and g11589 (n8334, n_3346, n_3347);
  not g11590 (n_3348, n8334);
  and g11591 (n8335, n_3122, n_3348);
  not g11592 (n_3349, n8062);
  not g11593 (n_3350, n8335);
  and g11594 (n8336, n_3349, n_3350);
  not g11595 (n_3351, n8336);
  and g11596 (n8337, n_3107, n_3351);
  not g11597 (n_3352, n7927);
  and g11598 (n8338, n7925, n_3352);
  not g11599 (n_3353, n8338);
  and g11600 (n8339, n_2998, n_3353);
  not g11601 (n_3354, n8337);
  and g11602 (n8340, n_3354, n8339);
  and g11603 (n8341, n_293, n5496);
  and g11604 (n8342, n_298, n4935);
  and g11605 (n8343, n_295, n5407);
  and g11611 (n8346, n4861, n4938);
  not g11614 (n_3359, n8347);
  and g11615 (n8348, \a[20] , n_3359);
  not g11616 (n_3360, n8348);
  and g11617 (n8349, n_3359, n_3360);
  and g11618 (n8350, \a[20] , n_3360);
  not g11619 (n_3361, n8349);
  not g11620 (n_3362, n8350);
  and g11621 (n8351, n_3361, n_3362);
  not g11622 (n_3363, n8339);
  and g11623 (n8352, n8337, n_3363);
  not g11624 (n_3364, n8340);
  not g11625 (n_3365, n8352);
  and g11626 (n8353, n_3364, n_3365);
  not g11627 (n_3366, n8351);
  and g11628 (n8354, n_3366, n8353);
  not g11629 (n_3367, n8354);
  and g11630 (n8355, n_3364, n_3367);
  not g11631 (n_3368, n8044);
  not g11632 (n_3369, n8355);
  and g11633 (n8356, n_3368, n_3369);
  and g11634 (n8357, n8044, n8355);
  not g11635 (n_3370, n8356);
  not g11636 (n_3371, n8357);
  and g11637 (n8358, n_3370, n_3371);
  and g11638 (n8359, n_260, n6233);
  and g11639 (n8360, n_281, n5663);
  and g11640 (n8361, n_275, n5939);
  and g11646 (n8364, n4179, n5666);
  not g11649 (n_3376, n8365);
  and g11650 (n8366, \a[17] , n_3376);
  not g11651 (n_3377, n8366);
  and g11652 (n8367, \a[17] , n_3377);
  and g11653 (n8368, n_3376, n_3377);
  not g11654 (n_3378, n8367);
  not g11655 (n_3379, n8368);
  and g11656 (n8369, n_3378, n_3379);
  not g11657 (n_3380, n8369);
  and g11658 (n8370, n8358, n_3380);
  not g11659 (n_3381, n8370);
  and g11660 (n8371, n_3370, n_3381);
  not g11661 (n_3382, n8041);
  not g11662 (n_3383, n8371);
  and g11663 (n8372, n_3382, n_3383);
  and g11664 (n8373, n8041, n8371);
  not g11665 (n_3384, n8372);
  not g11666 (n_3385, n8373);
  and g11667 (n8374, n_3384, n_3385);
  and g11668 (n8375, n_484, n7101);
  and g11669 (n8376, n_236, n6402);
  and g11670 (n8377, n_415, n6951);
  and g11676 (n8380, n3715, n6397);
  not g11679 (n_3390, n8381);
  and g11680 (n8382, \a[14] , n_3390);
  not g11681 (n_3391, n8382);
  and g11682 (n8383, \a[14] , n_3391);
  and g11683 (n8384, n_3390, n_3391);
  not g11684 (n_3392, n8383);
  not g11685 (n_3393, n8384);
  and g11686 (n8385, n_3392, n_3393);
  not g11687 (n_3394, n8385);
  and g11688 (n8386, n8374, n_3394);
  not g11689 (n_3395, n8386);
  and g11690 (n8387, n_3384, n_3395);
  not g11691 (n_3396, n8026);
  and g11692 (n8388, n_3396, n8037);
  not g11693 (n_3397, n8038);
  not g11694 (n_3398, n8388);
  and g11695 (n8389, n_3397, n_3398);
  not g11696 (n_3399, n8387);
  and g11697 (n8390, n_3399, n8389);
  not g11698 (n_3400, n8390);
  and g11699 (n8391, n_3397, n_3400);
  not g11700 (n_3401, n8024);
  not g11701 (n_3402, n8391);
  and g11702 (n8392, n_3401, n_3402);
  and g11703 (n8393, n8024, n8391);
  not g11704 (n_3403, n8392);
  not g11705 (n_3404, n8393);
  and g11706 (n8394, n_3403, n_3404);
  and g11707 (n8395, n_566, n7983);
  and g11708 (n8396, n_535, n7291);
  and g11709 (n8397, n_565, n7632);
  and g11715 (n8400, n4477, n7294);
  not g11718 (n_3409, n8401);
  and g11719 (n8402, \a[11] , n_3409);
  not g11720 (n_3410, n8402);
  and g11721 (n8403, \a[11] , n_3410);
  and g11722 (n8404, n_3409, n_3410);
  not g11723 (n_3411, n8403);
  not g11724 (n_3412, n8404);
  and g11725 (n8405, n_3411, n_3412);
  not g11726 (n_3413, n8405);
  and g11727 (n8406, n8394, n_3413);
  not g11728 (n_3414, n8406);
  and g11729 (n8407, n_3403, n_3414);
  not g11730 (n_3416, \a[6] );
  and g11731 (n8408, n_3416, \a[7] );
  not g11732 (n_3418, \a[7] );
  and g11733 (n8409, \a[6] , n_3418);
  not g11734 (n_3419, n8408);
  not g11735 (n_3420, n8409);
  and g11736 (n8410, n_3419, n_3420);
  and g11737 (n8411, \a[7] , n_1106);
  and g11738 (n8412, n_3418, \a[8] );
  not g11739 (n_3421, n8411);
  not g11740 (n_3422, n8412);
  and g11741 (n8413, n_3421, n_3422);
  and g11742 (n8414, \a[5] , n_3416);
  and g11743 (n8415, n_3, \a[6] );
  not g11744 (n_3423, n8414);
  not g11745 (n_3424, n8415);
  and g11746 (n8416, n_3423, n_3424);
  not g11747 (n_3425, n8413);
  and g11748 (n8417, n_3425, n8416);
  and g11749 (n8418, n8410, n8417);
  and g11750 (n8419, n_712, n8418);
  not g11751 (n_3426, n8419);
  and g11752 (n8420, n_729, n_3426);
  not g11753 (n_3427, n8416);
  and g11754 (n8421, n_3425, n_3427);
  not g11755 (n_3428, n8421);
  and g11756 (n8422, n_3426, n_3428);
  not g11757 (n_3429, n8420);
  not g11758 (n_3430, n8422);
  and g11759 (n8423, n_3429, n_3430);
  not g11760 (n_3431, n8423);
  and g11761 (n8424, \a[8] , n_3431);
  and g11762 (n8425, n_1106, n8423);
  not g11763 (n_3432, n8424);
  not g11764 (n_3433, n8425);
  and g11765 (n8426, n_3432, n_3433);
  not g11766 (n_3434, n8407);
  not g11767 (n_3435, n8426);
  and g11768 (n8427, n_3434, n_3435);
  and g11769 (n8428, n7982, n_3057);
  and g11770 (n8429, n_3056, n_3057);
  not g11771 (n_3436, n8428);
  not g11772 (n_3437, n8429);
  and g11773 (n8430, n_3436, n_3437);
  and g11774 (n8431, n8407, n8426);
  not g11775 (n_3438, n8427);
  not g11776 (n_3439, n8431);
  and g11777 (n8432, n_3438, n_3439);
  not g11778 (n_3440, n8430);
  and g11779 (n8433, n_3440, n8432);
  not g11780 (n_3441, n8433);
  and g11781 (n8434, n_3438, n_3441);
  not g11782 (n_3442, n8021);
  not g11783 (n_3443, n8434);
  and g11784 (n8435, n_3442, n_3443);
  and g11785 (n8436, n8021, n8434);
  not g11786 (n_3444, n8435);
  not g11787 (n_3445, n8436);
  and g11788 (n8437, n_3444, n_3445);
  and g11789 (n8438, n_3440, n_3441);
  and g11790 (n8439, n8432, n_3441);
  not g11791 (n_3446, n8438);
  not g11792 (n_3447, n8439);
  and g11793 (n8440, n_3446, n_3447);
  and g11794 (n8441, n8374, n_3395);
  and g11795 (n8442, n_3394, n_3395);
  not g11796 (n_3448, n8441);
  not g11797 (n_3449, n8442);
  and g11798 (n8443, n_3448, n_3449);
  and g11799 (n8444, n8358, n_3381);
  and g11800 (n8445, n_3380, n_3381);
  not g11801 (n_3450, n8444);
  not g11802 (n_3451, n8445);
  and g11803 (n8446, n_3450, n_3451);
  and g11804 (n8447, n8062, n8335);
  not g11805 (n_3452, n8447);
  and g11806 (n8448, n_3351, n_3452);
  and g11807 (n8449, n_295, n5496);
  and g11808 (n8450, n_299, n4935);
  and g11809 (n8451, n_298, n5407);
  not g11810 (n_3453, n8450);
  not g11811 (n_3454, n8451);
  and g11812 (n8452, n_3453, n_3454);
  not g11813 (n_3455, n8449);
  and g11814 (n8453, n_3455, n8452);
  and g11815 (n8454, n_1011, n8453);
  not g11816 (n_3456, n4848);
  and g11817 (n8455, n_3456, n8453);
  not g11818 (n_3457, n8454);
  not g11819 (n_3458, n8455);
  and g11820 (n8456, n_3457, n_3458);
  not g11821 (n_3459, n8456);
  and g11822 (n8457, \a[20] , n_3459);
  and g11823 (n8458, n_435, n8456);
  not g11824 (n_3460, n8457);
  not g11825 (n_3461, n8458);
  and g11826 (n8459, n_3460, n_3461);
  not g11827 (n_3462, n8459);
  and g11828 (n8460, n8448, n_3462);
  and g11829 (n8461, n8080, n8333);
  not g11830 (n_3463, n8461);
  and g11831 (n8462, n_3348, n_3463);
  and g11832 (n8463, n_298, n5496);
  and g11833 (n8464, n_300, n4935);
  and g11834 (n8465, n_299, n5407);
  not g11835 (n_3464, n8464);
  not g11836 (n_3465, n8465);
  and g11837 (n8466, n_3464, n_3465);
  not g11838 (n_3466, n8463);
  and g11839 (n8467, n_3466, n8466);
  and g11840 (n8468, n_1011, n8467);
  and g11841 (n8469, n_1505, n8467);
  not g11842 (n_3467, n8468);
  not g11843 (n_3468, n8469);
  and g11844 (n8470, n_3467, n_3468);
  not g11845 (n_3469, n8470);
  and g11846 (n8471, \a[20] , n_3469);
  and g11847 (n8472, n_435, n8470);
  not g11848 (n_3470, n8471);
  not g11849 (n_3471, n8472);
  and g11850 (n8473, n_3470, n_3471);
  not g11851 (n_3472, n8473);
  and g11852 (n8474, n8462, n_3472);
  and g11853 (n8475, n8098, n8331);
  not g11854 (n_3473, n8475);
  and g11855 (n8476, n_3345, n_3473);
  and g11856 (n8477, n_299, n5496);
  and g11857 (n8478, n_301, n4935);
  and g11858 (n8479, n_300, n5407);
  not g11859 (n_3474, n8478);
  not g11860 (n_3475, n8479);
  and g11861 (n8480, n_3474, n_3475);
  not g11862 (n_3476, n8477);
  and g11863 (n8481, n_3476, n8480);
  and g11864 (n8482, n_1011, n8481);
  and g11865 (n8483, n_2193, n8481);
  not g11866 (n_3477, n8482);
  not g11867 (n_3478, n8483);
  and g11868 (n8484, n_3477, n_3478);
  not g11869 (n_3479, n8484);
  and g11870 (n8485, \a[20] , n_3479);
  and g11871 (n8486, n_435, n8484);
  not g11872 (n_3480, n8485);
  not g11873 (n_3481, n8486);
  and g11874 (n8487, n_3480, n_3481);
  not g11875 (n_3482, n8487);
  and g11876 (n8488, n8476, n_3482);
  and g11877 (n8489, n8116, n8329);
  not g11878 (n_3483, n8489);
  and g11879 (n8490, n_3342, n_3483);
  and g11880 (n8491, n_300, n5496);
  and g11881 (n8492, n_302, n4935);
  and g11882 (n8493, n_301, n5407);
  not g11883 (n_3484, n8492);
  not g11884 (n_3485, n8493);
  and g11885 (n8494, n_3484, n_3485);
  not g11886 (n_3486, n8491);
  and g11887 (n8495, n_3486, n8494);
  and g11888 (n8496, n_1011, n8495);
  and g11889 (n8497, n_1801, n8495);
  not g11890 (n_3487, n8496);
  not g11891 (n_3488, n8497);
  and g11892 (n8498, n_3487, n_3488);
  not g11893 (n_3489, n8498);
  and g11894 (n8499, \a[20] , n_3489);
  and g11895 (n8500, n_435, n8498);
  not g11896 (n_3490, n8499);
  not g11897 (n_3491, n8500);
  and g11898 (n8501, n_3490, n_3491);
  not g11899 (n_3492, n8501);
  and g11900 (n8502, n8490, n_3492);
  and g11901 (n8503, n8134, n8327);
  not g11902 (n_3493, n8503);
  and g11903 (n8504, n_3339, n_3493);
  and g11904 (n8505, n_301, n5496);
  and g11905 (n8506, n_303, n4935);
  and g11906 (n8507, n_302, n5407);
  not g11907 (n_3494, n8506);
  not g11908 (n_3495, n8507);
  and g11909 (n8508, n_3494, n_3495);
  not g11910 (n_3496, n8505);
  and g11911 (n8509, n_3496, n8508);
  and g11912 (n8510, n_1011, n8509);
  and g11913 (n8511, n_1672, n8509);
  not g11914 (n_3497, n8510);
  not g11915 (n_3498, n8511);
  and g11916 (n8512, n_3497, n_3498);
  not g11917 (n_3499, n8512);
  and g11918 (n8513, \a[20] , n_3499);
  and g11919 (n8514, n_435, n8512);
  not g11920 (n_3500, n8513);
  not g11921 (n_3501, n8514);
  and g11922 (n8515, n_3500, n_3501);
  not g11923 (n_3502, n8515);
  and g11924 (n8516, n8504, n_3502);
  and g11925 (n8517, n8152, n8325);
  not g11926 (n_3503, n8517);
  and g11927 (n8518, n_3336, n_3503);
  and g11928 (n8519, n_302, n5496);
  and g11929 (n8520, n_304, n4935);
  and g11930 (n8521, n_303, n5407);
  not g11931 (n_3504, n8520);
  not g11932 (n_3505, n8521);
  and g11933 (n8522, n_3504, n_3505);
  not g11934 (n_3506, n8519);
  and g11935 (n8523, n_3506, n8522);
  and g11936 (n8524, n_1011, n8523);
  not g11937 (n_3507, n5851);
  and g11938 (n8525, n_3507, n8523);
  not g11939 (n_3508, n8524);
  not g11940 (n_3509, n8525);
  and g11941 (n8526, n_3508, n_3509);
  not g11942 (n_3510, n8526);
  and g11943 (n8527, \a[20] , n_3510);
  and g11944 (n8528, n_435, n8526);
  not g11945 (n_3511, n8527);
  not g11946 (n_3512, n8528);
  and g11947 (n8529, n_3511, n_3512);
  not g11948 (n_3513, n8529);
  and g11949 (n8530, n8518, n_3513);
  and g11950 (n8531, n8170, n8323);
  not g11951 (n_3514, n8531);
  and g11952 (n8532, n_3333, n_3514);
  and g11953 (n8533, n_303, n5496);
  and g11954 (n8534, n_305, n4935);
  and g11955 (n8535, n_304, n5407);
  not g11956 (n_3515, n8534);
  not g11957 (n_3516, n8535);
  and g11958 (n8536, n_3515, n_3516);
  not g11959 (n_3517, n8533);
  and g11960 (n8537, n_3517, n8536);
  and g11961 (n8538, n_1011, n8537);
  and g11962 (n8539, n_2206, n8537);
  not g11963 (n_3518, n8538);
  not g11964 (n_3519, n8539);
  and g11965 (n8540, n_3518, n_3519);
  not g11966 (n_3520, n8540);
  and g11967 (n8541, \a[20] , n_3520);
  and g11968 (n8542, n_435, n8540);
  not g11969 (n_3521, n8541);
  not g11970 (n_3522, n8542);
  and g11971 (n8543, n_3521, n_3522);
  not g11972 (n_3523, n8543);
  and g11973 (n8544, n8532, n_3523);
  and g11974 (n8545, n_304, n5496);
  and g11975 (n8546, n_306, n4935);
  and g11976 (n8547, n_305, n5407);
  and g11982 (n8550, n4938, n5834);
  not g11985 (n_3528, n8551);
  and g11986 (n8552, \a[20] , n_3528);
  not g11987 (n_3529, n8552);
  and g11988 (n8553, n_3528, n_3529);
  and g11989 (n8554, \a[20] , n_3529);
  not g11990 (n_3530, n8553);
  not g11991 (n_3531, n8554);
  and g11992 (n8555, n_3530, n_3531);
  not g11993 (n_3532, n8321);
  and g11994 (n8556, n8319, n_3532);
  not g11995 (n_3533, n8556);
  and g11996 (n8557, n_3330, n_3533);
  not g11997 (n_3534, n8555);
  and g11998 (n8558, n_3534, n8557);
  not g11999 (n_3535, n8558);
  and g12000 (n8559, n_3534, n_3535);
  and g12001 (n8560, n8557, n_3535);
  not g12002 (n_3536, n8559);
  not g12003 (n_3537, n8560);
  and g12004 (n8561, n_3536, n_3537);
  and g12005 (n8562, n_305, n5496);
  and g12006 (n8563, n_307, n4935);
  and g12007 (n8564, n_306, n5407);
  and g12013 (n8567, n4938, n6143);
  not g12016 (n_3542, n8568);
  and g12017 (n8569, \a[20] , n_3542);
  not g12018 (n_3543, n8569);
  and g12019 (n8570, n_3542, n_3543);
  and g12020 (n8571, \a[20] , n_3543);
  not g12021 (n_3544, n8570);
  not g12022 (n_3545, n8571);
  and g12023 (n8572, n_3544, n_3545);
  and g12024 (n8573, n_3323, n_3325);
  and g12025 (n8574, n_3324, n_3325);
  not g12026 (n_3546, n8573);
  not g12027 (n_3547, n8574);
  and g12028 (n8575, n_3546, n_3547);
  not g12029 (n_3548, n8572);
  not g12030 (n_3549, n8575);
  and g12031 (n8576, n_3548, n_3549);
  not g12032 (n_3550, n8576);
  and g12033 (n8577, n_3548, n_3550);
  and g12034 (n8578, n_3549, n_3550);
  not g12035 (n_3551, n8577);
  not g12036 (n_3552, n8578);
  and g12037 (n8579, n_3551, n_3552);
  and g12038 (n8580, n8215, n8312);
  not g12039 (n_3553, n8580);
  and g12040 (n8581, n_3319, n_3553);
  and g12041 (n8582, n_306, n5496);
  and g12042 (n8583, n_308, n4935);
  and g12043 (n8584, n_307, n5407);
  not g12044 (n_3554, n8583);
  not g12045 (n_3555, n8584);
  and g12046 (n8585, n_3554, n_3555);
  not g12047 (n_3556, n8582);
  and g12048 (n8586, n_3556, n8585);
  and g12049 (n8587, n_1011, n8586);
  and g12050 (n8588, n_2498, n8586);
  not g12051 (n_3557, n8587);
  not g12052 (n_3558, n8588);
  and g12053 (n8589, n_3557, n_3558);
  not g12054 (n_3559, n8589);
  and g12055 (n8590, \a[20] , n_3559);
  and g12056 (n8591, n_435, n8589);
  not g12057 (n_3560, n8590);
  not g12058 (n_3561, n8591);
  and g12059 (n8592, n_3560, n_3561);
  not g12060 (n_3562, n8592);
  and g12061 (n8593, n8581, n_3562);
  not g12062 (n_3563, n8310);
  and g12063 (n8594, n8308, n_3563);
  not g12064 (n_3564, n8594);
  and g12065 (n8595, n_3316, n_3564);
  and g12066 (n8596, n_307, n5496);
  and g12067 (n8597, n_309, n4935);
  and g12068 (n8598, n_308, n5407);
  not g12069 (n_3565, n8597);
  not g12070 (n_3566, n8598);
  and g12071 (n8599, n_3565, n_3566);
  not g12072 (n_3567, n8596);
  and g12073 (n8600, n_3567, n8599);
  and g12074 (n8601, n_1011, n8600);
  and g12075 (n8602, n_2511, n8600);
  not g12076 (n_3568, n8601);
  not g12077 (n_3569, n8602);
  and g12078 (n8603, n_3568, n_3569);
  not g12079 (n_3570, n8603);
  and g12080 (n8604, \a[20] , n_3570);
  and g12081 (n8605, n_435, n8603);
  not g12082 (n_3571, n8604);
  not g12083 (n_3572, n8605);
  and g12084 (n8606, n_3571, n_3572);
  not g12085 (n_3573, n8606);
  and g12086 (n8607, n8595, n_3573);
  and g12087 (n8608, n8247, n8306);
  not g12088 (n_3574, n8608);
  and g12089 (n8609, n_3312, n_3574);
  and g12090 (n8610, n_308, n5496);
  and g12091 (n8611, n_310, n4935);
  and g12092 (n8612, n_309, n5407);
  not g12093 (n_3575, n8611);
  not g12094 (n_3576, n8612);
  and g12095 (n8613, n_3575, n_3576);
  not g12096 (n_3577, n8610);
  and g12097 (n8614, n_3577, n8613);
  and g12098 (n8615, n_1011, n8614);
  and g12099 (n8616, n_2839, n8614);
  not g12100 (n_3578, n8615);
  not g12101 (n_3579, n8616);
  and g12102 (n8617, n_3578, n_3579);
  not g12103 (n_3580, n8617);
  and g12104 (n8618, \a[20] , n_3580);
  and g12105 (n8619, n_435, n8617);
  not g12106 (n_3581, n8618);
  not g12107 (n_3582, n8619);
  and g12108 (n8620, n_3581, n_3582);
  not g12109 (n_3583, n8620);
  and g12110 (n8621, n8609, n_3583);
  and g12111 (n8622, n_309, n5496);
  and g12112 (n8623, n_311, n4935);
  and g12113 (n8624, n_310, n5407);
  and g12119 (n8627, n4938, n6541);
  not g12122 (n_3588, n8628);
  and g12123 (n8629, \a[20] , n_3588);
  not g12124 (n_3589, n8629);
  and g12125 (n8630, n_3588, n_3589);
  and g12126 (n8631, \a[20] , n_3589);
  not g12127 (n_3590, n8630);
  not g12128 (n_3591, n8631);
  and g12129 (n8632, n_3590, n_3591);
  not g12130 (n_3592, n8304);
  and g12131 (n8633, n8302, n_3592);
  not g12132 (n_3593, n8633);
  and g12133 (n8634, n_3309, n_3593);
  not g12134 (n_3594, n8632);
  and g12135 (n8635, n_3594, n8634);
  not g12136 (n_3595, n8635);
  and g12137 (n8636, n_3594, n_3595);
  and g12138 (n8637, n8634, n_3595);
  not g12139 (n_3596, n8636);
  not g12140 (n_3597, n8637);
  and g12141 (n8638, n_3596, n_3597);
  and g12142 (n8639, n_3302, n_3304);
  and g12143 (n8640, n_3303, n_3304);
  not g12144 (n_3598, n8639);
  not g12145 (n_3599, n8640);
  and g12146 (n8641, n_3598, n_3599);
  and g12147 (n8642, n_310, n5496);
  and g12148 (n8643, n_312, n4935);
  and g12149 (n8644, n_311, n5407);
  not g12150 (n_3600, n8643);
  not g12151 (n_3601, n8644);
  and g12152 (n8645, n_3600, n_3601);
  not g12153 (n_3602, n8642);
  and g12154 (n8646, n_3602, n8645);
  and g12155 (n8647, n_1011, n8646);
  and g12156 (n8648, n_3239, n8646);
  not g12157 (n_3603, n8647);
  not g12158 (n_3604, n8648);
  and g12159 (n8649, n_3603, n_3604);
  not g12160 (n_3605, n8649);
  and g12161 (n8650, \a[20] , n_3605);
  and g12162 (n8651, n_435, n8649);
  not g12163 (n_3606, n8650);
  not g12164 (n_3607, n8651);
  and g12165 (n8652, n_3606, n_3607);
  not g12166 (n_3608, n8641);
  not g12167 (n_3609, n8652);
  and g12168 (n8653, n_3608, n_3609);
  and g12169 (n8654, n_311, n5496);
  and g12170 (n8655, n_313, n4935);
  and g12171 (n8656, n_312, n5407);
  and g12177 (n8659, n4938, n6646);
  not g12180 (n_3614, n8660);
  and g12181 (n8661, \a[20] , n_3614);
  not g12182 (n_3615, n8661);
  and g12183 (n8662, n_3614, n_3615);
  and g12184 (n8663, \a[20] , n_3615);
  not g12185 (n_3616, n8662);
  not g12186 (n_3617, n8663);
  and g12187 (n8664, n_3616, n_3617);
  not g12188 (n_3618, n8273);
  and g12189 (n8665, n_3618, n8284);
  not g12190 (n_3619, n8285);
  not g12191 (n_3620, n8665);
  and g12192 (n8666, n_3619, n_3620);
  not g12193 (n_3621, n8664);
  and g12194 (n8667, n_3621, n8666);
  not g12195 (n_3622, n8667);
  and g12196 (n8668, n_3621, n_3622);
  and g12197 (n8669, n8666, n_3622);
  not g12198 (n_3623, n8668);
  not g12199 (n_3624, n8669);
  and g12200 (n8670, n_3623, n_3624);
  not g12201 (n_3625, n8272);
  and g12202 (n8671, n8270, n_3625);
  not g12203 (n_3626, n8671);
  and g12204 (n8672, n_3618, n_3626);
  and g12205 (n8673, n_312, n5496);
  and g12206 (n8674, n_314, n4935);
  and g12207 (n8675, n_313, n5407);
  not g12208 (n_3627, n8674);
  not g12209 (n_3628, n8675);
  and g12210 (n8676, n_3627, n_3628);
  not g12211 (n_3629, n8673);
  and g12212 (n8677, n_3629, n8676);
  and g12213 (n8678, n_1011, n8677);
  and g12214 (n8679, n_2891, n8677);
  not g12215 (n_3630, n8678);
  not g12216 (n_3631, n8679);
  and g12217 (n8680, n_3630, n_3631);
  not g12218 (n_3632, n8680);
  and g12219 (n8681, \a[20] , n_3632);
  and g12220 (n8682, n_435, n8680);
  not g12221 (n_3633, n8681);
  not g12222 (n_3634, n8682);
  and g12223 (n8683, n_3633, n_3634);
  not g12224 (n_3635, n8683);
  and g12225 (n8684, n8672, n_3635);
  and g12226 (n8685, n_316, n5407);
  and g12227 (n8686, n_315, n5496);
  not g12228 (n_3636, n8685);
  not g12229 (n_3637, n8686);
  and g12230 (n8687, n_3636, n_3637);
  and g12231 (n8688, n4938, n_2588);
  not g12232 (n_3638, n8688);
  and g12233 (n8689, n8687, n_3638);
  not g12234 (n_3639, n8689);
  and g12235 (n8690, \a[20] , n_3639);
  not g12236 (n_3640, n8690);
  and g12237 (n8691, \a[20] , n_3640);
  and g12238 (n8692, n_3639, n_3640);
  not g12239 (n_3641, n8691);
  not g12240 (n_3642, n8692);
  and g12241 (n8693, n_3641, n_3642);
  and g12242 (n8694, n_316, n_1010);
  not g12243 (n_3643, n8694);
  and g12244 (n8695, \a[20] , n_3643);
  not g12245 (n_3644, n8693);
  and g12246 (n8696, n_3644, n8695);
  and g12247 (n8697, n_314, n5496);
  and g12248 (n8698, n_316, n4935);
  and g12249 (n8699, n_315, n5407);
  not g12250 (n_3645, n8698);
  not g12251 (n_3646, n8699);
  and g12252 (n8700, n_3645, n_3646);
  not g12253 (n_3647, n8697);
  and g12254 (n8701, n_3647, n8700);
  and g12255 (n8702, n_1011, n8701);
  and g12256 (n8703, n_2612, n8701);
  not g12257 (n_3648, n8702);
  not g12258 (n_3649, n8703);
  and g12259 (n8704, n_3648, n_3649);
  not g12260 (n_3650, n8704);
  and g12261 (n8705, \a[20] , n_3650);
  and g12262 (n8706, n_435, n8704);
  not g12263 (n_3651, n8705);
  not g12264 (n_3652, n8706);
  and g12265 (n8707, n_3651, n_3652);
  not g12266 (n_3653, n8707);
  and g12267 (n8708, n8696, n_3653);
  and g12268 (n8709, n8271, n8708);
  not g12269 (n_3654, n8709);
  and g12270 (n8710, n8708, n_3654);
  and g12271 (n8711, n8271, n_3654);
  not g12272 (n_3655, n8710);
  not g12273 (n_3656, n8711);
  and g12274 (n8712, n_3655, n_3656);
  and g12275 (n8713, n_313, n5496);
  and g12276 (n8714, n_315, n4935);
  and g12277 (n8715, n_314, n5407);
  and g12283 (n8718, n4938, n6806);
  not g12286 (n_3661, n8719);
  and g12287 (n8720, \a[20] , n_3661);
  not g12288 (n_3662, n8720);
  and g12289 (n8721, \a[20] , n_3662);
  and g12290 (n8722, n_3661, n_3662);
  not g12291 (n_3663, n8721);
  not g12292 (n_3664, n8722);
  and g12293 (n8723, n_3663, n_3664);
  not g12294 (n_3665, n8712);
  not g12295 (n_3666, n8723);
  and g12296 (n8724, n_3665, n_3666);
  not g12297 (n_3667, n8724);
  and g12298 (n8725, n_3654, n_3667);
  not g12299 (n_3668, n8672);
  and g12300 (n8726, n_3668, n8683);
  not g12301 (n_3669, n8684);
  not g12302 (n_3670, n8726);
  and g12303 (n8727, n_3669, n_3670);
  not g12304 (n_3671, n8725);
  and g12305 (n8728, n_3671, n8727);
  not g12306 (n_3672, n8728);
  and g12307 (n8729, n_3669, n_3672);
  not g12308 (n_3673, n8670);
  not g12309 (n_3674, n8729);
  and g12310 (n8730, n_3673, n_3674);
  not g12311 (n_3675, n8730);
  and g12312 (n8731, n_3622, n_3675);
  and g12313 (n8732, n8641, n8652);
  not g12314 (n_3676, n8653);
  not g12315 (n_3677, n8732);
  and g12316 (n8733, n_3676, n_3677);
  not g12317 (n_3678, n8731);
  and g12318 (n8734, n_3678, n8733);
  not g12319 (n_3679, n8734);
  and g12320 (n8735, n_3676, n_3679);
  not g12321 (n_3680, n8638);
  not g12322 (n_3681, n8735);
  and g12323 (n8736, n_3680, n_3681);
  not g12324 (n_3682, n8736);
  and g12325 (n8737, n_3595, n_3682);
  not g12326 (n_3683, n8621);
  and g12327 (n8738, n8609, n_3683);
  and g12328 (n8739, n_3583, n_3683);
  not g12329 (n_3684, n8738);
  not g12330 (n_3685, n8739);
  and g12331 (n8740, n_3684, n_3685);
  not g12332 (n_3686, n8737);
  not g12333 (n_3687, n8740);
  and g12334 (n8741, n_3686, n_3687);
  not g12335 (n_3688, n8741);
  and g12336 (n8742, n_3683, n_3688);
  not g12337 (n_3689, n8607);
  and g12338 (n8743, n8595, n_3689);
  and g12339 (n8744, n_3573, n_3689);
  not g12340 (n_3690, n8743);
  not g12341 (n_3691, n8744);
  and g12342 (n8745, n_3690, n_3691);
  not g12343 (n_3692, n8742);
  not g12344 (n_3693, n8745);
  and g12345 (n8746, n_3692, n_3693);
  not g12346 (n_3694, n8746);
  and g12347 (n8747, n_3689, n_3694);
  not g12348 (n_3695, n8581);
  and g12349 (n8748, n_3695, n8592);
  not g12350 (n_3696, n8593);
  not g12351 (n_3697, n8748);
  and g12352 (n8749, n_3696, n_3697);
  not g12353 (n_3698, n8747);
  and g12354 (n8750, n_3698, n8749);
  not g12355 (n_3699, n8750);
  and g12356 (n8751, n_3696, n_3699);
  not g12357 (n_3700, n8579);
  not g12358 (n_3701, n8751);
  and g12359 (n8752, n_3700, n_3701);
  not g12360 (n_3702, n8752);
  and g12361 (n8753, n_3550, n_3702);
  not g12362 (n_3703, n8561);
  not g12363 (n_3704, n8753);
  and g12364 (n8754, n_3703, n_3704);
  not g12365 (n_3705, n8754);
  and g12366 (n8755, n_3535, n_3705);
  not g12367 (n_3706, n8544);
  and g12368 (n8756, n8532, n_3706);
  and g12369 (n8757, n_3523, n_3706);
  not g12370 (n_3707, n8756);
  not g12371 (n_3708, n8757);
  and g12372 (n8758, n_3707, n_3708);
  not g12373 (n_3709, n8755);
  not g12374 (n_3710, n8758);
  and g12375 (n8759, n_3709, n_3710);
  not g12376 (n_3711, n8759);
  and g12377 (n8760, n_3706, n_3711);
  not g12378 (n_3712, n8530);
  and g12379 (n8761, n8518, n_3712);
  and g12380 (n8762, n_3513, n_3712);
  not g12381 (n_3713, n8761);
  not g12382 (n_3714, n8762);
  and g12383 (n8763, n_3713, n_3714);
  not g12384 (n_3715, n8760);
  not g12385 (n_3716, n8763);
  and g12386 (n8764, n_3715, n_3716);
  not g12387 (n_3717, n8764);
  and g12388 (n8765, n_3712, n_3717);
  not g12389 (n_3718, n8516);
  and g12390 (n8766, n8504, n_3718);
  and g12391 (n8767, n_3502, n_3718);
  not g12392 (n_3719, n8766);
  not g12393 (n_3720, n8767);
  and g12394 (n8768, n_3719, n_3720);
  not g12395 (n_3721, n8765);
  not g12396 (n_3722, n8768);
  and g12397 (n8769, n_3721, n_3722);
  not g12398 (n_3723, n8769);
  and g12399 (n8770, n_3718, n_3723);
  not g12400 (n_3724, n8502);
  and g12401 (n8771, n8490, n_3724);
  and g12402 (n8772, n_3492, n_3724);
  not g12403 (n_3725, n8771);
  not g12404 (n_3726, n8772);
  and g12405 (n8773, n_3725, n_3726);
  not g12406 (n_3727, n8770);
  not g12407 (n_3728, n8773);
  and g12408 (n8774, n_3727, n_3728);
  not g12409 (n_3729, n8774);
  and g12410 (n8775, n_3724, n_3729);
  not g12411 (n_3730, n8488);
  and g12412 (n8776, n8476, n_3730);
  and g12413 (n8777, n_3482, n_3730);
  not g12414 (n_3731, n8776);
  not g12415 (n_3732, n8777);
  and g12416 (n8778, n_3731, n_3732);
  not g12417 (n_3733, n8775);
  not g12418 (n_3734, n8778);
  and g12419 (n8779, n_3733, n_3734);
  not g12420 (n_3735, n8779);
  and g12421 (n8780, n_3730, n_3735);
  not g12422 (n_3736, n8474);
  and g12423 (n8781, n8462, n_3736);
  and g12424 (n8782, n_3472, n_3736);
  not g12425 (n_3737, n8781);
  not g12426 (n_3738, n8782);
  and g12427 (n8783, n_3737, n_3738);
  not g12428 (n_3739, n8780);
  not g12429 (n_3740, n8783);
  and g12430 (n8784, n_3739, n_3740);
  not g12431 (n_3741, n8784);
  and g12432 (n8785, n_3736, n_3741);
  not g12433 (n_3742, n8460);
  and g12434 (n8786, n8448, n_3742);
  and g12435 (n8787, n_3462, n_3742);
  not g12436 (n_3743, n8786);
  not g12437 (n_3744, n8787);
  and g12438 (n8788, n_3743, n_3744);
  not g12439 (n_3745, n8785);
  not g12440 (n_3746, n8788);
  and g12441 (n8789, n_3745, n_3746);
  not g12442 (n_3747, n8789);
  and g12443 (n8790, n_3742, n_3747);
  not g12444 (n_3748, n8353);
  and g12445 (n8791, n8351, n_3748);
  not g12446 (n_3749, n8791);
  and g12447 (n8792, n_3367, n_3749);
  not g12448 (n_3750, n8790);
  and g12449 (n8793, n_3750, n8792);
  and g12450 (n8794, n_275, n6233);
  and g12451 (n8795, n_286, n5663);
  and g12452 (n8796, n_281, n5939);
  and g12458 (n8799, n4204, n5666);
  not g12461 (n_3755, n8800);
  and g12462 (n8801, \a[17] , n_3755);
  not g12463 (n_3756, n8801);
  and g12464 (n8802, n_3755, n_3756);
  and g12465 (n8803, \a[17] , n_3756);
  not g12466 (n_3757, n8802);
  not g12467 (n_3758, n8803);
  and g12468 (n8804, n_3757, n_3758);
  not g12469 (n_3759, n8792);
  and g12470 (n8805, n8790, n_3759);
  not g12471 (n_3760, n8793);
  not g12472 (n_3761, n8805);
  and g12473 (n8806, n_3760, n_3761);
  not g12474 (n_3762, n8804);
  and g12475 (n8807, n_3762, n8806);
  not g12476 (n_3763, n8807);
  and g12477 (n8808, n_3760, n_3763);
  not g12478 (n_3764, n8446);
  not g12479 (n_3765, n8808);
  and g12480 (n8809, n_3764, n_3765);
  and g12481 (n8810, n8446, n8808);
  not g12482 (n_3766, n8809);
  not g12483 (n_3767, n8810);
  and g12484 (n8811, n_3766, n_3767);
  and g12485 (n8812, n_415, n7101);
  and g12486 (n8813, n_237, n6402);
  and g12487 (n8814, n_236, n6951);
  and g12493 (n8817, n3018, n6397);
  not g12496 (n_3772, n8818);
  and g12497 (n8819, \a[14] , n_3772);
  not g12498 (n_3773, n8819);
  and g12499 (n8820, \a[14] , n_3773);
  and g12500 (n8821, n_3772, n_3773);
  not g12501 (n_3774, n8820);
  not g12502 (n_3775, n8821);
  and g12503 (n8822, n_3774, n_3775);
  not g12504 (n_3776, n8822);
  and g12505 (n8823, n8811, n_3776);
  not g12506 (n_3777, n8823);
  and g12507 (n8824, n_3766, n_3777);
  not g12508 (n_3778, n8443);
  not g12509 (n_3779, n8824);
  and g12510 (n8825, n_3778, n_3779);
  and g12511 (n8826, n8443, n8824);
  not g12512 (n_3780, n8825);
  not g12513 (n_3781, n8826);
  and g12514 (n8827, n_3780, n_3781);
  and g12515 (n8828, n_535, n7983);
  and g12516 (n8829, n_485, n7291);
  and g12517 (n8830, n_480, n7632);
  and g12523 (n8833, n3818, n7294);
  not g12526 (n_3786, n8834);
  and g12527 (n8835, \a[11] , n_3786);
  not g12528 (n_3787, n8835);
  and g12529 (n8836, \a[11] , n_3787);
  and g12530 (n8837, n_3786, n_3787);
  not g12531 (n_3788, n8836);
  not g12532 (n_3789, n8837);
  and g12533 (n8838, n_3788, n_3789);
  not g12534 (n_3790, n8838);
  and g12535 (n8839, n8827, n_3790);
  not g12536 (n_3791, n8839);
  and g12537 (n8840, n_3780, n_3791);
  and g12538 (n8841, n_565, n7983);
  and g12539 (n8842, n_480, n7291);
  and g12540 (n8843, n_535, n7632);
  not g12541 (n_3792, n8842);
  not g12542 (n_3793, n8843);
  and g12543 (n8844, n_3792, n_3793);
  not g12544 (n_3794, n8841);
  and g12545 (n8845, n_3794, n8844);
  and g12546 (n8846, n_2446, n8845);
  and g12547 (n8847, n_753, n8845);
  not g12548 (n_3795, n8846);
  not g12549 (n_3796, n8847);
  and g12550 (n8848, n_3795, n_3796);
  not g12551 (n_3797, n8848);
  and g12552 (n8849, \a[11] , n_3797);
  and g12553 (n8850, n_1071, n8848);
  not g12554 (n_3798, n8849);
  not g12555 (n_3799, n8850);
  and g12556 (n8851, n_3798, n_3799);
  not g12557 (n_3800, n8840);
  not g12558 (n_3801, n8851);
  and g12559 (n8852, n_3800, n_3801);
  and g12560 (n8853, n8840, n8851);
  not g12561 (n_3802, n8852);
  not g12562 (n_3803, n8853);
  and g12563 (n8854, n_3802, n_3803);
  not g12564 (n_3804, n8389);
  and g12565 (n8855, n8387, n_3804);
  not g12566 (n_3805, n8855);
  and g12567 (n8856, n_3400, n_3805);
  and g12568 (n8857, n8854, n8856);
  not g12569 (n_3806, n8857);
  and g12570 (n8858, n_3802, n_3806);
  and g12571 (n8859, n_560, n8418);
  not g12572 (n_3807, n8410);
  and g12573 (n8860, n_3807, n8416);
  and g12574 (n8861, n_712, n8860);
  not g12575 (n_3808, n8859);
  not g12576 (n_3809, n8861);
  and g12577 (n8862, n_3808, n_3809);
  and g12578 (n8863, n_3428, n8862);
  and g12579 (n8864, n_2152, n8862);
  not g12580 (n_3810, n8863);
  not g12581 (n_3811, n8864);
  and g12582 (n8865, n_3810, n_3811);
  not g12583 (n_3812, n8865);
  and g12584 (n8866, \a[8] , n_3812);
  and g12585 (n8867, n_1106, n8865);
  not g12586 (n_3813, n8866);
  not g12587 (n_3814, n8867);
  and g12588 (n8868, n_3813, n_3814);
  not g12589 (n_3815, n8858);
  not g12590 (n_3816, n8868);
  and g12591 (n8869, n_3815, n_3816);
  and g12592 (n8870, n8394, n_3414);
  and g12593 (n8871, n_3413, n_3414);
  not g12594 (n_3817, n8870);
  not g12595 (n_3818, n8871);
  and g12596 (n8872, n_3817, n_3818);
  and g12597 (n8873, n8858, n8868);
  not g12598 (n_3819, n8869);
  not g12599 (n_3820, n8873);
  and g12600 (n8874, n_3819, n_3820);
  not g12601 (n_3821, n8872);
  and g12602 (n8875, n_3821, n8874);
  not g12603 (n_3822, n8875);
  and g12604 (n8876, n_3819, n_3822);
  not g12605 (n_3823, n8440);
  not g12606 (n_3824, n8876);
  and g12607 (n8877, n_3823, n_3824);
  and g12608 (n8878, n8440, n8876);
  not g12609 (n_3825, n8877);
  not g12610 (n_3826, n8878);
  and g12611 (n8879, n_3825, n_3826);
  and g12612 (n8880, n8827, n_3791);
  and g12613 (n8881, n_3790, n_3791);
  not g12614 (n_3827, n8880);
  not g12615 (n_3828, n8881);
  and g12616 (n8882, n_3827, n_3828);
  and g12617 (n8883, n8811, n_3777);
  and g12618 (n8884, n_3776, n_3777);
  not g12619 (n_3829, n8883);
  not g12620 (n_3830, n8884);
  and g12621 (n8885, n_3829, n_3830);
  and g12622 (n8886, n_281, n6233);
  and g12623 (n8887, n_293, n5663);
  and g12624 (n8888, n_286, n5939);
  and g12630 (n8891, n4633, n5666);
  not g12633 (n_3835, n8892);
  and g12634 (n8893, \a[17] , n_3835);
  not g12635 (n_3836, n8893);
  and g12636 (n8894, n_3835, n_3836);
  and g12637 (n8895, \a[17] , n_3836);
  not g12638 (n_3837, n8894);
  not g12639 (n_3838, n8895);
  and g12640 (n8896, n_3837, n_3838);
  and g12641 (n8897, n_3745, n_3747);
  and g12642 (n8898, n_3746, n_3747);
  not g12643 (n_3839, n8897);
  not g12644 (n_3840, n8898);
  and g12645 (n8899, n_3839, n_3840);
  not g12646 (n_3841, n8896);
  not g12647 (n_3842, n8899);
  and g12648 (n8900, n_3841, n_3842);
  not g12649 (n_3843, n8900);
  and g12650 (n8901, n_3841, n_3843);
  and g12651 (n8902, n_3842, n_3843);
  not g12652 (n_3844, n8901);
  not g12653 (n_3845, n8902);
  and g12654 (n8903, n_3844, n_3845);
  and g12655 (n8904, n_286, n6233);
  and g12656 (n8905, n_295, n5663);
  and g12657 (n8906, n_293, n5939);
  and g12663 (n8909, n4429, n5666);
  not g12666 (n_3850, n8910);
  and g12667 (n8911, \a[17] , n_3850);
  not g12668 (n_3851, n8911);
  and g12669 (n8912, n_3850, n_3851);
  and g12670 (n8913, \a[17] , n_3851);
  not g12671 (n_3852, n8912);
  not g12672 (n_3853, n8913);
  and g12673 (n8914, n_3852, n_3853);
  and g12674 (n8915, n_3739, n_3741);
  and g12675 (n8916, n_3740, n_3741);
  not g12676 (n_3854, n8915);
  not g12677 (n_3855, n8916);
  and g12678 (n8917, n_3854, n_3855);
  not g12679 (n_3856, n8914);
  not g12680 (n_3857, n8917);
  and g12681 (n8918, n_3856, n_3857);
  not g12682 (n_3858, n8918);
  and g12683 (n8919, n_3856, n_3858);
  and g12684 (n8920, n_3857, n_3858);
  not g12685 (n_3859, n8919);
  not g12686 (n_3860, n8920);
  and g12687 (n8921, n_3859, n_3860);
  and g12688 (n8922, n_293, n6233);
  and g12689 (n8923, n_298, n5663);
  and g12690 (n8924, n_295, n5939);
  and g12696 (n8927, n4861, n5666);
  not g12699 (n_3865, n8928);
  and g12700 (n8929, \a[17] , n_3865);
  not g12701 (n_3866, n8929);
  and g12702 (n8930, n_3865, n_3866);
  and g12703 (n8931, \a[17] , n_3866);
  not g12704 (n_3867, n8930);
  not g12705 (n_3868, n8931);
  and g12706 (n8932, n_3867, n_3868);
  and g12707 (n8933, n_3733, n_3735);
  and g12708 (n8934, n_3734, n_3735);
  not g12709 (n_3869, n8933);
  not g12710 (n_3870, n8934);
  and g12711 (n8935, n_3869, n_3870);
  not g12712 (n_3871, n8932);
  not g12713 (n_3872, n8935);
  and g12714 (n8936, n_3871, n_3872);
  not g12715 (n_3873, n8936);
  and g12716 (n8937, n_3871, n_3873);
  and g12717 (n8938, n_3872, n_3873);
  not g12718 (n_3874, n8937);
  not g12719 (n_3875, n8938);
  and g12720 (n8939, n_3874, n_3875);
  and g12721 (n8940, n_295, n6233);
  and g12722 (n8941, n_299, n5663);
  and g12723 (n8942, n_298, n5939);
  and g12729 (n8945, n4848, n5666);
  not g12732 (n_3880, n8946);
  and g12733 (n8947, \a[17] , n_3880);
  not g12734 (n_3881, n8947);
  and g12735 (n8948, n_3880, n_3881);
  and g12736 (n8949, \a[17] , n_3881);
  not g12737 (n_3882, n8948);
  not g12738 (n_3883, n8949);
  and g12739 (n8950, n_3882, n_3883);
  and g12740 (n8951, n_3727, n_3729);
  and g12741 (n8952, n_3728, n_3729);
  not g12742 (n_3884, n8951);
  not g12743 (n_3885, n8952);
  and g12744 (n8953, n_3884, n_3885);
  not g12745 (n_3886, n8950);
  not g12746 (n_3887, n8953);
  and g12747 (n8954, n_3886, n_3887);
  not g12748 (n_3888, n8954);
  and g12749 (n8955, n_3886, n_3888);
  and g12750 (n8956, n_3887, n_3888);
  not g12751 (n_3889, n8955);
  not g12752 (n_3890, n8956);
  and g12753 (n8957, n_3889, n_3890);
  and g12754 (n8958, n_298, n6233);
  and g12755 (n8959, n_300, n5663);
  and g12756 (n8960, n_299, n5939);
  and g12762 (n8963, n5114, n5666);
  not g12765 (n_3895, n8964);
  and g12766 (n8965, \a[17] , n_3895);
  not g12767 (n_3896, n8965);
  and g12768 (n8966, n_3895, n_3896);
  and g12769 (n8967, \a[17] , n_3896);
  not g12770 (n_3897, n8966);
  not g12771 (n_3898, n8967);
  and g12772 (n8968, n_3897, n_3898);
  and g12773 (n8969, n_3721, n_3723);
  and g12774 (n8970, n_3722, n_3723);
  not g12775 (n_3899, n8969);
  not g12776 (n_3900, n8970);
  and g12777 (n8971, n_3899, n_3900);
  not g12778 (n_3901, n8968);
  not g12779 (n_3902, n8971);
  and g12780 (n8972, n_3901, n_3902);
  not g12781 (n_3903, n8972);
  and g12782 (n8973, n_3901, n_3903);
  and g12783 (n8974, n_3902, n_3903);
  not g12784 (n_3904, n8973);
  not g12785 (n_3905, n8974);
  and g12786 (n8975, n_3904, n_3905);
  and g12787 (n8976, n_299, n6233);
  and g12788 (n8977, n_301, n5663);
  and g12789 (n8978, n_300, n5939);
  and g12795 (n8981, n5139, n5666);
  not g12798 (n_3910, n8982);
  and g12799 (n8983, \a[17] , n_3910);
  not g12800 (n_3911, n8983);
  and g12801 (n8984, n_3910, n_3911);
  and g12802 (n8985, \a[17] , n_3911);
  not g12803 (n_3912, n8984);
  not g12804 (n_3913, n8985);
  and g12805 (n8986, n_3912, n_3913);
  and g12806 (n8987, n_3715, n_3717);
  and g12807 (n8988, n_3716, n_3717);
  not g12808 (n_3914, n8987);
  not g12809 (n_3915, n8988);
  and g12810 (n8989, n_3914, n_3915);
  not g12811 (n_3916, n8986);
  not g12812 (n_3917, n8989);
  and g12813 (n8990, n_3916, n_3917);
  not g12814 (n_3918, n8990);
  and g12815 (n8991, n_3916, n_3918);
  and g12816 (n8992, n_3917, n_3918);
  not g12817 (n_3919, n8991);
  not g12818 (n_3920, n8992);
  and g12819 (n8993, n_3919, n_3920);
  and g12820 (n8994, n_300, n6233);
  and g12821 (n8995, n_302, n5663);
  and g12822 (n8996, n_301, n5939);
  and g12828 (n8999, n5561, n5666);
  not g12831 (n_3925, n9000);
  and g12832 (n9001, \a[17] , n_3925);
  not g12833 (n_3926, n9001);
  and g12834 (n9002, n_3925, n_3926);
  and g12835 (n9003, \a[17] , n_3926);
  not g12836 (n_3927, n9002);
  not g12837 (n_3928, n9003);
  and g12838 (n9004, n_3927, n_3928);
  and g12839 (n9005, n_3709, n_3711);
  and g12840 (n9006, n_3710, n_3711);
  not g12841 (n_3929, n9005);
  not g12842 (n_3930, n9006);
  and g12843 (n9007, n_3929, n_3930);
  not g12844 (n_3931, n9004);
  not g12845 (n_3932, n9007);
  and g12846 (n9008, n_3931, n_3932);
  not g12847 (n_3933, n9008);
  and g12848 (n9009, n_3931, n_3933);
  and g12849 (n9010, n_3932, n_3933);
  not g12850 (n_3934, n9009);
  not g12851 (n_3935, n9010);
  and g12852 (n9011, n_3934, n_3935);
  and g12853 (n9012, n8561, n8753);
  not g12854 (n_3936, n9012);
  and g12855 (n9013, n_3705, n_3936);
  and g12856 (n9014, n_301, n6233);
  and g12857 (n9015, n_303, n5663);
  and g12858 (n9016, n_302, n5939);
  not g12859 (n_3937, n9015);
  not g12860 (n_3938, n9016);
  and g12861 (n9017, n_3937, n_3938);
  not g12862 (n_3939, n9014);
  and g12863 (n9018, n_3939, n9017);
  and g12864 (n9019, n_1409, n9018);
  and g12865 (n9020, n_1672, n9018);
  not g12866 (n_3940, n9019);
  not g12867 (n_3941, n9020);
  and g12868 (n9021, n_3940, n_3941);
  not g12869 (n_3942, n9021);
  and g12870 (n9022, \a[17] , n_3942);
  and g12871 (n9023, n_617, n9021);
  not g12872 (n_3943, n9022);
  not g12873 (n_3944, n9023);
  and g12874 (n9024, n_3943, n_3944);
  not g12875 (n_3945, n9024);
  and g12876 (n9025, n9013, n_3945);
  and g12877 (n9026, n8579, n8751);
  not g12878 (n_3946, n9026);
  and g12879 (n9027, n_3702, n_3946);
  and g12880 (n9028, n_302, n6233);
  and g12881 (n9029, n_304, n5663);
  and g12882 (n9030, n_303, n5939);
  not g12883 (n_3947, n9029);
  not g12884 (n_3948, n9030);
  and g12885 (n9031, n_3947, n_3948);
  not g12886 (n_3949, n9028);
  and g12887 (n9032, n_3949, n9031);
  and g12888 (n9033, n_1409, n9032);
  and g12889 (n9034, n_3507, n9032);
  not g12890 (n_3950, n9033);
  not g12891 (n_3951, n9034);
  and g12892 (n9035, n_3950, n_3951);
  not g12893 (n_3952, n9035);
  and g12894 (n9036, \a[17] , n_3952);
  and g12895 (n9037, n_617, n9035);
  not g12896 (n_3953, n9036);
  not g12897 (n_3954, n9037);
  and g12898 (n9038, n_3953, n_3954);
  not g12899 (n_3955, n9038);
  and g12900 (n9039, n9027, n_3955);
  and g12901 (n9040, n_303, n6233);
  and g12902 (n9041, n_305, n5663);
  and g12903 (n9042, n_304, n5939);
  and g12909 (n9045, n5666, n6007);
  not g12912 (n_3960, n9046);
  and g12913 (n9047, \a[17] , n_3960);
  not g12914 (n_3961, n9047);
  and g12915 (n9048, n_3960, n_3961);
  and g12916 (n9049, \a[17] , n_3961);
  not g12917 (n_3962, n9048);
  not g12918 (n_3963, n9049);
  and g12919 (n9050, n_3962, n_3963);
  not g12920 (n_3964, n8749);
  and g12921 (n9051, n8747, n_3964);
  not g12922 (n_3965, n9051);
  and g12923 (n9052, n_3699, n_3965);
  not g12924 (n_3966, n9050);
  and g12925 (n9053, n_3966, n9052);
  not g12926 (n_3967, n9053);
  and g12927 (n9054, n_3966, n_3967);
  and g12928 (n9055, n9052, n_3967);
  not g12929 (n_3968, n9054);
  not g12930 (n_3969, n9055);
  and g12931 (n9056, n_3968, n_3969);
  and g12932 (n9057, n_304, n6233);
  and g12933 (n9058, n_306, n5663);
  and g12934 (n9059, n_305, n5939);
  and g12940 (n9062, n5666, n5834);
  not g12943 (n_3974, n9063);
  and g12944 (n9064, \a[17] , n_3974);
  not g12945 (n_3975, n9064);
  and g12946 (n9065, n_3974, n_3975);
  and g12947 (n9066, \a[17] , n_3975);
  not g12948 (n_3976, n9065);
  not g12949 (n_3977, n9066);
  and g12950 (n9067, n_3976, n_3977);
  and g12951 (n9068, n_3692, n_3694);
  and g12952 (n9069, n_3693, n_3694);
  not g12953 (n_3978, n9068);
  not g12954 (n_3979, n9069);
  and g12955 (n9070, n_3978, n_3979);
  not g12956 (n_3980, n9067);
  not g12957 (n_3981, n9070);
  and g12958 (n9071, n_3980, n_3981);
  not g12959 (n_3982, n9071);
  and g12960 (n9072, n_3980, n_3982);
  and g12961 (n9073, n_3981, n_3982);
  not g12962 (n_3983, n9072);
  not g12963 (n_3984, n9073);
  and g12964 (n9074, n_3983, n_3984);
  and g12965 (n9075, n_305, n6233);
  and g12966 (n9076, n_307, n5663);
  and g12967 (n9077, n_306, n5939);
  and g12973 (n9080, n5666, n6143);
  not g12976 (n_3989, n9081);
  and g12977 (n9082, \a[17] , n_3989);
  not g12978 (n_3990, n9082);
  and g12979 (n9083, n_3989, n_3990);
  and g12980 (n9084, \a[17] , n_3990);
  not g12981 (n_3991, n9083);
  not g12982 (n_3992, n9084);
  and g12983 (n9085, n_3991, n_3992);
  and g12984 (n9086, n_3686, n_3688);
  and g12985 (n9087, n_3687, n_3688);
  not g12986 (n_3993, n9086);
  not g12987 (n_3994, n9087);
  and g12988 (n9088, n_3993, n_3994);
  not g12989 (n_3995, n9085);
  not g12990 (n_3996, n9088);
  and g12991 (n9089, n_3995, n_3996);
  not g12992 (n_3997, n9089);
  and g12993 (n9090, n_3995, n_3997);
  and g12994 (n9091, n_3996, n_3997);
  not g12995 (n_3998, n9090);
  not g12996 (n_3999, n9091);
  and g12997 (n9092, n_3998, n_3999);
  and g12998 (n9093, n8638, n8735);
  not g12999 (n_4000, n9093);
  and g13000 (n9094, n_3682, n_4000);
  and g13001 (n9095, n_306, n6233);
  and g13002 (n9096, n_308, n5663);
  and g13003 (n9097, n_307, n5939);
  not g13004 (n_4001, n9096);
  not g13005 (n_4002, n9097);
  and g13006 (n9098, n_4001, n_4002);
  not g13007 (n_4003, n9095);
  and g13008 (n9099, n_4003, n9098);
  and g13009 (n9100, n_1409, n9099);
  and g13010 (n9101, n_2498, n9099);
  not g13011 (n_4004, n9100);
  not g13012 (n_4005, n9101);
  and g13013 (n9102, n_4004, n_4005);
  not g13014 (n_4006, n9102);
  and g13015 (n9103, \a[17] , n_4006);
  and g13016 (n9104, n_617, n9102);
  not g13017 (n_4007, n9103);
  not g13018 (n_4008, n9104);
  and g13019 (n9105, n_4007, n_4008);
  not g13020 (n_4009, n9105);
  and g13021 (n9106, n9094, n_4009);
  not g13022 (n_4010, n8733);
  and g13023 (n9107, n8731, n_4010);
  not g13024 (n_4011, n9107);
  and g13025 (n9108, n_3679, n_4011);
  and g13026 (n9109, n_307, n6233);
  and g13027 (n9110, n_309, n5663);
  and g13028 (n9111, n_308, n5939);
  not g13029 (n_4012, n9110);
  not g13030 (n_4013, n9111);
  and g13031 (n9112, n_4012, n_4013);
  not g13032 (n_4014, n9109);
  and g13033 (n9113, n_4014, n9112);
  and g13034 (n9114, n_1409, n9113);
  and g13035 (n9115, n_2511, n9113);
  not g13036 (n_4015, n9114);
  not g13037 (n_4016, n9115);
  and g13038 (n9116, n_4015, n_4016);
  not g13039 (n_4017, n9116);
  and g13040 (n9117, \a[17] , n_4017);
  and g13041 (n9118, n_617, n9116);
  not g13042 (n_4018, n9117);
  not g13043 (n_4019, n9118);
  and g13044 (n9119, n_4018, n_4019);
  not g13045 (n_4020, n9119);
  and g13046 (n9120, n9108, n_4020);
  and g13047 (n9121, n8670, n8729);
  not g13048 (n_4021, n9121);
  and g13049 (n9122, n_3675, n_4021);
  and g13050 (n9123, n_308, n6233);
  and g13051 (n9124, n_310, n5663);
  and g13052 (n9125, n_309, n5939);
  not g13053 (n_4022, n9124);
  not g13054 (n_4023, n9125);
  and g13055 (n9126, n_4022, n_4023);
  not g13056 (n_4024, n9123);
  and g13057 (n9127, n_4024, n9126);
  and g13058 (n9128, n_1409, n9127);
  and g13059 (n9129, n_2839, n9127);
  not g13060 (n_4025, n9128);
  not g13061 (n_4026, n9129);
  and g13062 (n9130, n_4025, n_4026);
  not g13063 (n_4027, n9130);
  and g13064 (n9131, \a[17] , n_4027);
  and g13065 (n9132, n_617, n9130);
  not g13066 (n_4028, n9131);
  not g13067 (n_4029, n9132);
  and g13068 (n9133, n_4028, n_4029);
  not g13069 (n_4030, n9133);
  and g13070 (n9134, n9122, n_4030);
  and g13071 (n9135, n_309, n6233);
  and g13072 (n9136, n_311, n5663);
  and g13073 (n9137, n_310, n5939);
  and g13079 (n9140, n5666, n6541);
  not g13082 (n_4035, n9141);
  and g13083 (n9142, \a[17] , n_4035);
  not g13084 (n_4036, n9142);
  and g13085 (n9143, n_4035, n_4036);
  and g13086 (n9144, \a[17] , n_4036);
  not g13087 (n_4037, n9143);
  not g13088 (n_4038, n9144);
  and g13089 (n9145, n_4037, n_4038);
  not g13090 (n_4039, n8727);
  and g13091 (n9146, n8725, n_4039);
  not g13092 (n_4040, n9146);
  and g13093 (n9147, n_3672, n_4040);
  not g13094 (n_4041, n9145);
  and g13095 (n9148, n_4041, n9147);
  not g13096 (n_4042, n9148);
  and g13097 (n9149, n_4041, n_4042);
  and g13098 (n9150, n9147, n_4042);
  not g13099 (n_4043, n9149);
  not g13100 (n_4044, n9150);
  and g13101 (n9151, n_4043, n_4044);
  and g13102 (n9152, n_3665, n_3667);
  and g13103 (n9153, n_3666, n_3667);
  not g13104 (n_4045, n9152);
  not g13105 (n_4046, n9153);
  and g13106 (n9154, n_4045, n_4046);
  and g13107 (n9155, n_310, n6233);
  and g13108 (n9156, n_312, n5663);
  and g13109 (n9157, n_311, n5939);
  not g13110 (n_4047, n9156);
  not g13111 (n_4048, n9157);
  and g13112 (n9158, n_4047, n_4048);
  not g13113 (n_4049, n9155);
  and g13114 (n9159, n_4049, n9158);
  and g13115 (n9160, n_1409, n9159);
  and g13116 (n9161, n_3239, n9159);
  not g13117 (n_4050, n9160);
  not g13118 (n_4051, n9161);
  and g13119 (n9162, n_4050, n_4051);
  not g13120 (n_4052, n9162);
  and g13121 (n9163, \a[17] , n_4052);
  and g13122 (n9164, n_617, n9162);
  not g13123 (n_4053, n9163);
  not g13124 (n_4054, n9164);
  and g13125 (n9165, n_4053, n_4054);
  not g13126 (n_4055, n9154);
  not g13127 (n_4056, n9165);
  and g13128 (n9166, n_4055, n_4056);
  and g13129 (n9167, n_311, n6233);
  and g13130 (n9168, n_313, n5663);
  and g13131 (n9169, n_312, n5939);
  and g13137 (n9172, n5666, n6646);
  not g13140 (n_4061, n9173);
  and g13141 (n9174, \a[17] , n_4061);
  not g13142 (n_4062, n9174);
  and g13143 (n9175, n_4061, n_4062);
  and g13144 (n9176, \a[17] , n_4062);
  not g13145 (n_4063, n9175);
  not g13146 (n_4064, n9176);
  and g13147 (n9177, n_4063, n_4064);
  not g13148 (n_4065, n8696);
  and g13149 (n9178, n_4065, n8707);
  not g13150 (n_4066, n8708);
  not g13151 (n_4067, n9178);
  and g13152 (n9179, n_4066, n_4067);
  not g13153 (n_4068, n9177);
  and g13154 (n9180, n_4068, n9179);
  not g13155 (n_4069, n9180);
  and g13156 (n9181, n_4068, n_4069);
  and g13157 (n9182, n9179, n_4069);
  not g13158 (n_4070, n9181);
  not g13159 (n_4071, n9182);
  and g13160 (n9183, n_4070, n_4071);
  not g13161 (n_4072, n8695);
  and g13162 (n9184, n8693, n_4072);
  not g13163 (n_4073, n9184);
  and g13164 (n9185, n_4065, n_4073);
  and g13165 (n9186, n_312, n6233);
  and g13166 (n9187, n_314, n5663);
  and g13167 (n9188, n_313, n5939);
  not g13168 (n_4074, n9187);
  not g13169 (n_4075, n9188);
  and g13170 (n9189, n_4074, n_4075);
  not g13171 (n_4076, n9186);
  and g13172 (n9190, n_4076, n9189);
  and g13173 (n9191, n_1409, n9190);
  and g13174 (n9192, n_2891, n9190);
  not g13175 (n_4077, n9191);
  not g13176 (n_4078, n9192);
  and g13177 (n9193, n_4077, n_4078);
  not g13178 (n_4079, n9193);
  and g13179 (n9194, \a[17] , n_4079);
  and g13180 (n9195, n_617, n9193);
  not g13181 (n_4080, n9194);
  not g13182 (n_4081, n9195);
  and g13183 (n9196, n_4080, n_4081);
  not g13184 (n_4082, n9196);
  and g13185 (n9197, n9185, n_4082);
  and g13186 (n9198, n_316, n5939);
  and g13187 (n9199, n_315, n6233);
  not g13188 (n_4083, n9198);
  not g13189 (n_4084, n9199);
  and g13190 (n9200, n_4083, n_4084);
  and g13191 (n9201, n5666, n_2588);
  not g13192 (n_4085, n9201);
  and g13193 (n9202, n9200, n_4085);
  not g13194 (n_4086, n9202);
  and g13195 (n9203, \a[17] , n_4086);
  not g13196 (n_4087, n9203);
  and g13197 (n9204, \a[17] , n_4087);
  and g13198 (n9205, n_4086, n_4087);
  not g13199 (n_4088, n9204);
  not g13200 (n_4089, n9205);
  and g13201 (n9206, n_4088, n_4089);
  and g13202 (n9207, n_316, n_1408);
  not g13203 (n_4090, n9207);
  and g13204 (n9208, \a[17] , n_4090);
  not g13205 (n_4091, n9206);
  and g13206 (n9209, n_4091, n9208);
  and g13207 (n9210, n_314, n6233);
  and g13208 (n9211, n_316, n5663);
  and g13209 (n9212, n_315, n5939);
  not g13210 (n_4092, n9211);
  not g13211 (n_4093, n9212);
  and g13212 (n9213, n_4092, n_4093);
  not g13213 (n_4094, n9210);
  and g13214 (n9214, n_4094, n9213);
  and g13215 (n9215, n_1409, n9214);
  and g13216 (n9216, n_2612, n9214);
  not g13217 (n_4095, n9215);
  not g13218 (n_4096, n9216);
  and g13219 (n9217, n_4095, n_4096);
  not g13220 (n_4097, n9217);
  and g13221 (n9218, \a[17] , n_4097);
  and g13222 (n9219, n_617, n9217);
  not g13223 (n_4098, n9218);
  not g13224 (n_4099, n9219);
  and g13225 (n9220, n_4098, n_4099);
  not g13226 (n_4100, n9220);
  and g13227 (n9221, n9209, n_4100);
  and g13228 (n9222, n8694, n9221);
  not g13229 (n_4101, n9222);
  and g13230 (n9223, n9221, n_4101);
  and g13231 (n9224, n8694, n_4101);
  not g13232 (n_4102, n9223);
  not g13233 (n_4103, n9224);
  and g13234 (n9225, n_4102, n_4103);
  and g13235 (n9226, n_313, n6233);
  and g13236 (n9227, n_315, n5663);
  and g13237 (n9228, n_314, n5939);
  and g13243 (n9231, n5666, n6806);
  not g13246 (n_4108, n9232);
  and g13247 (n9233, \a[17] , n_4108);
  not g13248 (n_4109, n9233);
  and g13249 (n9234, \a[17] , n_4109);
  and g13250 (n9235, n_4108, n_4109);
  not g13251 (n_4110, n9234);
  not g13252 (n_4111, n9235);
  and g13253 (n9236, n_4110, n_4111);
  not g13254 (n_4112, n9225);
  not g13255 (n_4113, n9236);
  and g13256 (n9237, n_4112, n_4113);
  not g13257 (n_4114, n9237);
  and g13258 (n9238, n_4101, n_4114);
  not g13259 (n_4115, n9185);
  and g13260 (n9239, n_4115, n9196);
  not g13261 (n_4116, n9197);
  not g13262 (n_4117, n9239);
  and g13263 (n9240, n_4116, n_4117);
  not g13264 (n_4118, n9238);
  and g13265 (n9241, n_4118, n9240);
  not g13266 (n_4119, n9241);
  and g13267 (n9242, n_4116, n_4119);
  not g13268 (n_4120, n9183);
  not g13269 (n_4121, n9242);
  and g13270 (n9243, n_4120, n_4121);
  not g13271 (n_4122, n9243);
  and g13272 (n9244, n_4069, n_4122);
  and g13273 (n9245, n9154, n9165);
  not g13274 (n_4123, n9166);
  not g13275 (n_4124, n9245);
  and g13276 (n9246, n_4123, n_4124);
  not g13277 (n_4125, n9244);
  and g13278 (n9247, n_4125, n9246);
  not g13279 (n_4126, n9247);
  and g13280 (n9248, n_4123, n_4126);
  not g13281 (n_4127, n9151);
  not g13282 (n_4128, n9248);
  and g13283 (n9249, n_4127, n_4128);
  not g13284 (n_4129, n9249);
  and g13285 (n9250, n_4042, n_4129);
  not g13286 (n_4130, n9134);
  and g13287 (n9251, n9122, n_4130);
  and g13288 (n9252, n_4030, n_4130);
  not g13289 (n_4131, n9251);
  not g13290 (n_4132, n9252);
  and g13291 (n9253, n_4131, n_4132);
  not g13292 (n_4133, n9250);
  not g13293 (n_4134, n9253);
  and g13294 (n9254, n_4133, n_4134);
  not g13295 (n_4135, n9254);
  and g13296 (n9255, n_4130, n_4135);
  not g13297 (n_4136, n9120);
  and g13298 (n9256, n9108, n_4136);
  and g13299 (n9257, n_4020, n_4136);
  not g13300 (n_4137, n9256);
  not g13301 (n_4138, n9257);
  and g13302 (n9258, n_4137, n_4138);
  not g13303 (n_4139, n9255);
  not g13304 (n_4140, n9258);
  and g13305 (n9259, n_4139, n_4140);
  not g13306 (n_4141, n9259);
  and g13307 (n9260, n_4136, n_4141);
  not g13308 (n_4142, n9094);
  and g13309 (n9261, n_4142, n9105);
  not g13310 (n_4143, n9106);
  not g13311 (n_4144, n9261);
  and g13312 (n9262, n_4143, n_4144);
  not g13313 (n_4145, n9260);
  and g13314 (n9263, n_4145, n9262);
  not g13315 (n_4146, n9263);
  and g13316 (n9264, n_4143, n_4146);
  not g13317 (n_4147, n9092);
  not g13318 (n_4148, n9264);
  and g13319 (n9265, n_4147, n_4148);
  not g13320 (n_4149, n9265);
  and g13321 (n9266, n_3997, n_4149);
  not g13322 (n_4150, n9074);
  not g13323 (n_4151, n9266);
  and g13324 (n9267, n_4150, n_4151);
  not g13325 (n_4152, n9267);
  and g13326 (n9268, n_3982, n_4152);
  not g13327 (n_4153, n9056);
  not g13328 (n_4154, n9268);
  and g13329 (n9269, n_4153, n_4154);
  not g13330 (n_4155, n9269);
  and g13331 (n9270, n_3967, n_4155);
  not g13332 (n_4156, n9039);
  and g13333 (n9271, n9027, n_4156);
  and g13334 (n9272, n_3955, n_4156);
  not g13335 (n_4157, n9271);
  not g13336 (n_4158, n9272);
  and g13337 (n9273, n_4157, n_4158);
  not g13338 (n_4159, n9270);
  not g13339 (n_4160, n9273);
  and g13340 (n9274, n_4159, n_4160);
  not g13341 (n_4161, n9274);
  and g13342 (n9275, n_4156, n_4161);
  not g13343 (n_4162, n9013);
  and g13344 (n9276, n_4162, n9024);
  not g13345 (n_4163, n9025);
  not g13346 (n_4164, n9276);
  and g13347 (n9277, n_4163, n_4164);
  not g13348 (n_4165, n9275);
  and g13349 (n9278, n_4165, n9277);
  not g13350 (n_4166, n9278);
  and g13351 (n9279, n_4163, n_4166);
  not g13352 (n_4167, n9011);
  not g13353 (n_4168, n9279);
  and g13354 (n9280, n_4167, n_4168);
  not g13355 (n_4169, n9280);
  and g13356 (n9281, n_3933, n_4169);
  not g13357 (n_4170, n8993);
  not g13358 (n_4171, n9281);
  and g13359 (n9282, n_4170, n_4171);
  not g13360 (n_4172, n9282);
  and g13361 (n9283, n_3918, n_4172);
  not g13362 (n_4173, n8975);
  not g13363 (n_4174, n9283);
  and g13364 (n9284, n_4173, n_4174);
  not g13365 (n_4175, n9284);
  and g13366 (n9285, n_3903, n_4175);
  not g13367 (n_4176, n8957);
  not g13368 (n_4177, n9285);
  and g13369 (n9286, n_4176, n_4177);
  not g13370 (n_4178, n9286);
  and g13371 (n9287, n_3888, n_4178);
  not g13372 (n_4179, n8939);
  not g13373 (n_4180, n9287);
  and g13374 (n9288, n_4179, n_4180);
  not g13375 (n_4181, n9288);
  and g13376 (n9289, n_3873, n_4181);
  not g13377 (n_4182, n8921);
  not g13378 (n_4183, n9289);
  and g13379 (n9290, n_4182, n_4183);
  not g13380 (n_4184, n9290);
  and g13381 (n9291, n_3858, n_4184);
  not g13382 (n_4185, n8903);
  not g13383 (n_4186, n9291);
  and g13384 (n9292, n_4185, n_4186);
  not g13385 (n_4187, n9292);
  and g13386 (n9293, n_3843, n_4187);
  not g13387 (n_4188, n8806);
  and g13388 (n9294, n8804, n_4188);
  not g13389 (n_4189, n9294);
  and g13390 (n9295, n_3763, n_4189);
  not g13391 (n_4190, n9293);
  and g13392 (n9296, n_4190, n9295);
  and g13393 (n9297, n_236, n7101);
  and g13394 (n9298, n_260, n6402);
  and g13395 (n9299, n_237, n6951);
  and g13401 (n9302, n3347, n6397);
  not g13404 (n_4195, n9303);
  and g13405 (n9304, \a[14] , n_4195);
  not g13406 (n_4196, n9304);
  and g13407 (n9305, n_4195, n_4196);
  and g13408 (n9306, \a[14] , n_4196);
  not g13409 (n_4197, n9305);
  not g13410 (n_4198, n9306);
  and g13411 (n9307, n_4197, n_4198);
  not g13412 (n_4199, n9295);
  and g13413 (n9308, n9293, n_4199);
  not g13414 (n_4200, n9296);
  not g13415 (n_4201, n9308);
  and g13416 (n9309, n_4200, n_4201);
  not g13417 (n_4202, n9307);
  and g13418 (n9310, n_4202, n9309);
  not g13419 (n_4203, n9310);
  and g13420 (n9311, n_4200, n_4203);
  not g13421 (n_4204, n8885);
  not g13422 (n_4205, n9311);
  and g13423 (n9312, n_4204, n_4205);
  and g13424 (n9313, n8885, n9311);
  not g13425 (n_4206, n9312);
  not g13426 (n_4207, n9313);
  and g13427 (n9314, n_4206, n_4207);
  and g13428 (n9315, n_480, n7983);
  and g13429 (n9316, n_484, n7291);
  and g13430 (n9317, n_485, n7632);
  and g13436 (n9320, n3627, n7294);
  not g13439 (n_4212, n9321);
  and g13440 (n9322, \a[11] , n_4212);
  not g13441 (n_4213, n9322);
  and g13442 (n9323, \a[11] , n_4213);
  and g13443 (n9324, n_4212, n_4213);
  not g13444 (n_4214, n9323);
  not g13445 (n_4215, n9324);
  and g13446 (n9325, n_4214, n_4215);
  not g13447 (n_4216, n9325);
  and g13448 (n9326, n9314, n_4216);
  not g13449 (n_4217, n9326);
  and g13450 (n9327, n_4206, n_4217);
  not g13451 (n_4218, n8882);
  not g13452 (n_4219, n9327);
  and g13453 (n9328, n_4218, n_4219);
  and g13454 (n9329, n8882, n9327);
  not g13455 (n_4220, n9328);
  not g13456 (n_4221, n9329);
  and g13457 (n9330, n_4220, n_4221);
  and g13458 (n9331, n8413, n_3427);
  and g13459 (n9332, n_560, n9331);
  and g13460 (n9333, n_565, n8418);
  and g13461 (n9334, n_566, n8860);
  and g13467 (n9337, n4067, n8421);
  not g13470 (n_4226, n9338);
  and g13471 (n9339, \a[8] , n_4226);
  not g13472 (n_4227, n9339);
  and g13473 (n9340, \a[8] , n_4227);
  and g13474 (n9341, n_4226, n_4227);
  not g13475 (n_4228, n9340);
  not g13476 (n_4229, n9341);
  and g13477 (n9342, n_4228, n_4229);
  not g13478 (n_4230, n9342);
  and g13479 (n9343, n9330, n_4230);
  not g13480 (n_4231, n9343);
  and g13481 (n9344, n_4220, n_4231);
  and g13482 (n9345, n_712, n9331);
  and g13483 (n9346, n_566, n8418);
  and g13484 (n9347, n_560, n8860);
  not g13485 (n_4232, n9346);
  not g13486 (n_4233, n9347);
  and g13487 (n9348, n_4232, n_4233);
  not g13488 (n_4234, n9345);
  and g13489 (n9349, n_4234, n9348);
  and g13490 (n9350, n_3428, n9349);
  and g13491 (n9351, n_888, n9349);
  not g13492 (n_4235, n9350);
  not g13493 (n_4236, n9351);
  and g13494 (n9352, n_4235, n_4236);
  not g13495 (n_4237, n9352);
  and g13496 (n9353, \a[8] , n_4237);
  and g13497 (n9354, n_1106, n9352);
  not g13498 (n_4238, n9353);
  not g13499 (n_4239, n9354);
  and g13500 (n9355, n_4238, n_4239);
  not g13501 (n_4240, n9344);
  not g13502 (n_4241, n9355);
  and g13503 (n9356, n_4240, n_4241);
  not g13504 (n_4242, n9356);
  and g13505 (n9357, n_4240, n_4242);
  and g13506 (n9358, n_4241, n_4242);
  not g13507 (n_4243, n9357);
  not g13508 (n_4244, n9358);
  and g13509 (n9359, n_4243, n_4244);
  not g13510 (n_4245, n8854);
  not g13511 (n_4246, n8856);
  and g13512 (n9360, n_4245, n_4246);
  not g13513 (n_4247, n9360);
  and g13514 (n9361, n_3806, n_4247);
  not g13515 (n_4248, n9359);
  and g13516 (n9362, n_4248, n9361);
  not g13517 (n_4249, n9362);
  and g13518 (n9363, n_4242, n_4249);
  not g13519 (n_4250, n8874);
  and g13520 (n9364, n8872, n_4250);
  not g13521 (n_4251, n9364);
  and g13522 (n9365, n_3822, n_4251);
  not g13523 (n_4252, n9363);
  and g13524 (n9366, n_4252, n9365);
  and g13525 (n9367, n9314, n_4217);
  and g13526 (n9368, n_4216, n_4217);
  not g13527 (n_4253, n9367);
  not g13528 (n_4254, n9368);
  and g13529 (n9369, n_4253, n_4254);
  and g13530 (n9370, n8903, n9291);
  not g13531 (n_4255, n9370);
  and g13532 (n9371, n_4187, n_4255);
  and g13533 (n9372, n_237, n7101);
  and g13534 (n9373, n_275, n6402);
  and g13535 (n9374, n_260, n6951);
  not g13536 (n_4256, n9373);
  not g13537 (n_4257, n9374);
  and g13538 (n9375, n_4256, n_4257);
  not g13539 (n_4258, n9372);
  and g13540 (n9376, n_4258, n9375);
  and g13541 (n9377, n_1885, n9376);
  not g13542 (n_4259, n3331);
  and g13543 (n9378, n_4259, n9376);
  not g13544 (n_4260, n9377);
  not g13545 (n_4261, n9378);
  and g13546 (n9379, n_4260, n_4261);
  not g13547 (n_4262, n9379);
  and g13548 (n9380, \a[14] , n_4262);
  and g13549 (n9381, n_652, n9379);
  not g13550 (n_4263, n9380);
  not g13551 (n_4264, n9381);
  and g13552 (n9382, n_4263, n_4264);
  not g13553 (n_4265, n9382);
  and g13554 (n9383, n9371, n_4265);
  and g13555 (n9384, n8921, n9289);
  not g13556 (n_4266, n9384);
  and g13557 (n9385, n_4184, n_4266);
  and g13558 (n9386, n_260, n7101);
  and g13559 (n9387, n_281, n6402);
  and g13560 (n9388, n_275, n6951);
  not g13561 (n_4267, n9387);
  not g13562 (n_4268, n9388);
  and g13563 (n9389, n_4267, n_4268);
  not g13564 (n_4269, n9386);
  and g13565 (n9390, n_4269, n9389);
  and g13566 (n9391, n_1885, n9390);
  and g13567 (n9392, n_958, n9390);
  not g13568 (n_4270, n9391);
  not g13569 (n_4271, n9392);
  and g13570 (n9393, n_4270, n_4271);
  not g13571 (n_4272, n9393);
  and g13572 (n9394, \a[14] , n_4272);
  and g13573 (n9395, n_652, n9393);
  not g13574 (n_4273, n9394);
  not g13575 (n_4274, n9395);
  and g13576 (n9396, n_4273, n_4274);
  not g13577 (n_4275, n9396);
  and g13578 (n9397, n9385, n_4275);
  and g13579 (n9398, n8939, n9287);
  not g13580 (n_4276, n9398);
  and g13581 (n9399, n_4181, n_4276);
  and g13582 (n9400, n_275, n7101);
  and g13583 (n9401, n_286, n6402);
  and g13584 (n9402, n_281, n6951);
  not g13585 (n_4277, n9401);
  not g13586 (n_4278, n9402);
  and g13587 (n9403, n_4277, n_4278);
  not g13588 (n_4279, n9400);
  and g13589 (n9404, n_4279, n9403);
  and g13590 (n9405, n_1885, n9404);
  and g13591 (n9406, n_1450, n9404);
  not g13592 (n_4280, n9405);
  not g13593 (n_4281, n9406);
  and g13594 (n9407, n_4280, n_4281);
  not g13595 (n_4282, n9407);
  and g13596 (n9408, \a[14] , n_4282);
  and g13597 (n9409, n_652, n9407);
  not g13598 (n_4283, n9408);
  not g13599 (n_4284, n9409);
  and g13600 (n9410, n_4283, n_4284);
  not g13601 (n_4285, n9410);
  and g13602 (n9411, n9399, n_4285);
  and g13603 (n9412, n8957, n9285);
  not g13604 (n_4286, n9412);
  and g13605 (n9413, n_4178, n_4286);
  and g13606 (n9414, n_281, n7101);
  and g13607 (n9415, n_293, n6402);
  and g13608 (n9416, n_286, n6951);
  not g13609 (n_4287, n9415);
  not g13610 (n_4288, n9416);
  and g13611 (n9417, n_4287, n_4288);
  not g13612 (n_4289, n9414);
  and g13613 (n9418, n_4289, n9417);
  and g13614 (n9419, n_1885, n9418);
  and g13615 (n9420, n_1228, n9418);
  not g13616 (n_4290, n9419);
  not g13617 (n_4291, n9420);
  and g13618 (n9421, n_4290, n_4291);
  not g13619 (n_4292, n9421);
  and g13620 (n9422, \a[14] , n_4292);
  and g13621 (n9423, n_652, n9421);
  not g13622 (n_4293, n9422);
  not g13623 (n_4294, n9423);
  and g13624 (n9424, n_4293, n_4294);
  not g13625 (n_4295, n9424);
  and g13626 (n9425, n9413, n_4295);
  and g13627 (n9426, n8975, n9283);
  not g13628 (n_4296, n9426);
  and g13629 (n9427, n_4175, n_4296);
  and g13630 (n9428, n_286, n7101);
  and g13631 (n9429, n_295, n6402);
  and g13632 (n9430, n_293, n6951);
  not g13633 (n_4297, n9429);
  not g13634 (n_4298, n9430);
  and g13635 (n9431, n_4297, n_4298);
  not g13636 (n_4299, n9428);
  and g13637 (n9432, n_4299, n9431);
  and g13638 (n9433, n_1885, n9432);
  and g13639 (n9434, n_1134, n9432);
  not g13640 (n_4300, n9433);
  not g13641 (n_4301, n9434);
  and g13642 (n9435, n_4300, n_4301);
  not g13643 (n_4302, n9435);
  and g13644 (n9436, \a[14] , n_4302);
  and g13645 (n9437, n_652, n9435);
  not g13646 (n_4303, n9436);
  not g13647 (n_4304, n9437);
  and g13648 (n9438, n_4303, n_4304);
  not g13649 (n_4305, n9438);
  and g13650 (n9439, n9427, n_4305);
  and g13651 (n9440, n8993, n9281);
  not g13652 (n_4306, n9440);
  and g13653 (n9441, n_4172, n_4306);
  and g13654 (n9442, n_293, n7101);
  and g13655 (n9443, n_298, n6402);
  and g13656 (n9444, n_295, n6951);
  not g13657 (n_4307, n9443);
  not g13658 (n_4308, n9444);
  and g13659 (n9445, n_4307, n_4308);
  not g13660 (n_4309, n9442);
  and g13661 (n9446, n_4309, n9445);
  and g13662 (n9447, n_1885, n9446);
  and g13663 (n9448, n_1789, n9446);
  not g13664 (n_4310, n9447);
  not g13665 (n_4311, n9448);
  and g13666 (n9449, n_4310, n_4311);
  not g13667 (n_4312, n9449);
  and g13668 (n9450, \a[14] , n_4312);
  and g13669 (n9451, n_652, n9449);
  not g13670 (n_4313, n9450);
  not g13671 (n_4314, n9451);
  and g13672 (n9452, n_4313, n_4314);
  not g13673 (n_4315, n9452);
  and g13674 (n9453, n9441, n_4315);
  and g13675 (n9454, n9011, n9279);
  not g13676 (n_4316, n9454);
  and g13677 (n9455, n_4169, n_4316);
  and g13678 (n9456, n_295, n7101);
  and g13679 (n9457, n_299, n6402);
  and g13680 (n9458, n_298, n6951);
  not g13681 (n_4317, n9457);
  not g13682 (n_4318, n9458);
  and g13683 (n9459, n_4317, n_4318);
  not g13684 (n_4319, n9456);
  and g13685 (n9460, n_4319, n9459);
  and g13686 (n9461, n_1885, n9460);
  and g13687 (n9462, n_3456, n9460);
  not g13688 (n_4320, n9461);
  not g13689 (n_4321, n9462);
  and g13690 (n9463, n_4320, n_4321);
  not g13691 (n_4322, n9463);
  and g13692 (n9464, \a[14] , n_4322);
  and g13693 (n9465, n_652, n9463);
  not g13694 (n_4323, n9464);
  not g13695 (n_4324, n9465);
  and g13696 (n9466, n_4323, n_4324);
  not g13697 (n_4325, n9466);
  and g13698 (n9467, n9455, n_4325);
  and g13699 (n9468, n_298, n7101);
  and g13700 (n9469, n_300, n6402);
  and g13701 (n9470, n_299, n6951);
  and g13707 (n9473, n5114, n6397);
  not g13710 (n_4330, n9474);
  and g13711 (n9475, \a[14] , n_4330);
  not g13712 (n_4331, n9475);
  and g13713 (n9476, n_4330, n_4331);
  and g13714 (n9477, \a[14] , n_4331);
  not g13715 (n_4332, n9476);
  not g13716 (n_4333, n9477);
  and g13717 (n9478, n_4332, n_4333);
  not g13718 (n_4334, n9277);
  and g13719 (n9479, n9275, n_4334);
  not g13720 (n_4335, n9479);
  and g13721 (n9480, n_4166, n_4335);
  not g13722 (n_4336, n9478);
  and g13723 (n9481, n_4336, n9480);
  not g13724 (n_4337, n9481);
  and g13725 (n9482, n_4336, n_4337);
  and g13726 (n9483, n9480, n_4337);
  not g13727 (n_4338, n9482);
  not g13728 (n_4339, n9483);
  and g13729 (n9484, n_4338, n_4339);
  and g13730 (n9485, n_299, n7101);
  and g13731 (n9486, n_301, n6402);
  and g13732 (n9487, n_300, n6951);
  and g13738 (n9490, n5139, n6397);
  not g13741 (n_4344, n9491);
  and g13742 (n9492, \a[14] , n_4344);
  not g13743 (n_4345, n9492);
  and g13744 (n9493, n_4344, n_4345);
  and g13745 (n9494, \a[14] , n_4345);
  not g13746 (n_4346, n9493);
  not g13747 (n_4347, n9494);
  and g13748 (n9495, n_4346, n_4347);
  and g13749 (n9496, n_4159, n_4161);
  and g13750 (n9497, n_4160, n_4161);
  not g13751 (n_4348, n9496);
  not g13752 (n_4349, n9497);
  and g13753 (n9498, n_4348, n_4349);
  not g13754 (n_4350, n9495);
  not g13755 (n_4351, n9498);
  and g13756 (n9499, n_4350, n_4351);
  not g13757 (n_4352, n9499);
  and g13758 (n9500, n_4350, n_4352);
  and g13759 (n9501, n_4351, n_4352);
  not g13760 (n_4353, n9500);
  not g13761 (n_4354, n9501);
  and g13762 (n9502, n_4353, n_4354);
  and g13763 (n9503, n9056, n9268);
  not g13764 (n_4355, n9503);
  and g13765 (n9504, n_4155, n_4355);
  and g13766 (n9505, n_300, n7101);
  and g13767 (n9506, n_302, n6402);
  and g13768 (n9507, n_301, n6951);
  not g13769 (n_4356, n9506);
  not g13770 (n_4357, n9507);
  and g13771 (n9508, n_4356, n_4357);
  not g13772 (n_4358, n9505);
  and g13773 (n9509, n_4358, n9508);
  and g13774 (n9510, n_1885, n9509);
  and g13775 (n9511, n_1801, n9509);
  not g13776 (n_4359, n9510);
  not g13777 (n_4360, n9511);
  and g13778 (n9512, n_4359, n_4360);
  not g13779 (n_4361, n9512);
  and g13780 (n9513, \a[14] , n_4361);
  and g13781 (n9514, n_652, n9512);
  not g13782 (n_4362, n9513);
  not g13783 (n_4363, n9514);
  and g13784 (n9515, n_4362, n_4363);
  not g13785 (n_4364, n9515);
  and g13786 (n9516, n9504, n_4364);
  and g13787 (n9517, n9074, n9266);
  not g13788 (n_4365, n9517);
  and g13789 (n9518, n_4152, n_4365);
  and g13790 (n9519, n_301, n7101);
  and g13791 (n9520, n_303, n6402);
  and g13792 (n9521, n_302, n6951);
  not g13793 (n_4366, n9520);
  not g13794 (n_4367, n9521);
  and g13795 (n9522, n_4366, n_4367);
  not g13796 (n_4368, n9519);
  and g13797 (n9523, n_4368, n9522);
  and g13798 (n9524, n_1885, n9523);
  and g13799 (n9525, n_1672, n9523);
  not g13800 (n_4369, n9524);
  not g13801 (n_4370, n9525);
  and g13802 (n9526, n_4369, n_4370);
  not g13803 (n_4371, n9526);
  and g13804 (n9527, \a[14] , n_4371);
  and g13805 (n9528, n_652, n9526);
  not g13806 (n_4372, n9527);
  not g13807 (n_4373, n9528);
  and g13808 (n9529, n_4372, n_4373);
  not g13809 (n_4374, n9529);
  and g13810 (n9530, n9518, n_4374);
  and g13811 (n9531, n9092, n9264);
  not g13812 (n_4375, n9531);
  and g13813 (n9532, n_4149, n_4375);
  and g13814 (n9533, n_302, n7101);
  and g13815 (n9534, n_304, n6402);
  and g13816 (n9535, n_303, n6951);
  not g13817 (n_4376, n9534);
  not g13818 (n_4377, n9535);
  and g13819 (n9536, n_4376, n_4377);
  not g13820 (n_4378, n9533);
  and g13821 (n9537, n_4378, n9536);
  and g13822 (n9538, n_1885, n9537);
  and g13823 (n9539, n_3507, n9537);
  not g13824 (n_4379, n9538);
  not g13825 (n_4380, n9539);
  and g13826 (n9540, n_4379, n_4380);
  not g13827 (n_4381, n9540);
  and g13828 (n9541, \a[14] , n_4381);
  and g13829 (n9542, n_652, n9540);
  not g13830 (n_4382, n9541);
  not g13831 (n_4383, n9542);
  and g13832 (n9543, n_4382, n_4383);
  not g13833 (n_4384, n9543);
  and g13834 (n9544, n9532, n_4384);
  and g13835 (n9545, n_303, n7101);
  and g13836 (n9546, n_305, n6402);
  and g13837 (n9547, n_304, n6951);
  and g13843 (n9550, n6007, n6397);
  not g13846 (n_4389, n9551);
  and g13847 (n9552, \a[14] , n_4389);
  not g13848 (n_4390, n9552);
  and g13849 (n9553, n_4389, n_4390);
  and g13850 (n9554, \a[14] , n_4390);
  not g13851 (n_4391, n9553);
  not g13852 (n_4392, n9554);
  and g13853 (n9555, n_4391, n_4392);
  not g13854 (n_4393, n9262);
  and g13855 (n9556, n9260, n_4393);
  not g13856 (n_4394, n9556);
  and g13857 (n9557, n_4146, n_4394);
  not g13858 (n_4395, n9555);
  and g13859 (n9558, n_4395, n9557);
  not g13860 (n_4396, n9558);
  and g13861 (n9559, n_4395, n_4396);
  and g13862 (n9560, n9557, n_4396);
  not g13863 (n_4397, n9559);
  not g13864 (n_4398, n9560);
  and g13865 (n9561, n_4397, n_4398);
  and g13866 (n9562, n_304, n7101);
  and g13867 (n9563, n_306, n6402);
  and g13868 (n9564, n_305, n6951);
  and g13874 (n9567, n5834, n6397);
  not g13877 (n_4403, n9568);
  and g13878 (n9569, \a[14] , n_4403);
  not g13879 (n_4404, n9569);
  and g13880 (n9570, n_4403, n_4404);
  and g13881 (n9571, \a[14] , n_4404);
  not g13882 (n_4405, n9570);
  not g13883 (n_4406, n9571);
  and g13884 (n9572, n_4405, n_4406);
  and g13885 (n9573, n_4139, n_4141);
  and g13886 (n9574, n_4140, n_4141);
  not g13887 (n_4407, n9573);
  not g13888 (n_4408, n9574);
  and g13889 (n9575, n_4407, n_4408);
  not g13890 (n_4409, n9572);
  not g13891 (n_4410, n9575);
  and g13892 (n9576, n_4409, n_4410);
  not g13893 (n_4411, n9576);
  and g13894 (n9577, n_4409, n_4411);
  and g13895 (n9578, n_4410, n_4411);
  not g13896 (n_4412, n9577);
  not g13897 (n_4413, n9578);
  and g13898 (n9579, n_4412, n_4413);
  and g13899 (n9580, n_305, n7101);
  and g13900 (n9581, n_307, n6402);
  and g13901 (n9582, n_306, n6951);
  and g13907 (n9585, n6143, n6397);
  not g13910 (n_4418, n9586);
  and g13911 (n9587, \a[14] , n_4418);
  not g13912 (n_4419, n9587);
  and g13913 (n9588, n_4418, n_4419);
  and g13914 (n9589, \a[14] , n_4419);
  not g13915 (n_4420, n9588);
  not g13916 (n_4421, n9589);
  and g13917 (n9590, n_4420, n_4421);
  and g13918 (n9591, n_4133, n_4135);
  and g13919 (n9592, n_4134, n_4135);
  not g13920 (n_4422, n9591);
  not g13921 (n_4423, n9592);
  and g13922 (n9593, n_4422, n_4423);
  not g13923 (n_4424, n9590);
  not g13924 (n_4425, n9593);
  and g13925 (n9594, n_4424, n_4425);
  not g13926 (n_4426, n9594);
  and g13927 (n9595, n_4424, n_4426);
  and g13928 (n9596, n_4425, n_4426);
  not g13929 (n_4427, n9595);
  not g13930 (n_4428, n9596);
  and g13931 (n9597, n_4427, n_4428);
  and g13932 (n9598, n9151, n9248);
  not g13933 (n_4429, n9598);
  and g13934 (n9599, n_4129, n_4429);
  and g13935 (n9600, n_306, n7101);
  and g13936 (n9601, n_308, n6402);
  and g13937 (n9602, n_307, n6951);
  not g13938 (n_4430, n9601);
  not g13939 (n_4431, n9602);
  and g13940 (n9603, n_4430, n_4431);
  not g13941 (n_4432, n9600);
  and g13942 (n9604, n_4432, n9603);
  and g13943 (n9605, n_1885, n9604);
  and g13944 (n9606, n_2498, n9604);
  not g13945 (n_4433, n9605);
  not g13946 (n_4434, n9606);
  and g13947 (n9607, n_4433, n_4434);
  not g13948 (n_4435, n9607);
  and g13949 (n9608, \a[14] , n_4435);
  and g13950 (n9609, n_652, n9607);
  not g13951 (n_4436, n9608);
  not g13952 (n_4437, n9609);
  and g13953 (n9610, n_4436, n_4437);
  not g13954 (n_4438, n9610);
  and g13955 (n9611, n9599, n_4438);
  not g13956 (n_4439, n9246);
  and g13957 (n9612, n9244, n_4439);
  not g13958 (n_4440, n9612);
  and g13959 (n9613, n_4126, n_4440);
  and g13960 (n9614, n_307, n7101);
  and g13961 (n9615, n_309, n6402);
  and g13962 (n9616, n_308, n6951);
  not g13963 (n_4441, n9615);
  not g13964 (n_4442, n9616);
  and g13965 (n9617, n_4441, n_4442);
  not g13966 (n_4443, n9614);
  and g13967 (n9618, n_4443, n9617);
  and g13968 (n9619, n_1885, n9618);
  and g13969 (n9620, n_2511, n9618);
  not g13970 (n_4444, n9619);
  not g13971 (n_4445, n9620);
  and g13972 (n9621, n_4444, n_4445);
  not g13973 (n_4446, n9621);
  and g13974 (n9622, \a[14] , n_4446);
  and g13975 (n9623, n_652, n9621);
  not g13976 (n_4447, n9622);
  not g13977 (n_4448, n9623);
  and g13978 (n9624, n_4447, n_4448);
  not g13979 (n_4449, n9624);
  and g13980 (n9625, n9613, n_4449);
  and g13981 (n9626, n9183, n9242);
  not g13982 (n_4450, n9626);
  and g13983 (n9627, n_4122, n_4450);
  and g13984 (n9628, n_308, n7101);
  and g13985 (n9629, n_310, n6402);
  and g13986 (n9630, n_309, n6951);
  not g13987 (n_4451, n9629);
  not g13988 (n_4452, n9630);
  and g13989 (n9631, n_4451, n_4452);
  not g13990 (n_4453, n9628);
  and g13991 (n9632, n_4453, n9631);
  and g13992 (n9633, n_1885, n9632);
  and g13993 (n9634, n_2839, n9632);
  not g13994 (n_4454, n9633);
  not g13995 (n_4455, n9634);
  and g13996 (n9635, n_4454, n_4455);
  not g13997 (n_4456, n9635);
  and g13998 (n9636, \a[14] , n_4456);
  and g13999 (n9637, n_652, n9635);
  not g14000 (n_4457, n9636);
  not g14001 (n_4458, n9637);
  and g14002 (n9638, n_4457, n_4458);
  not g14003 (n_4459, n9638);
  and g14004 (n9639, n9627, n_4459);
  and g14005 (n9640, n_309, n7101);
  and g14006 (n9641, n_311, n6402);
  and g14007 (n9642, n_310, n6951);
  and g14013 (n9645, n6397, n6541);
  not g14016 (n_4464, n9646);
  and g14017 (n9647, \a[14] , n_4464);
  not g14018 (n_4465, n9647);
  and g14019 (n9648, n_4464, n_4465);
  and g14020 (n9649, \a[14] , n_4465);
  not g14021 (n_4466, n9648);
  not g14022 (n_4467, n9649);
  and g14023 (n9650, n_4466, n_4467);
  not g14024 (n_4468, n9240);
  and g14025 (n9651, n9238, n_4468);
  not g14026 (n_4469, n9651);
  and g14027 (n9652, n_4119, n_4469);
  not g14028 (n_4470, n9650);
  and g14029 (n9653, n_4470, n9652);
  not g14030 (n_4471, n9653);
  and g14031 (n9654, n_4470, n_4471);
  and g14032 (n9655, n9652, n_4471);
  not g14033 (n_4472, n9654);
  not g14034 (n_4473, n9655);
  and g14035 (n9656, n_4472, n_4473);
  and g14036 (n9657, n_4112, n_4114);
  and g14037 (n9658, n_4113, n_4114);
  not g14038 (n_4474, n9657);
  not g14039 (n_4475, n9658);
  and g14040 (n9659, n_4474, n_4475);
  and g14041 (n9660, n_310, n7101);
  and g14042 (n9661, n_312, n6402);
  and g14043 (n9662, n_311, n6951);
  not g14044 (n_4476, n9661);
  not g14045 (n_4477, n9662);
  and g14046 (n9663, n_4476, n_4477);
  not g14047 (n_4478, n9660);
  and g14048 (n9664, n_4478, n9663);
  and g14049 (n9665, n_1885, n9664);
  and g14050 (n9666, n_3239, n9664);
  not g14051 (n_4479, n9665);
  not g14052 (n_4480, n9666);
  and g14053 (n9667, n_4479, n_4480);
  not g14054 (n_4481, n9667);
  and g14055 (n9668, \a[14] , n_4481);
  and g14056 (n9669, n_652, n9667);
  not g14057 (n_4482, n9668);
  not g14058 (n_4483, n9669);
  and g14059 (n9670, n_4482, n_4483);
  not g14060 (n_4484, n9659);
  not g14061 (n_4485, n9670);
  and g14062 (n9671, n_4484, n_4485);
  and g14063 (n9672, n_311, n7101);
  and g14064 (n9673, n_313, n6402);
  and g14065 (n9674, n_312, n6951);
  and g14071 (n9677, n6397, n6646);
  not g14074 (n_4490, n9678);
  and g14075 (n9679, \a[14] , n_4490);
  not g14076 (n_4491, n9679);
  and g14077 (n9680, n_4490, n_4491);
  and g14078 (n9681, \a[14] , n_4491);
  not g14079 (n_4492, n9680);
  not g14080 (n_4493, n9681);
  and g14081 (n9682, n_4492, n_4493);
  not g14082 (n_4494, n9209);
  and g14083 (n9683, n_4494, n9220);
  not g14084 (n_4495, n9221);
  not g14085 (n_4496, n9683);
  and g14086 (n9684, n_4495, n_4496);
  not g14087 (n_4497, n9682);
  and g14088 (n9685, n_4497, n9684);
  not g14089 (n_4498, n9685);
  and g14090 (n9686, n_4497, n_4498);
  and g14091 (n9687, n9684, n_4498);
  not g14092 (n_4499, n9686);
  not g14093 (n_4500, n9687);
  and g14094 (n9688, n_4499, n_4500);
  not g14095 (n_4501, n9208);
  and g14096 (n9689, n9206, n_4501);
  not g14097 (n_4502, n9689);
  and g14098 (n9690, n_4494, n_4502);
  and g14099 (n9691, n_312, n7101);
  and g14100 (n9692, n_314, n6402);
  and g14101 (n9693, n_313, n6951);
  not g14102 (n_4503, n9692);
  not g14103 (n_4504, n9693);
  and g14104 (n9694, n_4503, n_4504);
  not g14105 (n_4505, n9691);
  and g14106 (n9695, n_4505, n9694);
  and g14107 (n9696, n_1885, n9695);
  and g14108 (n9697, n_2891, n9695);
  not g14109 (n_4506, n9696);
  not g14110 (n_4507, n9697);
  and g14111 (n9698, n_4506, n_4507);
  not g14112 (n_4508, n9698);
  and g14113 (n9699, \a[14] , n_4508);
  and g14114 (n9700, n_652, n9698);
  not g14115 (n_4509, n9699);
  not g14116 (n_4510, n9700);
  and g14117 (n9701, n_4509, n_4510);
  not g14118 (n_4511, n9701);
  and g14119 (n9702, n9690, n_4511);
  and g14120 (n9703, n_316, n6951);
  and g14121 (n9704, n_315, n7101);
  not g14122 (n_4512, n9703);
  not g14123 (n_4513, n9704);
  and g14124 (n9705, n_4512, n_4513);
  and g14125 (n9706, n6397, n_2588);
  not g14126 (n_4514, n9706);
  and g14127 (n9707, n9705, n_4514);
  not g14128 (n_4515, n9707);
  and g14129 (n9708, \a[14] , n_4515);
  not g14130 (n_4516, n9708);
  and g14131 (n9709, \a[14] , n_4516);
  and g14132 (n9710, n_4515, n_4516);
  not g14133 (n_4517, n9709);
  not g14134 (n_4518, n9710);
  and g14135 (n9711, n_4517, n_4518);
  and g14136 (n9712, n_316, n_1881);
  not g14137 (n_4519, n9712);
  and g14138 (n9713, \a[14] , n_4519);
  not g14139 (n_4520, n9711);
  and g14140 (n9714, n_4520, n9713);
  and g14141 (n9715, n_314, n7101);
  and g14142 (n9716, n_316, n6402);
  and g14143 (n9717, n_315, n6951);
  not g14144 (n_4521, n9716);
  not g14145 (n_4522, n9717);
  and g14146 (n9718, n_4521, n_4522);
  not g14147 (n_4523, n9715);
  and g14148 (n9719, n_4523, n9718);
  and g14149 (n9720, n_1885, n9719);
  and g14150 (n9721, n_2612, n9719);
  not g14151 (n_4524, n9720);
  not g14152 (n_4525, n9721);
  and g14153 (n9722, n_4524, n_4525);
  not g14154 (n_4526, n9722);
  and g14155 (n9723, \a[14] , n_4526);
  and g14156 (n9724, n_652, n9722);
  not g14157 (n_4527, n9723);
  not g14158 (n_4528, n9724);
  and g14159 (n9725, n_4527, n_4528);
  not g14160 (n_4529, n9725);
  and g14161 (n9726, n9714, n_4529);
  and g14162 (n9727, n9207, n9726);
  not g14163 (n_4530, n9727);
  and g14164 (n9728, n9726, n_4530);
  and g14165 (n9729, n9207, n_4530);
  not g14166 (n_4531, n9728);
  not g14167 (n_4532, n9729);
  and g14168 (n9730, n_4531, n_4532);
  and g14169 (n9731, n_313, n7101);
  and g14170 (n9732, n_315, n6402);
  and g14171 (n9733, n_314, n6951);
  and g14177 (n9736, n6397, n6806);
  not g14180 (n_4537, n9737);
  and g14181 (n9738, \a[14] , n_4537);
  not g14182 (n_4538, n9738);
  and g14183 (n9739, \a[14] , n_4538);
  and g14184 (n9740, n_4537, n_4538);
  not g14185 (n_4539, n9739);
  not g14186 (n_4540, n9740);
  and g14187 (n9741, n_4539, n_4540);
  not g14188 (n_4541, n9730);
  not g14189 (n_4542, n9741);
  and g14190 (n9742, n_4541, n_4542);
  not g14191 (n_4543, n9742);
  and g14192 (n9743, n_4530, n_4543);
  not g14193 (n_4544, n9690);
  and g14194 (n9744, n_4544, n9701);
  not g14195 (n_4545, n9702);
  not g14196 (n_4546, n9744);
  and g14197 (n9745, n_4545, n_4546);
  not g14198 (n_4547, n9743);
  and g14199 (n9746, n_4547, n9745);
  not g14200 (n_4548, n9746);
  and g14201 (n9747, n_4545, n_4548);
  not g14202 (n_4549, n9688);
  not g14203 (n_4550, n9747);
  and g14204 (n9748, n_4549, n_4550);
  not g14205 (n_4551, n9748);
  and g14206 (n9749, n_4498, n_4551);
  and g14207 (n9750, n9659, n9670);
  not g14208 (n_4552, n9671);
  not g14209 (n_4553, n9750);
  and g14210 (n9751, n_4552, n_4553);
  not g14211 (n_4554, n9749);
  and g14212 (n9752, n_4554, n9751);
  not g14213 (n_4555, n9752);
  and g14214 (n9753, n_4552, n_4555);
  not g14215 (n_4556, n9656);
  not g14216 (n_4557, n9753);
  and g14217 (n9754, n_4556, n_4557);
  not g14218 (n_4558, n9754);
  and g14219 (n9755, n_4471, n_4558);
  not g14220 (n_4559, n9639);
  and g14221 (n9756, n9627, n_4559);
  and g14222 (n9757, n_4459, n_4559);
  not g14223 (n_4560, n9756);
  not g14224 (n_4561, n9757);
  and g14225 (n9758, n_4560, n_4561);
  not g14226 (n_4562, n9755);
  not g14227 (n_4563, n9758);
  and g14228 (n9759, n_4562, n_4563);
  not g14229 (n_4564, n9759);
  and g14230 (n9760, n_4559, n_4564);
  not g14231 (n_4565, n9625);
  and g14232 (n9761, n9613, n_4565);
  and g14233 (n9762, n_4449, n_4565);
  not g14234 (n_4566, n9761);
  not g14235 (n_4567, n9762);
  and g14236 (n9763, n_4566, n_4567);
  not g14237 (n_4568, n9760);
  not g14238 (n_4569, n9763);
  and g14239 (n9764, n_4568, n_4569);
  not g14240 (n_4570, n9764);
  and g14241 (n9765, n_4565, n_4570);
  not g14242 (n_4571, n9599);
  and g14243 (n9766, n_4571, n9610);
  not g14244 (n_4572, n9611);
  not g14245 (n_4573, n9766);
  and g14246 (n9767, n_4572, n_4573);
  not g14247 (n_4574, n9765);
  and g14248 (n9768, n_4574, n9767);
  not g14249 (n_4575, n9768);
  and g14250 (n9769, n_4572, n_4575);
  not g14251 (n_4576, n9597);
  not g14252 (n_4577, n9769);
  and g14253 (n9770, n_4576, n_4577);
  not g14254 (n_4578, n9770);
  and g14255 (n9771, n_4426, n_4578);
  not g14256 (n_4579, n9579);
  not g14257 (n_4580, n9771);
  and g14258 (n9772, n_4579, n_4580);
  not g14259 (n_4581, n9772);
  and g14260 (n9773, n_4411, n_4581);
  not g14261 (n_4582, n9561);
  not g14262 (n_4583, n9773);
  and g14263 (n9774, n_4582, n_4583);
  not g14264 (n_4584, n9774);
  and g14265 (n9775, n_4396, n_4584);
  not g14266 (n_4585, n9544);
  and g14267 (n9776, n9532, n_4585);
  and g14268 (n9777, n_4384, n_4585);
  not g14269 (n_4586, n9776);
  not g14270 (n_4587, n9777);
  and g14271 (n9778, n_4586, n_4587);
  not g14272 (n_4588, n9775);
  not g14273 (n_4589, n9778);
  and g14274 (n9779, n_4588, n_4589);
  not g14275 (n_4590, n9779);
  and g14276 (n9780, n_4585, n_4590);
  not g14277 (n_4591, n9530);
  and g14278 (n9781, n9518, n_4591);
  and g14279 (n9782, n_4374, n_4591);
  not g14280 (n_4592, n9781);
  not g14281 (n_4593, n9782);
  and g14282 (n9783, n_4592, n_4593);
  not g14283 (n_4594, n9780);
  not g14284 (n_4595, n9783);
  and g14285 (n9784, n_4594, n_4595);
  not g14286 (n_4596, n9784);
  and g14287 (n9785, n_4591, n_4596);
  not g14288 (n_4597, n9504);
  and g14289 (n9786, n_4597, n9515);
  not g14290 (n_4598, n9516);
  not g14291 (n_4599, n9786);
  and g14292 (n9787, n_4598, n_4599);
  not g14293 (n_4600, n9785);
  and g14294 (n9788, n_4600, n9787);
  not g14295 (n_4601, n9788);
  and g14296 (n9789, n_4598, n_4601);
  not g14297 (n_4602, n9502);
  not g14298 (n_4603, n9789);
  and g14299 (n9790, n_4602, n_4603);
  not g14300 (n_4604, n9790);
  and g14301 (n9791, n_4352, n_4604);
  not g14302 (n_4605, n9484);
  not g14303 (n_4606, n9791);
  and g14304 (n9792, n_4605, n_4606);
  not g14305 (n_4607, n9792);
  and g14306 (n9793, n_4337, n_4607);
  not g14307 (n_4608, n9467);
  and g14308 (n9794, n9455, n_4608);
  and g14309 (n9795, n_4325, n_4608);
  not g14310 (n_4609, n9794);
  not g14311 (n_4610, n9795);
  and g14312 (n9796, n_4609, n_4610);
  not g14313 (n_4611, n9793);
  not g14314 (n_4612, n9796);
  and g14315 (n9797, n_4611, n_4612);
  not g14316 (n_4613, n9797);
  and g14317 (n9798, n_4608, n_4613);
  not g14318 (n_4614, n9453);
  and g14319 (n9799, n9441, n_4614);
  and g14320 (n9800, n_4315, n_4614);
  not g14321 (n_4615, n9799);
  not g14322 (n_4616, n9800);
  and g14323 (n9801, n_4615, n_4616);
  not g14324 (n_4617, n9798);
  not g14325 (n_4618, n9801);
  and g14326 (n9802, n_4617, n_4618);
  not g14327 (n_4619, n9802);
  and g14328 (n9803, n_4614, n_4619);
  not g14329 (n_4620, n9439);
  and g14330 (n9804, n9427, n_4620);
  and g14331 (n9805, n_4305, n_4620);
  not g14332 (n_4621, n9804);
  not g14333 (n_4622, n9805);
  and g14334 (n9806, n_4621, n_4622);
  not g14335 (n_4623, n9803);
  not g14336 (n_4624, n9806);
  and g14337 (n9807, n_4623, n_4624);
  not g14338 (n_4625, n9807);
  and g14339 (n9808, n_4620, n_4625);
  not g14340 (n_4626, n9425);
  and g14341 (n9809, n9413, n_4626);
  and g14342 (n9810, n_4295, n_4626);
  not g14343 (n_4627, n9809);
  not g14344 (n_4628, n9810);
  and g14345 (n9811, n_4627, n_4628);
  not g14346 (n_4629, n9808);
  not g14347 (n_4630, n9811);
  and g14348 (n9812, n_4629, n_4630);
  not g14349 (n_4631, n9812);
  and g14350 (n9813, n_4626, n_4631);
  not g14351 (n_4632, n9411);
  and g14352 (n9814, n9399, n_4632);
  and g14353 (n9815, n_4285, n_4632);
  not g14354 (n_4633, n9814);
  not g14355 (n_4634, n9815);
  and g14356 (n9816, n_4633, n_4634);
  not g14357 (n_4635, n9813);
  not g14358 (n_4636, n9816);
  and g14359 (n9817, n_4635, n_4636);
  not g14360 (n_4637, n9817);
  and g14361 (n9818, n_4632, n_4637);
  not g14362 (n_4638, n9397);
  and g14363 (n9819, n9385, n_4638);
  and g14364 (n9820, n_4275, n_4638);
  not g14365 (n_4639, n9819);
  not g14366 (n_4640, n9820);
  and g14367 (n9821, n_4639, n_4640);
  not g14368 (n_4641, n9818);
  not g14369 (n_4642, n9821);
  and g14370 (n9822, n_4641, n_4642);
  not g14371 (n_4643, n9822);
  and g14372 (n9823, n_4638, n_4643);
  not g14373 (n_4644, n9383);
  and g14374 (n9824, n9371, n_4644);
  and g14375 (n9825, n_4265, n_4644);
  not g14376 (n_4645, n9824);
  not g14377 (n_4646, n9825);
  and g14378 (n9826, n_4645, n_4646);
  not g14379 (n_4647, n9823);
  not g14380 (n_4648, n9826);
  and g14381 (n9827, n_4647, n_4648);
  not g14382 (n_4649, n9827);
  and g14383 (n9828, n_4644, n_4649);
  not g14384 (n_4650, n9309);
  and g14385 (n9829, n9307, n_4650);
  not g14386 (n_4651, n9829);
  and g14387 (n9830, n_4203, n_4651);
  not g14388 (n_4652, n9828);
  and g14389 (n9831, n_4652, n9830);
  and g14390 (n9832, n_485, n7983);
  and g14391 (n9833, n_415, n7291);
  and g14392 (n9834, n_484, n7632);
  and g14398 (n9837, n4084, n7294);
  not g14401 (n_4657, n9838);
  and g14402 (n9839, \a[11] , n_4657);
  not g14403 (n_4658, n9839);
  and g14404 (n9840, n_4657, n_4658);
  and g14405 (n9841, \a[11] , n_4658);
  not g14406 (n_4659, n9840);
  not g14407 (n_4660, n9841);
  and g14408 (n9842, n_4659, n_4660);
  not g14409 (n_4661, n9830);
  and g14410 (n9843, n9828, n_4661);
  not g14411 (n_4662, n9831);
  not g14412 (n_4663, n9843);
  and g14413 (n9844, n_4662, n_4663);
  not g14414 (n_4664, n9842);
  and g14415 (n9845, n_4664, n9844);
  not g14416 (n_4665, n9845);
  and g14417 (n9846, n_4662, n_4665);
  not g14418 (n_4666, n9369);
  not g14419 (n_4667, n9846);
  and g14420 (n9847, n_4666, n_4667);
  and g14421 (n9848, n9369, n9846);
  not g14422 (n_4668, n9847);
  not g14423 (n_4669, n9848);
  and g14424 (n9849, n_4668, n_4669);
  and g14425 (n9850, n_566, n9331);
  and g14426 (n9851, n_535, n8418);
  and g14427 (n9852, n_565, n8860);
  and g14433 (n9855, n4477, n8421);
  not g14436 (n_4674, n9856);
  and g14437 (n9857, \a[8] , n_4674);
  not g14438 (n_4675, n9857);
  and g14439 (n9858, \a[8] , n_4675);
  and g14440 (n9859, n_4674, n_4675);
  not g14441 (n_4676, n9858);
  not g14442 (n_4677, n9859);
  and g14443 (n9860, n_4676, n_4677);
  not g14444 (n_4678, n9860);
  and g14445 (n9861, n9849, n_4678);
  not g14446 (n_4679, n9861);
  and g14447 (n9862, n_4668, n_4679);
  and g14448 (n9863, n_9, \a[4] );
  and g14449 (n9864, \a[3] , n_4);
  not g14450 (n_4680, n9863);
  not g14451 (n_4681, n9864);
  and g14452 (n9865, n_4680, n_4681);
  not g14453 (n_4682, n67);
  and g14454 (n9866, n_4682, n70);
  and g14455 (n9867, n9865, n9866);
  and g14456 (n9868, n_712, n9867);
  not g14457 (n_4683, n9868);
  and g14458 (n9869, n_729, n_4683);
  and g14459 (n9870, n_4682, n_13);
  not g14460 (n_4684, n9870);
  and g14461 (n9871, n_4683, n_4684);
  not g14462 (n_4685, n9869);
  not g14463 (n_4686, n9871);
  and g14464 (n9872, n_4685, n_4686);
  not g14465 (n_4687, n9872);
  and g14466 (n9873, \a[5] , n_4687);
  and g14467 (n9874, n_3, n9872);
  not g14468 (n_4688, n9873);
  not g14469 (n_4689, n9874);
  and g14470 (n9875, n_4688, n_4689);
  not g14471 (n_4690, n9862);
  not g14472 (n_4691, n9875);
  and g14473 (n9876, n_4690, n_4691);
  and g14474 (n9877, n9330, n_4231);
  and g14475 (n9878, n_4230, n_4231);
  not g14476 (n_4692, n9877);
  not g14477 (n_4693, n9878);
  and g14478 (n9879, n_4692, n_4693);
  and g14479 (n9880, n9862, n9875);
  not g14480 (n_4694, n9876);
  not g14481 (n_4695, n9880);
  and g14482 (n9881, n_4694, n_4695);
  not g14483 (n_4696, n9879);
  and g14484 (n9882, n_4696, n9881);
  not g14485 (n_4697, n9882);
  and g14486 (n9883, n_4694, n_4697);
  not g14487 (n_4698, n9361);
  and g14488 (n9884, n_4244, n_4698);
  and g14489 (n9885, n_4243, n9884);
  not g14490 (n_4699, n9885);
  and g14491 (n9886, n_4249, n_4699);
  not g14492 (n_4700, n9883);
  and g14493 (n9887, n_4700, n9886);
  and g14494 (n9888, n_4696, n_4697);
  and g14495 (n9889, n9881, n_4697);
  not g14496 (n_4701, n9888);
  not g14497 (n_4702, n9889);
  and g14498 (n9890, n_4701, n_4702);
  and g14499 (n9891, n_484, n7983);
  and g14500 (n9892, n_236, n7291);
  and g14501 (n9893, n_415, n7632);
  and g14507 (n9896, n3715, n7294);
  not g14510 (n_4707, n9897);
  and g14511 (n9898, \a[11] , n_4707);
  not g14512 (n_4708, n9898);
  and g14513 (n9899, n_4707, n_4708);
  and g14514 (n9900, \a[11] , n_4708);
  not g14515 (n_4709, n9899);
  not g14516 (n_4710, n9900);
  and g14517 (n9901, n_4709, n_4710);
  and g14518 (n9902, n_4647, n_4649);
  and g14519 (n9903, n_4648, n_4649);
  not g14520 (n_4711, n9902);
  not g14521 (n_4712, n9903);
  and g14522 (n9904, n_4711, n_4712);
  not g14523 (n_4713, n9901);
  not g14524 (n_4714, n9904);
  and g14525 (n9905, n_4713, n_4714);
  not g14526 (n_4715, n9905);
  and g14527 (n9906, n_4713, n_4715);
  and g14528 (n9907, n_4714, n_4715);
  not g14529 (n_4716, n9906);
  not g14530 (n_4717, n9907);
  and g14531 (n9908, n_4716, n_4717);
  and g14532 (n9909, n_415, n7983);
  and g14533 (n9910, n_237, n7291);
  and g14534 (n9911, n_236, n7632);
  and g14540 (n9914, n3018, n7294);
  not g14543 (n_4722, n9915);
  and g14544 (n9916, \a[11] , n_4722);
  not g14545 (n_4723, n9916);
  and g14546 (n9917, n_4722, n_4723);
  and g14547 (n9918, \a[11] , n_4723);
  not g14548 (n_4724, n9917);
  not g14549 (n_4725, n9918);
  and g14550 (n9919, n_4724, n_4725);
  and g14551 (n9920, n_4641, n_4643);
  and g14552 (n9921, n_4642, n_4643);
  not g14553 (n_4726, n9920);
  not g14554 (n_4727, n9921);
  and g14555 (n9922, n_4726, n_4727);
  not g14556 (n_4728, n9919);
  not g14557 (n_4729, n9922);
  and g14558 (n9923, n_4728, n_4729);
  not g14559 (n_4730, n9923);
  and g14560 (n9924, n_4728, n_4730);
  and g14561 (n9925, n_4729, n_4730);
  not g14562 (n_4731, n9924);
  not g14563 (n_4732, n9925);
  and g14564 (n9926, n_4731, n_4732);
  and g14565 (n9927, n_236, n7983);
  and g14566 (n9928, n_260, n7291);
  and g14567 (n9929, n_237, n7632);
  and g14573 (n9932, n3347, n7294);
  not g14576 (n_4737, n9933);
  and g14577 (n9934, \a[11] , n_4737);
  not g14578 (n_4738, n9934);
  and g14579 (n9935, n_4737, n_4738);
  and g14580 (n9936, \a[11] , n_4738);
  not g14581 (n_4739, n9935);
  not g14582 (n_4740, n9936);
  and g14583 (n9937, n_4739, n_4740);
  and g14584 (n9938, n_4635, n_4637);
  and g14585 (n9939, n_4636, n_4637);
  not g14586 (n_4741, n9938);
  not g14587 (n_4742, n9939);
  and g14588 (n9940, n_4741, n_4742);
  not g14589 (n_4743, n9937);
  not g14590 (n_4744, n9940);
  and g14591 (n9941, n_4743, n_4744);
  not g14592 (n_4745, n9941);
  and g14593 (n9942, n_4743, n_4745);
  and g14594 (n9943, n_4744, n_4745);
  not g14595 (n_4746, n9942);
  not g14596 (n_4747, n9943);
  and g14597 (n9944, n_4746, n_4747);
  and g14598 (n9945, n_237, n7983);
  and g14599 (n9946, n_275, n7291);
  and g14600 (n9947, n_260, n7632);
  and g14606 (n9950, n3331, n7294);
  not g14609 (n_4752, n9951);
  and g14610 (n9952, \a[11] , n_4752);
  not g14611 (n_4753, n9952);
  and g14612 (n9953, n_4752, n_4753);
  and g14613 (n9954, \a[11] , n_4753);
  not g14614 (n_4754, n9953);
  not g14615 (n_4755, n9954);
  and g14616 (n9955, n_4754, n_4755);
  and g14617 (n9956, n_4629, n_4631);
  and g14618 (n9957, n_4630, n_4631);
  not g14619 (n_4756, n9956);
  not g14620 (n_4757, n9957);
  and g14621 (n9958, n_4756, n_4757);
  not g14622 (n_4758, n9955);
  not g14623 (n_4759, n9958);
  and g14624 (n9959, n_4758, n_4759);
  not g14625 (n_4760, n9959);
  and g14626 (n9960, n_4758, n_4760);
  and g14627 (n9961, n_4759, n_4760);
  not g14628 (n_4761, n9960);
  not g14629 (n_4762, n9961);
  and g14630 (n9962, n_4761, n_4762);
  and g14631 (n9963, n_260, n7983);
  and g14632 (n9964, n_281, n7291);
  and g14633 (n9965, n_275, n7632);
  and g14639 (n9968, n4179, n7294);
  not g14642 (n_4767, n9969);
  and g14643 (n9970, \a[11] , n_4767);
  not g14644 (n_4768, n9970);
  and g14645 (n9971, n_4767, n_4768);
  and g14646 (n9972, \a[11] , n_4768);
  not g14647 (n_4769, n9971);
  not g14648 (n_4770, n9972);
  and g14649 (n9973, n_4769, n_4770);
  and g14650 (n9974, n_4623, n_4625);
  and g14651 (n9975, n_4624, n_4625);
  not g14652 (n_4771, n9974);
  not g14653 (n_4772, n9975);
  and g14654 (n9976, n_4771, n_4772);
  not g14655 (n_4773, n9973);
  not g14656 (n_4774, n9976);
  and g14657 (n9977, n_4773, n_4774);
  not g14658 (n_4775, n9977);
  and g14659 (n9978, n_4773, n_4775);
  and g14660 (n9979, n_4774, n_4775);
  not g14661 (n_4776, n9978);
  not g14662 (n_4777, n9979);
  and g14663 (n9980, n_4776, n_4777);
  and g14664 (n9981, n_275, n7983);
  and g14665 (n9982, n_286, n7291);
  and g14666 (n9983, n_281, n7632);
  and g14672 (n9986, n4204, n7294);
  not g14675 (n_4782, n9987);
  and g14676 (n9988, \a[11] , n_4782);
  not g14677 (n_4783, n9988);
  and g14678 (n9989, n_4782, n_4783);
  and g14679 (n9990, \a[11] , n_4783);
  not g14680 (n_4784, n9989);
  not g14681 (n_4785, n9990);
  and g14682 (n9991, n_4784, n_4785);
  and g14683 (n9992, n_4617, n_4619);
  and g14684 (n9993, n_4618, n_4619);
  not g14685 (n_4786, n9992);
  not g14686 (n_4787, n9993);
  and g14687 (n9994, n_4786, n_4787);
  not g14688 (n_4788, n9991);
  not g14689 (n_4789, n9994);
  and g14690 (n9995, n_4788, n_4789);
  not g14691 (n_4790, n9995);
  and g14692 (n9996, n_4788, n_4790);
  and g14693 (n9997, n_4789, n_4790);
  not g14694 (n_4791, n9996);
  not g14695 (n_4792, n9997);
  and g14696 (n9998, n_4791, n_4792);
  and g14697 (n9999, n_281, n7983);
  and g14698 (n10000, n_293, n7291);
  and g14699 (n10001, n_286, n7632);
  and g14705 (n10004, n4633, n7294);
  not g14708 (n_4797, n10005);
  and g14709 (n10006, \a[11] , n_4797);
  not g14710 (n_4798, n10006);
  and g14711 (n10007, n_4797, n_4798);
  and g14712 (n10008, \a[11] , n_4798);
  not g14713 (n_4799, n10007);
  not g14714 (n_4800, n10008);
  and g14715 (n10009, n_4799, n_4800);
  and g14716 (n10010, n_4611, n_4613);
  and g14717 (n10011, n_4612, n_4613);
  not g14718 (n_4801, n10010);
  not g14719 (n_4802, n10011);
  and g14720 (n10012, n_4801, n_4802);
  not g14721 (n_4803, n10009);
  not g14722 (n_4804, n10012);
  and g14723 (n10013, n_4803, n_4804);
  not g14724 (n_4805, n10013);
  and g14725 (n10014, n_4803, n_4805);
  and g14726 (n10015, n_4804, n_4805);
  not g14727 (n_4806, n10014);
  not g14728 (n_4807, n10015);
  and g14729 (n10016, n_4806, n_4807);
  and g14730 (n10017, n9484, n9791);
  not g14731 (n_4808, n10017);
  and g14732 (n10018, n_4607, n_4808);
  and g14733 (n10019, n_286, n7983);
  and g14734 (n10020, n_295, n7291);
  and g14735 (n10021, n_293, n7632);
  not g14736 (n_4809, n10020);
  not g14737 (n_4810, n10021);
  and g14738 (n10022, n_4809, n_4810);
  not g14739 (n_4811, n10019);
  and g14740 (n10023, n_4811, n10022);
  and g14741 (n10024, n_2446, n10023);
  and g14742 (n10025, n_1134, n10023);
  not g14743 (n_4812, n10024);
  not g14744 (n_4813, n10025);
  and g14745 (n10026, n_4812, n_4813);
  not g14746 (n_4814, n10026);
  and g14747 (n10027, \a[11] , n_4814);
  and g14748 (n10028, n_1071, n10026);
  not g14749 (n_4815, n10027);
  not g14750 (n_4816, n10028);
  and g14751 (n10029, n_4815, n_4816);
  not g14752 (n_4817, n10029);
  and g14753 (n10030, n10018, n_4817);
  and g14754 (n10031, n9502, n9789);
  not g14755 (n_4818, n10031);
  and g14756 (n10032, n_4604, n_4818);
  and g14757 (n10033, n_293, n7983);
  and g14758 (n10034, n_298, n7291);
  and g14759 (n10035, n_295, n7632);
  not g14760 (n_4819, n10034);
  not g14761 (n_4820, n10035);
  and g14762 (n10036, n_4819, n_4820);
  not g14763 (n_4821, n10033);
  and g14764 (n10037, n_4821, n10036);
  and g14765 (n10038, n_2446, n10037);
  and g14766 (n10039, n_1789, n10037);
  not g14767 (n_4822, n10038);
  not g14768 (n_4823, n10039);
  and g14769 (n10040, n_4822, n_4823);
  not g14770 (n_4824, n10040);
  and g14771 (n10041, \a[11] , n_4824);
  and g14772 (n10042, n_1071, n10040);
  not g14773 (n_4825, n10041);
  not g14774 (n_4826, n10042);
  and g14775 (n10043, n_4825, n_4826);
  not g14776 (n_4827, n10043);
  and g14777 (n10044, n10032, n_4827);
  and g14778 (n10045, n_295, n7983);
  and g14779 (n10046, n_299, n7291);
  and g14780 (n10047, n_298, n7632);
  and g14786 (n10050, n4848, n7294);
  not g14789 (n_4832, n10051);
  and g14790 (n10052, \a[11] , n_4832);
  not g14791 (n_4833, n10052);
  and g14792 (n10053, n_4832, n_4833);
  and g14793 (n10054, \a[11] , n_4833);
  not g14794 (n_4834, n10053);
  not g14795 (n_4835, n10054);
  and g14796 (n10055, n_4834, n_4835);
  not g14797 (n_4836, n9787);
  and g14798 (n10056, n9785, n_4836);
  not g14799 (n_4837, n10056);
  and g14800 (n10057, n_4601, n_4837);
  not g14801 (n_4838, n10055);
  and g14802 (n10058, n_4838, n10057);
  not g14803 (n_4839, n10058);
  and g14804 (n10059, n_4838, n_4839);
  and g14805 (n10060, n10057, n_4839);
  not g14806 (n_4840, n10059);
  not g14807 (n_4841, n10060);
  and g14808 (n10061, n_4840, n_4841);
  and g14809 (n10062, n_298, n7983);
  and g14810 (n10063, n_300, n7291);
  and g14811 (n10064, n_299, n7632);
  and g14817 (n10067, n5114, n7294);
  not g14820 (n_4846, n10068);
  and g14821 (n10069, \a[11] , n_4846);
  not g14822 (n_4847, n10069);
  and g14823 (n10070, n_4846, n_4847);
  and g14824 (n10071, \a[11] , n_4847);
  not g14825 (n_4848, n10070);
  not g14826 (n_4849, n10071);
  and g14827 (n10072, n_4848, n_4849);
  and g14828 (n10073, n_4594, n_4596);
  and g14829 (n10074, n_4595, n_4596);
  not g14830 (n_4850, n10073);
  not g14831 (n_4851, n10074);
  and g14832 (n10075, n_4850, n_4851);
  not g14833 (n_4852, n10072);
  not g14834 (n_4853, n10075);
  and g14835 (n10076, n_4852, n_4853);
  not g14836 (n_4854, n10076);
  and g14837 (n10077, n_4852, n_4854);
  and g14838 (n10078, n_4853, n_4854);
  not g14839 (n_4855, n10077);
  not g14840 (n_4856, n10078);
  and g14841 (n10079, n_4855, n_4856);
  and g14842 (n10080, n_299, n7983);
  and g14843 (n10081, n_301, n7291);
  and g14844 (n10082, n_300, n7632);
  and g14850 (n10085, n5139, n7294);
  not g14853 (n_4861, n10086);
  and g14854 (n10087, \a[11] , n_4861);
  not g14855 (n_4862, n10087);
  and g14856 (n10088, n_4861, n_4862);
  and g14857 (n10089, \a[11] , n_4862);
  not g14858 (n_4863, n10088);
  not g14859 (n_4864, n10089);
  and g14860 (n10090, n_4863, n_4864);
  and g14861 (n10091, n_4588, n_4590);
  and g14862 (n10092, n_4589, n_4590);
  not g14863 (n_4865, n10091);
  not g14864 (n_4866, n10092);
  and g14865 (n10093, n_4865, n_4866);
  not g14866 (n_4867, n10090);
  not g14867 (n_4868, n10093);
  and g14868 (n10094, n_4867, n_4868);
  not g14869 (n_4869, n10094);
  and g14870 (n10095, n_4867, n_4869);
  and g14871 (n10096, n_4868, n_4869);
  not g14872 (n_4870, n10095);
  not g14873 (n_4871, n10096);
  and g14874 (n10097, n_4870, n_4871);
  and g14875 (n10098, n9561, n9773);
  not g14876 (n_4872, n10098);
  and g14877 (n10099, n_4584, n_4872);
  and g14878 (n10100, n_300, n7983);
  and g14879 (n10101, n_302, n7291);
  and g14880 (n10102, n_301, n7632);
  not g14881 (n_4873, n10101);
  not g14882 (n_4874, n10102);
  and g14883 (n10103, n_4873, n_4874);
  not g14884 (n_4875, n10100);
  and g14885 (n10104, n_4875, n10103);
  and g14886 (n10105, n_2446, n10104);
  and g14887 (n10106, n_1801, n10104);
  not g14888 (n_4876, n10105);
  not g14889 (n_4877, n10106);
  and g14890 (n10107, n_4876, n_4877);
  not g14891 (n_4878, n10107);
  and g14892 (n10108, \a[11] , n_4878);
  and g14893 (n10109, n_1071, n10107);
  not g14894 (n_4879, n10108);
  not g14895 (n_4880, n10109);
  and g14896 (n10110, n_4879, n_4880);
  not g14897 (n_4881, n10110);
  and g14898 (n10111, n10099, n_4881);
  and g14899 (n10112, n9579, n9771);
  not g14900 (n_4882, n10112);
  and g14901 (n10113, n_4581, n_4882);
  and g14902 (n10114, n_301, n7983);
  and g14903 (n10115, n_303, n7291);
  and g14904 (n10116, n_302, n7632);
  not g14905 (n_4883, n10115);
  not g14906 (n_4884, n10116);
  and g14907 (n10117, n_4883, n_4884);
  not g14908 (n_4885, n10114);
  and g14909 (n10118, n_4885, n10117);
  and g14910 (n10119, n_2446, n10118);
  and g14911 (n10120, n_1672, n10118);
  not g14912 (n_4886, n10119);
  not g14913 (n_4887, n10120);
  and g14914 (n10121, n_4886, n_4887);
  not g14915 (n_4888, n10121);
  and g14916 (n10122, \a[11] , n_4888);
  and g14917 (n10123, n_1071, n10121);
  not g14918 (n_4889, n10122);
  not g14919 (n_4890, n10123);
  and g14920 (n10124, n_4889, n_4890);
  not g14921 (n_4891, n10124);
  and g14922 (n10125, n10113, n_4891);
  and g14923 (n10126, n9597, n9769);
  not g14924 (n_4892, n10126);
  and g14925 (n10127, n_4578, n_4892);
  and g14926 (n10128, n_302, n7983);
  and g14927 (n10129, n_304, n7291);
  and g14928 (n10130, n_303, n7632);
  not g14929 (n_4893, n10129);
  not g14930 (n_4894, n10130);
  and g14931 (n10131, n_4893, n_4894);
  not g14932 (n_4895, n10128);
  and g14933 (n10132, n_4895, n10131);
  and g14934 (n10133, n_2446, n10132);
  and g14935 (n10134, n_3507, n10132);
  not g14936 (n_4896, n10133);
  not g14937 (n_4897, n10134);
  and g14938 (n10135, n_4896, n_4897);
  not g14939 (n_4898, n10135);
  and g14940 (n10136, \a[11] , n_4898);
  and g14941 (n10137, n_1071, n10135);
  not g14942 (n_4899, n10136);
  not g14943 (n_4900, n10137);
  and g14944 (n10138, n_4899, n_4900);
  not g14945 (n_4901, n10138);
  and g14946 (n10139, n10127, n_4901);
  and g14947 (n10140, n_303, n7983);
  and g14948 (n10141, n_305, n7291);
  and g14949 (n10142, n_304, n7632);
  and g14955 (n10145, n6007, n7294);
  not g14958 (n_4906, n10146);
  and g14959 (n10147, \a[11] , n_4906);
  not g14960 (n_4907, n10147);
  and g14961 (n10148, n_4906, n_4907);
  and g14962 (n10149, \a[11] , n_4907);
  not g14963 (n_4908, n10148);
  not g14964 (n_4909, n10149);
  and g14965 (n10150, n_4908, n_4909);
  not g14966 (n_4910, n9767);
  and g14967 (n10151, n9765, n_4910);
  not g14968 (n_4911, n10151);
  and g14969 (n10152, n_4575, n_4911);
  not g14970 (n_4912, n10150);
  and g14971 (n10153, n_4912, n10152);
  not g14972 (n_4913, n10153);
  and g14973 (n10154, n_4912, n_4913);
  and g14974 (n10155, n10152, n_4913);
  not g14975 (n_4914, n10154);
  not g14976 (n_4915, n10155);
  and g14977 (n10156, n_4914, n_4915);
  and g14978 (n10157, n_304, n7983);
  and g14979 (n10158, n_306, n7291);
  and g14980 (n10159, n_305, n7632);
  and g14986 (n10162, n5834, n7294);
  not g14989 (n_4920, n10163);
  and g14990 (n10164, \a[11] , n_4920);
  not g14991 (n_4921, n10164);
  and g14992 (n10165, n_4920, n_4921);
  and g14993 (n10166, \a[11] , n_4921);
  not g14994 (n_4922, n10165);
  not g14995 (n_4923, n10166);
  and g14996 (n10167, n_4922, n_4923);
  and g14997 (n10168, n_4568, n_4570);
  and g14998 (n10169, n_4569, n_4570);
  not g14999 (n_4924, n10168);
  not g15000 (n_4925, n10169);
  and g15001 (n10170, n_4924, n_4925);
  not g15002 (n_4926, n10167);
  not g15003 (n_4927, n10170);
  and g15004 (n10171, n_4926, n_4927);
  not g15005 (n_4928, n10171);
  and g15006 (n10172, n_4926, n_4928);
  and g15007 (n10173, n_4927, n_4928);
  not g15008 (n_4929, n10172);
  not g15009 (n_4930, n10173);
  and g15010 (n10174, n_4929, n_4930);
  and g15011 (n10175, n_305, n7983);
  and g15012 (n10176, n_307, n7291);
  and g15013 (n10177, n_306, n7632);
  and g15019 (n10180, n6143, n7294);
  not g15022 (n_4935, n10181);
  and g15023 (n10182, \a[11] , n_4935);
  not g15024 (n_4936, n10182);
  and g15025 (n10183, n_4935, n_4936);
  and g15026 (n10184, \a[11] , n_4936);
  not g15027 (n_4937, n10183);
  not g15028 (n_4938, n10184);
  and g15029 (n10185, n_4937, n_4938);
  and g15030 (n10186, n_4562, n_4564);
  and g15031 (n10187, n_4563, n_4564);
  not g15032 (n_4939, n10186);
  not g15033 (n_4940, n10187);
  and g15034 (n10188, n_4939, n_4940);
  not g15035 (n_4941, n10185);
  not g15036 (n_4942, n10188);
  and g15037 (n10189, n_4941, n_4942);
  not g15038 (n_4943, n10189);
  and g15039 (n10190, n_4941, n_4943);
  and g15040 (n10191, n_4942, n_4943);
  not g15041 (n_4944, n10190);
  not g15042 (n_4945, n10191);
  and g15043 (n10192, n_4944, n_4945);
  and g15044 (n10193, n9656, n9753);
  not g15045 (n_4946, n10193);
  and g15046 (n10194, n_4558, n_4946);
  and g15047 (n10195, n_306, n7983);
  and g15048 (n10196, n_308, n7291);
  and g15049 (n10197, n_307, n7632);
  not g15050 (n_4947, n10196);
  not g15051 (n_4948, n10197);
  and g15052 (n10198, n_4947, n_4948);
  not g15053 (n_4949, n10195);
  and g15054 (n10199, n_4949, n10198);
  and g15055 (n10200, n_2446, n10199);
  and g15056 (n10201, n_2498, n10199);
  not g15057 (n_4950, n10200);
  not g15058 (n_4951, n10201);
  and g15059 (n10202, n_4950, n_4951);
  not g15060 (n_4952, n10202);
  and g15061 (n10203, \a[11] , n_4952);
  and g15062 (n10204, n_1071, n10202);
  not g15063 (n_4953, n10203);
  not g15064 (n_4954, n10204);
  and g15065 (n10205, n_4953, n_4954);
  not g15066 (n_4955, n10205);
  and g15067 (n10206, n10194, n_4955);
  not g15068 (n_4956, n9751);
  and g15069 (n10207, n9749, n_4956);
  not g15070 (n_4957, n10207);
  and g15071 (n10208, n_4555, n_4957);
  and g15072 (n10209, n_307, n7983);
  and g15073 (n10210, n_309, n7291);
  and g15074 (n10211, n_308, n7632);
  not g15075 (n_4958, n10210);
  not g15076 (n_4959, n10211);
  and g15077 (n10212, n_4958, n_4959);
  not g15078 (n_4960, n10209);
  and g15079 (n10213, n_4960, n10212);
  and g15080 (n10214, n_2446, n10213);
  and g15081 (n10215, n_2511, n10213);
  not g15082 (n_4961, n10214);
  not g15083 (n_4962, n10215);
  and g15084 (n10216, n_4961, n_4962);
  not g15085 (n_4963, n10216);
  and g15086 (n10217, \a[11] , n_4963);
  and g15087 (n10218, n_1071, n10216);
  not g15088 (n_4964, n10217);
  not g15089 (n_4965, n10218);
  and g15090 (n10219, n_4964, n_4965);
  not g15091 (n_4966, n10219);
  and g15092 (n10220, n10208, n_4966);
  and g15093 (n10221, n9688, n9747);
  not g15094 (n_4967, n10221);
  and g15095 (n10222, n_4551, n_4967);
  and g15096 (n10223, n_308, n7983);
  and g15097 (n10224, n_310, n7291);
  and g15098 (n10225, n_309, n7632);
  not g15099 (n_4968, n10224);
  not g15100 (n_4969, n10225);
  and g15101 (n10226, n_4968, n_4969);
  not g15102 (n_4970, n10223);
  and g15103 (n10227, n_4970, n10226);
  and g15104 (n10228, n_2446, n10227);
  and g15105 (n10229, n_2839, n10227);
  not g15106 (n_4971, n10228);
  not g15107 (n_4972, n10229);
  and g15108 (n10230, n_4971, n_4972);
  not g15109 (n_4973, n10230);
  and g15110 (n10231, \a[11] , n_4973);
  and g15111 (n10232, n_1071, n10230);
  not g15112 (n_4974, n10231);
  not g15113 (n_4975, n10232);
  and g15114 (n10233, n_4974, n_4975);
  not g15115 (n_4976, n10233);
  and g15116 (n10234, n10222, n_4976);
  and g15117 (n10235, n_309, n7983);
  and g15118 (n10236, n_311, n7291);
  and g15119 (n10237, n_310, n7632);
  and g15125 (n10240, n6541, n7294);
  not g15128 (n_4981, n10241);
  and g15129 (n10242, \a[11] , n_4981);
  not g15130 (n_4982, n10242);
  and g15131 (n10243, n_4981, n_4982);
  and g15132 (n10244, \a[11] , n_4982);
  not g15133 (n_4983, n10243);
  not g15134 (n_4984, n10244);
  and g15135 (n10245, n_4983, n_4984);
  not g15136 (n_4985, n9745);
  and g15137 (n10246, n9743, n_4985);
  not g15138 (n_4986, n10246);
  and g15139 (n10247, n_4548, n_4986);
  not g15140 (n_4987, n10245);
  and g15141 (n10248, n_4987, n10247);
  not g15142 (n_4988, n10248);
  and g15143 (n10249, n_4987, n_4988);
  and g15144 (n10250, n10247, n_4988);
  not g15145 (n_4989, n10249);
  not g15146 (n_4990, n10250);
  and g15147 (n10251, n_4989, n_4990);
  and g15148 (n10252, n_4541, n_4543);
  and g15149 (n10253, n_4542, n_4543);
  not g15150 (n_4991, n10252);
  not g15151 (n_4992, n10253);
  and g15152 (n10254, n_4991, n_4992);
  and g15153 (n10255, n_310, n7983);
  and g15154 (n10256, n_312, n7291);
  and g15155 (n10257, n_311, n7632);
  not g15156 (n_4993, n10256);
  not g15157 (n_4994, n10257);
  and g15158 (n10258, n_4993, n_4994);
  not g15159 (n_4995, n10255);
  and g15160 (n10259, n_4995, n10258);
  and g15161 (n10260, n_2446, n10259);
  and g15162 (n10261, n_3239, n10259);
  not g15163 (n_4996, n10260);
  not g15164 (n_4997, n10261);
  and g15165 (n10262, n_4996, n_4997);
  not g15166 (n_4998, n10262);
  and g15167 (n10263, \a[11] , n_4998);
  and g15168 (n10264, n_1071, n10262);
  not g15169 (n_4999, n10263);
  not g15170 (n_5000, n10264);
  and g15171 (n10265, n_4999, n_5000);
  not g15172 (n_5001, n10254);
  not g15173 (n_5002, n10265);
  and g15174 (n10266, n_5001, n_5002);
  and g15175 (n10267, n_311, n7983);
  and g15176 (n10268, n_313, n7291);
  and g15177 (n10269, n_312, n7632);
  and g15183 (n10272, n6646, n7294);
  not g15186 (n_5007, n10273);
  and g15187 (n10274, \a[11] , n_5007);
  not g15188 (n_5008, n10274);
  and g15189 (n10275, n_5007, n_5008);
  and g15190 (n10276, \a[11] , n_5008);
  not g15191 (n_5009, n10275);
  not g15192 (n_5010, n10276);
  and g15193 (n10277, n_5009, n_5010);
  not g15194 (n_5011, n9714);
  and g15195 (n10278, n_5011, n9725);
  not g15196 (n_5012, n9726);
  not g15197 (n_5013, n10278);
  and g15198 (n10279, n_5012, n_5013);
  not g15199 (n_5014, n10277);
  and g15200 (n10280, n_5014, n10279);
  not g15201 (n_5015, n10280);
  and g15202 (n10281, n_5014, n_5015);
  and g15203 (n10282, n10279, n_5015);
  not g15204 (n_5016, n10281);
  not g15205 (n_5017, n10282);
  and g15206 (n10283, n_5016, n_5017);
  not g15207 (n_5018, n9713);
  and g15208 (n10284, n9711, n_5018);
  not g15209 (n_5019, n10284);
  and g15210 (n10285, n_5011, n_5019);
  and g15211 (n10286, n_312, n7983);
  and g15212 (n10287, n_314, n7291);
  and g15213 (n10288, n_313, n7632);
  not g15214 (n_5020, n10287);
  not g15215 (n_5021, n10288);
  and g15216 (n10289, n_5020, n_5021);
  not g15217 (n_5022, n10286);
  and g15218 (n10290, n_5022, n10289);
  and g15219 (n10291, n_2446, n10290);
  and g15220 (n10292, n_2891, n10290);
  not g15221 (n_5023, n10291);
  not g15222 (n_5024, n10292);
  and g15223 (n10293, n_5023, n_5024);
  not g15224 (n_5025, n10293);
  and g15225 (n10294, \a[11] , n_5025);
  and g15226 (n10295, n_1071, n10293);
  not g15227 (n_5026, n10294);
  not g15228 (n_5027, n10295);
  and g15229 (n10296, n_5026, n_5027);
  not g15230 (n_5028, n10296);
  and g15231 (n10297, n10285, n_5028);
  and g15232 (n10298, n_316, n7632);
  and g15233 (n10299, n_315, n7983);
  not g15234 (n_5029, n10298);
  not g15235 (n_5030, n10299);
  and g15236 (n10300, n_5029, n_5030);
  and g15237 (n10301, n7294, n_2588);
  not g15238 (n_5031, n10301);
  and g15239 (n10302, n10300, n_5031);
  not g15240 (n_5032, n10302);
  and g15241 (n10303, \a[11] , n_5032);
  not g15242 (n_5033, n10303);
  and g15243 (n10304, \a[11] , n_5033);
  and g15244 (n10305, n_5032, n_5033);
  not g15245 (n_5034, n10304);
  not g15246 (n_5035, n10305);
  and g15247 (n10306, n_5034, n_5035);
  and g15248 (n10307, n_316, n_2445);
  not g15249 (n_5036, n10307);
  and g15250 (n10308, \a[11] , n_5036);
  not g15251 (n_5037, n10306);
  and g15252 (n10309, n_5037, n10308);
  and g15253 (n10310, n_314, n7983);
  and g15254 (n10311, n_316, n7291);
  and g15255 (n10312, n_315, n7632);
  not g15256 (n_5038, n10311);
  not g15257 (n_5039, n10312);
  and g15258 (n10313, n_5038, n_5039);
  not g15259 (n_5040, n10310);
  and g15260 (n10314, n_5040, n10313);
  and g15261 (n10315, n_2446, n10314);
  and g15262 (n10316, n_2612, n10314);
  not g15263 (n_5041, n10315);
  not g15264 (n_5042, n10316);
  and g15265 (n10317, n_5041, n_5042);
  not g15266 (n_5043, n10317);
  and g15267 (n10318, \a[11] , n_5043);
  and g15268 (n10319, n_1071, n10317);
  not g15269 (n_5044, n10318);
  not g15270 (n_5045, n10319);
  and g15271 (n10320, n_5044, n_5045);
  not g15272 (n_5046, n10320);
  and g15273 (n10321, n10309, n_5046);
  and g15274 (n10322, n9712, n10321);
  not g15275 (n_5047, n10322);
  and g15276 (n10323, n10321, n_5047);
  and g15277 (n10324, n9712, n_5047);
  not g15278 (n_5048, n10323);
  not g15279 (n_5049, n10324);
  and g15280 (n10325, n_5048, n_5049);
  and g15281 (n10326, n_313, n7983);
  and g15282 (n10327, n_315, n7291);
  and g15283 (n10328, n_314, n7632);
  and g15289 (n10331, n6806, n7294);
  not g15292 (n_5054, n10332);
  and g15293 (n10333, \a[11] , n_5054);
  not g15294 (n_5055, n10333);
  and g15295 (n10334, \a[11] , n_5055);
  and g15296 (n10335, n_5054, n_5055);
  not g15297 (n_5056, n10334);
  not g15298 (n_5057, n10335);
  and g15299 (n10336, n_5056, n_5057);
  not g15300 (n_5058, n10325);
  not g15301 (n_5059, n10336);
  and g15302 (n10337, n_5058, n_5059);
  not g15303 (n_5060, n10337);
  and g15304 (n10338, n_5047, n_5060);
  not g15305 (n_5061, n10285);
  and g15306 (n10339, n_5061, n10296);
  not g15307 (n_5062, n10297);
  not g15308 (n_5063, n10339);
  and g15309 (n10340, n_5062, n_5063);
  not g15310 (n_5064, n10338);
  and g15311 (n10341, n_5064, n10340);
  not g15312 (n_5065, n10341);
  and g15313 (n10342, n_5062, n_5065);
  not g15314 (n_5066, n10283);
  not g15315 (n_5067, n10342);
  and g15316 (n10343, n_5066, n_5067);
  not g15317 (n_5068, n10343);
  and g15318 (n10344, n_5015, n_5068);
  and g15319 (n10345, n10254, n10265);
  not g15320 (n_5069, n10266);
  not g15321 (n_5070, n10345);
  and g15322 (n10346, n_5069, n_5070);
  not g15323 (n_5071, n10344);
  and g15324 (n10347, n_5071, n10346);
  not g15325 (n_5072, n10347);
  and g15326 (n10348, n_5069, n_5072);
  not g15327 (n_5073, n10251);
  not g15328 (n_5074, n10348);
  and g15329 (n10349, n_5073, n_5074);
  not g15330 (n_5075, n10349);
  and g15331 (n10350, n_4988, n_5075);
  not g15332 (n_5076, n10234);
  and g15333 (n10351, n10222, n_5076);
  and g15334 (n10352, n_4976, n_5076);
  not g15335 (n_5077, n10351);
  not g15336 (n_5078, n10352);
  and g15337 (n10353, n_5077, n_5078);
  not g15338 (n_5079, n10350);
  not g15339 (n_5080, n10353);
  and g15340 (n10354, n_5079, n_5080);
  not g15341 (n_5081, n10354);
  and g15342 (n10355, n_5076, n_5081);
  not g15343 (n_5082, n10220);
  and g15344 (n10356, n10208, n_5082);
  and g15345 (n10357, n_4966, n_5082);
  not g15346 (n_5083, n10356);
  not g15347 (n_5084, n10357);
  and g15348 (n10358, n_5083, n_5084);
  not g15349 (n_5085, n10355);
  not g15350 (n_5086, n10358);
  and g15351 (n10359, n_5085, n_5086);
  not g15352 (n_5087, n10359);
  and g15353 (n10360, n_5082, n_5087);
  not g15354 (n_5088, n10194);
  and g15355 (n10361, n_5088, n10205);
  not g15356 (n_5089, n10206);
  not g15357 (n_5090, n10361);
  and g15358 (n10362, n_5089, n_5090);
  not g15359 (n_5091, n10360);
  and g15360 (n10363, n_5091, n10362);
  not g15361 (n_5092, n10363);
  and g15362 (n10364, n_5089, n_5092);
  not g15363 (n_5093, n10192);
  not g15364 (n_5094, n10364);
  and g15365 (n10365, n_5093, n_5094);
  not g15366 (n_5095, n10365);
  and g15367 (n10366, n_4943, n_5095);
  not g15368 (n_5096, n10174);
  not g15369 (n_5097, n10366);
  and g15370 (n10367, n_5096, n_5097);
  not g15371 (n_5098, n10367);
  and g15372 (n10368, n_4928, n_5098);
  not g15373 (n_5099, n10156);
  not g15374 (n_5100, n10368);
  and g15375 (n10369, n_5099, n_5100);
  not g15376 (n_5101, n10369);
  and g15377 (n10370, n_4913, n_5101);
  not g15378 (n_5102, n10139);
  and g15379 (n10371, n10127, n_5102);
  and g15380 (n10372, n_4901, n_5102);
  not g15381 (n_5103, n10371);
  not g15382 (n_5104, n10372);
  and g15383 (n10373, n_5103, n_5104);
  not g15384 (n_5105, n10370);
  not g15385 (n_5106, n10373);
  and g15386 (n10374, n_5105, n_5106);
  not g15387 (n_5107, n10374);
  and g15388 (n10375, n_5102, n_5107);
  not g15389 (n_5108, n10125);
  and g15390 (n10376, n10113, n_5108);
  and g15391 (n10377, n_4891, n_5108);
  not g15392 (n_5109, n10376);
  not g15393 (n_5110, n10377);
  and g15394 (n10378, n_5109, n_5110);
  not g15395 (n_5111, n10375);
  not g15396 (n_5112, n10378);
  and g15397 (n10379, n_5111, n_5112);
  not g15398 (n_5113, n10379);
  and g15399 (n10380, n_5108, n_5113);
  not g15400 (n_5114, n10099);
  and g15401 (n10381, n_5114, n10110);
  not g15402 (n_5115, n10111);
  not g15403 (n_5116, n10381);
  and g15404 (n10382, n_5115, n_5116);
  not g15405 (n_5117, n10380);
  and g15406 (n10383, n_5117, n10382);
  not g15407 (n_5118, n10383);
  and g15408 (n10384, n_5115, n_5118);
  not g15409 (n_5119, n10097);
  not g15410 (n_5120, n10384);
  and g15411 (n10385, n_5119, n_5120);
  not g15412 (n_5121, n10385);
  and g15413 (n10386, n_4869, n_5121);
  not g15414 (n_5122, n10079);
  not g15415 (n_5123, n10386);
  and g15416 (n10387, n_5122, n_5123);
  not g15417 (n_5124, n10387);
  and g15418 (n10388, n_4854, n_5124);
  not g15419 (n_5125, n10061);
  not g15420 (n_5126, n10388);
  and g15421 (n10389, n_5125, n_5126);
  not g15422 (n_5127, n10389);
  and g15423 (n10390, n_4839, n_5127);
  not g15424 (n_5128, n10044);
  and g15425 (n10391, n10032, n_5128);
  and g15426 (n10392, n_4827, n_5128);
  not g15427 (n_5129, n10391);
  not g15428 (n_5130, n10392);
  and g15429 (n10393, n_5129, n_5130);
  not g15430 (n_5131, n10390);
  not g15431 (n_5132, n10393);
  and g15432 (n10394, n_5131, n_5132);
  not g15433 (n_5133, n10394);
  and g15434 (n10395, n_5128, n_5133);
  not g15435 (n_5134, n10018);
  and g15436 (n10396, n_5134, n10029);
  not g15437 (n_5135, n10030);
  not g15438 (n_5136, n10396);
  and g15439 (n10397, n_5135, n_5136);
  not g15440 (n_5137, n10395);
  and g15441 (n10398, n_5137, n10397);
  not g15442 (n_5138, n10398);
  and g15443 (n10399, n_5135, n_5138);
  not g15444 (n_5139, n10016);
  not g15445 (n_5140, n10399);
  and g15446 (n10400, n_5139, n_5140);
  not g15447 (n_5141, n10400);
  and g15448 (n10401, n_4805, n_5141);
  not g15449 (n_5142, n9998);
  not g15450 (n_5143, n10401);
  and g15451 (n10402, n_5142, n_5143);
  not g15452 (n_5144, n10402);
  and g15453 (n10403, n_4790, n_5144);
  not g15454 (n_5145, n9980);
  not g15455 (n_5146, n10403);
  and g15456 (n10404, n_5145, n_5146);
  not g15457 (n_5147, n10404);
  and g15458 (n10405, n_4775, n_5147);
  not g15459 (n_5148, n9962);
  not g15460 (n_5149, n10405);
  and g15461 (n10406, n_5148, n_5149);
  not g15462 (n_5150, n10406);
  and g15463 (n10407, n_4760, n_5150);
  not g15464 (n_5151, n9944);
  not g15465 (n_5152, n10407);
  and g15466 (n10408, n_5151, n_5152);
  not g15467 (n_5153, n10408);
  and g15468 (n10409, n_4745, n_5153);
  not g15469 (n_5154, n9926);
  not g15470 (n_5155, n10409);
  and g15471 (n10410, n_5154, n_5155);
  not g15472 (n_5156, n10410);
  and g15473 (n10411, n_4730, n_5156);
  not g15474 (n_5157, n9908);
  not g15475 (n_5158, n10411);
  and g15476 (n10412, n_5157, n_5158);
  not g15477 (n_5159, n10412);
  and g15478 (n10413, n_4715, n_5159);
  not g15479 (n_5160, n9844);
  and g15480 (n10414, n9842, n_5160);
  not g15481 (n_5161, n10414);
  and g15482 (n10415, n_4665, n_5161);
  not g15483 (n_5162, n10413);
  and g15484 (n10416, n_5162, n10415);
  and g15485 (n10417, n_565, n9331);
  and g15486 (n10418, n_480, n8418);
  and g15487 (n10419, n_535, n8860);
  and g15493 (n10422, n4558, n8421);
  not g15496 (n_5167, n10423);
  and g15497 (n10424, \a[8] , n_5167);
  not g15498 (n_5168, n10424);
  and g15499 (n10425, n_5167, n_5168);
  and g15500 (n10426, \a[8] , n_5168);
  not g15501 (n_5169, n10425);
  not g15502 (n_5170, n10426);
  and g15503 (n10427, n_5169, n_5170);
  not g15504 (n_5171, n10416);
  and g15505 (n10428, n_5162, n_5171);
  and g15506 (n10429, n10415, n_5171);
  not g15507 (n_5172, n10428);
  not g15508 (n_5173, n10429);
  and g15509 (n10430, n_5172, n_5173);
  not g15510 (n_5174, n10427);
  not g15511 (n_5175, n10430);
  and g15512 (n10431, n_5174, n_5175);
  not g15513 (n_5176, n10431);
  and g15514 (n10432, n_5171, n_5176);
  and g15515 (n10433, n_560, n9867);
  not g15516 (n_5177, n9865);
  and g15517 (n10434, n70, n_5177);
  and g15518 (n10435, n_712, n10434);
  not g15519 (n_5178, n10433);
  not g15520 (n_5179, n10435);
  and g15521 (n10436, n_5178, n_5179);
  and g15522 (n10437, n_4684, n10436);
  and g15523 (n10438, n_2152, n10436);
  not g15524 (n_5180, n10437);
  not g15525 (n_5181, n10438);
  and g15526 (n10439, n_5180, n_5181);
  not g15527 (n_5182, n10439);
  and g15528 (n10440, \a[5] , n_5182);
  and g15529 (n10441, n_3, n10439);
  not g15530 (n_5183, n10440);
  not g15531 (n_5184, n10441);
  and g15532 (n10442, n_5183, n_5184);
  not g15533 (n_5185, n10432);
  not g15534 (n_5186, n10442);
  and g15535 (n10443, n_5185, n_5186);
  and g15536 (n10444, n9849, n_4679);
  and g15537 (n10445, n_4678, n_4679);
  not g15538 (n_5187, n10444);
  not g15539 (n_5188, n10445);
  and g15540 (n10446, n_5187, n_5188);
  and g15541 (n10447, n10432, n10442);
  not g15542 (n_5189, n10443);
  not g15543 (n_5190, n10447);
  and g15544 (n10448, n_5189, n_5190);
  not g15545 (n_5191, n10446);
  and g15546 (n10449, n_5191, n10448);
  not g15547 (n_5192, n10449);
  and g15548 (n10450, n_5189, n_5192);
  not g15549 (n_5193, n9890);
  not g15550 (n_5194, n10450);
  and g15551 (n10451, n_5193, n_5194);
  and g15552 (n10452, n9890, n10450);
  not g15553 (n_5195, n10451);
  not g15554 (n_5196, n10452);
  and g15555 (n10453, n_5195, n_5196);
  and g15556 (n10454, n9908, n10411);
  not g15557 (n_5197, n10454);
  and g15558 (n10455, n_5159, n_5197);
  and g15559 (n10456, n_535, n9331);
  and g15560 (n10457, n_485, n8418);
  and g15561 (n10458, n_480, n8860);
  not g15562 (n_5198, n10457);
  not g15563 (n_5199, n10458);
  and g15564 (n10459, n_5198, n_5199);
  not g15565 (n_5200, n10456);
  and g15566 (n10460, n_5200, n10459);
  and g15567 (n10461, n_3428, n10460);
  and g15568 (n10462, n_545, n10460);
  not g15569 (n_5201, n10461);
  not g15570 (n_5202, n10462);
  and g15571 (n10463, n_5201, n_5202);
  not g15572 (n_5203, n10463);
  and g15573 (n10464, \a[8] , n_5203);
  and g15574 (n10465, n_1106, n10463);
  not g15575 (n_5204, n10464);
  not g15576 (n_5205, n10465);
  and g15577 (n10466, n_5204, n_5205);
  not g15578 (n_5206, n10466);
  and g15579 (n10467, n10455, n_5206);
  and g15580 (n10468, n9926, n10409);
  not g15581 (n_5207, n10468);
  and g15582 (n10469, n_5156, n_5207);
  and g15583 (n10470, n_480, n9331);
  and g15584 (n10471, n_484, n8418);
  and g15585 (n10472, n_485, n8860);
  not g15586 (n_5208, n10471);
  not g15587 (n_5209, n10472);
  and g15588 (n10473, n_5208, n_5209);
  not g15589 (n_5210, n10470);
  and g15590 (n10474, n_5210, n10473);
  and g15591 (n10475, n_3428, n10474);
  and g15592 (n10476, n_504, n10474);
  not g15593 (n_5211, n10475);
  not g15594 (n_5212, n10476);
  and g15595 (n10477, n_5211, n_5212);
  not g15596 (n_5213, n10477);
  and g15597 (n10478, \a[8] , n_5213);
  and g15598 (n10479, n_1106, n10477);
  not g15599 (n_5214, n10478);
  not g15600 (n_5215, n10479);
  and g15601 (n10480, n_5214, n_5215);
  not g15602 (n_5216, n10480);
  and g15603 (n10481, n10469, n_5216);
  and g15604 (n10482, n9944, n10407);
  not g15605 (n_5217, n10482);
  and g15606 (n10483, n_5153, n_5217);
  and g15607 (n10484, n_485, n9331);
  and g15608 (n10485, n_415, n8418);
  and g15609 (n10486, n_484, n8860);
  not g15610 (n_5218, n10485);
  not g15611 (n_5219, n10486);
  and g15612 (n10487, n_5218, n_5219);
  not g15613 (n_5220, n10484);
  and g15614 (n10488, n_5220, n10487);
  and g15615 (n10489, n_3428, n10488);
  and g15616 (n10490, n_914, n10488);
  not g15617 (n_5221, n10489);
  not g15618 (n_5222, n10490);
  and g15619 (n10491, n_5221, n_5222);
  not g15620 (n_5223, n10491);
  and g15621 (n10492, \a[8] , n_5223);
  and g15622 (n10493, n_1106, n10491);
  not g15623 (n_5224, n10492);
  not g15624 (n_5225, n10493);
  and g15625 (n10494, n_5224, n_5225);
  not g15626 (n_5226, n10494);
  and g15627 (n10495, n10483, n_5226);
  and g15628 (n10496, n9962, n10405);
  not g15629 (n_5227, n10496);
  and g15630 (n10497, n_5150, n_5227);
  and g15631 (n10498, n_484, n9331);
  and g15632 (n10499, n_236, n8418);
  and g15633 (n10500, n_415, n8860);
  not g15634 (n_5228, n10499);
  not g15635 (n_5229, n10500);
  and g15636 (n10501, n_5228, n_5229);
  not g15637 (n_5230, n10498);
  and g15638 (n10502, n_5230, n10501);
  and g15639 (n10503, n_3428, n10502);
  and g15640 (n10504, n_773, n10502);
  not g15641 (n_5231, n10503);
  not g15642 (n_5232, n10504);
  and g15643 (n10505, n_5231, n_5232);
  not g15644 (n_5233, n10505);
  and g15645 (n10506, \a[8] , n_5233);
  and g15646 (n10507, n_1106, n10505);
  not g15647 (n_5234, n10506);
  not g15648 (n_5235, n10507);
  and g15649 (n10508, n_5234, n_5235);
  not g15650 (n_5236, n10508);
  and g15651 (n10509, n10497, n_5236);
  and g15652 (n10510, n9980, n10403);
  not g15653 (n_5237, n10510);
  and g15654 (n10511, n_5147, n_5237);
  and g15655 (n10512, n_415, n9331);
  and g15656 (n10513, n_237, n8418);
  and g15657 (n10514, n_236, n8860);
  not g15658 (n_5238, n10513);
  not g15659 (n_5239, n10514);
  and g15660 (n10515, n_5238, n_5239);
  not g15661 (n_5240, n10512);
  and g15662 (n10516, n_5240, n10515);
  and g15663 (n10517, n_3428, n10516);
  and g15664 (n10518, n_680, n10516);
  not g15665 (n_5241, n10517);
  not g15666 (n_5242, n10518);
  and g15667 (n10519, n_5241, n_5242);
  not g15668 (n_5243, n10519);
  and g15669 (n10520, \a[8] , n_5243);
  and g15670 (n10521, n_1106, n10519);
  not g15671 (n_5244, n10520);
  not g15672 (n_5245, n10521);
  and g15673 (n10522, n_5244, n_5245);
  not g15674 (n_5246, n10522);
  and g15675 (n10523, n10511, n_5246);
  and g15676 (n10524, n9998, n10401);
  not g15677 (n_5247, n10524);
  and g15678 (n10525, n_5144, n_5247);
  and g15679 (n10526, n_236, n9331);
  and g15680 (n10527, n_260, n8418);
  and g15681 (n10528, n_237, n8860);
  not g15682 (n_5248, n10527);
  not g15683 (n_5249, n10528);
  and g15684 (n10529, n_5248, n_5249);
  not g15685 (n_5250, n10526);
  and g15686 (n10530, n_5250, n10529);
  and g15687 (n10531, n_3428, n10530);
  and g15688 (n10532, n_1208, n10530);
  not g15689 (n_5251, n10531);
  not g15690 (n_5252, n10532);
  and g15691 (n10533, n_5251, n_5252);
  not g15692 (n_5253, n10533);
  and g15693 (n10534, \a[8] , n_5253);
  and g15694 (n10535, n_1106, n10533);
  not g15695 (n_5254, n10534);
  not g15696 (n_5255, n10535);
  and g15697 (n10536, n_5254, n_5255);
  not g15698 (n_5256, n10536);
  and g15699 (n10537, n10525, n_5256);
  and g15700 (n10538, n10016, n10399);
  not g15701 (n_5257, n10538);
  and g15702 (n10539, n_5141, n_5257);
  and g15703 (n10540, n_237, n9331);
  and g15704 (n10541, n_275, n8418);
  and g15705 (n10542, n_260, n8860);
  not g15706 (n_5258, n10541);
  not g15707 (n_5259, n10542);
  and g15708 (n10543, n_5258, n_5259);
  not g15709 (n_5260, n10540);
  and g15710 (n10544, n_5260, n10543);
  and g15711 (n10545, n_3428, n10544);
  and g15712 (n10546, n_4259, n10544);
  not g15713 (n_5261, n10545);
  not g15714 (n_5262, n10546);
  and g15715 (n10547, n_5261, n_5262);
  not g15716 (n_5263, n10547);
  and g15717 (n10548, \a[8] , n_5263);
  and g15718 (n10549, n_1106, n10547);
  not g15719 (n_5264, n10548);
  not g15720 (n_5265, n10549);
  and g15721 (n10550, n_5264, n_5265);
  not g15722 (n_5266, n10550);
  and g15723 (n10551, n10539, n_5266);
  and g15724 (n10552, n_260, n9331);
  and g15725 (n10553, n_281, n8418);
  and g15726 (n10554, n_275, n8860);
  and g15732 (n10557, n4179, n8421);
  not g15735 (n_5271, n10558);
  and g15736 (n10559, \a[8] , n_5271);
  not g15737 (n_5272, n10559);
  and g15738 (n10560, n_5271, n_5272);
  and g15739 (n10561, \a[8] , n_5272);
  not g15740 (n_5273, n10560);
  not g15741 (n_5274, n10561);
  and g15742 (n10562, n_5273, n_5274);
  not g15743 (n_5275, n10397);
  and g15744 (n10563, n10395, n_5275);
  not g15745 (n_5276, n10563);
  and g15746 (n10564, n_5138, n_5276);
  not g15747 (n_5277, n10562);
  and g15748 (n10565, n_5277, n10564);
  not g15749 (n_5278, n10565);
  and g15750 (n10566, n_5277, n_5278);
  and g15751 (n10567, n10564, n_5278);
  not g15752 (n_5279, n10566);
  not g15753 (n_5280, n10567);
  and g15754 (n10568, n_5279, n_5280);
  and g15755 (n10569, n_275, n9331);
  and g15756 (n10570, n_286, n8418);
  and g15757 (n10571, n_281, n8860);
  and g15763 (n10574, n4204, n8421);
  not g15766 (n_5285, n10575);
  and g15767 (n10576, \a[8] , n_5285);
  not g15768 (n_5286, n10576);
  and g15769 (n10577, n_5285, n_5286);
  and g15770 (n10578, \a[8] , n_5286);
  not g15771 (n_5287, n10577);
  not g15772 (n_5288, n10578);
  and g15773 (n10579, n_5287, n_5288);
  and g15774 (n10580, n_5131, n_5133);
  and g15775 (n10581, n_5132, n_5133);
  not g15776 (n_5289, n10580);
  not g15777 (n_5290, n10581);
  and g15778 (n10582, n_5289, n_5290);
  not g15779 (n_5291, n10579);
  not g15780 (n_5292, n10582);
  and g15781 (n10583, n_5291, n_5292);
  not g15782 (n_5293, n10583);
  and g15783 (n10584, n_5291, n_5293);
  and g15784 (n10585, n_5292, n_5293);
  not g15785 (n_5294, n10584);
  not g15786 (n_5295, n10585);
  and g15787 (n10586, n_5294, n_5295);
  and g15788 (n10587, n10061, n10388);
  not g15789 (n_5296, n10587);
  and g15790 (n10588, n_5127, n_5296);
  and g15791 (n10589, n_281, n9331);
  and g15792 (n10590, n_293, n8418);
  and g15793 (n10591, n_286, n8860);
  not g15794 (n_5297, n10590);
  not g15795 (n_5298, n10591);
  and g15796 (n10592, n_5297, n_5298);
  not g15797 (n_5299, n10589);
  and g15798 (n10593, n_5299, n10592);
  and g15799 (n10594, n_3428, n10593);
  and g15800 (n10595, n_1228, n10593);
  not g15801 (n_5300, n10594);
  not g15802 (n_5301, n10595);
  and g15803 (n10596, n_5300, n_5301);
  not g15804 (n_5302, n10596);
  and g15805 (n10597, \a[8] , n_5302);
  and g15806 (n10598, n_1106, n10596);
  not g15807 (n_5303, n10597);
  not g15808 (n_5304, n10598);
  and g15809 (n10599, n_5303, n_5304);
  not g15810 (n_5305, n10599);
  and g15811 (n10600, n10588, n_5305);
  and g15812 (n10601, n10079, n10386);
  not g15813 (n_5306, n10601);
  and g15814 (n10602, n_5124, n_5306);
  and g15815 (n10603, n_286, n9331);
  and g15816 (n10604, n_295, n8418);
  and g15817 (n10605, n_293, n8860);
  not g15818 (n_5307, n10604);
  not g15819 (n_5308, n10605);
  and g15820 (n10606, n_5307, n_5308);
  not g15821 (n_5309, n10603);
  and g15822 (n10607, n_5309, n10606);
  and g15823 (n10608, n_3428, n10607);
  and g15824 (n10609, n_1134, n10607);
  not g15825 (n_5310, n10608);
  not g15826 (n_5311, n10609);
  and g15827 (n10610, n_5310, n_5311);
  not g15828 (n_5312, n10610);
  and g15829 (n10611, \a[8] , n_5312);
  and g15830 (n10612, n_1106, n10610);
  not g15831 (n_5313, n10611);
  not g15832 (n_5314, n10612);
  and g15833 (n10613, n_5313, n_5314);
  not g15834 (n_5315, n10613);
  and g15835 (n10614, n10602, n_5315);
  and g15836 (n10615, n10097, n10384);
  not g15837 (n_5316, n10615);
  and g15838 (n10616, n_5121, n_5316);
  and g15839 (n10617, n_293, n9331);
  and g15840 (n10618, n_298, n8418);
  and g15841 (n10619, n_295, n8860);
  not g15842 (n_5317, n10618);
  not g15843 (n_5318, n10619);
  and g15844 (n10620, n_5317, n_5318);
  not g15845 (n_5319, n10617);
  and g15846 (n10621, n_5319, n10620);
  and g15847 (n10622, n_3428, n10621);
  and g15848 (n10623, n_1789, n10621);
  not g15849 (n_5320, n10622);
  not g15850 (n_5321, n10623);
  and g15851 (n10624, n_5320, n_5321);
  not g15852 (n_5322, n10624);
  and g15853 (n10625, \a[8] , n_5322);
  and g15854 (n10626, n_1106, n10624);
  not g15855 (n_5323, n10625);
  not g15856 (n_5324, n10626);
  and g15857 (n10627, n_5323, n_5324);
  not g15858 (n_5325, n10627);
  and g15859 (n10628, n10616, n_5325);
  and g15860 (n10629, n_295, n9331);
  and g15861 (n10630, n_299, n8418);
  and g15862 (n10631, n_298, n8860);
  and g15868 (n10634, n4848, n8421);
  not g15871 (n_5330, n10635);
  and g15872 (n10636, \a[8] , n_5330);
  not g15873 (n_5331, n10636);
  and g15874 (n10637, n_5330, n_5331);
  and g15875 (n10638, \a[8] , n_5331);
  not g15876 (n_5332, n10637);
  not g15877 (n_5333, n10638);
  and g15878 (n10639, n_5332, n_5333);
  not g15879 (n_5334, n10382);
  and g15880 (n10640, n10380, n_5334);
  not g15881 (n_5335, n10640);
  and g15882 (n10641, n_5118, n_5335);
  not g15883 (n_5336, n10639);
  and g15884 (n10642, n_5336, n10641);
  not g15885 (n_5337, n10642);
  and g15886 (n10643, n_5336, n_5337);
  and g15887 (n10644, n10641, n_5337);
  not g15888 (n_5338, n10643);
  not g15889 (n_5339, n10644);
  and g15890 (n10645, n_5338, n_5339);
  and g15891 (n10646, n_298, n9331);
  and g15892 (n10647, n_300, n8418);
  and g15893 (n10648, n_299, n8860);
  and g15899 (n10651, n5114, n8421);
  not g15902 (n_5344, n10652);
  and g15903 (n10653, \a[8] , n_5344);
  not g15904 (n_5345, n10653);
  and g15905 (n10654, n_5344, n_5345);
  and g15906 (n10655, \a[8] , n_5345);
  not g15907 (n_5346, n10654);
  not g15908 (n_5347, n10655);
  and g15909 (n10656, n_5346, n_5347);
  and g15910 (n10657, n_5111, n_5113);
  and g15911 (n10658, n_5112, n_5113);
  not g15912 (n_5348, n10657);
  not g15913 (n_5349, n10658);
  and g15914 (n10659, n_5348, n_5349);
  not g15915 (n_5350, n10656);
  not g15916 (n_5351, n10659);
  and g15917 (n10660, n_5350, n_5351);
  not g15918 (n_5352, n10660);
  and g15919 (n10661, n_5350, n_5352);
  and g15920 (n10662, n_5351, n_5352);
  not g15921 (n_5353, n10661);
  not g15922 (n_5354, n10662);
  and g15923 (n10663, n_5353, n_5354);
  and g15924 (n10664, n_299, n9331);
  and g15925 (n10665, n_301, n8418);
  and g15926 (n10666, n_300, n8860);
  and g15932 (n10669, n5139, n8421);
  not g15935 (n_5359, n10670);
  and g15936 (n10671, \a[8] , n_5359);
  not g15937 (n_5360, n10671);
  and g15938 (n10672, n_5359, n_5360);
  and g15939 (n10673, \a[8] , n_5360);
  not g15940 (n_5361, n10672);
  not g15941 (n_5362, n10673);
  and g15942 (n10674, n_5361, n_5362);
  and g15943 (n10675, n_5105, n_5107);
  and g15944 (n10676, n_5106, n_5107);
  not g15945 (n_5363, n10675);
  not g15946 (n_5364, n10676);
  and g15947 (n10677, n_5363, n_5364);
  not g15948 (n_5365, n10674);
  not g15949 (n_5366, n10677);
  and g15950 (n10678, n_5365, n_5366);
  not g15951 (n_5367, n10678);
  and g15952 (n10679, n_5365, n_5367);
  and g15953 (n10680, n_5366, n_5367);
  not g15954 (n_5368, n10679);
  not g15955 (n_5369, n10680);
  and g15956 (n10681, n_5368, n_5369);
  and g15957 (n10682, n10156, n10368);
  not g15958 (n_5370, n10682);
  and g15959 (n10683, n_5101, n_5370);
  and g15960 (n10684, n_300, n9331);
  and g15961 (n10685, n_302, n8418);
  and g15962 (n10686, n_301, n8860);
  not g15963 (n_5371, n10685);
  not g15964 (n_5372, n10686);
  and g15965 (n10687, n_5371, n_5372);
  not g15966 (n_5373, n10684);
  and g15967 (n10688, n_5373, n10687);
  and g15968 (n10689, n_3428, n10688);
  and g15969 (n10690, n_1801, n10688);
  not g15970 (n_5374, n10689);
  not g15971 (n_5375, n10690);
  and g15972 (n10691, n_5374, n_5375);
  not g15973 (n_5376, n10691);
  and g15974 (n10692, \a[8] , n_5376);
  and g15975 (n10693, n_1106, n10691);
  not g15976 (n_5377, n10692);
  not g15977 (n_5378, n10693);
  and g15978 (n10694, n_5377, n_5378);
  not g15979 (n_5379, n10694);
  and g15980 (n10695, n10683, n_5379);
  and g15981 (n10696, n10174, n10366);
  not g15982 (n_5380, n10696);
  and g15983 (n10697, n_5098, n_5380);
  and g15984 (n10698, n_301, n9331);
  and g15985 (n10699, n_303, n8418);
  and g15986 (n10700, n_302, n8860);
  not g15987 (n_5381, n10699);
  not g15988 (n_5382, n10700);
  and g15989 (n10701, n_5381, n_5382);
  not g15990 (n_5383, n10698);
  and g15991 (n10702, n_5383, n10701);
  and g15992 (n10703, n_3428, n10702);
  and g15993 (n10704, n_1672, n10702);
  not g15994 (n_5384, n10703);
  not g15995 (n_5385, n10704);
  and g15996 (n10705, n_5384, n_5385);
  not g15997 (n_5386, n10705);
  and g15998 (n10706, \a[8] , n_5386);
  and g15999 (n10707, n_1106, n10705);
  not g16000 (n_5387, n10706);
  not g16001 (n_5388, n10707);
  and g16002 (n10708, n_5387, n_5388);
  not g16003 (n_5389, n10708);
  and g16004 (n10709, n10697, n_5389);
  and g16005 (n10710, n10192, n10364);
  not g16006 (n_5390, n10710);
  and g16007 (n10711, n_5095, n_5390);
  and g16008 (n10712, n_302, n9331);
  and g16009 (n10713, n_304, n8418);
  and g16010 (n10714, n_303, n8860);
  not g16011 (n_5391, n10713);
  not g16012 (n_5392, n10714);
  and g16013 (n10715, n_5391, n_5392);
  not g16014 (n_5393, n10712);
  and g16015 (n10716, n_5393, n10715);
  and g16016 (n10717, n_3428, n10716);
  and g16017 (n10718, n_3507, n10716);
  not g16018 (n_5394, n10717);
  not g16019 (n_5395, n10718);
  and g16020 (n10719, n_5394, n_5395);
  not g16021 (n_5396, n10719);
  and g16022 (n10720, \a[8] , n_5396);
  and g16023 (n10721, n_1106, n10719);
  not g16024 (n_5397, n10720);
  not g16025 (n_5398, n10721);
  and g16026 (n10722, n_5397, n_5398);
  not g16027 (n_5399, n10722);
  and g16028 (n10723, n10711, n_5399);
  and g16029 (n10724, n_303, n9331);
  and g16030 (n10725, n_305, n8418);
  and g16031 (n10726, n_304, n8860);
  and g16037 (n10729, n6007, n8421);
  not g16040 (n_5404, n10730);
  and g16041 (n10731, \a[8] , n_5404);
  not g16042 (n_5405, n10731);
  and g16043 (n10732, n_5404, n_5405);
  and g16044 (n10733, \a[8] , n_5405);
  not g16045 (n_5406, n10732);
  not g16046 (n_5407, n10733);
  and g16047 (n10734, n_5406, n_5407);
  not g16048 (n_5408, n10362);
  and g16049 (n10735, n10360, n_5408);
  not g16050 (n_5409, n10735);
  and g16051 (n10736, n_5092, n_5409);
  not g16052 (n_5410, n10734);
  and g16053 (n10737, n_5410, n10736);
  not g16054 (n_5411, n10737);
  and g16055 (n10738, n_5410, n_5411);
  and g16056 (n10739, n10736, n_5411);
  not g16057 (n_5412, n10738);
  not g16058 (n_5413, n10739);
  and g16059 (n10740, n_5412, n_5413);
  and g16060 (n10741, n_304, n9331);
  and g16061 (n10742, n_306, n8418);
  and g16062 (n10743, n_305, n8860);
  and g16068 (n10746, n5834, n8421);
  not g16071 (n_5418, n10747);
  and g16072 (n10748, \a[8] , n_5418);
  not g16073 (n_5419, n10748);
  and g16074 (n10749, n_5418, n_5419);
  and g16075 (n10750, \a[8] , n_5419);
  not g16076 (n_5420, n10749);
  not g16077 (n_5421, n10750);
  and g16078 (n10751, n_5420, n_5421);
  and g16079 (n10752, n_5085, n_5087);
  and g16080 (n10753, n_5086, n_5087);
  not g16081 (n_5422, n10752);
  not g16082 (n_5423, n10753);
  and g16083 (n10754, n_5422, n_5423);
  not g16084 (n_5424, n10751);
  not g16085 (n_5425, n10754);
  and g16086 (n10755, n_5424, n_5425);
  not g16087 (n_5426, n10755);
  and g16088 (n10756, n_5424, n_5426);
  and g16089 (n10757, n_5425, n_5426);
  not g16090 (n_5427, n10756);
  not g16091 (n_5428, n10757);
  and g16092 (n10758, n_5427, n_5428);
  and g16093 (n10759, n_305, n9331);
  and g16094 (n10760, n_307, n8418);
  and g16095 (n10761, n_306, n8860);
  and g16101 (n10764, n6143, n8421);
  not g16104 (n_5433, n10765);
  and g16105 (n10766, \a[8] , n_5433);
  not g16106 (n_5434, n10766);
  and g16107 (n10767, n_5433, n_5434);
  and g16108 (n10768, \a[8] , n_5434);
  not g16109 (n_5435, n10767);
  not g16110 (n_5436, n10768);
  and g16111 (n10769, n_5435, n_5436);
  and g16112 (n10770, n_5079, n_5081);
  and g16113 (n10771, n_5080, n_5081);
  not g16114 (n_5437, n10770);
  not g16115 (n_5438, n10771);
  and g16116 (n10772, n_5437, n_5438);
  not g16117 (n_5439, n10769);
  not g16118 (n_5440, n10772);
  and g16119 (n10773, n_5439, n_5440);
  not g16120 (n_5441, n10773);
  and g16121 (n10774, n_5439, n_5441);
  and g16122 (n10775, n_5440, n_5441);
  not g16123 (n_5442, n10774);
  not g16124 (n_5443, n10775);
  and g16125 (n10776, n_5442, n_5443);
  and g16126 (n10777, n10251, n10348);
  not g16127 (n_5444, n10777);
  and g16128 (n10778, n_5075, n_5444);
  and g16129 (n10779, n_306, n9331);
  and g16130 (n10780, n_308, n8418);
  and g16131 (n10781, n_307, n8860);
  not g16132 (n_5445, n10780);
  not g16133 (n_5446, n10781);
  and g16134 (n10782, n_5445, n_5446);
  not g16135 (n_5447, n10779);
  and g16136 (n10783, n_5447, n10782);
  and g16137 (n10784, n_3428, n10783);
  and g16138 (n10785, n_2498, n10783);
  not g16139 (n_5448, n10784);
  not g16140 (n_5449, n10785);
  and g16141 (n10786, n_5448, n_5449);
  not g16142 (n_5450, n10786);
  and g16143 (n10787, \a[8] , n_5450);
  and g16144 (n10788, n_1106, n10786);
  not g16145 (n_5451, n10787);
  not g16146 (n_5452, n10788);
  and g16147 (n10789, n_5451, n_5452);
  not g16148 (n_5453, n10789);
  and g16149 (n10790, n10778, n_5453);
  not g16150 (n_5454, n10346);
  and g16151 (n10791, n10344, n_5454);
  not g16152 (n_5455, n10791);
  and g16153 (n10792, n_5072, n_5455);
  and g16154 (n10793, n_307, n9331);
  and g16155 (n10794, n_309, n8418);
  and g16156 (n10795, n_308, n8860);
  not g16157 (n_5456, n10794);
  not g16158 (n_5457, n10795);
  and g16159 (n10796, n_5456, n_5457);
  not g16160 (n_5458, n10793);
  and g16161 (n10797, n_5458, n10796);
  and g16162 (n10798, n_3428, n10797);
  and g16163 (n10799, n_2511, n10797);
  not g16164 (n_5459, n10798);
  not g16165 (n_5460, n10799);
  and g16166 (n10800, n_5459, n_5460);
  not g16167 (n_5461, n10800);
  and g16168 (n10801, \a[8] , n_5461);
  and g16169 (n10802, n_1106, n10800);
  not g16170 (n_5462, n10801);
  not g16171 (n_5463, n10802);
  and g16172 (n10803, n_5462, n_5463);
  not g16173 (n_5464, n10803);
  and g16174 (n10804, n10792, n_5464);
  and g16175 (n10805, n10283, n10342);
  not g16176 (n_5465, n10805);
  and g16177 (n10806, n_5068, n_5465);
  and g16178 (n10807, n_308, n9331);
  and g16179 (n10808, n_310, n8418);
  and g16180 (n10809, n_309, n8860);
  not g16181 (n_5466, n10808);
  not g16182 (n_5467, n10809);
  and g16183 (n10810, n_5466, n_5467);
  not g16184 (n_5468, n10807);
  and g16185 (n10811, n_5468, n10810);
  and g16186 (n10812, n_3428, n10811);
  and g16187 (n10813, n_2839, n10811);
  not g16188 (n_5469, n10812);
  not g16189 (n_5470, n10813);
  and g16190 (n10814, n_5469, n_5470);
  not g16191 (n_5471, n10814);
  and g16192 (n10815, \a[8] , n_5471);
  and g16193 (n10816, n_1106, n10814);
  not g16194 (n_5472, n10815);
  not g16195 (n_5473, n10816);
  and g16196 (n10817, n_5472, n_5473);
  not g16197 (n_5474, n10817);
  and g16198 (n10818, n10806, n_5474);
  and g16199 (n10819, n_309, n9331);
  and g16200 (n10820, n_311, n8418);
  and g16201 (n10821, n_310, n8860);
  and g16207 (n10824, n6541, n8421);
  not g16210 (n_5479, n10825);
  and g16211 (n10826, \a[8] , n_5479);
  not g16212 (n_5480, n10826);
  and g16213 (n10827, n_5479, n_5480);
  and g16214 (n10828, \a[8] , n_5480);
  not g16215 (n_5481, n10827);
  not g16216 (n_5482, n10828);
  and g16217 (n10829, n_5481, n_5482);
  not g16218 (n_5483, n10340);
  and g16219 (n10830, n10338, n_5483);
  not g16220 (n_5484, n10830);
  and g16221 (n10831, n_5065, n_5484);
  not g16222 (n_5485, n10829);
  and g16223 (n10832, n_5485, n10831);
  not g16224 (n_5486, n10832);
  and g16225 (n10833, n_5485, n_5486);
  and g16226 (n10834, n10831, n_5486);
  not g16227 (n_5487, n10833);
  not g16228 (n_5488, n10834);
  and g16229 (n10835, n_5487, n_5488);
  and g16230 (n10836, n_5058, n_5060);
  and g16231 (n10837, n_5059, n_5060);
  not g16232 (n_5489, n10836);
  not g16233 (n_5490, n10837);
  and g16234 (n10838, n_5489, n_5490);
  and g16235 (n10839, n_310, n9331);
  and g16236 (n10840, n_312, n8418);
  and g16237 (n10841, n_311, n8860);
  not g16238 (n_5491, n10840);
  not g16239 (n_5492, n10841);
  and g16240 (n10842, n_5491, n_5492);
  not g16241 (n_5493, n10839);
  and g16242 (n10843, n_5493, n10842);
  and g16243 (n10844, n_3428, n10843);
  and g16244 (n10845, n_3239, n10843);
  not g16245 (n_5494, n10844);
  not g16246 (n_5495, n10845);
  and g16247 (n10846, n_5494, n_5495);
  not g16248 (n_5496, n10846);
  and g16249 (n10847, \a[8] , n_5496);
  and g16250 (n10848, n_1106, n10846);
  not g16251 (n_5497, n10847);
  not g16252 (n_5498, n10848);
  and g16253 (n10849, n_5497, n_5498);
  not g16254 (n_5499, n10838);
  not g16255 (n_5500, n10849);
  and g16256 (n10850, n_5499, n_5500);
  and g16257 (n10851, n_311, n9331);
  and g16258 (n10852, n_313, n8418);
  and g16259 (n10853, n_312, n8860);
  and g16265 (n10856, n6646, n8421);
  not g16268 (n_5505, n10857);
  and g16269 (n10858, \a[8] , n_5505);
  not g16270 (n_5506, n10858);
  and g16271 (n10859, n_5505, n_5506);
  and g16272 (n10860, \a[8] , n_5506);
  not g16273 (n_5507, n10859);
  not g16274 (n_5508, n10860);
  and g16275 (n10861, n_5507, n_5508);
  not g16276 (n_5509, n10309);
  and g16277 (n10862, n_5509, n10320);
  not g16278 (n_5510, n10321);
  not g16279 (n_5511, n10862);
  and g16280 (n10863, n_5510, n_5511);
  not g16281 (n_5512, n10861);
  and g16282 (n10864, n_5512, n10863);
  not g16283 (n_5513, n10864);
  and g16284 (n10865, n_5512, n_5513);
  and g16285 (n10866, n10863, n_5513);
  not g16286 (n_5514, n10865);
  not g16287 (n_5515, n10866);
  and g16288 (n10867, n_5514, n_5515);
  not g16289 (n_5516, n10308);
  and g16290 (n10868, n10306, n_5516);
  not g16291 (n_5517, n10868);
  and g16292 (n10869, n_5509, n_5517);
  and g16293 (n10870, n_312, n9331);
  and g16294 (n10871, n_314, n8418);
  and g16295 (n10872, n_313, n8860);
  not g16296 (n_5518, n10871);
  not g16297 (n_5519, n10872);
  and g16298 (n10873, n_5518, n_5519);
  not g16299 (n_5520, n10870);
  and g16300 (n10874, n_5520, n10873);
  and g16301 (n10875, n_3428, n10874);
  and g16302 (n10876, n_2891, n10874);
  not g16303 (n_5521, n10875);
  not g16304 (n_5522, n10876);
  and g16305 (n10877, n_5521, n_5522);
  not g16306 (n_5523, n10877);
  and g16307 (n10878, \a[8] , n_5523);
  and g16308 (n10879, n_1106, n10877);
  not g16309 (n_5524, n10878);
  not g16310 (n_5525, n10879);
  and g16311 (n10880, n_5524, n_5525);
  not g16312 (n_5526, n10880);
  and g16313 (n10881, n10869, n_5526);
  and g16314 (n10882, n_316, n8860);
  and g16315 (n10883, n_315, n9331);
  not g16316 (n_5527, n10882);
  not g16317 (n_5528, n10883);
  and g16318 (n10884, n_5527, n_5528);
  and g16319 (n10885, n_2588, n8421);
  not g16320 (n_5529, n10885);
  and g16321 (n10886, n10884, n_5529);
  not g16322 (n_5530, n10886);
  and g16323 (n10887, \a[8] , n_5530);
  not g16324 (n_5531, n10887);
  and g16325 (n10888, \a[8] , n_5531);
  and g16326 (n10889, n_5530, n_5531);
  not g16327 (n_5532, n10888);
  not g16328 (n_5533, n10889);
  and g16329 (n10890, n_5532, n_5533);
  and g16330 (n10891, n_316, n_3427);
  not g16331 (n_5534, n10891);
  and g16332 (n10892, \a[8] , n_5534);
  not g16333 (n_5535, n10890);
  and g16334 (n10893, n_5535, n10892);
  and g16335 (n10894, n_314, n9331);
  and g16336 (n10895, n_316, n8418);
  and g16337 (n10896, n_315, n8860);
  not g16338 (n_5536, n10895);
  not g16339 (n_5537, n10896);
  and g16340 (n10897, n_5536, n_5537);
  not g16341 (n_5538, n10894);
  and g16342 (n10898, n_5538, n10897);
  and g16343 (n10899, n_3428, n10898);
  and g16344 (n10900, n_2612, n10898);
  not g16345 (n_5539, n10899);
  not g16346 (n_5540, n10900);
  and g16347 (n10901, n_5539, n_5540);
  not g16348 (n_5541, n10901);
  and g16349 (n10902, \a[8] , n_5541);
  and g16350 (n10903, n_1106, n10901);
  not g16351 (n_5542, n10902);
  not g16352 (n_5543, n10903);
  and g16353 (n10904, n_5542, n_5543);
  not g16354 (n_5544, n10904);
  and g16355 (n10905, n10893, n_5544);
  and g16356 (n10906, n10307, n10905);
  not g16357 (n_5545, n10906);
  and g16358 (n10907, n10905, n_5545);
  and g16359 (n10908, n10307, n_5545);
  not g16360 (n_5546, n10907);
  not g16361 (n_5547, n10908);
  and g16362 (n10909, n_5546, n_5547);
  and g16363 (n10910, n_313, n9331);
  and g16364 (n10911, n_315, n8418);
  and g16365 (n10912, n_314, n8860);
  and g16371 (n10915, n6806, n8421);
  not g16374 (n_5552, n10916);
  and g16375 (n10917, \a[8] , n_5552);
  not g16376 (n_5553, n10917);
  and g16377 (n10918, \a[8] , n_5553);
  and g16378 (n10919, n_5552, n_5553);
  not g16379 (n_5554, n10918);
  not g16380 (n_5555, n10919);
  and g16381 (n10920, n_5554, n_5555);
  not g16382 (n_5556, n10909);
  not g16383 (n_5557, n10920);
  and g16384 (n10921, n_5556, n_5557);
  not g16385 (n_5558, n10921);
  and g16386 (n10922, n_5545, n_5558);
  not g16387 (n_5559, n10869);
  and g16388 (n10923, n_5559, n10880);
  not g16389 (n_5560, n10881);
  not g16390 (n_5561, n10923);
  and g16391 (n10924, n_5560, n_5561);
  not g16392 (n_5562, n10922);
  and g16393 (n10925, n_5562, n10924);
  not g16394 (n_5563, n10925);
  and g16395 (n10926, n_5560, n_5563);
  not g16396 (n_5564, n10867);
  not g16397 (n_5565, n10926);
  and g16398 (n10927, n_5564, n_5565);
  not g16399 (n_5566, n10927);
  and g16400 (n10928, n_5513, n_5566);
  and g16401 (n10929, n10838, n10849);
  not g16402 (n_5567, n10850);
  not g16403 (n_5568, n10929);
  and g16404 (n10930, n_5567, n_5568);
  not g16405 (n_5569, n10928);
  and g16406 (n10931, n_5569, n10930);
  not g16407 (n_5570, n10931);
  and g16408 (n10932, n_5567, n_5570);
  not g16409 (n_5571, n10835);
  not g16410 (n_5572, n10932);
  and g16411 (n10933, n_5571, n_5572);
  not g16412 (n_5573, n10933);
  and g16413 (n10934, n_5486, n_5573);
  not g16414 (n_5574, n10818);
  and g16415 (n10935, n10806, n_5574);
  and g16416 (n10936, n_5474, n_5574);
  not g16417 (n_5575, n10935);
  not g16418 (n_5576, n10936);
  and g16419 (n10937, n_5575, n_5576);
  not g16420 (n_5577, n10934);
  not g16421 (n_5578, n10937);
  and g16422 (n10938, n_5577, n_5578);
  not g16423 (n_5579, n10938);
  and g16424 (n10939, n_5574, n_5579);
  not g16425 (n_5580, n10804);
  and g16426 (n10940, n10792, n_5580);
  and g16427 (n10941, n_5464, n_5580);
  not g16428 (n_5581, n10940);
  not g16429 (n_5582, n10941);
  and g16430 (n10942, n_5581, n_5582);
  not g16431 (n_5583, n10939);
  not g16432 (n_5584, n10942);
  and g16433 (n10943, n_5583, n_5584);
  not g16434 (n_5585, n10943);
  and g16435 (n10944, n_5580, n_5585);
  not g16436 (n_5586, n10778);
  and g16437 (n10945, n_5586, n10789);
  not g16438 (n_5587, n10790);
  not g16439 (n_5588, n10945);
  and g16440 (n10946, n_5587, n_5588);
  not g16441 (n_5589, n10944);
  and g16442 (n10947, n_5589, n10946);
  not g16443 (n_5590, n10947);
  and g16444 (n10948, n_5587, n_5590);
  not g16445 (n_5591, n10776);
  not g16446 (n_5592, n10948);
  and g16447 (n10949, n_5591, n_5592);
  not g16448 (n_5593, n10949);
  and g16449 (n10950, n_5441, n_5593);
  not g16450 (n_5594, n10758);
  not g16451 (n_5595, n10950);
  and g16452 (n10951, n_5594, n_5595);
  not g16453 (n_5596, n10951);
  and g16454 (n10952, n_5426, n_5596);
  not g16455 (n_5597, n10740);
  not g16456 (n_5598, n10952);
  and g16457 (n10953, n_5597, n_5598);
  not g16458 (n_5599, n10953);
  and g16459 (n10954, n_5411, n_5599);
  not g16460 (n_5600, n10723);
  and g16461 (n10955, n10711, n_5600);
  and g16462 (n10956, n_5399, n_5600);
  not g16463 (n_5601, n10955);
  not g16464 (n_5602, n10956);
  and g16465 (n10957, n_5601, n_5602);
  not g16466 (n_5603, n10954);
  not g16467 (n_5604, n10957);
  and g16468 (n10958, n_5603, n_5604);
  not g16469 (n_5605, n10958);
  and g16470 (n10959, n_5600, n_5605);
  not g16471 (n_5606, n10709);
  and g16472 (n10960, n10697, n_5606);
  and g16473 (n10961, n_5389, n_5606);
  not g16474 (n_5607, n10960);
  not g16475 (n_5608, n10961);
  and g16476 (n10962, n_5607, n_5608);
  not g16477 (n_5609, n10959);
  not g16478 (n_5610, n10962);
  and g16479 (n10963, n_5609, n_5610);
  not g16480 (n_5611, n10963);
  and g16481 (n10964, n_5606, n_5611);
  not g16482 (n_5612, n10683);
  and g16483 (n10965, n_5612, n10694);
  not g16484 (n_5613, n10695);
  not g16485 (n_5614, n10965);
  and g16486 (n10966, n_5613, n_5614);
  not g16487 (n_5615, n10964);
  and g16488 (n10967, n_5615, n10966);
  not g16489 (n_5616, n10967);
  and g16490 (n10968, n_5613, n_5616);
  not g16491 (n_5617, n10681);
  not g16492 (n_5618, n10968);
  and g16493 (n10969, n_5617, n_5618);
  not g16494 (n_5619, n10969);
  and g16495 (n10970, n_5367, n_5619);
  not g16496 (n_5620, n10663);
  not g16497 (n_5621, n10970);
  and g16498 (n10971, n_5620, n_5621);
  not g16499 (n_5622, n10971);
  and g16500 (n10972, n_5352, n_5622);
  not g16501 (n_5623, n10645);
  not g16502 (n_5624, n10972);
  and g16503 (n10973, n_5623, n_5624);
  not g16504 (n_5625, n10973);
  and g16505 (n10974, n_5337, n_5625);
  not g16506 (n_5626, n10628);
  and g16507 (n10975, n10616, n_5626);
  and g16508 (n10976, n_5325, n_5626);
  not g16509 (n_5627, n10975);
  not g16510 (n_5628, n10976);
  and g16511 (n10977, n_5627, n_5628);
  not g16512 (n_5629, n10974);
  not g16513 (n_5630, n10977);
  and g16514 (n10978, n_5629, n_5630);
  not g16515 (n_5631, n10978);
  and g16516 (n10979, n_5626, n_5631);
  not g16517 (n_5632, n10614);
  and g16518 (n10980, n10602, n_5632);
  and g16519 (n10981, n_5315, n_5632);
  not g16520 (n_5633, n10980);
  not g16521 (n_5634, n10981);
  and g16522 (n10982, n_5633, n_5634);
  not g16523 (n_5635, n10979);
  not g16524 (n_5636, n10982);
  and g16525 (n10983, n_5635, n_5636);
  not g16526 (n_5637, n10983);
  and g16527 (n10984, n_5632, n_5637);
  not g16528 (n_5638, n10588);
  and g16529 (n10985, n_5638, n10599);
  not g16530 (n_5639, n10600);
  not g16531 (n_5640, n10985);
  and g16532 (n10986, n_5639, n_5640);
  not g16533 (n_5641, n10984);
  and g16534 (n10987, n_5641, n10986);
  not g16535 (n_5642, n10987);
  and g16536 (n10988, n_5639, n_5642);
  not g16537 (n_5643, n10586);
  not g16538 (n_5644, n10988);
  and g16539 (n10989, n_5643, n_5644);
  not g16540 (n_5645, n10989);
  and g16541 (n10990, n_5293, n_5645);
  not g16542 (n_5646, n10568);
  not g16543 (n_5647, n10990);
  and g16544 (n10991, n_5646, n_5647);
  not g16545 (n_5648, n10991);
  and g16546 (n10992, n_5278, n_5648);
  not g16547 (n_5649, n10551);
  and g16548 (n10993, n10539, n_5649);
  and g16549 (n10994, n_5266, n_5649);
  not g16550 (n_5650, n10993);
  not g16551 (n_5651, n10994);
  and g16552 (n10995, n_5650, n_5651);
  not g16553 (n_5652, n10992);
  not g16554 (n_5653, n10995);
  and g16555 (n10996, n_5652, n_5653);
  not g16556 (n_5654, n10996);
  and g16557 (n10997, n_5649, n_5654);
  not g16558 (n_5655, n10537);
  and g16559 (n10998, n10525, n_5655);
  and g16560 (n10999, n_5256, n_5655);
  not g16561 (n_5656, n10998);
  not g16562 (n_5657, n10999);
  and g16563 (n11000, n_5656, n_5657);
  not g16564 (n_5658, n10997);
  not g16565 (n_5659, n11000);
  and g16566 (n11001, n_5658, n_5659);
  not g16567 (n_5660, n11001);
  and g16568 (n11002, n_5655, n_5660);
  not g16569 (n_5661, n10523);
  and g16570 (n11003, n10511, n_5661);
  and g16571 (n11004, n_5246, n_5661);
  not g16572 (n_5662, n11003);
  not g16573 (n_5663, n11004);
  and g16574 (n11005, n_5662, n_5663);
  not g16575 (n_5664, n11002);
  not g16576 (n_5665, n11005);
  and g16577 (n11006, n_5664, n_5665);
  not g16578 (n_5666, n11006);
  and g16579 (n11007, n_5661, n_5666);
  not g16580 (n_5667, n10509);
  and g16581 (n11008, n10497, n_5667);
  and g16582 (n11009, n_5236, n_5667);
  not g16583 (n_5668, n11008);
  not g16584 (n_5669, n11009);
  and g16585 (n11010, n_5668, n_5669);
  not g16586 (n_5670, n11007);
  not g16587 (n_5671, n11010);
  and g16588 (n11011, n_5670, n_5671);
  not g16589 (n_5672, n11011);
  and g16590 (n11012, n_5667, n_5672);
  not g16591 (n_5673, n10495);
  and g16592 (n11013, n10483, n_5673);
  and g16593 (n11014, n_5226, n_5673);
  not g16594 (n_5674, n11013);
  not g16595 (n_5675, n11014);
  and g16596 (n11015, n_5674, n_5675);
  not g16597 (n_5676, n11012);
  not g16598 (n_5677, n11015);
  and g16599 (n11016, n_5676, n_5677);
  not g16600 (n_5678, n11016);
  and g16601 (n11017, n_5673, n_5678);
  not g16602 (n_5679, n10481);
  and g16603 (n11018, n10469, n_5679);
  and g16604 (n11019, n_5216, n_5679);
  not g16605 (n_5680, n11018);
  not g16606 (n_5681, n11019);
  and g16607 (n11020, n_5680, n_5681);
  not g16608 (n_5682, n11017);
  not g16609 (n_5683, n11020);
  and g16610 (n11021, n_5682, n_5683);
  not g16611 (n_5684, n11021);
  and g16612 (n11022, n_5679, n_5684);
  not g16613 (n_5685, n10467);
  and g16614 (n11023, n10455, n_5685);
  and g16615 (n11024, n_5206, n_5685);
  not g16616 (n_5686, n11023);
  not g16617 (n_5687, n11024);
  and g16618 (n11025, n_5686, n_5687);
  not g16619 (n_5688, n11022);
  not g16620 (n_5689, n11025);
  and g16621 (n11026, n_5688, n_5689);
  not g16622 (n_5690, n11026);
  and g16623 (n11027, n_5685, n_5690);
  and g16624 (n11028, n10427, n_5173);
  and g16625 (n11029, n_5172, n11028);
  not g16626 (n_5691, n11029);
  and g16627 (n11030, n_5176, n_5691);
  not g16628 (n_5692, n11027);
  and g16629 (n11031, n_5692, n11030);
  and g16630 (n11032, n71, n_712);
  and g16631 (n11033, n_566, n9867);
  and g16632 (n11034, n_560, n10434);
  and g16638 (n11037, n4715, n9870);
  not g16641 (n_5697, n11038);
  and g16642 (n11039, \a[5] , n_5697);
  not g16643 (n_5698, n11039);
  and g16644 (n11040, n_5697, n_5698);
  and g16645 (n11041, \a[5] , n_5698);
  not g16646 (n_5699, n11040);
  not g16647 (n_5700, n11041);
  and g16648 (n11042, n_5699, n_5700);
  not g16649 (n_5701, n11031);
  and g16650 (n11043, n_5692, n_5701);
  and g16651 (n11044, n11030, n_5701);
  not g16652 (n_5702, n11043);
  not g16653 (n_5703, n11044);
  and g16654 (n11045, n_5702, n_5703);
  not g16655 (n_5704, n11042);
  not g16656 (n_5705, n11045);
  and g16657 (n11046, n_5704, n_5705);
  not g16658 (n_5706, n11046);
  and g16659 (n11047, n_5701, n_5706);
  not g16660 (n_5707, n10448);
  and g16661 (n11048, n10446, n_5707);
  not g16662 (n_5708, n11048);
  and g16663 (n11049, n_5192, n_5708);
  not g16664 (n_5709, n11047);
  and g16665 (n11050, n_5709, n11049);
  and g16666 (n11051, \a[1] , n_10);
  not g16667 (n_5711, \a[1] );
  and g16668 (n11052, n_5711, \a[2] );
  not g16669 (n_5712, n11051);
  not g16670 (n_5713, n11052);
  and g16671 (n11053, n_5712, n_5713);
  not g16672 (n_5715, \a[0] );
  and g16673 (n11054, n_5715, n_5711);
  not g16674 (n_5716, n11053);
  and g16675 (n11055, n_5716, n11054);
  and g16676 (n11056, n_712, n11055);
  and g16677 (n11057, \a[0] , n_5716);
  and g16678 (n11058, n4522, n11057);
  not g16679 (n_5717, n11056);
  not g16680 (n_5718, n11058);
  and g16681 (n11059, n_5717, n_5718);
  not g16682 (n_5719, n11059);
  and g16683 (n11060, \a[2] , n_5719);
  not g16684 (n_5720, n11060);
  and g16685 (n11061, n_5719, n_5720);
  and g16686 (n11062, \a[2] , n_5720);
  not g16687 (n_5721, n11061);
  not g16688 (n_5722, n11062);
  and g16689 (n11063, n_5721, n_5722);
  and g16690 (n11064, n71, n_560);
  and g16691 (n11065, n_565, n9867);
  and g16692 (n11066, n_566, n10434);
  and g16698 (n11069, n4067, n9870);
  not g16701 (n_5727, n11070);
  and g16702 (n11071, \a[5] , n_5727);
  not g16703 (n_5728, n11071);
  and g16704 (n11072, \a[5] , n_5728);
  and g16705 (n11073, n_5727, n_5728);
  not g16706 (n_5729, n11072);
  not g16707 (n_5730, n11073);
  and g16708 (n11074, n_5729, n_5730);
  not g16709 (n_5731, n11063);
  not g16710 (n_5732, n11074);
  and g16711 (n11075, n_5731, n_5732);
  not g16712 (n_5733, n11075);
  and g16713 (n11076, n_5731, n_5733);
  and g16714 (n11077, n_5732, n_5733);
  not g16715 (n_5734, n11076);
  not g16716 (n_5735, n11077);
  and g16717 (n11078, n_5734, n_5735);
  and g16718 (n11079, n_5688, n_5690);
  and g16719 (n11080, n_5689, n_5690);
  not g16720 (n_5736, n11079);
  not g16721 (n_5737, n11080);
  and g16722 (n11081, n_5736, n_5737);
  not g16723 (n_5738, n11078);
  not g16724 (n_5739, n11081);
  and g16725 (n11082, n_5738, n_5739);
  not g16726 (n_5740, n11082);
  and g16727 (n11083, n_5733, n_5740);
  and g16728 (n11084, n11042, n_5703);
  and g16729 (n11085, n_5702, n11084);
  not g16730 (n_5741, n11085);
  and g16731 (n11086, n_5706, n_5741);
  not g16732 (n_5742, n11083);
  and g16733 (n11087, n_5742, n11086);
  and g16734 (n11088, n_5738, n_5740);
  and g16735 (n11089, n_5739, n_5740);
  not g16736 (n_5743, n11088);
  not g16737 (n_5744, n11089);
  and g16738 (n11090, n_5743, n_5744);
  and g16739 (n11091, n71, n_566);
  and g16740 (n11092, n_535, n9867);
  and g16741 (n11093, n_565, n10434);
  and g16747 (n11096, n4477, n9870);
  not g16750 (n_5749, n11097);
  and g16751 (n11098, \a[5] , n_5749);
  not g16752 (n_5750, n11098);
  and g16753 (n11099, n_5749, n_5750);
  and g16754 (n11100, \a[5] , n_5750);
  not g16755 (n_5751, n11099);
  not g16756 (n_5752, n11100);
  and g16757 (n11101, n_5751, n_5752);
  and g16758 (n11102, n_5682, n_5684);
  and g16759 (n11103, n_5683, n_5684);
  not g16760 (n_5753, n11102);
  not g16761 (n_5754, n11103);
  and g16762 (n11104, n_5753, n_5754);
  not g16763 (n_5755, n11101);
  not g16764 (n_5756, n11104);
  and g16765 (n11105, n_5755, n_5756);
  not g16766 (n_5757, n11105);
  and g16767 (n11106, n_5755, n_5757);
  and g16768 (n11107, n_5756, n_5757);
  not g16769 (n_5758, n11106);
  not g16770 (n_5759, n11107);
  and g16771 (n11108, n_5758, n_5759);
  and g16772 (n11109, n71, n_565);
  and g16773 (n11110, n_480, n9867);
  and g16774 (n11111, n_535, n10434);
  and g16780 (n11114, n4558, n9870);
  not g16783 (n_5764, n11115);
  and g16784 (n11116, \a[5] , n_5764);
  not g16785 (n_5765, n11116);
  and g16786 (n11117, n_5764, n_5765);
  and g16787 (n11118, \a[5] , n_5765);
  not g16788 (n_5766, n11117);
  not g16789 (n_5767, n11118);
  and g16790 (n11119, n_5766, n_5767);
  and g16791 (n11120, n_5676, n_5678);
  and g16792 (n11121, n_5677, n_5678);
  not g16793 (n_5768, n11120);
  not g16794 (n_5769, n11121);
  and g16795 (n11122, n_5768, n_5769);
  not g16796 (n_5770, n11119);
  not g16797 (n_5771, n11122);
  and g16798 (n11123, n_5770, n_5771);
  not g16799 (n_5772, n11123);
  and g16800 (n11124, n_5770, n_5772);
  and g16801 (n11125, n_5771, n_5772);
  not g16802 (n_5773, n11124);
  not g16803 (n_5774, n11125);
  and g16804 (n11126, n_5773, n_5774);
  and g16805 (n11127, n71, n_535);
  and g16806 (n11128, n_485, n9867);
  and g16807 (n11129, n_480, n10434);
  and g16813 (n11132, n3818, n9870);
  not g16816 (n_5779, n11133);
  and g16817 (n11134, \a[5] , n_5779);
  not g16818 (n_5780, n11134);
  and g16819 (n11135, n_5779, n_5780);
  and g16820 (n11136, \a[5] , n_5780);
  not g16821 (n_5781, n11135);
  not g16822 (n_5782, n11136);
  and g16823 (n11137, n_5781, n_5782);
  and g16824 (n11138, n_5670, n_5672);
  and g16825 (n11139, n_5671, n_5672);
  not g16826 (n_5783, n11138);
  not g16827 (n_5784, n11139);
  and g16828 (n11140, n_5783, n_5784);
  not g16829 (n_5785, n11137);
  not g16830 (n_5786, n11140);
  and g16831 (n11141, n_5785, n_5786);
  not g16832 (n_5787, n11141);
  and g16833 (n11142, n_5785, n_5787);
  and g16834 (n11143, n_5786, n_5787);
  not g16835 (n_5788, n11142);
  not g16836 (n_5789, n11143);
  and g16837 (n11144, n_5788, n_5789);
  and g16838 (n11145, n71, n_480);
  and g16839 (n11146, n_484, n9867);
  and g16840 (n11147, n_485, n10434);
  and g16846 (n11150, n3627, n9870);
  not g16849 (n_5794, n11151);
  and g16850 (n11152, \a[5] , n_5794);
  not g16851 (n_5795, n11152);
  and g16852 (n11153, n_5794, n_5795);
  and g16853 (n11154, \a[5] , n_5795);
  not g16854 (n_5796, n11153);
  not g16855 (n_5797, n11154);
  and g16856 (n11155, n_5796, n_5797);
  and g16857 (n11156, n_5664, n_5666);
  and g16858 (n11157, n_5665, n_5666);
  not g16859 (n_5798, n11156);
  not g16860 (n_5799, n11157);
  and g16861 (n11158, n_5798, n_5799);
  not g16862 (n_5800, n11155);
  not g16863 (n_5801, n11158);
  and g16864 (n11159, n_5800, n_5801);
  not g16865 (n_5802, n11159);
  and g16866 (n11160, n_5800, n_5802);
  and g16867 (n11161, n_5801, n_5802);
  not g16868 (n_5803, n11160);
  not g16869 (n_5804, n11161);
  and g16870 (n11162, n_5803, n_5804);
  and g16871 (n11163, n71, n_485);
  and g16872 (n11164, n_415, n9867);
  and g16873 (n11165, n_484, n10434);
  and g16879 (n11168, n4084, n9870);
  not g16882 (n_5809, n11169);
  and g16883 (n11170, \a[5] , n_5809);
  not g16884 (n_5810, n11170);
  and g16885 (n11171, n_5809, n_5810);
  and g16886 (n11172, \a[5] , n_5810);
  not g16887 (n_5811, n11171);
  not g16888 (n_5812, n11172);
  and g16889 (n11173, n_5811, n_5812);
  and g16890 (n11174, n_5658, n_5660);
  and g16891 (n11175, n_5659, n_5660);
  not g16892 (n_5813, n11174);
  not g16893 (n_5814, n11175);
  and g16894 (n11176, n_5813, n_5814);
  not g16895 (n_5815, n11173);
  not g16896 (n_5816, n11176);
  and g16897 (n11177, n_5815, n_5816);
  not g16898 (n_5817, n11177);
  and g16899 (n11178, n_5815, n_5817);
  and g16900 (n11179, n_5816, n_5817);
  not g16901 (n_5818, n11178);
  not g16902 (n_5819, n11179);
  and g16903 (n11180, n_5818, n_5819);
  and g16904 (n11181, n71, n_484);
  and g16905 (n11182, n_236, n9867);
  and g16906 (n11183, n_415, n10434);
  and g16912 (n11186, n3715, n9870);
  not g16915 (n_5824, n11187);
  and g16916 (n11188, \a[5] , n_5824);
  not g16917 (n_5825, n11188);
  and g16918 (n11189, n_5824, n_5825);
  and g16919 (n11190, \a[5] , n_5825);
  not g16920 (n_5826, n11189);
  not g16921 (n_5827, n11190);
  and g16922 (n11191, n_5826, n_5827);
  and g16923 (n11192, n_5652, n_5654);
  and g16924 (n11193, n_5653, n_5654);
  not g16925 (n_5828, n11192);
  not g16926 (n_5829, n11193);
  and g16927 (n11194, n_5828, n_5829);
  not g16928 (n_5830, n11191);
  not g16929 (n_5831, n11194);
  and g16930 (n11195, n_5830, n_5831);
  not g16931 (n_5832, n11195);
  and g16932 (n11196, n_5830, n_5832);
  and g16933 (n11197, n_5831, n_5832);
  not g16934 (n_5833, n11196);
  not g16935 (n_5834, n11197);
  and g16936 (n11198, n_5833, n_5834);
  and g16937 (n11199, n10568, n10990);
  not g16938 (n_5835, n11199);
  and g16939 (n11200, n_5648, n_5835);
  and g16940 (n11201, n71, n_415);
  and g16941 (n11202, n_237, n9867);
  and g16942 (n11203, n_236, n10434);
  not g16943 (n_5836, n11202);
  not g16944 (n_5837, n11203);
  and g16945 (n11204, n_5836, n_5837);
  not g16946 (n_5838, n11201);
  and g16947 (n11205, n_5838, n11204);
  and g16948 (n11206, n_4684, n11205);
  and g16949 (n11207, n_680, n11205);
  not g16950 (n_5839, n11206);
  not g16951 (n_5840, n11207);
  and g16952 (n11208, n_5839, n_5840);
  not g16953 (n_5841, n11208);
  and g16954 (n11209, \a[5] , n_5841);
  and g16955 (n11210, n_3, n11208);
  not g16956 (n_5842, n11209);
  not g16957 (n_5843, n11210);
  and g16958 (n11211, n_5842, n_5843);
  not g16959 (n_5844, n11211);
  and g16960 (n11212, n11200, n_5844);
  and g16961 (n11213, n10586, n10988);
  not g16962 (n_5845, n11213);
  and g16963 (n11214, n_5645, n_5845);
  and g16964 (n11215, n71, n_236);
  and g16965 (n11216, n_260, n9867);
  and g16966 (n11217, n_237, n10434);
  not g16967 (n_5846, n11216);
  not g16968 (n_5847, n11217);
  and g16969 (n11218, n_5846, n_5847);
  not g16970 (n_5848, n11215);
  and g16971 (n11219, n_5848, n11218);
  and g16972 (n11220, n_4684, n11219);
  and g16973 (n11221, n_1208, n11219);
  not g16974 (n_5849, n11220);
  not g16975 (n_5850, n11221);
  and g16976 (n11222, n_5849, n_5850);
  not g16977 (n_5851, n11222);
  and g16978 (n11223, \a[5] , n_5851);
  and g16979 (n11224, n_3, n11222);
  not g16980 (n_5852, n11223);
  not g16981 (n_5853, n11224);
  and g16982 (n11225, n_5852, n_5853);
  not g16983 (n_5854, n11225);
  and g16984 (n11226, n11214, n_5854);
  and g16985 (n11227, n71, n_237);
  and g16986 (n11228, n_275, n9867);
  and g16987 (n11229, n_260, n10434);
  and g16993 (n11232, n3331, n9870);
  not g16996 (n_5859, n11233);
  and g16997 (n11234, \a[5] , n_5859);
  not g16998 (n_5860, n11234);
  and g16999 (n11235, n_5859, n_5860);
  and g17000 (n11236, \a[5] , n_5860);
  not g17001 (n_5861, n11235);
  not g17002 (n_5862, n11236);
  and g17003 (n11237, n_5861, n_5862);
  not g17004 (n_5863, n10986);
  and g17005 (n11238, n10984, n_5863);
  not g17006 (n_5864, n11238);
  and g17007 (n11239, n_5642, n_5864);
  not g17008 (n_5865, n11237);
  and g17009 (n11240, n_5865, n11239);
  not g17010 (n_5866, n11240);
  and g17011 (n11241, n_5865, n_5866);
  and g17012 (n11242, n11239, n_5866);
  not g17013 (n_5867, n11241);
  not g17014 (n_5868, n11242);
  and g17015 (n11243, n_5867, n_5868);
  and g17016 (n11244, n71, n_260);
  and g17017 (n11245, n_281, n9867);
  and g17018 (n11246, n_275, n10434);
  and g17024 (n11249, n4179, n9870);
  not g17027 (n_5873, n11250);
  and g17028 (n11251, \a[5] , n_5873);
  not g17029 (n_5874, n11251);
  and g17030 (n11252, n_5873, n_5874);
  and g17031 (n11253, \a[5] , n_5874);
  not g17032 (n_5875, n11252);
  not g17033 (n_5876, n11253);
  and g17034 (n11254, n_5875, n_5876);
  and g17035 (n11255, n_5635, n_5637);
  and g17036 (n11256, n_5636, n_5637);
  not g17037 (n_5877, n11255);
  not g17038 (n_5878, n11256);
  and g17039 (n11257, n_5877, n_5878);
  not g17040 (n_5879, n11254);
  not g17041 (n_5880, n11257);
  and g17042 (n11258, n_5879, n_5880);
  not g17043 (n_5881, n11258);
  and g17044 (n11259, n_5879, n_5881);
  and g17045 (n11260, n_5880, n_5881);
  not g17046 (n_5882, n11259);
  not g17047 (n_5883, n11260);
  and g17048 (n11261, n_5882, n_5883);
  and g17049 (n11262, n71, n_275);
  and g17050 (n11263, n_286, n9867);
  and g17051 (n11264, n_281, n10434);
  and g17057 (n11267, n4204, n9870);
  not g17060 (n_5888, n11268);
  and g17061 (n11269, \a[5] , n_5888);
  not g17062 (n_5889, n11269);
  and g17063 (n11270, n_5888, n_5889);
  and g17064 (n11271, \a[5] , n_5889);
  not g17065 (n_5890, n11270);
  not g17066 (n_5891, n11271);
  and g17067 (n11272, n_5890, n_5891);
  and g17068 (n11273, n_5629, n_5631);
  and g17069 (n11274, n_5630, n_5631);
  not g17070 (n_5892, n11273);
  not g17071 (n_5893, n11274);
  and g17072 (n11275, n_5892, n_5893);
  not g17073 (n_5894, n11272);
  not g17074 (n_5895, n11275);
  and g17075 (n11276, n_5894, n_5895);
  not g17076 (n_5896, n11276);
  and g17077 (n11277, n_5894, n_5896);
  and g17078 (n11278, n_5895, n_5896);
  not g17079 (n_5897, n11277);
  not g17080 (n_5898, n11278);
  and g17081 (n11279, n_5897, n_5898);
  and g17082 (n11280, n10645, n10972);
  not g17083 (n_5899, n11280);
  and g17084 (n11281, n_5625, n_5899);
  and g17085 (n11282, n71, n_281);
  and g17086 (n11283, n_293, n9867);
  and g17087 (n11284, n_286, n10434);
  not g17088 (n_5900, n11283);
  not g17089 (n_5901, n11284);
  and g17090 (n11285, n_5900, n_5901);
  not g17091 (n_5902, n11282);
  and g17092 (n11286, n_5902, n11285);
  and g17093 (n11287, n_4684, n11286);
  and g17094 (n11288, n_1228, n11286);
  not g17095 (n_5903, n11287);
  not g17096 (n_5904, n11288);
  and g17097 (n11289, n_5903, n_5904);
  not g17098 (n_5905, n11289);
  and g17099 (n11290, \a[5] , n_5905);
  and g17100 (n11291, n_3, n11289);
  not g17101 (n_5906, n11290);
  not g17102 (n_5907, n11291);
  and g17103 (n11292, n_5906, n_5907);
  not g17104 (n_5908, n11292);
  and g17105 (n11293, n11281, n_5908);
  and g17106 (n11294, n10663, n10970);
  not g17107 (n_5909, n11294);
  and g17108 (n11295, n_5622, n_5909);
  and g17109 (n11296, n71, n_286);
  and g17110 (n11297, n_295, n9867);
  and g17111 (n11298, n_293, n10434);
  not g17112 (n_5910, n11297);
  not g17113 (n_5911, n11298);
  and g17114 (n11299, n_5910, n_5911);
  not g17115 (n_5912, n11296);
  and g17116 (n11300, n_5912, n11299);
  and g17117 (n11301, n_4684, n11300);
  and g17118 (n11302, n_1134, n11300);
  not g17119 (n_5913, n11301);
  not g17120 (n_5914, n11302);
  and g17121 (n11303, n_5913, n_5914);
  not g17122 (n_5915, n11303);
  and g17123 (n11304, \a[5] , n_5915);
  and g17124 (n11305, n_3, n11303);
  not g17125 (n_5916, n11304);
  not g17126 (n_5917, n11305);
  and g17127 (n11306, n_5916, n_5917);
  not g17128 (n_5918, n11306);
  and g17129 (n11307, n11295, n_5918);
  and g17130 (n11308, n10681, n10968);
  not g17131 (n_5919, n11308);
  and g17132 (n11309, n_5619, n_5919);
  and g17133 (n11310, n71, n_293);
  and g17134 (n11311, n_298, n9867);
  and g17135 (n11312, n_295, n10434);
  not g17136 (n_5920, n11311);
  not g17137 (n_5921, n11312);
  and g17138 (n11313, n_5920, n_5921);
  not g17139 (n_5922, n11310);
  and g17140 (n11314, n_5922, n11313);
  and g17141 (n11315, n_4684, n11314);
  and g17142 (n11316, n_1789, n11314);
  not g17143 (n_5923, n11315);
  not g17144 (n_5924, n11316);
  and g17145 (n11317, n_5923, n_5924);
  not g17146 (n_5925, n11317);
  and g17147 (n11318, \a[5] , n_5925);
  and g17148 (n11319, n_3, n11317);
  not g17149 (n_5926, n11318);
  not g17150 (n_5927, n11319);
  and g17151 (n11320, n_5926, n_5927);
  not g17152 (n_5928, n11320);
  and g17153 (n11321, n11309, n_5928);
  and g17154 (n11322, n71, n_295);
  and g17155 (n11323, n_299, n9867);
  and g17156 (n11324, n_298, n10434);
  and g17162 (n11327, n4848, n9870);
  not g17165 (n_5933, n11328);
  and g17166 (n11329, \a[5] , n_5933);
  not g17167 (n_5934, n11329);
  and g17168 (n11330, n_5933, n_5934);
  and g17169 (n11331, \a[5] , n_5934);
  not g17170 (n_5935, n11330);
  not g17171 (n_5936, n11331);
  and g17172 (n11332, n_5935, n_5936);
  not g17173 (n_5937, n10966);
  and g17174 (n11333, n10964, n_5937);
  not g17175 (n_5938, n11333);
  and g17176 (n11334, n_5616, n_5938);
  not g17177 (n_5939, n11332);
  and g17178 (n11335, n_5939, n11334);
  not g17179 (n_5940, n11335);
  and g17180 (n11336, n_5939, n_5940);
  and g17181 (n11337, n11334, n_5940);
  not g17182 (n_5941, n11336);
  not g17183 (n_5942, n11337);
  and g17184 (n11338, n_5941, n_5942);
  and g17185 (n11339, n71, n_298);
  and g17186 (n11340, n_300, n9867);
  and g17187 (n11341, n_299, n10434);
  and g17193 (n11344, n5114, n9870);
  not g17196 (n_5947, n11345);
  and g17197 (n11346, \a[5] , n_5947);
  not g17198 (n_5948, n11346);
  and g17199 (n11347, n_5947, n_5948);
  and g17200 (n11348, \a[5] , n_5948);
  not g17201 (n_5949, n11347);
  not g17202 (n_5950, n11348);
  and g17203 (n11349, n_5949, n_5950);
  and g17204 (n11350, n_5609, n_5611);
  and g17205 (n11351, n_5610, n_5611);
  not g17206 (n_5951, n11350);
  not g17207 (n_5952, n11351);
  and g17208 (n11352, n_5951, n_5952);
  not g17209 (n_5953, n11349);
  not g17210 (n_5954, n11352);
  and g17211 (n11353, n_5953, n_5954);
  not g17212 (n_5955, n11353);
  and g17213 (n11354, n_5953, n_5955);
  and g17214 (n11355, n_5954, n_5955);
  not g17215 (n_5956, n11354);
  not g17216 (n_5957, n11355);
  and g17217 (n11356, n_5956, n_5957);
  and g17218 (n11357, n71, n_299);
  and g17219 (n11358, n_301, n9867);
  and g17220 (n11359, n_300, n10434);
  and g17226 (n11362, n5139, n9870);
  not g17229 (n_5962, n11363);
  and g17230 (n11364, \a[5] , n_5962);
  not g17231 (n_5963, n11364);
  and g17232 (n11365, n_5962, n_5963);
  and g17233 (n11366, \a[5] , n_5963);
  not g17234 (n_5964, n11365);
  not g17235 (n_5965, n11366);
  and g17236 (n11367, n_5964, n_5965);
  and g17237 (n11368, n_5603, n_5605);
  and g17238 (n11369, n_5604, n_5605);
  not g17239 (n_5966, n11368);
  not g17240 (n_5967, n11369);
  and g17241 (n11370, n_5966, n_5967);
  not g17242 (n_5968, n11367);
  not g17243 (n_5969, n11370);
  and g17244 (n11371, n_5968, n_5969);
  not g17245 (n_5970, n11371);
  and g17246 (n11372, n_5968, n_5970);
  and g17247 (n11373, n_5969, n_5970);
  not g17248 (n_5971, n11372);
  not g17249 (n_5972, n11373);
  and g17250 (n11374, n_5971, n_5972);
  and g17251 (n11375, n10740, n10952);
  not g17252 (n_5973, n11375);
  and g17253 (n11376, n_5599, n_5973);
  and g17254 (n11377, n71, n_300);
  and g17255 (n11378, n_302, n9867);
  and g17256 (n11379, n_301, n10434);
  not g17257 (n_5974, n11378);
  not g17258 (n_5975, n11379);
  and g17259 (n11380, n_5974, n_5975);
  not g17260 (n_5976, n11377);
  and g17261 (n11381, n_5976, n11380);
  and g17262 (n11382, n_4684, n11381);
  and g17263 (n11383, n_1801, n11381);
  not g17264 (n_5977, n11382);
  not g17265 (n_5978, n11383);
  and g17266 (n11384, n_5977, n_5978);
  not g17267 (n_5979, n11384);
  and g17268 (n11385, \a[5] , n_5979);
  and g17269 (n11386, n_3, n11384);
  not g17270 (n_5980, n11385);
  not g17271 (n_5981, n11386);
  and g17272 (n11387, n_5980, n_5981);
  not g17273 (n_5982, n11387);
  and g17274 (n11388, n11376, n_5982);
  and g17275 (n11389, n10758, n10950);
  not g17276 (n_5983, n11389);
  and g17277 (n11390, n_5596, n_5983);
  and g17278 (n11391, n71, n_301);
  and g17279 (n11392, n_303, n9867);
  and g17280 (n11393, n_302, n10434);
  not g17281 (n_5984, n11392);
  not g17282 (n_5985, n11393);
  and g17283 (n11394, n_5984, n_5985);
  not g17284 (n_5986, n11391);
  and g17285 (n11395, n_5986, n11394);
  and g17286 (n11396, n_4684, n11395);
  and g17287 (n11397, n_1672, n11395);
  not g17288 (n_5987, n11396);
  not g17289 (n_5988, n11397);
  and g17290 (n11398, n_5987, n_5988);
  not g17291 (n_5989, n11398);
  and g17292 (n11399, \a[5] , n_5989);
  and g17293 (n11400, n_3, n11398);
  not g17294 (n_5990, n11399);
  not g17295 (n_5991, n11400);
  and g17296 (n11401, n_5990, n_5991);
  not g17297 (n_5992, n11401);
  and g17298 (n11402, n11390, n_5992);
  and g17299 (n11403, n10776, n10948);
  not g17300 (n_5993, n11403);
  and g17301 (n11404, n_5593, n_5993);
  and g17302 (n11405, n71, n_302);
  and g17303 (n11406, n_304, n9867);
  and g17304 (n11407, n_303, n10434);
  not g17305 (n_5994, n11406);
  not g17306 (n_5995, n11407);
  and g17307 (n11408, n_5994, n_5995);
  not g17308 (n_5996, n11405);
  and g17309 (n11409, n_5996, n11408);
  and g17310 (n11410, n_4684, n11409);
  and g17311 (n11411, n_3507, n11409);
  not g17312 (n_5997, n11410);
  not g17313 (n_5998, n11411);
  and g17314 (n11412, n_5997, n_5998);
  not g17315 (n_5999, n11412);
  and g17316 (n11413, \a[5] , n_5999);
  and g17317 (n11414, n_3, n11412);
  not g17318 (n_6000, n11413);
  not g17319 (n_6001, n11414);
  and g17320 (n11415, n_6000, n_6001);
  not g17321 (n_6002, n11415);
  and g17322 (n11416, n11404, n_6002);
  and g17323 (n11417, n71, n_303);
  and g17324 (n11418, n_305, n9867);
  and g17325 (n11419, n_304, n10434);
  and g17331 (n11422, n6007, n9870);
  not g17334 (n_6007, n11423);
  and g17335 (n11424, \a[5] , n_6007);
  not g17336 (n_6008, n11424);
  and g17337 (n11425, n_6007, n_6008);
  and g17338 (n11426, \a[5] , n_6008);
  not g17339 (n_6009, n11425);
  not g17340 (n_6010, n11426);
  and g17341 (n11427, n_6009, n_6010);
  not g17342 (n_6011, n10946);
  and g17343 (n11428, n10944, n_6011);
  not g17344 (n_6012, n11428);
  and g17345 (n11429, n_5590, n_6012);
  not g17346 (n_6013, n11427);
  and g17347 (n11430, n_6013, n11429);
  not g17348 (n_6014, n11430);
  and g17349 (n11431, n_6013, n_6014);
  and g17350 (n11432, n11429, n_6014);
  not g17351 (n_6015, n11431);
  not g17352 (n_6016, n11432);
  and g17353 (n11433, n_6015, n_6016);
  and g17354 (n11434, n71, n_304);
  and g17355 (n11435, n_306, n9867);
  and g17356 (n11436, n_305, n10434);
  and g17362 (n11439, n5834, n9870);
  not g17365 (n_6021, n11440);
  and g17366 (n11441, \a[5] , n_6021);
  not g17367 (n_6022, n11441);
  and g17368 (n11442, n_6021, n_6022);
  and g17369 (n11443, \a[5] , n_6022);
  not g17370 (n_6023, n11442);
  not g17371 (n_6024, n11443);
  and g17372 (n11444, n_6023, n_6024);
  and g17373 (n11445, n_5583, n_5585);
  and g17374 (n11446, n_5584, n_5585);
  not g17375 (n_6025, n11445);
  not g17376 (n_6026, n11446);
  and g17377 (n11447, n_6025, n_6026);
  not g17378 (n_6027, n11444);
  not g17379 (n_6028, n11447);
  and g17380 (n11448, n_6027, n_6028);
  not g17381 (n_6029, n11448);
  and g17382 (n11449, n_6027, n_6029);
  and g17383 (n11450, n_6028, n_6029);
  not g17384 (n_6030, n11449);
  not g17385 (n_6031, n11450);
  and g17386 (n11451, n_6030, n_6031);
  and g17387 (n11452, n71, n_305);
  and g17388 (n11453, n_307, n9867);
  and g17389 (n11454, n_306, n10434);
  and g17395 (n11457, n6143, n9870);
  not g17398 (n_6036, n11458);
  and g17399 (n11459, \a[5] , n_6036);
  not g17400 (n_6037, n11459);
  and g17401 (n11460, n_6036, n_6037);
  and g17402 (n11461, \a[5] , n_6037);
  not g17403 (n_6038, n11460);
  not g17404 (n_6039, n11461);
  and g17405 (n11462, n_6038, n_6039);
  and g17406 (n11463, n_5577, n_5579);
  and g17407 (n11464, n_5578, n_5579);
  not g17408 (n_6040, n11463);
  not g17409 (n_6041, n11464);
  and g17410 (n11465, n_6040, n_6041);
  not g17411 (n_6042, n11462);
  not g17412 (n_6043, n11465);
  and g17413 (n11466, n_6042, n_6043);
  not g17414 (n_6044, n11466);
  and g17415 (n11467, n_6042, n_6044);
  and g17416 (n11468, n_6043, n_6044);
  not g17417 (n_6045, n11467);
  not g17418 (n_6046, n11468);
  and g17419 (n11469, n_6045, n_6046);
  and g17420 (n11470, n10835, n10932);
  not g17421 (n_6047, n11470);
  and g17422 (n11471, n_5573, n_6047);
  and g17423 (n11472, n71, n_306);
  and g17424 (n11473, n_308, n9867);
  and g17425 (n11474, n_307, n10434);
  not g17426 (n_6048, n11473);
  not g17427 (n_6049, n11474);
  and g17428 (n11475, n_6048, n_6049);
  not g17429 (n_6050, n11472);
  and g17430 (n11476, n_6050, n11475);
  and g17431 (n11477, n_4684, n11476);
  and g17432 (n11478, n_2498, n11476);
  not g17433 (n_6051, n11477);
  not g17434 (n_6052, n11478);
  and g17435 (n11479, n_6051, n_6052);
  not g17436 (n_6053, n11479);
  and g17437 (n11480, \a[5] , n_6053);
  and g17438 (n11481, n_3, n11479);
  not g17439 (n_6054, n11480);
  not g17440 (n_6055, n11481);
  and g17441 (n11482, n_6054, n_6055);
  not g17442 (n_6056, n11482);
  and g17443 (n11483, n11471, n_6056);
  not g17444 (n_6057, n10930);
  and g17445 (n11484, n10928, n_6057);
  not g17446 (n_6058, n11484);
  and g17447 (n11485, n_5570, n_6058);
  and g17448 (n11486, n71, n_307);
  and g17449 (n11487, n_309, n9867);
  and g17450 (n11488, n_308, n10434);
  not g17451 (n_6059, n11487);
  not g17452 (n_6060, n11488);
  and g17453 (n11489, n_6059, n_6060);
  not g17454 (n_6061, n11486);
  and g17455 (n11490, n_6061, n11489);
  and g17456 (n11491, n_4684, n11490);
  and g17457 (n11492, n_2511, n11490);
  not g17458 (n_6062, n11491);
  not g17459 (n_6063, n11492);
  and g17460 (n11493, n_6062, n_6063);
  not g17461 (n_6064, n11493);
  and g17462 (n11494, \a[5] , n_6064);
  and g17463 (n11495, n_3, n11493);
  not g17464 (n_6065, n11494);
  not g17465 (n_6066, n11495);
  and g17466 (n11496, n_6065, n_6066);
  not g17467 (n_6067, n11496);
  and g17468 (n11497, n11485, n_6067);
  and g17469 (n11498, n10867, n10926);
  not g17470 (n_6068, n11498);
  and g17471 (n11499, n_5566, n_6068);
  and g17472 (n11500, n71, n_308);
  and g17473 (n11501, n_310, n9867);
  and g17474 (n11502, n_309, n10434);
  not g17475 (n_6069, n11501);
  not g17476 (n_6070, n11502);
  and g17477 (n11503, n_6069, n_6070);
  not g17478 (n_6071, n11500);
  and g17479 (n11504, n_6071, n11503);
  and g17480 (n11505, n_4684, n11504);
  and g17481 (n11506, n_2839, n11504);
  not g17482 (n_6072, n11505);
  not g17483 (n_6073, n11506);
  and g17484 (n11507, n_6072, n_6073);
  not g17485 (n_6074, n11507);
  and g17486 (n11508, \a[5] , n_6074);
  and g17487 (n11509, n_3, n11507);
  not g17488 (n_6075, n11508);
  not g17489 (n_6076, n11509);
  and g17490 (n11510, n_6075, n_6076);
  not g17491 (n_6077, n11510);
  and g17492 (n11511, n11499, n_6077);
  and g17493 (n11512, n71, n_309);
  and g17494 (n11513, n_311, n9867);
  and g17495 (n11514, n_310, n10434);
  and g17501 (n11517, n6541, n9870);
  not g17504 (n_6082, n11518);
  and g17505 (n11519, \a[5] , n_6082);
  not g17506 (n_6083, n11519);
  and g17507 (n11520, n_6082, n_6083);
  and g17508 (n11521, \a[5] , n_6083);
  not g17509 (n_6084, n11520);
  not g17510 (n_6085, n11521);
  and g17511 (n11522, n_6084, n_6085);
  not g17512 (n_6086, n10924);
  and g17513 (n11523, n10922, n_6086);
  not g17514 (n_6087, n11523);
  and g17515 (n11524, n_5563, n_6087);
  not g17516 (n_6088, n11522);
  and g17517 (n11525, n_6088, n11524);
  not g17518 (n_6089, n11525);
  and g17519 (n11526, n_6088, n_6089);
  and g17520 (n11527, n11524, n_6089);
  not g17521 (n_6090, n11526);
  not g17522 (n_6091, n11527);
  and g17523 (n11528, n_6090, n_6091);
  and g17524 (n11529, n_5556, n_5558);
  and g17525 (n11530, n_5557, n_5558);
  not g17526 (n_6092, n11529);
  not g17527 (n_6093, n11530);
  and g17528 (n11531, n_6092, n_6093);
  and g17529 (n11532, n71, n_310);
  and g17530 (n11533, n_312, n9867);
  and g17531 (n11534, n_311, n10434);
  not g17532 (n_6094, n11533);
  not g17533 (n_6095, n11534);
  and g17534 (n11535, n_6094, n_6095);
  not g17535 (n_6096, n11532);
  and g17536 (n11536, n_6096, n11535);
  and g17537 (n11537, n_4684, n11536);
  and g17538 (n11538, n_3239, n11536);
  not g17539 (n_6097, n11537);
  not g17540 (n_6098, n11538);
  and g17541 (n11539, n_6097, n_6098);
  not g17542 (n_6099, n11539);
  and g17543 (n11540, \a[5] , n_6099);
  and g17544 (n11541, n_3, n11539);
  not g17545 (n_6100, n11540);
  not g17546 (n_6101, n11541);
  and g17547 (n11542, n_6100, n_6101);
  not g17548 (n_6102, n11531);
  not g17549 (n_6103, n11542);
  and g17550 (n11543, n_6102, n_6103);
  and g17551 (n11544, n71, n_311);
  and g17552 (n11545, n_313, n9867);
  and g17553 (n11546, n_312, n10434);
  and g17559 (n11549, n6646, n9870);
  not g17562 (n_6108, n11550);
  and g17563 (n11551, \a[5] , n_6108);
  not g17564 (n_6109, n11551);
  and g17565 (n11552, n_6108, n_6109);
  and g17566 (n11553, \a[5] , n_6109);
  not g17567 (n_6110, n11552);
  not g17568 (n_6111, n11553);
  and g17569 (n11554, n_6110, n_6111);
  not g17570 (n_6112, n10893);
  and g17571 (n11555, n_6112, n10904);
  not g17572 (n_6113, n10905);
  not g17573 (n_6114, n11555);
  and g17574 (n11556, n_6113, n_6114);
  not g17575 (n_6115, n11554);
  and g17576 (n11557, n_6115, n11556);
  not g17577 (n_6116, n11557);
  and g17578 (n11558, n_6115, n_6116);
  and g17579 (n11559, n11556, n_6116);
  not g17580 (n_6117, n11558);
  not g17581 (n_6118, n11559);
  and g17582 (n11560, n_6117, n_6118);
  not g17583 (n_6119, n10892);
  and g17584 (n11561, n10890, n_6119);
  not g17585 (n_6120, n11561);
  and g17586 (n11562, n_6112, n_6120);
  and g17587 (n11563, n71, n_312);
  and g17588 (n11564, n_314, n9867);
  and g17589 (n11565, n_313, n10434);
  not g17590 (n_6121, n11564);
  not g17591 (n_6122, n11565);
  and g17592 (n11566, n_6121, n_6122);
  not g17593 (n_6123, n11563);
  and g17594 (n11567, n_6123, n11566);
  and g17595 (n11568, n_4684, n11567);
  and g17596 (n11569, n_2891, n11567);
  not g17597 (n_6124, n11568);
  not g17598 (n_6125, n11569);
  and g17599 (n11570, n_6124, n_6125);
  not g17600 (n_6126, n11570);
  and g17601 (n11571, \a[5] , n_6126);
  and g17602 (n11572, n_3, n11570);
  not g17603 (n_6127, n11571);
  not g17604 (n_6128, n11572);
  and g17605 (n11573, n_6127, n_6128);
  not g17606 (n_6129, n11573);
  and g17607 (n11574, n11562, n_6129);
  and g17608 (n11575, n_316, n10434);
  and g17609 (n11576, n71, n_315);
  not g17610 (n_6130, n11575);
  not g17611 (n_6131, n11576);
  and g17612 (n11577, n_6130, n_6131);
  and g17613 (n11578, n_2588, n9870);
  not g17614 (n_6132, n11578);
  and g17615 (n11579, n11577, n_6132);
  not g17616 (n_6133, n11579);
  and g17617 (n11580, \a[5] , n_6133);
  not g17618 (n_6134, n11580);
  and g17619 (n11581, \a[5] , n_6134);
  and g17620 (n11582, n_6133, n_6134);
  not g17621 (n_6135, n11581);
  not g17622 (n_6136, n11582);
  and g17623 (n11583, n_6135, n_6136);
  and g17624 (n11584, n_13, n_316);
  not g17625 (n_6137, n11584);
  and g17626 (n11585, \a[5] , n_6137);
  not g17627 (n_6138, n11583);
  and g17628 (n11586, n_6138, n11585);
  and g17629 (n11587, n71, n_314);
  and g17630 (n11588, n_316, n9867);
  and g17631 (n11589, n_315, n10434);
  not g17632 (n_6139, n11588);
  not g17633 (n_6140, n11589);
  and g17634 (n11590, n_6139, n_6140);
  not g17635 (n_6141, n11587);
  and g17636 (n11591, n_6141, n11590);
  and g17637 (n11592, n_4684, n11591);
  and g17638 (n11593, n_2612, n11591);
  not g17639 (n_6142, n11592);
  not g17640 (n_6143, n11593);
  and g17641 (n11594, n_6142, n_6143);
  not g17642 (n_6144, n11594);
  and g17643 (n11595, \a[5] , n_6144);
  and g17644 (n11596, n_3, n11594);
  not g17645 (n_6145, n11595);
  not g17646 (n_6146, n11596);
  and g17647 (n11597, n_6145, n_6146);
  not g17648 (n_6147, n11597);
  and g17649 (n11598, n11586, n_6147);
  and g17650 (n11599, n10891, n11598);
  not g17651 (n_6148, n11599);
  and g17652 (n11600, n11598, n_6148);
  and g17653 (n11601, n10891, n_6148);
  not g17654 (n_6149, n11600);
  not g17655 (n_6150, n11601);
  and g17656 (n11602, n_6149, n_6150);
  and g17657 (n11603, n71, n_313);
  and g17658 (n11604, n_315, n9867);
  and g17659 (n11605, n_314, n10434);
  and g17665 (n11608, n6806, n9870);
  not g17668 (n_6155, n11609);
  and g17669 (n11610, \a[5] , n_6155);
  not g17670 (n_6156, n11610);
  and g17671 (n11611, \a[5] , n_6156);
  and g17672 (n11612, n_6155, n_6156);
  not g17673 (n_6157, n11611);
  not g17674 (n_6158, n11612);
  and g17675 (n11613, n_6157, n_6158);
  not g17676 (n_6159, n11602);
  not g17677 (n_6160, n11613);
  and g17678 (n11614, n_6159, n_6160);
  not g17679 (n_6161, n11614);
  and g17680 (n11615, n_6148, n_6161);
  not g17681 (n_6162, n11562);
  and g17682 (n11616, n_6162, n11573);
  not g17683 (n_6163, n11574);
  not g17684 (n_6164, n11616);
  and g17685 (n11617, n_6163, n_6164);
  not g17686 (n_6165, n11615);
  and g17687 (n11618, n_6165, n11617);
  not g17688 (n_6166, n11618);
  and g17689 (n11619, n_6163, n_6166);
  not g17690 (n_6167, n11560);
  not g17691 (n_6168, n11619);
  and g17692 (n11620, n_6167, n_6168);
  not g17693 (n_6169, n11620);
  and g17694 (n11621, n_6116, n_6169);
  and g17695 (n11622, n11531, n11542);
  not g17696 (n_6170, n11543);
  not g17697 (n_6171, n11622);
  and g17698 (n11623, n_6170, n_6171);
  not g17699 (n_6172, n11621);
  and g17700 (n11624, n_6172, n11623);
  not g17701 (n_6173, n11624);
  and g17702 (n11625, n_6170, n_6173);
  not g17703 (n_6174, n11528);
  not g17704 (n_6175, n11625);
  and g17705 (n11626, n_6174, n_6175);
  not g17706 (n_6176, n11626);
  and g17707 (n11627, n_6089, n_6176);
  not g17708 (n_6177, n11511);
  and g17709 (n11628, n11499, n_6177);
  and g17710 (n11629, n_6077, n_6177);
  not g17711 (n_6178, n11628);
  not g17712 (n_6179, n11629);
  and g17713 (n11630, n_6178, n_6179);
  not g17714 (n_6180, n11627);
  not g17715 (n_6181, n11630);
  and g17716 (n11631, n_6180, n_6181);
  not g17717 (n_6182, n11631);
  and g17718 (n11632, n_6177, n_6182);
  not g17719 (n_6183, n11497);
  and g17720 (n11633, n11485, n_6183);
  and g17721 (n11634, n_6067, n_6183);
  not g17722 (n_6184, n11633);
  not g17723 (n_6185, n11634);
  and g17724 (n11635, n_6184, n_6185);
  not g17725 (n_6186, n11632);
  not g17726 (n_6187, n11635);
  and g17727 (n11636, n_6186, n_6187);
  not g17728 (n_6188, n11636);
  and g17729 (n11637, n_6183, n_6188);
  not g17730 (n_6189, n11471);
  and g17731 (n11638, n_6189, n11482);
  not g17732 (n_6190, n11483);
  not g17733 (n_6191, n11638);
  and g17734 (n11639, n_6190, n_6191);
  not g17735 (n_6192, n11637);
  and g17736 (n11640, n_6192, n11639);
  not g17737 (n_6193, n11640);
  and g17738 (n11641, n_6190, n_6193);
  not g17739 (n_6194, n11469);
  not g17740 (n_6195, n11641);
  and g17741 (n11642, n_6194, n_6195);
  not g17742 (n_6196, n11642);
  and g17743 (n11643, n_6044, n_6196);
  not g17744 (n_6197, n11451);
  not g17745 (n_6198, n11643);
  and g17746 (n11644, n_6197, n_6198);
  not g17747 (n_6199, n11644);
  and g17748 (n11645, n_6029, n_6199);
  not g17749 (n_6200, n11433);
  not g17750 (n_6201, n11645);
  and g17751 (n11646, n_6200, n_6201);
  not g17752 (n_6202, n11646);
  and g17753 (n11647, n_6014, n_6202);
  not g17754 (n_6203, n11416);
  and g17755 (n11648, n11404, n_6203);
  and g17756 (n11649, n_6002, n_6203);
  not g17757 (n_6204, n11648);
  not g17758 (n_6205, n11649);
  and g17759 (n11650, n_6204, n_6205);
  not g17760 (n_6206, n11647);
  not g17761 (n_6207, n11650);
  and g17762 (n11651, n_6206, n_6207);
  not g17763 (n_6208, n11651);
  and g17764 (n11652, n_6203, n_6208);
  not g17765 (n_6209, n11402);
  and g17766 (n11653, n11390, n_6209);
  and g17767 (n11654, n_5992, n_6209);
  not g17768 (n_6210, n11653);
  not g17769 (n_6211, n11654);
  and g17770 (n11655, n_6210, n_6211);
  not g17771 (n_6212, n11652);
  not g17772 (n_6213, n11655);
  and g17773 (n11656, n_6212, n_6213);
  not g17774 (n_6214, n11656);
  and g17775 (n11657, n_6209, n_6214);
  not g17776 (n_6215, n11376);
  and g17777 (n11658, n_6215, n11387);
  not g17778 (n_6216, n11388);
  not g17779 (n_6217, n11658);
  and g17780 (n11659, n_6216, n_6217);
  not g17781 (n_6218, n11657);
  and g17782 (n11660, n_6218, n11659);
  not g17783 (n_6219, n11660);
  and g17784 (n11661, n_6216, n_6219);
  not g17785 (n_6220, n11374);
  not g17786 (n_6221, n11661);
  and g17787 (n11662, n_6220, n_6221);
  not g17788 (n_6222, n11662);
  and g17789 (n11663, n_5970, n_6222);
  not g17790 (n_6223, n11356);
  not g17791 (n_6224, n11663);
  and g17792 (n11664, n_6223, n_6224);
  not g17793 (n_6225, n11664);
  and g17794 (n11665, n_5955, n_6225);
  not g17795 (n_6226, n11338);
  not g17796 (n_6227, n11665);
  and g17797 (n11666, n_6226, n_6227);
  not g17798 (n_6228, n11666);
  and g17799 (n11667, n_5940, n_6228);
  not g17800 (n_6229, n11321);
  and g17801 (n11668, n11309, n_6229);
  and g17802 (n11669, n_5928, n_6229);
  not g17803 (n_6230, n11668);
  not g17804 (n_6231, n11669);
  and g17805 (n11670, n_6230, n_6231);
  not g17806 (n_6232, n11667);
  not g17807 (n_6233, n11670);
  and g17808 (n11671, n_6232, n_6233);
  not g17809 (n_6234, n11671);
  and g17810 (n11672, n_6229, n_6234);
  not g17811 (n_6235, n11307);
  and g17812 (n11673, n11295, n_6235);
  and g17813 (n11674, n_5918, n_6235);
  not g17814 (n_6236, n11673);
  not g17815 (n_6237, n11674);
  and g17816 (n11675, n_6236, n_6237);
  not g17817 (n_6238, n11672);
  not g17818 (n_6239, n11675);
  and g17819 (n11676, n_6238, n_6239);
  not g17820 (n_6240, n11676);
  and g17821 (n11677, n_6235, n_6240);
  not g17822 (n_6241, n11281);
  and g17823 (n11678, n_6241, n11292);
  not g17824 (n_6242, n11293);
  not g17825 (n_6243, n11678);
  and g17826 (n11679, n_6242, n_6243);
  not g17827 (n_6244, n11677);
  and g17828 (n11680, n_6244, n11679);
  not g17829 (n_6245, n11680);
  and g17830 (n11681, n_6242, n_6245);
  not g17831 (n_6246, n11279);
  not g17832 (n_6247, n11681);
  and g17833 (n11682, n_6246, n_6247);
  not g17834 (n_6248, n11682);
  and g17835 (n11683, n_5896, n_6248);
  not g17836 (n_6249, n11261);
  not g17837 (n_6250, n11683);
  and g17838 (n11684, n_6249, n_6250);
  not g17839 (n_6251, n11684);
  and g17840 (n11685, n_5881, n_6251);
  not g17841 (n_6252, n11243);
  not g17842 (n_6253, n11685);
  and g17843 (n11686, n_6252, n_6253);
  not g17844 (n_6254, n11686);
  and g17845 (n11687, n_5866, n_6254);
  not g17846 (n_6255, n11226);
  and g17847 (n11688, n11214, n_6255);
  and g17848 (n11689, n_5854, n_6255);
  not g17849 (n_6256, n11688);
  not g17850 (n_6257, n11689);
  and g17851 (n11690, n_6256, n_6257);
  not g17852 (n_6258, n11687);
  not g17853 (n_6259, n11690);
  and g17854 (n11691, n_6258, n_6259);
  not g17855 (n_6260, n11691);
  and g17856 (n11692, n_6255, n_6260);
  not g17857 (n_6261, n11200);
  and g17858 (n11693, n_6261, n11211);
  not g17859 (n_6262, n11212);
  not g17860 (n_6263, n11693);
  and g17861 (n11694, n_6262, n_6263);
  not g17862 (n_6264, n11692);
  and g17863 (n11695, n_6264, n11694);
  not g17864 (n_6265, n11695);
  and g17865 (n11696, n_6262, n_6265);
  not g17866 (n_6266, n11198);
  not g17867 (n_6267, n11696);
  and g17868 (n11697, n_6266, n_6267);
  not g17869 (n_6268, n11697);
  and g17870 (n11698, n_5832, n_6268);
  not g17871 (n_6269, n11180);
  not g17872 (n_6270, n11698);
  and g17873 (n11699, n_6269, n_6270);
  not g17874 (n_6271, n11699);
  and g17875 (n11700, n_5817, n_6271);
  not g17876 (n_6272, n11162);
  not g17877 (n_6273, n11700);
  and g17878 (n11701, n_6272, n_6273);
  not g17879 (n_6274, n11701);
  and g17880 (n11702, n_5802, n_6274);
  not g17881 (n_6275, n11144);
  not g17882 (n_6276, n11702);
  and g17883 (n11703, n_6275, n_6276);
  not g17884 (n_6277, n11703);
  and g17885 (n11704, n_5787, n_6277);
  not g17886 (n_6278, n11126);
  not g17887 (n_6279, n11704);
  and g17888 (n11705, n_6278, n_6279);
  not g17889 (n_6280, n11705);
  and g17890 (n11706, n_5772, n_6280);
  not g17891 (n_6281, n11108);
  not g17892 (n_6282, n11706);
  and g17893 (n11707, n_6281, n_6282);
  not g17894 (n_6283, n11707);
  and g17895 (n11708, n_5757, n_6283);
  not g17896 (n_6284, n11090);
  not g17897 (n_6285, n11708);
  and g17898 (n11709, n_6284, n_6285);
  and g17899 (n11710, n11090, n11708);
  not g17900 (n_6286, n11709);
  not g17901 (n_6287, n11710);
  and g17902 (n11711, n_6286, n_6287);
  and g17903 (n11712, n11108, n11706);
  not g17904 (n_6288, n11712);
  and g17905 (n11713, n_6283, n_6288);
  and g17906 (n11714, n_560, n11055);
  and g17907 (n11715, n_5715, \a[1] );
  and g17908 (n11716, n_712, n11715);
  not g17909 (n_6289, n11714);
  not g17910 (n_6290, n11716);
  and g17911 (n11717, n_6289, n_6290);
  not g17912 (n_6291, n11057);
  and g17913 (n11718, n_6291, n11717);
  and g17914 (n11719, n_2152, n11717);
  not g17915 (n_6292, n11718);
  not g17916 (n_6293, n11719);
  and g17917 (n11720, n_6292, n_6293);
  not g17918 (n_6294, n11720);
  and g17919 (n11721, \a[2] , n_6294);
  and g17920 (n11722, n_10, n11720);
  not g17921 (n_6295, n11721);
  not g17922 (n_6296, n11722);
  and g17923 (n11723, n_6295, n_6296);
  not g17924 (n_6297, n11723);
  and g17925 (n11724, n11713, n_6297);
  and g17926 (n11725, n11126, n11704);
  not g17927 (n_6298, n11725);
  and g17928 (n11726, n_6280, n_6298);
  and g17929 (n11727, \a[0] , n11053);
  and g17930 (n11728, n_712, n11727);
  and g17931 (n11729, n_566, n11055);
  and g17932 (n11730, n_560, n11715);
  not g17933 (n_6299, n11729);
  not g17934 (n_6300, n11730);
  and g17935 (n11731, n_6299, n_6300);
  not g17936 (n_6301, n11728);
  and g17937 (n11732, n_6301, n11731);
  and g17938 (n11733, n_6291, n11732);
  and g17939 (n11734, n_888, n11732);
  not g17940 (n_6302, n11733);
  not g17941 (n_6303, n11734);
  and g17942 (n11735, n_6302, n_6303);
  not g17943 (n_6304, n11735);
  and g17944 (n11736, \a[2] , n_6304);
  and g17945 (n11737, n_10, n11735);
  not g17946 (n_6305, n11736);
  not g17947 (n_6306, n11737);
  and g17948 (n11738, n_6305, n_6306);
  not g17949 (n_6307, n11738);
  and g17950 (n11739, n11726, n_6307);
  and g17951 (n11740, n11144, n11702);
  not g17952 (n_6308, n11740);
  and g17953 (n11741, n_6277, n_6308);
  and g17954 (n11742, n_560, n11727);
  and g17955 (n11743, n_565, n11055);
  and g17956 (n11744, n_566, n11715);
  not g17957 (n_6309, n11743);
  not g17958 (n_6310, n11744);
  and g17959 (n11745, n_6309, n_6310);
  not g17960 (n_6311, n11742);
  and g17961 (n11746, n_6311, n11745);
  and g17962 (n11747, n_6291, n11746);
  not g17963 (n_6312, n4067);
  and g17964 (n11748, n_6312, n11746);
  not g17965 (n_6313, n11747);
  not g17966 (n_6314, n11748);
  and g17967 (n11749, n_6313, n_6314);
  not g17968 (n_6315, n11749);
  and g17969 (n11750, \a[2] , n_6315);
  and g17970 (n11751, n_10, n11749);
  not g17971 (n_6316, n11750);
  not g17972 (n_6317, n11751);
  and g17973 (n11752, n_6316, n_6317);
  not g17974 (n_6318, n11752);
  and g17975 (n11753, n11741, n_6318);
  and g17976 (n11754, n11162, n11700);
  not g17977 (n_6319, n11754);
  and g17978 (n11755, n_6274, n_6319);
  and g17979 (n11756, n_566, n11727);
  and g17980 (n11757, n_535, n11055);
  and g17981 (n11758, n_565, n11715);
  not g17982 (n_6320, n11757);
  not g17983 (n_6321, n11758);
  and g17984 (n11759, n_6320, n_6321);
  not g17985 (n_6322, n11756);
  and g17986 (n11760, n_6322, n11759);
  and g17987 (n11761, n_6291, n11760);
  not g17988 (n_6323, n4477);
  and g17989 (n11762, n_6323, n11760);
  not g17990 (n_6324, n11761);
  not g17991 (n_6325, n11762);
  and g17992 (n11763, n_6324, n_6325);
  not g17993 (n_6326, n11763);
  and g17994 (n11764, \a[2] , n_6326);
  and g17995 (n11765, n_10, n11763);
  not g17996 (n_6327, n11764);
  not g17997 (n_6328, n11765);
  and g17998 (n11766, n_6327, n_6328);
  not g17999 (n_6329, n11766);
  and g18000 (n11767, n11755, n_6329);
  and g18001 (n11768, n11180, n11698);
  not g18002 (n_6330, n11768);
  and g18003 (n11769, n_6271, n_6330);
  and g18004 (n11770, n_565, n11727);
  and g18005 (n11771, n_480, n11055);
  and g18006 (n11772, n_535, n11715);
  not g18007 (n_6331, n11771);
  not g18008 (n_6332, n11772);
  and g18009 (n11773, n_6331, n_6332);
  not g18010 (n_6333, n11770);
  and g18011 (n11774, n_6333, n11773);
  and g18012 (n11775, n_6291, n11774);
  and g18013 (n11776, n_753, n11774);
  not g18014 (n_6334, n11775);
  not g18015 (n_6335, n11776);
  and g18016 (n11777, n_6334, n_6335);
  not g18017 (n_6336, n11777);
  and g18018 (n11778, \a[2] , n_6336);
  and g18019 (n11779, n_10, n11777);
  not g18020 (n_6337, n11778);
  not g18021 (n_6338, n11779);
  and g18022 (n11780, n_6337, n_6338);
  not g18023 (n_6339, n11780);
  and g18024 (n11781, n11769, n_6339);
  not g18025 (n_6340, n11694);
  and g18026 (n11782, n11692, n_6340);
  not g18027 (n_6341, n11782);
  and g18028 (n11783, n_6265, n_6341);
  not g18029 (n_6342, n11679);
  and g18030 (n11784, n11677, n_6342);
  not g18031 (n_6343, n11784);
  and g18032 (n11785, n_6245, n_6343);
  not g18033 (n_6344, n11659);
  and g18034 (n11786, n11657, n_6344);
  not g18035 (n_6345, n11786);
  and g18036 (n11787, n_6219, n_6345);
  not g18037 (n_6346, n11639);
  and g18038 (n11788, n11637, n_6346);
  not g18039 (n_6347, n11788);
  and g18040 (n11789, n_6193, n_6347);
  not g18041 (n_6348, n11617);
  and g18042 (n11790, n11615, n_6348);
  not g18043 (n_6349, n11790);
  and g18044 (n11791, n_6166, n_6349);
  not g18045 (n_6350, n11586);
  and g18046 (n11792, n_6350, n11597);
  not g18047 (n_6351, n11598);
  not g18048 (n_6352, n11792);
  and g18049 (n11793, n_6351, n_6352);
  not g18050 (n_6353, n11727);
  and g18051 (n11794, n_6291, n_6353);
  not g18052 (n_6354, n11794);
  and g18053 (n11795, n_316, n_6354);
  and g18054 (n11796, \a[2] , n11057);
  and g18055 (n11797, n6798, n11796);
  and g18056 (n11798, n_314, n11727);
  and g18057 (n11799, n_316, n11055);
  and g18058 (n11800, n_315, n11715);
  not g18059 (n_6355, n11799);
  not g18060 (n_6356, n11800);
  and g18061 (n11801, n_6355, n_6356);
  not g18062 (n_6357, n11798);
  and g18063 (n11802, n_6357, n11801);
  not g18064 (n_6358, n11802);
  and g18065 (n11803, \a[2] , n_6358);
  and g18066 (n11804, n_2588, n11796);
  and g18067 (n11805, \a[2] , n11715);
  and g18068 (n11806, n_316, n11805);
  and g18069 (n11807, \a[2] , n11727);
  and g18070 (n11808, n_315, n11807);
  and g18083 (n11815, n11584, n11814);
  not g18084 (n_6365, n11814);
  and g18085 (n11816, n_6137, n_6365);
  and g18086 (n11817, n_313, n11727);
  and g18087 (n11818, n_315, n11055);
  and g18088 (n11819, n_314, n11715);
  and g18094 (n11822, n6806, n11057);
  not g18097 (n_6370, n11823);
  and g18098 (n11824, n_10, n_6370);
  and g18099 (n11825, \a[2] , n11823);
  not g18100 (n_6371, n11824);
  not g18101 (n_6372, n11825);
  and g18102 (n11826, n_6371, n_6372);
  not g18103 (n_6373, n11816);
  not g18104 (n_6374, n11826);
  and g18105 (n11827, n_6373, n_6374);
  not g18106 (n_6375, n11815);
  not g18107 (n_6376, n11827);
  and g18108 (n11828, n_6375, n_6376);
  and g18109 (n11829, n_312, n11727);
  and g18110 (n11830, n_314, n11055);
  and g18111 (n11831, n_313, n11715);
  not g18112 (n_6377, n11830);
  not g18113 (n_6378, n11831);
  and g18114 (n11832, n_6377, n_6378);
  not g18115 (n_6379, n11829);
  and g18116 (n11833, n_6379, n11832);
  and g18117 (n11834, n_6291, n11833);
  and g18118 (n11835, n_2891, n11833);
  not g18119 (n_6380, n11834);
  not g18120 (n_6381, n11835);
  and g18121 (n11836, n_6380, n_6381);
  not g18122 (n_6382, n11836);
  and g18123 (n11837, \a[2] , n_6382);
  and g18124 (n11838, n_10, n11836);
  not g18125 (n_6383, n11837);
  not g18126 (n_6384, n11838);
  and g18127 (n11839, n_6383, n_6384);
  and g18128 (n11840, n11828, n11839);
  not g18129 (n_6385, n11585);
  and g18130 (n11841, n11583, n_6385);
  not g18131 (n_6386, n11841);
  and g18132 (n11842, n_6350, n_6386);
  not g18133 (n_6387, n11840);
  and g18134 (n11843, n_6387, n11842);
  not g18135 (n_6388, n11828);
  not g18136 (n_6389, n11839);
  and g18137 (n11844, n_6388, n_6389);
  not g18138 (n_6390, n11843);
  not g18139 (n_6391, n11844);
  and g18140 (n11845, n_6390, n_6391);
  not g18141 (n_6392, n11845);
  and g18142 (n11846, n11793, n_6392);
  not g18143 (n_6393, n11793);
  and g18144 (n11847, n_6393, n11845);
  and g18145 (n11848, n_311, n11727);
  and g18146 (n11849, n_313, n11055);
  and g18147 (n11850, n_312, n11715);
  and g18153 (n11853, n6646, n11057);
  not g18156 (n_6398, n11854);
  and g18157 (n11855, n_10, n_6398);
  and g18158 (n11856, \a[2] , n11854);
  not g18159 (n_6399, n11855);
  not g18160 (n_6400, n11856);
  and g18161 (n11857, n_6399, n_6400);
  not g18162 (n_6401, n11847);
  not g18163 (n_6402, n11857);
  and g18164 (n11858, n_6401, n_6402);
  not g18165 (n_6403, n11846);
  not g18166 (n_6404, n11858);
  and g18167 (n11859, n_6403, n_6404);
  and g18168 (n11860, n_310, n11727);
  and g18169 (n11861, n_312, n11055);
  and g18170 (n11862, n_311, n11715);
  not g18171 (n_6405, n11861);
  not g18172 (n_6406, n11862);
  and g18173 (n11863, n_6405, n_6406);
  not g18174 (n_6407, n11860);
  and g18175 (n11864, n_6407, n11863);
  and g18176 (n11865, n_6291, n11864);
  and g18177 (n11866, n_3239, n11864);
  not g18178 (n_6408, n11865);
  not g18179 (n_6409, n11866);
  and g18180 (n11867, n_6408, n_6409);
  not g18181 (n_6410, n11867);
  and g18182 (n11868, \a[2] , n_6410);
  and g18183 (n11869, n_10, n11867);
  not g18184 (n_6411, n11868);
  not g18185 (n_6412, n11869);
  and g18186 (n11870, n_6411, n_6412);
  not g18187 (n_6413, n11859);
  not g18188 (n_6414, n11870);
  and g18189 (n11871, n_6413, n_6414);
  and g18190 (n11872, n11859, n11870);
  and g18191 (n11873, n11602, n11613);
  not g18192 (n_6415, n11873);
  and g18193 (n11874, n_6161, n_6415);
  not g18194 (n_6416, n11872);
  and g18195 (n11875, n_6416, n11874);
  not g18196 (n_6417, n11871);
  not g18197 (n_6418, n11875);
  and g18198 (n11876, n_6417, n_6418);
  not g18199 (n_6419, n11876);
  and g18200 (n11877, n11791, n_6419);
  not g18201 (n_6420, n11791);
  and g18202 (n11878, n_6420, n11876);
  and g18203 (n11879, n_309, n11727);
  and g18204 (n11880, n_311, n11055);
  and g18205 (n11881, n_310, n11715);
  and g18211 (n11884, n6541, n11057);
  not g18214 (n_6425, n11885);
  and g18215 (n11886, n_10, n_6425);
  and g18216 (n11887, \a[2] , n11885);
  not g18217 (n_6426, n11886);
  not g18218 (n_6427, n11887);
  and g18219 (n11888, n_6426, n_6427);
  not g18220 (n_6428, n11878);
  not g18221 (n_6429, n11888);
  and g18222 (n11889, n_6428, n_6429);
  not g18223 (n_6430, n11877);
  not g18224 (n_6431, n11889);
  and g18225 (n11890, n_6430, n_6431);
  and g18226 (n11891, n_308, n11727);
  and g18227 (n11892, n_310, n11055);
  and g18228 (n11893, n_309, n11715);
  not g18229 (n_6432, n11892);
  not g18230 (n_6433, n11893);
  and g18231 (n11894, n_6432, n_6433);
  not g18232 (n_6434, n11891);
  and g18233 (n11895, n_6434, n11894);
  and g18234 (n11896, n_6291, n11895);
  and g18235 (n11897, n_2839, n11895);
  not g18236 (n_6435, n11896);
  not g18237 (n_6436, n11897);
  and g18238 (n11898, n_6435, n_6436);
  not g18239 (n_6437, n11898);
  and g18240 (n11899, \a[2] , n_6437);
  and g18241 (n11900, n_10, n11898);
  not g18242 (n_6438, n11899);
  not g18243 (n_6439, n11900);
  and g18244 (n11901, n_6438, n_6439);
  and g18245 (n11902, n11890, n11901);
  and g18246 (n11903, n11560, n11619);
  not g18247 (n_6440, n11903);
  and g18248 (n11904, n_6169, n_6440);
  not g18249 (n_6441, n11902);
  and g18250 (n11905, n_6441, n11904);
  not g18251 (n_6442, n11890);
  not g18252 (n_6443, n11901);
  and g18253 (n11906, n_6442, n_6443);
  not g18254 (n_6444, n11905);
  not g18255 (n_6445, n11906);
  and g18256 (n11907, n_6444, n_6445);
  and g18257 (n11908, n_307, n11727);
  and g18258 (n11909, n_309, n11055);
  and g18259 (n11910, n_308, n11715);
  not g18260 (n_6446, n11909);
  not g18261 (n_6447, n11910);
  and g18262 (n11911, n_6446, n_6447);
  not g18263 (n_6448, n11908);
  and g18264 (n11912, n_6448, n11911);
  and g18265 (n11913, n_6291, n11912);
  and g18266 (n11914, n_2511, n11912);
  not g18267 (n_6449, n11913);
  not g18268 (n_6450, n11914);
  and g18269 (n11915, n_6449, n_6450);
  not g18270 (n_6451, n11915);
  and g18271 (n11916, \a[2] , n_6451);
  and g18272 (n11917, n_10, n11915);
  not g18273 (n_6452, n11916);
  not g18274 (n_6453, n11917);
  and g18275 (n11918, n_6452, n_6453);
  and g18276 (n11919, n11907, n11918);
  not g18277 (n_6454, n11623);
  and g18278 (n11920, n11621, n_6454);
  not g18279 (n_6455, n11920);
  and g18280 (n11921, n_6173, n_6455);
  not g18281 (n_6456, n11919);
  and g18282 (n11922, n_6456, n11921);
  not g18283 (n_6457, n11907);
  not g18284 (n_6458, n11918);
  and g18285 (n11923, n_6457, n_6458);
  not g18286 (n_6459, n11922);
  not g18287 (n_6460, n11923);
  and g18288 (n11924, n_6459, n_6460);
  and g18289 (n11925, n_306, n11727);
  and g18290 (n11926, n_308, n11055);
  and g18291 (n11927, n_307, n11715);
  not g18292 (n_6461, n11926);
  not g18293 (n_6462, n11927);
  and g18294 (n11928, n_6461, n_6462);
  not g18295 (n_6463, n11925);
  and g18296 (n11929, n_6463, n11928);
  and g18297 (n11930, n_6291, n11929);
  and g18298 (n11931, n_2498, n11929);
  not g18299 (n_6464, n11930);
  not g18300 (n_6465, n11931);
  and g18301 (n11932, n_6464, n_6465);
  not g18302 (n_6466, n11932);
  and g18303 (n11933, \a[2] , n_6466);
  and g18304 (n11934, n_10, n11932);
  not g18305 (n_6467, n11933);
  not g18306 (n_6468, n11934);
  and g18307 (n11935, n_6467, n_6468);
  and g18308 (n11936, n11924, n11935);
  and g18309 (n11937, n11528, n11625);
  not g18310 (n_6469, n11937);
  and g18311 (n11938, n_6176, n_6469);
  not g18312 (n_6470, n11936);
  and g18313 (n11939, n_6470, n11938);
  not g18314 (n_6471, n11924);
  not g18315 (n_6472, n11935);
  and g18316 (n11940, n_6471, n_6472);
  not g18317 (n_6473, n11939);
  not g18318 (n_6474, n11940);
  and g18319 (n11941, n_6473, n_6474);
  and g18320 (n11942, n11627, n_6179);
  and g18321 (n11943, n_6178, n11942);
  not g18322 (n_6475, n11943);
  and g18323 (n11944, n_6182, n_6475);
  not g18324 (n_6476, n11941);
  and g18325 (n11945, n_6476, n11944);
  not g18326 (n_6477, n11944);
  and g18327 (n11946, n11941, n_6477);
  and g18328 (n11947, n_305, n11727);
  and g18329 (n11948, n_307, n11055);
  and g18330 (n11949, n_306, n11715);
  and g18336 (n11952, n6143, n11057);
  not g18339 (n_6482, n11953);
  and g18340 (n11954, n_10, n_6482);
  and g18341 (n11955, \a[2] , n11953);
  not g18342 (n_6483, n11954);
  not g18343 (n_6484, n11955);
  and g18344 (n11956, n_6483, n_6484);
  not g18345 (n_6485, n11946);
  not g18346 (n_6486, n11956);
  and g18347 (n11957, n_6485, n_6486);
  not g18348 (n_6487, n11945);
  not g18349 (n_6488, n11957);
  and g18350 (n11958, n_6487, n_6488);
  and g18351 (n11959, n11632, n_6185);
  and g18352 (n11960, n_6184, n11959);
  not g18353 (n_6489, n11960);
  and g18354 (n11961, n_6188, n_6489);
  not g18355 (n_6490, n11958);
  and g18356 (n11962, n_6490, n11961);
  not g18357 (n_6491, n11961);
  and g18358 (n11963, n11958, n_6491);
  and g18359 (n11964, n_304, n11727);
  and g18360 (n11965, n_306, n11055);
  and g18361 (n11966, n_305, n11715);
  and g18367 (n11969, n5834, n11057);
  not g18370 (n_6496, n11970);
  and g18371 (n11971, n_10, n_6496);
  and g18372 (n11972, \a[2] , n11970);
  not g18373 (n_6497, n11971);
  not g18374 (n_6498, n11972);
  and g18375 (n11973, n_6497, n_6498);
  not g18376 (n_6499, n11963);
  not g18377 (n_6500, n11973);
  and g18378 (n11974, n_6499, n_6500);
  not g18379 (n_6501, n11962);
  not g18380 (n_6502, n11974);
  and g18381 (n11975, n_6501, n_6502);
  not g18382 (n_6503, n11975);
  and g18383 (n11976, n11789, n_6503);
  not g18384 (n_6504, n11789);
  and g18385 (n11977, n_6504, n11975);
  and g18386 (n11978, n_303, n11727);
  and g18387 (n11979, n_305, n11055);
  and g18388 (n11980, n_304, n11715);
  and g18394 (n11983, n6007, n11057);
  not g18397 (n_6509, n11984);
  and g18398 (n11985, n_10, n_6509);
  and g18399 (n11986, \a[2] , n11984);
  not g18400 (n_6510, n11985);
  not g18401 (n_6511, n11986);
  and g18402 (n11987, n_6510, n_6511);
  not g18403 (n_6512, n11977);
  not g18404 (n_6513, n11987);
  and g18405 (n11988, n_6512, n_6513);
  not g18406 (n_6514, n11976);
  not g18407 (n_6515, n11988);
  and g18408 (n11989, n_6514, n_6515);
  and g18409 (n11990, n_302, n11727);
  and g18410 (n11991, n_304, n11055);
  and g18411 (n11992, n_303, n11715);
  not g18412 (n_6516, n11991);
  not g18413 (n_6517, n11992);
  and g18414 (n11993, n_6516, n_6517);
  not g18415 (n_6518, n11990);
  and g18416 (n11994, n_6518, n11993);
  and g18417 (n11995, n_6291, n11994);
  and g18418 (n11996, n_3507, n11994);
  not g18419 (n_6519, n11995);
  not g18420 (n_6520, n11996);
  and g18421 (n11997, n_6519, n_6520);
  not g18422 (n_6521, n11997);
  and g18423 (n11998, \a[2] , n_6521);
  and g18424 (n11999, n_10, n11997);
  not g18425 (n_6522, n11998);
  not g18426 (n_6523, n11999);
  and g18427 (n12000, n_6522, n_6523);
  and g18428 (n12001, n11989, n12000);
  and g18429 (n12002, n11469, n11641);
  not g18430 (n_6524, n12002);
  and g18431 (n12003, n_6196, n_6524);
  not g18432 (n_6525, n12001);
  and g18433 (n12004, n_6525, n12003);
  not g18434 (n_6526, n11989);
  not g18435 (n_6527, n12000);
  and g18436 (n12005, n_6526, n_6527);
  not g18437 (n_6528, n12004);
  not g18438 (n_6529, n12005);
  and g18439 (n12006, n_6528, n_6529);
  and g18440 (n12007, n_301, n11727);
  and g18441 (n12008, n_303, n11055);
  and g18442 (n12009, n_302, n11715);
  not g18443 (n_6530, n12008);
  not g18444 (n_6531, n12009);
  and g18445 (n12010, n_6530, n_6531);
  not g18446 (n_6532, n12007);
  and g18447 (n12011, n_6532, n12010);
  and g18448 (n12012, n_6291, n12011);
  and g18449 (n12013, n_1672, n12011);
  not g18450 (n_6533, n12012);
  not g18451 (n_6534, n12013);
  and g18452 (n12014, n_6533, n_6534);
  not g18453 (n_6535, n12014);
  and g18454 (n12015, \a[2] , n_6535);
  and g18455 (n12016, n_10, n12014);
  not g18456 (n_6536, n12015);
  not g18457 (n_6537, n12016);
  and g18458 (n12017, n_6536, n_6537);
  and g18459 (n12018, n12006, n12017);
  and g18460 (n12019, n11451, n11643);
  not g18461 (n_6538, n12019);
  and g18462 (n12020, n_6199, n_6538);
  not g18463 (n_6539, n12018);
  and g18464 (n12021, n_6539, n12020);
  not g18465 (n_6540, n12006);
  not g18466 (n_6541, n12017);
  and g18467 (n12022, n_6540, n_6541);
  not g18468 (n_6542, n12021);
  not g18469 (n_6543, n12022);
  and g18470 (n12023, n_6542, n_6543);
  and g18471 (n12024, n_300, n11727);
  and g18472 (n12025, n_302, n11055);
  and g18473 (n12026, n_301, n11715);
  not g18474 (n_6544, n12025);
  not g18475 (n_6545, n12026);
  and g18476 (n12027, n_6544, n_6545);
  not g18477 (n_6546, n12024);
  and g18478 (n12028, n_6546, n12027);
  and g18479 (n12029, n_6291, n12028);
  and g18480 (n12030, n_1801, n12028);
  not g18481 (n_6547, n12029);
  not g18482 (n_6548, n12030);
  and g18483 (n12031, n_6547, n_6548);
  not g18484 (n_6549, n12031);
  and g18485 (n12032, \a[2] , n_6549);
  and g18486 (n12033, n_10, n12031);
  not g18487 (n_6550, n12032);
  not g18488 (n_6551, n12033);
  and g18489 (n12034, n_6550, n_6551);
  and g18490 (n12035, n12023, n12034);
  and g18491 (n12036, n11433, n11645);
  not g18492 (n_6552, n12036);
  and g18493 (n12037, n_6202, n_6552);
  not g18494 (n_6553, n12035);
  and g18495 (n12038, n_6553, n12037);
  not g18496 (n_6554, n12023);
  not g18497 (n_6555, n12034);
  and g18498 (n12039, n_6554, n_6555);
  not g18499 (n_6556, n12038);
  not g18500 (n_6557, n12039);
  and g18501 (n12040, n_6556, n_6557);
  and g18502 (n12041, n11647, n_6205);
  and g18503 (n12042, n_6204, n12041);
  not g18504 (n_6558, n12042);
  and g18505 (n12043, n_6208, n_6558);
  not g18506 (n_6559, n12040);
  and g18507 (n12044, n_6559, n12043);
  not g18508 (n_6560, n12043);
  and g18509 (n12045, n12040, n_6560);
  and g18510 (n12046, n_299, n11727);
  and g18511 (n12047, n_301, n11055);
  and g18512 (n12048, n_300, n11715);
  and g18518 (n12051, n5139, n11057);
  not g18521 (n_6565, n12052);
  and g18522 (n12053, n_10, n_6565);
  and g18523 (n12054, \a[2] , n12052);
  not g18524 (n_6566, n12053);
  not g18525 (n_6567, n12054);
  and g18526 (n12055, n_6566, n_6567);
  not g18527 (n_6568, n12045);
  not g18528 (n_6569, n12055);
  and g18529 (n12056, n_6568, n_6569);
  not g18530 (n_6570, n12044);
  not g18531 (n_6571, n12056);
  and g18532 (n12057, n_6570, n_6571);
  and g18533 (n12058, n11652, n_6211);
  and g18534 (n12059, n_6210, n12058);
  not g18535 (n_6572, n12059);
  and g18536 (n12060, n_6214, n_6572);
  not g18537 (n_6573, n12057);
  and g18538 (n12061, n_6573, n12060);
  not g18539 (n_6574, n12060);
  and g18540 (n12062, n12057, n_6574);
  and g18541 (n12063, n_298, n11727);
  and g18542 (n12064, n_300, n11055);
  and g18543 (n12065, n_299, n11715);
  and g18549 (n12068, n5114, n11057);
  not g18552 (n_6579, n12069);
  and g18553 (n12070, n_10, n_6579);
  and g18554 (n12071, \a[2] , n12069);
  not g18555 (n_6580, n12070);
  not g18556 (n_6581, n12071);
  and g18557 (n12072, n_6580, n_6581);
  not g18558 (n_6582, n12062);
  not g18559 (n_6583, n12072);
  and g18560 (n12073, n_6582, n_6583);
  not g18561 (n_6584, n12061);
  not g18562 (n_6585, n12073);
  and g18563 (n12074, n_6584, n_6585);
  not g18564 (n_6586, n12074);
  and g18565 (n12075, n11787, n_6586);
  not g18566 (n_6587, n11787);
  and g18567 (n12076, n_6587, n12074);
  and g18568 (n12077, n_295, n11727);
  and g18569 (n12078, n_299, n11055);
  and g18570 (n12079, n_298, n11715);
  and g18576 (n12082, n4848, n11057);
  not g18579 (n_6592, n12083);
  and g18580 (n12084, n_10, n_6592);
  and g18581 (n12085, \a[2] , n12083);
  not g18582 (n_6593, n12084);
  not g18583 (n_6594, n12085);
  and g18584 (n12086, n_6593, n_6594);
  not g18585 (n_6595, n12076);
  not g18586 (n_6596, n12086);
  and g18587 (n12087, n_6595, n_6596);
  not g18588 (n_6597, n12075);
  not g18589 (n_6598, n12087);
  and g18590 (n12088, n_6597, n_6598);
  and g18591 (n12089, n_293, n11727);
  and g18592 (n12090, n_298, n11055);
  and g18593 (n12091, n_295, n11715);
  not g18594 (n_6599, n12090);
  not g18595 (n_6600, n12091);
  and g18596 (n12092, n_6599, n_6600);
  not g18597 (n_6601, n12089);
  and g18598 (n12093, n_6601, n12092);
  and g18599 (n12094, n_6291, n12093);
  and g18600 (n12095, n_1789, n12093);
  not g18601 (n_6602, n12094);
  not g18602 (n_6603, n12095);
  and g18603 (n12096, n_6602, n_6603);
  not g18604 (n_6604, n12096);
  and g18605 (n12097, \a[2] , n_6604);
  and g18606 (n12098, n_10, n12096);
  not g18607 (n_6605, n12097);
  not g18608 (n_6606, n12098);
  and g18609 (n12099, n_6605, n_6606);
  and g18610 (n12100, n12088, n12099);
  and g18611 (n12101, n11374, n11661);
  not g18612 (n_6607, n12101);
  and g18613 (n12102, n_6222, n_6607);
  not g18614 (n_6608, n12100);
  and g18615 (n12103, n_6608, n12102);
  not g18616 (n_6609, n12088);
  not g18617 (n_6610, n12099);
  and g18618 (n12104, n_6609, n_6610);
  not g18619 (n_6611, n12103);
  not g18620 (n_6612, n12104);
  and g18621 (n12105, n_6611, n_6612);
  and g18622 (n12106, n_286, n11727);
  and g18623 (n12107, n_295, n11055);
  and g18624 (n12108, n_293, n11715);
  not g18625 (n_6613, n12107);
  not g18626 (n_6614, n12108);
  and g18627 (n12109, n_6613, n_6614);
  not g18628 (n_6615, n12106);
  and g18629 (n12110, n_6615, n12109);
  and g18630 (n12111, n_6291, n12110);
  and g18631 (n12112, n_1134, n12110);
  not g18632 (n_6616, n12111);
  not g18633 (n_6617, n12112);
  and g18634 (n12113, n_6616, n_6617);
  not g18635 (n_6618, n12113);
  and g18636 (n12114, \a[2] , n_6618);
  and g18637 (n12115, n_10, n12113);
  not g18638 (n_6619, n12114);
  not g18639 (n_6620, n12115);
  and g18640 (n12116, n_6619, n_6620);
  and g18641 (n12117, n12105, n12116);
  and g18642 (n12118, n11356, n11663);
  not g18643 (n_6621, n12118);
  and g18644 (n12119, n_6225, n_6621);
  not g18645 (n_6622, n12117);
  and g18646 (n12120, n_6622, n12119);
  not g18647 (n_6623, n12105);
  not g18648 (n_6624, n12116);
  and g18649 (n12121, n_6623, n_6624);
  not g18650 (n_6625, n12120);
  not g18651 (n_6626, n12121);
  and g18652 (n12122, n_6625, n_6626);
  and g18653 (n12123, n_281, n11727);
  and g18654 (n12124, n_293, n11055);
  and g18655 (n12125, n_286, n11715);
  not g18656 (n_6627, n12124);
  not g18657 (n_6628, n12125);
  and g18658 (n12126, n_6627, n_6628);
  not g18659 (n_6629, n12123);
  and g18660 (n12127, n_6629, n12126);
  and g18661 (n12128, n_6291, n12127);
  and g18662 (n12129, n_1228, n12127);
  not g18663 (n_6630, n12128);
  not g18664 (n_6631, n12129);
  and g18665 (n12130, n_6630, n_6631);
  not g18666 (n_6632, n12130);
  and g18667 (n12131, \a[2] , n_6632);
  and g18668 (n12132, n_10, n12130);
  not g18669 (n_6633, n12131);
  not g18670 (n_6634, n12132);
  and g18671 (n12133, n_6633, n_6634);
  and g18672 (n12134, n12122, n12133);
  and g18673 (n12135, n11338, n11665);
  not g18674 (n_6635, n12135);
  and g18675 (n12136, n_6228, n_6635);
  not g18676 (n_6636, n12134);
  and g18677 (n12137, n_6636, n12136);
  not g18678 (n_6637, n12122);
  not g18679 (n_6638, n12133);
  and g18680 (n12138, n_6637, n_6638);
  not g18681 (n_6639, n12137);
  not g18682 (n_6640, n12138);
  and g18683 (n12139, n_6639, n_6640);
  and g18684 (n12140, n11667, n_6231);
  and g18685 (n12141, n_6230, n12140);
  not g18686 (n_6641, n12141);
  and g18687 (n12142, n_6234, n_6641);
  not g18688 (n_6642, n12139);
  and g18689 (n12143, n_6642, n12142);
  not g18690 (n_6643, n12142);
  and g18691 (n12144, n12139, n_6643);
  and g18692 (n12145, n_275, n11727);
  and g18693 (n12146, n_286, n11055);
  and g18694 (n12147, n_281, n11715);
  and g18700 (n12150, n4204, n11057);
  not g18703 (n_6648, n12151);
  and g18704 (n12152, n_10, n_6648);
  and g18705 (n12153, \a[2] , n12151);
  not g18706 (n_6649, n12152);
  not g18707 (n_6650, n12153);
  and g18708 (n12154, n_6649, n_6650);
  not g18709 (n_6651, n12144);
  not g18710 (n_6652, n12154);
  and g18711 (n12155, n_6651, n_6652);
  not g18712 (n_6653, n12143);
  not g18713 (n_6654, n12155);
  and g18714 (n12156, n_6653, n_6654);
  and g18715 (n12157, n11672, n_6237);
  and g18716 (n12158, n_6236, n12157);
  not g18717 (n_6655, n12158);
  and g18718 (n12159, n_6240, n_6655);
  not g18719 (n_6656, n12156);
  and g18720 (n12160, n_6656, n12159);
  not g18721 (n_6657, n12159);
  and g18722 (n12161, n12156, n_6657);
  and g18723 (n12162, n_260, n11727);
  and g18724 (n12163, n_281, n11055);
  and g18725 (n12164, n_275, n11715);
  and g18731 (n12167, n4179, n11057);
  not g18734 (n_6662, n12168);
  and g18735 (n12169, n_10, n_6662);
  and g18736 (n12170, \a[2] , n12168);
  not g18737 (n_6663, n12169);
  not g18738 (n_6664, n12170);
  and g18739 (n12171, n_6663, n_6664);
  not g18740 (n_6665, n12161);
  not g18741 (n_6666, n12171);
  and g18742 (n12172, n_6665, n_6666);
  not g18743 (n_6667, n12160);
  not g18744 (n_6668, n12172);
  and g18745 (n12173, n_6667, n_6668);
  not g18746 (n_6669, n12173);
  and g18747 (n12174, n11785, n_6669);
  not g18748 (n_6670, n11785);
  and g18749 (n12175, n_6670, n12173);
  and g18750 (n12176, n_237, n11727);
  and g18751 (n12177, n_275, n11055);
  and g18752 (n12178, n_260, n11715);
  and g18758 (n12181, n3331, n11057);
  not g18761 (n_6675, n12182);
  and g18762 (n12183, n_10, n_6675);
  and g18763 (n12184, \a[2] , n12182);
  not g18764 (n_6676, n12183);
  not g18765 (n_6677, n12184);
  and g18766 (n12185, n_6676, n_6677);
  not g18767 (n_6678, n12175);
  not g18768 (n_6679, n12185);
  and g18769 (n12186, n_6678, n_6679);
  not g18770 (n_6680, n12174);
  not g18771 (n_6681, n12186);
  and g18772 (n12187, n_6680, n_6681);
  and g18773 (n12188, n_236, n11727);
  and g18774 (n12189, n_260, n11055);
  and g18775 (n12190, n_237, n11715);
  not g18776 (n_6682, n12189);
  not g18777 (n_6683, n12190);
  and g18778 (n12191, n_6682, n_6683);
  not g18779 (n_6684, n12188);
  and g18780 (n12192, n_6684, n12191);
  and g18781 (n12193, n_6291, n12192);
  and g18782 (n12194, n_1208, n12192);
  not g18783 (n_6685, n12193);
  not g18784 (n_6686, n12194);
  and g18785 (n12195, n_6685, n_6686);
  not g18786 (n_6687, n12195);
  and g18787 (n12196, \a[2] , n_6687);
  and g18788 (n12197, n_10, n12195);
  not g18789 (n_6688, n12196);
  not g18790 (n_6689, n12197);
  and g18791 (n12198, n_6688, n_6689);
  and g18792 (n12199, n12187, n12198);
  and g18793 (n12200, n11279, n11681);
  not g18794 (n_6690, n12200);
  and g18795 (n12201, n_6248, n_6690);
  not g18796 (n_6691, n12199);
  and g18797 (n12202, n_6691, n12201);
  not g18798 (n_6692, n12187);
  not g18799 (n_6693, n12198);
  and g18800 (n12203, n_6692, n_6693);
  not g18801 (n_6694, n12202);
  not g18802 (n_6695, n12203);
  and g18803 (n12204, n_6694, n_6695);
  and g18804 (n12205, n_415, n11727);
  and g18805 (n12206, n_237, n11055);
  and g18806 (n12207, n_236, n11715);
  not g18807 (n_6696, n12206);
  not g18808 (n_6697, n12207);
  and g18809 (n12208, n_6696, n_6697);
  not g18810 (n_6698, n12205);
  and g18811 (n12209, n_6698, n12208);
  and g18812 (n12210, n_6291, n12209);
  and g18813 (n12211, n_680, n12209);
  not g18814 (n_6699, n12210);
  not g18815 (n_6700, n12211);
  and g18816 (n12212, n_6699, n_6700);
  not g18817 (n_6701, n12212);
  and g18818 (n12213, \a[2] , n_6701);
  and g18819 (n12214, n_10, n12212);
  not g18820 (n_6702, n12213);
  not g18821 (n_6703, n12214);
  and g18822 (n12215, n_6702, n_6703);
  and g18823 (n12216, n12204, n12215);
  and g18824 (n12217, n11261, n11683);
  not g18825 (n_6704, n12217);
  and g18826 (n12218, n_6251, n_6704);
  not g18827 (n_6705, n12216);
  and g18828 (n12219, n_6705, n12218);
  not g18829 (n_6706, n12204);
  not g18830 (n_6707, n12215);
  and g18831 (n12220, n_6706, n_6707);
  not g18832 (n_6708, n12219);
  not g18833 (n_6709, n12220);
  and g18834 (n12221, n_6708, n_6709);
  and g18835 (n12222, n_484, n11727);
  and g18836 (n12223, n_236, n11055);
  and g18837 (n12224, n_415, n11715);
  not g18838 (n_6710, n12223);
  not g18839 (n_6711, n12224);
  and g18840 (n12225, n_6710, n_6711);
  not g18841 (n_6712, n12222);
  and g18842 (n12226, n_6712, n12225);
  and g18843 (n12227, n_6291, n12226);
  and g18844 (n12228, n_773, n12226);
  not g18845 (n_6713, n12227);
  not g18846 (n_6714, n12228);
  and g18847 (n12229, n_6713, n_6714);
  not g18848 (n_6715, n12229);
  and g18849 (n12230, \a[2] , n_6715);
  and g18850 (n12231, n_10, n12229);
  not g18851 (n_6716, n12230);
  not g18852 (n_6717, n12231);
  and g18853 (n12232, n_6716, n_6717);
  and g18854 (n12233, n12221, n12232);
  and g18855 (n12234, n11243, n11685);
  not g18856 (n_6718, n12234);
  and g18857 (n12235, n_6254, n_6718);
  not g18858 (n_6719, n12233);
  and g18859 (n12236, n_6719, n12235);
  not g18860 (n_6720, n12221);
  not g18861 (n_6721, n12232);
  and g18862 (n12237, n_6720, n_6721);
  not g18863 (n_6722, n12236);
  not g18864 (n_6723, n12237);
  and g18865 (n12238, n_6722, n_6723);
  and g18866 (n12239, n11687, n_6257);
  and g18867 (n12240, n_6256, n12239);
  not g18868 (n_6724, n12240);
  and g18869 (n12241, n_6260, n_6724);
  not g18870 (n_6725, n12238);
  and g18871 (n12242, n_6725, n12241);
  not g18872 (n_6726, n12241);
  and g18873 (n12243, n12238, n_6726);
  and g18874 (n12244, n_485, n11727);
  and g18875 (n12245, n_415, n11055);
  and g18876 (n12246, n_484, n11715);
  and g18882 (n12249, n4084, n11057);
  not g18885 (n_6731, n12250);
  and g18886 (n12251, n_10, n_6731);
  and g18887 (n12252, \a[2] , n12250);
  not g18888 (n_6732, n12251);
  not g18889 (n_6733, n12252);
  and g18890 (n12253, n_6732, n_6733);
  not g18891 (n_6734, n12243);
  not g18892 (n_6735, n12253);
  and g18893 (n12254, n_6734, n_6735);
  not g18894 (n_6736, n12242);
  not g18895 (n_6737, n12254);
  and g18896 (n12255, n_6736, n_6737);
  not g18897 (n_6738, n12255);
  and g18898 (n12256, n11783, n_6738);
  not g18899 (n_6739, n11783);
  and g18900 (n12257, n_6739, n12255);
  and g18901 (n12258, n_480, n11727);
  and g18902 (n12259, n_484, n11055);
  and g18903 (n12260, n_485, n11715);
  and g18909 (n12263, n3627, n11057);
  not g18912 (n_6744, n12264);
  and g18913 (n12265, n_10, n_6744);
  and g18914 (n12266, \a[2] , n12264);
  not g18915 (n_6745, n12265);
  not g18916 (n_6746, n12266);
  and g18917 (n12267, n_6745, n_6746);
  not g18918 (n_6747, n12257);
  not g18919 (n_6748, n12267);
  and g18920 (n12268, n_6747, n_6748);
  not g18921 (n_6749, n12256);
  not g18922 (n_6750, n12268);
  and g18923 (n12269, n_6749, n_6750);
  and g18924 (n12270, n_535, n11727);
  and g18925 (n12271, n_485, n11055);
  and g18926 (n12272, n_480, n11715);
  not g18927 (n_6751, n12271);
  not g18928 (n_6752, n12272);
  and g18929 (n12273, n_6751, n_6752);
  not g18930 (n_6753, n12270);
  and g18931 (n12274, n_6753, n12273);
  and g18932 (n12275, n_6291, n12274);
  and g18933 (n12276, n_545, n12274);
  not g18934 (n_6754, n12275);
  not g18935 (n_6755, n12276);
  and g18936 (n12277, n_6754, n_6755);
  not g18937 (n_6756, n12277);
  and g18938 (n12278, \a[2] , n_6756);
  and g18939 (n12279, n_10, n12277);
  not g18940 (n_6757, n12278);
  not g18941 (n_6758, n12279);
  and g18942 (n12280, n_6757, n_6758);
  and g18943 (n12281, n12269, n12280);
  and g18944 (n12282, n11198, n11696);
  not g18945 (n_6759, n12282);
  and g18946 (n12283, n_6268, n_6759);
  not g18947 (n_6760, n12281);
  and g18948 (n12284, n_6760, n12283);
  not g18949 (n_6761, n12269);
  not g18950 (n_6762, n12280);
  and g18951 (n12285, n_6761, n_6762);
  not g18952 (n_6763, n12284);
  not g18953 (n_6764, n12285);
  and g18954 (n12286, n_6763, n_6764);
  not g18955 (n_6765, n11781);
  and g18956 (n12287, n11769, n_6765);
  and g18957 (n12288, n_6339, n_6765);
  not g18958 (n_6766, n12287);
  not g18959 (n_6767, n12288);
  and g18960 (n12289, n_6766, n_6767);
  not g18961 (n_6768, n12286);
  not g18962 (n_6769, n12289);
  and g18963 (n12290, n_6768, n_6769);
  not g18964 (n_6770, n12290);
  and g18965 (n12291, n_6765, n_6770);
  not g18966 (n_6771, n11755);
  and g18967 (n12292, n_6771, n11766);
  not g18968 (n_6772, n11767);
  not g18969 (n_6773, n12292);
  and g18970 (n12293, n_6772, n_6773);
  not g18971 (n_6774, n12291);
  and g18972 (n12294, n_6774, n12293);
  not g18973 (n_6775, n12294);
  and g18974 (n12295, n_6772, n_6775);
  not g18975 (n_6776, n11741);
  and g18976 (n12296, n_6776, n11752);
  not g18977 (n_6777, n11753);
  not g18978 (n_6778, n12296);
  and g18979 (n12297, n_6777, n_6778);
  not g18980 (n_6779, n12295);
  and g18981 (n12298, n_6779, n12297);
  not g18982 (n_6780, n12298);
  and g18983 (n12299, n_6777, n_6780);
  not g18984 (n_6781, n11726);
  and g18985 (n12300, n_6781, n11738);
  not g18986 (n_6782, n11739);
  not g18987 (n_6783, n12300);
  and g18988 (n12301, n_6782, n_6783);
  not g18989 (n_6784, n12299);
  and g18990 (n12302, n_6784, n12301);
  not g18991 (n_6785, n12302);
  and g18992 (n12303, n_6782, n_6785);
  not g18993 (n_6786, n11713);
  and g18994 (n12304, n_6786, n11723);
  not g18995 (n_6787, n11724);
  not g18996 (n_6788, n12304);
  and g18997 (n12305, n_6787, n_6788);
  not g18998 (n_6789, n12303);
  and g18999 (n12306, n_6789, n12305);
  not g19000 (n_6790, n12306);
  and g19001 (n12307, n_6787, n_6790);
  not g19002 (n_6791, n12307);
  and g19003 (n12308, n11711, n_6791);
  not g19004 (n_6792, n12308);
  and g19005 (n12309, n_6286, n_6792);
  not g19006 (n_6793, n11086);
  and g19007 (n12310, n11083, n_6793);
  not g19008 (n_6794, n11087);
  not g19009 (n_6795, n12310);
  and g19010 (n12311, n_6794, n_6795);
  not g19011 (n_6796, n12309);
  and g19012 (n12312, n_6796, n12311);
  not g19013 (n_6797, n12312);
  and g19014 (n12313, n_6794, n_6797);
  not g19015 (n_6798, n11049);
  and g19016 (n12314, n11047, n_6798);
  not g19017 (n_6799, n11050);
  not g19018 (n_6800, n12314);
  and g19019 (n12315, n_6799, n_6800);
  not g19020 (n_6801, n12313);
  and g19021 (n12316, n_6801, n12315);
  not g19022 (n_6802, n12316);
  and g19023 (n12317, n_6799, n_6802);
  not g19024 (n_6803, n12317);
  and g19025 (n12318, n10453, n_6803);
  not g19026 (n_6804, n12318);
  and g19027 (n12319, n_5195, n_6804);
  not g19028 (n_6805, n9886);
  and g19029 (n12320, n9883, n_6805);
  not g19030 (n_6806, n9887);
  not g19031 (n_6807, n12320);
  and g19032 (n12321, n_6806, n_6807);
  not g19033 (n_6808, n12319);
  and g19034 (n12322, n_6808, n12321);
  not g19035 (n_6809, n12322);
  and g19036 (n12323, n_6806, n_6809);
  not g19037 (n_6810, n9365);
  and g19038 (n12324, n9363, n_6810);
  not g19039 (n_6811, n9366);
  not g19040 (n_6812, n12324);
  and g19041 (n12325, n_6811, n_6812);
  not g19042 (n_6813, n12323);
  and g19043 (n12326, n_6813, n12325);
  not g19044 (n_6814, n12326);
  and g19045 (n12327, n_6811, n_6814);
  not g19046 (n_6815, n12327);
  and g19047 (n12328, n8879, n_6815);
  not g19048 (n_6816, n12328);
  and g19049 (n12329, n_3825, n_6816);
  not g19050 (n_6817, n12329);
  and g19051 (n12330, n8437, n_6817);
  not g19052 (n_6818, n12330);
  and g19053 (n12331, n_3444, n_6818);
  not g19054 (n_6819, n8017);
  and g19055 (n12332, n8015, n_6819);
  not g19056 (n_6820, n8018);
  not g19057 (n_6821, n12332);
  and g19058 (n12333, n_6820, n_6821);
  not g19059 (n_6822, n12331);
  and g19060 (n12334, n_6822, n12333);
  not g19061 (n_6823, n12334);
  and g19062 (n12335, n_6820, n_6823);
  not g19063 (n_6824, n12335);
  and g19064 (n12336, n7651, n_6824);
  not g19065 (n_6825, n12336);
  and g19066 (n12337, n_2759, n_6825);
  not g19067 (n_6826, n7310);
  and g19068 (n12338, n7307, n_6826);
  not g19069 (n_6827, n7311);
  not g19070 (n_6828, n12338);
  and g19071 (n12339, n_6827, n_6828);
  not g19072 (n_6829, n12337);
  and g19073 (n12340, n_6829, n12339);
  not g19074 (n_6830, n12340);
  and g19075 (n12341, n_6827, n_6830);
  not g19076 (n_6831, n7135);
  and g19077 (n12342, n7133, n_6831);
  not g19078 (n_6832, n7136);
  not g19079 (n_6833, n12342);
  and g19080 (n12343, n_6832, n_6833);
  not g19081 (n_6834, n12341);
  and g19082 (n12344, n_6834, n12343);
  not g19083 (n_6835, n12344);
  and g19084 (n12345, n_6832, n_6835);
  not g19085 (n_6836, n12345);
  and g19086 (n12346, n6970, n_6836);
  not g19087 (n_6837, n12346);
  and g19088 (n12347, n_2168, n_6837);
  not g19089 (n_6838, n12347);
  and g19090 (n12348, n6422, n_6838);
  not g19091 (n_6839, n12348);
  and g19092 (n12349, n_1905, n_6839);
  not g19093 (n_6840, n12349);
  and g19094 (n12350, n6267, n_6840);
  not g19095 (n_6841, n12350);
  and g19096 (n12351, n_1767, n_6841);
  not g19097 (n_6842, n12351);
  and g19098 (n12352, n5952, n_6842);
  not g19099 (n_6843, n12352);
  and g19100 (n12353, n_1580, n_6843);
  not g19101 (n_6844, n5681);
  and g19102 (n12354, n5679, n_6844);
  not g19103 (n_6845, n5682);
  not g19104 (n_6846, n12354);
  and g19105 (n12355, n_6845, n_6846);
  not g19106 (n_6847, n12353);
  and g19107 (n12356, n_6847, n12355);
  not g19108 (n_6848, n12356);
  and g19109 (n12357, n_6845, n_6848);
  not g19110 (n_6849, n12357);
  and g19111 (n12358, n5530, n_6849);
  not g19112 (n_6850, n12358);
  and g19113 (n12359, n_1289, n_6850);
  not g19114 (n_6851, n12359);
  and g19115 (n12360, n5420, n_6851);
  not g19116 (n_6852, n12360);
  and g19117 (n12361, n_1196, n_6852);
  not g19118 (n_6853, n12361);
  and g19119 (n12362, n4954, n_6853);
  not g19120 (n_6854, n12362);
  and g19121 (n12363, n_1027, n_6854);
  not g19122 (n_6855, n4730);
  and g19123 (n12364, n4728, n_6855);
  not g19124 (n_6856, n4731);
  not g19125 (n_6857, n12364);
  and g19126 (n12365, n_6856, n_6857);
  not g19127 (n_6858, n12363);
  and g19128 (n12366, n_6858, n12365);
  not g19129 (n_6859, n12366);
  and g19130 (n12367, n_6856, n_6859);
  not g19131 (n_6860, n12367);
  and g19132 (n12368, n4622, n_6860);
  not g19133 (n_6861, n4622);
  and g19134 (n12369, n_6861, n12367);
  not g19135 (n_6862, n12368);
  not g19136 (n_6863, n12369);
  and g19137 (n12370, n_6862, n_6863);
  and g19138 (n12371, n_810, n_6862);
  and g19139 (n12372, n_740, n_743);
  and g19140 (n12373, n3457, n_565);
  and g19141 (n12374, n_480, n3542);
  and g19142 (n12375, n3606, n_535);
  and g19148 (n12378, n3368, n4558);
  not g19151 (n_6868, n12379);
  and g19152 (n12380, \a[29] , n_6868);
  not g19153 (n_6869, n12380);
  and g19154 (n12381, \a[29] , n_6869);
  and g19155 (n12382, n_6868, n_6869);
  not g19156 (n_6870, n12381);
  not g19157 (n_6871, n12382);
  and g19158 (n12383, n_6870, n_6871);
  and g19159 (n12384, n_527, n_532);
  and g19172 (n12397, n_171, n_294);
  not g19224 (n_6872, n12448);
  and g19225 (n12449, n_512, n_6872);
  and g19226 (n12450, n3702, n12448);
  not g19227 (n_6873, n12449);
  not g19228 (n_6874, n12450);
  and g19229 (n12451, n_6873, n_6874);
  and g19230 (n12452, n_27, n12451);
  not g19231 (n_6875, n12452);
  and g19232 (n12453, n_27, n_6875);
  and g19233 (n12454, n_6873, n_6875);
  and g19234 (n12455, n_6874, n12454);
  not g19235 (n_6876, n12453);
  not g19236 (n_6877, n12455);
  and g19237 (n12456, n_6876, n_6877);
  and g19238 (n12457, n3020, n_485);
  and g19239 (n12458, n3028, n_484);
  and g19240 (n12459, n_415, n3023);
  and g19241 (n12460, n75, n4084);
  not g19249 (n_6882, n12456);
  not g19250 (n_6883, n12463);
  and g19251 (n12464, n_6882, n_6883);
  and g19252 (n12465, n12456, n12463);
  not g19253 (n_6884, n12464);
  not g19254 (n_6885, n12465);
  and g19255 (n12466, n_6884, n_6885);
  not g19256 (n_6886, n3708);
  and g19257 (n12467, n_6886, n12466);
  not g19258 (n_6887, n12466);
  and g19259 (n12468, n3708, n_6887);
  not g19260 (n_6888, n12467);
  not g19261 (n_6889, n12468);
  and g19262 (n12469, n_6888, n_6889);
  not g19263 (n_6890, n12384);
  and g19264 (n12470, n_6890, n12469);
  not g19265 (n_6891, n12469);
  and g19266 (n12471, n12384, n_6891);
  not g19267 (n_6892, n12470);
  not g19268 (n_6893, n12471);
  and g19269 (n12472, n_6892, n_6893);
  not g19270 (n_6894, n12383);
  and g19271 (n12473, n_6894, n12472);
  not g19272 (n_6895, n12473);
  and g19273 (n12474, n12472, n_6895);
  and g19274 (n12475, n_6894, n_6895);
  not g19275 (n_6896, n12474);
  not g19276 (n_6897, n12475);
  and g19277 (n12476, n_6896, n_6897);
  and g19278 (n12477, n_554, n_590);
  and g19279 (n12478, n3884, n_712);
  and g19280 (n12479, n3967, n_566);
  and g19281 (n12480, n_560, n4046);
  not g19282 (n_6898, n12479);
  not g19283 (n_6899, n12480);
  and g19284 (n12481, n_6898, n_6899);
  not g19285 (n_6900, n12478);
  and g19286 (n12482, n_6900, n12481);
  and g19287 (n12483, n_750, n12482);
  and g19288 (n12484, n_888, n12482);
  not g19289 (n_6901, n12483);
  not g19290 (n_6902, n12484);
  and g19291 (n12485, n_6901, n_6902);
  not g19292 (n_6903, n12485);
  and g19293 (n12486, \a[26] , n_6903);
  and g19294 (n12487, n_33, n12485);
  not g19295 (n_6904, n12486);
  not g19296 (n_6905, n12487);
  and g19297 (n12488, n_6904, n_6905);
  not g19298 (n_6906, n12477);
  not g19299 (n_6907, n12488);
  and g19300 (n12489, n_6906, n_6907);
  not g19301 (n_6908, n12489);
  and g19302 (n12490, n_6906, n_6908);
  and g19303 (n12491, n_6907, n_6908);
  not g19304 (n_6909, n12490);
  not g19305 (n_6910, n12491);
  and g19306 (n12492, n_6909, n_6910);
  not g19307 (n_6911, n12476);
  not g19308 (n_6912, n12492);
  and g19309 (n12493, n_6911, n_6912);
  and g19310 (n12494, n12476, n_6910);
  and g19311 (n12495, n_6909, n12494);
  not g19312 (n_6913, n12493);
  not g19313 (n_6914, n12495);
  and g19314 (n12496, n_6913, n_6914);
  not g19315 (n_6915, n12372);
  and g19316 (n12497, n_6915, n12496);
  not g19317 (n_6916, n12496);
  and g19318 (n12498, n12372, n_6916);
  not g19319 (n_6917, n12497);
  not g19320 (n_6918, n12498);
  and g19321 (n12499, n_6917, n_6918);
  not g19322 (n_6919, n12371);
  and g19323 (n12500, n_6919, n12499);
  not g19324 (n_6920, n12499);
  and g19325 (n12501, n12371, n_6920);
  not g19326 (n_6921, n12500);
  not g19327 (n_6922, n12501);
  and g19328 (n12502, n_6921, n_6922);
  and g19329 (n12503, n12370, n12502);
  not g19330 (n_6923, n12365);
  and g19331 (n12504, n12363, n_6923);
  not g19332 (n_6924, n12504);
  and g19333 (n12505, n_6859, n_6924);
  and g19334 (n12506, n12370, n12505);
  not g19335 (n_6925, n4954);
  and g19336 (n12507, n_6925, n12361);
  not g19337 (n_6926, n12507);
  and g19338 (n12508, n_6854, n_6926);
  and g19339 (n12509, n12505, n12508);
  not g19340 (n_6927, n5530);
  and g19341 (n12510, n_6927, n12357);
  not g19342 (n_6928, n12510);
  and g19343 (n12511, n_6850, n_6928);
  not g19344 (n_6929, n5420);
  and g19345 (n12512, n_6929, n12359);
  not g19346 (n_6930, n12512);
  and g19347 (n12513, n_6852, n_6930);
  and g19348 (n12514, n12511, n12513);
  not g19349 (n_6931, n12355);
  and g19350 (n12515, n12353, n_6931);
  not g19351 (n_6932, n12515);
  and g19352 (n12516, n_6848, n_6932);
  and g19353 (n12517, n12511, n12516);
  not g19354 (n_6933, n5952);
  and g19355 (n12518, n_6933, n12351);
  not g19356 (n_6934, n12518);
  and g19357 (n12519, n_6843, n_6934);
  and g19358 (n12520, n12516, n12519);
  not g19359 (n_6935, n6267);
  and g19360 (n12521, n_6935, n12349);
  not g19361 (n_6936, n12521);
  and g19362 (n12522, n_6841, n_6936);
  and g19363 (n12523, n12519, n12522);
  not g19364 (n_6937, n6422);
  and g19365 (n12524, n_6937, n12347);
  not g19366 (n_6938, n12524);
  and g19367 (n12525, n_6839, n_6938);
  and g19368 (n12526, n12522, n12525);
  not g19369 (n_6939, n6970);
  and g19370 (n12527, n_6939, n12345);
  not g19371 (n_6940, n12527);
  and g19372 (n12528, n_6837, n_6940);
  and g19373 (n12529, n12525, n12528);
  not g19374 (n_6941, n12343);
  and g19375 (n12530, n12341, n_6941);
  not g19376 (n_6942, n12530);
  and g19377 (n12531, n_6835, n_6942);
  and g19378 (n12532, n12528, n12531);
  not g19379 (n_6943, n12339);
  and g19380 (n12533, n12337, n_6943);
  not g19381 (n_6944, n12533);
  and g19382 (n12534, n_6830, n_6944);
  and g19383 (n12535, n12531, n12534);
  not g19384 (n_6945, n7651);
  and g19385 (n12536, n_6945, n12335);
  not g19386 (n_6946, n12536);
  and g19387 (n12537, n_6825, n_6946);
  and g19388 (n12538, n12534, n12537);
  not g19389 (n_6947, n12333);
  and g19390 (n12539, n12331, n_6947);
  not g19391 (n_6948, n12539);
  and g19392 (n12540, n_6823, n_6948);
  and g19393 (n12541, n12537, n12540);
  not g19394 (n_6949, n8437);
  and g19395 (n12542, n_6949, n12329);
  not g19396 (n_6950, n12542);
  and g19397 (n12543, n_6818, n_6950);
  and g19398 (n12544, n12540, n12543);
  not g19399 (n_6951, n8879);
  and g19400 (n12545, n_6951, n12327);
  not g19401 (n_6952, n12545);
  and g19402 (n12546, n_6816, n_6952);
  and g19403 (n12547, n12543, n12546);
  not g19404 (n_6953, n12325);
  and g19405 (n12548, n12323, n_6953);
  not g19406 (n_6954, n12548);
  and g19407 (n12549, n_6814, n_6954);
  and g19408 (n12550, n12546, n12549);
  not g19409 (n_6955, n12321);
  and g19410 (n12551, n12319, n_6955);
  not g19411 (n_6956, n12551);
  and g19412 (n12552, n_6809, n_6956);
  and g19413 (n12553, n12549, n12552);
  not g19414 (n_6957, n10453);
  and g19415 (n12554, n_6957, n12317);
  not g19416 (n_6958, n12554);
  and g19417 (n12555, n_6804, n_6958);
  and g19418 (n12556, n12552, n12555);
  not g19419 (n_6959, n12315);
  and g19420 (n12557, n12313, n_6959);
  not g19421 (n_6960, n12557);
  and g19422 (n12558, n_6802, n_6960);
  and g19423 (n12559, n12555, n12558);
  not g19424 (n_6961, n12311);
  and g19425 (n12560, n12309, n_6961);
  not g19426 (n_6962, n12560);
  and g19427 (n12561, n_6797, n_6962);
  and g19428 (n12562, n12558, n12561);
  not g19429 (n_6963, n11711);
  and g19430 (n12563, n_6963, n12307);
  not g19431 (n_6964, n12563);
  and g19432 (n12564, n_6792, n_6964);
  and g19433 (n12565, n12561, n12564);
  not g19434 (n_6965, n12305);
  and g19435 (n12566, n12303, n_6965);
  not g19436 (n_6966, n12566);
  and g19437 (n12567, n_6790, n_6966);
  and g19438 (n12568, n12564, n12567);
  not g19439 (n_6967, n12564);
  not g19440 (n_6968, n12567);
  and g19441 (n12569, n_6967, n_6968);
  not g19442 (n_6969, n12301);
  and g19443 (n12570, n12299, n_6969);
  not g19444 (n_6970, n12570);
  and g19445 (n12571, n_6785, n_6970);
  and g19446 (n12572, n12567, n12571);
  not g19447 (n_6971, n12297);
  and g19448 (n12573, n12295, n_6971);
  not g19449 (n_6972, n12573);
  and g19450 (n12574, n_6780, n_6972);
  and g19451 (n12575, n12571, n12574);
  not g19452 (n_6973, n12293);
  and g19453 (n12576, n12291, n_6973);
  not g19454 (n_6974, n12576);
  and g19455 (n12577, n_6775, n_6974);
  and g19456 (n12578, n12574, n12577);
  and g19457 (n12579, n_6768, n_6770);
  and g19458 (n12580, n_6769, n_6770);
  not g19459 (n_6975, n12579);
  not g19460 (n_6976, n12580);
  and g19461 (n12581, n_6975, n_6976);
  not g19462 (n_6977, n12581);
  and g19463 (n12582, n12577, n_6977);
  not g19464 (n_6978, n12574);
  and g19465 (n12583, n_6978, n12582);
  not g19466 (n_6979, n12578);
  not g19467 (n_6980, n12583);
  and g19468 (n12584, n_6979, n_6980);
  not g19469 (n_6981, n12571);
  and g19470 (n12585, n_6981, n_6978);
  not g19471 (n_6982, n12575);
  not g19472 (n_6983, n12585);
  and g19473 (n12586, n_6982, n_6983);
  not g19474 (n_6984, n12584);
  and g19475 (n12587, n_6984, n12586);
  not g19476 (n_6985, n12587);
  and g19477 (n12588, n_6982, n_6985);
  and g19478 (n12589, n_6968, n_6981);
  not g19479 (n_6986, n12572);
  not g19480 (n_6987, n12589);
  and g19481 (n12590, n_6986, n_6987);
  not g19482 (n_6988, n12588);
  and g19483 (n12591, n_6988, n12590);
  not g19484 (n_6989, n12591);
  and g19485 (n12592, n_6986, n_6989);
  not g19486 (n_6990, n12568);
  not g19487 (n_6991, n12592);
  and g19488 (n12593, n_6990, n_6991);
  not g19489 (n_6992, n12569);
  and g19490 (n12594, n_6992, n12593);
  not g19491 (n_6993, n12594);
  and g19492 (n12595, n_6990, n_6993);
  not g19493 (n_6994, n12561);
  and g19494 (n12596, n_6994, n_6967);
  not g19495 (n_6995, n12595);
  not g19496 (n_6996, n12596);
  and g19497 (n12597, n_6995, n_6996);
  not g19498 (n_6997, n12565);
  and g19499 (n12598, n_6997, n12597);
  not g19500 (n_6998, n12598);
  and g19501 (n12599, n_6997, n_6998);
  not g19502 (n_6999, n12558);
  and g19503 (n12600, n_6999, n_6994);
  not g19504 (n_7000, n12562);
  not g19505 (n_7001, n12600);
  and g19506 (n12601, n_7000, n_7001);
  not g19507 (n_7002, n12599);
  and g19508 (n12602, n_7002, n12601);
  not g19509 (n_7003, n12602);
  and g19510 (n12603, n_7000, n_7003);
  not g19511 (n_7004, n12555);
  and g19512 (n12604, n_7004, n_6999);
  not g19513 (n_7005, n12603);
  not g19514 (n_7006, n12604);
  and g19515 (n12605, n_7005, n_7006);
  not g19516 (n_7007, n12559);
  and g19517 (n12606, n_7007, n12605);
  not g19518 (n_7008, n12606);
  and g19519 (n12607, n_7007, n_7008);
  not g19520 (n_7009, n12552);
  and g19521 (n12608, n_7009, n_7004);
  not g19522 (n_7010, n12607);
  not g19523 (n_7011, n12608);
  and g19524 (n12609, n_7010, n_7011);
  not g19525 (n_7012, n12556);
  and g19526 (n12610, n_7012, n12609);
  not g19527 (n_7013, n12610);
  and g19528 (n12611, n_7012, n_7013);
  not g19529 (n_7014, n12549);
  and g19530 (n12612, n_7014, n_7009);
  not g19531 (n_7015, n12553);
  not g19532 (n_7016, n12612);
  and g19533 (n12613, n_7015, n_7016);
  not g19534 (n_7017, n12611);
  and g19535 (n12614, n_7017, n12613);
  not g19536 (n_7018, n12614);
  and g19537 (n12615, n_7015, n_7018);
  not g19538 (n_7019, n12546);
  and g19539 (n12616, n_7019, n_7014);
  not g19540 (n_7020, n12615);
  not g19541 (n_7021, n12616);
  and g19542 (n12617, n_7020, n_7021);
  not g19543 (n_7022, n12550);
  and g19544 (n12618, n_7022, n12617);
  not g19545 (n_7023, n12618);
  and g19546 (n12619, n_7022, n_7023);
  not g19547 (n_7024, n12543);
  and g19548 (n12620, n_7024, n_7019);
  not g19549 (n_7025, n12547);
  not g19550 (n_7026, n12620);
  and g19551 (n12621, n_7025, n_7026);
  not g19552 (n_7027, n12619);
  and g19553 (n12622, n_7027, n12621);
  not g19554 (n_7028, n12622);
  and g19555 (n12623, n_7025, n_7028);
  not g19556 (n_7029, n12540);
  and g19557 (n12624, n_7029, n_7024);
  not g19558 (n_7030, n12623);
  not g19559 (n_7031, n12624);
  and g19560 (n12625, n_7030, n_7031);
  not g19561 (n_7032, n12544);
  and g19562 (n12626, n_7032, n12625);
  not g19563 (n_7033, n12626);
  and g19564 (n12627, n_7032, n_7033);
  not g19565 (n_7034, n12537);
  and g19566 (n12628, n_7034, n_7029);
  not g19567 (n_7035, n12627);
  not g19568 (n_7036, n12628);
  and g19569 (n12629, n_7035, n_7036);
  not g19570 (n_7037, n12541);
  and g19571 (n12630, n_7037, n12629);
  not g19572 (n_7038, n12630);
  and g19573 (n12631, n_7037, n_7038);
  not g19574 (n_7039, n12534);
  and g19575 (n12632, n_7039, n_7034);
  not g19576 (n_7040, n12631);
  not g19577 (n_7041, n12632);
  and g19578 (n12633, n_7040, n_7041);
  not g19579 (n_7042, n12538);
  and g19580 (n12634, n_7042, n12633);
  not g19581 (n_7043, n12634);
  and g19582 (n12635, n_7042, n_7043);
  not g19583 (n_7044, n12531);
  and g19584 (n12636, n_7044, n_7039);
  not g19585 (n_7045, n12535);
  not g19586 (n_7046, n12636);
  and g19587 (n12637, n_7045, n_7046);
  not g19588 (n_7047, n12635);
  and g19589 (n12638, n_7047, n12637);
  not g19590 (n_7048, n12638);
  and g19591 (n12639, n_7045, n_7048);
  not g19592 (n_7049, n12528);
  and g19593 (n12640, n_7049, n_7044);
  not g19594 (n_7050, n12639);
  not g19595 (n_7051, n12640);
  and g19596 (n12641, n_7050, n_7051);
  not g19597 (n_7052, n12532);
  and g19598 (n12642, n_7052, n12641);
  not g19599 (n_7053, n12642);
  and g19600 (n12643, n_7052, n_7053);
  not g19601 (n_7054, n12525);
  and g19602 (n12644, n_7054, n_7049);
  not g19603 (n_7055, n12529);
  not g19604 (n_7056, n12644);
  and g19605 (n12645, n_7055, n_7056);
  not g19606 (n_7057, n12643);
  and g19607 (n12646, n_7057, n12645);
  not g19608 (n_7058, n12646);
  and g19609 (n12647, n_7055, n_7058);
  not g19610 (n_7059, n12522);
  and g19611 (n12648, n_7059, n_7054);
  not g19612 (n_7060, n12526);
  not g19613 (n_7061, n12648);
  and g19614 (n12649, n_7060, n_7061);
  not g19615 (n_7062, n12647);
  and g19616 (n12650, n_7062, n12649);
  not g19617 (n_7063, n12650);
  and g19618 (n12651, n_7060, n_7063);
  not g19619 (n_7064, n12519);
  and g19620 (n12652, n_7064, n_7059);
  not g19621 (n_7065, n12523);
  not g19622 (n_7066, n12652);
  and g19623 (n12653, n_7065, n_7066);
  not g19624 (n_7067, n12651);
  and g19625 (n12654, n_7067, n12653);
  not g19626 (n_7068, n12654);
  and g19627 (n12655, n_7065, n_7068);
  not g19628 (n_7069, n12516);
  and g19629 (n12656, n_7069, n_7064);
  not g19630 (n_7070, n12655);
  not g19631 (n_7071, n12656);
  and g19632 (n12657, n_7070, n_7071);
  not g19633 (n_7072, n12520);
  and g19634 (n12658, n_7072, n12657);
  not g19635 (n_7073, n12658);
  and g19636 (n12659, n_7072, n_7073);
  not g19637 (n_7074, n12511);
  and g19638 (n12660, n_7074, n_7069);
  not g19639 (n_7075, n12659);
  not g19640 (n_7076, n12660);
  and g19641 (n12661, n_7075, n_7076);
  not g19642 (n_7077, n12517);
  and g19643 (n12662, n_7077, n12661);
  not g19644 (n_7078, n12662);
  and g19645 (n12663, n_7077, n_7078);
  not g19646 (n_7079, n12513);
  and g19647 (n12664, n_7074, n_7079);
  not g19648 (n_7080, n12514);
  not g19649 (n_7081, n12664);
  and g19650 (n12665, n_7080, n_7081);
  not g19651 (n_7082, n12663);
  and g19652 (n12666, n_7082, n12665);
  not g19653 (n_7083, n12666);
  and g19654 (n12667, n_7080, n_7083);
  not g19655 (n_7084, n12508);
  and g19656 (n12668, n_7084, n_7079);
  and g19657 (n12669, n12508, n12513);
  not g19658 (n_7085, n12668);
  not g19659 (n_7086, n12669);
  and g19660 (n12670, n_7085, n_7086);
  not g19661 (n_7087, n12667);
  and g19662 (n12671, n_7087, n12670);
  not g19663 (n_7088, n12671);
  and g19664 (n12672, n_7086, n_7088);
  not g19665 (n_7089, n12505);
  and g19666 (n12673, n_7089, n_7084);
  not g19667 (n_7090, n12672);
  not g19668 (n_7091, n12673);
  and g19669 (n12674, n_7090, n_7091);
  not g19670 (n_7092, n12509);
  and g19671 (n12675, n_7092, n12674);
  not g19672 (n_7093, n12675);
  and g19673 (n12676, n_7092, n_7093);
  not g19674 (n_7094, n12370);
  and g19675 (n12677, n_7094, n_7089);
  not g19676 (n_7095, n12676);
  not g19677 (n_7096, n12677);
  and g19678 (n12678, n_7095, n_7096);
  not g19679 (n_7097, n12506);
  and g19680 (n12679, n_7097, n12678);
  not g19681 (n_7098, n12679);
  and g19682 (n12680, n_7097, n_7098);
  not g19683 (n_7099, n12502);
  and g19684 (n12681, n_7094, n_7099);
  not g19685 (n_7100, n12680);
  not g19686 (n_7101, n12681);
  and g19687 (n12682, n_7100, n_7101);
  not g19688 (n_7102, n12503);
  and g19689 (n12683, n_7102, n12682);
  not g19690 (n_7103, n12683);
  and g19691 (n12684, n_7102, n_7103);
  and g19692 (n12685, n_6917, n_6921);
  and g19693 (n12686, n_6908, n_6913);
  and g19694 (n12687, n_560, n3967);
  and g19695 (n12688, n4046, n_712);
  not g19696 (n_7104, n12687);
  not g19697 (n_7105, n12688);
  and g19698 (n12689, n_7104, n_7105);
  and g19699 (n12690, n4050, n4609);
  not g19700 (n_7106, n12690);
  and g19701 (n12691, n12689, n_7106);
  not g19702 (n_7107, n12691);
  and g19703 (n12692, \a[26] , n_7107);
  not g19704 (n_7108, n12692);
  and g19705 (n12693, n_7107, n_7108);
  and g19706 (n12694, \a[26] , n_7108);
  not g19707 (n_7109, n12693);
  not g19708 (n_7110, n12694);
  and g19709 (n12695, n_7109, n_7110);
  and g19710 (n12696, n_6892, n_6895);
  and g19711 (n12697, n75, n3627);
  and g19712 (n12698, n3020, n_480);
  and g19713 (n12699, n3023, n_484);
  and g19714 (n12700, n3028, n_485);
  and g19729 (n12711, n_90, n_235);
  and g19730 (n12712, n_73, n12711);
  not g19749 (n_7115, n12454);
  and g19750 (n12731, n_7115, n12730);
  not g19751 (n_7116, n12730);
  and g19752 (n12732, n12454, n_7116);
  not g19753 (n_7117, n12731);
  not g19754 (n_7118, n12732);
  and g19755 (n12733, n_7117, n_7118);
  not g19756 (n_7119, n12703);
  and g19757 (n12734, n_7119, n12733);
  not g19758 (n_7120, n12734);
  and g19759 (n12735, n_7119, n_7120);
  and g19760 (n12736, n12733, n_7120);
  not g19761 (n_7121, n12735);
  not g19762 (n_7122, n12736);
  and g19763 (n12737, n_7121, n_7122);
  and g19764 (n12738, n_6884, n_6888);
  and g19765 (n12739, n12737, n12738);
  not g19766 (n_7123, n12737);
  not g19767 (n_7124, n12738);
  and g19768 (n12740, n_7123, n_7124);
  not g19769 (n_7125, n12739);
  not g19770 (n_7126, n12740);
  and g19771 (n12741, n_7125, n_7126);
  and g19772 (n12742, n3457, n_566);
  and g19773 (n12743, n3542, n_535);
  and g19774 (n12744, n3606, n_565);
  not g19775 (n_7127, n12743);
  not g19776 (n_7128, n12744);
  and g19777 (n12745, n_7127, n_7128);
  not g19778 (n_7129, n12742);
  and g19779 (n12746, n_7129, n12745);
  and g19780 (n12747, n_489, n12746);
  and g19781 (n12748, n_6323, n12746);
  not g19782 (n_7130, n12747);
  not g19783 (n_7131, n12748);
  and g19784 (n12749, n_7130, n_7131);
  not g19785 (n_7132, n12749);
  and g19786 (n12750, \a[29] , n_7132);
  and g19787 (n12751, n_15, n12749);
  not g19788 (n_7133, n12750);
  not g19789 (n_7134, n12751);
  and g19790 (n12752, n_7133, n_7134);
  not g19791 (n_7135, n12752);
  and g19792 (n12753, n12741, n_7135);
  not g19793 (n_7136, n12741);
  and g19794 (n12754, n_7136, n12752);
  not g19795 (n_7137, n12753);
  not g19796 (n_7138, n12754);
  and g19797 (n12755, n_7137, n_7138);
  not g19798 (n_7139, n12696);
  and g19799 (n12756, n_7139, n12755);
  not g19800 (n_7140, n12756);
  and g19801 (n12757, n_7139, n_7140);
  and g19802 (n12758, n12755, n_7140);
  not g19803 (n_7141, n12757);
  not g19804 (n_7142, n12758);
  and g19805 (n12759, n_7141, n_7142);
  not g19806 (n_7143, n12695);
  not g19807 (n_7144, n12759);
  and g19808 (n12760, n_7143, n_7144);
  and g19809 (n12761, n12695, n_7142);
  and g19810 (n12762, n_7141, n12761);
  not g19811 (n_7145, n12760);
  not g19812 (n_7146, n12762);
  and g19813 (n12763, n_7145, n_7146);
  not g19814 (n_7147, n12686);
  and g19815 (n12764, n_7147, n12763);
  not g19816 (n_7148, n12763);
  and g19817 (n12765, n12686, n_7148);
  not g19818 (n_7149, n12764);
  not g19819 (n_7150, n12765);
  and g19820 (n12766, n_7149, n_7150);
  not g19821 (n_7151, n12685);
  and g19822 (n12767, n_7151, n12766);
  not g19823 (n_7152, n12766);
  and g19824 (n12768, n12685, n_7152);
  not g19825 (n_7153, n12767);
  not g19826 (n_7154, n12768);
  and g19827 (n12769, n_7153, n_7154);
  not g19828 (n_7155, n12769);
  and g19829 (n12770, n_7099, n_7155);
  and g19830 (n12771, n12502, n12769);
  not g19831 (n_7156, n12770);
  not g19832 (n_7157, n12771);
  and g19833 (n12772, n_7156, n_7157);
  not g19834 (n_7158, n12684);
  and g19835 (n12773, n_7158, n12772);
  not g19836 (n_7159, n12773);
  and g19837 (n12774, n_7157, n_7159);
  and g19838 (n12775, n_7149, n_7153);
  and g19839 (n12776, n_7140, n_7145);
  and g19840 (n12777, n75, n3818);
  and g19841 (n12778, n3020, n_535);
  and g19842 (n12779, n3023, n_485);
  and g19843 (n12780, n3028, n_480);
  and g19851 (n12784, n_107, n_128);
  and g19852 (n12785, n_265, n12784);
  and g19878 (n12811, n_173, n_210);
  and g19879 (n12812, n_242, n12811);
  and g19896 (n12829, n_140, n_184);
  and g19897 (n12830, n_104, n12829);
  and g19910 (n12843, n_7116, n12842);
  not g19911 (n_7164, n12842);
  and g19912 (n12844, n12730, n_7164);
  not g19913 (n_7165, n12783);
  not g19914 (n_7166, n12844);
  and g19915 (n12845, n_7165, n_7166);
  not g19916 (n_7167, n12843);
  and g19917 (n12846, n_7167, n12845);
  not g19918 (n_7168, n12846);
  and g19919 (n12847, n_7165, n_7168);
  and g19920 (n12848, n_7166, n_7168);
  and g19921 (n12849, n_7167, n12848);
  not g19922 (n_7169, n12847);
  not g19923 (n_7170, n12849);
  and g19924 (n12850, n_7169, n_7170);
  and g19925 (n12851, n_7117, n_7120);
  and g19926 (n12852, n12850, n12851);
  not g19927 (n_7171, n12850);
  not g19928 (n_7172, n12851);
  and g19929 (n12853, n_7171, n_7172);
  not g19930 (n_7173, n12852);
  not g19931 (n_7174, n12853);
  and g19932 (n12854, n_7173, n_7174);
  and g19933 (n12855, n_7126, n_7137);
  not g19934 (n_7175, n12855);
  and g19935 (n12856, n12854, n_7175);
  not g19936 (n_7176, n12854);
  and g19937 (n12857, n_7176, n12855);
  not g19938 (n_7177, n12856);
  not g19939 (n_7178, n12857);
  and g19940 (n12858, n_7177, n_7178);
  and g19941 (n12859, n4050, n4522);
  and g19942 (n12860, n3967, n_712);
  not g19943 (n_7179, n12859);
  not g19944 (n_7180, n12860);
  and g19945 (n12861, n_7179, n_7180);
  not g19946 (n_7181, n12861);
  and g19947 (n12862, \a[26] , n_7181);
  not g19948 (n_7182, n12862);
  and g19949 (n12863, n_7181, n_7182);
  and g19950 (n12864, \a[26] , n_7182);
  not g19951 (n_7183, n12863);
  not g19952 (n_7184, n12864);
  and g19953 (n12865, n_7183, n_7184);
  and g19954 (n12866, n3457, n_560);
  and g19955 (n12867, n3542, n_565);
  and g19956 (n12868, n3606, n_566);
  and g19962 (n12871, n3368, n4067);
  not g19965 (n_7189, n12872);
  and g19966 (n12873, \a[29] , n_7189);
  not g19967 (n_7190, n12873);
  and g19968 (n12874, \a[29] , n_7190);
  and g19969 (n12875, n_7189, n_7190);
  not g19970 (n_7191, n12874);
  not g19971 (n_7192, n12875);
  and g19972 (n12876, n_7191, n_7192);
  not g19973 (n_7193, n12865);
  not g19974 (n_7194, n12876);
  and g19975 (n12877, n_7193, n_7194);
  not g19976 (n_7195, n12877);
  and g19977 (n12878, n_7193, n_7195);
  and g19978 (n12879, n_7194, n_7195);
  not g19979 (n_7196, n12878);
  not g19980 (n_7197, n12879);
  and g19981 (n12880, n_7196, n_7197);
  not g19982 (n_7198, n12880);
  and g19983 (n12881, n12858, n_7198);
  not g19984 (n_7199, n12858);
  and g19985 (n12882, n_7199, n12880);
  not g19986 (n_7200, n12881);
  not g19987 (n_7201, n12882);
  and g19988 (n12883, n_7200, n_7201);
  not g19989 (n_7202, n12776);
  and g19990 (n12884, n_7202, n12883);
  not g19991 (n_7203, n12883);
  and g19992 (n12885, n12776, n_7203);
  not g19993 (n_7204, n12884);
  not g19994 (n_7205, n12885);
  and g19995 (n12886, n_7204, n_7205);
  not g19996 (n_7206, n12775);
  and g19997 (n12887, n_7206, n12886);
  not g19998 (n_7207, n12886);
  and g19999 (n12888, n12775, n_7207);
  not g20000 (n_7208, n12887);
  not g20001 (n_7209, n12888);
  and g20002 (n12889, n_7208, n_7209);
  not g20003 (n_7210, n12889);
  and g20004 (n12890, n_7155, n_7210);
  and g20005 (n12891, n12769, n12889);
  not g20006 (n_7211, n12890);
  not g20007 (n_7212, n12891);
  and g20008 (n12892, n_7211, n_7212);
  not g20009 (n_7213, n12774);
  and g20010 (n12893, n_7213, n12892);
  not g20011 (n_7214, n12892);
  and g20012 (n12894, n12774, n_7214);
  not g20013 (n_7215, n12893);
  not g20014 (n_7216, n12894);
  and g20015 (n12895, n_7215, n_7216);
  and g20016 (n12896, n75, n12895);
  and g20017 (n12897, n3020, n12889);
  and g20018 (n12898, n3023, n12502);
  and g20019 (n12899, n3028, n12769);
  and g20034 (n12910, n230, n_129);
  and g20035 (n12911, n_135, n12910);
  and g20064 (n12940, n_153, n_284);
  and g20065 (n12941, n_55, n12940);
  not g20120 (n_7221, n12995);
  and g20121 (n12996, n12958, n_7221);
  not g20122 (n_7222, n12958);
  and g20123 (n12997, n_7222, n12995);
  not g20124 (n_7223, n12772);
  and g20125 (n12998, n12684, n_7223);
  not g20126 (n_7224, n12998);
  and g20127 (n12999, n_7159, n_7224);
  and g20128 (n13000, n75, n12999);
  and g20129 (n13001, n3020, n12769);
  and g20130 (n13002, n3023, n12370);
  and g20131 (n13003, n3028, n12502);
  not g20139 (n_7229, n12996);
  not g20140 (n_7230, n13006);
  and g20141 (n13007, n_7229, n_7230);
  not g20142 (n_7231, n12997);
  and g20143 (n13008, n_7231, n13007);
  not g20144 (n_7232, n13008);
  and g20145 (n13009, n_7229, n_7232);
  and g20149 (n13013, n_156, n_272);
  and g20150 (n13014, n_150, n13013);
  and g20151 (n13015, n_178, n_258);
  and g20152 (n13016, n_206, n13015);
  and g20211 (n13075, n3569, n3906);
  and g20218 (n13082, n13074, n13081);
  not g20219 (n_7233, n13059);
  and g20220 (n13083, n_7233, n13082);
  not g20233 (n_7234, n13095);
  and g20234 (n13096, n13074, n_7234);
  not g20235 (n_7235, n13074);
  and g20236 (n13097, n_7235, n13095);
  and g20237 (n13098, n75, n4522);
  and g20238 (n13099, n3023, n_712);
  not g20239 (n_7236, n13098);
  not g20240 (n_7237, n13099);
  and g20241 (n13100, n_7236, n_7237);
  not g20242 (n_7238, n13096);
  not g20243 (n_7239, n13100);
  and g20244 (n13101, n_7238, n_7239);
  not g20245 (n_7240, n13097);
  and g20246 (n13102, n_7240, n13101);
  not g20247 (n_7241, n13102);
  and g20248 (n13103, n_7238, n_7241);
  not g20249 (n_7242, n13081);
  and g20250 (n13104, n_7235, n_7242);
  not g20251 (n_7243, n13082);
  not g20252 (n_7244, n13104);
  and g20253 (n13105, n_7243, n_7244);
  not g20254 (n_7245, n13103);
  not g20255 (n_7246, n13105);
  and g20256 (n13106, n_7245, n_7246);
  not g20257 (n_7247, n13106);
  and g20258 (n13107, n_7245, n_7247);
  and g20259 (n13108, n_7246, n_7247);
  not g20260 (n_7248, n13107);
  not g20261 (n_7249, n13108);
  and g20262 (n13109, n_7248, n_7249);
  and g20263 (n13110, n_7239, n_7241);
  and g20264 (n13111, n_7240, n13103);
  not g20265 (n_7250, n13110);
  not g20266 (n_7251, n13111);
  and g20267 (n13112, n_7250, n_7251);
  and g20268 (n13113, n_114, n_297);
  and g20269 (n13114, n_102, n13113);
  not g20328 (n_7252, n13158);
  not g20329 (n_7253, n13172);
  and g20330 (n13173, n_7252, n_7253);
  and g20331 (n13174, n13158, n13172);
  not g20332 (n_7254, n13173);
  not g20333 (n_7255, n13174);
  and g20334 (n13175, n_7254, n_7255);
  and g20335 (n13176, n_15, n13175);
  not g20336 (n_7256, n13176);
  and g20337 (n13177, n_7254, n_7256);
  not g20338 (n_7257, n13177);
  and g20339 (n13178, n13074, n_7257);
  and g20340 (n13179, n75, n4609);
  and g20341 (n13180, n3023, n_560);
  and g20342 (n13181, n3028, n_712);
  not g20343 (n_7258, n13180);
  not g20344 (n_7259, n13181);
  and g20345 (n13182, n_7258, n_7259);
  not g20346 (n_7260, n13179);
  and g20347 (n13183, n_7260, n13182);
  and g20348 (n13184, n_7235, n13177);
  not g20349 (n_7261, n13178);
  not g20350 (n_7262, n13184);
  and g20351 (n13185, n_7261, n_7262);
  not g20352 (n_7263, n13183);
  and g20353 (n13186, n_7263, n13185);
  not g20354 (n_7264, n13186);
  and g20355 (n13187, n_7261, n_7264);
  not g20356 (n_7265, n13112);
  not g20357 (n_7266, n13187);
  and g20358 (n13188, n_7265, n_7266);
  and g20359 (n13189, n13112, n13187);
  not g20360 (n_7267, n13188);
  not g20361 (n_7268, n13189);
  and g20362 (n13190, n_7267, n_7268);
  and g20363 (n13191, n_7263, n_7264);
  and g20364 (n13192, n13185, n_7264);
  not g20365 (n_7269, n13191);
  not g20366 (n_7270, n13192);
  and g20367 (n13193, n_7269, n_7270);
  and g20368 (n13194, n_15, n_7256);
  and g20369 (n13195, n_7255, n13177);
  not g20370 (n_7271, n13194);
  not g20371 (n_7272, n13195);
  and g20372 (n13196, n_7271, n_7272);
  not g20415 (n_7273, n13238);
  and g20416 (n13239, n13158, n_7273);
  and g20417 (n13240, n_7252, n13238);
  and g20425 (n13248, n_82, n_273);
  and g20426 (n13249, n_43, n13248);
  not g20461 (n_7274, n13283);
  and g20462 (n13284, n_7116, n_7274);
  and g20463 (n13285, n12730, n13283);
  not g20464 (n_7275, n13284);
  not g20465 (n_7276, n13285);
  and g20466 (n13286, n_7275, n_7276);
  and g20467 (n13287, n_33, n13286);
  not g20468 (n_7277, n13287);
  and g20469 (n13288, n_7275, n_7277);
  not g20470 (n_7278, n13288);
  and g20471 (n13289, n13238, n_7278);
  and g20472 (n13290, n75, n4477);
  and g20473 (n13291, n3020, n_566);
  and g20474 (n13292, n3023, n_535);
  and g20475 (n13293, n3028, n_565);
  and g20483 (n13297, n_7273, n13288);
  not g20484 (n_7283, n13289);
  not g20485 (n_7284, n13297);
  and g20486 (n13298, n_7283, n_7284);
  not g20487 (n_7285, n13296);
  and g20488 (n13299, n_7285, n13298);
  not g20489 (n_7286, n13299);
  and g20490 (n13300, n_7283, n_7286);
  not g20491 (n_7287, n13239);
  not g20492 (n_7288, n13300);
  and g20493 (n13301, n_7287, n_7288);
  not g20494 (n_7289, n13240);
  and g20495 (n13302, n_7289, n13301);
  not g20496 (n_7290, n13302);
  and g20497 (n13303, n_7287, n_7290);
  not g20498 (n_7291, n13196);
  not g20499 (n_7292, n13303);
  and g20500 (n13304, n_7291, n_7292);
  and g20501 (n13305, n75, n4715);
  and g20502 (n13306, n3020, n_712);
  and g20503 (n13307, n3023, n_566);
  and g20504 (n13308, n3028, n_560);
  and g20512 (n13312, n13196, n13303);
  not g20513 (n_7297, n13304);
  not g20514 (n_7298, n13312);
  and g20515 (n13313, n_7297, n_7298);
  not g20516 (n_7299, n13311);
  and g20517 (n13314, n_7299, n13313);
  not g20518 (n_7300, n13314);
  and g20519 (n13315, n_7297, n_7300);
  not g20520 (n_7301, n13193);
  not g20521 (n_7302, n13315);
  and g20522 (n13316, n_7301, n_7302);
  and g20523 (n13317, n13193, n13315);
  not g20524 (n_7303, n13316);
  not g20525 (n_7304, n13317);
  and g20526 (n13318, n_7303, n_7304);
  and g20527 (n13319, n3542, n_712);
  and g20528 (n13320, n3368, n4522);
  not g20529 (n_7305, n13319);
  not g20530 (n_7306, n13320);
  and g20531 (n13321, n_7305, n_7306);
  not g20532 (n_7307, n13321);
  and g20533 (n13322, \a[29] , n_7307);
  not g20534 (n_7308, n13322);
  and g20535 (n13323, n_7307, n_7308);
  and g20536 (n13324, \a[29] , n_7308);
  not g20537 (n_7309, n13323);
  not g20538 (n_7310, n13324);
  and g20539 (n13325, n_7309, n_7310);
  and g20540 (n13326, n75, n4067);
  and g20541 (n13327, n3020, n_560);
  and g20542 (n13328, n3023, n_565);
  and g20543 (n13329, n3028, n_566);
  not g20551 (n_7315, n13325);
  not g20552 (n_7316, n13332);
  and g20553 (n13333, n_7315, n_7316);
  not g20554 (n_7317, n13333);
  and g20555 (n13334, n_7315, n_7317);
  and g20556 (n13335, n_7316, n_7317);
  not g20557 (n_7318, n13334);
  not g20558 (n_7319, n13335);
  and g20559 (n13336, n_7318, n_7319);
  and g20560 (n13337, n_7288, n_7290);
  and g20561 (n13338, n_7289, n13303);
  not g20562 (n_7320, n13337);
  not g20563 (n_7321, n13338);
  and g20564 (n13339, n_7320, n_7321);
  not g20565 (n_7322, n13336);
  not g20566 (n_7323, n13339);
  and g20567 (n13340, n_7322, n_7323);
  not g20568 (n_7324, n13340);
  and g20569 (n13341, n_7317, n_7324);
  not g20570 (n_7325, n13313);
  and g20571 (n13342, n13311, n_7325);
  not g20572 (n_7326, n13342);
  and g20573 (n13343, n_7300, n_7326);
  not g20574 (n_7327, n13341);
  and g20575 (n13344, n_7327, n13343);
  and g20576 (n13345, n_7285, n_7286);
  and g20577 (n13346, n13298, n_7286);
  not g20578 (n_7328, n13345);
  not g20579 (n_7329, n13346);
  and g20580 (n13347, n_7328, n_7329);
  and g20581 (n13348, n_33, n_7277);
  and g20582 (n13349, n_7276, n13288);
  not g20583 (n_7330, n13348);
  not g20584 (n_7331, n13349);
  and g20585 (n13350, n_7330, n_7331);
  not g20586 (n_7332, n12848);
  not g20587 (n_7333, n13350);
  and g20588 (n13351, n_7332, n_7333);
  and g20589 (n13352, n75, n4558);
  and g20590 (n13353, n3020, n_565);
  and g20591 (n13354, n3023, n_480);
  and g20592 (n13355, n3028, n_535);
  and g20600 (n13359, n12848, n13350);
  not g20601 (n_7338, n13351);
  not g20602 (n_7339, n13359);
  and g20603 (n13360, n_7338, n_7339);
  not g20604 (n_7340, n13358);
  and g20605 (n13361, n_7340, n13360);
  not g20606 (n_7341, n13361);
  and g20607 (n13362, n_7338, n_7341);
  not g20608 (n_7342, n13347);
  not g20609 (n_7343, n13362);
  and g20610 (n13363, n_7342, n_7343);
  and g20611 (n13364, n13347, n13362);
  not g20612 (n_7344, n13363);
  not g20613 (n_7345, n13364);
  and g20614 (n13365, n_7344, n_7345);
  and g20615 (n13366, n3542, n_560);
  and g20616 (n13367, n3606, n_712);
  not g20617 (n_7346, n13366);
  not g20618 (n_7347, n13367);
  and g20619 (n13368, n_7346, n_7347);
  and g20620 (n13369, n3368, n4609);
  not g20621 (n_7348, n13369);
  and g20622 (n13370, n13368, n_7348);
  not g20623 (n_7349, n13370);
  and g20624 (n13371, \a[29] , n_7349);
  not g20625 (n_7350, n13371);
  and g20626 (n13372, \a[29] , n_7350);
  and g20627 (n13373, n_7349, n_7350);
  not g20628 (n_7351, n13372);
  not g20629 (n_7352, n13373);
  and g20630 (n13374, n_7351, n_7352);
  not g20631 (n_7353, n13374);
  and g20632 (n13375, n13365, n_7353);
  not g20633 (n_7354, n13375);
  and g20634 (n13376, n_7344, n_7354);
  and g20635 (n13377, n_7322, n13339);
  and g20636 (n13378, n13336, n_7323);
  not g20637 (n_7355, n13377);
  not g20638 (n_7356, n13378);
  and g20639 (n13379, n_7355, n_7356);
  not g20640 (n_7357, n13376);
  not g20641 (n_7358, n13379);
  and g20642 (n13380, n_7357, n_7358);
  and g20643 (n13381, n13365, n_7354);
  and g20644 (n13382, n_7353, n_7354);
  not g20645 (n_7359, n13381);
  not g20646 (n_7360, n13382);
  and g20647 (n13383, n_7359, n_7360);
  and g20648 (n13384, n_7174, n_7177);
  and g20649 (n13385, n_7340, n_7341);
  and g20650 (n13386, n13360, n_7341);
  not g20651 (n_7361, n13385);
  not g20652 (n_7362, n13386);
  and g20653 (n13387, n_7361, n_7362);
  not g20654 (n_7363, n13384);
  not g20655 (n_7364, n13387);
  and g20656 (n13388, n_7363, n_7364);
  not g20657 (n_7365, n13388);
  and g20658 (n13389, n_7363, n_7365);
  and g20659 (n13390, n_7364, n_7365);
  not g20660 (n_7366, n13389);
  not g20661 (n_7367, n13390);
  and g20662 (n13391, n_7366, n_7367);
  and g20663 (n13392, n3457, n_712);
  and g20664 (n13393, n3542, n_566);
  and g20665 (n13394, n3606, n_560);
  and g20671 (n13397, n3368, n4715);
  not g20674 (n_7372, n13398);
  and g20675 (n13399, \a[29] , n_7372);
  not g20676 (n_7373, n13399);
  and g20677 (n13400, \a[29] , n_7373);
  and g20678 (n13401, n_7372, n_7373);
  not g20679 (n_7374, n13400);
  not g20680 (n_7375, n13401);
  and g20681 (n13402, n_7374, n_7375);
  not g20682 (n_7376, n13391);
  not g20683 (n_7377, n13402);
  and g20684 (n13403, n_7376, n_7377);
  not g20685 (n_7378, n13403);
  and g20686 (n13404, n_7365, n_7378);
  not g20687 (n_7379, n13383);
  not g20688 (n_7380, n13404);
  and g20689 (n13405, n_7379, n_7380);
  and g20690 (n13406, n13383, n13404);
  not g20691 (n_7381, n13405);
  not g20692 (n_7382, n13406);
  and g20693 (n13407, n_7381, n_7382);
  and g20694 (n13408, n_7376, n_7378);
  and g20695 (n13409, n_7377, n_7378);
  not g20696 (n_7383, n13408);
  not g20697 (n_7384, n13409);
  and g20698 (n13410, n_7383, n_7384);
  and g20699 (n13411, n_7195, n_7200);
  not g20700 (n_7385, n13410);
  not g20701 (n_7386, n13411);
  and g20702 (n13412, n_7385, n_7386);
  not g20703 (n_7387, n13412);
  and g20704 (n13413, n_7385, n_7387);
  and g20705 (n13414, n_7386, n_7387);
  not g20706 (n_7388, n13413);
  not g20707 (n_7389, n13414);
  and g20708 (n13415, n_7388, n_7389);
  and g20709 (n13416, n_7204, n_7208);
  not g20710 (n_7390, n13415);
  not g20711 (n_7391, n13416);
  and g20712 (n13417, n_7390, n_7391);
  not g20713 (n_7392, n13417);
  and g20714 (n13418, n_7387, n_7392);
  not g20715 (n_7393, n13418);
  and g20716 (n13419, n13407, n_7393);
  not g20717 (n_7394, n13419);
  and g20718 (n13420, n_7381, n_7394);
  and g20719 (n13421, n13376, n13379);
  not g20720 (n_7395, n13380);
  not g20721 (n_7396, n13421);
  and g20722 (n13422, n_7395, n_7396);
  not g20723 (n_7397, n13420);
  and g20724 (n13423, n_7397, n13422);
  not g20725 (n_7398, n13423);
  and g20726 (n13424, n_7395, n_7398);
  not g20727 (n_7399, n13343);
  and g20728 (n13425, n13341, n_7399);
  not g20729 (n_7400, n13344);
  not g20730 (n_7401, n13425);
  and g20731 (n13426, n_7400, n_7401);
  not g20732 (n_7402, n13424);
  and g20733 (n13427, n_7402, n13426);
  not g20734 (n_7403, n13427);
  and g20735 (n13428, n_7400, n_7403);
  not g20736 (n_7404, n13428);
  and g20737 (n13429, n13318, n_7404);
  not g20738 (n_7405, n13429);
  and g20739 (n13430, n_7303, n_7405);
  not g20740 (n_7406, n13430);
  and g20741 (n13431, n13190, n_7406);
  not g20742 (n_7407, n13431);
  and g20743 (n13432, n_7267, n_7407);
  not g20744 (n_7408, n13109);
  not g20745 (n_7409, n13432);
  and g20746 (n13433, n_7408, n_7409);
  not g20747 (n_7410, n13433);
  and g20748 (n13434, n_7247, n_7410);
  and g20749 (n13435, n13059, n_7243);
  not g20750 (n_7411, n13434);
  not g20751 (n_7412, n13435);
  and g20752 (n13436, n_7411, n_7412);
  not g20753 (n_7413, n13083);
  and g20754 (n13437, n_7413, n13436);
  and g20755 (n13438, n_7233, n13437);
  not g20756 (n_7414, n5407);
  not g20757 (n_7415, n5496);
  and g20758 (n13439, n_7414, n_7415);
  not g20759 (n_7416, n4935);
  and g20760 (n13440, n_7416, n13439);
  and g20761 (n13441, n_1011, n13440);
  not g20762 (n_7417, n13438);
  not g20763 (n_7418, n13441);
  and g20764 (n13442, n_7417, n_7418);
  not g20765 (n_7419, n13442);
  and g20766 (n13443, \a[20] , n_7419);
  and g20767 (n13444, n_435, n13442);
  not g20768 (n_7420, n13443);
  not g20769 (n_7421, n13444);
  and g20770 (n13445, n_7420, n_7421);
  and g20800 (n13475, n12958, n13474);
  not g20801 (n_7422, n13474);
  and g20802 (n13476, n_7222, n_7422);
  not g20803 (n_7423, n13475);
  not g20804 (n_7424, n13476);
  and g20805 (n13477, n_7423, n_7424);
  and g20806 (n13478, n13445, n13477);
  not g20807 (n_7425, n13445);
  not g20808 (n_7426, n13477);
  and g20809 (n13479, n_7425, n_7426);
  not g20810 (n_7427, n13478);
  not g20811 (n_7428, n13479);
  and g20812 (n13480, n_7427, n_7428);
  not g20813 (n_7429, n13009);
  and g20814 (n13481, n_7429, n13480);
  not g20815 (n_7430, n13480);
  and g20816 (n13482, n13009, n_7430);
  not g20817 (n_7431, n13481);
  not g20818 (n_7432, n13482);
  and g20819 (n13483, n_7431, n_7432);
  not g20820 (n_7433, n12902);
  and g20821 (n13484, n_7433, n13483);
  not g20822 (n_7434, n13484);
  and g20823 (n13485, n_7431, n_7434);
  and g20824 (n13486, n_7424, n_7427);
  not g20825 (n_7435, n13486);
  and g20826 (n13487, n13031, n_7435);
  not g20827 (n_7436, n13031);
  and g20828 (n13488, n_7436, n13486);
  not g20829 (n_7437, n13487);
  not g20830 (n_7438, n13488);
  and g20831 (n13489, n_7437, n_7438);
  and g20832 (n13490, n13415, n13416);
  not g20833 (n_7439, n13490);
  and g20834 (n13491, n_7392, n_7439);
  and g20835 (n13492, n3020, n13491);
  and g20836 (n13493, n3028, n12889);
  and g20837 (n13494, n3023, n12769);
  and g20838 (n13495, n_7212, n_7215);
  and g20839 (n13496, n12889, n13491);
  not g20840 (n_7440, n13491);
  and g20841 (n13497, n_7210, n_7440);
  not g20842 (n_7441, n13495);
  not g20843 (n_7442, n13497);
  and g20844 (n13498, n_7441, n_7442);
  not g20845 (n_7443, n13496);
  and g20846 (n13499, n_7443, n13498);
  not g20847 (n_7444, n13499);
  and g20848 (n13500, n_7441, n_7444);
  and g20849 (n13501, n_7443, n_7444);
  and g20850 (n13502, n_7442, n13501);
  not g20851 (n_7445, n13500);
  not g20852 (n_7446, n13502);
  and g20853 (n13503, n_7445, n_7446);
  not g20854 (n_7447, n13503);
  and g20855 (n13504, n75, n_7447);
  not g20863 (n_7452, n13507);
  and g20864 (n13508, n13489, n_7452);
  not g20865 (n_7453, n13489);
  and g20866 (n13509, n_7453, n13507);
  not g20867 (n_7454, n13508);
  not g20868 (n_7455, n13509);
  and g20869 (n13510, n_7454, n_7455);
  not g20870 (n_7456, n13485);
  and g20871 (n13511, n_7456, n13510);
  not g20872 (n_7457, n13510);
  and g20873 (n13512, n13485, n_7457);
  not g20874 (n_7458, n13511);
  not g20875 (n_7459, n13512);
  and g20876 (n13513, n_7458, n_7459);
  not g20877 (n_7460, n13426);
  and g20878 (n13514, n13424, n_7460);
  not g20879 (n_7461, n13514);
  and g20880 (n13515, n_7403, n_7461);
  and g20881 (n13516, n3457, n13515);
  not g20882 (n_7462, n13407);
  and g20883 (n13517, n_7462, n13418);
  not g20884 (n_7463, n13517);
  and g20885 (n13518, n_7394, n_7463);
  and g20886 (n13519, n3542, n13518);
  not g20887 (n_7464, n13422);
  and g20888 (n13520, n13420, n_7464);
  not g20889 (n_7465, n13520);
  and g20890 (n13521, n_7398, n_7465);
  and g20891 (n13522, n3606, n13521);
  not g20892 (n_7466, n13519);
  not g20893 (n_7467, n13522);
  and g20894 (n13523, n_7466, n_7467);
  not g20895 (n_7468, n13516);
  and g20896 (n13524, n_7468, n13523);
  and g20897 (n13525, n_489, n13524);
  and g20898 (n13526, n13518, n13521);
  and g20899 (n13527, n13491, n13518);
  not g20900 (n_7469, n13518);
  and g20901 (n13528, n_7440, n_7469);
  not g20902 (n_7470, n13527);
  not g20903 (n_7471, n13528);
  and g20904 (n13529, n_7470, n_7471);
  not g20905 (n_7472, n13501);
  and g20906 (n13530, n_7472, n13529);
  not g20907 (n_7473, n13530);
  and g20908 (n13531, n_7470, n_7473);
  not g20909 (n_7474, n13521);
  and g20910 (n13532, n_7469, n_7474);
  not g20911 (n_7475, n13531);
  not g20912 (n_7476, n13532);
  and g20913 (n13533, n_7475, n_7476);
  not g20914 (n_7477, n13526);
  and g20915 (n13534, n_7477, n13533);
  not g20916 (n_7478, n13534);
  and g20917 (n13535, n_7477, n_7478);
  not g20918 (n_7479, n13515);
  and g20919 (n13536, n_7479, n_7474);
  and g20920 (n13537, n13515, n13521);
  not g20921 (n_7480, n13536);
  not g20922 (n_7481, n13537);
  and g20923 (n13538, n_7480, n_7481);
  not g20924 (n_7482, n13535);
  and g20925 (n13539, n_7482, n13538);
  not g20926 (n_7483, n13538);
  and g20927 (n13540, n13535, n_7483);
  not g20928 (n_7484, n13539);
  not g20929 (n_7485, n13540);
  and g20930 (n13541, n_7484, n_7485);
  not g20931 (n_7486, n13541);
  and g20932 (n13542, n13524, n_7486);
  not g20933 (n_7487, n13525);
  not g20934 (n_7488, n13542);
  and g20935 (n13543, n_7487, n_7488);
  not g20936 (n_7489, n13543);
  and g20937 (n13544, \a[29] , n_7489);
  and g20938 (n13545, n_15, n13543);
  not g20939 (n_7490, n13544);
  not g20940 (n_7491, n13545);
  and g20941 (n13546, n_7490, n_7491);
  not g20942 (n_7492, n13546);
  and g20943 (n13547, n13513, n_7492);
  not g20944 (n_7493, n13547);
  and g20945 (n13548, n_7458, n_7493);
  and g20946 (n13549, n_7437, n_7454);
  and g20972 (n13575, n_7436, n13574);
  not g20973 (n_7494, n13574);
  and g20974 (n13576, n13031, n_7494);
  not g20975 (n_7495, n13549);
  not g20976 (n_7496, n13576);
  and g20977 (n13577, n_7495, n_7496);
  not g20978 (n_7497, n13575);
  and g20979 (n13578, n_7497, n13577);
  not g20980 (n_7498, n13578);
  and g20981 (n13579, n_7495, n_7498);
  and g20982 (n13580, n_7497, n_7498);
  and g20983 (n13581, n_7496, n13580);
  not g20984 (n_7499, n13579);
  not g20985 (n_7500, n13581);
  and g20986 (n13582, n_7499, n_7500);
  not g20987 (n_7501, n13529);
  and g20988 (n13583, n13501, n_7501);
  not g20989 (n_7502, n13583);
  and g20990 (n13584, n_7473, n_7502);
  and g20991 (n13585, n75, n13584);
  and g20992 (n13586, n3020, n13518);
  and g20993 (n13587, n3023, n12889);
  and g20994 (n13588, n3028, n13491);
  not g21002 (n_7507, n13582);
  not g21003 (n_7508, n13591);
  and g21004 (n13592, n_7507, n_7508);
  not g21005 (n_7509, n13592);
  and g21006 (n13593, n_7507, n_7509);
  and g21007 (n13594, n_7508, n_7509);
  not g21008 (n_7510, n13593);
  not g21009 (n_7511, n13594);
  and g21010 (n13595, n_7510, n_7511);
  not g21011 (n_7512, n13318);
  and g21012 (n13596, n_7512, n13428);
  not g21013 (n_7513, n13596);
  and g21014 (n13597, n_7405, n_7513);
  and g21015 (n13598, n3457, n13597);
  and g21016 (n13599, n3542, n13521);
  and g21017 (n13600, n3606, n13515);
  not g21018 (n_7514, n13599);
  not g21019 (n_7515, n13600);
  and g21020 (n13601, n_7514, n_7515);
  not g21021 (n_7516, n13598);
  and g21022 (n13602, n_7516, n13601);
  and g21023 (n13603, n_489, n13602);
  and g21024 (n13604, n_7481, n_7484);
  and g21025 (n13605, n13515, n13597);
  not g21026 (n_7517, n13597);
  and g21027 (n13606, n_7479, n_7517);
  not g21028 (n_7518, n13604);
  not g21029 (n_7519, n13606);
  and g21030 (n13607, n_7518, n_7519);
  not g21031 (n_7520, n13605);
  and g21032 (n13608, n_7520, n13607);
  not g21033 (n_7521, n13608);
  and g21034 (n13609, n_7518, n_7521);
  and g21035 (n13610, n_7520, n_7521);
  and g21036 (n13611, n_7519, n13610);
  not g21037 (n_7522, n13609);
  not g21038 (n_7523, n13611);
  and g21039 (n13612, n_7522, n_7523);
  and g21040 (n13613, n13602, n13612);
  not g21041 (n_7524, n13603);
  not g21042 (n_7525, n13613);
  and g21043 (n13614, n_7524, n_7525);
  not g21044 (n_7526, n13614);
  and g21045 (n13615, \a[29] , n_7526);
  and g21046 (n13616, n_15, n13614);
  not g21047 (n_7527, n13615);
  not g21048 (n_7528, n13616);
  and g21049 (n13617, n_7527, n_7528);
  not g21050 (n_7529, n13595);
  not g21051 (n_7530, n13617);
  and g21052 (n13618, n_7529, n_7530);
  and g21053 (n13619, n13595, n13617);
  not g21054 (n_7531, n13618);
  not g21055 (n_7532, n13619);
  and g21056 (n13620, n_7531, n_7532);
  not g21057 (n_7533, n13548);
  and g21058 (n13621, n_7533, n13620);
  not g21059 (n_7534, n13620);
  and g21060 (n13622, n13548, n_7534);
  not g21061 (n_7535, n13621);
  not g21062 (n_7536, n13622);
  and g21063 (n13623, n_7535, n_7536);
  not g21064 (n_7537, n13437);
  and g21065 (n13624, n_7411, n_7537);
  and g21066 (n13625, n_7412, n_7537);
  and g21067 (n13626, n_7413, n13625);
  not g21068 (n_7538, n13624);
  not g21069 (n_7539, n13626);
  and g21070 (n13627, n_7538, n_7539);
  not g21071 (n_7540, n13627);
  and g21072 (n13628, n3884, n_7540);
  not g21073 (n_7541, n13190);
  and g21074 (n13629, n_7541, n13430);
  not g21075 (n_7542, n13629);
  and g21076 (n13630, n_7407, n_7542);
  and g21077 (n13631, n3967, n13630);
  and g21078 (n13632, n13109, n13432);
  not g21079 (n_7543, n13632);
  and g21080 (n13633, n_7410, n_7543);
  and g21081 (n13634, n4046, n13633);
  and g21087 (n13637, n13630, n13633);
  and g21088 (n13638, n13597, n13630);
  not g21089 (n_7547, n13630);
  and g21090 (n13639, n_7517, n_7547);
  not g21091 (n_7548, n13638);
  not g21092 (n_7549, n13639);
  and g21093 (n13640, n_7548, n_7549);
  not g21094 (n_7550, n13610);
  and g21095 (n13641, n_7550, n13640);
  not g21096 (n_7551, n13641);
  and g21097 (n13642, n_7548, n_7551);
  not g21098 (n_7552, n13633);
  and g21099 (n13643, n_7547, n_7552);
  not g21100 (n_7553, n13637);
  not g21101 (n_7554, n13643);
  and g21102 (n13644, n_7553, n_7554);
  not g21103 (n_7555, n13642);
  and g21104 (n13645, n_7555, n13644);
  not g21105 (n_7556, n13645);
  and g21106 (n13646, n_7553, n_7556);
  and g21107 (n13647, n_7540, n13633);
  and g21108 (n13648, n13627, n_7552);
  not g21109 (n_7557, n13646);
  not g21110 (n_7558, n13648);
  and g21111 (n13649, n_7557, n_7558);
  not g21112 (n_7559, n13647);
  and g21113 (n13650, n_7559, n13649);
  not g21114 (n_7560, n13650);
  and g21115 (n13651, n_7557, n_7560);
  and g21116 (n13652, n_7559, n_7560);
  and g21117 (n13653, n_7558, n13652);
  not g21118 (n_7561, n13651);
  not g21119 (n_7562, n13653);
  and g21120 (n13654, n_7561, n_7562);
  not g21121 (n_7563, n13654);
  and g21122 (n13655, n4050, n_7563);
  not g21125 (n_7565, n13656);
  and g21126 (n13657, \a[26] , n_7565);
  not g21127 (n_7566, n13657);
  and g21128 (n13658, \a[26] , n_7566);
  and g21129 (n13659, n_7565, n_7566);
  not g21130 (n_7567, n13658);
  not g21131 (n_7568, n13659);
  and g21132 (n13660, n_7567, n_7568);
  not g21133 (n_7569, n13660);
  and g21134 (n13661, n13623, n_7569);
  not g21135 (n_7570, n13661);
  and g21136 (n13662, n13623, n_7570);
  and g21137 (n13663, n_7569, n_7570);
  not g21138 (n_7571, n13662);
  not g21139 (n_7572, n13663);
  and g21140 (n13664, n_7571, n_7572);
  and g21141 (n13665, n13483, n_7434);
  and g21142 (n13666, n_7433, n_7434);
  not g21143 (n_7573, n13665);
  not g21144 (n_7574, n13666);
  and g21145 (n13667, n_7573, n_7574);
  and g21146 (n13668, n_7230, n_7232);
  and g21147 (n13669, n_7231, n13009);
  not g21148 (n_7575, n13668);
  not g21149 (n_7576, n13669);
  and g21150 (n13670, n_7575, n_7576);
  and g21151 (n13671, n_146, n_157);
  and g21179 (n13699, n421, n_249);
  and g21180 (n13700, n_238, n13699);
  not g21196 (n_7577, n13695);
  not g21197 (n_7578, n13715);
  and g21198 (n13716, n_7577, n_7578);
  not g21199 (n_7579, n5939);
  not g21200 (n_7580, n6233);
  and g21201 (n13717, n_7579, n_7580);
  not g21202 (n_7581, n5663);
  and g21203 (n13718, n_7581, n13717);
  and g21204 (n13719, n_1409, n13718);
  not g21205 (n_7582, n13719);
  and g21206 (n13720, n_7417, n_7582);
  not g21207 (n_7583, n13720);
  and g21208 (n13721, \a[17] , n_7583);
  and g21209 (n13722, n_617, n13720);
  not g21210 (n_7584, n13721);
  not g21211 (n_7585, n13722);
  and g21212 (n13723, n_7584, n_7585);
  and g21213 (n13724, n13695, n13715);
  not g21214 (n_7586, n13716);
  not g21215 (n_7587, n13724);
  and g21216 (n13725, n_7586, n_7587);
  and g21217 (n13726, n13723, n13725);
  not g21218 (n_7588, n13726);
  and g21219 (n13727, n_7586, n_7588);
  not g21220 (n_7589, n13727);
  and g21221 (n13728, n12958, n_7589);
  and g21222 (n13729, n_7222, n13727);
  not g21223 (n_7590, n13728);
  not g21224 (n_7591, n13729);
  and g21225 (n13730, n_7590, n_7591);
  and g21226 (n13731, n3020, n12502);
  and g21227 (n13732, n3028, n12370);
  and g21228 (n13733, n3023, n12505);
  and g21229 (n13734, n_7100, n_7103);
  and g21230 (n13735, n_7101, n12684);
  not g21231 (n_7592, n13734);
  not g21232 (n_7593, n13735);
  and g21233 (n13736, n_7592, n_7593);
  not g21234 (n_7594, n13736);
  and g21235 (n13737, n75, n_7594);
  not g21243 (n_7599, n13740);
  and g21244 (n13741, n13730, n_7599);
  not g21245 (n_7600, n13741);
  and g21246 (n13742, n_7590, n_7600);
  not g21247 (n_7601, n13670);
  not g21248 (n_7602, n13742);
  and g21249 (n13743, n_7601, n_7602);
  and g21250 (n13744, n13670, n13742);
  not g21251 (n_7603, n13743);
  not g21252 (n_7604, n13744);
  and g21253 (n13745, n_7603, n_7604);
  and g21254 (n13746, n_7095, n_7098);
  and g21255 (n13747, n_7096, n12680);
  not g21256 (n_7605, n13746);
  not g21257 (n_7606, n13747);
  and g21258 (n13748, n_7605, n_7606);
  not g21259 (n_7607, n13748);
  and g21260 (n13749, n75, n_7607);
  and g21261 (n13750, n3020, n12370);
  and g21262 (n13751, n3023, n12508);
  and g21263 (n13752, n3028, n12505);
  not g21271 (n_7612, n13723);
  not g21272 (n_7613, n13725);
  and g21273 (n13756, n_7612, n_7613);
  not g21274 (n_7614, n13756);
  and g21275 (n13757, n_7588, n_7614);
  not g21276 (n_7615, n13755);
  and g21277 (n13758, n_7615, n13757);
  and g21293 (n13774, n_44, n_84);
  and g21307 (n13788, n2683, n13787);
  and g21308 (n13789, n_60, n13788);
  not g21325 (n_7616, n13805);
  and g21326 (n13806, n13695, n_7616);
  and g21327 (n13807, n_47, n5082);
  and g21328 (n13808, n_278, n13807);
  and g21347 (n13827, n773, n1528);
  not g21364 (n_7617, n13821);
  not g21365 (n_7618, n13843);
  and g21366 (n13844, n_7617, n_7618);
  not g21367 (n_7619, n6951);
  not g21368 (n_7620, n7101);
  and g21369 (n13845, n_7619, n_7620);
  not g21370 (n_7621, n6402);
  and g21371 (n13846, n_7621, n13845);
  and g21372 (n13847, n_1885, n13846);
  not g21373 (n_7622, n13847);
  and g21374 (n13848, n_7417, n_7622);
  not g21375 (n_7623, n13848);
  and g21376 (n13849, \a[14] , n_7623);
  and g21377 (n13850, n_652, n13848);
  not g21378 (n_7624, n13849);
  not g21379 (n_7625, n13850);
  and g21380 (n13851, n_7624, n_7625);
  and g21381 (n13852, n13821, n13843);
  not g21382 (n_7626, n13844);
  not g21383 (n_7627, n13852);
  and g21384 (n13853, n_7626, n_7627);
  and g21385 (n13854, n13851, n13853);
  not g21386 (n_7628, n13854);
  and g21387 (n13855, n_7626, n_7628);
  not g21388 (n_7629, n13855);
  and g21389 (n13856, n13805, n_7629);
  and g21390 (n13857, n_7616, n13855);
  not g21391 (n_7630, n13856);
  not g21392 (n_7631, n13857);
  and g21393 (n13858, n_7630, n_7631);
  and g21394 (n13859, n3020, n12508);
  and g21395 (n13860, n3028, n12513);
  and g21396 (n13861, n3023, n12511);
  not g21397 (n_7632, n12670);
  and g21398 (n13862, n12667, n_7632);
  not g21399 (n_7633, n13862);
  and g21400 (n13863, n_7088, n_7633);
  and g21401 (n13864, n75, n13863);
  not g21409 (n_7638, n13867);
  and g21410 (n13868, n13858, n_7638);
  not g21411 (n_7639, n13868);
  and g21412 (n13869, n_7630, n_7639);
  and g21413 (n13870, n_7577, n13805);
  not g21414 (n_7640, n13869);
  not g21415 (n_7641, n13870);
  and g21416 (n13871, n_7640, n_7641);
  not g21417 (n_7642, n13806);
  and g21418 (n13872, n_7642, n13871);
  not g21419 (n_7643, n13872);
  and g21420 (n13873, n_7642, n_7643);
  not g21421 (n_7644, n13758);
  and g21422 (n13874, n13757, n_7644);
  and g21423 (n13875, n_7615, n_7644);
  not g21424 (n_7645, n13874);
  not g21425 (n_7646, n13875);
  and g21426 (n13876, n_7645, n_7646);
  not g21427 (n_7647, n13873);
  not g21428 (n_7648, n13876);
  and g21429 (n13877, n_7647, n_7648);
  not g21430 (n_7649, n13877);
  and g21431 (n13878, n_7644, n_7649);
  not g21432 (n_7650, n13730);
  and g21433 (n13879, n_7650, n13740);
  not g21434 (n_7651, n13879);
  and g21435 (n13880, n_7600, n_7651);
  not g21436 (n_7652, n13878);
  and g21437 (n13881, n_7652, n13880);
  not g21438 (n_7653, n13880);
  and g21439 (n13882, n13878, n_7653);
  not g21440 (n_7654, n13881);
  not g21441 (n_7655, n13882);
  and g21442 (n13883, n_7654, n_7655);
  and g21443 (n13884, n3457, n13491);
  and g21444 (n13885, n3542, n12769);
  and g21445 (n13886, n3606, n12889);
  not g21446 (n_7656, n13885);
  not g21447 (n_7657, n13886);
  and g21448 (n13887, n_7656, n_7657);
  not g21449 (n_7658, n13884);
  and g21450 (n13888, n_7658, n13887);
  and g21451 (n13889, n_489, n13888);
  and g21452 (n13890, n13503, n13888);
  not g21453 (n_7659, n13889);
  not g21454 (n_7660, n13890);
  and g21455 (n13891, n_7659, n_7660);
  not g21456 (n_7661, n13891);
  and g21457 (n13892, \a[29] , n_7661);
  and g21458 (n13893, n_15, n13891);
  not g21459 (n_7662, n13892);
  not g21460 (n_7663, n13893);
  and g21461 (n13894, n_7662, n_7663);
  not g21462 (n_7664, n13894);
  and g21463 (n13895, n13883, n_7664);
  not g21464 (n_7665, n13895);
  and g21465 (n13896, n_7654, n_7665);
  not g21466 (n_7666, n13896);
  and g21467 (n13897, n13745, n_7666);
  not g21468 (n_7667, n13897);
  and g21469 (n13898, n_7603, n_7667);
  not g21470 (n_7668, n13667);
  not g21471 (n_7669, n13898);
  and g21472 (n13899, n_7668, n_7669);
  and g21473 (n13900, n13667, n13898);
  not g21474 (n_7670, n13899);
  not g21475 (n_7671, n13900);
  and g21476 (n13901, n_7670, n_7671);
  and g21477 (n13902, n3457, n13521);
  and g21478 (n13903, n3542, n13491);
  and g21479 (n13904, n3606, n13518);
  and g21485 (n13907, n_7475, n_7478);
  and g21486 (n13908, n_7476, n13535);
  not g21487 (n_7675, n13907);
  not g21488 (n_7676, n13908);
  and g21489 (n13909, n_7675, n_7676);
  not g21490 (n_7677, n13909);
  and g21491 (n13910, n3368, n_7677);
  not g21494 (n_7679, n13911);
  and g21495 (n13912, \a[29] , n_7679);
  not g21496 (n_7680, n13912);
  and g21497 (n13913, \a[29] , n_7680);
  and g21498 (n13914, n_7679, n_7680);
  not g21499 (n_7681, n13913);
  not g21500 (n_7682, n13914);
  and g21501 (n13915, n_7681, n_7682);
  not g21502 (n_7683, n13915);
  and g21503 (n13916, n13901, n_7683);
  not g21504 (n_7684, n13916);
  and g21505 (n13917, n_7670, n_7684);
  not g21506 (n_7685, n13513);
  and g21507 (n13918, n_7685, n13546);
  not g21508 (n_7686, n13918);
  and g21509 (n13919, n_7493, n_7686);
  not g21510 (n_7687, n13917);
  and g21511 (n13920, n_7687, n13919);
  not g21512 (n_7688, n13919);
  and g21513 (n13921, n13917, n_7688);
  not g21514 (n_7689, n13920);
  not g21515 (n_7690, n13921);
  and g21516 (n13922, n_7689, n_7690);
  and g21517 (n13923, n3884, n13633);
  and g21518 (n13924, n3967, n13597);
  and g21519 (n13925, n4046, n13630);
  not g21525 (n_7694, n13644);
  and g21526 (n13928, n13642, n_7694);
  not g21527 (n_7695, n13928);
  and g21528 (n13929, n_7556, n_7695);
  and g21529 (n13930, n4050, n13929);
  not g21532 (n_7697, n13931);
  and g21533 (n13932, \a[26] , n_7697);
  not g21534 (n_7698, n13932);
  and g21535 (n13933, \a[26] , n_7698);
  and g21536 (n13934, n_7697, n_7698);
  not g21537 (n_7699, n13933);
  not g21538 (n_7700, n13934);
  and g21539 (n13935, n_7699, n_7700);
  not g21540 (n_7701, n13935);
  and g21541 (n13936, n13922, n_7701);
  not g21542 (n_7702, n13936);
  and g21543 (n13937, n_7689, n_7702);
  not g21544 (n_7703, n4604);
  not g21545 (n_7704, n4694);
  and g21546 (n13938, n_7703, n_7704);
  not g21547 (n_7705, n13938);
  and g21548 (n13939, n_7417, n_7705);
  and g21549 (n13940, n13059, n13625);
  not g21550 (n_7706, n13940);
  and g21551 (n13941, n_7417, n_7706);
  and g21552 (n13942, n4533, n13941);
  not g21553 (n_7707, n13939);
  not g21554 (n_7708, n13942);
  and g21555 (n13943, n_7707, n_7708);
  and g21556 (n13944, n_732, n13943);
  and g21557 (n13945, n_7540, n13941);
  not g21558 (n_7709, n13941);
  and g21559 (n13946, n13627, n_7709);
  not g21560 (n_7710, n13945);
  not g21561 (n_7711, n13946);
  and g21562 (n13947, n_7710, n_7711);
  not g21563 (n_7712, n13652);
  and g21564 (n13948, n_7712, n13947);
  not g21565 (n_7713, n13948);
  and g21566 (n13949, n_7710, n_7713);
  not g21567 (n_7714, n13949);
  and g21568 (n13950, n13940, n_7714);
  not g21569 (n_7715, n13950);
  and g21570 (n13951, n_7709, n_7715);
  and g21571 (n13952, n13943, n13951);
  not g21572 (n_7716, n13944);
  not g21573 (n_7717, n13952);
  and g21574 (n13953, n_7716, n_7717);
  not g21575 (n_7718, n13953);
  and g21576 (n13954, \a[23] , n_7718);
  and g21577 (n13955, n_27, n13953);
  not g21578 (n_7719, n13954);
  not g21579 (n_7720, n13955);
  and g21580 (n13956, n_7719, n_7720);
  not g21581 (n_7721, n13937);
  not g21582 (n_7722, n13956);
  and g21583 (n13957, n_7721, n_7722);
  and g21584 (n13958, n13937, n13956);
  not g21585 (n_7723, n13957);
  not g21586 (n_7724, n13958);
  and g21587 (n13959, n_7723, n_7724);
  not g21588 (n_7725, n13664);
  and g21589 (n13960, n_7725, n13959);
  not g21590 (n_7726, n13960);
  and g21591 (n13961, n_7725, n_7726);
  and g21592 (n13962, n13959, n_7726);
  not g21593 (n_7727, n13961);
  not g21594 (n_7728, n13962);
  and g21595 (n13963, n_7727, n_7728);
  and g21596 (n13964, n13922, n_7702);
  and g21597 (n13965, n_7701, n_7702);
  not g21598 (n_7729, n13964);
  not g21599 (n_7730, n13965);
  and g21600 (n13966, n_7729, n_7730);
  and g21601 (n13967, n13901, n_7684);
  and g21602 (n13968, n_7683, n_7684);
  not g21603 (n_7731, n13967);
  not g21604 (n_7732, n13968);
  and g21605 (n13969, n_7731, n_7732);
  and g21606 (n13970, n3884, n13630);
  and g21607 (n13971, n3967, n13515);
  and g21608 (n13972, n4046, n13597);
  not g21614 (n_7736, n13640);
  and g21615 (n13975, n13610, n_7736);
  not g21616 (n_7737, n13975);
  and g21617 (n13976, n_7551, n_7737);
  and g21618 (n13977, n4050, n13976);
  not g21621 (n_7739, n13978);
  and g21622 (n13979, \a[26] , n_7739);
  not g21623 (n_7740, n13979);
  and g21624 (n13980, \a[26] , n_7740);
  and g21625 (n13981, n_7739, n_7740);
  not g21626 (n_7741, n13980);
  not g21627 (n_7742, n13981);
  and g21628 (n13982, n_7741, n_7742);
  not g21629 (n_7743, n13969);
  not g21630 (n_7744, n13982);
  and g21631 (n13983, n_7743, n_7744);
  not g21632 (n_7745, n13983);
  and g21633 (n13984, n_7743, n_7745);
  and g21634 (n13985, n_7744, n_7745);
  not g21635 (n_7746, n13984);
  not g21636 (n_7747, n13985);
  and g21637 (n13986, n_7746, n_7747);
  not g21638 (n_7748, n13745);
  and g21639 (n13987, n_7748, n13896);
  not g21640 (n_7749, n13987);
  and g21641 (n13988, n_7667, n_7749);
  and g21642 (n13989, n3457, n13518);
  and g21643 (n13990, n3542, n12889);
  and g21644 (n13991, n3606, n13491);
  and g21650 (n13994, n3368, n13584);
  not g21653 (n_7754, n13995);
  and g21654 (n13996, \a[29] , n_7754);
  not g21655 (n_7755, n13996);
  and g21656 (n13997, \a[29] , n_7755);
  and g21657 (n13998, n_7754, n_7755);
  not g21658 (n_7756, n13997);
  not g21659 (n_7757, n13998);
  and g21660 (n13999, n_7756, n_7757);
  not g21661 (n_7758, n13999);
  and g21662 (n14000, n13988, n_7758);
  not g21663 (n_7759, n14000);
  and g21664 (n14001, n13988, n_7759);
  and g21665 (n14002, n_7758, n_7759);
  not g21666 (n_7760, n14001);
  not g21667 (n_7761, n14002);
  and g21668 (n14003, n_7760, n_7761);
  and g21669 (n14004, n3884, n13597);
  and g21670 (n14005, n3967, n13521);
  and g21671 (n14006, n4046, n13515);
  not g21677 (n_7765, n13612);
  and g21678 (n14009, n4050, n_7765);
  not g21681 (n_7767, n14010);
  and g21682 (n14011, \a[26] , n_7767);
  not g21683 (n_7768, n14011);
  and g21684 (n14012, \a[26] , n_7768);
  and g21685 (n14013, n_7767, n_7768);
  not g21686 (n_7769, n14012);
  not g21687 (n_7770, n14013);
  and g21688 (n14014, n_7769, n_7770);
  not g21689 (n_7771, n14003);
  not g21690 (n_7772, n14014);
  and g21691 (n14015, n_7771, n_7772);
  not g21692 (n_7773, n14015);
  and g21693 (n14016, n_7759, n_7773);
  not g21694 (n_7774, n13986);
  not g21695 (n_7775, n14016);
  and g21696 (n14017, n_7774, n_7775);
  not g21697 (n_7776, n14017);
  and g21698 (n14018, n_7745, n_7776);
  not g21699 (n_7777, n13966);
  not g21700 (n_7778, n14018);
  and g21701 (n14019, n_7777, n_7778);
  and g21702 (n14020, n13966, n14018);
  not g21703 (n_7779, n14019);
  not g21704 (n_7780, n14020);
  and g21705 (n14021, n_7779, n_7780);
  and g21706 (n14022, n4694, n_7417);
  and g21707 (n14023, n4533, n_7540);
  and g21708 (n14024, n4604, n13941);
  and g21714 (n14027, n_7706, n13949);
  not g21715 (n_7784, n14027);
  and g21716 (n14028, n_7715, n_7784);
  and g21717 (n14029, n4536, n14028);
  not g21720 (n_7786, n14030);
  and g21721 (n14031, \a[23] , n_7786);
  not g21722 (n_7787, n14031);
  and g21723 (n14032, \a[23] , n_7787);
  and g21724 (n14033, n_7786, n_7787);
  not g21725 (n_7788, n14032);
  not g21726 (n_7789, n14033);
  and g21727 (n14034, n_7788, n_7789);
  not g21728 (n_7790, n14034);
  and g21729 (n14035, n14021, n_7790);
  not g21730 (n_7791, n14035);
  and g21731 (n14036, n_7779, n_7791);
  not g21732 (n_7792, n13963);
  not g21733 (n_7793, n14036);
  and g21734 (n14037, n_7792, n_7793);
  and g21735 (n14038, n13963, n14036);
  not g21736 (n_7794, n14037);
  not g21737 (n_7795, n14038);
  and g21738 (n14039, n_7794, n_7795);
  and g21739 (n14040, n14021, n_7791);
  and g21740 (n14041, n_7790, n_7791);
  not g21741 (n_7796, n14040);
  not g21742 (n_7797, n14041);
  and g21743 (n14042, n_7796, n_7797);
  and g21744 (n14043, n_7771, n_7773);
  and g21745 (n14044, n_7772, n_7773);
  not g21746 (n_7798, n14043);
  not g21747 (n_7799, n14044);
  and g21748 (n14045, n_7798, n_7799);
  and g21749 (n14046, n_7640, n_7643);
  and g21750 (n14047, n_7641, n13873);
  not g21751 (n_7800, n14046);
  not g21752 (n_7801, n14047);
  and g21753 (n14048, n_7800, n_7801);
  and g21754 (n14049, n_7090, n_7093);
  and g21755 (n14050, n_7091, n12676);
  not g21756 (n_7802, n14049);
  not g21757 (n_7803, n14050);
  and g21758 (n14051, n_7802, n_7803);
  not g21759 (n_7804, n14051);
  and g21760 (n14052, n75, n_7804);
  and g21761 (n14053, n3020, n12505);
  and g21762 (n14054, n3023, n12513);
  and g21763 (n14055, n3028, n12508);
  not g21771 (n_7809, n14048);
  not g21772 (n_7810, n14058);
  and g21773 (n14059, n_7809, n_7810);
  not g21774 (n_7811, n14059);
  and g21775 (n14060, n_7809, n_7811);
  and g21776 (n14061, n_7810, n_7811);
  not g21777 (n_7812, n14060);
  not g21778 (n_7813, n14061);
  and g21779 (n14062, n_7812, n_7813);
  and g21780 (n14063, n3457, n12769);
  and g21781 (n14064, n3542, n12370);
  and g21782 (n14065, n3606, n12502);
  not g21783 (n_7814, n14064);
  not g21784 (n_7815, n14065);
  and g21785 (n14066, n_7814, n_7815);
  not g21786 (n_7816, n14063);
  and g21787 (n14067, n_7816, n14066);
  and g21788 (n14068, n_489, n14067);
  not g21789 (n_7817, n12999);
  and g21790 (n14069, n_7817, n14067);
  not g21791 (n_7818, n14068);
  not g21792 (n_7819, n14069);
  and g21793 (n14070, n_7818, n_7819);
  not g21794 (n_7820, n14070);
  and g21795 (n14071, \a[29] , n_7820);
  and g21796 (n14072, n_15, n14070);
  not g21797 (n_7821, n14071);
  not g21798 (n_7822, n14072);
  and g21799 (n14073, n_7821, n_7822);
  not g21800 (n_7823, n14062);
  not g21801 (n_7824, n14073);
  and g21802 (n14074, n_7823, n_7824);
  not g21803 (n_7825, n14074);
  and g21804 (n14075, n_7811, n_7825);
  and g21805 (n14076, n_7648, n_7649);
  and g21806 (n14077, n_7647, n_7649);
  not g21807 (n_7826, n14076);
  not g21808 (n_7827, n14077);
  and g21809 (n14078, n_7826, n_7827);
  not g21810 (n_7828, n14075);
  not g21811 (n_7829, n14078);
  and g21812 (n14079, n_7828, n_7829);
  not g21813 (n_7830, n14079);
  and g21814 (n14080, n_7828, n_7830);
  and g21815 (n14081, n_7829, n_7830);
  not g21816 (n_7831, n14080);
  not g21817 (n_7832, n14081);
  and g21818 (n14082, n_7831, n_7832);
  and g21819 (n14083, n3457, n12889);
  and g21820 (n14084, n3542, n12502);
  and g21821 (n14085, n3606, n12769);
  and g21827 (n14088, n3368, n12895);
  not g21830 (n_7837, n14089);
  and g21831 (n14090, \a[29] , n_7837);
  not g21832 (n_7838, n14090);
  and g21833 (n14091, \a[29] , n_7838);
  and g21834 (n14092, n_7837, n_7838);
  not g21835 (n_7839, n14091);
  not g21836 (n_7840, n14092);
  and g21837 (n14093, n_7839, n_7840);
  not g21838 (n_7841, n14082);
  not g21839 (n_7842, n14093);
  and g21840 (n14094, n_7841, n_7842);
  not g21841 (n_7843, n14094);
  and g21842 (n14095, n_7830, n_7843);
  not g21843 (n_7844, n13883);
  and g21844 (n14096, n_7844, n13894);
  not g21845 (n_7845, n14096);
  and g21846 (n14097, n_7665, n_7845);
  not g21847 (n_7846, n14095);
  and g21848 (n14098, n_7846, n14097);
  not g21849 (n_7847, n14097);
  and g21850 (n14099, n14095, n_7847);
  not g21851 (n_7848, n14098);
  not g21852 (n_7849, n14099);
  and g21853 (n14100, n_7848, n_7849);
  and g21854 (n14101, n3884, n13515);
  and g21855 (n14102, n3967, n13518);
  and g21856 (n14103, n4046, n13521);
  and g21862 (n14106, n4050, n13541);
  not g21865 (n_7854, n14107);
  and g21866 (n14108, \a[26] , n_7854);
  not g21867 (n_7855, n14108);
  and g21868 (n14109, \a[26] , n_7855);
  and g21869 (n14110, n_7854, n_7855);
  not g21870 (n_7856, n14109);
  not g21871 (n_7857, n14110);
  and g21872 (n14111, n_7856, n_7857);
  not g21873 (n_7858, n14111);
  and g21874 (n14112, n14100, n_7858);
  not g21875 (n_7859, n14112);
  and g21876 (n14113, n_7848, n_7859);
  not g21877 (n_7860, n14045);
  not g21878 (n_7861, n14113);
  and g21879 (n14114, n_7860, n_7861);
  and g21880 (n14115, n14045, n14113);
  not g21881 (n_7862, n14114);
  not g21882 (n_7863, n14115);
  and g21883 (n14116, n_7862, n_7863);
  and g21884 (n14117, n4694, n_7540);
  and g21885 (n14118, n4533, n13630);
  and g21886 (n14119, n4604, n13633);
  and g21892 (n14122, n4536, n_7563);
  not g21895 (n_7868, n14123);
  and g21896 (n14124, \a[23] , n_7868);
  not g21897 (n_7869, n14124);
  and g21898 (n14125, \a[23] , n_7869);
  and g21899 (n14126, n_7868, n_7869);
  not g21900 (n_7870, n14125);
  not g21901 (n_7871, n14126);
  and g21902 (n14127, n_7870, n_7871);
  not g21903 (n_7872, n14127);
  and g21904 (n14128, n14116, n_7872);
  not g21905 (n_7873, n14128);
  and g21906 (n14129, n_7862, n_7873);
  and g21907 (n14130, n4694, n13941);
  and g21908 (n14131, n4533, n13633);
  and g21909 (n14132, n4604, n_7540);
  not g21915 (n_7877, n13947);
  and g21916 (n14135, n13652, n_7877);
  not g21917 (n_7878, n14135);
  and g21918 (n14136, n_7713, n_7878);
  and g21919 (n14137, n4536, n14136);
  not g21922 (n_7880, n14138);
  and g21923 (n14139, \a[23] , n_7880);
  not g21924 (n_7881, n14139);
  and g21925 (n14140, \a[23] , n_7881);
  and g21926 (n14141, n_7880, n_7881);
  not g21927 (n_7882, n14140);
  not g21928 (n_7883, n14141);
  and g21929 (n14142, n_7882, n_7883);
  not g21930 (n_7884, n14129);
  not g21931 (n_7885, n14142);
  and g21932 (n14143, n_7884, n_7885);
  and g21933 (n14144, n13986, n14016);
  not g21934 (n_7886, n14144);
  and g21935 (n14145, n_7776, n_7886);
  not g21936 (n_7887, n14143);
  and g21937 (n14146, n_7884, n_7887);
  and g21938 (n14147, n_7885, n_7887);
  not g21939 (n_7888, n14146);
  not g21940 (n_7889, n14147);
  and g21941 (n14148, n_7888, n_7889);
  not g21942 (n_7890, n14148);
  and g21943 (n14149, n14145, n_7890);
  not g21944 (n_7891, n14149);
  and g21945 (n14150, n_7887, n_7891);
  not g21946 (n_7892, n14042);
  not g21947 (n_7893, n14150);
  and g21948 (n14151, n_7892, n_7893);
  not g21949 (n_7894, n14151);
  and g21950 (n14152, n_7892, n_7894);
  and g21951 (n14153, n_7893, n_7894);
  not g21952 (n_7895, n14152);
  not g21953 (n_7896, n14153);
  and g21954 (n14154, n_7895, n_7896);
  and g21955 (n14155, n14100, n_7859);
  and g21956 (n14156, n_7858, n_7859);
  not g21957 (n_7897, n14155);
  not g21958 (n_7898, n14156);
  and g21959 (n14157, n_7897, n_7898);
  and g21960 (n14158, n_7841, n_7843);
  and g21961 (n14159, n_7842, n_7843);
  not g21962 (n_7899, n14158);
  not g21963 (n_7900, n14159);
  and g21964 (n14160, n_7899, n_7900);
  and g21965 (n14161, n3884, n13521);
  and g21966 (n14162, n3967, n13491);
  and g21967 (n14163, n4046, n13518);
  and g21973 (n14166, n4050, n_7677);
  not g21976 (n_7905, n14167);
  and g21977 (n14168, \a[26] , n_7905);
  not g21978 (n_7906, n14168);
  and g21979 (n14169, \a[26] , n_7906);
  and g21980 (n14170, n_7905, n_7906);
  not g21981 (n_7907, n14169);
  not g21982 (n_7908, n14170);
  and g21983 (n14171, n_7907, n_7908);
  not g21984 (n_7909, n14160);
  not g21985 (n_7910, n14171);
  and g21986 (n14172, n_7909, n_7910);
  not g21987 (n_7911, n14172);
  and g21988 (n14173, n_7909, n_7911);
  and g21989 (n14174, n_7910, n_7911);
  not g21990 (n_7912, n14173);
  not g21991 (n_7913, n14174);
  and g21992 (n14175, n_7912, n_7913);
  not g21993 (n_7914, n12665);
  and g21994 (n14176, n12663, n_7914);
  not g21995 (n_7915, n14176);
  and g21996 (n14177, n_7083, n_7915);
  and g21997 (n14178, n75, n14177);
  and g21998 (n14179, n3020, n12513);
  and g21999 (n14180, n3023, n12516);
  and g22000 (n14181, n3028, n12511);
  not g22052 (n_7920, n14228);
  and g22053 (n14229, n13821, n_7920);
  and g22054 (n14230, n_7617, n14228);
  and g22055 (n14231, n_7075, n_7078);
  and g22056 (n14232, n_7076, n12663);
  not g22057 (n_7921, n14231);
  not g22058 (n_7922, n14232);
  and g22059 (n14233, n_7921, n_7922);
  not g22060 (n_7923, n14233);
  and g22061 (n14234, n75, n_7923);
  and g22062 (n14235, n3020, n12511);
  and g22063 (n14236, n3023, n12519);
  and g22064 (n14237, n3028, n12516);
  not g22072 (n_7928, n14229);
  not g22073 (n_7929, n14240);
  and g22074 (n14241, n_7928, n_7929);
  not g22075 (n_7930, n14230);
  and g22076 (n14242, n_7930, n14241);
  not g22077 (n_7931, n14242);
  and g22078 (n14243, n_7928, n_7931);
  not g22079 (n_7932, n13851);
  not g22080 (n_7933, n13853);
  and g22081 (n14244, n_7932, n_7933);
  not g22082 (n_7934, n14244);
  and g22083 (n14245, n_7628, n_7934);
  not g22084 (n_7935, n14243);
  and g22085 (n14246, n_7935, n14245);
  not g22086 (n_7936, n14245);
  and g22087 (n14247, n14243, n_7936);
  not g22088 (n_7937, n14246);
  not g22089 (n_7938, n14247);
  and g22090 (n14248, n_7937, n_7938);
  not g22091 (n_7939, n14184);
  and g22092 (n14249, n_7939, n14248);
  not g22093 (n_7940, n14249);
  and g22094 (n14250, n_7937, n_7940);
  not g22095 (n_7941, n13858);
  and g22096 (n14251, n_7941, n13867);
  not g22097 (n_7942, n14251);
  and g22098 (n14252, n_7639, n_7942);
  not g22099 (n_7943, n14250);
  and g22100 (n14253, n_7943, n14252);
  not g22101 (n_7944, n14252);
  and g22102 (n14254, n14250, n_7944);
  not g22103 (n_7945, n14253);
  not g22104 (n_7946, n14254);
  and g22105 (n14255, n_7945, n_7946);
  and g22106 (n14256, n3457, n12502);
  and g22107 (n14257, n3542, n12505);
  and g22108 (n14258, n3606, n12370);
  not g22109 (n_7947, n14257);
  not g22110 (n_7948, n14258);
  and g22111 (n14259, n_7947, n_7948);
  not g22112 (n_7949, n14256);
  and g22113 (n14260, n_7949, n14259);
  and g22114 (n14261, n_489, n14260);
  and g22115 (n14262, n13736, n14260);
  not g22116 (n_7950, n14261);
  not g22117 (n_7951, n14262);
  and g22118 (n14263, n_7950, n_7951);
  not g22119 (n_7952, n14263);
  and g22120 (n14264, \a[29] , n_7952);
  and g22121 (n14265, n_15, n14263);
  not g22122 (n_7953, n14264);
  not g22123 (n_7954, n14265);
  and g22124 (n14266, n_7953, n_7954);
  not g22125 (n_7955, n14266);
  and g22126 (n14267, n14255, n_7955);
  not g22127 (n_7956, n14267);
  and g22128 (n14268, n_7945, n_7956);
  and g22129 (n14269, n14062, n14073);
  not g22130 (n_7957, n14269);
  and g22131 (n14270, n_7825, n_7957);
  not g22132 (n_7958, n14268);
  and g22133 (n14271, n_7958, n14270);
  not g22134 (n_7959, n14270);
  and g22135 (n14272, n14268, n_7959);
  not g22136 (n_7960, n14271);
  not g22137 (n_7961, n14272);
  and g22138 (n14273, n_7960, n_7961);
  and g22139 (n14274, n3884, n13518);
  and g22140 (n14275, n3967, n12889);
  and g22141 (n14276, n4046, n13491);
  and g22147 (n14279, n4050, n13584);
  not g22150 (n_7966, n14280);
  and g22151 (n14281, \a[26] , n_7966);
  not g22152 (n_7967, n14281);
  and g22153 (n14282, \a[26] , n_7967);
  and g22154 (n14283, n_7966, n_7967);
  not g22155 (n_7968, n14282);
  not g22156 (n_7969, n14283);
  and g22157 (n14284, n_7968, n_7969);
  not g22158 (n_7970, n14284);
  and g22159 (n14285, n14273, n_7970);
  not g22160 (n_7971, n14285);
  and g22161 (n14286, n_7960, n_7971);
  not g22162 (n_7972, n14175);
  not g22163 (n_7973, n14286);
  and g22164 (n14287, n_7972, n_7973);
  not g22165 (n_7974, n14287);
  and g22166 (n14288, n_7911, n_7974);
  not g22167 (n_7975, n14157);
  not g22168 (n_7976, n14288);
  and g22169 (n14289, n_7975, n_7976);
  and g22170 (n14290, n14157, n14288);
  not g22171 (n_7977, n14289);
  not g22172 (n_7978, n14290);
  and g22173 (n14291, n_7977, n_7978);
  and g22174 (n14292, n4694, n13633);
  and g22175 (n14293, n4533, n13597);
  and g22176 (n14294, n4604, n13630);
  and g22182 (n14297, n4536, n13929);
  not g22185 (n_7983, n14298);
  and g22186 (n14299, \a[23] , n_7983);
  not g22187 (n_7984, n14299);
  and g22188 (n14300, \a[23] , n_7984);
  and g22189 (n14301, n_7983, n_7984);
  not g22190 (n_7985, n14300);
  not g22191 (n_7986, n14301);
  and g22192 (n14302, n_7985, n_7986);
  not g22193 (n_7987, n14302);
  and g22194 (n14303, n14291, n_7987);
  not g22195 (n_7988, n14303);
  and g22196 (n14304, n_7977, n_7988);
  not g22197 (n_7989, n13439);
  and g22198 (n14305, n_7417, n_7989);
  and g22199 (n14306, n4935, n13941);
  not g22200 (n_7990, n14305);
  not g22201 (n_7991, n14306);
  and g22202 (n14307, n_7990, n_7991);
  and g22203 (n14308, n_1011, n14307);
  and g22204 (n14309, n13951, n14307);
  not g22205 (n_7992, n14308);
  not g22206 (n_7993, n14309);
  and g22207 (n14310, n_7992, n_7993);
  not g22208 (n_7994, n14310);
  and g22209 (n14311, \a[20] , n_7994);
  and g22210 (n14312, n_435, n14310);
  not g22211 (n_7995, n14311);
  not g22212 (n_7996, n14312);
  and g22213 (n14313, n_7995, n_7996);
  not g22214 (n_7997, n14304);
  not g22215 (n_7998, n14313);
  and g22216 (n14314, n_7997, n_7998);
  and g22217 (n14315, n14116, n_7873);
  and g22218 (n14316, n_7872, n_7873);
  not g22219 (n_7999, n14315);
  not g22220 (n_8000, n14316);
  and g22221 (n14317, n_7999, n_8000);
  and g22222 (n14318, n14304, n14313);
  not g22223 (n_8001, n14314);
  not g22224 (n_8002, n14318);
  and g22225 (n14319, n_8001, n_8002);
  not g22226 (n_8003, n14317);
  and g22227 (n14320, n_8003, n14319);
  not g22228 (n_8004, n14320);
  and g22229 (n14321, n_8001, n_8004);
  not g22230 (n_8005, n14145);
  and g22231 (n14322, n_8005, n14148);
  not g22232 (n_8006, n14322);
  and g22233 (n14323, n_7891, n_8006);
  not g22234 (n_8007, n14321);
  and g22235 (n14324, n_8007, n14323);
  and g22236 (n14325, n_8003, n_8004);
  and g22237 (n14326, n14319, n_8004);
  not g22238 (n_8008, n14325);
  not g22239 (n_8009, n14326);
  and g22240 (n14327, n_8008, n_8009);
  and g22241 (n14328, n14291, n_7988);
  and g22242 (n14329, n_7987, n_7988);
  not g22243 (n_8010, n14328);
  not g22244 (n_8011, n14329);
  and g22245 (n14330, n_8010, n_8011);
  and g22246 (n14331, n14175, n14286);
  not g22247 (n_8012, n14331);
  and g22248 (n14332, n_7974, n_8012);
  and g22249 (n14333, n4694, n13630);
  and g22250 (n14334, n4533, n13515);
  and g22251 (n14335, n4604, n13597);
  and g22257 (n14338, n4536, n13976);
  not g22260 (n_8017, n14339);
  and g22261 (n14340, \a[23] , n_8017);
  not g22262 (n_8018, n14340);
  and g22263 (n14341, \a[23] , n_8018);
  and g22264 (n14342, n_8017, n_8018);
  not g22265 (n_8019, n14341);
  not g22266 (n_8020, n14342);
  and g22267 (n14343, n_8019, n_8020);
  not g22268 (n_8021, n14343);
  and g22269 (n14344, n14332, n_8021);
  not g22270 (n_8022, n14344);
  and g22271 (n14345, n14332, n_8022);
  and g22272 (n14346, n_8021, n_8022);
  not g22273 (n_8023, n14345);
  not g22274 (n_8024, n14346);
  and g22275 (n14347, n_8023, n_8024);
  and g22276 (n14348, n14273, n_7971);
  and g22277 (n14349, n_7970, n_7971);
  not g22278 (n_8025, n14348);
  not g22279 (n_8026, n14349);
  and g22280 (n14350, n_8025, n_8026);
  and g22281 (n14351, n14248, n_7940);
  and g22282 (n14352, n_7939, n_7940);
  not g22283 (n_8027, n14351);
  not g22284 (n_8028, n14352);
  and g22285 (n14353, n_8027, n_8028);
  and g22286 (n14354, n3457, n12370);
  and g22287 (n14355, n3542, n12508);
  and g22288 (n14356, n3606, n12505);
  and g22294 (n14359, n3368, n_7607);
  not g22297 (n_8033, n14360);
  and g22298 (n14361, \a[29] , n_8033);
  not g22299 (n_8034, n14361);
  and g22300 (n14362, \a[29] , n_8034);
  and g22301 (n14363, n_8033, n_8034);
  not g22302 (n_8035, n14362);
  not g22303 (n_8036, n14363);
  and g22304 (n14364, n_8035, n_8036);
  not g22305 (n_8037, n14353);
  not g22306 (n_8038, n14364);
  and g22307 (n14365, n_8037, n_8038);
  not g22308 (n_8039, n14365);
  and g22309 (n14366, n_8037, n_8039);
  and g22310 (n14367, n_8038, n_8039);
  not g22311 (n_8040, n14366);
  not g22312 (n_8041, n14367);
  and g22313 (n14368, n_8040, n_8041);
  and g22314 (n14369, n_7929, n_7931);
  and g22315 (n14370, n_7930, n14243);
  not g22316 (n_8042, n14369);
  not g22317 (n_8043, n14370);
  and g22318 (n14371, n_8042, n_8043);
  not g22370 (n_8044, n14403);
  not g22371 (n_8045, n14422);
  and g22372 (n14423, n_8044, n_8045);
  not g22373 (n_8046, n7632);
  not g22374 (n_8047, n7983);
  and g22375 (n14424, n_8046, n_8047);
  not g22376 (n_8048, n7291);
  and g22377 (n14425, n_8048, n14424);
  and g22378 (n14426, n_2446, n14425);
  not g22379 (n_8049, n14426);
  and g22380 (n14427, n_7417, n_8049);
  not g22381 (n_8050, n14427);
  and g22382 (n14428, \a[11] , n_8050);
  and g22383 (n14429, n_1071, n14427);
  not g22384 (n_8051, n14428);
  not g22385 (n_8052, n14429);
  and g22386 (n14430, n_8051, n_8052);
  and g22387 (n14431, n14403, n14422);
  not g22388 (n_8053, n14423);
  not g22389 (n_8054, n14431);
  and g22390 (n14432, n_8053, n_8054);
  and g22391 (n14433, n14430, n14432);
  not g22392 (n_8055, n14433);
  and g22393 (n14434, n_8053, n_8055);
  not g22394 (n_8056, n14434);
  and g22395 (n14435, n13821, n_8056);
  and g22396 (n14436, n_7617, n14434);
  not g22397 (n_8057, n14435);
  not g22398 (n_8058, n14436);
  and g22399 (n14437, n_8057, n_8058);
  and g22400 (n14438, n3020, n12516);
  and g22401 (n14439, n3028, n12519);
  and g22402 (n14440, n3023, n12522);
  and g22403 (n14441, n_7070, n_7073);
  and g22404 (n14442, n_7071, n12659);
  not g22405 (n_8059, n14441);
  not g22406 (n_8060, n14442);
  and g22407 (n14443, n_8059, n_8060);
  not g22408 (n_8061, n14443);
  and g22409 (n14444, n75, n_8061);
  not g22417 (n_8066, n14447);
  and g22418 (n14448, n14437, n_8066);
  not g22419 (n_8067, n14448);
  and g22420 (n14449, n_8057, n_8067);
  not g22421 (n_8068, n14371);
  not g22422 (n_8069, n14449);
  and g22423 (n14450, n_8068, n_8069);
  and g22424 (n14451, n14371, n14449);
  not g22425 (n_8070, n14450);
  not g22426 (n_8071, n14451);
  and g22427 (n14452, n_8070, n_8071);
  not g22428 (n_8072, n12653);
  and g22429 (n14453, n12651, n_8072);
  not g22430 (n_8073, n14453);
  and g22431 (n14454, n_7068, n_8073);
  and g22432 (n14455, n75, n14454);
  and g22433 (n14456, n3020, n12519);
  and g22434 (n14457, n3023, n12525);
  and g22435 (n14458, n3028, n12522);
  not g22443 (n_8078, n14430);
  not g22444 (n_8079, n14432);
  and g22445 (n14462, n_8078, n_8079);
  not g22446 (n_8080, n14462);
  and g22447 (n14463, n_8055, n_8080);
  not g22448 (n_8081, n14461);
  and g22449 (n14464, n_8081, n14463);
  not g22450 (n_8082, n14464);
  and g22451 (n14465, n14463, n_8082);
  and g22452 (n14466, n_8081, n_8082);
  not g22453 (n_8083, n14465);
  not g22454 (n_8084, n14466);
  and g22455 (n14467, n_8083, n_8084);
  not g22503 (n_8085, n14514);
  and g22504 (n14515, n14403, n_8085);
  and g22505 (n14516, n_8044, n14514);
  and g22506 (n14517, n_40, n454);
  and g22507 (n14518, n_62, n14517);
  and g22549 (n14560, n_239, n_261);
  and g22550 (n14561, n_138, n14560);
  not g22578 (n_8086, n14559);
  not g22579 (n_8087, n14588);
  and g22580 (n14589, n_8086, n_8087);
  not g22581 (n_8088, n8860);
  not g22582 (n_8089, n9331);
  and g22583 (n14590, n_8088, n_8089);
  not g22584 (n_8090, n8418);
  and g22585 (n14591, n_8090, n14590);
  and g22586 (n14592, n_3428, n14591);
  not g22587 (n_8091, n14592);
  and g22588 (n14593, n_7417, n_8091);
  not g22589 (n_8092, n14593);
  and g22590 (n14594, \a[8] , n_8092);
  and g22591 (n14595, n_1106, n14593);
  not g22592 (n_8093, n14594);
  not g22593 (n_8094, n14595);
  and g22594 (n14596, n_8093, n_8094);
  and g22595 (n14597, n14559, n14588);
  not g22596 (n_8095, n14589);
  not g22597 (n_8096, n14597);
  and g22598 (n14598, n_8095, n_8096);
  and g22599 (n14599, n14596, n14598);
  not g22600 (n_8097, n14599);
  and g22601 (n14600, n_8095, n_8097);
  not g22602 (n_8098, n14600);
  and g22603 (n14601, n14403, n_8098);
  and g22604 (n14602, n_8044, n14600);
  not g22605 (n_8099, n14601);
  not g22606 (n_8100, n14602);
  and g22607 (n14603, n_8099, n_8100);
  and g22608 (n14604, n3020, n12525);
  and g22609 (n14605, n3028, n12528);
  and g22610 (n14606, n3023, n12531);
  not g22611 (n_8101, n12645);
  and g22612 (n14607, n12643, n_8101);
  not g22613 (n_8102, n14607);
  and g22614 (n14608, n_7058, n_8102);
  and g22615 (n14609, n75, n14608);
  not g22623 (n_8107, n14612);
  and g22624 (n14613, n14603, n_8107);
  not g22625 (n_8108, n14613);
  and g22626 (n14614, n_8099, n_8108);
  not g22627 (n_8109, n14515);
  not g22628 (n_8110, n14614);
  and g22629 (n14615, n_8109, n_8110);
  not g22630 (n_8111, n14516);
  and g22631 (n14616, n_8111, n14615);
  not g22632 (n_8112, n14616);
  and g22633 (n14617, n_8109, n_8112);
  not g22634 (n_8113, n14467);
  not g22635 (n_8114, n14617);
  and g22636 (n14618, n_8113, n_8114);
  not g22637 (n_8115, n14618);
  and g22638 (n14619, n_8082, n_8115);
  not g22639 (n_8116, n14437);
  and g22640 (n14620, n_8116, n14447);
  not g22641 (n_8117, n14620);
  and g22642 (n14621, n_8067, n_8117);
  not g22643 (n_8118, n14619);
  and g22644 (n14622, n_8118, n14621);
  not g22645 (n_8119, n14621);
  and g22646 (n14623, n14619, n_8119);
  not g22647 (n_8120, n14622);
  not g22648 (n_8121, n14623);
  and g22649 (n14624, n_8120, n_8121);
  and g22650 (n14625, n3457, n12508);
  and g22651 (n14626, n3542, n12511);
  and g22652 (n14627, n3606, n12513);
  not g22653 (n_8122, n14626);
  not g22654 (n_8123, n14627);
  and g22655 (n14628, n_8122, n_8123);
  not g22656 (n_8124, n14625);
  and g22657 (n14629, n_8124, n14628);
  and g22658 (n14630, n_489, n14629);
  not g22659 (n_8125, n13863);
  and g22660 (n14631, n_8125, n14629);
  not g22661 (n_8126, n14630);
  not g22662 (n_8127, n14631);
  and g22663 (n14632, n_8126, n_8127);
  not g22664 (n_8128, n14632);
  and g22665 (n14633, \a[29] , n_8128);
  and g22666 (n14634, n_15, n14632);
  not g22667 (n_8129, n14633);
  not g22668 (n_8130, n14634);
  and g22669 (n14635, n_8129, n_8130);
  not g22670 (n_8131, n14635);
  and g22671 (n14636, n14624, n_8131);
  not g22672 (n_8132, n14636);
  and g22673 (n14637, n_8120, n_8132);
  not g22674 (n_8133, n14637);
  and g22675 (n14638, n14452, n_8133);
  not g22676 (n_8134, n14638);
  and g22677 (n14639, n_8070, n_8134);
  not g22678 (n_8135, n14368);
  not g22679 (n_8136, n14639);
  and g22680 (n14640, n_8135, n_8136);
  not g22681 (n_8137, n14640);
  and g22682 (n14641, n_8039, n_8137);
  not g22683 (n_8138, n14255);
  and g22684 (n14642, n_8138, n14266);
  not g22685 (n_8139, n14642);
  and g22686 (n14643, n_7956, n_8139);
  not g22687 (n_8140, n14641);
  and g22688 (n14644, n_8140, n14643);
  not g22689 (n_8141, n14643);
  and g22690 (n14645, n14641, n_8141);
  not g22691 (n_8142, n14644);
  not g22692 (n_8143, n14645);
  and g22693 (n14646, n_8142, n_8143);
  and g22694 (n14647, n3884, n13491);
  and g22695 (n14648, n3967, n12769);
  and g22696 (n14649, n4046, n12889);
  and g22702 (n14652, n4050, n_7447);
  not g22705 (n_8148, n14653);
  and g22706 (n14654, \a[26] , n_8148);
  not g22707 (n_8149, n14654);
  and g22708 (n14655, \a[26] , n_8149);
  and g22709 (n14656, n_8148, n_8149);
  not g22710 (n_8150, n14655);
  not g22711 (n_8151, n14656);
  and g22712 (n14657, n_8150, n_8151);
  not g22713 (n_8152, n14657);
  and g22714 (n14658, n14646, n_8152);
  not g22715 (n_8153, n14658);
  and g22716 (n14659, n_8142, n_8153);
  not g22717 (n_8154, n14350);
  not g22718 (n_8155, n14659);
  and g22719 (n14660, n_8154, n_8155);
  and g22720 (n14661, n14350, n14659);
  not g22721 (n_8156, n14660);
  not g22722 (n_8157, n14661);
  and g22723 (n14662, n_8156, n_8157);
  and g22724 (n14663, n4694, n13597);
  and g22725 (n14664, n4533, n13521);
  and g22726 (n14665, n4604, n13515);
  and g22732 (n14668, n4536, n_7765);
  not g22735 (n_8162, n14669);
  and g22736 (n14670, \a[23] , n_8162);
  not g22737 (n_8163, n14670);
  and g22738 (n14671, \a[23] , n_8163);
  and g22739 (n14672, n_8162, n_8163);
  not g22740 (n_8164, n14671);
  not g22741 (n_8165, n14672);
  and g22742 (n14673, n_8164, n_8165);
  not g22743 (n_8166, n14673);
  and g22744 (n14674, n14662, n_8166);
  not g22745 (n_8167, n14674);
  and g22746 (n14675, n_8156, n_8167);
  not g22747 (n_8168, n14347);
  not g22748 (n_8169, n14675);
  and g22749 (n14676, n_8168, n_8169);
  not g22750 (n_8170, n14676);
  and g22751 (n14677, n_8022, n_8170);
  not g22752 (n_8171, n14330);
  not g22753 (n_8172, n14677);
  and g22754 (n14678, n_8171, n_8172);
  and g22755 (n14679, n14330, n14677);
  not g22756 (n_8173, n14678);
  not g22757 (n_8174, n14679);
  and g22758 (n14680, n_8173, n_8174);
  and g22759 (n14681, n5496, n_7417);
  and g22760 (n14682, n4935, n_7540);
  and g22761 (n14683, n5407, n13941);
  and g22767 (n14686, n4938, n14028);
  not g22770 (n_8179, n14687);
  and g22771 (n14688, \a[20] , n_8179);
  not g22772 (n_8180, n14688);
  and g22773 (n14689, \a[20] , n_8180);
  and g22774 (n14690, n_8179, n_8180);
  not g22775 (n_8181, n14689);
  not g22776 (n_8182, n14690);
  and g22777 (n14691, n_8181, n_8182);
  not g22778 (n_8183, n14691);
  and g22779 (n14692, n14680, n_8183);
  not g22780 (n_8184, n14692);
  and g22781 (n14693, n_8173, n_8184);
  not g22782 (n_8185, n14327);
  not g22783 (n_8186, n14693);
  and g22784 (n14694, n_8185, n_8186);
  and g22785 (n14695, n14327, n14693);
  not g22786 (n_8187, n14694);
  not g22787 (n_8188, n14695);
  and g22788 (n14696, n_8187, n_8188);
  and g22789 (n14697, n14680, n_8184);
  and g22790 (n14698, n_8183, n_8184);
  not g22791 (n_8189, n14697);
  not g22792 (n_8190, n14698);
  and g22793 (n14699, n_8189, n_8190);
  and g22794 (n14700, n14662, n_8167);
  and g22795 (n14701, n_8166, n_8167);
  not g22796 (n_8191, n14700);
  not g22797 (n_8192, n14701);
  and g22798 (n14702, n_8191, n_8192);
  and g22799 (n14703, n14646, n_8153);
  and g22800 (n14704, n_8152, n_8153);
  not g22801 (n_8193, n14703);
  not g22802 (n_8194, n14704);
  and g22803 (n14705, n_8193, n_8194);
  and g22804 (n14706, n14368, n14639);
  not g22805 (n_8195, n14706);
  and g22806 (n14707, n_8137, n_8195);
  and g22807 (n14708, n3884, n12889);
  and g22808 (n14709, n3967, n12502);
  and g22809 (n14710, n4046, n12769);
  and g22815 (n14713, n4050, n12895);
  not g22818 (n_8200, n14714);
  and g22819 (n14715, \a[26] , n_8200);
  not g22820 (n_8201, n14715);
  and g22821 (n14716, \a[26] , n_8201);
  and g22822 (n14717, n_8200, n_8201);
  not g22823 (n_8202, n14716);
  not g22824 (n_8203, n14717);
  and g22825 (n14718, n_8202, n_8203);
  not g22826 (n_8204, n14718);
  and g22827 (n14719, n14707, n_8204);
  not g22828 (n_8205, n14719);
  and g22829 (n14720, n14707, n_8205);
  and g22830 (n14721, n_8204, n_8205);
  not g22831 (n_8206, n14720);
  not g22832 (n_8207, n14721);
  and g22833 (n14722, n_8206, n_8207);
  not g22834 (n_8208, n14452);
  and g22835 (n14723, n_8208, n14637);
  not g22836 (n_8209, n14723);
  and g22837 (n14724, n_8134, n_8209);
  and g22838 (n14725, n3457, n12505);
  and g22839 (n14726, n3542, n12513);
  and g22840 (n14727, n3606, n12508);
  and g22846 (n14730, n3368, n_7804);
  not g22849 (n_8214, n14731);
  and g22850 (n14732, \a[29] , n_8214);
  not g22851 (n_8215, n14732);
  and g22852 (n14733, \a[29] , n_8215);
  and g22853 (n14734, n_8214, n_8215);
  not g22854 (n_8216, n14733);
  not g22855 (n_8217, n14734);
  and g22856 (n14735, n_8216, n_8217);
  not g22857 (n_8218, n14735);
  and g22858 (n14736, n14724, n_8218);
  not g22859 (n_8219, n14736);
  and g22860 (n14737, n14724, n_8219);
  and g22861 (n14738, n_8218, n_8219);
  not g22862 (n_8220, n14737);
  not g22863 (n_8221, n14738);
  and g22864 (n14739, n_8220, n_8221);
  and g22865 (n14740, n3884, n12769);
  and g22866 (n14741, n3967, n12370);
  and g22867 (n14742, n4046, n12502);
  and g22873 (n14745, n4050, n12999);
  not g22876 (n_8226, n14746);
  and g22877 (n14747, \a[26] , n_8226);
  not g22878 (n_8227, n14747);
  and g22879 (n14748, \a[26] , n_8227);
  and g22880 (n14749, n_8226, n_8227);
  not g22881 (n_8228, n14748);
  not g22882 (n_8229, n14749);
  and g22883 (n14750, n_8228, n_8229);
  not g22884 (n_8230, n14739);
  not g22885 (n_8231, n14750);
  and g22886 (n14751, n_8230, n_8231);
  not g22887 (n_8232, n14751);
  and g22888 (n14752, n_8219, n_8232);
  not g22889 (n_8233, n14722);
  not g22890 (n_8234, n14752);
  and g22891 (n14753, n_8233, n_8234);
  not g22892 (n_8235, n14753);
  and g22893 (n14754, n_8205, n_8235);
  not g22894 (n_8236, n14705);
  not g22895 (n_8237, n14754);
  and g22896 (n14755, n_8236, n_8237);
  and g22897 (n14756, n14705, n14754);
  not g22898 (n_8238, n14755);
  not g22899 (n_8239, n14756);
  and g22900 (n14757, n_8238, n_8239);
  and g22901 (n14758, n4694, n13515);
  and g22902 (n14759, n4533, n13518);
  and g22903 (n14760, n4604, n13521);
  and g22909 (n14763, n4536, n13541);
  not g22912 (n_8244, n14764);
  and g22913 (n14765, \a[23] , n_8244);
  not g22914 (n_8245, n14765);
  and g22915 (n14766, \a[23] , n_8245);
  and g22916 (n14767, n_8244, n_8245);
  not g22917 (n_8246, n14766);
  not g22918 (n_8247, n14767);
  and g22919 (n14768, n_8246, n_8247);
  not g22920 (n_8248, n14768);
  and g22921 (n14769, n14757, n_8248);
  not g22922 (n_8249, n14769);
  and g22923 (n14770, n_8238, n_8249);
  not g22924 (n_8250, n14702);
  not g22925 (n_8251, n14770);
  and g22926 (n14771, n_8250, n_8251);
  and g22927 (n14772, n14702, n14770);
  not g22928 (n_8252, n14771);
  not g22929 (n_8253, n14772);
  and g22930 (n14773, n_8252, n_8253);
  and g22931 (n14774, n5496, n_7540);
  and g22932 (n14775, n4935, n13630);
  and g22933 (n14776, n5407, n13633);
  and g22939 (n14779, n4938, n_7563);
  not g22942 (n_8258, n14780);
  and g22943 (n14781, \a[20] , n_8258);
  not g22944 (n_8259, n14781);
  and g22945 (n14782, \a[20] , n_8259);
  and g22946 (n14783, n_8258, n_8259);
  not g22947 (n_8260, n14782);
  not g22948 (n_8261, n14783);
  and g22949 (n14784, n_8260, n_8261);
  not g22950 (n_8262, n14784);
  and g22951 (n14785, n14773, n_8262);
  not g22952 (n_8263, n14785);
  and g22953 (n14786, n_8252, n_8263);
  and g22954 (n14787, n5496, n13941);
  and g22955 (n14788, n4935, n13633);
  and g22956 (n14789, n5407, n_7540);
  and g22962 (n14792, n4938, n14136);
  not g22965 (n_8268, n14793);
  and g22966 (n14794, \a[20] , n_8268);
  not g22967 (n_8269, n14794);
  and g22968 (n14795, \a[20] , n_8269);
  and g22969 (n14796, n_8268, n_8269);
  not g22970 (n_8270, n14795);
  not g22971 (n_8271, n14796);
  and g22972 (n14797, n_8270, n_8271);
  not g22973 (n_8272, n14786);
  not g22974 (n_8273, n14797);
  and g22975 (n14798, n_8272, n_8273);
  and g22976 (n14799, n14347, n14675);
  not g22977 (n_8274, n14799);
  and g22978 (n14800, n_8170, n_8274);
  not g22979 (n_8275, n14798);
  and g22980 (n14801, n_8272, n_8275);
  and g22981 (n14802, n_8273, n_8275);
  not g22982 (n_8276, n14801);
  not g22983 (n_8277, n14802);
  and g22984 (n14803, n_8276, n_8277);
  not g22985 (n_8278, n14803);
  and g22986 (n14804, n14800, n_8278);
  not g22987 (n_8279, n14804);
  and g22988 (n14805, n_8275, n_8279);
  not g22989 (n_8280, n14699);
  not g22990 (n_8281, n14805);
  and g22991 (n14806, n_8280, n_8281);
  not g22992 (n_8282, n14806);
  and g22993 (n14807, n_8280, n_8282);
  and g22994 (n14808, n_8281, n_8282);
  not g22995 (n_8283, n14807);
  not g22996 (n_8284, n14808);
  and g22997 (n14809, n_8283, n_8284);
  and g22998 (n14810, n14757, n_8249);
  and g22999 (n14811, n_8248, n_8249);
  not g23000 (n_8285, n14810);
  not g23001 (n_8286, n14811);
  and g23002 (n14812, n_8285, n_8286);
  and g23003 (n14813, n14722, n14752);
  not g23004 (n_8287, n14813);
  and g23005 (n14814, n_8235, n_8287);
  and g23006 (n14815, n4694, n13521);
  and g23007 (n14816, n4533, n13491);
  and g23008 (n14817, n4604, n13518);
  and g23014 (n14820, n4536, n_7677);
  not g23017 (n_8292, n14821);
  and g23018 (n14822, \a[23] , n_8292);
  not g23019 (n_8293, n14822);
  and g23020 (n14823, \a[23] , n_8293);
  and g23021 (n14824, n_8292, n_8293);
  not g23022 (n_8294, n14823);
  not g23023 (n_8295, n14824);
  and g23024 (n14825, n_8294, n_8295);
  not g23025 (n_8296, n14825);
  and g23026 (n14826, n14814, n_8296);
  not g23027 (n_8297, n14826);
  and g23028 (n14827, n14814, n_8297);
  and g23029 (n14828, n_8296, n_8297);
  not g23030 (n_8298, n14827);
  not g23031 (n_8299, n14828);
  and g23032 (n14829, n_8298, n_8299);
  and g23033 (n14830, n_8230, n_8232);
  and g23034 (n14831, n_8231, n_8232);
  not g23035 (n_8300, n14830);
  not g23036 (n_8301, n14831);
  and g23037 (n14832, n_8300, n_8301);
  and g23038 (n14833, n_8110, n_8112);
  and g23039 (n14834, n_8111, n14617);
  not g23040 (n_8302, n14833);
  not g23041 (n_8303, n14834);
  and g23042 (n14835, n_8302, n_8303);
  not g23043 (n_8304, n12649);
  and g23044 (n14836, n12647, n_8304);
  not g23045 (n_8305, n14836);
  and g23046 (n14837, n_7063, n_8305);
  and g23047 (n14838, n75, n14837);
  and g23048 (n14839, n3020, n12522);
  and g23049 (n14840, n3023, n12528);
  and g23050 (n14841, n3028, n12525);
  not g23058 (n_8310, n14835);
  not g23059 (n_8311, n14844);
  and g23060 (n14845, n_8310, n_8311);
  not g23061 (n_8312, n14845);
  and g23062 (n14846, n_8310, n_8312);
  and g23063 (n14847, n_8311, n_8312);
  not g23064 (n_8313, n14846);
  not g23065 (n_8314, n14847);
  and g23066 (n14848, n_8313, n_8314);
  and g23067 (n14849, n3457, n12511);
  and g23068 (n14850, n3542, n12519);
  and g23069 (n14851, n3606, n12516);
  not g23070 (n_8315, n14850);
  not g23071 (n_8316, n14851);
  and g23072 (n14852, n_8315, n_8316);
  not g23073 (n_8317, n14849);
  and g23074 (n14853, n_8317, n14852);
  and g23075 (n14854, n_489, n14853);
  and g23076 (n14855, n14233, n14853);
  not g23077 (n_8318, n14854);
  not g23078 (n_8319, n14855);
  and g23079 (n14856, n_8318, n_8319);
  not g23080 (n_8320, n14856);
  and g23081 (n14857, \a[29] , n_8320);
  and g23082 (n14858, n_15, n14856);
  not g23083 (n_8321, n14857);
  not g23084 (n_8322, n14858);
  and g23085 (n14859, n_8321, n_8322);
  not g23086 (n_8323, n14848);
  not g23087 (n_8324, n14859);
  and g23088 (n14860, n_8323, n_8324);
  not g23089 (n_8325, n14860);
  and g23090 (n14861, n_8312, n_8325);
  and g23091 (n14862, n_8113, n_8115);
  and g23092 (n14863, n_8114, n_8115);
  not g23093 (n_8326, n14862);
  not g23094 (n_8327, n14863);
  and g23095 (n14864, n_8326, n_8327);
  not g23096 (n_8328, n14861);
  not g23097 (n_8329, n14864);
  and g23098 (n14865, n_8328, n_8329);
  not g23099 (n_8330, n14865);
  and g23100 (n14866, n_8328, n_8330);
  and g23101 (n14867, n_8329, n_8330);
  not g23102 (n_8331, n14866);
  not g23103 (n_8332, n14867);
  and g23104 (n14868, n_8331, n_8332);
  and g23105 (n14869, n3457, n12513);
  and g23106 (n14870, n3542, n12516);
  and g23107 (n14871, n3606, n12511);
  and g23113 (n14874, n3368, n14177);
  not g23116 (n_8337, n14875);
  and g23117 (n14876, \a[29] , n_8337);
  not g23118 (n_8338, n14876);
  and g23119 (n14877, \a[29] , n_8338);
  and g23120 (n14878, n_8337, n_8338);
  not g23121 (n_8339, n14877);
  not g23122 (n_8340, n14878);
  and g23123 (n14879, n_8339, n_8340);
  not g23124 (n_8341, n14868);
  not g23125 (n_8342, n14879);
  and g23126 (n14880, n_8341, n_8342);
  not g23127 (n_8343, n14880);
  and g23128 (n14881, n_8330, n_8343);
  not g23129 (n_8344, n14624);
  and g23130 (n14882, n_8344, n14635);
  not g23131 (n_8345, n14882);
  and g23132 (n14883, n_8132, n_8345);
  not g23133 (n_8346, n14881);
  and g23134 (n14884, n_8346, n14883);
  not g23135 (n_8347, n14883);
  and g23136 (n14885, n14881, n_8347);
  not g23137 (n_8348, n14884);
  not g23138 (n_8349, n14885);
  and g23139 (n14886, n_8348, n_8349);
  and g23140 (n14887, n3884, n12502);
  and g23141 (n14888, n3967, n12505);
  and g23142 (n14889, n4046, n12370);
  and g23148 (n14892, n4050, n_7594);
  not g23151 (n_8354, n14893);
  and g23152 (n14894, \a[26] , n_8354);
  not g23153 (n_8355, n14894);
  and g23154 (n14895, \a[26] , n_8355);
  and g23155 (n14896, n_8354, n_8355);
  not g23156 (n_8356, n14895);
  not g23157 (n_8357, n14896);
  and g23158 (n14897, n_8356, n_8357);
  not g23159 (n_8358, n14897);
  and g23160 (n14898, n14886, n_8358);
  not g23161 (n_8359, n14898);
  and g23162 (n14899, n_8348, n_8359);
  not g23163 (n_8360, n14832);
  not g23164 (n_8361, n14899);
  and g23165 (n14900, n_8360, n_8361);
  and g23166 (n14901, n14832, n14899);
  not g23167 (n_8362, n14900);
  not g23168 (n_8363, n14901);
  and g23169 (n14902, n_8362, n_8363);
  and g23170 (n14903, n4694, n13518);
  and g23171 (n14904, n4533, n12889);
  and g23172 (n14905, n4604, n13491);
  and g23178 (n14908, n4536, n13584);
  not g23181 (n_8368, n14909);
  and g23182 (n14910, \a[23] , n_8368);
  not g23183 (n_8369, n14910);
  and g23184 (n14911, \a[23] , n_8369);
  and g23185 (n14912, n_8368, n_8369);
  not g23186 (n_8370, n14911);
  not g23187 (n_8371, n14912);
  and g23188 (n14913, n_8370, n_8371);
  not g23189 (n_8372, n14913);
  and g23190 (n14914, n14902, n_8372);
  not g23191 (n_8373, n14914);
  and g23192 (n14915, n_8362, n_8373);
  not g23193 (n_8374, n14829);
  not g23194 (n_8375, n14915);
  and g23195 (n14916, n_8374, n_8375);
  not g23196 (n_8376, n14916);
  and g23197 (n14917, n_8297, n_8376);
  not g23198 (n_8377, n14812);
  not g23199 (n_8378, n14917);
  and g23200 (n14918, n_8377, n_8378);
  and g23201 (n14919, n14812, n14917);
  not g23202 (n_8379, n14918);
  not g23203 (n_8380, n14919);
  and g23204 (n14920, n_8379, n_8380);
  and g23205 (n14921, n5496, n13633);
  and g23206 (n14922, n4935, n13597);
  and g23207 (n14923, n5407, n13630);
  and g23213 (n14926, n4938, n13929);
  not g23216 (n_8385, n14927);
  and g23217 (n14928, \a[20] , n_8385);
  not g23218 (n_8386, n14928);
  and g23219 (n14929, \a[20] , n_8386);
  and g23220 (n14930, n_8385, n_8386);
  not g23221 (n_8387, n14929);
  not g23222 (n_8388, n14930);
  and g23223 (n14931, n_8387, n_8388);
  not g23224 (n_8389, n14931);
  and g23225 (n14932, n14920, n_8389);
  not g23226 (n_8390, n14932);
  and g23227 (n14933, n_8379, n_8390);
  not g23228 (n_8391, n13717);
  and g23229 (n14934, n_7417, n_8391);
  and g23230 (n14935, n5663, n13941);
  not g23231 (n_8392, n14934);
  not g23232 (n_8393, n14935);
  and g23233 (n14936, n_8392, n_8393);
  and g23234 (n14937, n_1409, n14936);
  and g23235 (n14938, n13951, n14936);
  not g23236 (n_8394, n14937);
  not g23237 (n_8395, n14938);
  and g23238 (n14939, n_8394, n_8395);
  not g23239 (n_8396, n14939);
  and g23240 (n14940, \a[17] , n_8396);
  and g23241 (n14941, n_617, n14939);
  not g23242 (n_8397, n14940);
  not g23243 (n_8398, n14941);
  and g23244 (n14942, n_8397, n_8398);
  not g23245 (n_8399, n14933);
  not g23246 (n_8400, n14942);
  and g23247 (n14943, n_8399, n_8400);
  and g23248 (n14944, n14773, n_8263);
  and g23249 (n14945, n_8262, n_8263);
  not g23250 (n_8401, n14944);
  not g23251 (n_8402, n14945);
  and g23252 (n14946, n_8401, n_8402);
  and g23253 (n14947, n14933, n14942);
  not g23254 (n_8403, n14943);
  not g23255 (n_8404, n14947);
  and g23256 (n14948, n_8403, n_8404);
  not g23257 (n_8405, n14946);
  and g23258 (n14949, n_8405, n14948);
  not g23259 (n_8406, n14949);
  and g23260 (n14950, n_8403, n_8406);
  not g23261 (n_8407, n14800);
  and g23262 (n14951, n_8407, n14803);
  not g23263 (n_8408, n14951);
  and g23264 (n14952, n_8279, n_8408);
  not g23265 (n_8409, n14950);
  and g23266 (n14953, n_8409, n14952);
  and g23267 (n14954, n_8405, n_8406);
  and g23268 (n14955, n14948, n_8406);
  not g23269 (n_8410, n14954);
  not g23270 (n_8411, n14955);
  and g23271 (n14956, n_8410, n_8411);
  and g23272 (n14957, n14920, n_8390);
  and g23273 (n14958, n_8389, n_8390);
  not g23274 (n_8412, n14957);
  not g23275 (n_8413, n14958);
  and g23276 (n14959, n_8412, n_8413);
  and g23277 (n14960, n14829, n14915);
  not g23278 (n_8414, n14960);
  and g23279 (n14961, n_8376, n_8414);
  and g23280 (n14962, n5496, n13630);
  and g23281 (n14963, n4935, n13515);
  and g23282 (n14964, n5407, n13597);
  and g23288 (n14967, n4938, n13976);
  not g23291 (n_8419, n14968);
  and g23292 (n14969, \a[20] , n_8419);
  not g23293 (n_8420, n14969);
  and g23294 (n14970, \a[20] , n_8420);
  and g23295 (n14971, n_8419, n_8420);
  not g23296 (n_8421, n14970);
  not g23297 (n_8422, n14971);
  and g23298 (n14972, n_8421, n_8422);
  not g23299 (n_8423, n14972);
  and g23300 (n14973, n14961, n_8423);
  not g23301 (n_8424, n14973);
  and g23302 (n14974, n14961, n_8424);
  and g23303 (n14975, n_8423, n_8424);
  not g23304 (n_8425, n14974);
  not g23305 (n_8426, n14975);
  and g23306 (n14976, n_8425, n_8426);
  and g23307 (n14977, n14902, n_8373);
  and g23308 (n14978, n_8372, n_8373);
  not g23309 (n_8427, n14977);
  not g23310 (n_8428, n14978);
  and g23311 (n14979, n_8427, n_8428);
  and g23312 (n14980, n14886, n_8359);
  and g23313 (n14981, n_8358, n_8359);
  not g23314 (n_8429, n14980);
  not g23315 (n_8430, n14981);
  and g23316 (n14982, n_8429, n_8430);
  and g23317 (n14983, n_8341, n_8343);
  and g23318 (n14984, n_8342, n_8343);
  not g23319 (n_8431, n14983);
  not g23320 (n_8432, n14984);
  and g23321 (n14985, n_8431, n_8432);
  and g23322 (n14986, n3884, n12370);
  and g23323 (n14987, n3967, n12508);
  and g23324 (n14988, n4046, n12505);
  and g23330 (n14991, n4050, n_7607);
  not g23333 (n_8437, n14992);
  and g23334 (n14993, \a[26] , n_8437);
  not g23335 (n_8438, n14993);
  and g23336 (n14994, \a[26] , n_8438);
  and g23337 (n14995, n_8437, n_8438);
  not g23338 (n_8439, n14994);
  not g23339 (n_8440, n14995);
  and g23340 (n14996, n_8439, n_8440);
  not g23341 (n_8441, n14985);
  not g23342 (n_8442, n14996);
  and g23343 (n14997, n_8441, n_8442);
  not g23344 (n_8443, n14997);
  and g23345 (n14998, n_8441, n_8443);
  and g23346 (n14999, n_8442, n_8443);
  not g23347 (n_8444, n14998);
  not g23348 (n_8445, n14999);
  and g23349 (n15000, n_8444, n_8445);
  and g23350 (n15001, n_7050, n_7053);
  and g23351 (n15002, n_7051, n12643);
  not g23352 (n_8446, n15001);
  not g23353 (n_8447, n15002);
  and g23354 (n15003, n_8446, n_8447);
  not g23355 (n_8448, n15003);
  and g23356 (n15004, n75, n_8448);
  and g23357 (n15005, n3020, n12528);
  and g23358 (n15006, n3023, n12534);
  and g23359 (n15007, n3028, n12531);
  and g23367 (n15011, n_254, n1139);
  and g23368 (n15012, n_277, n15011);
  not g23385 (n_8453, n15028);
  and g23386 (n15029, n14559, n_8453);
  and g23387 (n15030, n_8086, n15028);
  and g23388 (n15031, n11053, n11054);
  not g23389 (n_8454, n15031);
  and g23390 (n15032, n_7417, n_8454);
  not g23391 (n_8455, n15032);
  and g23392 (n15033, \a[2] , n_8455);
  and g23393 (n15034, n_10, n15032);
  not g23394 (n_8456, n15033);
  not g23395 (n_8457, n15034);
  and g23396 (n15035, n_8456, n_8457);
  not g23436 (n_8458, n15074);
  and g23437 (n15075, n15035, n_8458);
  not g23438 (n_8459, n71);
  not g23439 (n_8460, n10434);
  and g23440 (n15076, n_8459, n_8460);
  not g23441 (n_8461, n9867);
  and g23442 (n15077, n_8461, n15076);
  and g23443 (n15078, n_4684, n15077);
  not g23444 (n_8462, n15078);
  and g23445 (n15079, n_7417, n_8462);
  and g23446 (n15080, n_3, n15079);
  and g23447 (n15081, n15035, n15074);
  not g23448 (n_8463, n15035);
  and g23449 (n15082, n_8463, n_8458);
  not g23450 (n_8464, n15081);
  not g23451 (n_8465, n15082);
  and g23452 (n15083, n_8464, n_8465);
  not g23453 (n_8466, n15079);
  and g23454 (n15084, \a[5] , n_8466);
  not g23455 (n_8467, n15083);
  not g23456 (n_8468, n15084);
  and g23457 (n15085, n_8467, n_8468);
  not g23458 (n_8469, n15080);
  and g23459 (n15086, n_8469, n15085);
  not g23460 (n_8470, n15075);
  not g23461 (n_8471, n15086);
  and g23462 (n15087, n_8470, n_8471);
  not g23463 (n_8472, n15087);
  and g23464 (n15088, n14559, n_8472);
  and g23465 (n15089, n_8086, n15087);
  not g23466 (n_8473, n15088);
  not g23467 (n_8474, n15089);
  and g23468 (n15090, n_8473, n_8474);
  and g23469 (n15091, n3020, n12534);
  and g23470 (n15092, n3028, n12537);
  and g23471 (n15093, n3023, n12540);
  and g23472 (n15094, n_7040, n_7043);
  and g23473 (n15095, n_7041, n12635);
  not g23474 (n_8475, n15094);
  not g23475 (n_8476, n15095);
  and g23476 (n15096, n_8475, n_8476);
  not g23477 (n_8477, n15096);
  and g23478 (n15097, n75, n_8477);
  not g23486 (n_8482, n15100);
  and g23487 (n15101, n15090, n_8482);
  not g23488 (n_8483, n15101);
  and g23489 (n15102, n_8473, n_8483);
  not g23490 (n_8484, n15029);
  not g23491 (n_8485, n15102);
  and g23492 (n15103, n_8484, n_8485);
  not g23493 (n_8486, n15030);
  and g23494 (n15104, n_8486, n15103);
  not g23495 (n_8487, n15104);
  and g23496 (n15105, n_8484, n_8487);
  not g23497 (n_8488, n14596);
  not g23498 (n_8489, n14598);
  and g23499 (n15106, n_8488, n_8489);
  not g23500 (n_8490, n15106);
  and g23501 (n15107, n_8097, n_8490);
  not g23502 (n_8491, n15105);
  and g23503 (n15108, n_8491, n15107);
  not g23504 (n_8492, n15107);
  and g23505 (n15109, n15105, n_8492);
  not g23506 (n_8493, n15108);
  not g23507 (n_8494, n15109);
  and g23508 (n15110, n_8493, n_8494);
  not g23509 (n_8495, n15010);
  and g23510 (n15111, n_8495, n15110);
  not g23511 (n_8496, n15111);
  and g23512 (n15112, n_8493, n_8496);
  not g23513 (n_8497, n14603);
  and g23514 (n15113, n_8497, n14612);
  not g23515 (n_8498, n15113);
  and g23516 (n15114, n_8108, n_8498);
  not g23517 (n_8499, n15112);
  and g23518 (n15115, n_8499, n15114);
  not g23519 (n_8500, n15114);
  and g23520 (n15116, n15112, n_8500);
  not g23521 (n_8501, n15115);
  not g23522 (n_8502, n15116);
  and g23523 (n15117, n_8501, n_8502);
  and g23524 (n15118, n3457, n12516);
  and g23525 (n15119, n3542, n12522);
  and g23526 (n15120, n3606, n12519);
  not g23527 (n_8503, n15119);
  not g23528 (n_8504, n15120);
  and g23529 (n15121, n_8503, n_8504);
  not g23530 (n_8505, n15118);
  and g23531 (n15122, n_8505, n15121);
  and g23532 (n15123, n_489, n15122);
  and g23533 (n15124, n14443, n15122);
  not g23534 (n_8506, n15123);
  not g23535 (n_8507, n15124);
  and g23536 (n15125, n_8506, n_8507);
  not g23537 (n_8508, n15125);
  and g23538 (n15126, \a[29] , n_8508);
  and g23539 (n15127, n_15, n15125);
  not g23540 (n_8509, n15126);
  not g23541 (n_8510, n15127);
  and g23542 (n15128, n_8509, n_8510);
  not g23543 (n_8511, n15128);
  and g23544 (n15129, n15117, n_8511);
  not g23545 (n_8512, n15129);
  and g23546 (n15130, n_8501, n_8512);
  and g23547 (n15131, n14848, n14859);
  not g23548 (n_8513, n15131);
  and g23549 (n15132, n_8325, n_8513);
  not g23550 (n_8514, n15130);
  and g23551 (n15133, n_8514, n15132);
  not g23552 (n_8515, n15132);
  and g23553 (n15134, n15130, n_8515);
  not g23554 (n_8516, n15133);
  not g23555 (n_8517, n15134);
  and g23556 (n15135, n_8516, n_8517);
  and g23557 (n15136, n3884, n12505);
  and g23558 (n15137, n3967, n12513);
  and g23559 (n15138, n4046, n12508);
  and g23565 (n15141, n4050, n_7804);
  not g23568 (n_8522, n15142);
  and g23569 (n15143, \a[26] , n_8522);
  not g23570 (n_8523, n15143);
  and g23571 (n15144, \a[26] , n_8523);
  and g23572 (n15145, n_8522, n_8523);
  not g23573 (n_8524, n15144);
  not g23574 (n_8525, n15145);
  and g23575 (n15146, n_8524, n_8525);
  not g23576 (n_8526, n15146);
  and g23577 (n15147, n15135, n_8526);
  not g23578 (n_8527, n15147);
  and g23579 (n15148, n_8516, n_8527);
  not g23580 (n_8528, n15000);
  not g23581 (n_8529, n15148);
  and g23582 (n15149, n_8528, n_8529);
  not g23583 (n_8530, n15149);
  and g23584 (n15150, n_8443, n_8530);
  not g23585 (n_8531, n14982);
  not g23586 (n_8532, n15150);
  and g23587 (n15151, n_8531, n_8532);
  and g23588 (n15152, n14982, n15150);
  not g23589 (n_8533, n15151);
  not g23590 (n_8534, n15152);
  and g23591 (n15153, n_8533, n_8534);
  and g23592 (n15154, n4694, n13491);
  and g23593 (n15155, n4533, n12769);
  and g23594 (n15156, n4604, n12889);
  and g23600 (n15159, n4536, n_7447);
  not g23603 (n_8539, n15160);
  and g23604 (n15161, \a[23] , n_8539);
  not g23605 (n_8540, n15161);
  and g23606 (n15162, \a[23] , n_8540);
  and g23607 (n15163, n_8539, n_8540);
  not g23608 (n_8541, n15162);
  not g23609 (n_8542, n15163);
  and g23610 (n15164, n_8541, n_8542);
  not g23611 (n_8543, n15164);
  and g23612 (n15165, n15153, n_8543);
  not g23613 (n_8544, n15165);
  and g23614 (n15166, n_8533, n_8544);
  not g23615 (n_8545, n14979);
  not g23616 (n_8546, n15166);
  and g23617 (n15167, n_8545, n_8546);
  and g23618 (n15168, n14979, n15166);
  not g23619 (n_8547, n15167);
  not g23620 (n_8548, n15168);
  and g23621 (n15169, n_8547, n_8548);
  and g23622 (n15170, n5496, n13597);
  and g23623 (n15171, n4935, n13521);
  and g23624 (n15172, n5407, n13515);
  and g23630 (n15175, n4938, n_7765);
  not g23633 (n_8553, n15176);
  and g23634 (n15177, \a[20] , n_8553);
  not g23635 (n_8554, n15177);
  and g23636 (n15178, \a[20] , n_8554);
  and g23637 (n15179, n_8553, n_8554);
  not g23638 (n_8555, n15178);
  not g23639 (n_8556, n15179);
  and g23640 (n15180, n_8555, n_8556);
  not g23641 (n_8557, n15180);
  and g23642 (n15181, n15169, n_8557);
  not g23643 (n_8558, n15181);
  and g23644 (n15182, n_8547, n_8558);
  not g23645 (n_8559, n14976);
  not g23646 (n_8560, n15182);
  and g23647 (n15183, n_8559, n_8560);
  not g23648 (n_8561, n15183);
  and g23649 (n15184, n_8424, n_8561);
  not g23650 (n_8562, n14959);
  not g23651 (n_8563, n15184);
  and g23652 (n15185, n_8562, n_8563);
  and g23653 (n15186, n14959, n15184);
  not g23654 (n_8564, n15185);
  not g23655 (n_8565, n15186);
  and g23656 (n15187, n_8564, n_8565);
  and g23657 (n15188, n6233, n_7417);
  and g23658 (n15189, n5663, n_7540);
  and g23659 (n15190, n5939, n13941);
  and g23665 (n15193, n5666, n14028);
  not g23668 (n_8570, n15194);
  and g23669 (n15195, \a[17] , n_8570);
  not g23670 (n_8571, n15195);
  and g23671 (n15196, \a[17] , n_8571);
  and g23672 (n15197, n_8570, n_8571);
  not g23673 (n_8572, n15196);
  not g23674 (n_8573, n15197);
  and g23675 (n15198, n_8572, n_8573);
  not g23676 (n_8574, n15198);
  and g23677 (n15199, n15187, n_8574);
  not g23678 (n_8575, n15199);
  and g23679 (n15200, n_8564, n_8575);
  not g23680 (n_8576, n14956);
  not g23681 (n_8577, n15200);
  and g23682 (n15201, n_8576, n_8577);
  and g23683 (n15202, n14956, n15200);
  not g23684 (n_8578, n15201);
  not g23685 (n_8579, n15202);
  and g23686 (n15203, n_8578, n_8579);
  and g23687 (n15204, n15187, n_8575);
  and g23688 (n15205, n_8574, n_8575);
  not g23689 (n_8580, n15204);
  not g23690 (n_8581, n15205);
  and g23691 (n15206, n_8580, n_8581);
  and g23692 (n15207, n15169, n_8558);
  and g23693 (n15208, n_8557, n_8558);
  not g23694 (n_8582, n15207);
  not g23695 (n_8583, n15208);
  and g23696 (n15209, n_8582, n_8583);
  and g23697 (n15210, n15153, n_8544);
  and g23698 (n15211, n_8543, n_8544);
  not g23699 (n_8584, n15210);
  not g23700 (n_8585, n15211);
  and g23701 (n15212, n_8584, n_8585);
  and g23702 (n15213, n15000, n15148);
  not g23703 (n_8586, n15213);
  and g23704 (n15214, n_8530, n_8586);
  and g23705 (n15215, n4694, n12889);
  and g23706 (n15216, n4533, n12502);
  and g23707 (n15217, n4604, n12769);
  and g23713 (n15220, n4536, n12895);
  not g23716 (n_8591, n15221);
  and g23717 (n15222, \a[23] , n_8591);
  not g23718 (n_8592, n15222);
  and g23719 (n15223, \a[23] , n_8592);
  and g23720 (n15224, n_8591, n_8592);
  not g23721 (n_8593, n15223);
  not g23722 (n_8594, n15224);
  and g23723 (n15225, n_8593, n_8594);
  not g23724 (n_8595, n15225);
  and g23725 (n15226, n15214, n_8595);
  not g23726 (n_8596, n15226);
  and g23727 (n15227, n15214, n_8596);
  and g23728 (n15228, n_8595, n_8596);
  not g23729 (n_8597, n15227);
  not g23730 (n_8598, n15228);
  and g23731 (n15229, n_8597, n_8598);
  and g23732 (n15230, n15135, n_8527);
  and g23733 (n15231, n_8526, n_8527);
  not g23734 (n_8599, n15230);
  not g23735 (n_8600, n15231);
  and g23736 (n15232, n_8599, n_8600);
  and g23737 (n15233, n15110, n_8496);
  and g23738 (n15234, n_8495, n_8496);
  not g23739 (n_8601, n15233);
  not g23740 (n_8602, n15234);
  and g23741 (n15235, n_8601, n_8602);
  and g23742 (n15236, n3457, n12519);
  and g23743 (n15237, n3542, n12525);
  and g23744 (n15238, n3606, n12522);
  and g23750 (n15241, n3368, n14454);
  not g23753 (n_8607, n15242);
  and g23754 (n15243, \a[29] , n_8607);
  not g23755 (n_8608, n15243);
  and g23756 (n15244, \a[29] , n_8608);
  and g23757 (n15245, n_8607, n_8608);
  not g23758 (n_8609, n15244);
  not g23759 (n_8610, n15245);
  and g23760 (n15246, n_8609, n_8610);
  not g23761 (n_8611, n15235);
  not g23762 (n_8612, n15246);
  and g23763 (n15247, n_8611, n_8612);
  not g23764 (n_8613, n15247);
  and g23765 (n15248, n_8611, n_8613);
  and g23766 (n15249, n_8612, n_8613);
  not g23767 (n_8614, n15248);
  not g23768 (n_8615, n15249);
  and g23769 (n15250, n_8614, n_8615);
  and g23770 (n15251, n_8485, n_8487);
  and g23771 (n15252, n_8486, n15105);
  not g23772 (n_8616, n15251);
  not g23773 (n_8617, n15252);
  and g23774 (n15253, n_8616, n_8617);
  not g23775 (n_8618, n12637);
  and g23776 (n15254, n12635, n_8618);
  not g23777 (n_8619, n15254);
  and g23778 (n15255, n_7048, n_8619);
  and g23779 (n15256, n75, n15255);
  and g23780 (n15257, n3020, n12531);
  and g23781 (n15258, n3023, n12537);
  and g23782 (n15259, n3028, n12534);
  not g23790 (n_8624, n15253);
  not g23791 (n_8625, n15262);
  and g23792 (n15263, n_8624, n_8625);
  not g23793 (n_8626, n15263);
  and g23794 (n15264, n_8624, n_8626);
  and g23795 (n15265, n_8625, n_8626);
  not g23796 (n_8627, n15264);
  not g23797 (n_8628, n15265);
  and g23798 (n15266, n_8627, n_8628);
  not g23816 (n_8629, n15283);
  and g23817 (n15284, n_8463, n_8629);
  and g23818 (n15285, n634, n13774);
  and g23819 (n15286, n_148, n15285);
  not g23839 (n_8630, n15305);
  and g23840 (n15306, n_8463, n_8630);
  not g23887 (n_8631, n15352);
  and g23888 (n15353, n_8463, n_8631);
  and g23889 (n15354, n_7020, n_7023);
  and g23890 (n15355, n_7021, n12619);
  not g23891 (n_8632, n15354);
  not g23892 (n_8633, n15355);
  and g23893 (n15356, n_8632, n_8633);
  not g23894 (n_8634, n15356);
  and g23895 (n15357, n75, n_8634);
  and g23896 (n15358, n3020, n12546);
  and g23897 (n15359, n3023, n12552);
  and g23898 (n15360, n3028, n12549);
  and g23906 (n15364, n15035, n15352);
  not g23907 (n_8639, n15363);
  not g23908 (n_8640, n15364);
  and g23909 (n15365, n_8639, n_8640);
  not g23910 (n_8641, n15353);
  and g23911 (n15366, n_8641, n15365);
  not g23912 (n_8642, n15366);
  and g23913 (n15367, n_8641, n_8642);
  and g23914 (n15368, n15035, n15305);
  not g23915 (n_8643, n15367);
  not g23916 (n_8644, n15368);
  and g23917 (n15369, n_8643, n_8644);
  not g23918 (n_8645, n15306);
  and g23919 (n15370, n_8645, n15369);
  not g23920 (n_8646, n15370);
  and g23921 (n15371, n_8645, n_8646);
  and g23922 (n15372, n15035, n15283);
  not g23923 (n_8647, n15371);
  not g23924 (n_8648, n15372);
  and g23925 (n15373, n_8647, n_8648);
  not g23926 (n_8649, n15284);
  and g23927 (n15374, n_8649, n15373);
  not g23928 (n_8650, n15374);
  and g23929 (n15375, n_8649, n_8650);
  and g23930 (n15376, n_8467, n_8471);
  and g23931 (n15377, n_8468, n_8471);
  and g23932 (n15378, n_8469, n15377);
  not g23933 (n_8651, n15376);
  not g23934 (n_8652, n15378);
  and g23935 (n15379, n_8651, n_8652);
  not g23936 (n_8653, n15375);
  and g23937 (n15380, n_8653, n15379);
  not g23938 (n_8654, n15379);
  and g23939 (n15381, n15375, n_8654);
  not g23940 (n_8655, n15380);
  not g23941 (n_8656, n15381);
  and g23942 (n15382, n_8655, n_8656);
  and g23943 (n15383, n_7035, n_7038);
  and g23944 (n15384, n_7036, n12631);
  not g23945 (n_8657, n15383);
  not g23946 (n_8658, n15384);
  and g23947 (n15385, n_8657, n_8658);
  not g23948 (n_8659, n15385);
  and g23949 (n15386, n75, n_8659);
  and g23950 (n15387, n3020, n12537);
  and g23951 (n15388, n3023, n12543);
  and g23952 (n15389, n3028, n12540);
  not g23960 (n_8664, n15382);
  not g23961 (n_8665, n15392);
  and g23962 (n15393, n_8664, n_8665);
  and g23963 (n15394, n_8653, n_8654);
  not g23964 (n_8666, n15393);
  not g23965 (n_8667, n15394);
  and g23966 (n15395, n_8666, n_8667);
  not g23967 (n_8668, n15090);
  and g23968 (n15396, n_8668, n15100);
  not g23969 (n_8669, n15396);
  and g23970 (n15397, n_8483, n_8669);
  not g23971 (n_8670, n15395);
  and g23972 (n15398, n_8670, n15397);
  not g23973 (n_8671, n15397);
  and g23974 (n15399, n15395, n_8671);
  not g23975 (n_8672, n15398);
  not g23976 (n_8673, n15399);
  and g23977 (n15400, n_8672, n_8673);
  and g23978 (n15401, n3457, n12525);
  and g23979 (n15402, n3542, n12531);
  and g23980 (n15403, n3606, n12528);
  not g23981 (n_8674, n15402);
  not g23982 (n_8675, n15403);
  and g23983 (n15404, n_8674, n_8675);
  not g23984 (n_8676, n15401);
  and g23985 (n15405, n_8676, n15404);
  and g23986 (n15406, n_489, n15405);
  not g23987 (n_8677, n14608);
  and g23988 (n15407, n_8677, n15405);
  not g23989 (n_8678, n15406);
  not g23990 (n_8679, n15407);
  and g23991 (n15408, n_8678, n_8679);
  not g23992 (n_8680, n15408);
  and g23993 (n15409, \a[29] , n_8680);
  and g23994 (n15410, n_15, n15408);
  not g23995 (n_8681, n15409);
  not g23996 (n_8682, n15410);
  and g23997 (n15411, n_8681, n_8682);
  not g23998 (n_8683, n15411);
  and g23999 (n15412, n15400, n_8683);
  not g24000 (n_8684, n15412);
  and g24001 (n15413, n_8672, n_8684);
  not g24002 (n_8685, n15266);
  not g24003 (n_8686, n15413);
  and g24004 (n15414, n_8685, n_8686);
  not g24005 (n_8687, n15414);
  and g24006 (n15415, n_8626, n_8687);
  not g24007 (n_8688, n15250);
  not g24008 (n_8689, n15415);
  and g24009 (n15416, n_8688, n_8689);
  not g24010 (n_8690, n15416);
  and g24011 (n15417, n_8613, n_8690);
  not g24012 (n_8691, n15117);
  and g24013 (n15418, n_8691, n15128);
  not g24014 (n_8692, n15418);
  and g24015 (n15419, n_8512, n_8692);
  not g24016 (n_8693, n15417);
  and g24017 (n15420, n_8693, n15419);
  not g24018 (n_8694, n15419);
  and g24019 (n15421, n15417, n_8694);
  not g24020 (n_8695, n15420);
  not g24021 (n_8696, n15421);
  and g24022 (n15422, n_8695, n_8696);
  and g24023 (n15423, n3884, n12508);
  and g24024 (n15424, n3967, n12511);
  and g24025 (n15425, n4046, n12513);
  and g24031 (n15428, n4050, n13863);
  not g24034 (n_8701, n15429);
  and g24035 (n15430, \a[26] , n_8701);
  not g24036 (n_8702, n15430);
  and g24037 (n15431, \a[26] , n_8702);
  and g24038 (n15432, n_8701, n_8702);
  not g24039 (n_8703, n15431);
  not g24040 (n_8704, n15432);
  and g24041 (n15433, n_8703, n_8704);
  not g24042 (n_8705, n15433);
  and g24043 (n15434, n15422, n_8705);
  not g24044 (n_8706, n15434);
  and g24045 (n15435, n_8695, n_8706);
  not g24046 (n_8707, n15232);
  not g24047 (n_8708, n15435);
  and g24048 (n15436, n_8707, n_8708);
  and g24049 (n15437, n15232, n15435);
  not g24050 (n_8709, n15436);
  not g24051 (n_8710, n15437);
  and g24052 (n15438, n_8709, n_8710);
  and g24053 (n15439, n4694, n12769);
  and g24054 (n15440, n4533, n12370);
  and g24055 (n15441, n4604, n12502);
  and g24061 (n15444, n4536, n12999);
  not g24064 (n_8715, n15445);
  and g24065 (n15446, \a[23] , n_8715);
  not g24066 (n_8716, n15446);
  and g24067 (n15447, \a[23] , n_8716);
  and g24068 (n15448, n_8715, n_8716);
  not g24069 (n_8717, n15447);
  not g24070 (n_8718, n15448);
  and g24071 (n15449, n_8717, n_8718);
  not g24072 (n_8719, n15449);
  and g24073 (n15450, n15438, n_8719);
  not g24074 (n_8720, n15450);
  and g24075 (n15451, n_8709, n_8720);
  not g24076 (n_8721, n15229);
  not g24077 (n_8722, n15451);
  and g24078 (n15452, n_8721, n_8722);
  not g24079 (n_8723, n15452);
  and g24080 (n15453, n_8596, n_8723);
  not g24081 (n_8724, n15212);
  not g24082 (n_8725, n15453);
  and g24083 (n15454, n_8724, n_8725);
  and g24084 (n15455, n15212, n15453);
  not g24085 (n_8726, n15454);
  not g24086 (n_8727, n15455);
  and g24087 (n15456, n_8726, n_8727);
  and g24088 (n15457, n5496, n13515);
  and g24089 (n15458, n4935, n13518);
  and g24090 (n15459, n5407, n13521);
  and g24096 (n15462, n4938, n13541);
  not g24099 (n_8732, n15463);
  and g24100 (n15464, \a[20] , n_8732);
  not g24101 (n_8733, n15464);
  and g24102 (n15465, \a[20] , n_8733);
  and g24103 (n15466, n_8732, n_8733);
  not g24104 (n_8734, n15465);
  not g24105 (n_8735, n15466);
  and g24106 (n15467, n_8734, n_8735);
  not g24107 (n_8736, n15467);
  and g24108 (n15468, n15456, n_8736);
  not g24109 (n_8737, n15468);
  and g24110 (n15469, n_8726, n_8737);
  not g24111 (n_8738, n15209);
  not g24112 (n_8739, n15469);
  and g24113 (n15470, n_8738, n_8739);
  and g24114 (n15471, n15209, n15469);
  not g24115 (n_8740, n15470);
  not g24116 (n_8741, n15471);
  and g24117 (n15472, n_8740, n_8741);
  and g24118 (n15473, n6233, n_7540);
  and g24119 (n15474, n5663, n13630);
  and g24120 (n15475, n5939, n13633);
  and g24126 (n15478, n5666, n_7563);
  not g24129 (n_8746, n15479);
  and g24130 (n15480, \a[17] , n_8746);
  not g24131 (n_8747, n15480);
  and g24132 (n15481, \a[17] , n_8747);
  and g24133 (n15482, n_8746, n_8747);
  not g24134 (n_8748, n15481);
  not g24135 (n_8749, n15482);
  and g24136 (n15483, n_8748, n_8749);
  not g24137 (n_8750, n15483);
  and g24138 (n15484, n15472, n_8750);
  not g24139 (n_8751, n15484);
  and g24140 (n15485, n_8740, n_8751);
  and g24141 (n15486, n6233, n13941);
  and g24142 (n15487, n5663, n13633);
  and g24143 (n15488, n5939, n_7540);
  and g24149 (n15491, n5666, n14136);
  not g24152 (n_8756, n15492);
  and g24153 (n15493, \a[17] , n_8756);
  not g24154 (n_8757, n15493);
  and g24155 (n15494, \a[17] , n_8757);
  and g24156 (n15495, n_8756, n_8757);
  not g24157 (n_8758, n15494);
  not g24158 (n_8759, n15495);
  and g24159 (n15496, n_8758, n_8759);
  not g24160 (n_8760, n15485);
  not g24161 (n_8761, n15496);
  and g24162 (n15497, n_8760, n_8761);
  and g24163 (n15498, n14976, n15182);
  not g24164 (n_8762, n15498);
  and g24165 (n15499, n_8561, n_8762);
  not g24166 (n_8763, n15497);
  and g24167 (n15500, n_8760, n_8763);
  and g24168 (n15501, n_8761, n_8763);
  not g24169 (n_8764, n15500);
  not g24170 (n_8765, n15501);
  and g24171 (n15502, n_8764, n_8765);
  not g24172 (n_8766, n15502);
  and g24173 (n15503, n15499, n_8766);
  not g24174 (n_8767, n15503);
  and g24175 (n15504, n_8763, n_8767);
  not g24176 (n_8768, n15206);
  not g24177 (n_8769, n15504);
  and g24178 (n15505, n_8768, n_8769);
  not g24179 (n_8770, n15505);
  and g24180 (n15506, n_8768, n_8770);
  and g24181 (n15507, n_8769, n_8770);
  not g24182 (n_8771, n15506);
  not g24183 (n_8772, n15507);
  and g24184 (n15508, n_8771, n_8772);
  and g24185 (n15509, n15456, n_8737);
  and g24186 (n15510, n_8736, n_8737);
  not g24187 (n_8773, n15509);
  not g24188 (n_8774, n15510);
  and g24189 (n15511, n_8773, n_8774);
  and g24190 (n15512, n15229, n15451);
  not g24191 (n_8775, n15512);
  and g24192 (n15513, n_8723, n_8775);
  and g24193 (n15514, n5496, n13521);
  and g24194 (n15515, n4935, n13491);
  and g24195 (n15516, n5407, n13518);
  and g24201 (n15519, n4938, n_7677);
  not g24204 (n_8780, n15520);
  and g24205 (n15521, \a[20] , n_8780);
  not g24206 (n_8781, n15521);
  and g24207 (n15522, \a[20] , n_8781);
  and g24208 (n15523, n_8780, n_8781);
  not g24209 (n_8782, n15522);
  not g24210 (n_8783, n15523);
  and g24211 (n15524, n_8782, n_8783);
  not g24212 (n_8784, n15524);
  and g24213 (n15525, n15513, n_8784);
  not g24214 (n_8785, n15525);
  and g24215 (n15526, n15513, n_8785);
  and g24216 (n15527, n_8784, n_8785);
  not g24217 (n_8786, n15526);
  not g24218 (n_8787, n15527);
  and g24219 (n15528, n_8786, n_8787);
  and g24220 (n15529, n15438, n_8720);
  and g24221 (n15530, n_8719, n_8720);
  not g24222 (n_8788, n15529);
  not g24223 (n_8789, n15530);
  and g24224 (n15531, n_8788, n_8789);
  and g24225 (n15532, n15422, n_8706);
  and g24226 (n15533, n_8705, n_8706);
  not g24227 (n_8790, n15532);
  not g24228 (n_8791, n15533);
  and g24229 (n15534, n_8790, n_8791);
  and g24230 (n15535, n15250, n15415);
  not g24231 (n_8792, n15535);
  and g24232 (n15536, n_8690, n_8792);
  and g24233 (n15537, n3884, n12513);
  and g24234 (n15538, n3967, n12516);
  and g24235 (n15539, n4046, n12511);
  and g24241 (n15542, n4050, n14177);
  not g24244 (n_8797, n15543);
  and g24245 (n15544, \a[26] , n_8797);
  not g24246 (n_8798, n15544);
  and g24247 (n15545, \a[26] , n_8798);
  and g24248 (n15546, n_8797, n_8798);
  not g24249 (n_8799, n15545);
  not g24250 (n_8800, n15546);
  and g24251 (n15547, n_8799, n_8800);
  not g24252 (n_8801, n15547);
  and g24253 (n15548, n15536, n_8801);
  not g24254 (n_8802, n15548);
  and g24255 (n15549, n15536, n_8802);
  and g24256 (n15550, n_8801, n_8802);
  not g24257 (n_8803, n15549);
  not g24258 (n_8804, n15550);
  and g24259 (n15551, n_8803, n_8804);
  and g24260 (n15552, n15266, n15413);
  not g24261 (n_8805, n15552);
  and g24262 (n15553, n_8687, n_8805);
  and g24263 (n15554, n3457, n12522);
  and g24264 (n15555, n3542, n12528);
  and g24265 (n15556, n3606, n12525);
  and g24271 (n15559, n3368, n14837);
  not g24274 (n_8810, n15560);
  and g24275 (n15561, \a[29] , n_8810);
  not g24276 (n_8811, n15561);
  and g24277 (n15562, \a[29] , n_8811);
  and g24278 (n15563, n_8810, n_8811);
  not g24279 (n_8812, n15562);
  not g24280 (n_8813, n15563);
  and g24281 (n15564, n_8812, n_8813);
  not g24282 (n_8814, n15564);
  and g24283 (n15565, n15553, n_8814);
  not g24284 (n_8815, n15565);
  and g24285 (n15566, n15553, n_8815);
  and g24286 (n15567, n_8814, n_8815);
  not g24287 (n_8816, n15566);
  not g24288 (n_8817, n15567);
  and g24289 (n15568, n_8816, n_8817);
  and g24290 (n15569, n3884, n12511);
  and g24291 (n15570, n3967, n12519);
  and g24292 (n15571, n4046, n12516);
  and g24298 (n15574, n4050, n_7923);
  not g24301 (n_8822, n15575);
  and g24302 (n15576, \a[26] , n_8822);
  not g24303 (n_8823, n15576);
  and g24304 (n15577, \a[26] , n_8823);
  and g24305 (n15578, n_8822, n_8823);
  not g24306 (n_8824, n15577);
  not g24307 (n_8825, n15578);
  and g24308 (n15579, n_8824, n_8825);
  not g24309 (n_8826, n15568);
  not g24310 (n_8827, n15579);
  and g24311 (n15580, n_8826, n_8827);
  not g24312 (n_8828, n15580);
  and g24313 (n15581, n_8815, n_8828);
  not g24314 (n_8829, n15551);
  not g24315 (n_8830, n15581);
  and g24316 (n15582, n_8829, n_8830);
  not g24317 (n_8831, n15582);
  and g24318 (n15583, n_8802, n_8831);
  not g24319 (n_8832, n15534);
  not g24320 (n_8833, n15583);
  and g24321 (n15584, n_8832, n_8833);
  and g24322 (n15585, n15534, n15583);
  not g24323 (n_8834, n15584);
  not g24324 (n_8835, n15585);
  and g24325 (n15586, n_8834, n_8835);
  and g24326 (n15587, n4694, n12502);
  and g24327 (n15588, n4533, n12505);
  and g24328 (n15589, n4604, n12370);
  and g24334 (n15592, n4536, n_7594);
  not g24337 (n_8840, n15593);
  and g24338 (n15594, \a[23] , n_8840);
  not g24339 (n_8841, n15594);
  and g24340 (n15595, \a[23] , n_8841);
  and g24341 (n15596, n_8840, n_8841);
  not g24342 (n_8842, n15595);
  not g24343 (n_8843, n15596);
  and g24344 (n15597, n_8842, n_8843);
  not g24345 (n_8844, n15597);
  and g24346 (n15598, n15586, n_8844);
  not g24347 (n_8845, n15598);
  and g24348 (n15599, n_8834, n_8845);
  not g24349 (n_8846, n15531);
  not g24350 (n_8847, n15599);
  and g24351 (n15600, n_8846, n_8847);
  and g24352 (n15601, n15531, n15599);
  not g24353 (n_8848, n15600);
  not g24354 (n_8849, n15601);
  and g24355 (n15602, n_8848, n_8849);
  and g24356 (n15603, n5496, n13518);
  and g24357 (n15604, n4935, n12889);
  and g24358 (n15605, n5407, n13491);
  and g24364 (n15608, n4938, n13584);
  not g24367 (n_8854, n15609);
  and g24368 (n15610, \a[20] , n_8854);
  not g24369 (n_8855, n15610);
  and g24370 (n15611, \a[20] , n_8855);
  and g24371 (n15612, n_8854, n_8855);
  not g24372 (n_8856, n15611);
  not g24373 (n_8857, n15612);
  and g24374 (n15613, n_8856, n_8857);
  not g24375 (n_8858, n15613);
  and g24376 (n15614, n15602, n_8858);
  not g24377 (n_8859, n15614);
  and g24378 (n15615, n_8848, n_8859);
  not g24379 (n_8860, n15528);
  not g24380 (n_8861, n15615);
  and g24381 (n15616, n_8860, n_8861);
  not g24382 (n_8862, n15616);
  and g24383 (n15617, n_8785, n_8862);
  not g24384 (n_8863, n15511);
  not g24385 (n_8864, n15617);
  and g24386 (n15618, n_8863, n_8864);
  and g24387 (n15619, n15511, n15617);
  not g24388 (n_8865, n15618);
  not g24389 (n_8866, n15619);
  and g24390 (n15620, n_8865, n_8866);
  and g24391 (n15621, n6233, n13633);
  and g24392 (n15622, n5663, n13597);
  and g24393 (n15623, n5939, n13630);
  and g24399 (n15626, n5666, n13929);
  not g24402 (n_8871, n15627);
  and g24403 (n15628, \a[17] , n_8871);
  not g24404 (n_8872, n15628);
  and g24405 (n15629, \a[17] , n_8872);
  and g24406 (n15630, n_8871, n_8872);
  not g24407 (n_8873, n15629);
  not g24408 (n_8874, n15630);
  and g24409 (n15631, n_8873, n_8874);
  not g24410 (n_8875, n15631);
  and g24411 (n15632, n15620, n_8875);
  not g24412 (n_8876, n15632);
  and g24413 (n15633, n_8865, n_8876);
  not g24414 (n_8877, n13845);
  and g24415 (n15634, n_7417, n_8877);
  and g24416 (n15635, n6402, n13941);
  not g24417 (n_8878, n15634);
  not g24418 (n_8879, n15635);
  and g24419 (n15636, n_8878, n_8879);
  and g24420 (n15637, n_1885, n15636);
  and g24421 (n15638, n13951, n15636);
  not g24422 (n_8880, n15637);
  not g24423 (n_8881, n15638);
  and g24424 (n15639, n_8880, n_8881);
  not g24425 (n_8882, n15639);
  and g24426 (n15640, \a[14] , n_8882);
  and g24427 (n15641, n_652, n15639);
  not g24428 (n_8883, n15640);
  not g24429 (n_8884, n15641);
  and g24430 (n15642, n_8883, n_8884);
  not g24431 (n_8885, n15633);
  not g24432 (n_8886, n15642);
  and g24433 (n15643, n_8885, n_8886);
  and g24434 (n15644, n15472, n_8751);
  and g24435 (n15645, n_8750, n_8751);
  not g24436 (n_8887, n15644);
  not g24437 (n_8888, n15645);
  and g24438 (n15646, n_8887, n_8888);
  and g24439 (n15647, n15633, n15642);
  not g24440 (n_8889, n15643);
  not g24441 (n_8890, n15647);
  and g24442 (n15648, n_8889, n_8890);
  not g24443 (n_8891, n15646);
  and g24444 (n15649, n_8891, n15648);
  not g24445 (n_8892, n15649);
  and g24446 (n15650, n_8889, n_8892);
  not g24447 (n_8893, n15499);
  and g24448 (n15651, n_8893, n15502);
  not g24449 (n_8894, n15651);
  and g24450 (n15652, n_8767, n_8894);
  not g24451 (n_8895, n15650);
  and g24452 (n15653, n_8895, n15652);
  and g24453 (n15654, n_8891, n_8892);
  and g24454 (n15655, n15648, n_8892);
  not g24455 (n_8896, n15654);
  not g24456 (n_8897, n15655);
  and g24457 (n15656, n_8896, n_8897);
  and g24458 (n15657, n15620, n_8876);
  and g24459 (n15658, n_8875, n_8876);
  not g24460 (n_8898, n15657);
  not g24461 (n_8899, n15658);
  and g24462 (n15659, n_8898, n_8899);
  and g24463 (n15660, n15528, n15615);
  not g24464 (n_8900, n15660);
  and g24465 (n15661, n_8862, n_8900);
  and g24466 (n15662, n6233, n13630);
  and g24467 (n15663, n5663, n13515);
  and g24468 (n15664, n5939, n13597);
  and g24474 (n15667, n5666, n13976);
  not g24477 (n_8905, n15668);
  and g24478 (n15669, \a[17] , n_8905);
  not g24479 (n_8906, n15669);
  and g24480 (n15670, \a[17] , n_8906);
  and g24481 (n15671, n_8905, n_8906);
  not g24482 (n_8907, n15670);
  not g24483 (n_8908, n15671);
  and g24484 (n15672, n_8907, n_8908);
  not g24485 (n_8909, n15672);
  and g24486 (n15673, n15661, n_8909);
  not g24487 (n_8910, n15673);
  and g24488 (n15674, n15661, n_8910);
  and g24489 (n15675, n_8909, n_8910);
  not g24490 (n_8911, n15674);
  not g24491 (n_8912, n15675);
  and g24492 (n15676, n_8911, n_8912);
  and g24493 (n15677, n15602, n_8859);
  and g24494 (n15678, n_8858, n_8859);
  not g24495 (n_8913, n15677);
  not g24496 (n_8914, n15678);
  and g24497 (n15679, n_8913, n_8914);
  and g24498 (n15680, n15586, n_8845);
  and g24499 (n15681, n_8844, n_8845);
  not g24500 (n_8915, n15680);
  not g24501 (n_8916, n15681);
  and g24502 (n15682, n_8915, n_8916);
  and g24503 (n15683, n15551, n15581);
  not g24504 (n_8917, n15683);
  and g24505 (n15684, n_8831, n_8917);
  and g24506 (n15685, n4694, n12370);
  and g24507 (n15686, n4533, n12508);
  and g24508 (n15687, n4604, n12505);
  and g24514 (n15690, n4536, n_7607);
  not g24517 (n_8922, n15691);
  and g24518 (n15692, \a[23] , n_8922);
  not g24519 (n_8923, n15692);
  and g24520 (n15693, \a[23] , n_8923);
  and g24521 (n15694, n_8922, n_8923);
  not g24522 (n_8924, n15693);
  not g24523 (n_8925, n15694);
  and g24524 (n15695, n_8924, n_8925);
  not g24525 (n_8926, n15695);
  and g24526 (n15696, n15684, n_8926);
  not g24527 (n_8927, n15696);
  and g24528 (n15697, n15684, n_8927);
  and g24529 (n15698, n_8926, n_8927);
  not g24530 (n_8928, n15697);
  not g24531 (n_8929, n15698);
  and g24532 (n15699, n_8928, n_8929);
  and g24533 (n15700, n_8826, n_8828);
  and g24534 (n15701, n_8827, n_8828);
  not g24535 (n_8930, n15700);
  not g24536 (n_8931, n15701);
  and g24537 (n15702, n_8930, n_8931);
  and g24538 (n15703, n_8647, n_8650);
  and g24539 (n15704, n_8648, n15375);
  not g24540 (n_8932, n15703);
  not g24541 (n_8933, n15704);
  and g24542 (n15705, n_8932, n_8933);
  and g24543 (n15706, n_7030, n_7033);
  and g24544 (n15707, n_7031, n12627);
  not g24545 (n_8934, n15706);
  not g24546 (n_8935, n15707);
  and g24547 (n15708, n_8934, n_8935);
  not g24548 (n_8936, n15708);
  and g24549 (n15709, n75, n_8936);
  and g24550 (n15710, n3020, n12540);
  and g24551 (n15711, n3023, n12546);
  and g24552 (n15712, n3028, n12543);
  not g24560 (n_8941, n15705);
  not g24561 (n_8942, n15715);
  and g24562 (n15716, n_8941, n_8942);
  not g24563 (n_8943, n15716);
  and g24564 (n15717, n_8941, n_8943);
  and g24565 (n15718, n_8942, n_8943);
  not g24566 (n_8944, n15717);
  not g24567 (n_8945, n15718);
  and g24568 (n15719, n_8944, n_8945);
  and g24569 (n15720, n_8643, n_8646);
  and g24570 (n15721, n_8644, n15371);
  not g24571 (n_8946, n15720);
  not g24572 (n_8947, n15721);
  and g24573 (n15722, n_8946, n_8947);
  not g24574 (n_8948, n12621);
  and g24575 (n15723, n12619, n_8948);
  not g24576 (n_8949, n15723);
  and g24577 (n15724, n_7028, n_8949);
  and g24578 (n15725, n75, n15724);
  and g24579 (n15726, n3020, n12543);
  and g24580 (n15727, n3023, n12549);
  and g24581 (n15728, n3028, n12546);
  not g24589 (n_8954, n15722);
  not g24590 (n_8955, n15731);
  and g24591 (n15732, n_8954, n_8955);
  not g24592 (n_8956, n15732);
  and g24593 (n15733, n_8954, n_8956);
  and g24594 (n15734, n_8955, n_8956);
  not g24595 (n_8957, n15733);
  not g24596 (n_8958, n15734);
  and g24597 (n15735, n_8957, n_8958);
  and g24598 (n15736, n_8639, n_8642);
  and g24599 (n15737, n_8640, n15367);
  not g24600 (n_8959, n15736);
  not g24601 (n_8960, n15737);
  and g24602 (n15738, n_8959, n_8960);
  and g24624 (n15760, n3020, n12549);
  and g24625 (n15761, n3028, n12552);
  and g24626 (n15762, n3023, n12555);
  not g24627 (n_8961, n12613);
  and g24628 (n15763, n12611, n_8961);
  not g24629 (n_8962, n15763);
  and g24630 (n15764, n_7018, n_8962);
  and g24631 (n15765, n75, n15764);
  not g24639 (n_8967, n15759);
  not g24640 (n_8968, n15768);
  and g24641 (n15769, n_8967, n_8968);
  and g24658 (n15786, n3020, n12552);
  and g24659 (n15787, n3028, n12555);
  and g24660 (n15788, n3023, n12558);
  and g24661 (n15789, n_7010, n_7013);
  and g24662 (n15790, n_7011, n12611);
  not g24663 (n_8969, n15789);
  not g24664 (n_8970, n15790);
  and g24665 (n15791, n_8969, n_8970);
  not g24666 (n_8971, n15791);
  and g24667 (n15792, n75, n_8971);
  not g24675 (n_8976, n15785);
  not g24676 (n_8977, n15795);
  and g24677 (n15796, n_8976, n_8977);
  and g24692 (n15811, n3020, n12555);
  and g24693 (n15812, n3028, n12558);
  and g24694 (n15813, n3023, n12561);
  and g24695 (n15814, n_7005, n_7008);
  and g24696 (n15815, n_7006, n12607);
  not g24697 (n_8978, n15814);
  not g24698 (n_8979, n15815);
  and g24699 (n15816, n_8978, n_8979);
  not g24700 (n_8980, n15816);
  and g24701 (n15817, n75, n_8980);
  not g24709 (n_8985, n15810);
  not g24710 (n_8986, n15820);
  and g24711 (n15821, n_8985, n_8986);
  and g24733 (n15843, n3020, n12558);
  and g24734 (n15844, n3028, n12561);
  and g24735 (n15845, n3023, n12564);
  not g24736 (n_8987, n12601);
  and g24737 (n15846, n12599, n_8987);
  not g24738 (n_8988, n15846);
  and g24739 (n15847, n_7003, n_8988);
  and g24740 (n15848, n75, n15847);
  not g24748 (n_8993, n15842);
  not g24749 (n_8994, n15851);
  and g24750 (n15852, n_8993, n_8994);
  and g24751 (n15853, n_165, n_223);
  and g24752 (n15854, n_294, n15853);
  and g24779 (n15881, n_267, n12711);
  and g24780 (n15882, n_169, n15881);
  and g24798 (n15900, n3020, n12561);
  and g24799 (n15901, n3028, n12564);
  and g24800 (n15902, n3023, n12567);
  and g24801 (n15903, n_6995, n_6998);
  and g24802 (n15904, n_6996, n12599);
  not g24803 (n_8995, n15903);
  not g24804 (n_8996, n15904);
  and g24805 (n15905, n_8995, n_8996);
  not g24806 (n_8997, n15905);
  and g24807 (n15906, n75, n_8997);
  not g24815 (n_9002, n15899);
  not g24816 (n_9003, n15909);
  and g24817 (n15910, n_9002, n_9003);
  and g24846 (n15939, n3020, n12564);
  and g24847 (n15940, n3028, n12567);
  and g24848 (n15941, n3023, n12571);
  and g24849 (n15942, n_6991, n_6993);
  and g24850 (n15943, n_6992, n12595);
  not g24851 (n_9004, n15942);
  not g24852 (n_9005, n15943);
  and g24853 (n15944, n_9004, n_9005);
  not g24854 (n_9006, n15944);
  and g24855 (n15945, n75, n_9006);
  not g24863 (n_9011, n15938);
  not g24864 (n_9012, n15948);
  and g24865 (n15949, n_9011, n_9012);
  and g24901 (n15985, n3020, n12567);
  and g24902 (n15986, n3028, n12571);
  and g24903 (n15987, n3023, n12574);
  not g24904 (n_9013, n12590);
  and g24905 (n15988, n12588, n_9013);
  not g24906 (n_9014, n15988);
  and g24907 (n15989, n_6989, n_9014);
  and g24908 (n15990, n75, n15989);
  not g24916 (n_9019, n15984);
  not g24917 (n_9020, n15993);
  and g24918 (n15994, n_9019, n_9020);
  and g24933 (n16009, n3020, n12571);
  and g24934 (n16010, n3028, n12574);
  and g24935 (n16011, n3023, n12577);
  not g24936 (n_9021, n12586);
  and g24937 (n16012, n12584, n_9021);
  not g24938 (n_9022, n16012);
  and g24939 (n16013, n_6985, n_9022);
  and g24940 (n16014, n75, n16013);
  not g24948 (n_9027, n16008);
  not g24949 (n_9028, n16017);
  and g24950 (n16018, n_9027, n_9028);
  and g24951 (n16019, n_79, n_273);
  and g24952 (n16020, n_259, n16019);
  and g25014 (n16082, n3020, n12577);
  and g25015 (n16083, n12577, n12581);
  not g25016 (n_9029, n12577);
  and g25017 (n16084, n_9029, n_6977);
  not g25018 (n_9030, n16083);
  not g25019 (n_9031, n16084);
  and g25020 (n16085, n_9030, n_9031);
  not g25021 (n_9032, n16085);
  and g25022 (n16086, n75, n_9032);
  and g25023 (n16087, n3028, n_6977);
  not g25024 (n_9033, n16086);
  not g25025 (n_9034, n16087);
  and g25026 (n16088, n_9033, n_9034);
  not g25027 (n_9035, n16082);
  and g25028 (n16089, n_9035, n16088);
  not g25029 (n_9036, n16081);
  not g25030 (n_9037, n16089);
  and g25031 (n16090, n_9036, n_9037);
  not g25032 (n_9038, n16049);
  and g25033 (n16091, n_9038, n16090);
  and g25034 (n16092, n_6978, n16083);
  and g25035 (n16093, n12574, n_9030);
  not g25036 (n_9039, n16092);
  not g25037 (n_9040, n16093);
  and g25038 (n16094, n_9039, n_9040);
  not g25039 (n_9041, n16094);
  and g25040 (n16095, n75, n_9041);
  and g25041 (n16096, n3020, n12574);
  and g25042 (n16097, n3023, n_6977);
  and g25043 (n16098, n3028, n12577);
  not g25051 (n_9046, n16090);
  and g25052 (n16102, n16049, n_9046);
  not g25053 (n_9047, n16091);
  not g25054 (n_9048, n16102);
  and g25055 (n16103, n_9047, n_9048);
  not g25056 (n_9049, n16101);
  and g25057 (n16104, n_9049, n16103);
  not g25058 (n_9050, n16104);
  and g25059 (n16105, n_9047, n_9050);
  not g25060 (n_9051, n16018);
  and g25061 (n16106, n_9027, n_9051);
  and g25062 (n16107, n_9028, n_9051);
  not g25063 (n_9052, n16106);
  not g25064 (n_9053, n16107);
  and g25065 (n16108, n_9052, n_9053);
  not g25066 (n_9054, n16105);
  not g25067 (n_9055, n16108);
  and g25068 (n16109, n_9054, n_9055);
  not g25069 (n_9056, n16109);
  and g25070 (n16110, n_9051, n_9056);
  not g25071 (n_9057, n15994);
  and g25072 (n16111, n_9019, n_9057);
  and g25073 (n16112, n_9020, n_9057);
  not g25074 (n_9058, n16111);
  not g25075 (n_9059, n16112);
  and g25076 (n16113, n_9058, n_9059);
  not g25077 (n_9060, n16110);
  not g25078 (n_9061, n16113);
  and g25079 (n16114, n_9060, n_9061);
  not g25080 (n_9062, n16114);
  and g25081 (n16115, n_9057, n_9062);
  not g25082 (n_9063, n15949);
  and g25083 (n16116, n_9011, n_9063);
  and g25084 (n16117, n_9012, n_9063);
  not g25085 (n_9064, n16116);
  not g25086 (n_9065, n16117);
  and g25087 (n16118, n_9064, n_9065);
  not g25088 (n_9066, n16115);
  not g25089 (n_9067, n16118);
  and g25090 (n16119, n_9066, n_9067);
  not g25091 (n_9068, n16119);
  and g25092 (n16120, n_9063, n_9068);
  not g25093 (n_9069, n15910);
  and g25094 (n16121, n_9002, n_9069);
  and g25095 (n16122, n_9003, n_9069);
  not g25096 (n_9070, n16121);
  not g25097 (n_9071, n16122);
  and g25098 (n16123, n_9070, n_9071);
  not g25099 (n_9072, n16120);
  not g25100 (n_9073, n16123);
  and g25101 (n16124, n_9072, n_9073);
  not g25102 (n_9074, n16124);
  and g25103 (n16125, n_9069, n_9074);
  not g25104 (n_9075, n15852);
  and g25105 (n16126, n_8993, n_9075);
  and g25106 (n16127, n_8994, n_9075);
  not g25107 (n_9076, n16126);
  not g25108 (n_9077, n16127);
  and g25109 (n16128, n_9076, n_9077);
  not g25110 (n_9078, n16125);
  not g25111 (n_9079, n16128);
  and g25112 (n16129, n_9078, n_9079);
  not g25113 (n_9080, n16129);
  and g25114 (n16130, n_9075, n_9080);
  not g25115 (n_9081, n15821);
  and g25116 (n16131, n_8985, n_9081);
  and g25117 (n16132, n_8986, n_9081);
  not g25118 (n_9082, n16131);
  not g25119 (n_9083, n16132);
  and g25120 (n16133, n_9082, n_9083);
  not g25121 (n_9084, n16130);
  not g25122 (n_9085, n16133);
  and g25123 (n16134, n_9084, n_9085);
  not g25124 (n_9086, n16134);
  and g25125 (n16135, n_9081, n_9086);
  not g25126 (n_9087, n15796);
  and g25127 (n16136, n_8976, n_9087);
  and g25128 (n16137, n_8977, n_9087);
  not g25129 (n_9088, n16136);
  not g25130 (n_9089, n16137);
  and g25131 (n16138, n_9088, n_9089);
  not g25132 (n_9090, n16135);
  not g25133 (n_9091, n16138);
  and g25134 (n16139, n_9090, n_9091);
  not g25135 (n_9092, n16139);
  and g25136 (n16140, n_9087, n_9092);
  not g25137 (n_9093, n15769);
  and g25138 (n16141, n_8967, n_9093);
  and g25139 (n16142, n_8968, n_9093);
  not g25140 (n_9094, n16141);
  not g25141 (n_9095, n16142);
  and g25142 (n16143, n_9094, n_9095);
  not g25143 (n_9096, n16140);
  not g25144 (n_9097, n16143);
  and g25145 (n16144, n_9096, n_9097);
  not g25146 (n_9098, n16144);
  and g25147 (n16145, n_9093, n_9098);
  not g25148 (n_9099, n15738);
  not g25149 (n_9100, n16145);
  and g25150 (n16146, n_9099, n_9100);
  and g25151 (n16147, n15738, n16145);
  not g25152 (n_9101, n16146);
  not g25153 (n_9102, n16147);
  and g25154 (n16148, n_9101, n_9102);
  and g25155 (n16149, n3457, n12537);
  and g25156 (n16150, n3542, n12543);
  and g25157 (n16151, n3606, n12540);
  not g25158 (n_9103, n16150);
  not g25159 (n_9104, n16151);
  and g25160 (n16152, n_9103, n_9104);
  not g25161 (n_9105, n16149);
  and g25162 (n16153, n_9105, n16152);
  and g25163 (n16154, n_489, n16153);
  and g25164 (n16155, n15385, n16153);
  not g25165 (n_9106, n16154);
  not g25166 (n_9107, n16155);
  and g25167 (n16156, n_9106, n_9107);
  not g25168 (n_9108, n16156);
  and g25169 (n16157, \a[29] , n_9108);
  and g25170 (n16158, n_15, n16156);
  not g25171 (n_9109, n16157);
  not g25172 (n_9110, n16158);
  and g25173 (n16159, n_9109, n_9110);
  not g25174 (n_9111, n16159);
  and g25175 (n16160, n16148, n_9111);
  not g25176 (n_9112, n16160);
  and g25177 (n16161, n_9101, n_9112);
  not g25178 (n_9113, n15735);
  not g25179 (n_9114, n16161);
  and g25180 (n16162, n_9113, n_9114);
  not g25181 (n_9115, n16162);
  and g25182 (n16163, n_8956, n_9115);
  not g25183 (n_9116, n15719);
  not g25184 (n_9117, n16163);
  and g25185 (n16164, n_9116, n_9117);
  not g25186 (n_9118, n16164);
  and g25187 (n16165, n_8943, n_9118);
  and g25188 (n16166, n15382, n15392);
  not g25189 (n_9119, n16166);
  and g25190 (n16167, n_8666, n_9119);
  not g25191 (n_9120, n16165);
  and g25192 (n16168, n_9120, n16167);
  not g25193 (n_9121, n16167);
  and g25194 (n16169, n16165, n_9121);
  not g25195 (n_9122, n16168);
  not g25196 (n_9123, n16169);
  and g25197 (n16170, n_9122, n_9123);
  and g25198 (n16171, n3457, n12528);
  and g25199 (n16172, n3542, n12534);
  and g25200 (n16173, n3606, n12531);
  and g25206 (n16176, n3368, n_8448);
  not g25209 (n_9128, n16177);
  and g25210 (n16178, \a[29] , n_9128);
  not g25211 (n_9129, n16178);
  and g25212 (n16179, \a[29] , n_9129);
  and g25213 (n16180, n_9128, n_9129);
  not g25214 (n_9130, n16179);
  not g25215 (n_9131, n16180);
  and g25216 (n16181, n_9130, n_9131);
  not g25217 (n_9132, n16181);
  and g25218 (n16182, n16170, n_9132);
  not g25219 (n_9133, n16182);
  and g25220 (n16183, n_9122, n_9133);
  not g25221 (n_9134, n15400);
  and g25222 (n16184, n_9134, n15411);
  not g25223 (n_9135, n16184);
  and g25224 (n16185, n_8684, n_9135);
  not g25225 (n_9136, n16183);
  and g25226 (n16186, n_9136, n16185);
  not g25227 (n_9137, n16185);
  and g25228 (n16187, n16183, n_9137);
  not g25229 (n_9138, n16186);
  not g25230 (n_9139, n16187);
  and g25231 (n16188, n_9138, n_9139);
  and g25232 (n16189, n3884, n12516);
  and g25233 (n16190, n3967, n12522);
  and g25234 (n16191, n4046, n12519);
  and g25240 (n16194, n4050, n_8061);
  not g25243 (n_9144, n16195);
  and g25244 (n16196, \a[26] , n_9144);
  not g25245 (n_9145, n16196);
  and g25246 (n16197, \a[26] , n_9145);
  and g25247 (n16198, n_9144, n_9145);
  not g25248 (n_9146, n16197);
  not g25249 (n_9147, n16198);
  and g25250 (n16199, n_9146, n_9147);
  not g25251 (n_9148, n16199);
  and g25252 (n16200, n16188, n_9148);
  not g25253 (n_9149, n16200);
  and g25254 (n16201, n_9138, n_9149);
  not g25255 (n_9150, n15702);
  not g25256 (n_9151, n16201);
  and g25257 (n16202, n_9150, n_9151);
  and g25258 (n16203, n15702, n16201);
  not g25259 (n_9152, n16202);
  not g25260 (n_9153, n16203);
  and g25261 (n16204, n_9152, n_9153);
  and g25262 (n16205, n4694, n12505);
  and g25263 (n16206, n4533, n12513);
  and g25264 (n16207, n4604, n12508);
  and g25270 (n16210, n4536, n_7804);
  not g25273 (n_9158, n16211);
  and g25274 (n16212, \a[23] , n_9158);
  not g25275 (n_9159, n16212);
  and g25276 (n16213, \a[23] , n_9159);
  and g25277 (n16214, n_9158, n_9159);
  not g25278 (n_9160, n16213);
  not g25279 (n_9161, n16214);
  and g25280 (n16215, n_9160, n_9161);
  not g25281 (n_9162, n16215);
  and g25282 (n16216, n16204, n_9162);
  not g25283 (n_9163, n16216);
  and g25284 (n16217, n_9152, n_9163);
  not g25285 (n_9164, n15699);
  not g25286 (n_9165, n16217);
  and g25287 (n16218, n_9164, n_9165);
  not g25288 (n_9166, n16218);
  and g25289 (n16219, n_8927, n_9166);
  not g25290 (n_9167, n15682);
  not g25291 (n_9168, n16219);
  and g25292 (n16220, n_9167, n_9168);
  and g25293 (n16221, n15682, n16219);
  not g25294 (n_9169, n16220);
  not g25295 (n_9170, n16221);
  and g25296 (n16222, n_9169, n_9170);
  and g25297 (n16223, n5496, n13491);
  and g25298 (n16224, n4935, n12769);
  and g25299 (n16225, n5407, n12889);
  and g25305 (n16228, n4938, n_7447);
  not g25308 (n_9175, n16229);
  and g25309 (n16230, \a[20] , n_9175);
  not g25310 (n_9176, n16230);
  and g25311 (n16231, \a[20] , n_9176);
  and g25312 (n16232, n_9175, n_9176);
  not g25313 (n_9177, n16231);
  not g25314 (n_9178, n16232);
  and g25315 (n16233, n_9177, n_9178);
  not g25316 (n_9179, n16233);
  and g25317 (n16234, n16222, n_9179);
  not g25318 (n_9180, n16234);
  and g25319 (n16235, n_9169, n_9180);
  not g25320 (n_9181, n15679);
  not g25321 (n_9182, n16235);
  and g25322 (n16236, n_9181, n_9182);
  and g25323 (n16237, n15679, n16235);
  not g25324 (n_9183, n16236);
  not g25325 (n_9184, n16237);
  and g25326 (n16238, n_9183, n_9184);
  and g25327 (n16239, n6233, n13597);
  and g25328 (n16240, n5663, n13521);
  and g25329 (n16241, n5939, n13515);
  and g25335 (n16244, n5666, n_7765);
  not g25338 (n_9189, n16245);
  and g25339 (n16246, \a[17] , n_9189);
  not g25340 (n_9190, n16246);
  and g25341 (n16247, \a[17] , n_9190);
  and g25342 (n16248, n_9189, n_9190);
  not g25343 (n_9191, n16247);
  not g25344 (n_9192, n16248);
  and g25345 (n16249, n_9191, n_9192);
  not g25346 (n_9193, n16249);
  and g25347 (n16250, n16238, n_9193);
  not g25348 (n_9194, n16250);
  and g25349 (n16251, n_9183, n_9194);
  not g25350 (n_9195, n15676);
  not g25351 (n_9196, n16251);
  and g25352 (n16252, n_9195, n_9196);
  not g25353 (n_9197, n16252);
  and g25354 (n16253, n_8910, n_9197);
  not g25355 (n_9198, n15659);
  not g25356 (n_9199, n16253);
  and g25357 (n16254, n_9198, n_9199);
  and g25358 (n16255, n15659, n16253);
  not g25359 (n_9200, n16254);
  not g25360 (n_9201, n16255);
  and g25361 (n16256, n_9200, n_9201);
  and g25362 (n16257, n7101, n_7417);
  and g25363 (n16258, n6402, n_7540);
  and g25364 (n16259, n6951, n13941);
  and g25370 (n16262, n6397, n14028);
  not g25373 (n_9206, n16263);
  and g25374 (n16264, \a[14] , n_9206);
  not g25375 (n_9207, n16264);
  and g25376 (n16265, \a[14] , n_9207);
  and g25377 (n16266, n_9206, n_9207);
  not g25378 (n_9208, n16265);
  not g25379 (n_9209, n16266);
  and g25380 (n16267, n_9208, n_9209);
  not g25381 (n_9210, n16267);
  and g25382 (n16268, n16256, n_9210);
  not g25383 (n_9211, n16268);
  and g25384 (n16269, n_9200, n_9211);
  not g25385 (n_9212, n15656);
  not g25386 (n_9213, n16269);
  and g25387 (n16270, n_9212, n_9213);
  and g25388 (n16271, n15656, n16269);
  not g25389 (n_9214, n16270);
  not g25390 (n_9215, n16271);
  and g25391 (n16272, n_9214, n_9215);
  and g25392 (n16273, n16256, n_9211);
  and g25393 (n16274, n_9210, n_9211);
  not g25394 (n_9216, n16273);
  not g25395 (n_9217, n16274);
  and g25396 (n16275, n_9216, n_9217);
  and g25397 (n16276, n16238, n_9194);
  and g25398 (n16277, n_9193, n_9194);
  not g25399 (n_9218, n16276);
  not g25400 (n_9219, n16277);
  and g25401 (n16278, n_9218, n_9219);
  and g25402 (n16279, n16222, n_9180);
  and g25403 (n16280, n_9179, n_9180);
  not g25404 (n_9220, n16279);
  not g25405 (n_9221, n16280);
  and g25406 (n16281, n_9220, n_9221);
  and g25407 (n16282, n15699, n16217);
  not g25408 (n_9222, n16282);
  and g25409 (n16283, n_9166, n_9222);
  and g25410 (n16284, n5496, n12889);
  and g25411 (n16285, n4935, n12502);
  and g25412 (n16286, n5407, n12769);
  and g25418 (n16289, n4938, n12895);
  not g25421 (n_9227, n16290);
  and g25422 (n16291, \a[20] , n_9227);
  not g25423 (n_9228, n16291);
  and g25424 (n16292, \a[20] , n_9228);
  and g25425 (n16293, n_9227, n_9228);
  not g25426 (n_9229, n16292);
  not g25427 (n_9230, n16293);
  and g25428 (n16294, n_9229, n_9230);
  not g25429 (n_9231, n16294);
  and g25430 (n16295, n16283, n_9231);
  not g25431 (n_9232, n16295);
  and g25432 (n16296, n16283, n_9232);
  and g25433 (n16297, n_9231, n_9232);
  not g25434 (n_9233, n16296);
  not g25435 (n_9234, n16297);
  and g25436 (n16298, n_9233, n_9234);
  and g25437 (n16299, n16204, n_9163);
  and g25438 (n16300, n_9162, n_9163);
  not g25439 (n_9235, n16299);
  not g25440 (n_9236, n16300);
  and g25441 (n16301, n_9235, n_9236);
  and g25442 (n16302, n16188, n_9149);
  and g25443 (n16303, n_9148, n_9149);
  not g25444 (n_9237, n16302);
  not g25445 (n_9238, n16303);
  and g25446 (n16304, n_9237, n_9238);
  and g25447 (n16305, n16170, n_9133);
  and g25448 (n16306, n_9132, n_9133);
  not g25449 (n_9239, n16305);
  not g25450 (n_9240, n16306);
  and g25451 (n16307, n_9239, n_9240);
  and g25452 (n16308, n3884, n12519);
  and g25453 (n16309, n3967, n12525);
  and g25454 (n16310, n4046, n12522);
  and g25460 (n16313, n4050, n14454);
  not g25463 (n_9245, n16314);
  and g25464 (n16315, \a[26] , n_9245);
  not g25465 (n_9246, n16315);
  and g25466 (n16316, \a[26] , n_9246);
  and g25467 (n16317, n_9245, n_9246);
  not g25468 (n_9247, n16316);
  not g25469 (n_9248, n16317);
  and g25470 (n16318, n_9247, n_9248);
  not g25471 (n_9249, n16307);
  not g25472 (n_9250, n16318);
  and g25473 (n16319, n_9249, n_9250);
  not g25474 (n_9251, n16319);
  and g25475 (n16320, n_9249, n_9251);
  and g25476 (n16321, n_9250, n_9251);
  not g25477 (n_9252, n16320);
  not g25478 (n_9253, n16321);
  and g25479 (n16322, n_9252, n_9253);
  and g25480 (n16323, n15719, n16163);
  not g25481 (n_9254, n16323);
  and g25482 (n16324, n_9118, n_9254);
  and g25483 (n16325, n3457, n12531);
  and g25484 (n16326, n3542, n12537);
  and g25485 (n16327, n3606, n12534);
  and g25491 (n16330, n3368, n15255);
  not g25494 (n_9259, n16331);
  and g25495 (n16332, \a[29] , n_9259);
  not g25496 (n_9260, n16332);
  and g25497 (n16333, \a[29] , n_9260);
  and g25498 (n16334, n_9259, n_9260);
  not g25499 (n_9261, n16333);
  not g25500 (n_9262, n16334);
  and g25501 (n16335, n_9261, n_9262);
  not g25502 (n_9263, n16335);
  and g25503 (n16336, n16324, n_9263);
  not g25504 (n_9264, n16336);
  and g25505 (n16337, n16324, n_9264);
  and g25506 (n16338, n_9263, n_9264);
  not g25507 (n_9265, n16337);
  not g25508 (n_9266, n16338);
  and g25509 (n16339, n_9265, n_9266);
  and g25510 (n16340, n3967, n12528);
  and g25511 (n16341, n4046, n12525);
  and g25512 (n16342, n3884, n12522);
  and g25518 (n16345, n4050, n14837);
  not g25521 (n_9271, n16346);
  and g25522 (n16347, \a[26] , n_9271);
  not g25523 (n_9272, n16347);
  and g25524 (n16348, \a[26] , n_9272);
  and g25525 (n16349, n_9271, n_9272);
  not g25526 (n_9273, n16348);
  not g25527 (n_9274, n16349);
  and g25528 (n16350, n_9273, n_9274);
  not g25529 (n_9275, n16339);
  not g25530 (n_9276, n16350);
  and g25531 (n16351, n_9275, n_9276);
  not g25532 (n_9277, n16351);
  and g25533 (n16352, n_9264, n_9277);
  not g25534 (n_9278, n16322);
  not g25535 (n_9279, n16352);
  and g25536 (n16353, n_9278, n_9279);
  not g25537 (n_9280, n16353);
  and g25538 (n16354, n_9251, n_9280);
  not g25539 (n_9281, n16304);
  not g25540 (n_9282, n16354);
  and g25541 (n16355, n_9281, n_9282);
  and g25542 (n16356, n16304, n16354);
  not g25543 (n_9283, n16355);
  not g25544 (n_9284, n16356);
  and g25545 (n16357, n_9283, n_9284);
  and g25546 (n16358, n4694, n12508);
  and g25547 (n16359, n4533, n12511);
  and g25548 (n16360, n4604, n12513);
  and g25554 (n16363, n4536, n13863);
  not g25557 (n_9289, n16364);
  and g25558 (n16365, \a[23] , n_9289);
  not g25559 (n_9290, n16365);
  and g25560 (n16366, \a[23] , n_9290);
  and g25561 (n16367, n_9289, n_9290);
  not g25562 (n_9291, n16366);
  not g25563 (n_9292, n16367);
  and g25564 (n16368, n_9291, n_9292);
  not g25565 (n_9293, n16368);
  and g25566 (n16369, n16357, n_9293);
  not g25567 (n_9294, n16369);
  and g25568 (n16370, n_9283, n_9294);
  not g25569 (n_9295, n16301);
  not g25570 (n_9296, n16370);
  and g25571 (n16371, n_9295, n_9296);
  and g25572 (n16372, n16301, n16370);
  not g25573 (n_9297, n16371);
  not g25574 (n_9298, n16372);
  and g25575 (n16373, n_9297, n_9298);
  and g25576 (n16374, n5496, n12769);
  and g25577 (n16375, n4935, n12370);
  and g25578 (n16376, n5407, n12502);
  and g25584 (n16379, n4938, n12999);
  not g25587 (n_9303, n16380);
  and g25588 (n16381, \a[20] , n_9303);
  not g25589 (n_9304, n16381);
  and g25590 (n16382, \a[20] , n_9304);
  and g25591 (n16383, n_9303, n_9304);
  not g25592 (n_9305, n16382);
  not g25593 (n_9306, n16383);
  and g25594 (n16384, n_9305, n_9306);
  not g25595 (n_9307, n16384);
  and g25596 (n16385, n16373, n_9307);
  not g25597 (n_9308, n16385);
  and g25598 (n16386, n_9297, n_9308);
  not g25599 (n_9309, n16298);
  not g25600 (n_9310, n16386);
  and g25601 (n16387, n_9309, n_9310);
  not g25602 (n_9311, n16387);
  and g25603 (n16388, n_9232, n_9311);
  not g25604 (n_9312, n16281);
  not g25605 (n_9313, n16388);
  and g25606 (n16389, n_9312, n_9313);
  and g25607 (n16390, n16281, n16388);
  not g25608 (n_9314, n16389);
  not g25609 (n_9315, n16390);
  and g25610 (n16391, n_9314, n_9315);
  and g25611 (n16392, n6233, n13515);
  and g25612 (n16393, n5663, n13518);
  and g25613 (n16394, n5939, n13521);
  and g25619 (n16397, n5666, n13541);
  not g25622 (n_9320, n16398);
  and g25623 (n16399, \a[17] , n_9320);
  not g25624 (n_9321, n16399);
  and g25625 (n16400, \a[17] , n_9321);
  and g25626 (n16401, n_9320, n_9321);
  not g25627 (n_9322, n16400);
  not g25628 (n_9323, n16401);
  and g25629 (n16402, n_9322, n_9323);
  not g25630 (n_9324, n16402);
  and g25631 (n16403, n16391, n_9324);
  not g25632 (n_9325, n16403);
  and g25633 (n16404, n_9314, n_9325);
  not g25634 (n_9326, n16278);
  not g25635 (n_9327, n16404);
  and g25636 (n16405, n_9326, n_9327);
  and g25637 (n16406, n16278, n16404);
  not g25638 (n_9328, n16405);
  not g25639 (n_9329, n16406);
  and g25640 (n16407, n_9328, n_9329);
  and g25641 (n16408, n7101, n_7540);
  and g25642 (n16409, n6402, n13630);
  and g25643 (n16410, n6951, n13633);
  and g25649 (n16413, n6397, n_7563);
  not g25652 (n_9334, n16414);
  and g25653 (n16415, \a[14] , n_9334);
  not g25654 (n_9335, n16415);
  and g25655 (n16416, \a[14] , n_9335);
  and g25656 (n16417, n_9334, n_9335);
  not g25657 (n_9336, n16416);
  not g25658 (n_9337, n16417);
  and g25659 (n16418, n_9336, n_9337);
  not g25660 (n_9338, n16418);
  and g25661 (n16419, n16407, n_9338);
  not g25662 (n_9339, n16419);
  and g25663 (n16420, n_9328, n_9339);
  and g25664 (n16421, n7101, n13941);
  and g25665 (n16422, n6402, n13633);
  and g25666 (n16423, n6951, n_7540);
  and g25672 (n16426, n6397, n14136);
  not g25675 (n_9344, n16427);
  and g25676 (n16428, \a[14] , n_9344);
  not g25677 (n_9345, n16428);
  and g25678 (n16429, \a[14] , n_9345);
  and g25679 (n16430, n_9344, n_9345);
  not g25680 (n_9346, n16429);
  not g25681 (n_9347, n16430);
  and g25682 (n16431, n_9346, n_9347);
  not g25683 (n_9348, n16420);
  not g25684 (n_9349, n16431);
  and g25685 (n16432, n_9348, n_9349);
  and g25686 (n16433, n15676, n16251);
  not g25687 (n_9350, n16433);
  and g25688 (n16434, n_9197, n_9350);
  not g25689 (n_9351, n16432);
  and g25690 (n16435, n_9348, n_9351);
  and g25691 (n16436, n_9349, n_9351);
  not g25692 (n_9352, n16435);
  not g25693 (n_9353, n16436);
  and g25694 (n16437, n_9352, n_9353);
  not g25695 (n_9354, n16437);
  and g25696 (n16438, n16434, n_9354);
  not g25697 (n_9355, n16438);
  and g25698 (n16439, n_9351, n_9355);
  not g25699 (n_9356, n16275);
  not g25700 (n_9357, n16439);
  and g25701 (n16440, n_9356, n_9357);
  not g25702 (n_9358, n16440);
  and g25703 (n16441, n_9356, n_9358);
  and g25704 (n16442, n_9357, n_9358);
  not g25705 (n_9359, n16441);
  not g25706 (n_9360, n16442);
  and g25707 (n16443, n_9359, n_9360);
  and g25708 (n16444, n16391, n_9325);
  and g25709 (n16445, n_9324, n_9325);
  not g25710 (n_9361, n16444);
  not g25711 (n_9362, n16445);
  and g25712 (n16446, n_9361, n_9362);
  and g25713 (n16447, n16298, n16386);
  not g25714 (n_9363, n16447);
  and g25715 (n16448, n_9311, n_9363);
  and g25716 (n16449, n6233, n13521);
  and g25717 (n16450, n5663, n13491);
  and g25718 (n16451, n5939, n13518);
  and g25724 (n16454, n5666, n_7677);
  not g25727 (n_9368, n16455);
  and g25728 (n16456, \a[17] , n_9368);
  not g25729 (n_9369, n16456);
  and g25730 (n16457, \a[17] , n_9369);
  and g25731 (n16458, n_9368, n_9369);
  not g25732 (n_9370, n16457);
  not g25733 (n_9371, n16458);
  and g25734 (n16459, n_9370, n_9371);
  not g25735 (n_9372, n16459);
  and g25736 (n16460, n16448, n_9372);
  not g25737 (n_9373, n16460);
  and g25738 (n16461, n16448, n_9373);
  and g25739 (n16462, n_9372, n_9373);
  not g25740 (n_9374, n16461);
  not g25741 (n_9375, n16462);
  and g25742 (n16463, n_9374, n_9375);
  and g25743 (n16464, n16373, n_9308);
  and g25744 (n16465, n_9307, n_9308);
  not g25745 (n_9376, n16464);
  not g25746 (n_9377, n16465);
  and g25747 (n16466, n_9376, n_9377);
  and g25748 (n16467, n16357, n_9294);
  and g25749 (n16468, n_9293, n_9294);
  not g25750 (n_9378, n16467);
  not g25751 (n_9379, n16468);
  and g25752 (n16469, n_9378, n_9379);
  and g25753 (n16470, n16322, n16352);
  not g25754 (n_9380, n16470);
  and g25755 (n16471, n_9280, n_9380);
  and g25756 (n16472, n4694, n12513);
  and g25757 (n16473, n4533, n12516);
  and g25758 (n16474, n4604, n12511);
  and g25764 (n16477, n4536, n14177);
  not g25767 (n_9385, n16478);
  and g25768 (n16479, \a[23] , n_9385);
  not g25769 (n_9386, n16479);
  and g25770 (n16480, \a[23] , n_9386);
  and g25771 (n16481, n_9385, n_9386);
  not g25772 (n_9387, n16480);
  not g25773 (n_9388, n16481);
  and g25774 (n16482, n_9387, n_9388);
  not g25775 (n_9389, n16482);
  and g25776 (n16483, n16471, n_9389);
  not g25777 (n_9390, n16483);
  and g25778 (n16484, n16471, n_9390);
  and g25779 (n16485, n_9389, n_9390);
  not g25780 (n_9391, n16484);
  not g25781 (n_9392, n16485);
  and g25782 (n16486, n_9391, n_9392);
  and g25783 (n16487, n_9275, n_9277);
  and g25784 (n16488, n_9276, n_9277);
  not g25785 (n_9393, n16487);
  not g25786 (n_9394, n16488);
  and g25787 (n16489, n_9393, n_9394);
  and g25788 (n16490, n15735, n16161);
  not g25789 (n_9395, n16490);
  and g25790 (n16491, n_9115, n_9395);
  and g25791 (n16492, n3457, n12534);
  and g25792 (n16493, n3542, n12540);
  and g25793 (n16494, n3606, n12537);
  and g25799 (n16497, n3368, n_8477);
  not g25802 (n_9400, n16498);
  and g25803 (n16499, \a[29] , n_9400);
  not g25804 (n_9401, n16499);
  and g25805 (n16500, \a[29] , n_9401);
  and g25806 (n16501, n_9400, n_9401);
  not g25807 (n_9402, n16500);
  not g25808 (n_9403, n16501);
  and g25809 (n16502, n_9402, n_9403);
  not g25810 (n_9404, n16502);
  and g25811 (n16503, n16491, n_9404);
  not g25812 (n_9405, n16503);
  and g25813 (n16504, n16491, n_9405);
  and g25814 (n16505, n_9404, n_9405);
  not g25815 (n_9406, n16504);
  not g25816 (n_9407, n16505);
  and g25817 (n16506, n_9406, n_9407);
  and g25818 (n16507, n4046, n12528);
  and g25819 (n16508, n3884, n12525);
  and g25820 (n16509, n3967, n12531);
  and g25826 (n16512, n4050, n14608);
  not g25829 (n_9412, n16513);
  and g25830 (n16514, \a[26] , n_9412);
  not g25831 (n_9413, n16514);
  and g25832 (n16515, \a[26] , n_9413);
  and g25833 (n16516, n_9412, n_9413);
  not g25834 (n_9414, n16515);
  not g25835 (n_9415, n16516);
  and g25836 (n16517, n_9414, n_9415);
  not g25837 (n_9416, n16506);
  not g25838 (n_9417, n16517);
  and g25839 (n16518, n_9416, n_9417);
  not g25840 (n_9418, n16518);
  and g25841 (n16519, n_9405, n_9418);
  not g25842 (n_9419, n16489);
  not g25843 (n_9420, n16519);
  and g25844 (n16520, n_9419, n_9420);
  and g25845 (n16521, n16489, n16519);
  not g25846 (n_9421, n16520);
  not g25847 (n_9422, n16521);
  and g25848 (n16522, n_9421, n_9422);
  and g25849 (n16523, n4694, n12511);
  and g25850 (n16524, n4533, n12519);
  and g25851 (n16525, n4604, n12516);
  and g25857 (n16528, n4536, n_7923);
  not g25860 (n_9427, n16529);
  and g25861 (n16530, \a[23] , n_9427);
  not g25862 (n_9428, n16530);
  and g25863 (n16531, \a[23] , n_9428);
  and g25864 (n16532, n_9427, n_9428);
  not g25865 (n_9429, n16531);
  not g25866 (n_9430, n16532);
  and g25867 (n16533, n_9429, n_9430);
  not g25868 (n_9431, n16533);
  and g25869 (n16534, n16522, n_9431);
  not g25870 (n_9432, n16534);
  and g25871 (n16535, n_9421, n_9432);
  not g25872 (n_9433, n16486);
  not g25873 (n_9434, n16535);
  and g25874 (n16536, n_9433, n_9434);
  not g25875 (n_9435, n16536);
  and g25876 (n16537, n_9390, n_9435);
  not g25877 (n_9436, n16469);
  not g25878 (n_9437, n16537);
  and g25879 (n16538, n_9436, n_9437);
  and g25880 (n16539, n16469, n16537);
  not g25881 (n_9438, n16538);
  not g25882 (n_9439, n16539);
  and g25883 (n16540, n_9438, n_9439);
  and g25884 (n16541, n5496, n12502);
  and g25885 (n16542, n4935, n12505);
  and g25886 (n16543, n5407, n12370);
  and g25892 (n16546, n4938, n_7594);
  not g25895 (n_9444, n16547);
  and g25896 (n16548, \a[20] , n_9444);
  not g25897 (n_9445, n16548);
  and g25898 (n16549, \a[20] , n_9445);
  and g25899 (n16550, n_9444, n_9445);
  not g25900 (n_9446, n16549);
  not g25901 (n_9447, n16550);
  and g25902 (n16551, n_9446, n_9447);
  not g25903 (n_9448, n16551);
  and g25904 (n16552, n16540, n_9448);
  not g25905 (n_9449, n16552);
  and g25906 (n16553, n_9438, n_9449);
  not g25907 (n_9450, n16466);
  not g25908 (n_9451, n16553);
  and g25909 (n16554, n_9450, n_9451);
  and g25910 (n16555, n16466, n16553);
  not g25911 (n_9452, n16554);
  not g25912 (n_9453, n16555);
  and g25913 (n16556, n_9452, n_9453);
  and g25914 (n16557, n6233, n13518);
  and g25915 (n16558, n5663, n12889);
  and g25916 (n16559, n5939, n13491);
  and g25922 (n16562, n5666, n13584);
  not g25925 (n_9458, n16563);
  and g25926 (n16564, \a[17] , n_9458);
  not g25927 (n_9459, n16564);
  and g25928 (n16565, \a[17] , n_9459);
  and g25929 (n16566, n_9458, n_9459);
  not g25930 (n_9460, n16565);
  not g25931 (n_9461, n16566);
  and g25932 (n16567, n_9460, n_9461);
  not g25933 (n_9462, n16567);
  and g25934 (n16568, n16556, n_9462);
  not g25935 (n_9463, n16568);
  and g25936 (n16569, n_9452, n_9463);
  not g25937 (n_9464, n16463);
  not g25938 (n_9465, n16569);
  and g25939 (n16570, n_9464, n_9465);
  not g25940 (n_9466, n16570);
  and g25941 (n16571, n_9373, n_9466);
  not g25942 (n_9467, n16446);
  not g25943 (n_9468, n16571);
  and g25944 (n16572, n_9467, n_9468);
  and g25945 (n16573, n16446, n16571);
  not g25946 (n_9469, n16572);
  not g25947 (n_9470, n16573);
  and g25948 (n16574, n_9469, n_9470);
  and g25949 (n16575, n7101, n13633);
  and g25950 (n16576, n6402, n13597);
  and g25951 (n16577, n6951, n13630);
  and g25957 (n16580, n6397, n13929);
  not g25960 (n_9475, n16581);
  and g25961 (n16582, \a[14] , n_9475);
  not g25962 (n_9476, n16582);
  and g25963 (n16583, \a[14] , n_9476);
  and g25964 (n16584, n_9475, n_9476);
  not g25965 (n_9477, n16583);
  not g25966 (n_9478, n16584);
  and g25967 (n16585, n_9477, n_9478);
  not g25968 (n_9479, n16585);
  and g25969 (n16586, n16574, n_9479);
  not g25970 (n_9480, n16586);
  and g25971 (n16587, n_9469, n_9480);
  not g25972 (n_9481, n14424);
  and g25973 (n16588, n_7417, n_9481);
  and g25974 (n16589, n7291, n13941);
  not g25975 (n_9482, n16588);
  not g25976 (n_9483, n16589);
  and g25977 (n16590, n_9482, n_9483);
  and g25978 (n16591, n_2446, n16590);
  and g25979 (n16592, n13951, n16590);
  not g25980 (n_9484, n16591);
  not g25981 (n_9485, n16592);
  and g25982 (n16593, n_9484, n_9485);
  not g25983 (n_9486, n16593);
  and g25984 (n16594, \a[11] , n_9486);
  and g25985 (n16595, n_1071, n16593);
  not g25986 (n_9487, n16594);
  not g25987 (n_9488, n16595);
  and g25988 (n16596, n_9487, n_9488);
  not g25989 (n_9489, n16587);
  not g25990 (n_9490, n16596);
  and g25991 (n16597, n_9489, n_9490);
  and g25992 (n16598, n16407, n_9339);
  and g25993 (n16599, n_9338, n_9339);
  not g25994 (n_9491, n16598);
  not g25995 (n_9492, n16599);
  and g25996 (n16600, n_9491, n_9492);
  and g25997 (n16601, n16587, n16596);
  not g25998 (n_9493, n16597);
  not g25999 (n_9494, n16601);
  and g26000 (n16602, n_9493, n_9494);
  not g26001 (n_9495, n16600);
  and g26002 (n16603, n_9495, n16602);
  not g26003 (n_9496, n16603);
  and g26004 (n16604, n_9493, n_9496);
  not g26005 (n_9497, n16434);
  and g26006 (n16605, n_9497, n16437);
  not g26007 (n_9498, n16605);
  and g26008 (n16606, n_9355, n_9498);
  not g26009 (n_9499, n16604);
  and g26010 (n16607, n_9499, n16606);
  and g26011 (n16608, n_9495, n_9496);
  and g26012 (n16609, n16602, n_9496);
  not g26013 (n_9500, n16608);
  not g26014 (n_9501, n16609);
  and g26015 (n16610, n_9500, n_9501);
  and g26016 (n16611, n16574, n_9480);
  and g26017 (n16612, n_9479, n_9480);
  not g26018 (n_9502, n16611);
  not g26019 (n_9503, n16612);
  and g26020 (n16613, n_9502, n_9503);
  and g26021 (n16614, n16463, n16569);
  not g26022 (n_9504, n16614);
  and g26023 (n16615, n_9466, n_9504);
  and g26024 (n16616, n7101, n13630);
  and g26025 (n16617, n6402, n13515);
  and g26026 (n16618, n6951, n13597);
  and g26032 (n16621, n6397, n13976);
  not g26035 (n_9509, n16622);
  and g26036 (n16623, \a[14] , n_9509);
  not g26037 (n_9510, n16623);
  and g26038 (n16624, \a[14] , n_9510);
  and g26039 (n16625, n_9509, n_9510);
  not g26040 (n_9511, n16624);
  not g26041 (n_9512, n16625);
  and g26042 (n16626, n_9511, n_9512);
  not g26043 (n_9513, n16626);
  and g26044 (n16627, n16615, n_9513);
  not g26045 (n_9514, n16627);
  and g26046 (n16628, n16615, n_9514);
  and g26047 (n16629, n_9513, n_9514);
  not g26048 (n_9515, n16628);
  not g26049 (n_9516, n16629);
  and g26050 (n16630, n_9515, n_9516);
  and g26051 (n16631, n16556, n_9463);
  and g26052 (n16632, n_9462, n_9463);
  not g26053 (n_9517, n16631);
  not g26054 (n_9518, n16632);
  and g26055 (n16633, n_9517, n_9518);
  and g26056 (n16634, n16540, n_9449);
  and g26057 (n16635, n_9448, n_9449);
  not g26058 (n_9519, n16634);
  not g26059 (n_9520, n16635);
  and g26060 (n16636, n_9519, n_9520);
  and g26061 (n16637, n16486, n16535);
  not g26062 (n_9521, n16637);
  and g26063 (n16638, n_9435, n_9521);
  and g26064 (n16639, n5496, n12370);
  and g26065 (n16640, n4935, n12508);
  and g26066 (n16641, n5407, n12505);
  and g26072 (n16644, n4938, n_7607);
  not g26075 (n_9526, n16645);
  and g26076 (n16646, \a[20] , n_9526);
  not g26077 (n_9527, n16646);
  and g26078 (n16647, \a[20] , n_9527);
  and g26079 (n16648, n_9526, n_9527);
  not g26080 (n_9528, n16647);
  not g26081 (n_9529, n16648);
  and g26082 (n16649, n_9528, n_9529);
  not g26083 (n_9530, n16649);
  and g26084 (n16650, n16638, n_9530);
  not g26085 (n_9531, n16650);
  and g26086 (n16651, n16638, n_9531);
  and g26087 (n16652, n_9530, n_9531);
  not g26088 (n_9532, n16651);
  not g26089 (n_9533, n16652);
  and g26090 (n16653, n_9532, n_9533);
  and g26091 (n16654, n16522, n_9432);
  and g26092 (n16655, n_9431, n_9432);
  not g26093 (n_9534, n16654);
  not g26094 (n_9535, n16655);
  and g26095 (n16656, n_9534, n_9535);
  and g26096 (n16657, n_9416, n_9418);
  and g26097 (n16658, n_9417, n_9418);
  not g26098 (n_9536, n16657);
  not g26099 (n_9537, n16658);
  and g26100 (n16659, n_9536, n_9537);
  and g26101 (n16660, n_9096, n_9098);
  and g26102 (n16661, n_9097, n_9098);
  not g26103 (n_9538, n16660);
  not g26104 (n_9539, n16661);
  and g26105 (n16662, n_9538, n_9539);
  and g26106 (n16663, n3457, n12540);
  and g26107 (n16664, n3542, n12546);
  and g26108 (n16665, n3606, n12543);
  not g26109 (n_9540, n16664);
  not g26110 (n_9541, n16665);
  and g26111 (n16666, n_9540, n_9541);
  not g26112 (n_9542, n16663);
  and g26113 (n16667, n_9542, n16666);
  and g26114 (n16668, n_489, n16667);
  and g26115 (n16669, n15708, n16667);
  not g26116 (n_9543, n16668);
  not g26117 (n_9544, n16669);
  and g26118 (n16670, n_9543, n_9544);
  not g26119 (n_9545, n16670);
  and g26120 (n16671, \a[29] , n_9545);
  and g26121 (n16672, n_15, n16670);
  not g26122 (n_9546, n16671);
  not g26123 (n_9547, n16672);
  and g26124 (n16673, n_9546, n_9547);
  not g26125 (n_9548, n16662);
  not g26126 (n_9549, n16673);
  and g26127 (n16674, n_9548, n_9549);
  and g26128 (n16675, n_9090, n_9092);
  and g26129 (n16676, n_9091, n_9092);
  not g26130 (n_9550, n16675);
  not g26131 (n_9551, n16676);
  and g26132 (n16677, n_9550, n_9551);
  and g26133 (n16678, n3457, n12543);
  and g26134 (n16679, n3542, n12549);
  and g26135 (n16680, n3606, n12546);
  not g26136 (n_9552, n16679);
  not g26137 (n_9553, n16680);
  and g26138 (n16681, n_9552, n_9553);
  not g26139 (n_9554, n16678);
  and g26140 (n16682, n_9554, n16681);
  and g26141 (n16683, n_489, n16682);
  not g26142 (n_9555, n15724);
  and g26143 (n16684, n_9555, n16682);
  not g26144 (n_9556, n16683);
  not g26145 (n_9557, n16684);
  and g26146 (n16685, n_9556, n_9557);
  not g26147 (n_9558, n16685);
  and g26148 (n16686, \a[29] , n_9558);
  and g26149 (n16687, n_15, n16685);
  not g26150 (n_9559, n16686);
  not g26151 (n_9560, n16687);
  and g26152 (n16688, n_9559, n_9560);
  not g26153 (n_9561, n16677);
  not g26154 (n_9562, n16688);
  and g26155 (n16689, n_9561, n_9562);
  and g26156 (n16690, n_9084, n_9086);
  and g26157 (n16691, n_9085, n_9086);
  not g26158 (n_9563, n16690);
  not g26159 (n_9564, n16691);
  and g26160 (n16692, n_9563, n_9564);
  and g26161 (n16693, n3457, n12546);
  and g26162 (n16694, n3542, n12552);
  and g26163 (n16695, n3606, n12549);
  not g26164 (n_9565, n16694);
  not g26165 (n_9566, n16695);
  and g26166 (n16696, n_9565, n_9566);
  not g26167 (n_9567, n16693);
  and g26168 (n16697, n_9567, n16696);
  and g26169 (n16698, n_489, n16697);
  and g26170 (n16699, n15356, n16697);
  not g26171 (n_9568, n16698);
  not g26172 (n_9569, n16699);
  and g26173 (n16700, n_9568, n_9569);
  not g26174 (n_9570, n16700);
  and g26175 (n16701, \a[29] , n_9570);
  and g26176 (n16702, n_15, n16700);
  not g26177 (n_9571, n16701);
  not g26178 (n_9572, n16702);
  and g26179 (n16703, n_9571, n_9572);
  not g26180 (n_9573, n16692);
  not g26181 (n_9574, n16703);
  and g26182 (n16704, n_9573, n_9574);
  and g26183 (n16705, n_9078, n_9080);
  and g26184 (n16706, n_9079, n_9080);
  not g26185 (n_9575, n16705);
  not g26186 (n_9576, n16706);
  and g26187 (n16707, n_9575, n_9576);
  and g26188 (n16708, n3457, n12549);
  and g26189 (n16709, n3542, n12555);
  and g26190 (n16710, n3606, n12552);
  not g26191 (n_9577, n16709);
  not g26192 (n_9578, n16710);
  and g26193 (n16711, n_9577, n_9578);
  not g26194 (n_9579, n16708);
  and g26195 (n16712, n_9579, n16711);
  and g26196 (n16713, n_489, n16712);
  not g26197 (n_9580, n15764);
  and g26198 (n16714, n_9580, n16712);
  not g26199 (n_9581, n16713);
  not g26200 (n_9582, n16714);
  and g26201 (n16715, n_9581, n_9582);
  not g26202 (n_9583, n16715);
  and g26203 (n16716, \a[29] , n_9583);
  and g26204 (n16717, n_15, n16715);
  not g26205 (n_9584, n16716);
  not g26206 (n_9585, n16717);
  and g26207 (n16718, n_9584, n_9585);
  not g26208 (n_9586, n16707);
  not g26209 (n_9587, n16718);
  and g26210 (n16719, n_9586, n_9587);
  and g26211 (n16720, n_9072, n_9074);
  and g26212 (n16721, n_9073, n_9074);
  not g26213 (n_9588, n16720);
  not g26214 (n_9589, n16721);
  and g26215 (n16722, n_9588, n_9589);
  and g26216 (n16723, n3457, n12552);
  and g26217 (n16724, n3542, n12558);
  and g26218 (n16725, n3606, n12555);
  not g26219 (n_9590, n16724);
  not g26220 (n_9591, n16725);
  and g26221 (n16726, n_9590, n_9591);
  not g26222 (n_9592, n16723);
  and g26223 (n16727, n_9592, n16726);
  and g26224 (n16728, n_489, n16727);
  and g26225 (n16729, n15791, n16727);
  not g26226 (n_9593, n16728);
  not g26227 (n_9594, n16729);
  and g26228 (n16730, n_9593, n_9594);
  not g26229 (n_9595, n16730);
  and g26230 (n16731, \a[29] , n_9595);
  and g26231 (n16732, n_15, n16730);
  not g26232 (n_9596, n16731);
  not g26233 (n_9597, n16732);
  and g26234 (n16733, n_9596, n_9597);
  not g26235 (n_9598, n16722);
  not g26236 (n_9599, n16733);
  and g26237 (n16734, n_9598, n_9599);
  and g26238 (n16735, n3457, n12555);
  and g26239 (n16736, n3542, n12561);
  and g26240 (n16737, n3606, n12558);
  and g26246 (n16740, n3368, n_8980);
  not g26249 (n_9604, n16741);
  and g26250 (n16742, \a[29] , n_9604);
  not g26251 (n_9605, n16742);
  and g26252 (n16743, n_9604, n_9605);
  and g26253 (n16744, \a[29] , n_9605);
  not g26254 (n_9606, n16743);
  not g26255 (n_9607, n16744);
  and g26256 (n16745, n_9606, n_9607);
  and g26257 (n16746, n_9066, n_9068);
  and g26258 (n16747, n_9067, n_9068);
  not g26259 (n_9608, n16746);
  not g26260 (n_9609, n16747);
  and g26261 (n16748, n_9608, n_9609);
  not g26262 (n_9610, n16745);
  not g26263 (n_9611, n16748);
  and g26264 (n16749, n_9610, n_9611);
  not g26265 (n_9612, n16749);
  and g26266 (n16750, n_9610, n_9612);
  and g26267 (n16751, n_9611, n_9612);
  not g26268 (n_9613, n16750);
  not g26269 (n_9614, n16751);
  and g26270 (n16752, n_9613, n_9614);
  and g26271 (n16753, n3457, n12558);
  and g26272 (n16754, n3542, n12564);
  and g26273 (n16755, n3606, n12561);
  and g26279 (n16758, n3368, n15847);
  not g26282 (n_9619, n16759);
  and g26283 (n16760, \a[29] , n_9619);
  not g26284 (n_9620, n16760);
  and g26285 (n16761, n_9619, n_9620);
  and g26286 (n16762, \a[29] , n_9620);
  not g26287 (n_9621, n16761);
  not g26288 (n_9622, n16762);
  and g26289 (n16763, n_9621, n_9622);
  and g26290 (n16764, n_9060, n_9062);
  and g26291 (n16765, n_9061, n_9062);
  not g26292 (n_9623, n16764);
  not g26293 (n_9624, n16765);
  and g26294 (n16766, n_9623, n_9624);
  not g26295 (n_9625, n16763);
  not g26296 (n_9626, n16766);
  and g26297 (n16767, n_9625, n_9626);
  not g26298 (n_9627, n16767);
  and g26299 (n16768, n_9625, n_9627);
  and g26300 (n16769, n_9626, n_9627);
  not g26301 (n_9628, n16768);
  not g26302 (n_9629, n16769);
  and g26303 (n16770, n_9628, n_9629);
  and g26304 (n16771, n3457, n12561);
  and g26305 (n16772, n3542, n12567);
  and g26306 (n16773, n3606, n12564);
  and g26312 (n16776, n3368, n_8997);
  not g26315 (n_9634, n16777);
  and g26316 (n16778, \a[29] , n_9634);
  not g26317 (n_9635, n16778);
  and g26318 (n16779, n_9634, n_9635);
  and g26319 (n16780, \a[29] , n_9635);
  not g26320 (n_9636, n16779);
  not g26321 (n_9637, n16780);
  and g26322 (n16781, n_9636, n_9637);
  and g26323 (n16782, n_9054, n_9056);
  and g26324 (n16783, n_9055, n_9056);
  not g26325 (n_9638, n16782);
  not g26326 (n_9639, n16783);
  and g26327 (n16784, n_9638, n_9639);
  not g26328 (n_9640, n16781);
  not g26329 (n_9641, n16784);
  and g26330 (n16785, n_9640, n_9641);
  not g26331 (n_9642, n16785);
  and g26332 (n16786, n_9640, n_9642);
  and g26333 (n16787, n_9641, n_9642);
  not g26334 (n_9643, n16786);
  not g26335 (n_9644, n16787);
  and g26336 (n16788, n_9643, n_9644);
  and g26337 (n16789, n3457, n12564);
  and g26338 (n16790, n3542, n12571);
  and g26339 (n16791, n3606, n12567);
  and g26345 (n16794, n3368, n_9006);
  not g26348 (n_9649, n16795);
  and g26349 (n16796, \a[29] , n_9649);
  not g26350 (n_9650, n16796);
  and g26351 (n16797, n_9649, n_9650);
  and g26352 (n16798, \a[29] , n_9650);
  not g26353 (n_9651, n16797);
  not g26354 (n_9652, n16798);
  and g26355 (n16799, n_9651, n_9652);
  and g26356 (n16800, n_9049, n_9050);
  and g26357 (n16801, n16103, n_9050);
  not g26358 (n_9653, n16800);
  not g26359 (n_9654, n16801);
  and g26360 (n16802, n_9653, n_9654);
  not g26361 (n_9655, n16799);
  not g26362 (n_9656, n16802);
  and g26363 (n16803, n_9655, n_9656);
  not g26364 (n_9657, n16803);
  and g26365 (n16804, n_9655, n_9657);
  and g26366 (n16805, n_9656, n_9657);
  not g26367 (n_9658, n16804);
  not g26368 (n_9659, n16805);
  and g26369 (n16806, n_9658, n_9659);
  and g26370 (n16807, n3457, n12567);
  and g26371 (n16808, n3542, n12574);
  and g26372 (n16809, n3606, n12571);
  and g26378 (n16812, n3368, n15989);
  not g26381 (n_9664, n16813);
  and g26382 (n16814, \a[29] , n_9664);
  not g26383 (n_9665, n16814);
  and g26384 (n16815, n_9664, n_9665);
  and g26385 (n16816, \a[29] , n_9665);
  not g26386 (n_9666, n16815);
  not g26387 (n_9667, n16816);
  and g26388 (n16817, n_9666, n_9667);
  and g26389 (n16818, n_9036, n_9046);
  and g26390 (n16819, n_9037, n_9046);
  not g26391 (n_9668, n16818);
  not g26392 (n_9669, n16819);
  and g26393 (n16820, n_9668, n_9669);
  not g26394 (n_9670, n16817);
  not g26395 (n_9671, n16820);
  and g26396 (n16821, n_9670, n_9671);
  not g26397 (n_9672, n16821);
  and g26398 (n16822, n_9670, n_9672);
  and g26399 (n16823, n_9671, n_9672);
  not g26400 (n_9673, n16822);
  not g26401 (n_9674, n16823);
  and g26402 (n16824, n_9673, n_9674);
  and g26403 (n16825, n_2599, n_6977);
  and g26404 (n16826, n3606, n_6977);
  and g26405 (n16827, n3457, n12577);
  not g26406 (n_9675, n16826);
  not g26407 (n_9676, n16827);
  and g26408 (n16828, n_9675, n_9676);
  and g26409 (n16829, n3368, n_9032);
  not g26410 (n_9677, n16829);
  and g26411 (n16830, n16828, n_9677);
  not g26412 (n_9678, n16830);
  and g26413 (n16831, \a[29] , n_9678);
  not g26414 (n_9679, n16831);
  and g26415 (n16832, \a[29] , n_9679);
  and g26416 (n16833, n_9678, n_9679);
  not g26417 (n_9680, n16832);
  not g26418 (n_9681, n16833);
  and g26419 (n16834, n_9680, n_9681);
  and g26420 (n16835, n_479, n_6977);
  not g26421 (n_9682, n16835);
  and g26422 (n16836, \a[29] , n_9682);
  not g26423 (n_9683, n16834);
  and g26424 (n16837, n_9683, n16836);
  and g26425 (n16838, n3457, n12574);
  and g26426 (n16839, n3542, n_6977);
  and g26427 (n16840, n3606, n12577);
  not g26428 (n_9684, n16839);
  not g26429 (n_9685, n16840);
  and g26430 (n16841, n_9684, n_9685);
  not g26431 (n_9686, n16838);
  and g26432 (n16842, n_9686, n16841);
  and g26433 (n16843, n_489, n16842);
  and g26434 (n16844, n16094, n16842);
  not g26435 (n_9687, n16843);
  not g26436 (n_9688, n16844);
  and g26437 (n16845, n_9687, n_9688);
  not g26438 (n_9689, n16845);
  and g26439 (n16846, \a[29] , n_9689);
  and g26440 (n16847, n_15, n16845);
  not g26441 (n_9690, n16846);
  not g26442 (n_9691, n16847);
  and g26443 (n16848, n_9690, n_9691);
  not g26444 (n_9692, n16848);
  and g26445 (n16849, n16837, n_9692);
  and g26446 (n16850, n16825, n16849);
  and g26447 (n16851, n3457, n12571);
  and g26448 (n16852, n3542, n12577);
  and g26449 (n16853, n3606, n12574);
  and g26455 (n16856, n3368, n16013);
  not g26458 (n_9697, n16857);
  and g26459 (n16858, \a[29] , n_9697);
  not g26460 (n_9698, n16858);
  and g26461 (n16859, n_9697, n_9698);
  and g26462 (n16860, \a[29] , n_9698);
  not g26463 (n_9699, n16859);
  not g26464 (n_9700, n16860);
  and g26465 (n16861, n_9699, n_9700);
  not g26466 (n_9701, n16825);
  and g26467 (n16862, n_9701, n16849);
  not g26468 (n_9702, n16849);
  and g26469 (n16863, n16825, n_9702);
  not g26470 (n_9703, n16862);
  not g26471 (n_9704, n16863);
  and g26472 (n16864, n_9703, n_9704);
  not g26473 (n_9705, n16861);
  not g26474 (n_9706, n16864);
  and g26475 (n16865, n_9705, n_9706);
  not g26476 (n_9707, n16850);
  not g26477 (n_9708, n16865);
  and g26478 (n16866, n_9707, n_9708);
  not g26479 (n_9709, n16824);
  not g26480 (n_9710, n16866);
  and g26481 (n16867, n_9709, n_9710);
  not g26482 (n_9711, n16867);
  and g26483 (n16868, n_9672, n_9711);
  not g26484 (n_9712, n16806);
  not g26485 (n_9713, n16868);
  and g26486 (n16869, n_9712, n_9713);
  not g26487 (n_9714, n16869);
  and g26488 (n16870, n_9657, n_9714);
  not g26489 (n_9715, n16788);
  not g26490 (n_9716, n16870);
  and g26491 (n16871, n_9715, n_9716);
  not g26492 (n_9717, n16871);
  and g26493 (n16872, n_9642, n_9717);
  not g26494 (n_9718, n16770);
  not g26495 (n_9719, n16872);
  and g26496 (n16873, n_9718, n_9719);
  not g26497 (n_9720, n16873);
  and g26498 (n16874, n_9627, n_9720);
  not g26499 (n_9721, n16752);
  not g26500 (n_9722, n16874);
  and g26501 (n16875, n_9721, n_9722);
  not g26502 (n_9723, n16875);
  and g26503 (n16876, n_9612, n_9723);
  and g26504 (n16877, n16722, n16733);
  not g26505 (n_9724, n16734);
  not g26506 (n_9725, n16877);
  and g26507 (n16878, n_9724, n_9725);
  not g26508 (n_9726, n16876);
  and g26509 (n16879, n_9726, n16878);
  not g26510 (n_9727, n16879);
  and g26511 (n16880, n_9724, n_9727);
  and g26512 (n16881, n16707, n16718);
  not g26513 (n_9728, n16719);
  not g26514 (n_9729, n16881);
  and g26515 (n16882, n_9728, n_9729);
  not g26516 (n_9730, n16880);
  and g26517 (n16883, n_9730, n16882);
  not g26518 (n_9731, n16883);
  and g26519 (n16884, n_9728, n_9731);
  and g26520 (n16885, n16692, n16703);
  not g26521 (n_9732, n16704);
  not g26522 (n_9733, n16885);
  and g26523 (n16886, n_9732, n_9733);
  not g26524 (n_9734, n16884);
  and g26525 (n16887, n_9734, n16886);
  not g26526 (n_9735, n16887);
  and g26527 (n16888, n_9732, n_9735);
  and g26528 (n16889, n16677, n16688);
  not g26529 (n_9736, n16689);
  not g26530 (n_9737, n16889);
  and g26531 (n16890, n_9736, n_9737);
  not g26532 (n_9738, n16888);
  and g26533 (n16891, n_9738, n16890);
  not g26534 (n_9739, n16891);
  and g26535 (n16892, n_9736, n_9739);
  and g26536 (n16893, n16662, n16673);
  not g26537 (n_9740, n16674);
  not g26538 (n_9741, n16893);
  and g26539 (n16894, n_9740, n_9741);
  not g26540 (n_9742, n16892);
  and g26541 (n16895, n_9742, n16894);
  not g26542 (n_9743, n16895);
  and g26543 (n16896, n_9740, n_9743);
  not g26544 (n_9744, n16148);
  and g26545 (n16897, n_9744, n16159);
  not g26546 (n_9745, n16897);
  and g26547 (n16898, n_9112, n_9745);
  not g26548 (n_9746, n16896);
  and g26549 (n16899, n_9746, n16898);
  not g26550 (n_9747, n16898);
  and g26551 (n16900, n16896, n_9747);
  not g26552 (n_9748, n16899);
  not g26553 (n_9749, n16900);
  and g26554 (n16901, n_9748, n_9749);
  and g26555 (n16902, n3884, n12528);
  and g26556 (n16903, n3967, n12534);
  and g26557 (n16904, n4046, n12531);
  and g26563 (n16907, n4050, n_8448);
  not g26566 (n_9754, n16908);
  and g26567 (n16909, \a[26] , n_9754);
  not g26568 (n_9755, n16909);
  and g26569 (n16910, \a[26] , n_9755);
  and g26570 (n16911, n_9754, n_9755);
  not g26571 (n_9756, n16910);
  not g26572 (n_9757, n16911);
  and g26573 (n16912, n_9756, n_9757);
  not g26574 (n_9758, n16912);
  and g26575 (n16913, n16901, n_9758);
  not g26576 (n_9759, n16913);
  and g26577 (n16914, n_9748, n_9759);
  not g26578 (n_9760, n16659);
  not g26579 (n_9761, n16914);
  and g26580 (n16915, n_9760, n_9761);
  and g26581 (n16916, n16659, n16914);
  not g26582 (n_9762, n16915);
  not g26583 (n_9763, n16916);
  and g26584 (n16917, n_9762, n_9763);
  and g26585 (n16918, n4694, n12516);
  and g26586 (n16919, n4533, n12522);
  and g26587 (n16920, n4604, n12519);
  and g26593 (n16923, n4536, n_8061);
  not g26596 (n_9768, n16924);
  and g26597 (n16925, \a[23] , n_9768);
  not g26598 (n_9769, n16925);
  and g26599 (n16926, \a[23] , n_9769);
  and g26600 (n16927, n_9768, n_9769);
  not g26601 (n_9770, n16926);
  not g26602 (n_9771, n16927);
  and g26603 (n16928, n_9770, n_9771);
  not g26604 (n_9772, n16928);
  and g26605 (n16929, n16917, n_9772);
  not g26606 (n_9773, n16929);
  and g26607 (n16930, n_9762, n_9773);
  not g26608 (n_9774, n16656);
  not g26609 (n_9775, n16930);
  and g26610 (n16931, n_9774, n_9775);
  and g26611 (n16932, n16656, n16930);
  not g26612 (n_9776, n16931);
  not g26613 (n_9777, n16932);
  and g26614 (n16933, n_9776, n_9777);
  and g26615 (n16934, n5496, n12505);
  and g26616 (n16935, n4935, n12513);
  and g26617 (n16936, n5407, n12508);
  and g26623 (n16939, n4938, n_7804);
  not g26626 (n_9782, n16940);
  and g26627 (n16941, \a[20] , n_9782);
  not g26628 (n_9783, n16941);
  and g26629 (n16942, \a[20] , n_9783);
  and g26630 (n16943, n_9782, n_9783);
  not g26631 (n_9784, n16942);
  not g26632 (n_9785, n16943);
  and g26633 (n16944, n_9784, n_9785);
  not g26634 (n_9786, n16944);
  and g26635 (n16945, n16933, n_9786);
  not g26636 (n_9787, n16945);
  and g26637 (n16946, n_9776, n_9787);
  not g26638 (n_9788, n16653);
  not g26639 (n_9789, n16946);
  and g26640 (n16947, n_9788, n_9789);
  not g26641 (n_9790, n16947);
  and g26642 (n16948, n_9531, n_9790);
  not g26643 (n_9791, n16636);
  not g26644 (n_9792, n16948);
  and g26645 (n16949, n_9791, n_9792);
  and g26646 (n16950, n16636, n16948);
  not g26647 (n_9793, n16949);
  not g26648 (n_9794, n16950);
  and g26649 (n16951, n_9793, n_9794);
  and g26650 (n16952, n6233, n13491);
  and g26651 (n16953, n5663, n12769);
  and g26652 (n16954, n5939, n12889);
  and g26658 (n16957, n5666, n_7447);
  not g26661 (n_9799, n16958);
  and g26662 (n16959, \a[17] , n_9799);
  not g26663 (n_9800, n16959);
  and g26664 (n16960, \a[17] , n_9800);
  and g26665 (n16961, n_9799, n_9800);
  not g26666 (n_9801, n16960);
  not g26667 (n_9802, n16961);
  and g26668 (n16962, n_9801, n_9802);
  not g26669 (n_9803, n16962);
  and g26670 (n16963, n16951, n_9803);
  not g26671 (n_9804, n16963);
  and g26672 (n16964, n_9793, n_9804);
  not g26673 (n_9805, n16633);
  not g26674 (n_9806, n16964);
  and g26675 (n16965, n_9805, n_9806);
  and g26676 (n16966, n16633, n16964);
  not g26677 (n_9807, n16965);
  not g26678 (n_9808, n16966);
  and g26679 (n16967, n_9807, n_9808);
  and g26680 (n16968, n7101, n13597);
  and g26681 (n16969, n6402, n13521);
  and g26682 (n16970, n6951, n13515);
  and g26688 (n16973, n6397, n_7765);
  not g26691 (n_9813, n16974);
  and g26692 (n16975, \a[14] , n_9813);
  not g26693 (n_9814, n16975);
  and g26694 (n16976, \a[14] , n_9814);
  and g26695 (n16977, n_9813, n_9814);
  not g26696 (n_9815, n16976);
  not g26697 (n_9816, n16977);
  and g26698 (n16978, n_9815, n_9816);
  not g26699 (n_9817, n16978);
  and g26700 (n16979, n16967, n_9817);
  not g26701 (n_9818, n16979);
  and g26702 (n16980, n_9807, n_9818);
  not g26703 (n_9819, n16630);
  not g26704 (n_9820, n16980);
  and g26705 (n16981, n_9819, n_9820);
  not g26706 (n_9821, n16981);
  and g26707 (n16982, n_9514, n_9821);
  not g26708 (n_9822, n16613);
  not g26709 (n_9823, n16982);
  and g26710 (n16983, n_9822, n_9823);
  and g26711 (n16984, n16613, n16982);
  not g26712 (n_9824, n16983);
  not g26713 (n_9825, n16984);
  and g26714 (n16985, n_9824, n_9825);
  and g26715 (n16986, n7983, n_7417);
  and g26716 (n16987, n7291, n_7540);
  and g26717 (n16988, n7632, n13941);
  and g26723 (n16991, n7294, n14028);
  not g26726 (n_9830, n16992);
  and g26727 (n16993, \a[11] , n_9830);
  not g26728 (n_9831, n16993);
  and g26729 (n16994, \a[11] , n_9831);
  and g26730 (n16995, n_9830, n_9831);
  not g26731 (n_9832, n16994);
  not g26732 (n_9833, n16995);
  and g26733 (n16996, n_9832, n_9833);
  not g26734 (n_9834, n16996);
  and g26735 (n16997, n16985, n_9834);
  not g26736 (n_9835, n16997);
  and g26737 (n16998, n_9824, n_9835);
  not g26738 (n_9836, n16610);
  not g26739 (n_9837, n16998);
  and g26740 (n16999, n_9836, n_9837);
  and g26741 (n17000, n16610, n16998);
  not g26742 (n_9838, n16999);
  not g26743 (n_9839, n17000);
  and g26744 (n17001, n_9838, n_9839);
  and g26745 (n17002, n16985, n_9835);
  and g26746 (n17003, n_9834, n_9835);
  not g26747 (n_9840, n17002);
  not g26748 (n_9841, n17003);
  and g26749 (n17004, n_9840, n_9841);
  and g26750 (n17005, n16967, n_9818);
  and g26751 (n17006, n_9817, n_9818);
  not g26752 (n_9842, n17005);
  not g26753 (n_9843, n17006);
  and g26754 (n17007, n_9842, n_9843);
  and g26755 (n17008, n16951, n_9804);
  and g26756 (n17009, n_9803, n_9804);
  not g26757 (n_9844, n17008);
  not g26758 (n_9845, n17009);
  and g26759 (n17010, n_9844, n_9845);
  and g26760 (n17011, n16653, n16946);
  not g26761 (n_9846, n17011);
  and g26762 (n17012, n_9790, n_9846);
  and g26763 (n17013, n6233, n12889);
  and g26764 (n17014, n5663, n12502);
  and g26765 (n17015, n5939, n12769);
  and g26771 (n17018, n5666, n12895);
  not g26774 (n_9851, n17019);
  and g26775 (n17020, \a[17] , n_9851);
  not g26776 (n_9852, n17020);
  and g26777 (n17021, \a[17] , n_9852);
  and g26778 (n17022, n_9851, n_9852);
  not g26779 (n_9853, n17021);
  not g26780 (n_9854, n17022);
  and g26781 (n17023, n_9853, n_9854);
  not g26782 (n_9855, n17023);
  and g26783 (n17024, n17012, n_9855);
  not g26784 (n_9856, n17024);
  and g26785 (n17025, n17012, n_9856);
  and g26786 (n17026, n_9855, n_9856);
  not g26787 (n_9857, n17025);
  not g26788 (n_9858, n17026);
  and g26789 (n17027, n_9857, n_9858);
  and g26790 (n17028, n16933, n_9787);
  and g26791 (n17029, n_9786, n_9787);
  not g26792 (n_9859, n17028);
  not g26793 (n_9860, n17029);
  and g26794 (n17030, n_9859, n_9860);
  and g26795 (n17031, n16917, n_9773);
  and g26796 (n17032, n_9772, n_9773);
  not g26797 (n_9861, n17031);
  not g26798 (n_9862, n17032);
  and g26799 (n17033, n_9861, n_9862);
  and g26800 (n17034, n16901, n_9759);
  and g26801 (n17035, n_9758, n_9759);
  not g26802 (n_9863, n17034);
  not g26803 (n_9864, n17035);
  and g26804 (n17036, n_9863, n_9864);
  not g26805 (n_9865, n16894);
  and g26806 (n17037, n16892, n_9865);
  not g26807 (n_9866, n17037);
  and g26808 (n17038, n_9743, n_9866);
  and g26809 (n17039, n3884, n12531);
  and g26810 (n17040, n3967, n12537);
  and g26811 (n17041, n4046, n12534);
  not g26812 (n_9867, n17040);
  not g26813 (n_9868, n17041);
  and g26814 (n17042, n_9867, n_9868);
  not g26815 (n_9869, n17039);
  and g26816 (n17043, n_9869, n17042);
  and g26817 (n17044, n_750, n17043);
  not g26818 (n_9870, n15255);
  and g26819 (n17045, n_9870, n17043);
  not g26820 (n_9871, n17044);
  not g26821 (n_9872, n17045);
  and g26822 (n17046, n_9871, n_9872);
  not g26823 (n_9873, n17046);
  and g26824 (n17047, \a[26] , n_9873);
  and g26825 (n17048, n_33, n17046);
  not g26826 (n_9874, n17047);
  not g26827 (n_9875, n17048);
  and g26828 (n17049, n_9874, n_9875);
  not g26829 (n_9876, n17049);
  and g26830 (n17050, n17038, n_9876);
  not g26831 (n_9877, n16890);
  and g26832 (n17051, n16888, n_9877);
  not g26833 (n_9878, n17051);
  and g26834 (n17052, n_9739, n_9878);
  and g26835 (n17053, n3884, n12534);
  and g26836 (n17054, n3967, n12540);
  and g26837 (n17055, n4046, n12537);
  not g26838 (n_9879, n17054);
  not g26839 (n_9880, n17055);
  and g26840 (n17056, n_9879, n_9880);
  not g26841 (n_9881, n17053);
  and g26842 (n17057, n_9881, n17056);
  and g26843 (n17058, n_750, n17057);
  and g26844 (n17059, n15096, n17057);
  not g26845 (n_9882, n17058);
  not g26846 (n_9883, n17059);
  and g26847 (n17060, n_9882, n_9883);
  not g26848 (n_9884, n17060);
  and g26849 (n17061, \a[26] , n_9884);
  and g26850 (n17062, n_33, n17060);
  not g26851 (n_9885, n17061);
  not g26852 (n_9886, n17062);
  and g26853 (n17063, n_9885, n_9886);
  not g26854 (n_9887, n17063);
  and g26855 (n17064, n17052, n_9887);
  not g26856 (n_9888, n16886);
  and g26857 (n17065, n16884, n_9888);
  not g26858 (n_9889, n17065);
  and g26859 (n17066, n_9735, n_9889);
  and g26860 (n17067, n3884, n12537);
  and g26861 (n17068, n3967, n12543);
  and g26862 (n17069, n4046, n12540);
  not g26863 (n_9890, n17068);
  not g26864 (n_9891, n17069);
  and g26865 (n17070, n_9890, n_9891);
  not g26866 (n_9892, n17067);
  and g26867 (n17071, n_9892, n17070);
  and g26868 (n17072, n_750, n17071);
  and g26869 (n17073, n15385, n17071);
  not g26870 (n_9893, n17072);
  not g26871 (n_9894, n17073);
  and g26872 (n17074, n_9893, n_9894);
  not g26873 (n_9895, n17074);
  and g26874 (n17075, \a[26] , n_9895);
  and g26875 (n17076, n_33, n17074);
  not g26876 (n_9896, n17075);
  not g26877 (n_9897, n17076);
  and g26878 (n17077, n_9896, n_9897);
  not g26879 (n_9898, n17077);
  and g26880 (n17078, n17066, n_9898);
  not g26881 (n_9899, n16882);
  and g26882 (n17079, n16880, n_9899);
  not g26883 (n_9900, n17079);
  and g26884 (n17080, n_9731, n_9900);
  and g26885 (n17081, n3884, n12540);
  and g26886 (n17082, n3967, n12546);
  and g26887 (n17083, n4046, n12543);
  not g26888 (n_9901, n17082);
  not g26889 (n_9902, n17083);
  and g26890 (n17084, n_9901, n_9902);
  not g26891 (n_9903, n17081);
  and g26892 (n17085, n_9903, n17084);
  and g26893 (n17086, n_750, n17085);
  and g26894 (n17087, n15708, n17085);
  not g26895 (n_9904, n17086);
  not g26896 (n_9905, n17087);
  and g26897 (n17088, n_9904, n_9905);
  not g26898 (n_9906, n17088);
  and g26899 (n17089, \a[26] , n_9906);
  and g26900 (n17090, n_33, n17088);
  not g26901 (n_9907, n17089);
  not g26902 (n_9908, n17090);
  and g26903 (n17091, n_9907, n_9908);
  not g26904 (n_9909, n17091);
  and g26905 (n17092, n17080, n_9909);
  not g26906 (n_9910, n16878);
  and g26907 (n17093, n16876, n_9910);
  not g26908 (n_9911, n17093);
  and g26909 (n17094, n_9727, n_9911);
  and g26910 (n17095, n3884, n12543);
  and g26911 (n17096, n3967, n12549);
  and g26912 (n17097, n4046, n12546);
  not g26913 (n_9912, n17096);
  not g26914 (n_9913, n17097);
  and g26915 (n17098, n_9912, n_9913);
  not g26916 (n_9914, n17095);
  and g26917 (n17099, n_9914, n17098);
  and g26918 (n17100, n_750, n17099);
  and g26919 (n17101, n_9555, n17099);
  not g26920 (n_9915, n17100);
  not g26921 (n_9916, n17101);
  and g26922 (n17102, n_9915, n_9916);
  not g26923 (n_9917, n17102);
  and g26924 (n17103, \a[26] , n_9917);
  and g26925 (n17104, n_33, n17102);
  not g26926 (n_9918, n17103);
  not g26927 (n_9919, n17104);
  and g26928 (n17105, n_9918, n_9919);
  not g26929 (n_9920, n17105);
  and g26930 (n17106, n17094, n_9920);
  and g26931 (n17107, n16752, n16874);
  not g26932 (n_9921, n17107);
  and g26933 (n17108, n_9723, n_9921);
  and g26934 (n17109, n3884, n12546);
  and g26935 (n17110, n3967, n12552);
  and g26936 (n17111, n4046, n12549);
  not g26937 (n_9922, n17110);
  not g26938 (n_9923, n17111);
  and g26939 (n17112, n_9922, n_9923);
  not g26940 (n_9924, n17109);
  and g26941 (n17113, n_9924, n17112);
  and g26942 (n17114, n_750, n17113);
  and g26943 (n17115, n15356, n17113);
  not g26944 (n_9925, n17114);
  not g26945 (n_9926, n17115);
  and g26946 (n17116, n_9925, n_9926);
  not g26947 (n_9927, n17116);
  and g26948 (n17117, \a[26] , n_9927);
  and g26949 (n17118, n_33, n17116);
  not g26950 (n_9928, n17117);
  not g26951 (n_9929, n17118);
  and g26952 (n17119, n_9928, n_9929);
  not g26953 (n_9930, n17119);
  and g26954 (n17120, n17108, n_9930);
  and g26955 (n17121, n16770, n16872);
  not g26956 (n_9931, n17121);
  and g26957 (n17122, n_9720, n_9931);
  and g26958 (n17123, n3967, n12555);
  and g26959 (n17124, n4046, n12552);
  and g26960 (n17125, n3884, n12549);
  not g26961 (n_9932, n17124);
  not g26962 (n_9933, n17125);
  and g26963 (n17126, n_9932, n_9933);
  not g26964 (n_9934, n17123);
  and g26965 (n17127, n_9934, n17126);
  and g26966 (n17128, n_750, n17127);
  and g26967 (n17129, n_9580, n17127);
  not g26968 (n_9935, n17128);
  not g26969 (n_9936, n17129);
  and g26970 (n17130, n_9935, n_9936);
  not g26971 (n_9937, n17130);
  and g26972 (n17131, \a[26] , n_9937);
  and g26973 (n17132, n_33, n17130);
  not g26974 (n_9938, n17131);
  not g26975 (n_9939, n17132);
  and g26976 (n17133, n_9938, n_9939);
  not g26977 (n_9940, n17133);
  and g26978 (n17134, n17122, n_9940);
  and g26979 (n17135, n16788, n16870);
  not g26980 (n_9941, n17135);
  and g26981 (n17136, n_9717, n_9941);
  and g26982 (n17137, n3967, n12558);
  and g26983 (n17138, n3884, n12552);
  and g26984 (n17139, n4046, n12555);
  not g26985 (n_9942, n17138);
  not g26986 (n_9943, n17139);
  and g26987 (n17140, n_9942, n_9943);
  not g26988 (n_9944, n17137);
  and g26989 (n17141, n_9944, n17140);
  and g26990 (n17142, n_750, n17141);
  and g26991 (n17143, n15791, n17141);
  not g26992 (n_9945, n17142);
  not g26993 (n_9946, n17143);
  and g26994 (n17144, n_9945, n_9946);
  not g26995 (n_9947, n17144);
  and g26996 (n17145, \a[26] , n_9947);
  and g26997 (n17146, n_33, n17144);
  not g26998 (n_9948, n17145);
  not g26999 (n_9949, n17146);
  and g27000 (n17147, n_9948, n_9949);
  not g27001 (n_9950, n17147);
  and g27002 (n17148, n17136, n_9950);
  and g27003 (n17149, n16806, n16868);
  not g27004 (n_9951, n17149);
  and g27005 (n17150, n_9714, n_9951);
  and g27006 (n17151, n4046, n12558);
  and g27007 (n17152, n3884, n12555);
  and g27008 (n17153, n3967, n12561);
  not g27009 (n_9952, n17152);
  not g27010 (n_9953, n17153);
  and g27011 (n17154, n_9952, n_9953);
  not g27012 (n_9954, n17151);
  and g27013 (n17155, n_9954, n17154);
  and g27014 (n17156, n_750, n17155);
  and g27015 (n17157, n15816, n17155);
  not g27016 (n_9955, n17156);
  not g27017 (n_9956, n17157);
  and g27018 (n17158, n_9955, n_9956);
  not g27019 (n_9957, n17158);
  and g27020 (n17159, \a[26] , n_9957);
  and g27021 (n17160, n_33, n17158);
  not g27022 (n_9958, n17159);
  not g27023 (n_9959, n17160);
  and g27024 (n17161, n_9958, n_9959);
  not g27025 (n_9960, n17161);
  and g27026 (n17162, n17150, n_9960);
  and g27027 (n17163, n_9709, n_9711);
  and g27028 (n17164, n_9710, n_9711);
  not g27029 (n_9961, n17163);
  not g27030 (n_9962, n17164);
  and g27031 (n17165, n_9961, n_9962);
  and g27032 (n17166, n3967, n12564);
  and g27033 (n17167, n4046, n12561);
  and g27034 (n17168, n3884, n12558);
  not g27035 (n_9963, n17167);
  not g27036 (n_9964, n17168);
  and g27037 (n17169, n_9963, n_9964);
  not g27038 (n_9965, n17166);
  and g27039 (n17170, n_9965, n17169);
  and g27040 (n17171, n_750, n17170);
  not g27041 (n_9966, n15847);
  and g27042 (n17172, n_9966, n17170);
  not g27043 (n_9967, n17171);
  not g27044 (n_9968, n17172);
  and g27045 (n17173, n_9967, n_9968);
  not g27046 (n_9969, n17173);
  and g27047 (n17174, \a[26] , n_9969);
  and g27048 (n17175, n_33, n17173);
  not g27049 (n_9970, n17174);
  not g27050 (n_9971, n17175);
  and g27051 (n17176, n_9970, n_9971);
  not g27052 (n_9972, n17165);
  not g27053 (n_9973, n17176);
  and g27054 (n17177, n_9972, n_9973);
  and g27055 (n17178, n4046, n12564);
  and g27056 (n17179, n3884, n12561);
  and g27057 (n17180, n3967, n12567);
  and g27063 (n17183, n4050, n_8997);
  not g27066 (n_9978, n17184);
  and g27067 (n17185, \a[26] , n_9978);
  not g27068 (n_9979, n17185);
  and g27069 (n17186, n_9978, n_9979);
  and g27070 (n17187, \a[26] , n_9979);
  not g27071 (n_9980, n17186);
  not g27072 (n_9981, n17187);
  and g27073 (n17188, n_9980, n_9981);
  and g27074 (n17189, n16861, n16864);
  not g27075 (n_9982, n17189);
  and g27076 (n17190, n_9708, n_9982);
  not g27077 (n_9983, n17188);
  and g27078 (n17191, n_9983, n17190);
  not g27079 (n_9984, n17191);
  and g27080 (n17192, n_9983, n_9984);
  and g27081 (n17193, n17190, n_9984);
  not g27082 (n_9985, n17192);
  not g27083 (n_9986, n17193);
  and g27084 (n17194, n_9985, n_9986);
  and g27085 (n17195, n3967, n12571);
  and g27086 (n17196, n4046, n12567);
  and g27087 (n17197, n3884, n12564);
  and g27093 (n17200, n4050, n_9006);
  not g27096 (n_9991, n17201);
  and g27097 (n17202, \a[26] , n_9991);
  not g27098 (n_9992, n17202);
  and g27099 (n17203, n_9991, n_9992);
  and g27100 (n17204, \a[26] , n_9992);
  not g27101 (n_9993, n17203);
  not g27102 (n_9994, n17204);
  and g27103 (n17205, n_9993, n_9994);
  not g27104 (n_9995, n16837);
  and g27105 (n17206, n_9995, n16848);
  not g27106 (n_9996, n17206);
  and g27107 (n17207, n_9702, n_9996);
  not g27108 (n_9997, n17205);
  and g27109 (n17208, n_9997, n17207);
  not g27110 (n_9998, n17208);
  and g27111 (n17209, n_9997, n_9998);
  and g27112 (n17210, n17207, n_9998);
  not g27113 (n_9999, n17209);
  not g27114 (n_10000, n17210);
  and g27115 (n17211, n_9999, n_10000);
  not g27116 (n_10001, n16836);
  and g27117 (n17212, n16834, n_10001);
  not g27118 (n_10002, n17212);
  and g27119 (n17213, n_9995, n_10002);
  and g27120 (n17214, n3967, n12574);
  and g27121 (n17215, n3884, n12567);
  and g27122 (n17216, n4046, n12571);
  not g27123 (n_10003, n17215);
  not g27124 (n_10004, n17216);
  and g27125 (n17217, n_10003, n_10004);
  not g27126 (n_10005, n17214);
  and g27127 (n17218, n_10005, n17217);
  and g27128 (n17219, n_750, n17218);
  not g27129 (n_10006, n15989);
  and g27130 (n17220, n_10006, n17218);
  not g27131 (n_10007, n17219);
  not g27132 (n_10008, n17220);
  and g27133 (n17221, n_10007, n_10008);
  not g27134 (n_10009, n17221);
  and g27135 (n17222, \a[26] , n_10009);
  and g27136 (n17223, n_33, n17221);
  not g27137 (n_10010, n17222);
  not g27138 (n_10011, n17223);
  and g27139 (n17224, n_10010, n_10011);
  not g27140 (n_10012, n17224);
  and g27141 (n17225, n17213, n_10012);
  and g27142 (n17226, n3884, n12577);
  and g27143 (n17227, n4046, n_6977);
  not g27144 (n_10013, n17226);
  not g27145 (n_10014, n17227);
  and g27146 (n17228, n_10013, n_10014);
  and g27147 (n17229, n4050, n_9032);
  not g27148 (n_10015, n17229);
  and g27149 (n17230, n17228, n_10015);
  not g27150 (n_10016, n17230);
  and g27151 (n17231, \a[26] , n_10016);
  not g27152 (n_10017, n17231);
  and g27153 (n17232, \a[26] , n_10017);
  and g27154 (n17233, n_10016, n_10017);
  not g27155 (n_10018, n17232);
  not g27156 (n_10019, n17233);
  and g27157 (n17234, n_10018, n_10019);
  and g27158 (n17235, n_559, n_6977);
  not g27159 (n_10020, n17235);
  and g27160 (n17236, \a[26] , n_10020);
  not g27161 (n_10021, n17234);
  and g27162 (n17237, n_10021, n17236);
  and g27163 (n17238, n3967, n_6977);
  and g27164 (n17239, n3884, n12574);
  and g27165 (n17240, n4046, n12577);
  not g27166 (n_10022, n17239);
  not g27167 (n_10023, n17240);
  and g27168 (n17241, n_10022, n_10023);
  not g27169 (n_10024, n17238);
  and g27170 (n17242, n_10024, n17241);
  and g27171 (n17243, n_750, n17242);
  and g27172 (n17244, n16094, n17242);
  not g27173 (n_10025, n17243);
  not g27174 (n_10026, n17244);
  and g27175 (n17245, n_10025, n_10026);
  not g27176 (n_10027, n17245);
  and g27177 (n17246, \a[26] , n_10027);
  and g27178 (n17247, n_33, n17245);
  not g27179 (n_10028, n17246);
  not g27180 (n_10029, n17247);
  and g27181 (n17248, n_10028, n_10029);
  not g27182 (n_10030, n17248);
  and g27183 (n17249, n17237, n_10030);
  and g27184 (n17250, n16835, n17249);
  not g27185 (n_10031, n17250);
  and g27186 (n17251, n17249, n_10031);
  and g27187 (n17252, n16835, n_10031);
  not g27188 (n_10032, n17251);
  not g27189 (n_10033, n17252);
  and g27190 (n17253, n_10032, n_10033);
  and g27191 (n17254, n3967, n12577);
  and g27192 (n17255, n3884, n12571);
  and g27193 (n17256, n4046, n12574);
  and g27199 (n17259, n4050, n16013);
  not g27202 (n_10038, n17260);
  and g27203 (n17261, \a[26] , n_10038);
  not g27204 (n_10039, n17261);
  and g27205 (n17262, \a[26] , n_10039);
  and g27206 (n17263, n_10038, n_10039);
  not g27207 (n_10040, n17262);
  not g27208 (n_10041, n17263);
  and g27209 (n17264, n_10040, n_10041);
  not g27210 (n_10042, n17253);
  not g27211 (n_10043, n17264);
  and g27212 (n17265, n_10042, n_10043);
  not g27213 (n_10044, n17265);
  and g27214 (n17266, n_10031, n_10044);
  not g27215 (n_10045, n17213);
  and g27216 (n17267, n_10045, n17224);
  not g27217 (n_10046, n17225);
  not g27218 (n_10047, n17267);
  and g27219 (n17268, n_10046, n_10047);
  not g27220 (n_10048, n17266);
  and g27221 (n17269, n_10048, n17268);
  not g27222 (n_10049, n17269);
  and g27223 (n17270, n_10046, n_10049);
  not g27224 (n_10050, n17211);
  not g27225 (n_10051, n17270);
  and g27226 (n17271, n_10050, n_10051);
  not g27227 (n_10052, n17271);
  and g27228 (n17272, n_9998, n_10052);
  not g27229 (n_10053, n17194);
  not g27230 (n_10054, n17272);
  and g27231 (n17273, n_10053, n_10054);
  not g27232 (n_10055, n17273);
  and g27233 (n17274, n_9984, n_10055);
  not g27234 (n_10056, n17177);
  and g27235 (n17275, n_9972, n_10056);
  and g27236 (n17276, n_9973, n_10056);
  not g27237 (n_10057, n17275);
  not g27238 (n_10058, n17276);
  and g27239 (n17277, n_10057, n_10058);
  not g27240 (n_10059, n17274);
  not g27241 (n_10060, n17277);
  and g27242 (n17278, n_10059, n_10060);
  not g27243 (n_10061, n17278);
  and g27244 (n17279, n_10056, n_10061);
  not g27245 (n_10062, n17162);
  and g27246 (n17280, n17150, n_10062);
  and g27247 (n17281, n_9960, n_10062);
  not g27248 (n_10063, n17280);
  not g27249 (n_10064, n17281);
  and g27250 (n17282, n_10063, n_10064);
  not g27251 (n_10065, n17279);
  not g27252 (n_10066, n17282);
  and g27253 (n17283, n_10065, n_10066);
  not g27254 (n_10067, n17283);
  and g27255 (n17284, n_10062, n_10067);
  not g27256 (n_10068, n17148);
  and g27257 (n17285, n17136, n_10068);
  and g27258 (n17286, n_9950, n_10068);
  not g27259 (n_10069, n17285);
  not g27260 (n_10070, n17286);
  and g27261 (n17287, n_10069, n_10070);
  not g27262 (n_10071, n17284);
  not g27263 (n_10072, n17287);
  and g27264 (n17288, n_10071, n_10072);
  not g27265 (n_10073, n17288);
  and g27266 (n17289, n_10068, n_10073);
  not g27267 (n_10074, n17134);
  and g27268 (n17290, n17122, n_10074);
  and g27269 (n17291, n_9940, n_10074);
  not g27270 (n_10075, n17290);
  not g27271 (n_10076, n17291);
  and g27272 (n17292, n_10075, n_10076);
  not g27273 (n_10077, n17289);
  not g27274 (n_10078, n17292);
  and g27275 (n17293, n_10077, n_10078);
  not g27276 (n_10079, n17293);
  and g27277 (n17294, n_10074, n_10079);
  not g27278 (n_10080, n17120);
  and g27279 (n17295, n17108, n_10080);
  and g27280 (n17296, n_9930, n_10080);
  not g27281 (n_10081, n17295);
  not g27282 (n_10082, n17296);
  and g27283 (n17297, n_10081, n_10082);
  not g27284 (n_10083, n17294);
  not g27285 (n_10084, n17297);
  and g27286 (n17298, n_10083, n_10084);
  not g27287 (n_10085, n17298);
  and g27288 (n17299, n_10080, n_10085);
  not g27289 (n_10086, n17106);
  and g27290 (n17300, n17094, n_10086);
  and g27291 (n17301, n_9920, n_10086);
  not g27292 (n_10087, n17300);
  not g27293 (n_10088, n17301);
  and g27294 (n17302, n_10087, n_10088);
  not g27295 (n_10089, n17299);
  not g27296 (n_10090, n17302);
  and g27297 (n17303, n_10089, n_10090);
  not g27298 (n_10091, n17303);
  and g27299 (n17304, n_10086, n_10091);
  not g27300 (n_10092, n17092);
  and g27301 (n17305, n17080, n_10092);
  and g27302 (n17306, n_9909, n_10092);
  not g27303 (n_10093, n17305);
  not g27304 (n_10094, n17306);
  and g27305 (n17307, n_10093, n_10094);
  not g27306 (n_10095, n17304);
  not g27307 (n_10096, n17307);
  and g27308 (n17308, n_10095, n_10096);
  not g27309 (n_10097, n17308);
  and g27310 (n17309, n_10092, n_10097);
  not g27311 (n_10098, n17078);
  and g27312 (n17310, n17066, n_10098);
  and g27313 (n17311, n_9898, n_10098);
  not g27314 (n_10099, n17310);
  not g27315 (n_10100, n17311);
  and g27316 (n17312, n_10099, n_10100);
  not g27317 (n_10101, n17309);
  not g27318 (n_10102, n17312);
  and g27319 (n17313, n_10101, n_10102);
  not g27320 (n_10103, n17313);
  and g27321 (n17314, n_10098, n_10103);
  not g27322 (n_10104, n17064);
  and g27323 (n17315, n17052, n_10104);
  and g27324 (n17316, n_9887, n_10104);
  not g27325 (n_10105, n17315);
  not g27326 (n_10106, n17316);
  and g27327 (n17317, n_10105, n_10106);
  not g27328 (n_10107, n17314);
  not g27329 (n_10108, n17317);
  and g27330 (n17318, n_10107, n_10108);
  not g27331 (n_10109, n17318);
  and g27332 (n17319, n_10104, n_10109);
  not g27333 (n_10110, n17038);
  and g27334 (n17320, n_10110, n17049);
  not g27335 (n_10111, n17050);
  not g27336 (n_10112, n17320);
  and g27337 (n17321, n_10111, n_10112);
  not g27338 (n_10113, n17319);
  and g27339 (n17322, n_10113, n17321);
  not g27340 (n_10114, n17322);
  and g27341 (n17323, n_10111, n_10114);
  not g27342 (n_10115, n17036);
  not g27343 (n_10116, n17323);
  and g27344 (n17324, n_10115, n_10116);
  and g27345 (n17325, n17036, n17323);
  not g27346 (n_10117, n17324);
  not g27347 (n_10118, n17325);
  and g27348 (n17326, n_10117, n_10118);
  and g27349 (n17327, n4694, n12519);
  and g27350 (n17328, n4533, n12525);
  and g27351 (n17329, n4604, n12522);
  and g27357 (n17332, n4536, n14454);
  not g27360 (n_10123, n17333);
  and g27361 (n17334, \a[23] , n_10123);
  not g27362 (n_10124, n17334);
  and g27363 (n17335, \a[23] , n_10124);
  and g27364 (n17336, n_10123, n_10124);
  not g27365 (n_10125, n17335);
  not g27366 (n_10126, n17336);
  and g27367 (n17337, n_10125, n_10126);
  not g27368 (n_10127, n17337);
  and g27369 (n17338, n17326, n_10127);
  not g27370 (n_10128, n17338);
  and g27371 (n17339, n_10117, n_10128);
  not g27372 (n_10129, n17033);
  not g27373 (n_10130, n17339);
  and g27374 (n17340, n_10129, n_10130);
  and g27375 (n17341, n17033, n17339);
  not g27376 (n_10131, n17340);
  not g27377 (n_10132, n17341);
  and g27378 (n17342, n_10131, n_10132);
  and g27379 (n17343, n5496, n12508);
  and g27380 (n17344, n4935, n12511);
  and g27381 (n17345, n5407, n12513);
  and g27387 (n17348, n4938, n13863);
  not g27390 (n_10137, n17349);
  and g27391 (n17350, \a[20] , n_10137);
  not g27392 (n_10138, n17350);
  and g27393 (n17351, \a[20] , n_10138);
  and g27394 (n17352, n_10137, n_10138);
  not g27395 (n_10139, n17351);
  not g27396 (n_10140, n17352);
  and g27397 (n17353, n_10139, n_10140);
  not g27398 (n_10141, n17353);
  and g27399 (n17354, n17342, n_10141);
  not g27400 (n_10142, n17354);
  and g27401 (n17355, n_10131, n_10142);
  not g27402 (n_10143, n17030);
  not g27403 (n_10144, n17355);
  and g27404 (n17356, n_10143, n_10144);
  and g27405 (n17357, n17030, n17355);
  not g27406 (n_10145, n17356);
  not g27407 (n_10146, n17357);
  and g27408 (n17358, n_10145, n_10146);
  and g27409 (n17359, n6233, n12769);
  and g27410 (n17360, n5663, n12370);
  and g27411 (n17361, n5939, n12502);
  and g27417 (n17364, n5666, n12999);
  not g27420 (n_10151, n17365);
  and g27421 (n17366, \a[17] , n_10151);
  not g27422 (n_10152, n17366);
  and g27423 (n17367, \a[17] , n_10152);
  and g27424 (n17368, n_10151, n_10152);
  not g27425 (n_10153, n17367);
  not g27426 (n_10154, n17368);
  and g27427 (n17369, n_10153, n_10154);
  not g27428 (n_10155, n17369);
  and g27429 (n17370, n17358, n_10155);
  not g27430 (n_10156, n17370);
  and g27431 (n17371, n_10145, n_10156);
  not g27432 (n_10157, n17027);
  not g27433 (n_10158, n17371);
  and g27434 (n17372, n_10157, n_10158);
  not g27435 (n_10159, n17372);
  and g27436 (n17373, n_9856, n_10159);
  not g27437 (n_10160, n17010);
  not g27438 (n_10161, n17373);
  and g27439 (n17374, n_10160, n_10161);
  and g27440 (n17375, n17010, n17373);
  not g27441 (n_10162, n17374);
  not g27442 (n_10163, n17375);
  and g27443 (n17376, n_10162, n_10163);
  and g27444 (n17377, n7101, n13515);
  and g27445 (n17378, n6402, n13518);
  and g27446 (n17379, n6951, n13521);
  and g27452 (n17382, n6397, n13541);
  not g27455 (n_10168, n17383);
  and g27456 (n17384, \a[14] , n_10168);
  not g27457 (n_10169, n17384);
  and g27458 (n17385, \a[14] , n_10169);
  and g27459 (n17386, n_10168, n_10169);
  not g27460 (n_10170, n17385);
  not g27461 (n_10171, n17386);
  and g27462 (n17387, n_10170, n_10171);
  not g27463 (n_10172, n17387);
  and g27464 (n17388, n17376, n_10172);
  not g27465 (n_10173, n17388);
  and g27466 (n17389, n_10162, n_10173);
  not g27467 (n_10174, n17007);
  not g27468 (n_10175, n17389);
  and g27469 (n17390, n_10174, n_10175);
  and g27470 (n17391, n17007, n17389);
  not g27471 (n_10176, n17390);
  not g27472 (n_10177, n17391);
  and g27473 (n17392, n_10176, n_10177);
  and g27474 (n17393, n7983, n_7540);
  and g27475 (n17394, n7291, n13630);
  and g27476 (n17395, n7632, n13633);
  and g27482 (n17398, n7294, n_7563);
  not g27485 (n_10182, n17399);
  and g27486 (n17400, \a[11] , n_10182);
  not g27487 (n_10183, n17400);
  and g27488 (n17401, \a[11] , n_10183);
  and g27489 (n17402, n_10182, n_10183);
  not g27490 (n_10184, n17401);
  not g27491 (n_10185, n17402);
  and g27492 (n17403, n_10184, n_10185);
  not g27493 (n_10186, n17403);
  and g27494 (n17404, n17392, n_10186);
  not g27495 (n_10187, n17404);
  and g27496 (n17405, n_10176, n_10187);
  and g27497 (n17406, n7983, n13941);
  and g27498 (n17407, n7291, n13633);
  and g27499 (n17408, n7632, n_7540);
  and g27505 (n17411, n7294, n14136);
  not g27508 (n_10192, n17412);
  and g27509 (n17413, \a[11] , n_10192);
  not g27510 (n_10193, n17413);
  and g27511 (n17414, \a[11] , n_10193);
  and g27512 (n17415, n_10192, n_10193);
  not g27513 (n_10194, n17414);
  not g27514 (n_10195, n17415);
  and g27515 (n17416, n_10194, n_10195);
  not g27516 (n_10196, n17405);
  not g27517 (n_10197, n17416);
  and g27518 (n17417, n_10196, n_10197);
  and g27519 (n17418, n16630, n16980);
  not g27520 (n_10198, n17418);
  and g27521 (n17419, n_9821, n_10198);
  not g27522 (n_10199, n17417);
  and g27523 (n17420, n_10196, n_10199);
  and g27524 (n17421, n_10197, n_10199);
  not g27525 (n_10200, n17420);
  not g27526 (n_10201, n17421);
  and g27527 (n17422, n_10200, n_10201);
  not g27528 (n_10202, n17422);
  and g27529 (n17423, n17419, n_10202);
  not g27530 (n_10203, n17423);
  and g27531 (n17424, n_10199, n_10203);
  not g27532 (n_10204, n17004);
  not g27533 (n_10205, n17424);
  and g27534 (n17425, n_10204, n_10205);
  not g27535 (n_10206, n17425);
  and g27536 (n17426, n_10204, n_10206);
  and g27537 (n17427, n_10205, n_10206);
  not g27538 (n_10207, n17426);
  not g27539 (n_10208, n17427);
  and g27540 (n17428, n_10207, n_10208);
  and g27541 (n17429, n17376, n_10173);
  and g27542 (n17430, n_10172, n_10173);
  not g27543 (n_10209, n17429);
  not g27544 (n_10210, n17430);
  and g27545 (n17431, n_10209, n_10210);
  and g27546 (n17432, n17027, n17371);
  not g27547 (n_10211, n17432);
  and g27548 (n17433, n_10159, n_10211);
  and g27549 (n17434, n7101, n13521);
  and g27550 (n17435, n6402, n13491);
  and g27551 (n17436, n6951, n13518);
  and g27557 (n17439, n6397, n_7677);
  not g27560 (n_10216, n17440);
  and g27561 (n17441, \a[14] , n_10216);
  not g27562 (n_10217, n17441);
  and g27563 (n17442, \a[14] , n_10217);
  and g27564 (n17443, n_10216, n_10217);
  not g27565 (n_10218, n17442);
  not g27566 (n_10219, n17443);
  and g27567 (n17444, n_10218, n_10219);
  not g27568 (n_10220, n17444);
  and g27569 (n17445, n17433, n_10220);
  not g27570 (n_10221, n17445);
  and g27571 (n17446, n17433, n_10221);
  and g27572 (n17447, n_10220, n_10221);
  not g27573 (n_10222, n17446);
  not g27574 (n_10223, n17447);
  and g27575 (n17448, n_10222, n_10223);
  and g27576 (n17449, n17358, n_10156);
  and g27577 (n17450, n_10155, n_10156);
  not g27578 (n_10224, n17449);
  not g27579 (n_10225, n17450);
  and g27580 (n17451, n_10224, n_10225);
  and g27581 (n17452, n17342, n_10142);
  and g27582 (n17453, n_10141, n_10142);
  not g27583 (n_10226, n17452);
  not g27584 (n_10227, n17453);
  and g27585 (n17454, n_10226, n_10227);
  and g27586 (n17455, n17326, n_10128);
  and g27587 (n17456, n_10127, n_10128);
  not g27588 (n_10228, n17455);
  not g27589 (n_10229, n17456);
  and g27590 (n17457, n_10228, n_10229);
  and g27591 (n17458, n4694, n12522);
  and g27592 (n17459, n4533, n12528);
  and g27593 (n17460, n4604, n12525);
  and g27599 (n17463, n4536, n14837);
  not g27602 (n_10234, n17464);
  and g27603 (n17465, \a[23] , n_10234);
  not g27604 (n_10235, n17465);
  and g27605 (n17466, n_10234, n_10235);
  and g27606 (n17467, \a[23] , n_10235);
  not g27607 (n_10236, n17466);
  not g27608 (n_10237, n17467);
  and g27609 (n17468, n_10236, n_10237);
  not g27610 (n_10238, n17321);
  and g27611 (n17469, n17319, n_10238);
  not g27612 (n_10239, n17469);
  and g27613 (n17470, n_10114, n_10239);
  not g27614 (n_10240, n17468);
  and g27615 (n17471, n_10240, n17470);
  not g27616 (n_10241, n17471);
  and g27617 (n17472, n_10240, n_10241);
  and g27618 (n17473, n17470, n_10241);
  not g27619 (n_10242, n17472);
  not g27620 (n_10243, n17473);
  and g27621 (n17474, n_10242, n_10243);
  and g27622 (n17475, n4694, n12525);
  and g27623 (n17476, n4533, n12531);
  and g27624 (n17477, n4604, n12528);
  and g27630 (n17480, n4536, n14608);
  not g27633 (n_10248, n17481);
  and g27634 (n17482, \a[23] , n_10248);
  not g27635 (n_10249, n17482);
  and g27636 (n17483, n_10248, n_10249);
  and g27637 (n17484, \a[23] , n_10249);
  not g27638 (n_10250, n17483);
  not g27639 (n_10251, n17484);
  and g27640 (n17485, n_10250, n_10251);
  and g27641 (n17486, n_10107, n_10109);
  and g27642 (n17487, n_10108, n_10109);
  not g27643 (n_10252, n17486);
  not g27644 (n_10253, n17487);
  and g27645 (n17488, n_10252, n_10253);
  not g27646 (n_10254, n17485);
  not g27647 (n_10255, n17488);
  and g27648 (n17489, n_10254, n_10255);
  not g27649 (n_10256, n17489);
  and g27650 (n17490, n_10254, n_10256);
  and g27651 (n17491, n_10255, n_10256);
  not g27652 (n_10257, n17490);
  not g27653 (n_10258, n17491);
  and g27654 (n17492, n_10257, n_10258);
  and g27655 (n17493, n4694, n12528);
  and g27656 (n17494, n4533, n12534);
  and g27657 (n17495, n4604, n12531);
  and g27663 (n17498, n4536, n_8448);
  not g27666 (n_10263, n17499);
  and g27667 (n17500, \a[23] , n_10263);
  not g27668 (n_10264, n17500);
  and g27669 (n17501, n_10263, n_10264);
  and g27670 (n17502, \a[23] , n_10264);
  not g27671 (n_10265, n17501);
  not g27672 (n_10266, n17502);
  and g27673 (n17503, n_10265, n_10266);
  and g27674 (n17504, n_10101, n_10103);
  and g27675 (n17505, n_10102, n_10103);
  not g27676 (n_10267, n17504);
  not g27677 (n_10268, n17505);
  and g27678 (n17506, n_10267, n_10268);
  not g27679 (n_10269, n17503);
  not g27680 (n_10270, n17506);
  and g27681 (n17507, n_10269, n_10270);
  not g27682 (n_10271, n17507);
  and g27683 (n17508, n_10269, n_10271);
  and g27684 (n17509, n_10270, n_10271);
  not g27685 (n_10272, n17508);
  not g27686 (n_10273, n17509);
  and g27687 (n17510, n_10272, n_10273);
  and g27688 (n17511, n4694, n12531);
  and g27689 (n17512, n4533, n12537);
  and g27690 (n17513, n4604, n12534);
  and g27696 (n17516, n4536, n15255);
  not g27699 (n_10278, n17517);
  and g27700 (n17518, \a[23] , n_10278);
  not g27701 (n_10279, n17518);
  and g27702 (n17519, n_10278, n_10279);
  and g27703 (n17520, \a[23] , n_10279);
  not g27704 (n_10280, n17519);
  not g27705 (n_10281, n17520);
  and g27706 (n17521, n_10280, n_10281);
  and g27707 (n17522, n_10095, n_10097);
  and g27708 (n17523, n_10096, n_10097);
  not g27709 (n_10282, n17522);
  not g27710 (n_10283, n17523);
  and g27711 (n17524, n_10282, n_10283);
  not g27712 (n_10284, n17521);
  not g27713 (n_10285, n17524);
  and g27714 (n17525, n_10284, n_10285);
  not g27715 (n_10286, n17525);
  and g27716 (n17526, n_10284, n_10286);
  and g27717 (n17527, n_10285, n_10286);
  not g27718 (n_10287, n17526);
  not g27719 (n_10288, n17527);
  and g27720 (n17528, n_10287, n_10288);
  and g27721 (n17529, n4694, n12534);
  and g27722 (n17530, n4533, n12540);
  and g27723 (n17531, n4604, n12537);
  and g27729 (n17534, n4536, n_8477);
  not g27732 (n_10293, n17535);
  and g27733 (n17536, \a[23] , n_10293);
  not g27734 (n_10294, n17536);
  and g27735 (n17537, n_10293, n_10294);
  and g27736 (n17538, \a[23] , n_10294);
  not g27737 (n_10295, n17537);
  not g27738 (n_10296, n17538);
  and g27739 (n17539, n_10295, n_10296);
  and g27740 (n17540, n_10089, n_10091);
  and g27741 (n17541, n_10090, n_10091);
  not g27742 (n_10297, n17540);
  not g27743 (n_10298, n17541);
  and g27744 (n17542, n_10297, n_10298);
  not g27745 (n_10299, n17539);
  not g27746 (n_10300, n17542);
  and g27747 (n17543, n_10299, n_10300);
  not g27748 (n_10301, n17543);
  and g27749 (n17544, n_10299, n_10301);
  and g27750 (n17545, n_10300, n_10301);
  not g27751 (n_10302, n17544);
  not g27752 (n_10303, n17545);
  and g27753 (n17546, n_10302, n_10303);
  and g27754 (n17547, n4694, n12537);
  and g27755 (n17548, n4533, n12543);
  and g27756 (n17549, n4604, n12540);
  and g27762 (n17552, n4536, n_8659);
  not g27765 (n_10308, n17553);
  and g27766 (n17554, \a[23] , n_10308);
  not g27767 (n_10309, n17554);
  and g27768 (n17555, n_10308, n_10309);
  and g27769 (n17556, \a[23] , n_10309);
  not g27770 (n_10310, n17555);
  not g27771 (n_10311, n17556);
  and g27772 (n17557, n_10310, n_10311);
  and g27773 (n17558, n_10083, n_10085);
  and g27774 (n17559, n_10084, n_10085);
  not g27775 (n_10312, n17558);
  not g27776 (n_10313, n17559);
  and g27777 (n17560, n_10312, n_10313);
  not g27778 (n_10314, n17557);
  not g27779 (n_10315, n17560);
  and g27780 (n17561, n_10314, n_10315);
  not g27781 (n_10316, n17561);
  and g27782 (n17562, n_10314, n_10316);
  and g27783 (n17563, n_10315, n_10316);
  not g27784 (n_10317, n17562);
  not g27785 (n_10318, n17563);
  and g27786 (n17564, n_10317, n_10318);
  and g27787 (n17565, n4694, n12540);
  and g27788 (n17566, n4533, n12546);
  and g27789 (n17567, n4604, n12543);
  and g27795 (n17570, n4536, n_8936);
  not g27798 (n_10323, n17571);
  and g27799 (n17572, \a[23] , n_10323);
  not g27800 (n_10324, n17572);
  and g27801 (n17573, n_10323, n_10324);
  and g27802 (n17574, \a[23] , n_10324);
  not g27803 (n_10325, n17573);
  not g27804 (n_10326, n17574);
  and g27805 (n17575, n_10325, n_10326);
  and g27806 (n17576, n_10077, n_10079);
  and g27807 (n17577, n_10078, n_10079);
  not g27808 (n_10327, n17576);
  not g27809 (n_10328, n17577);
  and g27810 (n17578, n_10327, n_10328);
  not g27811 (n_10329, n17575);
  not g27812 (n_10330, n17578);
  and g27813 (n17579, n_10329, n_10330);
  not g27814 (n_10331, n17579);
  and g27815 (n17580, n_10329, n_10331);
  and g27816 (n17581, n_10330, n_10331);
  not g27817 (n_10332, n17580);
  not g27818 (n_10333, n17581);
  and g27819 (n17582, n_10332, n_10333);
  and g27820 (n17583, n4694, n12543);
  and g27821 (n17584, n4533, n12549);
  and g27822 (n17585, n4604, n12546);
  and g27828 (n17588, n4536, n15724);
  not g27831 (n_10338, n17589);
  and g27832 (n17590, \a[23] , n_10338);
  not g27833 (n_10339, n17590);
  and g27834 (n17591, n_10338, n_10339);
  and g27835 (n17592, \a[23] , n_10339);
  not g27836 (n_10340, n17591);
  not g27837 (n_10341, n17592);
  and g27838 (n17593, n_10340, n_10341);
  and g27839 (n17594, n_10071, n_10073);
  and g27840 (n17595, n_10072, n_10073);
  not g27841 (n_10342, n17594);
  not g27842 (n_10343, n17595);
  and g27843 (n17596, n_10342, n_10343);
  not g27844 (n_10344, n17593);
  not g27845 (n_10345, n17596);
  and g27846 (n17597, n_10344, n_10345);
  not g27847 (n_10346, n17597);
  and g27848 (n17598, n_10344, n_10346);
  and g27849 (n17599, n_10345, n_10346);
  not g27850 (n_10347, n17598);
  not g27851 (n_10348, n17599);
  and g27852 (n17600, n_10347, n_10348);
  and g27853 (n17601, n4694, n12546);
  and g27854 (n17602, n4533, n12552);
  and g27855 (n17603, n4604, n12549);
  and g27861 (n17606, n4536, n_8634);
  not g27864 (n_10353, n17607);
  and g27865 (n17608, \a[23] , n_10353);
  not g27866 (n_10354, n17608);
  and g27867 (n17609, n_10353, n_10354);
  and g27868 (n17610, \a[23] , n_10354);
  not g27869 (n_10355, n17609);
  not g27870 (n_10356, n17610);
  and g27871 (n17611, n_10355, n_10356);
  and g27872 (n17612, n_10065, n_10067);
  and g27873 (n17613, n_10066, n_10067);
  not g27874 (n_10357, n17612);
  not g27875 (n_10358, n17613);
  and g27876 (n17614, n_10357, n_10358);
  not g27877 (n_10359, n17611);
  not g27878 (n_10360, n17614);
  and g27879 (n17615, n_10359, n_10360);
  not g27880 (n_10361, n17615);
  and g27881 (n17616, n_10359, n_10361);
  and g27882 (n17617, n_10360, n_10361);
  not g27883 (n_10362, n17616);
  not g27884 (n_10363, n17617);
  and g27885 (n17618, n_10362, n_10363);
  and g27886 (n17619, n4694, n12549);
  and g27887 (n17620, n4533, n12555);
  and g27888 (n17621, n4604, n12552);
  and g27894 (n17624, n4536, n15764);
  not g27897 (n_10368, n17625);
  and g27898 (n17626, \a[23] , n_10368);
  not g27899 (n_10369, n17626);
  and g27900 (n17627, n_10368, n_10369);
  and g27901 (n17628, \a[23] , n_10369);
  not g27902 (n_10370, n17627);
  not g27903 (n_10371, n17628);
  and g27904 (n17629, n_10370, n_10371);
  and g27905 (n17630, n_10059, n_10061);
  and g27906 (n17631, n_10060, n_10061);
  not g27907 (n_10372, n17630);
  not g27908 (n_10373, n17631);
  and g27909 (n17632, n_10372, n_10373);
  not g27910 (n_10374, n17629);
  not g27911 (n_10375, n17632);
  and g27912 (n17633, n_10374, n_10375);
  not g27913 (n_10376, n17633);
  and g27914 (n17634, n_10374, n_10376);
  and g27915 (n17635, n_10375, n_10376);
  not g27916 (n_10377, n17634);
  not g27917 (n_10378, n17635);
  and g27918 (n17636, n_10377, n_10378);
  and g27919 (n17637, n17194, n17272);
  not g27920 (n_10379, n17637);
  and g27921 (n17638, n_10055, n_10379);
  and g27922 (n17639, n4694, n12552);
  and g27923 (n17640, n4533, n12558);
  and g27924 (n17641, n4604, n12555);
  not g27925 (n_10380, n17640);
  not g27926 (n_10381, n17641);
  and g27927 (n17642, n_10380, n_10381);
  not g27928 (n_10382, n17639);
  and g27929 (n17643, n_10382, n17642);
  and g27930 (n17644, n_732, n17643);
  and g27931 (n17645, n15791, n17643);
  not g27932 (n_10383, n17644);
  not g27933 (n_10384, n17645);
  and g27934 (n17646, n_10383, n_10384);
  not g27935 (n_10385, n17646);
  and g27936 (n17647, \a[23] , n_10385);
  and g27937 (n17648, n_27, n17646);
  not g27938 (n_10386, n17647);
  not g27939 (n_10387, n17648);
  and g27940 (n17649, n_10386, n_10387);
  not g27941 (n_10388, n17649);
  and g27942 (n17650, n17638, n_10388);
  and g27943 (n17651, n17211, n17270);
  not g27944 (n_10389, n17651);
  and g27945 (n17652, n_10052, n_10389);
  and g27946 (n17653, n4694, n12555);
  and g27947 (n17654, n4533, n12561);
  and g27948 (n17655, n4604, n12558);
  not g27949 (n_10390, n17654);
  not g27950 (n_10391, n17655);
  and g27951 (n17656, n_10390, n_10391);
  not g27952 (n_10392, n17653);
  and g27953 (n17657, n_10392, n17656);
  and g27954 (n17658, n_732, n17657);
  and g27955 (n17659, n15816, n17657);
  not g27956 (n_10393, n17658);
  not g27957 (n_10394, n17659);
  and g27958 (n17660, n_10393, n_10394);
  not g27959 (n_10395, n17660);
  and g27960 (n17661, \a[23] , n_10395);
  and g27961 (n17662, n_27, n17660);
  not g27962 (n_10396, n17661);
  not g27963 (n_10397, n17662);
  and g27964 (n17663, n_10396, n_10397);
  not g27965 (n_10398, n17663);
  and g27966 (n17664, n17652, n_10398);
  and g27967 (n17665, n4694, n12558);
  and g27968 (n17666, n4533, n12564);
  and g27969 (n17667, n4604, n12561);
  and g27975 (n17670, n4536, n15847);
  not g27978 (n_10403, n17671);
  and g27979 (n17672, \a[23] , n_10403);
  not g27980 (n_10404, n17672);
  and g27981 (n17673, n_10403, n_10404);
  and g27982 (n17674, \a[23] , n_10404);
  not g27983 (n_10405, n17673);
  not g27984 (n_10406, n17674);
  and g27985 (n17675, n_10405, n_10406);
  not g27986 (n_10407, n17268);
  and g27987 (n17676, n17266, n_10407);
  not g27988 (n_10408, n17676);
  and g27989 (n17677, n_10049, n_10408);
  not g27990 (n_10409, n17675);
  and g27991 (n17678, n_10409, n17677);
  not g27992 (n_10410, n17678);
  and g27993 (n17679, n_10409, n_10410);
  and g27994 (n17680, n17677, n_10410);
  not g27995 (n_10411, n17679);
  not g27996 (n_10412, n17680);
  and g27997 (n17681, n_10411, n_10412);
  and g27998 (n17682, n_10042, n_10044);
  and g27999 (n17683, n_10043, n_10044);
  not g28000 (n_10413, n17682);
  not g28001 (n_10414, n17683);
  and g28002 (n17684, n_10413, n_10414);
  and g28003 (n17685, n4694, n12561);
  and g28004 (n17686, n4533, n12567);
  and g28005 (n17687, n4604, n12564);
  not g28006 (n_10415, n17686);
  not g28007 (n_10416, n17687);
  and g28008 (n17688, n_10415, n_10416);
  not g28009 (n_10417, n17685);
  and g28010 (n17689, n_10417, n17688);
  and g28011 (n17690, n_732, n17689);
  and g28012 (n17691, n15905, n17689);
  not g28013 (n_10418, n17690);
  not g28014 (n_10419, n17691);
  and g28015 (n17692, n_10418, n_10419);
  not g28016 (n_10420, n17692);
  and g28017 (n17693, \a[23] , n_10420);
  and g28018 (n17694, n_27, n17692);
  not g28019 (n_10421, n17693);
  not g28020 (n_10422, n17694);
  and g28021 (n17695, n_10421, n_10422);
  not g28022 (n_10423, n17684);
  not g28023 (n_10424, n17695);
  and g28024 (n17696, n_10423, n_10424);
  and g28025 (n17697, n4694, n12564);
  and g28026 (n17698, n4533, n12571);
  and g28027 (n17699, n4604, n12567);
  and g28033 (n17702, n4536, n_9006);
  not g28036 (n_10429, n17703);
  and g28037 (n17704, \a[23] , n_10429);
  not g28038 (n_10430, n17704);
  and g28039 (n17705, n_10429, n_10430);
  and g28040 (n17706, \a[23] , n_10430);
  not g28041 (n_10431, n17705);
  not g28042 (n_10432, n17706);
  and g28043 (n17707, n_10431, n_10432);
  not g28044 (n_10433, n17237);
  and g28045 (n17708, n_10433, n17248);
  not g28046 (n_10434, n17249);
  not g28047 (n_10435, n17708);
  and g28048 (n17709, n_10434, n_10435);
  not g28049 (n_10436, n17707);
  and g28050 (n17710, n_10436, n17709);
  not g28051 (n_10437, n17710);
  and g28052 (n17711, n_10436, n_10437);
  and g28053 (n17712, n17709, n_10437);
  not g28054 (n_10438, n17711);
  not g28055 (n_10439, n17712);
  and g28056 (n17713, n_10438, n_10439);
  not g28057 (n_10440, n17236);
  and g28058 (n17714, n17234, n_10440);
  not g28059 (n_10441, n17714);
  and g28060 (n17715, n_10433, n_10441);
  and g28061 (n17716, n4694, n12567);
  and g28062 (n17717, n4533, n12574);
  and g28063 (n17718, n4604, n12571);
  not g28064 (n_10442, n17717);
  not g28065 (n_10443, n17718);
  and g28066 (n17719, n_10442, n_10443);
  not g28067 (n_10444, n17716);
  and g28068 (n17720, n_10444, n17719);
  and g28069 (n17721, n_732, n17720);
  and g28070 (n17722, n_10006, n17720);
  not g28071 (n_10445, n17721);
  not g28072 (n_10446, n17722);
  and g28073 (n17723, n_10445, n_10446);
  not g28074 (n_10447, n17723);
  and g28075 (n17724, \a[23] , n_10447);
  and g28076 (n17725, n_27, n17723);
  not g28077 (n_10448, n17724);
  not g28078 (n_10449, n17725);
  and g28079 (n17726, n_10448, n_10449);
  not g28080 (n_10450, n17726);
  and g28081 (n17727, n17715, n_10450);
  and g28082 (n17728, n4604, n_6977);
  and g28083 (n17729, n4694, n12577);
  not g28084 (n_10451, n17728);
  not g28085 (n_10452, n17729);
  and g28086 (n17730, n_10451, n_10452);
  and g28087 (n17731, n4536, n_9032);
  not g28088 (n_10453, n17731);
  and g28089 (n17732, n17730, n_10453);
  not g28090 (n_10454, n17732);
  and g28091 (n17733, \a[23] , n_10454);
  not g28092 (n_10455, n17733);
  and g28093 (n17734, \a[23] , n_10455);
  and g28094 (n17735, n_10454, n_10455);
  not g28095 (n_10456, n17734);
  not g28096 (n_10457, n17735);
  and g28097 (n17736, n_10456, n_10457);
  and g28098 (n17737, n_731, n_6977);
  not g28099 (n_10458, n17737);
  and g28100 (n17738, \a[23] , n_10458);
  not g28101 (n_10459, n17736);
  and g28102 (n17739, n_10459, n17738);
  and g28103 (n17740, n4694, n12574);
  and g28104 (n17741, n4533, n_6977);
  and g28105 (n17742, n4604, n12577);
  not g28106 (n_10460, n17741);
  not g28107 (n_10461, n17742);
  and g28108 (n17743, n_10460, n_10461);
  not g28109 (n_10462, n17740);
  and g28110 (n17744, n_10462, n17743);
  and g28111 (n17745, n_732, n17744);
  and g28112 (n17746, n16094, n17744);
  not g28113 (n_10463, n17745);
  not g28114 (n_10464, n17746);
  and g28115 (n17747, n_10463, n_10464);
  not g28116 (n_10465, n17747);
  and g28117 (n17748, \a[23] , n_10465);
  and g28118 (n17749, n_27, n17747);
  not g28119 (n_10466, n17748);
  not g28120 (n_10467, n17749);
  and g28121 (n17750, n_10466, n_10467);
  not g28122 (n_10468, n17750);
  and g28123 (n17751, n17739, n_10468);
  and g28124 (n17752, n17235, n17751);
  not g28125 (n_10469, n17752);
  and g28126 (n17753, n17751, n_10469);
  and g28127 (n17754, n17235, n_10469);
  not g28128 (n_10470, n17753);
  not g28129 (n_10471, n17754);
  and g28130 (n17755, n_10470, n_10471);
  and g28131 (n17756, n4694, n12571);
  and g28132 (n17757, n4533, n12577);
  and g28133 (n17758, n4604, n12574);
  and g28139 (n17761, n4536, n16013);
  not g28142 (n_10476, n17762);
  and g28143 (n17763, \a[23] , n_10476);
  not g28144 (n_10477, n17763);
  and g28145 (n17764, \a[23] , n_10477);
  and g28146 (n17765, n_10476, n_10477);
  not g28147 (n_10478, n17764);
  not g28148 (n_10479, n17765);
  and g28149 (n17766, n_10478, n_10479);
  not g28150 (n_10480, n17755);
  not g28151 (n_10481, n17766);
  and g28152 (n17767, n_10480, n_10481);
  not g28153 (n_10482, n17767);
  and g28154 (n17768, n_10469, n_10482);
  not g28155 (n_10483, n17715);
  and g28156 (n17769, n_10483, n17726);
  not g28157 (n_10484, n17727);
  not g28158 (n_10485, n17769);
  and g28159 (n17770, n_10484, n_10485);
  not g28160 (n_10486, n17768);
  and g28161 (n17771, n_10486, n17770);
  not g28162 (n_10487, n17771);
  and g28163 (n17772, n_10484, n_10487);
  not g28164 (n_10488, n17713);
  not g28165 (n_10489, n17772);
  and g28166 (n17773, n_10488, n_10489);
  not g28167 (n_10490, n17773);
  and g28168 (n17774, n_10437, n_10490);
  and g28169 (n17775, n17684, n17695);
  not g28170 (n_10491, n17696);
  not g28171 (n_10492, n17775);
  and g28172 (n17776, n_10491, n_10492);
  not g28173 (n_10493, n17774);
  and g28174 (n17777, n_10493, n17776);
  not g28175 (n_10494, n17777);
  and g28176 (n17778, n_10491, n_10494);
  not g28177 (n_10495, n17681);
  not g28178 (n_10496, n17778);
  and g28179 (n17779, n_10495, n_10496);
  not g28180 (n_10497, n17779);
  and g28181 (n17780, n_10410, n_10497);
  not g28182 (n_10498, n17664);
  and g28183 (n17781, n17652, n_10498);
  and g28184 (n17782, n_10398, n_10498);
  not g28185 (n_10499, n17781);
  not g28186 (n_10500, n17782);
  and g28187 (n17783, n_10499, n_10500);
  not g28188 (n_10501, n17780);
  not g28189 (n_10502, n17783);
  and g28190 (n17784, n_10501, n_10502);
  not g28191 (n_10503, n17784);
  and g28192 (n17785, n_10498, n_10503);
  not g28193 (n_10504, n17638);
  and g28194 (n17786, n_10504, n17649);
  not g28195 (n_10505, n17650);
  not g28196 (n_10506, n17786);
  and g28197 (n17787, n_10505, n_10506);
  not g28198 (n_10507, n17785);
  and g28199 (n17788, n_10507, n17787);
  not g28200 (n_10508, n17788);
  and g28201 (n17789, n_10505, n_10508);
  not g28202 (n_10509, n17636);
  not g28203 (n_10510, n17789);
  and g28204 (n17790, n_10509, n_10510);
  not g28205 (n_10511, n17790);
  and g28206 (n17791, n_10376, n_10511);
  not g28207 (n_10512, n17618);
  not g28208 (n_10513, n17791);
  and g28209 (n17792, n_10512, n_10513);
  not g28210 (n_10514, n17792);
  and g28211 (n17793, n_10361, n_10514);
  not g28212 (n_10515, n17600);
  not g28213 (n_10516, n17793);
  and g28214 (n17794, n_10515, n_10516);
  not g28215 (n_10517, n17794);
  and g28216 (n17795, n_10346, n_10517);
  not g28217 (n_10518, n17582);
  not g28218 (n_10519, n17795);
  and g28219 (n17796, n_10518, n_10519);
  not g28220 (n_10520, n17796);
  and g28221 (n17797, n_10331, n_10520);
  not g28222 (n_10521, n17564);
  not g28223 (n_10522, n17797);
  and g28224 (n17798, n_10521, n_10522);
  not g28225 (n_10523, n17798);
  and g28226 (n17799, n_10316, n_10523);
  not g28227 (n_10524, n17546);
  not g28228 (n_10525, n17799);
  and g28229 (n17800, n_10524, n_10525);
  not g28230 (n_10526, n17800);
  and g28231 (n17801, n_10301, n_10526);
  not g28232 (n_10527, n17528);
  not g28233 (n_10528, n17801);
  and g28234 (n17802, n_10527, n_10528);
  not g28235 (n_10529, n17802);
  and g28236 (n17803, n_10286, n_10529);
  not g28237 (n_10530, n17510);
  not g28238 (n_10531, n17803);
  and g28239 (n17804, n_10530, n_10531);
  not g28240 (n_10532, n17804);
  and g28241 (n17805, n_10271, n_10532);
  not g28242 (n_10533, n17492);
  not g28243 (n_10534, n17805);
  and g28244 (n17806, n_10533, n_10534);
  not g28245 (n_10535, n17806);
  and g28246 (n17807, n_10256, n_10535);
  not g28247 (n_10536, n17474);
  not g28248 (n_10537, n17807);
  and g28249 (n17808, n_10536, n_10537);
  not g28250 (n_10538, n17808);
  and g28251 (n17809, n_10241, n_10538);
  not g28252 (n_10539, n17457);
  not g28253 (n_10540, n17809);
  and g28254 (n17810, n_10539, n_10540);
  and g28255 (n17811, n17457, n17809);
  not g28256 (n_10541, n17810);
  not g28257 (n_10542, n17811);
  and g28258 (n17812, n_10541, n_10542);
  and g28259 (n17813, n5496, n12513);
  and g28260 (n17814, n4935, n12516);
  and g28261 (n17815, n5407, n12511);
  and g28267 (n17818, n4938, n14177);
  not g28270 (n_10547, n17819);
  and g28271 (n17820, \a[20] , n_10547);
  not g28272 (n_10548, n17820);
  and g28273 (n17821, \a[20] , n_10548);
  and g28274 (n17822, n_10547, n_10548);
  not g28275 (n_10549, n17821);
  not g28276 (n_10550, n17822);
  and g28277 (n17823, n_10549, n_10550);
  not g28278 (n_10551, n17823);
  and g28279 (n17824, n17812, n_10551);
  not g28280 (n_10552, n17824);
  and g28281 (n17825, n_10541, n_10552);
  not g28282 (n_10553, n17454);
  not g28283 (n_10554, n17825);
  and g28284 (n17826, n_10553, n_10554);
  and g28285 (n17827, n17454, n17825);
  not g28286 (n_10555, n17826);
  not g28287 (n_10556, n17827);
  and g28288 (n17828, n_10555, n_10556);
  and g28289 (n17829, n6233, n12502);
  and g28290 (n17830, n5663, n12505);
  and g28291 (n17831, n5939, n12370);
  and g28297 (n17834, n5666, n_7594);
  not g28300 (n_10561, n17835);
  and g28301 (n17836, \a[17] , n_10561);
  not g28302 (n_10562, n17836);
  and g28303 (n17837, \a[17] , n_10562);
  and g28304 (n17838, n_10561, n_10562);
  not g28305 (n_10563, n17837);
  not g28306 (n_10564, n17838);
  and g28307 (n17839, n_10563, n_10564);
  not g28308 (n_10565, n17839);
  and g28309 (n17840, n17828, n_10565);
  not g28310 (n_10566, n17840);
  and g28311 (n17841, n_10555, n_10566);
  not g28312 (n_10567, n17451);
  not g28313 (n_10568, n17841);
  and g28314 (n17842, n_10567, n_10568);
  and g28315 (n17843, n17451, n17841);
  not g28316 (n_10569, n17842);
  not g28317 (n_10570, n17843);
  and g28318 (n17844, n_10569, n_10570);
  and g28319 (n17845, n7101, n13518);
  and g28320 (n17846, n6402, n12889);
  and g28321 (n17847, n6951, n13491);
  and g28327 (n17850, n6397, n13584);
  not g28330 (n_10575, n17851);
  and g28331 (n17852, \a[14] , n_10575);
  not g28332 (n_10576, n17852);
  and g28333 (n17853, \a[14] , n_10576);
  and g28334 (n17854, n_10575, n_10576);
  not g28335 (n_10577, n17853);
  not g28336 (n_10578, n17854);
  and g28337 (n17855, n_10577, n_10578);
  not g28338 (n_10579, n17855);
  and g28339 (n17856, n17844, n_10579);
  not g28340 (n_10580, n17856);
  and g28341 (n17857, n_10569, n_10580);
  not g28342 (n_10581, n17448);
  not g28343 (n_10582, n17857);
  and g28344 (n17858, n_10581, n_10582);
  not g28345 (n_10583, n17858);
  and g28346 (n17859, n_10221, n_10583);
  not g28347 (n_10584, n17431);
  not g28348 (n_10585, n17859);
  and g28349 (n17860, n_10584, n_10585);
  and g28350 (n17861, n17431, n17859);
  not g28351 (n_10586, n17860);
  not g28352 (n_10587, n17861);
  and g28353 (n17862, n_10586, n_10587);
  and g28354 (n17863, n7983, n13633);
  and g28355 (n17864, n7291, n13597);
  and g28356 (n17865, n7632, n13630);
  and g28362 (n17868, n7294, n13929);
  not g28365 (n_10592, n17869);
  and g28366 (n17870, \a[11] , n_10592);
  not g28367 (n_10593, n17870);
  and g28368 (n17871, \a[11] , n_10593);
  and g28369 (n17872, n_10592, n_10593);
  not g28370 (n_10594, n17871);
  not g28371 (n_10595, n17872);
  and g28372 (n17873, n_10594, n_10595);
  not g28373 (n_10596, n17873);
  and g28374 (n17874, n17862, n_10596);
  not g28375 (n_10597, n17874);
  and g28376 (n17875, n_10586, n_10597);
  not g28377 (n_10598, n14590);
  and g28378 (n17876, n_7417, n_10598);
  and g28379 (n17877, n8418, n13941);
  not g28380 (n_10599, n17876);
  not g28381 (n_10600, n17877);
  and g28382 (n17878, n_10599, n_10600);
  and g28383 (n17879, n_3428, n17878);
  and g28384 (n17880, n13951, n17878);
  not g28385 (n_10601, n17879);
  not g28386 (n_10602, n17880);
  and g28387 (n17881, n_10601, n_10602);
  not g28388 (n_10603, n17881);
  and g28389 (n17882, \a[8] , n_10603);
  and g28390 (n17883, n_1106, n17881);
  not g28391 (n_10604, n17882);
  not g28392 (n_10605, n17883);
  and g28393 (n17884, n_10604, n_10605);
  not g28394 (n_10606, n17875);
  not g28395 (n_10607, n17884);
  and g28396 (n17885, n_10606, n_10607);
  and g28397 (n17886, n17392, n_10187);
  and g28398 (n17887, n_10186, n_10187);
  not g28399 (n_10608, n17886);
  not g28400 (n_10609, n17887);
  and g28401 (n17888, n_10608, n_10609);
  and g28402 (n17889, n17875, n17884);
  not g28403 (n_10610, n17885);
  not g28404 (n_10611, n17889);
  and g28405 (n17890, n_10610, n_10611);
  not g28406 (n_10612, n17888);
  and g28407 (n17891, n_10612, n17890);
  not g28408 (n_10613, n17891);
  and g28409 (n17892, n_10610, n_10613);
  not g28410 (n_10614, n17419);
  and g28411 (n17893, n_10614, n17422);
  not g28412 (n_10615, n17893);
  and g28413 (n17894, n_10203, n_10615);
  not g28414 (n_10616, n17892);
  and g28415 (n17895, n_10616, n17894);
  and g28416 (n17896, n_10612, n_10613);
  and g28417 (n17897, n17890, n_10613);
  not g28418 (n_10617, n17896);
  not g28419 (n_10618, n17897);
  and g28420 (n17898, n_10617, n_10618);
  and g28421 (n17899, n17862, n_10597);
  and g28422 (n17900, n_10596, n_10597);
  not g28423 (n_10619, n17899);
  not g28424 (n_10620, n17900);
  and g28425 (n17901, n_10619, n_10620);
  and g28426 (n17902, n17448, n17857);
  not g28427 (n_10621, n17902);
  and g28428 (n17903, n_10583, n_10621);
  and g28429 (n17904, n7983, n13630);
  and g28430 (n17905, n7291, n13515);
  and g28431 (n17906, n7632, n13597);
  and g28437 (n17909, n7294, n13976);
  not g28440 (n_10626, n17910);
  and g28441 (n17911, \a[11] , n_10626);
  not g28442 (n_10627, n17911);
  and g28443 (n17912, \a[11] , n_10627);
  and g28444 (n17913, n_10626, n_10627);
  not g28445 (n_10628, n17912);
  not g28446 (n_10629, n17913);
  and g28447 (n17914, n_10628, n_10629);
  not g28448 (n_10630, n17914);
  and g28449 (n17915, n17903, n_10630);
  not g28450 (n_10631, n17915);
  and g28451 (n17916, n17903, n_10631);
  and g28452 (n17917, n_10630, n_10631);
  not g28453 (n_10632, n17916);
  not g28454 (n_10633, n17917);
  and g28455 (n17918, n_10632, n_10633);
  and g28456 (n17919, n17844, n_10580);
  and g28457 (n17920, n_10579, n_10580);
  not g28458 (n_10634, n17919);
  not g28459 (n_10635, n17920);
  and g28460 (n17921, n_10634, n_10635);
  and g28461 (n17922, n17828, n_10566);
  and g28462 (n17923, n_10565, n_10566);
  not g28463 (n_10636, n17922);
  not g28464 (n_10637, n17923);
  and g28465 (n17924, n_10636, n_10637);
  and g28466 (n17925, n17812, n_10552);
  and g28467 (n17926, n_10551, n_10552);
  not g28468 (n_10638, n17925);
  not g28469 (n_10639, n17926);
  and g28470 (n17927, n_10638, n_10639);
  and g28471 (n17928, n17474, n17807);
  not g28472 (n_10640, n17928);
  and g28473 (n17929, n_10538, n_10640);
  and g28474 (n17930, n5496, n12511);
  and g28475 (n17931, n4935, n12519);
  and g28476 (n17932, n5407, n12516);
  not g28477 (n_10641, n17931);
  not g28478 (n_10642, n17932);
  and g28479 (n17933, n_10641, n_10642);
  not g28480 (n_10643, n17930);
  and g28481 (n17934, n_10643, n17933);
  and g28482 (n17935, n_1011, n17934);
  and g28483 (n17936, n14233, n17934);
  not g28484 (n_10644, n17935);
  not g28485 (n_10645, n17936);
  and g28486 (n17937, n_10644, n_10645);
  not g28487 (n_10646, n17937);
  and g28488 (n17938, \a[20] , n_10646);
  and g28489 (n17939, n_435, n17937);
  not g28490 (n_10647, n17938);
  not g28491 (n_10648, n17939);
  and g28492 (n17940, n_10647, n_10648);
  not g28493 (n_10649, n17940);
  and g28494 (n17941, n17929, n_10649);
  and g28495 (n17942, n17492, n17805);
  not g28496 (n_10650, n17942);
  and g28497 (n17943, n_10535, n_10650);
  and g28498 (n17944, n5496, n12516);
  and g28499 (n17945, n4935, n12522);
  and g28500 (n17946, n5407, n12519);
  not g28501 (n_10651, n17945);
  not g28502 (n_10652, n17946);
  and g28503 (n17947, n_10651, n_10652);
  not g28504 (n_10653, n17944);
  and g28505 (n17948, n_10653, n17947);
  and g28506 (n17949, n_1011, n17948);
  and g28507 (n17950, n14443, n17948);
  not g28508 (n_10654, n17949);
  not g28509 (n_10655, n17950);
  and g28510 (n17951, n_10654, n_10655);
  not g28511 (n_10656, n17951);
  and g28512 (n17952, \a[20] , n_10656);
  and g28513 (n17953, n_435, n17951);
  not g28514 (n_10657, n17952);
  not g28515 (n_10658, n17953);
  and g28516 (n17954, n_10657, n_10658);
  not g28517 (n_10659, n17954);
  and g28518 (n17955, n17943, n_10659);
  and g28519 (n17956, n17510, n17803);
  not g28520 (n_10660, n17956);
  and g28521 (n17957, n_10532, n_10660);
  and g28522 (n17958, n5496, n12519);
  and g28523 (n17959, n4935, n12525);
  and g28524 (n17960, n5407, n12522);
  not g28525 (n_10661, n17959);
  not g28526 (n_10662, n17960);
  and g28527 (n17961, n_10661, n_10662);
  not g28528 (n_10663, n17958);
  and g28529 (n17962, n_10663, n17961);
  and g28530 (n17963, n_1011, n17962);
  not g28531 (n_10664, n14454);
  and g28532 (n17964, n_10664, n17962);
  not g28533 (n_10665, n17963);
  not g28534 (n_10666, n17964);
  and g28535 (n17965, n_10665, n_10666);
  not g28536 (n_10667, n17965);
  and g28537 (n17966, \a[20] , n_10667);
  and g28538 (n17967, n_435, n17965);
  not g28539 (n_10668, n17966);
  not g28540 (n_10669, n17967);
  and g28541 (n17968, n_10668, n_10669);
  not g28542 (n_10670, n17968);
  and g28543 (n17969, n17957, n_10670);
  and g28544 (n17970, n17528, n17801);
  not g28545 (n_10671, n17970);
  and g28546 (n17971, n_10529, n_10671);
  and g28547 (n17972, n5496, n12522);
  and g28548 (n17973, n4935, n12528);
  and g28549 (n17974, n5407, n12525);
  not g28550 (n_10672, n17973);
  not g28551 (n_10673, n17974);
  and g28552 (n17975, n_10672, n_10673);
  not g28553 (n_10674, n17972);
  and g28554 (n17976, n_10674, n17975);
  and g28555 (n17977, n_1011, n17976);
  not g28556 (n_10675, n14837);
  and g28557 (n17978, n_10675, n17976);
  not g28558 (n_10676, n17977);
  not g28559 (n_10677, n17978);
  and g28560 (n17979, n_10676, n_10677);
  not g28561 (n_10678, n17979);
  and g28562 (n17980, \a[20] , n_10678);
  and g28563 (n17981, n_435, n17979);
  not g28564 (n_10679, n17980);
  not g28565 (n_10680, n17981);
  and g28566 (n17982, n_10679, n_10680);
  not g28567 (n_10681, n17982);
  and g28568 (n17983, n17971, n_10681);
  and g28569 (n17984, n17546, n17799);
  not g28570 (n_10682, n17984);
  and g28571 (n17985, n_10526, n_10682);
  and g28572 (n17986, n5496, n12525);
  and g28573 (n17987, n4935, n12531);
  and g28574 (n17988, n5407, n12528);
  not g28575 (n_10683, n17987);
  not g28576 (n_10684, n17988);
  and g28577 (n17989, n_10683, n_10684);
  not g28578 (n_10685, n17986);
  and g28579 (n17990, n_10685, n17989);
  and g28580 (n17991, n_1011, n17990);
  and g28581 (n17992, n_8677, n17990);
  not g28582 (n_10686, n17991);
  not g28583 (n_10687, n17992);
  and g28584 (n17993, n_10686, n_10687);
  not g28585 (n_10688, n17993);
  and g28586 (n17994, \a[20] , n_10688);
  and g28587 (n17995, n_435, n17993);
  not g28588 (n_10689, n17994);
  not g28589 (n_10690, n17995);
  and g28590 (n17996, n_10689, n_10690);
  not g28591 (n_10691, n17996);
  and g28592 (n17997, n17985, n_10691);
  and g28593 (n17998, n17564, n17797);
  not g28594 (n_10692, n17998);
  and g28595 (n17999, n_10523, n_10692);
  and g28596 (n18000, n5496, n12528);
  and g28597 (n18001, n4935, n12534);
  and g28598 (n18002, n5407, n12531);
  not g28599 (n_10693, n18001);
  not g28600 (n_10694, n18002);
  and g28601 (n18003, n_10693, n_10694);
  not g28602 (n_10695, n18000);
  and g28603 (n18004, n_10695, n18003);
  and g28604 (n18005, n_1011, n18004);
  and g28605 (n18006, n15003, n18004);
  not g28606 (n_10696, n18005);
  not g28607 (n_10697, n18006);
  and g28608 (n18007, n_10696, n_10697);
  not g28609 (n_10698, n18007);
  and g28610 (n18008, \a[20] , n_10698);
  and g28611 (n18009, n_435, n18007);
  not g28612 (n_10699, n18008);
  not g28613 (n_10700, n18009);
  and g28614 (n18010, n_10699, n_10700);
  not g28615 (n_10701, n18010);
  and g28616 (n18011, n17999, n_10701);
  and g28617 (n18012, n17582, n17795);
  not g28618 (n_10702, n18012);
  and g28619 (n18013, n_10520, n_10702);
  and g28620 (n18014, n5496, n12531);
  and g28621 (n18015, n4935, n12537);
  and g28622 (n18016, n5407, n12534);
  not g28623 (n_10703, n18015);
  not g28624 (n_10704, n18016);
  and g28625 (n18017, n_10703, n_10704);
  not g28626 (n_10705, n18014);
  and g28627 (n18018, n_10705, n18017);
  and g28628 (n18019, n_1011, n18018);
  and g28629 (n18020, n_9870, n18018);
  not g28630 (n_10706, n18019);
  not g28631 (n_10707, n18020);
  and g28632 (n18021, n_10706, n_10707);
  not g28633 (n_10708, n18021);
  and g28634 (n18022, \a[20] , n_10708);
  and g28635 (n18023, n_435, n18021);
  not g28636 (n_10709, n18022);
  not g28637 (n_10710, n18023);
  and g28638 (n18024, n_10709, n_10710);
  not g28639 (n_10711, n18024);
  and g28640 (n18025, n18013, n_10711);
  and g28641 (n18026, n17600, n17793);
  not g28642 (n_10712, n18026);
  and g28643 (n18027, n_10517, n_10712);
  and g28644 (n18028, n5496, n12534);
  and g28645 (n18029, n4935, n12540);
  and g28646 (n18030, n5407, n12537);
  not g28647 (n_10713, n18029);
  not g28648 (n_10714, n18030);
  and g28649 (n18031, n_10713, n_10714);
  not g28650 (n_10715, n18028);
  and g28651 (n18032, n_10715, n18031);
  and g28652 (n18033, n_1011, n18032);
  and g28653 (n18034, n15096, n18032);
  not g28654 (n_10716, n18033);
  not g28655 (n_10717, n18034);
  and g28656 (n18035, n_10716, n_10717);
  not g28657 (n_10718, n18035);
  and g28658 (n18036, \a[20] , n_10718);
  and g28659 (n18037, n_435, n18035);
  not g28660 (n_10719, n18036);
  not g28661 (n_10720, n18037);
  and g28662 (n18038, n_10719, n_10720);
  not g28663 (n_10721, n18038);
  and g28664 (n18039, n18027, n_10721);
  and g28665 (n18040, n17618, n17791);
  not g28666 (n_10722, n18040);
  and g28667 (n18041, n_10514, n_10722);
  and g28668 (n18042, n5496, n12537);
  and g28669 (n18043, n4935, n12543);
  and g28670 (n18044, n5407, n12540);
  not g28671 (n_10723, n18043);
  not g28672 (n_10724, n18044);
  and g28673 (n18045, n_10723, n_10724);
  not g28674 (n_10725, n18042);
  and g28675 (n18046, n_10725, n18045);
  and g28676 (n18047, n_1011, n18046);
  and g28677 (n18048, n15385, n18046);
  not g28678 (n_10726, n18047);
  not g28679 (n_10727, n18048);
  and g28680 (n18049, n_10726, n_10727);
  not g28681 (n_10728, n18049);
  and g28682 (n18050, \a[20] , n_10728);
  and g28683 (n18051, n_435, n18049);
  not g28684 (n_10729, n18050);
  not g28685 (n_10730, n18051);
  and g28686 (n18052, n_10729, n_10730);
  not g28687 (n_10731, n18052);
  and g28688 (n18053, n18041, n_10731);
  and g28689 (n18054, n17636, n17789);
  not g28690 (n_10732, n18054);
  and g28691 (n18055, n_10511, n_10732);
  and g28692 (n18056, n5496, n12540);
  and g28693 (n18057, n4935, n12546);
  and g28694 (n18058, n5407, n12543);
  not g28695 (n_10733, n18057);
  not g28696 (n_10734, n18058);
  and g28697 (n18059, n_10733, n_10734);
  not g28698 (n_10735, n18056);
  and g28699 (n18060, n_10735, n18059);
  and g28700 (n18061, n_1011, n18060);
  and g28701 (n18062, n15708, n18060);
  not g28702 (n_10736, n18061);
  not g28703 (n_10737, n18062);
  and g28704 (n18063, n_10736, n_10737);
  not g28705 (n_10738, n18063);
  and g28706 (n18064, \a[20] , n_10738);
  and g28707 (n18065, n_435, n18063);
  not g28708 (n_10739, n18064);
  not g28709 (n_10740, n18065);
  and g28710 (n18066, n_10739, n_10740);
  not g28711 (n_10741, n18066);
  and g28712 (n18067, n18055, n_10741);
  and g28713 (n18068, n5496, n12543);
  and g28714 (n18069, n4935, n12549);
  and g28715 (n18070, n5407, n12546);
  and g28721 (n18073, n4938, n15724);
  not g28724 (n_10746, n18074);
  and g28725 (n18075, \a[20] , n_10746);
  not g28726 (n_10747, n18075);
  and g28727 (n18076, n_10746, n_10747);
  and g28728 (n18077, \a[20] , n_10747);
  not g28729 (n_10748, n18076);
  not g28730 (n_10749, n18077);
  and g28731 (n18078, n_10748, n_10749);
  not g28732 (n_10750, n17787);
  and g28733 (n18079, n17785, n_10750);
  not g28734 (n_10751, n18079);
  and g28735 (n18080, n_10508, n_10751);
  not g28736 (n_10752, n18078);
  and g28737 (n18081, n_10752, n18080);
  not g28738 (n_10753, n18081);
  and g28739 (n18082, n_10752, n_10753);
  and g28740 (n18083, n18080, n_10753);
  not g28741 (n_10754, n18082);
  not g28742 (n_10755, n18083);
  and g28743 (n18084, n_10754, n_10755);
  and g28744 (n18085, n5496, n12546);
  and g28745 (n18086, n4935, n12552);
  and g28746 (n18087, n5407, n12549);
  and g28752 (n18090, n4938, n_8634);
  not g28755 (n_10760, n18091);
  and g28756 (n18092, \a[20] , n_10760);
  not g28757 (n_10761, n18092);
  and g28758 (n18093, n_10760, n_10761);
  and g28759 (n18094, \a[20] , n_10761);
  not g28760 (n_10762, n18093);
  not g28761 (n_10763, n18094);
  and g28762 (n18095, n_10762, n_10763);
  and g28763 (n18096, n_10501, n_10503);
  and g28764 (n18097, n_10502, n_10503);
  not g28765 (n_10764, n18096);
  not g28766 (n_10765, n18097);
  and g28767 (n18098, n_10764, n_10765);
  not g28768 (n_10766, n18095);
  not g28769 (n_10767, n18098);
  and g28770 (n18099, n_10766, n_10767);
  not g28771 (n_10768, n18099);
  and g28772 (n18100, n_10766, n_10768);
  and g28773 (n18101, n_10767, n_10768);
  not g28774 (n_10769, n18100);
  not g28775 (n_10770, n18101);
  and g28776 (n18102, n_10769, n_10770);
  and g28777 (n18103, n17681, n17778);
  not g28778 (n_10771, n18103);
  and g28779 (n18104, n_10497, n_10771);
  and g28780 (n18105, n5496, n12549);
  and g28781 (n18106, n4935, n12555);
  and g28782 (n18107, n5407, n12552);
  not g28783 (n_10772, n18106);
  not g28784 (n_10773, n18107);
  and g28785 (n18108, n_10772, n_10773);
  not g28786 (n_10774, n18105);
  and g28787 (n18109, n_10774, n18108);
  and g28788 (n18110, n_1011, n18109);
  and g28789 (n18111, n_9580, n18109);
  not g28790 (n_10775, n18110);
  not g28791 (n_10776, n18111);
  and g28792 (n18112, n_10775, n_10776);
  not g28793 (n_10777, n18112);
  and g28794 (n18113, \a[20] , n_10777);
  and g28795 (n18114, n_435, n18112);
  not g28796 (n_10778, n18113);
  not g28797 (n_10779, n18114);
  and g28798 (n18115, n_10778, n_10779);
  not g28799 (n_10780, n18115);
  and g28800 (n18116, n18104, n_10780);
  not g28801 (n_10781, n17776);
  and g28802 (n18117, n17774, n_10781);
  not g28803 (n_10782, n18117);
  and g28804 (n18118, n_10494, n_10782);
  and g28805 (n18119, n5496, n12552);
  and g28806 (n18120, n4935, n12558);
  and g28807 (n18121, n5407, n12555);
  not g28808 (n_10783, n18120);
  not g28809 (n_10784, n18121);
  and g28810 (n18122, n_10783, n_10784);
  not g28811 (n_10785, n18119);
  and g28812 (n18123, n_10785, n18122);
  and g28813 (n18124, n_1011, n18123);
  and g28814 (n18125, n15791, n18123);
  not g28815 (n_10786, n18124);
  not g28816 (n_10787, n18125);
  and g28817 (n18126, n_10786, n_10787);
  not g28818 (n_10788, n18126);
  and g28819 (n18127, \a[20] , n_10788);
  and g28820 (n18128, n_435, n18126);
  not g28821 (n_10789, n18127);
  not g28822 (n_10790, n18128);
  and g28823 (n18129, n_10789, n_10790);
  not g28824 (n_10791, n18129);
  and g28825 (n18130, n18118, n_10791);
  and g28826 (n18131, n17713, n17772);
  not g28827 (n_10792, n18131);
  and g28828 (n18132, n_10490, n_10792);
  and g28829 (n18133, n5496, n12555);
  and g28830 (n18134, n4935, n12561);
  and g28831 (n18135, n5407, n12558);
  not g28832 (n_10793, n18134);
  not g28833 (n_10794, n18135);
  and g28834 (n18136, n_10793, n_10794);
  not g28835 (n_10795, n18133);
  and g28836 (n18137, n_10795, n18136);
  and g28837 (n18138, n_1011, n18137);
  and g28838 (n18139, n15816, n18137);
  not g28839 (n_10796, n18138);
  not g28840 (n_10797, n18139);
  and g28841 (n18140, n_10796, n_10797);
  not g28842 (n_10798, n18140);
  and g28843 (n18141, \a[20] , n_10798);
  and g28844 (n18142, n_435, n18140);
  not g28845 (n_10799, n18141);
  not g28846 (n_10800, n18142);
  and g28847 (n18143, n_10799, n_10800);
  not g28848 (n_10801, n18143);
  and g28849 (n18144, n18132, n_10801);
  and g28850 (n18145, n5496, n12558);
  and g28851 (n18146, n4935, n12564);
  and g28852 (n18147, n5407, n12561);
  and g28858 (n18150, n4938, n15847);
  not g28861 (n_10806, n18151);
  and g28862 (n18152, \a[20] , n_10806);
  not g28863 (n_10807, n18152);
  and g28864 (n18153, n_10806, n_10807);
  and g28865 (n18154, \a[20] , n_10807);
  not g28866 (n_10808, n18153);
  not g28867 (n_10809, n18154);
  and g28868 (n18155, n_10808, n_10809);
  not g28869 (n_10810, n17770);
  and g28870 (n18156, n17768, n_10810);
  not g28871 (n_10811, n18156);
  and g28872 (n18157, n_10487, n_10811);
  not g28873 (n_10812, n18155);
  and g28874 (n18158, n_10812, n18157);
  not g28875 (n_10813, n18158);
  and g28876 (n18159, n_10812, n_10813);
  and g28877 (n18160, n18157, n_10813);
  not g28878 (n_10814, n18159);
  not g28879 (n_10815, n18160);
  and g28880 (n18161, n_10814, n_10815);
  and g28881 (n18162, n_10480, n_10482);
  and g28882 (n18163, n_10481, n_10482);
  not g28883 (n_10816, n18162);
  not g28884 (n_10817, n18163);
  and g28885 (n18164, n_10816, n_10817);
  and g28886 (n18165, n5496, n12561);
  and g28887 (n18166, n4935, n12567);
  and g28888 (n18167, n5407, n12564);
  not g28889 (n_10818, n18166);
  not g28890 (n_10819, n18167);
  and g28891 (n18168, n_10818, n_10819);
  not g28892 (n_10820, n18165);
  and g28893 (n18169, n_10820, n18168);
  and g28894 (n18170, n_1011, n18169);
  and g28895 (n18171, n15905, n18169);
  not g28896 (n_10821, n18170);
  not g28897 (n_10822, n18171);
  and g28898 (n18172, n_10821, n_10822);
  not g28899 (n_10823, n18172);
  and g28900 (n18173, \a[20] , n_10823);
  and g28901 (n18174, n_435, n18172);
  not g28902 (n_10824, n18173);
  not g28903 (n_10825, n18174);
  and g28904 (n18175, n_10824, n_10825);
  not g28905 (n_10826, n18164);
  not g28906 (n_10827, n18175);
  and g28907 (n18176, n_10826, n_10827);
  and g28908 (n18177, n5496, n12564);
  and g28909 (n18178, n4935, n12571);
  and g28910 (n18179, n5407, n12567);
  and g28916 (n18182, n4938, n_9006);
  not g28919 (n_10832, n18183);
  and g28920 (n18184, \a[20] , n_10832);
  not g28921 (n_10833, n18184);
  and g28922 (n18185, n_10832, n_10833);
  and g28923 (n18186, \a[20] , n_10833);
  not g28924 (n_10834, n18185);
  not g28925 (n_10835, n18186);
  and g28926 (n18187, n_10834, n_10835);
  not g28927 (n_10836, n17739);
  and g28928 (n18188, n_10836, n17750);
  not g28929 (n_10837, n17751);
  not g28930 (n_10838, n18188);
  and g28931 (n18189, n_10837, n_10838);
  not g28932 (n_10839, n18187);
  and g28933 (n18190, n_10839, n18189);
  not g28934 (n_10840, n18190);
  and g28935 (n18191, n_10839, n_10840);
  and g28936 (n18192, n18189, n_10840);
  not g28937 (n_10841, n18191);
  not g28938 (n_10842, n18192);
  and g28939 (n18193, n_10841, n_10842);
  not g28940 (n_10843, n17738);
  and g28941 (n18194, n17736, n_10843);
  not g28942 (n_10844, n18194);
  and g28943 (n18195, n_10836, n_10844);
  and g28944 (n18196, n5496, n12567);
  and g28945 (n18197, n4935, n12574);
  and g28946 (n18198, n5407, n12571);
  not g28947 (n_10845, n18197);
  not g28948 (n_10846, n18198);
  and g28949 (n18199, n_10845, n_10846);
  not g28950 (n_10847, n18196);
  and g28951 (n18200, n_10847, n18199);
  and g28952 (n18201, n_1011, n18200);
  and g28953 (n18202, n_10006, n18200);
  not g28954 (n_10848, n18201);
  not g28955 (n_10849, n18202);
  and g28956 (n18203, n_10848, n_10849);
  not g28957 (n_10850, n18203);
  and g28958 (n18204, \a[20] , n_10850);
  and g28959 (n18205, n_435, n18203);
  not g28960 (n_10851, n18204);
  not g28961 (n_10852, n18205);
  and g28962 (n18206, n_10851, n_10852);
  not g28963 (n_10853, n18206);
  and g28964 (n18207, n18195, n_10853);
  and g28965 (n18208, n5407, n_6977);
  and g28966 (n18209, n5496, n12577);
  not g28967 (n_10854, n18208);
  not g28968 (n_10855, n18209);
  and g28969 (n18210, n_10854, n_10855);
  and g28970 (n18211, n4938, n_9032);
  not g28971 (n_10856, n18211);
  and g28972 (n18212, n18210, n_10856);
  not g28973 (n_10857, n18212);
  and g28974 (n18213, \a[20] , n_10857);
  not g28975 (n_10858, n18213);
  and g28976 (n18214, \a[20] , n_10858);
  and g28977 (n18215, n_10857, n_10858);
  not g28978 (n_10859, n18214);
  not g28979 (n_10860, n18215);
  and g28980 (n18216, n_10859, n_10860);
  and g28981 (n18217, n_1010, n_6977);
  not g28982 (n_10861, n18217);
  and g28983 (n18218, \a[20] , n_10861);
  not g28984 (n_10862, n18216);
  and g28985 (n18219, n_10862, n18218);
  and g28986 (n18220, n5496, n12574);
  and g28987 (n18221, n4935, n_6977);
  and g28988 (n18222, n5407, n12577);
  not g28989 (n_10863, n18221);
  not g28990 (n_10864, n18222);
  and g28991 (n18223, n_10863, n_10864);
  not g28992 (n_10865, n18220);
  and g28993 (n18224, n_10865, n18223);
  and g28994 (n18225, n_1011, n18224);
  and g28995 (n18226, n16094, n18224);
  not g28996 (n_10866, n18225);
  not g28997 (n_10867, n18226);
  and g28998 (n18227, n_10866, n_10867);
  not g28999 (n_10868, n18227);
  and g29000 (n18228, \a[20] , n_10868);
  and g29001 (n18229, n_435, n18227);
  not g29002 (n_10869, n18228);
  not g29003 (n_10870, n18229);
  and g29004 (n18230, n_10869, n_10870);
  not g29005 (n_10871, n18230);
  and g29006 (n18231, n18219, n_10871);
  and g29007 (n18232, n17737, n18231);
  not g29008 (n_10872, n18232);
  and g29009 (n18233, n18231, n_10872);
  and g29010 (n18234, n17737, n_10872);
  not g29011 (n_10873, n18233);
  not g29012 (n_10874, n18234);
  and g29013 (n18235, n_10873, n_10874);
  and g29014 (n18236, n5496, n12571);
  and g29015 (n18237, n4935, n12577);
  and g29016 (n18238, n5407, n12574);
  and g29022 (n18241, n4938, n16013);
  not g29025 (n_10879, n18242);
  and g29026 (n18243, \a[20] , n_10879);
  not g29027 (n_10880, n18243);
  and g29028 (n18244, \a[20] , n_10880);
  and g29029 (n18245, n_10879, n_10880);
  not g29030 (n_10881, n18244);
  not g29031 (n_10882, n18245);
  and g29032 (n18246, n_10881, n_10882);
  not g29033 (n_10883, n18235);
  not g29034 (n_10884, n18246);
  and g29035 (n18247, n_10883, n_10884);
  not g29036 (n_10885, n18247);
  and g29037 (n18248, n_10872, n_10885);
  not g29038 (n_10886, n18195);
  and g29039 (n18249, n_10886, n18206);
  not g29040 (n_10887, n18207);
  not g29041 (n_10888, n18249);
  and g29042 (n18250, n_10887, n_10888);
  not g29043 (n_10889, n18248);
  and g29044 (n18251, n_10889, n18250);
  not g29045 (n_10890, n18251);
  and g29046 (n18252, n_10887, n_10890);
  not g29047 (n_10891, n18193);
  not g29048 (n_10892, n18252);
  and g29049 (n18253, n_10891, n_10892);
  not g29050 (n_10893, n18253);
  and g29051 (n18254, n_10840, n_10893);
  and g29052 (n18255, n18164, n18175);
  not g29053 (n_10894, n18176);
  not g29054 (n_10895, n18255);
  and g29055 (n18256, n_10894, n_10895);
  not g29056 (n_10896, n18254);
  and g29057 (n18257, n_10896, n18256);
  not g29058 (n_10897, n18257);
  and g29059 (n18258, n_10894, n_10897);
  not g29060 (n_10898, n18161);
  not g29061 (n_10899, n18258);
  and g29062 (n18259, n_10898, n_10899);
  not g29063 (n_10900, n18259);
  and g29064 (n18260, n_10813, n_10900);
  not g29065 (n_10901, n18144);
  and g29066 (n18261, n18132, n_10901);
  and g29067 (n18262, n_10801, n_10901);
  not g29068 (n_10902, n18261);
  not g29069 (n_10903, n18262);
  and g29070 (n18263, n_10902, n_10903);
  not g29071 (n_10904, n18260);
  not g29072 (n_10905, n18263);
  and g29073 (n18264, n_10904, n_10905);
  not g29074 (n_10906, n18264);
  and g29075 (n18265, n_10901, n_10906);
  not g29076 (n_10907, n18130);
  and g29077 (n18266, n18118, n_10907);
  and g29078 (n18267, n_10791, n_10907);
  not g29079 (n_10908, n18266);
  not g29080 (n_10909, n18267);
  and g29081 (n18268, n_10908, n_10909);
  not g29082 (n_10910, n18265);
  not g29083 (n_10911, n18268);
  and g29084 (n18269, n_10910, n_10911);
  not g29085 (n_10912, n18269);
  and g29086 (n18270, n_10907, n_10912);
  not g29087 (n_10913, n18104);
  and g29088 (n18271, n_10913, n18115);
  not g29089 (n_10914, n18116);
  not g29090 (n_10915, n18271);
  and g29091 (n18272, n_10914, n_10915);
  not g29092 (n_10916, n18270);
  and g29093 (n18273, n_10916, n18272);
  not g29094 (n_10917, n18273);
  and g29095 (n18274, n_10914, n_10917);
  not g29096 (n_10918, n18102);
  not g29097 (n_10919, n18274);
  and g29098 (n18275, n_10918, n_10919);
  not g29099 (n_10920, n18275);
  and g29100 (n18276, n_10768, n_10920);
  not g29101 (n_10921, n18084);
  not g29102 (n_10922, n18276);
  and g29103 (n18277, n_10921, n_10922);
  not g29104 (n_10923, n18277);
  and g29105 (n18278, n_10753, n_10923);
  not g29106 (n_10924, n18067);
  and g29107 (n18279, n18055, n_10924);
  and g29108 (n18280, n_10741, n_10924);
  not g29109 (n_10925, n18279);
  not g29110 (n_10926, n18280);
  and g29111 (n18281, n_10925, n_10926);
  not g29112 (n_10927, n18278);
  not g29113 (n_10928, n18281);
  and g29114 (n18282, n_10927, n_10928);
  not g29115 (n_10929, n18282);
  and g29116 (n18283, n_10924, n_10929);
  not g29117 (n_10930, n18053);
  and g29118 (n18284, n18041, n_10930);
  and g29119 (n18285, n_10731, n_10930);
  not g29120 (n_10931, n18284);
  not g29121 (n_10932, n18285);
  and g29122 (n18286, n_10931, n_10932);
  not g29123 (n_10933, n18283);
  not g29124 (n_10934, n18286);
  and g29125 (n18287, n_10933, n_10934);
  not g29126 (n_10935, n18287);
  and g29127 (n18288, n_10930, n_10935);
  not g29128 (n_10936, n18039);
  and g29129 (n18289, n18027, n_10936);
  and g29130 (n18290, n_10721, n_10936);
  not g29131 (n_10937, n18289);
  not g29132 (n_10938, n18290);
  and g29133 (n18291, n_10937, n_10938);
  not g29134 (n_10939, n18288);
  not g29135 (n_10940, n18291);
  and g29136 (n18292, n_10939, n_10940);
  not g29137 (n_10941, n18292);
  and g29138 (n18293, n_10936, n_10941);
  not g29139 (n_10942, n18025);
  and g29140 (n18294, n18013, n_10942);
  and g29141 (n18295, n_10711, n_10942);
  not g29142 (n_10943, n18294);
  not g29143 (n_10944, n18295);
  and g29144 (n18296, n_10943, n_10944);
  not g29145 (n_10945, n18293);
  not g29146 (n_10946, n18296);
  and g29147 (n18297, n_10945, n_10946);
  not g29148 (n_10947, n18297);
  and g29149 (n18298, n_10942, n_10947);
  not g29150 (n_10948, n18011);
  and g29151 (n18299, n17999, n_10948);
  and g29152 (n18300, n_10701, n_10948);
  not g29153 (n_10949, n18299);
  not g29154 (n_10950, n18300);
  and g29155 (n18301, n_10949, n_10950);
  not g29156 (n_10951, n18298);
  not g29157 (n_10952, n18301);
  and g29158 (n18302, n_10951, n_10952);
  not g29159 (n_10953, n18302);
  and g29160 (n18303, n_10948, n_10953);
  not g29161 (n_10954, n17997);
  and g29162 (n18304, n17985, n_10954);
  and g29163 (n18305, n_10691, n_10954);
  not g29164 (n_10955, n18304);
  not g29165 (n_10956, n18305);
  and g29166 (n18306, n_10955, n_10956);
  not g29167 (n_10957, n18303);
  not g29168 (n_10958, n18306);
  and g29169 (n18307, n_10957, n_10958);
  not g29170 (n_10959, n18307);
  and g29171 (n18308, n_10954, n_10959);
  not g29172 (n_10960, n17983);
  and g29173 (n18309, n17971, n_10960);
  and g29174 (n18310, n_10681, n_10960);
  not g29175 (n_10961, n18309);
  not g29176 (n_10962, n18310);
  and g29177 (n18311, n_10961, n_10962);
  not g29178 (n_10963, n18308);
  not g29179 (n_10964, n18311);
  and g29180 (n18312, n_10963, n_10964);
  not g29181 (n_10965, n18312);
  and g29182 (n18313, n_10960, n_10965);
  not g29183 (n_10966, n17969);
  and g29184 (n18314, n17957, n_10966);
  and g29185 (n18315, n_10670, n_10966);
  not g29186 (n_10967, n18314);
  not g29187 (n_10968, n18315);
  and g29188 (n18316, n_10967, n_10968);
  not g29189 (n_10969, n18313);
  not g29190 (n_10970, n18316);
  and g29191 (n18317, n_10969, n_10970);
  not g29192 (n_10971, n18317);
  and g29193 (n18318, n_10966, n_10971);
  not g29194 (n_10972, n17955);
  and g29195 (n18319, n17943, n_10972);
  and g29196 (n18320, n_10659, n_10972);
  not g29197 (n_10973, n18319);
  not g29198 (n_10974, n18320);
  and g29199 (n18321, n_10973, n_10974);
  not g29200 (n_10975, n18318);
  not g29201 (n_10976, n18321);
  and g29202 (n18322, n_10975, n_10976);
  not g29203 (n_10977, n18322);
  and g29204 (n18323, n_10972, n_10977);
  not g29205 (n_10978, n17929);
  and g29206 (n18324, n_10978, n17940);
  not g29207 (n_10979, n17941);
  not g29208 (n_10980, n18324);
  and g29209 (n18325, n_10979, n_10980);
  not g29210 (n_10981, n18323);
  and g29211 (n18326, n_10981, n18325);
  not g29212 (n_10982, n18326);
  and g29213 (n18327, n_10979, n_10982);
  not g29214 (n_10983, n17927);
  not g29215 (n_10984, n18327);
  and g29216 (n18328, n_10983, n_10984);
  and g29217 (n18329, n17927, n18327);
  not g29218 (n_10985, n18328);
  not g29219 (n_10986, n18329);
  and g29220 (n18330, n_10985, n_10986);
  and g29221 (n18331, n6233, n12370);
  and g29222 (n18332, n5663, n12508);
  and g29223 (n18333, n5939, n12505);
  and g29229 (n18336, n5666, n_7607);
  not g29232 (n_10991, n18337);
  and g29233 (n18338, \a[17] , n_10991);
  not g29234 (n_10992, n18338);
  and g29235 (n18339, \a[17] , n_10992);
  and g29236 (n18340, n_10991, n_10992);
  not g29237 (n_10993, n18339);
  not g29238 (n_10994, n18340);
  and g29239 (n18341, n_10993, n_10994);
  not g29240 (n_10995, n18341);
  and g29241 (n18342, n18330, n_10995);
  not g29242 (n_10996, n18342);
  and g29243 (n18343, n_10985, n_10996);
  not g29244 (n_10997, n17924);
  not g29245 (n_10998, n18343);
  and g29246 (n18344, n_10997, n_10998);
  and g29247 (n18345, n17924, n18343);
  not g29248 (n_10999, n18344);
  not g29249 (n_11000, n18345);
  and g29250 (n18346, n_10999, n_11000);
  and g29251 (n18347, n7101, n13491);
  and g29252 (n18348, n6402, n12769);
  and g29253 (n18349, n6951, n12889);
  and g29259 (n18352, n6397, n_7447);
  not g29262 (n_11005, n18353);
  and g29263 (n18354, \a[14] , n_11005);
  not g29264 (n_11006, n18354);
  and g29265 (n18355, \a[14] , n_11006);
  and g29266 (n18356, n_11005, n_11006);
  not g29267 (n_11007, n18355);
  not g29268 (n_11008, n18356);
  and g29269 (n18357, n_11007, n_11008);
  not g29270 (n_11009, n18357);
  and g29271 (n18358, n18346, n_11009);
  not g29272 (n_11010, n18358);
  and g29273 (n18359, n_10999, n_11010);
  not g29274 (n_11011, n17921);
  not g29275 (n_11012, n18359);
  and g29276 (n18360, n_11011, n_11012);
  and g29277 (n18361, n17921, n18359);
  not g29278 (n_11013, n18360);
  not g29279 (n_11014, n18361);
  and g29280 (n18362, n_11013, n_11014);
  and g29281 (n18363, n7983, n13597);
  and g29282 (n18364, n7291, n13521);
  and g29283 (n18365, n7632, n13515);
  and g29289 (n18368, n7294, n_7765);
  not g29292 (n_11019, n18369);
  and g29293 (n18370, \a[11] , n_11019);
  not g29294 (n_11020, n18370);
  and g29295 (n18371, \a[11] , n_11020);
  and g29296 (n18372, n_11019, n_11020);
  not g29297 (n_11021, n18371);
  not g29298 (n_11022, n18372);
  and g29299 (n18373, n_11021, n_11022);
  not g29300 (n_11023, n18373);
  and g29301 (n18374, n18362, n_11023);
  not g29302 (n_11024, n18374);
  and g29303 (n18375, n_11013, n_11024);
  not g29304 (n_11025, n17918);
  not g29305 (n_11026, n18375);
  and g29306 (n18376, n_11025, n_11026);
  not g29307 (n_11027, n18376);
  and g29308 (n18377, n_10631, n_11027);
  not g29309 (n_11028, n17901);
  not g29310 (n_11029, n18377);
  and g29311 (n18378, n_11028, n_11029);
  and g29312 (n18379, n17901, n18377);
  not g29313 (n_11030, n18378);
  not g29314 (n_11031, n18379);
  and g29315 (n18380, n_11030, n_11031);
  and g29316 (n18381, n9331, n_7417);
  and g29317 (n18382, n8418, n_7540);
  and g29318 (n18383, n8860, n13941);
  and g29324 (n18386, n8421, n14028);
  not g29327 (n_11036, n18387);
  and g29328 (n18388, \a[8] , n_11036);
  not g29329 (n_11037, n18388);
  and g29330 (n18389, \a[8] , n_11037);
  and g29331 (n18390, n_11036, n_11037);
  not g29332 (n_11038, n18389);
  not g29333 (n_11039, n18390);
  and g29334 (n18391, n_11038, n_11039);
  not g29335 (n_11040, n18391);
  and g29336 (n18392, n18380, n_11040);
  not g29337 (n_11041, n18392);
  and g29338 (n18393, n_11030, n_11041);
  not g29339 (n_11042, n17898);
  not g29340 (n_11043, n18393);
  and g29341 (n18394, n_11042, n_11043);
  and g29342 (n18395, n17898, n18393);
  not g29343 (n_11044, n18394);
  not g29344 (n_11045, n18395);
  and g29345 (n18396, n_11044, n_11045);
  and g29346 (n18397, n18380, n_11041);
  and g29347 (n18398, n_11040, n_11041);
  not g29348 (n_11046, n18397);
  not g29349 (n_11047, n18398);
  and g29350 (n18399, n_11046, n_11047);
  and g29351 (n18400, n18362, n_11024);
  and g29352 (n18401, n_11023, n_11024);
  not g29353 (n_11048, n18400);
  not g29354 (n_11049, n18401);
  and g29355 (n18402, n_11048, n_11049);
  and g29356 (n18403, n18346, n_11010);
  and g29357 (n18404, n_11009, n_11010);
  not g29358 (n_11050, n18403);
  not g29359 (n_11051, n18404);
  and g29360 (n18405, n_11050, n_11051);
  and g29361 (n18406, n18330, n_10996);
  and g29362 (n18407, n_10995, n_10996);
  not g29363 (n_11052, n18406);
  not g29364 (n_11053, n18407);
  and g29365 (n18408, n_11052, n_11053);
  and g29366 (n18409, n6233, n12505);
  and g29367 (n18410, n5663, n12513);
  and g29368 (n18411, n5939, n12508);
  and g29374 (n18414, n5666, n_7804);
  not g29377 (n_11058, n18415);
  and g29378 (n18416, \a[17] , n_11058);
  not g29379 (n_11059, n18416);
  and g29380 (n18417, n_11058, n_11059);
  and g29381 (n18418, \a[17] , n_11059);
  not g29382 (n_11060, n18417);
  not g29383 (n_11061, n18418);
  and g29384 (n18419, n_11060, n_11061);
  not g29385 (n_11062, n18325);
  and g29386 (n18420, n18323, n_11062);
  not g29387 (n_11063, n18420);
  and g29388 (n18421, n_10982, n_11063);
  not g29389 (n_11064, n18419);
  and g29390 (n18422, n_11064, n18421);
  not g29391 (n_11065, n18422);
  and g29392 (n18423, n_11064, n_11065);
  and g29393 (n18424, n18421, n_11065);
  not g29394 (n_11066, n18423);
  not g29395 (n_11067, n18424);
  and g29396 (n18425, n_11066, n_11067);
  and g29397 (n18426, n6233, n12508);
  and g29398 (n18427, n5663, n12511);
  and g29399 (n18428, n5939, n12513);
  and g29405 (n18431, n5666, n13863);
  not g29408 (n_11072, n18432);
  and g29409 (n18433, \a[17] , n_11072);
  not g29410 (n_11073, n18433);
  and g29411 (n18434, n_11072, n_11073);
  and g29412 (n18435, \a[17] , n_11073);
  not g29413 (n_11074, n18434);
  not g29414 (n_11075, n18435);
  and g29415 (n18436, n_11074, n_11075);
  and g29416 (n18437, n_10975, n_10977);
  and g29417 (n18438, n_10976, n_10977);
  not g29418 (n_11076, n18437);
  not g29419 (n_11077, n18438);
  and g29420 (n18439, n_11076, n_11077);
  not g29421 (n_11078, n18436);
  not g29422 (n_11079, n18439);
  and g29423 (n18440, n_11078, n_11079);
  not g29424 (n_11080, n18440);
  and g29425 (n18441, n_11078, n_11080);
  and g29426 (n18442, n_11079, n_11080);
  not g29427 (n_11081, n18441);
  not g29428 (n_11082, n18442);
  and g29429 (n18443, n_11081, n_11082);
  and g29430 (n18444, n6233, n12513);
  and g29431 (n18445, n5663, n12516);
  and g29432 (n18446, n5939, n12511);
  and g29438 (n18449, n5666, n14177);
  not g29441 (n_11087, n18450);
  and g29442 (n18451, \a[17] , n_11087);
  not g29443 (n_11088, n18451);
  and g29444 (n18452, n_11087, n_11088);
  and g29445 (n18453, \a[17] , n_11088);
  not g29446 (n_11089, n18452);
  not g29447 (n_11090, n18453);
  and g29448 (n18454, n_11089, n_11090);
  and g29449 (n18455, n_10969, n_10971);
  and g29450 (n18456, n_10970, n_10971);
  not g29451 (n_11091, n18455);
  not g29452 (n_11092, n18456);
  and g29453 (n18457, n_11091, n_11092);
  not g29454 (n_11093, n18454);
  not g29455 (n_11094, n18457);
  and g29456 (n18458, n_11093, n_11094);
  not g29457 (n_11095, n18458);
  and g29458 (n18459, n_11093, n_11095);
  and g29459 (n18460, n_11094, n_11095);
  not g29460 (n_11096, n18459);
  not g29461 (n_11097, n18460);
  and g29462 (n18461, n_11096, n_11097);
  and g29463 (n18462, n6233, n12511);
  and g29464 (n18463, n5663, n12519);
  and g29465 (n18464, n5939, n12516);
  and g29471 (n18467, n5666, n_7923);
  not g29474 (n_11102, n18468);
  and g29475 (n18469, \a[17] , n_11102);
  not g29476 (n_11103, n18469);
  and g29477 (n18470, n_11102, n_11103);
  and g29478 (n18471, \a[17] , n_11103);
  not g29479 (n_11104, n18470);
  not g29480 (n_11105, n18471);
  and g29481 (n18472, n_11104, n_11105);
  and g29482 (n18473, n_10963, n_10965);
  and g29483 (n18474, n_10964, n_10965);
  not g29484 (n_11106, n18473);
  not g29485 (n_11107, n18474);
  and g29486 (n18475, n_11106, n_11107);
  not g29487 (n_11108, n18472);
  not g29488 (n_11109, n18475);
  and g29489 (n18476, n_11108, n_11109);
  not g29490 (n_11110, n18476);
  and g29491 (n18477, n_11108, n_11110);
  and g29492 (n18478, n_11109, n_11110);
  not g29493 (n_11111, n18477);
  not g29494 (n_11112, n18478);
  and g29495 (n18479, n_11111, n_11112);
  and g29496 (n18480, n6233, n12516);
  and g29497 (n18481, n5663, n12522);
  and g29498 (n18482, n5939, n12519);
  and g29504 (n18485, n5666, n_8061);
  not g29507 (n_11117, n18486);
  and g29508 (n18487, \a[17] , n_11117);
  not g29509 (n_11118, n18487);
  and g29510 (n18488, n_11117, n_11118);
  and g29511 (n18489, \a[17] , n_11118);
  not g29512 (n_11119, n18488);
  not g29513 (n_11120, n18489);
  and g29514 (n18490, n_11119, n_11120);
  and g29515 (n18491, n_10957, n_10959);
  and g29516 (n18492, n_10958, n_10959);
  not g29517 (n_11121, n18491);
  not g29518 (n_11122, n18492);
  and g29519 (n18493, n_11121, n_11122);
  not g29520 (n_11123, n18490);
  not g29521 (n_11124, n18493);
  and g29522 (n18494, n_11123, n_11124);
  not g29523 (n_11125, n18494);
  and g29524 (n18495, n_11123, n_11125);
  and g29525 (n18496, n_11124, n_11125);
  not g29526 (n_11126, n18495);
  not g29527 (n_11127, n18496);
  and g29528 (n18497, n_11126, n_11127);
  and g29529 (n18498, n6233, n12519);
  and g29530 (n18499, n5663, n12525);
  and g29531 (n18500, n5939, n12522);
  and g29537 (n18503, n5666, n14454);
  not g29540 (n_11132, n18504);
  and g29541 (n18505, \a[17] , n_11132);
  not g29542 (n_11133, n18505);
  and g29543 (n18506, n_11132, n_11133);
  and g29544 (n18507, \a[17] , n_11133);
  not g29545 (n_11134, n18506);
  not g29546 (n_11135, n18507);
  and g29547 (n18508, n_11134, n_11135);
  and g29548 (n18509, n_10951, n_10953);
  and g29549 (n18510, n_10952, n_10953);
  not g29550 (n_11136, n18509);
  not g29551 (n_11137, n18510);
  and g29552 (n18511, n_11136, n_11137);
  not g29553 (n_11138, n18508);
  not g29554 (n_11139, n18511);
  and g29555 (n18512, n_11138, n_11139);
  not g29556 (n_11140, n18512);
  and g29557 (n18513, n_11138, n_11140);
  and g29558 (n18514, n_11139, n_11140);
  not g29559 (n_11141, n18513);
  not g29560 (n_11142, n18514);
  and g29561 (n18515, n_11141, n_11142);
  and g29562 (n18516, n6233, n12522);
  and g29563 (n18517, n5663, n12528);
  and g29564 (n18518, n5939, n12525);
  and g29570 (n18521, n5666, n14837);
  not g29573 (n_11147, n18522);
  and g29574 (n18523, \a[17] , n_11147);
  not g29575 (n_11148, n18523);
  and g29576 (n18524, n_11147, n_11148);
  and g29577 (n18525, \a[17] , n_11148);
  not g29578 (n_11149, n18524);
  not g29579 (n_11150, n18525);
  and g29580 (n18526, n_11149, n_11150);
  and g29581 (n18527, n_10945, n_10947);
  and g29582 (n18528, n_10946, n_10947);
  not g29583 (n_11151, n18527);
  not g29584 (n_11152, n18528);
  and g29585 (n18529, n_11151, n_11152);
  not g29586 (n_11153, n18526);
  not g29587 (n_11154, n18529);
  and g29588 (n18530, n_11153, n_11154);
  not g29589 (n_11155, n18530);
  and g29590 (n18531, n_11153, n_11155);
  and g29591 (n18532, n_11154, n_11155);
  not g29592 (n_11156, n18531);
  not g29593 (n_11157, n18532);
  and g29594 (n18533, n_11156, n_11157);
  and g29595 (n18534, n6233, n12525);
  and g29596 (n18535, n5663, n12531);
  and g29597 (n18536, n5939, n12528);
  and g29603 (n18539, n5666, n14608);
  not g29606 (n_11162, n18540);
  and g29607 (n18541, \a[17] , n_11162);
  not g29608 (n_11163, n18541);
  and g29609 (n18542, n_11162, n_11163);
  and g29610 (n18543, \a[17] , n_11163);
  not g29611 (n_11164, n18542);
  not g29612 (n_11165, n18543);
  and g29613 (n18544, n_11164, n_11165);
  and g29614 (n18545, n_10939, n_10941);
  and g29615 (n18546, n_10940, n_10941);
  not g29616 (n_11166, n18545);
  not g29617 (n_11167, n18546);
  and g29618 (n18547, n_11166, n_11167);
  not g29619 (n_11168, n18544);
  not g29620 (n_11169, n18547);
  and g29621 (n18548, n_11168, n_11169);
  not g29622 (n_11170, n18548);
  and g29623 (n18549, n_11168, n_11170);
  and g29624 (n18550, n_11169, n_11170);
  not g29625 (n_11171, n18549);
  not g29626 (n_11172, n18550);
  and g29627 (n18551, n_11171, n_11172);
  and g29628 (n18552, n6233, n12528);
  and g29629 (n18553, n5663, n12534);
  and g29630 (n18554, n5939, n12531);
  and g29636 (n18557, n5666, n_8448);
  not g29639 (n_11177, n18558);
  and g29640 (n18559, \a[17] , n_11177);
  not g29641 (n_11178, n18559);
  and g29642 (n18560, n_11177, n_11178);
  and g29643 (n18561, \a[17] , n_11178);
  not g29644 (n_11179, n18560);
  not g29645 (n_11180, n18561);
  and g29646 (n18562, n_11179, n_11180);
  and g29647 (n18563, n_10933, n_10935);
  and g29648 (n18564, n_10934, n_10935);
  not g29649 (n_11181, n18563);
  not g29650 (n_11182, n18564);
  and g29651 (n18565, n_11181, n_11182);
  not g29652 (n_11183, n18562);
  not g29653 (n_11184, n18565);
  and g29654 (n18566, n_11183, n_11184);
  not g29655 (n_11185, n18566);
  and g29656 (n18567, n_11183, n_11185);
  and g29657 (n18568, n_11184, n_11185);
  not g29658 (n_11186, n18567);
  not g29659 (n_11187, n18568);
  and g29660 (n18569, n_11186, n_11187);
  and g29661 (n18570, n6233, n12531);
  and g29662 (n18571, n5663, n12537);
  and g29663 (n18572, n5939, n12534);
  and g29669 (n18575, n5666, n15255);
  not g29672 (n_11192, n18576);
  and g29673 (n18577, \a[17] , n_11192);
  not g29674 (n_11193, n18577);
  and g29675 (n18578, n_11192, n_11193);
  and g29676 (n18579, \a[17] , n_11193);
  not g29677 (n_11194, n18578);
  not g29678 (n_11195, n18579);
  and g29679 (n18580, n_11194, n_11195);
  and g29680 (n18581, n_10927, n_10929);
  and g29681 (n18582, n_10928, n_10929);
  not g29682 (n_11196, n18581);
  not g29683 (n_11197, n18582);
  and g29684 (n18583, n_11196, n_11197);
  not g29685 (n_11198, n18580);
  not g29686 (n_11199, n18583);
  and g29687 (n18584, n_11198, n_11199);
  not g29688 (n_11200, n18584);
  and g29689 (n18585, n_11198, n_11200);
  and g29690 (n18586, n_11199, n_11200);
  not g29691 (n_11201, n18585);
  not g29692 (n_11202, n18586);
  and g29693 (n18587, n_11201, n_11202);
  and g29694 (n18588, n18084, n18276);
  not g29695 (n_11203, n18588);
  and g29696 (n18589, n_10923, n_11203);
  and g29697 (n18590, n6233, n12534);
  and g29698 (n18591, n5663, n12540);
  and g29699 (n18592, n5939, n12537);
  not g29700 (n_11204, n18591);
  not g29701 (n_11205, n18592);
  and g29702 (n18593, n_11204, n_11205);
  not g29703 (n_11206, n18590);
  and g29704 (n18594, n_11206, n18593);
  and g29705 (n18595, n_1409, n18594);
  and g29706 (n18596, n15096, n18594);
  not g29707 (n_11207, n18595);
  not g29708 (n_11208, n18596);
  and g29709 (n18597, n_11207, n_11208);
  not g29710 (n_11209, n18597);
  and g29711 (n18598, \a[17] , n_11209);
  and g29712 (n18599, n_617, n18597);
  not g29713 (n_11210, n18598);
  not g29714 (n_11211, n18599);
  and g29715 (n18600, n_11210, n_11211);
  not g29716 (n_11212, n18600);
  and g29717 (n18601, n18589, n_11212);
  and g29718 (n18602, n18102, n18274);
  not g29719 (n_11213, n18602);
  and g29720 (n18603, n_10920, n_11213);
  and g29721 (n18604, n6233, n12537);
  and g29722 (n18605, n5663, n12543);
  and g29723 (n18606, n5939, n12540);
  not g29724 (n_11214, n18605);
  not g29725 (n_11215, n18606);
  and g29726 (n18607, n_11214, n_11215);
  not g29727 (n_11216, n18604);
  and g29728 (n18608, n_11216, n18607);
  and g29729 (n18609, n_1409, n18608);
  and g29730 (n18610, n15385, n18608);
  not g29731 (n_11217, n18609);
  not g29732 (n_11218, n18610);
  and g29733 (n18611, n_11217, n_11218);
  not g29734 (n_11219, n18611);
  and g29735 (n18612, \a[17] , n_11219);
  and g29736 (n18613, n_617, n18611);
  not g29737 (n_11220, n18612);
  not g29738 (n_11221, n18613);
  and g29739 (n18614, n_11220, n_11221);
  not g29740 (n_11222, n18614);
  and g29741 (n18615, n18603, n_11222);
  and g29742 (n18616, n6233, n12540);
  and g29743 (n18617, n5663, n12546);
  and g29744 (n18618, n5939, n12543);
  and g29750 (n18621, n5666, n_8936);
  not g29753 (n_11227, n18622);
  and g29754 (n18623, \a[17] , n_11227);
  not g29755 (n_11228, n18623);
  and g29756 (n18624, n_11227, n_11228);
  and g29757 (n18625, \a[17] , n_11228);
  not g29758 (n_11229, n18624);
  not g29759 (n_11230, n18625);
  and g29760 (n18626, n_11229, n_11230);
  not g29761 (n_11231, n18272);
  and g29762 (n18627, n18270, n_11231);
  not g29763 (n_11232, n18627);
  and g29764 (n18628, n_10917, n_11232);
  not g29765 (n_11233, n18626);
  and g29766 (n18629, n_11233, n18628);
  not g29767 (n_11234, n18629);
  and g29768 (n18630, n_11233, n_11234);
  and g29769 (n18631, n18628, n_11234);
  not g29770 (n_11235, n18630);
  not g29771 (n_11236, n18631);
  and g29772 (n18632, n_11235, n_11236);
  and g29773 (n18633, n6233, n12543);
  and g29774 (n18634, n5663, n12549);
  and g29775 (n18635, n5939, n12546);
  and g29781 (n18638, n5666, n15724);
  not g29784 (n_11241, n18639);
  and g29785 (n18640, \a[17] , n_11241);
  not g29786 (n_11242, n18640);
  and g29787 (n18641, n_11241, n_11242);
  and g29788 (n18642, \a[17] , n_11242);
  not g29789 (n_11243, n18641);
  not g29790 (n_11244, n18642);
  and g29791 (n18643, n_11243, n_11244);
  and g29792 (n18644, n_10910, n_10912);
  and g29793 (n18645, n_10911, n_10912);
  not g29794 (n_11245, n18644);
  not g29795 (n_11246, n18645);
  and g29796 (n18646, n_11245, n_11246);
  not g29797 (n_11247, n18643);
  not g29798 (n_11248, n18646);
  and g29799 (n18647, n_11247, n_11248);
  not g29800 (n_11249, n18647);
  and g29801 (n18648, n_11247, n_11249);
  and g29802 (n18649, n_11248, n_11249);
  not g29803 (n_11250, n18648);
  not g29804 (n_11251, n18649);
  and g29805 (n18650, n_11250, n_11251);
  and g29806 (n18651, n6233, n12546);
  and g29807 (n18652, n5663, n12552);
  and g29808 (n18653, n5939, n12549);
  and g29814 (n18656, n5666, n_8634);
  not g29817 (n_11256, n18657);
  and g29818 (n18658, \a[17] , n_11256);
  not g29819 (n_11257, n18658);
  and g29820 (n18659, n_11256, n_11257);
  and g29821 (n18660, \a[17] , n_11257);
  not g29822 (n_11258, n18659);
  not g29823 (n_11259, n18660);
  and g29824 (n18661, n_11258, n_11259);
  and g29825 (n18662, n_10904, n_10906);
  and g29826 (n18663, n_10905, n_10906);
  not g29827 (n_11260, n18662);
  not g29828 (n_11261, n18663);
  and g29829 (n18664, n_11260, n_11261);
  not g29830 (n_11262, n18661);
  not g29831 (n_11263, n18664);
  and g29832 (n18665, n_11262, n_11263);
  not g29833 (n_11264, n18665);
  and g29834 (n18666, n_11262, n_11264);
  and g29835 (n18667, n_11263, n_11264);
  not g29836 (n_11265, n18666);
  not g29837 (n_11266, n18667);
  and g29838 (n18668, n_11265, n_11266);
  and g29839 (n18669, n18161, n18258);
  not g29840 (n_11267, n18669);
  and g29841 (n18670, n_10900, n_11267);
  and g29842 (n18671, n6233, n12549);
  and g29843 (n18672, n5663, n12555);
  and g29844 (n18673, n5939, n12552);
  not g29845 (n_11268, n18672);
  not g29846 (n_11269, n18673);
  and g29847 (n18674, n_11268, n_11269);
  not g29848 (n_11270, n18671);
  and g29849 (n18675, n_11270, n18674);
  and g29850 (n18676, n_1409, n18675);
  and g29851 (n18677, n_9580, n18675);
  not g29852 (n_11271, n18676);
  not g29853 (n_11272, n18677);
  and g29854 (n18678, n_11271, n_11272);
  not g29855 (n_11273, n18678);
  and g29856 (n18679, \a[17] , n_11273);
  and g29857 (n18680, n_617, n18678);
  not g29858 (n_11274, n18679);
  not g29859 (n_11275, n18680);
  and g29860 (n18681, n_11274, n_11275);
  not g29861 (n_11276, n18681);
  and g29862 (n18682, n18670, n_11276);
  not g29863 (n_11277, n18256);
  and g29864 (n18683, n18254, n_11277);
  not g29865 (n_11278, n18683);
  and g29866 (n18684, n_10897, n_11278);
  and g29867 (n18685, n6233, n12552);
  and g29868 (n18686, n5663, n12558);
  and g29869 (n18687, n5939, n12555);
  not g29870 (n_11279, n18686);
  not g29871 (n_11280, n18687);
  and g29872 (n18688, n_11279, n_11280);
  not g29873 (n_11281, n18685);
  and g29874 (n18689, n_11281, n18688);
  and g29875 (n18690, n_1409, n18689);
  and g29876 (n18691, n15791, n18689);
  not g29877 (n_11282, n18690);
  not g29878 (n_11283, n18691);
  and g29879 (n18692, n_11282, n_11283);
  not g29880 (n_11284, n18692);
  and g29881 (n18693, \a[17] , n_11284);
  and g29882 (n18694, n_617, n18692);
  not g29883 (n_11285, n18693);
  not g29884 (n_11286, n18694);
  and g29885 (n18695, n_11285, n_11286);
  not g29886 (n_11287, n18695);
  and g29887 (n18696, n18684, n_11287);
  and g29888 (n18697, n18193, n18252);
  not g29889 (n_11288, n18697);
  and g29890 (n18698, n_10893, n_11288);
  and g29891 (n18699, n6233, n12555);
  and g29892 (n18700, n5663, n12561);
  and g29893 (n18701, n5939, n12558);
  not g29894 (n_11289, n18700);
  not g29895 (n_11290, n18701);
  and g29896 (n18702, n_11289, n_11290);
  not g29897 (n_11291, n18699);
  and g29898 (n18703, n_11291, n18702);
  and g29899 (n18704, n_1409, n18703);
  and g29900 (n18705, n15816, n18703);
  not g29901 (n_11292, n18704);
  not g29902 (n_11293, n18705);
  and g29903 (n18706, n_11292, n_11293);
  not g29904 (n_11294, n18706);
  and g29905 (n18707, \a[17] , n_11294);
  and g29906 (n18708, n_617, n18706);
  not g29907 (n_11295, n18707);
  not g29908 (n_11296, n18708);
  and g29909 (n18709, n_11295, n_11296);
  not g29910 (n_11297, n18709);
  and g29911 (n18710, n18698, n_11297);
  and g29912 (n18711, n6233, n12558);
  and g29913 (n18712, n5663, n12564);
  and g29914 (n18713, n5939, n12561);
  and g29920 (n18716, n5666, n15847);
  not g29923 (n_11302, n18717);
  and g29924 (n18718, \a[17] , n_11302);
  not g29925 (n_11303, n18718);
  and g29926 (n18719, n_11302, n_11303);
  and g29927 (n18720, \a[17] , n_11303);
  not g29928 (n_11304, n18719);
  not g29929 (n_11305, n18720);
  and g29930 (n18721, n_11304, n_11305);
  not g29931 (n_11306, n18250);
  and g29932 (n18722, n18248, n_11306);
  not g29933 (n_11307, n18722);
  and g29934 (n18723, n_10890, n_11307);
  not g29935 (n_11308, n18721);
  and g29936 (n18724, n_11308, n18723);
  not g29937 (n_11309, n18724);
  and g29938 (n18725, n_11308, n_11309);
  and g29939 (n18726, n18723, n_11309);
  not g29940 (n_11310, n18725);
  not g29941 (n_11311, n18726);
  and g29942 (n18727, n_11310, n_11311);
  and g29943 (n18728, n_10883, n_10885);
  and g29944 (n18729, n_10884, n_10885);
  not g29945 (n_11312, n18728);
  not g29946 (n_11313, n18729);
  and g29947 (n18730, n_11312, n_11313);
  and g29948 (n18731, n6233, n12561);
  and g29949 (n18732, n5663, n12567);
  and g29950 (n18733, n5939, n12564);
  not g29951 (n_11314, n18732);
  not g29952 (n_11315, n18733);
  and g29953 (n18734, n_11314, n_11315);
  not g29954 (n_11316, n18731);
  and g29955 (n18735, n_11316, n18734);
  and g29956 (n18736, n_1409, n18735);
  and g29957 (n18737, n15905, n18735);
  not g29958 (n_11317, n18736);
  not g29959 (n_11318, n18737);
  and g29960 (n18738, n_11317, n_11318);
  not g29961 (n_11319, n18738);
  and g29962 (n18739, \a[17] , n_11319);
  and g29963 (n18740, n_617, n18738);
  not g29964 (n_11320, n18739);
  not g29965 (n_11321, n18740);
  and g29966 (n18741, n_11320, n_11321);
  not g29967 (n_11322, n18730);
  not g29968 (n_11323, n18741);
  and g29969 (n18742, n_11322, n_11323);
  and g29970 (n18743, n6233, n12564);
  and g29971 (n18744, n5663, n12571);
  and g29972 (n18745, n5939, n12567);
  and g29978 (n18748, n5666, n_9006);
  not g29981 (n_11328, n18749);
  and g29982 (n18750, \a[17] , n_11328);
  not g29983 (n_11329, n18750);
  and g29984 (n18751, n_11328, n_11329);
  and g29985 (n18752, \a[17] , n_11329);
  not g29986 (n_11330, n18751);
  not g29987 (n_11331, n18752);
  and g29988 (n18753, n_11330, n_11331);
  not g29989 (n_11332, n18219);
  and g29990 (n18754, n_11332, n18230);
  not g29991 (n_11333, n18231);
  not g29992 (n_11334, n18754);
  and g29993 (n18755, n_11333, n_11334);
  not g29994 (n_11335, n18753);
  and g29995 (n18756, n_11335, n18755);
  not g29996 (n_11336, n18756);
  and g29997 (n18757, n_11335, n_11336);
  and g29998 (n18758, n18755, n_11336);
  not g29999 (n_11337, n18757);
  not g30000 (n_11338, n18758);
  and g30001 (n18759, n_11337, n_11338);
  not g30002 (n_11339, n18218);
  and g30003 (n18760, n18216, n_11339);
  not g30004 (n_11340, n18760);
  and g30005 (n18761, n_11332, n_11340);
  and g30006 (n18762, n6233, n12567);
  and g30007 (n18763, n5663, n12574);
  and g30008 (n18764, n5939, n12571);
  not g30009 (n_11341, n18763);
  not g30010 (n_11342, n18764);
  and g30011 (n18765, n_11341, n_11342);
  not g30012 (n_11343, n18762);
  and g30013 (n18766, n_11343, n18765);
  and g30014 (n18767, n_1409, n18766);
  and g30015 (n18768, n_10006, n18766);
  not g30016 (n_11344, n18767);
  not g30017 (n_11345, n18768);
  and g30018 (n18769, n_11344, n_11345);
  not g30019 (n_11346, n18769);
  and g30020 (n18770, \a[17] , n_11346);
  and g30021 (n18771, n_617, n18769);
  not g30022 (n_11347, n18770);
  not g30023 (n_11348, n18771);
  and g30024 (n18772, n_11347, n_11348);
  not g30025 (n_11349, n18772);
  and g30026 (n18773, n18761, n_11349);
  and g30027 (n18774, n5939, n_6977);
  and g30028 (n18775, n6233, n12577);
  not g30029 (n_11350, n18774);
  not g30030 (n_11351, n18775);
  and g30031 (n18776, n_11350, n_11351);
  and g30032 (n18777, n5666, n_9032);
  not g30033 (n_11352, n18777);
  and g30034 (n18778, n18776, n_11352);
  not g30035 (n_11353, n18778);
  and g30036 (n18779, \a[17] , n_11353);
  not g30037 (n_11354, n18779);
  and g30038 (n18780, \a[17] , n_11354);
  and g30039 (n18781, n_11353, n_11354);
  not g30040 (n_11355, n18780);
  not g30041 (n_11356, n18781);
  and g30042 (n18782, n_11355, n_11356);
  and g30043 (n18783, n_1408, n_6977);
  not g30044 (n_11357, n18783);
  and g30045 (n18784, \a[17] , n_11357);
  not g30046 (n_11358, n18782);
  and g30047 (n18785, n_11358, n18784);
  and g30048 (n18786, n6233, n12574);
  and g30049 (n18787, n5663, n_6977);
  and g30050 (n18788, n5939, n12577);
  not g30051 (n_11359, n18787);
  not g30052 (n_11360, n18788);
  and g30053 (n18789, n_11359, n_11360);
  not g30054 (n_11361, n18786);
  and g30055 (n18790, n_11361, n18789);
  and g30056 (n18791, n_1409, n18790);
  and g30057 (n18792, n16094, n18790);
  not g30058 (n_11362, n18791);
  not g30059 (n_11363, n18792);
  and g30060 (n18793, n_11362, n_11363);
  not g30061 (n_11364, n18793);
  and g30062 (n18794, \a[17] , n_11364);
  and g30063 (n18795, n_617, n18793);
  not g30064 (n_11365, n18794);
  not g30065 (n_11366, n18795);
  and g30066 (n18796, n_11365, n_11366);
  not g30067 (n_11367, n18796);
  and g30068 (n18797, n18785, n_11367);
  and g30069 (n18798, n18217, n18797);
  not g30070 (n_11368, n18798);
  and g30071 (n18799, n18797, n_11368);
  and g30072 (n18800, n18217, n_11368);
  not g30073 (n_11369, n18799);
  not g30074 (n_11370, n18800);
  and g30075 (n18801, n_11369, n_11370);
  and g30076 (n18802, n6233, n12571);
  and g30077 (n18803, n5663, n12577);
  and g30078 (n18804, n5939, n12574);
  and g30084 (n18807, n5666, n16013);
  not g30087 (n_11375, n18808);
  and g30088 (n18809, \a[17] , n_11375);
  not g30089 (n_11376, n18809);
  and g30090 (n18810, \a[17] , n_11376);
  and g30091 (n18811, n_11375, n_11376);
  not g30092 (n_11377, n18810);
  not g30093 (n_11378, n18811);
  and g30094 (n18812, n_11377, n_11378);
  not g30095 (n_11379, n18801);
  not g30096 (n_11380, n18812);
  and g30097 (n18813, n_11379, n_11380);
  not g30098 (n_11381, n18813);
  and g30099 (n18814, n_11368, n_11381);
  not g30100 (n_11382, n18761);
  and g30101 (n18815, n_11382, n18772);
  not g30102 (n_11383, n18773);
  not g30103 (n_11384, n18815);
  and g30104 (n18816, n_11383, n_11384);
  not g30105 (n_11385, n18814);
  and g30106 (n18817, n_11385, n18816);
  not g30107 (n_11386, n18817);
  and g30108 (n18818, n_11383, n_11386);
  not g30109 (n_11387, n18759);
  not g30110 (n_11388, n18818);
  and g30111 (n18819, n_11387, n_11388);
  not g30112 (n_11389, n18819);
  and g30113 (n18820, n_11336, n_11389);
  and g30114 (n18821, n18730, n18741);
  not g30115 (n_11390, n18742);
  not g30116 (n_11391, n18821);
  and g30117 (n18822, n_11390, n_11391);
  not g30118 (n_11392, n18820);
  and g30119 (n18823, n_11392, n18822);
  not g30120 (n_11393, n18823);
  and g30121 (n18824, n_11390, n_11393);
  not g30122 (n_11394, n18727);
  not g30123 (n_11395, n18824);
  and g30124 (n18825, n_11394, n_11395);
  not g30125 (n_11396, n18825);
  and g30126 (n18826, n_11309, n_11396);
  not g30127 (n_11397, n18710);
  and g30128 (n18827, n18698, n_11397);
  and g30129 (n18828, n_11297, n_11397);
  not g30130 (n_11398, n18827);
  not g30131 (n_11399, n18828);
  and g30132 (n18829, n_11398, n_11399);
  not g30133 (n_11400, n18826);
  not g30134 (n_11401, n18829);
  and g30135 (n18830, n_11400, n_11401);
  not g30136 (n_11402, n18830);
  and g30137 (n18831, n_11397, n_11402);
  not g30138 (n_11403, n18696);
  and g30139 (n18832, n18684, n_11403);
  and g30140 (n18833, n_11287, n_11403);
  not g30141 (n_11404, n18832);
  not g30142 (n_11405, n18833);
  and g30143 (n18834, n_11404, n_11405);
  not g30144 (n_11406, n18831);
  not g30145 (n_11407, n18834);
  and g30146 (n18835, n_11406, n_11407);
  not g30147 (n_11408, n18835);
  and g30148 (n18836, n_11403, n_11408);
  not g30149 (n_11409, n18670);
  and g30150 (n18837, n_11409, n18681);
  not g30151 (n_11410, n18682);
  not g30152 (n_11411, n18837);
  and g30153 (n18838, n_11410, n_11411);
  not g30154 (n_11412, n18836);
  and g30155 (n18839, n_11412, n18838);
  not g30156 (n_11413, n18839);
  and g30157 (n18840, n_11410, n_11413);
  not g30158 (n_11414, n18668);
  not g30159 (n_11415, n18840);
  and g30160 (n18841, n_11414, n_11415);
  not g30161 (n_11416, n18841);
  and g30162 (n18842, n_11264, n_11416);
  not g30163 (n_11417, n18650);
  not g30164 (n_11418, n18842);
  and g30165 (n18843, n_11417, n_11418);
  not g30166 (n_11419, n18843);
  and g30167 (n18844, n_11249, n_11419);
  not g30168 (n_11420, n18632);
  not g30169 (n_11421, n18844);
  and g30170 (n18845, n_11420, n_11421);
  not g30171 (n_11422, n18845);
  and g30172 (n18846, n_11234, n_11422);
  not g30173 (n_11423, n18615);
  and g30174 (n18847, n18603, n_11423);
  and g30175 (n18848, n_11222, n_11423);
  not g30176 (n_11424, n18847);
  not g30177 (n_11425, n18848);
  and g30178 (n18849, n_11424, n_11425);
  not g30179 (n_11426, n18846);
  not g30180 (n_11427, n18849);
  and g30181 (n18850, n_11426, n_11427);
  not g30182 (n_11428, n18850);
  and g30183 (n18851, n_11423, n_11428);
  not g30184 (n_11429, n18589);
  and g30185 (n18852, n_11429, n18600);
  not g30186 (n_11430, n18601);
  not g30187 (n_11431, n18852);
  and g30188 (n18853, n_11430, n_11431);
  not g30189 (n_11432, n18851);
  and g30190 (n18854, n_11432, n18853);
  not g30191 (n_11433, n18854);
  and g30192 (n18855, n_11430, n_11433);
  not g30193 (n_11434, n18587);
  not g30194 (n_11435, n18855);
  and g30195 (n18856, n_11434, n_11435);
  not g30196 (n_11436, n18856);
  and g30197 (n18857, n_11200, n_11436);
  not g30198 (n_11437, n18569);
  not g30199 (n_11438, n18857);
  and g30200 (n18858, n_11437, n_11438);
  not g30201 (n_11439, n18858);
  and g30202 (n18859, n_11185, n_11439);
  not g30203 (n_11440, n18551);
  not g30204 (n_11441, n18859);
  and g30205 (n18860, n_11440, n_11441);
  not g30206 (n_11442, n18860);
  and g30207 (n18861, n_11170, n_11442);
  not g30208 (n_11443, n18533);
  not g30209 (n_11444, n18861);
  and g30210 (n18862, n_11443, n_11444);
  not g30211 (n_11445, n18862);
  and g30212 (n18863, n_11155, n_11445);
  not g30213 (n_11446, n18515);
  not g30214 (n_11447, n18863);
  and g30215 (n18864, n_11446, n_11447);
  not g30216 (n_11448, n18864);
  and g30217 (n18865, n_11140, n_11448);
  not g30218 (n_11449, n18497);
  not g30219 (n_11450, n18865);
  and g30220 (n18866, n_11449, n_11450);
  not g30221 (n_11451, n18866);
  and g30222 (n18867, n_11125, n_11451);
  not g30223 (n_11452, n18479);
  not g30224 (n_11453, n18867);
  and g30225 (n18868, n_11452, n_11453);
  not g30226 (n_11454, n18868);
  and g30227 (n18869, n_11110, n_11454);
  not g30228 (n_11455, n18461);
  not g30229 (n_11456, n18869);
  and g30230 (n18870, n_11455, n_11456);
  not g30231 (n_11457, n18870);
  and g30232 (n18871, n_11095, n_11457);
  not g30233 (n_11458, n18443);
  not g30234 (n_11459, n18871);
  and g30235 (n18872, n_11458, n_11459);
  not g30236 (n_11460, n18872);
  and g30237 (n18873, n_11080, n_11460);
  not g30238 (n_11461, n18425);
  not g30239 (n_11462, n18873);
  and g30240 (n18874, n_11461, n_11462);
  not g30241 (n_11463, n18874);
  and g30242 (n18875, n_11065, n_11463);
  not g30243 (n_11464, n18408);
  not g30244 (n_11465, n18875);
  and g30245 (n18876, n_11464, n_11465);
  and g30246 (n18877, n18408, n18875);
  not g30247 (n_11466, n18876);
  not g30248 (n_11467, n18877);
  and g30249 (n18878, n_11466, n_11467);
  and g30250 (n18879, n7101, n12889);
  and g30251 (n18880, n6402, n12502);
  and g30252 (n18881, n6951, n12769);
  and g30258 (n18884, n6397, n12895);
  not g30261 (n_11472, n18885);
  and g30262 (n18886, \a[14] , n_11472);
  not g30263 (n_11473, n18886);
  and g30264 (n18887, \a[14] , n_11473);
  and g30265 (n18888, n_11472, n_11473);
  not g30266 (n_11474, n18887);
  not g30267 (n_11475, n18888);
  and g30268 (n18889, n_11474, n_11475);
  not g30269 (n_11476, n18889);
  and g30270 (n18890, n18878, n_11476);
  not g30271 (n_11477, n18890);
  and g30272 (n18891, n_11466, n_11477);
  not g30273 (n_11478, n18405);
  not g30274 (n_11479, n18891);
  and g30275 (n18892, n_11478, n_11479);
  and g30276 (n18893, n18405, n18891);
  not g30277 (n_11480, n18892);
  not g30278 (n_11481, n18893);
  and g30279 (n18894, n_11480, n_11481);
  and g30280 (n18895, n7983, n13515);
  and g30281 (n18896, n7291, n13518);
  and g30282 (n18897, n7632, n13521);
  and g30288 (n18900, n7294, n13541);
  not g30291 (n_11486, n18901);
  and g30292 (n18902, \a[11] , n_11486);
  not g30293 (n_11487, n18902);
  and g30294 (n18903, \a[11] , n_11487);
  and g30295 (n18904, n_11486, n_11487);
  not g30296 (n_11488, n18903);
  not g30297 (n_11489, n18904);
  and g30298 (n18905, n_11488, n_11489);
  not g30299 (n_11490, n18905);
  and g30300 (n18906, n18894, n_11490);
  not g30301 (n_11491, n18906);
  and g30302 (n18907, n_11480, n_11491);
  not g30303 (n_11492, n18402);
  not g30304 (n_11493, n18907);
  and g30305 (n18908, n_11492, n_11493);
  and g30306 (n18909, n18402, n18907);
  not g30307 (n_11494, n18908);
  not g30308 (n_11495, n18909);
  and g30309 (n18910, n_11494, n_11495);
  and g30310 (n18911, n9331, n_7540);
  and g30311 (n18912, n8418, n13630);
  and g30312 (n18913, n8860, n13633);
  and g30318 (n18916, n8421, n_7563);
  not g30321 (n_11500, n18917);
  and g30322 (n18918, \a[8] , n_11500);
  not g30323 (n_11501, n18918);
  and g30324 (n18919, \a[8] , n_11501);
  and g30325 (n18920, n_11500, n_11501);
  not g30326 (n_11502, n18919);
  not g30327 (n_11503, n18920);
  and g30328 (n18921, n_11502, n_11503);
  not g30329 (n_11504, n18921);
  and g30330 (n18922, n18910, n_11504);
  not g30331 (n_11505, n18922);
  and g30332 (n18923, n_11494, n_11505);
  and g30333 (n18924, n9331, n13941);
  and g30334 (n18925, n8418, n13633);
  and g30335 (n18926, n8860, n_7540);
  and g30341 (n18929, n8421, n14136);
  not g30344 (n_11510, n18930);
  and g30345 (n18931, \a[8] , n_11510);
  not g30346 (n_11511, n18931);
  and g30347 (n18932, \a[8] , n_11511);
  and g30348 (n18933, n_11510, n_11511);
  not g30349 (n_11512, n18932);
  not g30350 (n_11513, n18933);
  and g30351 (n18934, n_11512, n_11513);
  not g30352 (n_11514, n18923);
  not g30353 (n_11515, n18934);
  and g30354 (n18935, n_11514, n_11515);
  not g30355 (n_11516, n18935);
  and g30356 (n18936, n_11514, n_11516);
  and g30357 (n18937, n_11515, n_11516);
  not g30358 (n_11517, n18936);
  not g30359 (n_11518, n18937);
  and g30360 (n18938, n_11517, n_11518);
  and g30361 (n18939, n17918, n18375);
  not g30362 (n_11519, n18939);
  and g30363 (n18940, n_11027, n_11519);
  not g30364 (n_11520, n18938);
  and g30365 (n18941, n_11520, n18940);
  not g30366 (n_11521, n18941);
  and g30367 (n18942, n_11516, n_11521);
  not g30368 (n_11522, n18399);
  not g30369 (n_11523, n18942);
  and g30370 (n18943, n_11522, n_11523);
  not g30371 (n_11524, n18943);
  and g30372 (n18944, n_11522, n_11524);
  and g30373 (n18945, n_11523, n_11524);
  not g30374 (n_11525, n18944);
  not g30375 (n_11526, n18945);
  and g30376 (n18946, n_11525, n_11526);
  and g30377 (n18947, n18894, n_11491);
  and g30378 (n18948, n_11490, n_11491);
  not g30379 (n_11527, n18947);
  not g30380 (n_11528, n18948);
  and g30381 (n18949, n_11527, n_11528);
  and g30382 (n18950, n18878, n_11477);
  and g30383 (n18951, n_11476, n_11477);
  not g30384 (n_11529, n18950);
  not g30385 (n_11530, n18951);
  and g30386 (n18952, n_11529, n_11530);
  and g30387 (n18953, n18425, n18873);
  not g30388 (n_11531, n18953);
  and g30389 (n18954, n_11463, n_11531);
  and g30390 (n18955, n7101, n12769);
  and g30391 (n18956, n6402, n12370);
  and g30392 (n18957, n6951, n12502);
  not g30393 (n_11532, n18956);
  not g30394 (n_11533, n18957);
  and g30395 (n18958, n_11532, n_11533);
  not g30396 (n_11534, n18955);
  and g30397 (n18959, n_11534, n18958);
  and g30398 (n18960, n_1885, n18959);
  and g30399 (n18961, n_7817, n18959);
  not g30400 (n_11535, n18960);
  not g30401 (n_11536, n18961);
  and g30402 (n18962, n_11535, n_11536);
  not g30403 (n_11537, n18962);
  and g30404 (n18963, \a[14] , n_11537);
  and g30405 (n18964, n_652, n18962);
  not g30406 (n_11538, n18963);
  not g30407 (n_11539, n18964);
  and g30408 (n18965, n_11538, n_11539);
  not g30409 (n_11540, n18965);
  and g30410 (n18966, n18954, n_11540);
  and g30411 (n18967, n18443, n18871);
  not g30412 (n_11541, n18967);
  and g30413 (n18968, n_11460, n_11541);
  and g30414 (n18969, n7101, n12502);
  and g30415 (n18970, n6402, n12505);
  and g30416 (n18971, n6951, n12370);
  not g30417 (n_11542, n18970);
  not g30418 (n_11543, n18971);
  and g30419 (n18972, n_11542, n_11543);
  not g30420 (n_11544, n18969);
  and g30421 (n18973, n_11544, n18972);
  and g30422 (n18974, n_1885, n18973);
  and g30423 (n18975, n13736, n18973);
  not g30424 (n_11545, n18974);
  not g30425 (n_11546, n18975);
  and g30426 (n18976, n_11545, n_11546);
  not g30427 (n_11547, n18976);
  and g30428 (n18977, \a[14] , n_11547);
  and g30429 (n18978, n_652, n18976);
  not g30430 (n_11548, n18977);
  not g30431 (n_11549, n18978);
  and g30432 (n18979, n_11548, n_11549);
  not g30433 (n_11550, n18979);
  and g30434 (n18980, n18968, n_11550);
  and g30435 (n18981, n18461, n18869);
  not g30436 (n_11551, n18981);
  and g30437 (n18982, n_11457, n_11551);
  and g30438 (n18983, n7101, n12370);
  and g30439 (n18984, n6402, n12508);
  and g30440 (n18985, n6951, n12505);
  not g30441 (n_11552, n18984);
  not g30442 (n_11553, n18985);
  and g30443 (n18986, n_11552, n_11553);
  not g30444 (n_11554, n18983);
  and g30445 (n18987, n_11554, n18986);
  and g30446 (n18988, n_1885, n18987);
  and g30447 (n18989, n13748, n18987);
  not g30448 (n_11555, n18988);
  not g30449 (n_11556, n18989);
  and g30450 (n18990, n_11555, n_11556);
  not g30451 (n_11557, n18990);
  and g30452 (n18991, \a[14] , n_11557);
  and g30453 (n18992, n_652, n18990);
  not g30454 (n_11558, n18991);
  not g30455 (n_11559, n18992);
  and g30456 (n18993, n_11558, n_11559);
  not g30457 (n_11560, n18993);
  and g30458 (n18994, n18982, n_11560);
  and g30459 (n18995, n18479, n18867);
  not g30460 (n_11561, n18995);
  and g30461 (n18996, n_11454, n_11561);
  and g30462 (n18997, n7101, n12505);
  and g30463 (n18998, n6402, n12513);
  and g30464 (n18999, n6951, n12508);
  not g30465 (n_11562, n18998);
  not g30466 (n_11563, n18999);
  and g30467 (n19000, n_11562, n_11563);
  not g30468 (n_11564, n18997);
  and g30469 (n19001, n_11564, n19000);
  and g30470 (n19002, n_1885, n19001);
  and g30471 (n19003, n14051, n19001);
  not g30472 (n_11565, n19002);
  not g30473 (n_11566, n19003);
  and g30474 (n19004, n_11565, n_11566);
  not g30475 (n_11567, n19004);
  and g30476 (n19005, \a[14] , n_11567);
  and g30477 (n19006, n_652, n19004);
  not g30478 (n_11568, n19005);
  not g30479 (n_11569, n19006);
  and g30480 (n19007, n_11568, n_11569);
  not g30481 (n_11570, n19007);
  and g30482 (n19008, n18996, n_11570);
  and g30483 (n19009, n18497, n18865);
  not g30484 (n_11571, n19009);
  and g30485 (n19010, n_11451, n_11571);
  and g30486 (n19011, n7101, n12508);
  and g30487 (n19012, n6402, n12511);
  and g30488 (n19013, n6951, n12513);
  not g30489 (n_11572, n19012);
  not g30490 (n_11573, n19013);
  and g30491 (n19014, n_11572, n_11573);
  not g30492 (n_11574, n19011);
  and g30493 (n19015, n_11574, n19014);
  and g30494 (n19016, n_1885, n19015);
  and g30495 (n19017, n_8125, n19015);
  not g30496 (n_11575, n19016);
  not g30497 (n_11576, n19017);
  and g30498 (n19018, n_11575, n_11576);
  not g30499 (n_11577, n19018);
  and g30500 (n19019, \a[14] , n_11577);
  and g30501 (n19020, n_652, n19018);
  not g30502 (n_11578, n19019);
  not g30503 (n_11579, n19020);
  and g30504 (n19021, n_11578, n_11579);
  not g30505 (n_11580, n19021);
  and g30506 (n19022, n19010, n_11580);
  and g30507 (n19023, n18515, n18863);
  not g30508 (n_11581, n19023);
  and g30509 (n19024, n_11448, n_11581);
  and g30510 (n19025, n7101, n12513);
  and g30511 (n19026, n6402, n12516);
  and g30512 (n19027, n6951, n12511);
  not g30513 (n_11582, n19026);
  not g30514 (n_11583, n19027);
  and g30515 (n19028, n_11582, n_11583);
  not g30516 (n_11584, n19025);
  and g30517 (n19029, n_11584, n19028);
  and g30518 (n19030, n_1885, n19029);
  not g30519 (n_11585, n14177);
  and g30520 (n19031, n_11585, n19029);
  not g30521 (n_11586, n19030);
  not g30522 (n_11587, n19031);
  and g30523 (n19032, n_11586, n_11587);
  not g30524 (n_11588, n19032);
  and g30525 (n19033, \a[14] , n_11588);
  and g30526 (n19034, n_652, n19032);
  not g30527 (n_11589, n19033);
  not g30528 (n_11590, n19034);
  and g30529 (n19035, n_11589, n_11590);
  not g30530 (n_11591, n19035);
  and g30531 (n19036, n19024, n_11591);
  and g30532 (n19037, n18533, n18861);
  not g30533 (n_11592, n19037);
  and g30534 (n19038, n_11445, n_11592);
  and g30535 (n19039, n7101, n12511);
  and g30536 (n19040, n6402, n12519);
  and g30537 (n19041, n6951, n12516);
  not g30538 (n_11593, n19040);
  not g30539 (n_11594, n19041);
  and g30540 (n19042, n_11593, n_11594);
  not g30541 (n_11595, n19039);
  and g30542 (n19043, n_11595, n19042);
  and g30543 (n19044, n_1885, n19043);
  and g30544 (n19045, n14233, n19043);
  not g30545 (n_11596, n19044);
  not g30546 (n_11597, n19045);
  and g30547 (n19046, n_11596, n_11597);
  not g30548 (n_11598, n19046);
  and g30549 (n19047, \a[14] , n_11598);
  and g30550 (n19048, n_652, n19046);
  not g30551 (n_11599, n19047);
  not g30552 (n_11600, n19048);
  and g30553 (n19049, n_11599, n_11600);
  not g30554 (n_11601, n19049);
  and g30555 (n19050, n19038, n_11601);
  and g30556 (n19051, n18551, n18859);
  not g30557 (n_11602, n19051);
  and g30558 (n19052, n_11442, n_11602);
  and g30559 (n19053, n7101, n12516);
  and g30560 (n19054, n6402, n12522);
  and g30561 (n19055, n6951, n12519);
  not g30562 (n_11603, n19054);
  not g30563 (n_11604, n19055);
  and g30564 (n19056, n_11603, n_11604);
  not g30565 (n_11605, n19053);
  and g30566 (n19057, n_11605, n19056);
  and g30567 (n19058, n_1885, n19057);
  and g30568 (n19059, n14443, n19057);
  not g30569 (n_11606, n19058);
  not g30570 (n_11607, n19059);
  and g30571 (n19060, n_11606, n_11607);
  not g30572 (n_11608, n19060);
  and g30573 (n19061, \a[14] , n_11608);
  and g30574 (n19062, n_652, n19060);
  not g30575 (n_11609, n19061);
  not g30576 (n_11610, n19062);
  and g30577 (n19063, n_11609, n_11610);
  not g30578 (n_11611, n19063);
  and g30579 (n19064, n19052, n_11611);
  and g30580 (n19065, n18569, n18857);
  not g30581 (n_11612, n19065);
  and g30582 (n19066, n_11439, n_11612);
  and g30583 (n19067, n7101, n12519);
  and g30584 (n19068, n6402, n12525);
  and g30585 (n19069, n6951, n12522);
  not g30586 (n_11613, n19068);
  not g30587 (n_11614, n19069);
  and g30588 (n19070, n_11613, n_11614);
  not g30589 (n_11615, n19067);
  and g30590 (n19071, n_11615, n19070);
  and g30591 (n19072, n_1885, n19071);
  and g30592 (n19073, n_10664, n19071);
  not g30593 (n_11616, n19072);
  not g30594 (n_11617, n19073);
  and g30595 (n19074, n_11616, n_11617);
  not g30596 (n_11618, n19074);
  and g30597 (n19075, \a[14] , n_11618);
  and g30598 (n19076, n_652, n19074);
  not g30599 (n_11619, n19075);
  not g30600 (n_11620, n19076);
  and g30601 (n19077, n_11619, n_11620);
  not g30602 (n_11621, n19077);
  and g30603 (n19078, n19066, n_11621);
  and g30604 (n19079, n18587, n18855);
  not g30605 (n_11622, n19079);
  and g30606 (n19080, n_11436, n_11622);
  and g30607 (n19081, n7101, n12522);
  and g30608 (n19082, n6402, n12528);
  and g30609 (n19083, n6951, n12525);
  not g30610 (n_11623, n19082);
  not g30611 (n_11624, n19083);
  and g30612 (n19084, n_11623, n_11624);
  not g30613 (n_11625, n19081);
  and g30614 (n19085, n_11625, n19084);
  and g30615 (n19086, n_1885, n19085);
  and g30616 (n19087, n_10675, n19085);
  not g30617 (n_11626, n19086);
  not g30618 (n_11627, n19087);
  and g30619 (n19088, n_11626, n_11627);
  not g30620 (n_11628, n19088);
  and g30621 (n19089, \a[14] , n_11628);
  and g30622 (n19090, n_652, n19088);
  not g30623 (n_11629, n19089);
  not g30624 (n_11630, n19090);
  and g30625 (n19091, n_11629, n_11630);
  not g30626 (n_11631, n19091);
  and g30627 (n19092, n19080, n_11631);
  and g30628 (n19093, n7101, n12525);
  and g30629 (n19094, n6402, n12531);
  and g30630 (n19095, n6951, n12528);
  and g30636 (n19098, n6397, n14608);
  not g30639 (n_11636, n19099);
  and g30640 (n19100, \a[14] , n_11636);
  not g30641 (n_11637, n19100);
  and g30642 (n19101, n_11636, n_11637);
  and g30643 (n19102, \a[14] , n_11637);
  not g30644 (n_11638, n19101);
  not g30645 (n_11639, n19102);
  and g30646 (n19103, n_11638, n_11639);
  not g30647 (n_11640, n18853);
  and g30648 (n19104, n18851, n_11640);
  not g30649 (n_11641, n19104);
  and g30650 (n19105, n_11433, n_11641);
  not g30651 (n_11642, n19103);
  and g30652 (n19106, n_11642, n19105);
  not g30653 (n_11643, n19106);
  and g30654 (n19107, n_11642, n_11643);
  and g30655 (n19108, n19105, n_11643);
  not g30656 (n_11644, n19107);
  not g30657 (n_11645, n19108);
  and g30658 (n19109, n_11644, n_11645);
  and g30659 (n19110, n7101, n12528);
  and g30660 (n19111, n6402, n12534);
  and g30661 (n19112, n6951, n12531);
  and g30667 (n19115, n6397, n_8448);
  not g30670 (n_11650, n19116);
  and g30671 (n19117, \a[14] , n_11650);
  not g30672 (n_11651, n19117);
  and g30673 (n19118, n_11650, n_11651);
  and g30674 (n19119, \a[14] , n_11651);
  not g30675 (n_11652, n19118);
  not g30676 (n_11653, n19119);
  and g30677 (n19120, n_11652, n_11653);
  and g30678 (n19121, n_11426, n_11428);
  and g30679 (n19122, n_11427, n_11428);
  not g30680 (n_11654, n19121);
  not g30681 (n_11655, n19122);
  and g30682 (n19123, n_11654, n_11655);
  not g30683 (n_11656, n19120);
  not g30684 (n_11657, n19123);
  and g30685 (n19124, n_11656, n_11657);
  not g30686 (n_11658, n19124);
  and g30687 (n19125, n_11656, n_11658);
  and g30688 (n19126, n_11657, n_11658);
  not g30689 (n_11659, n19125);
  not g30690 (n_11660, n19126);
  and g30691 (n19127, n_11659, n_11660);
  and g30692 (n19128, n18632, n18844);
  not g30693 (n_11661, n19128);
  and g30694 (n19129, n_11422, n_11661);
  and g30695 (n19130, n7101, n12531);
  and g30696 (n19131, n6402, n12537);
  and g30697 (n19132, n6951, n12534);
  not g30698 (n_11662, n19131);
  not g30699 (n_11663, n19132);
  and g30700 (n19133, n_11662, n_11663);
  not g30701 (n_11664, n19130);
  and g30702 (n19134, n_11664, n19133);
  and g30703 (n19135, n_1885, n19134);
  and g30704 (n19136, n_9870, n19134);
  not g30705 (n_11665, n19135);
  not g30706 (n_11666, n19136);
  and g30707 (n19137, n_11665, n_11666);
  not g30708 (n_11667, n19137);
  and g30709 (n19138, \a[14] , n_11667);
  and g30710 (n19139, n_652, n19137);
  not g30711 (n_11668, n19138);
  not g30712 (n_11669, n19139);
  and g30713 (n19140, n_11668, n_11669);
  not g30714 (n_11670, n19140);
  and g30715 (n19141, n19129, n_11670);
  and g30716 (n19142, n18650, n18842);
  not g30717 (n_11671, n19142);
  and g30718 (n19143, n_11419, n_11671);
  and g30719 (n19144, n7101, n12534);
  and g30720 (n19145, n6402, n12540);
  and g30721 (n19146, n6951, n12537);
  not g30722 (n_11672, n19145);
  not g30723 (n_11673, n19146);
  and g30724 (n19147, n_11672, n_11673);
  not g30725 (n_11674, n19144);
  and g30726 (n19148, n_11674, n19147);
  and g30727 (n19149, n_1885, n19148);
  and g30728 (n19150, n15096, n19148);
  not g30729 (n_11675, n19149);
  not g30730 (n_11676, n19150);
  and g30731 (n19151, n_11675, n_11676);
  not g30732 (n_11677, n19151);
  and g30733 (n19152, \a[14] , n_11677);
  and g30734 (n19153, n_652, n19151);
  not g30735 (n_11678, n19152);
  not g30736 (n_11679, n19153);
  and g30737 (n19154, n_11678, n_11679);
  not g30738 (n_11680, n19154);
  and g30739 (n19155, n19143, n_11680);
  and g30740 (n19156, n18668, n18840);
  not g30741 (n_11681, n19156);
  and g30742 (n19157, n_11416, n_11681);
  and g30743 (n19158, n7101, n12537);
  and g30744 (n19159, n6402, n12543);
  and g30745 (n19160, n6951, n12540);
  not g30746 (n_11682, n19159);
  not g30747 (n_11683, n19160);
  and g30748 (n19161, n_11682, n_11683);
  not g30749 (n_11684, n19158);
  and g30750 (n19162, n_11684, n19161);
  and g30751 (n19163, n_1885, n19162);
  and g30752 (n19164, n15385, n19162);
  not g30753 (n_11685, n19163);
  not g30754 (n_11686, n19164);
  and g30755 (n19165, n_11685, n_11686);
  not g30756 (n_11687, n19165);
  and g30757 (n19166, \a[14] , n_11687);
  and g30758 (n19167, n_652, n19165);
  not g30759 (n_11688, n19166);
  not g30760 (n_11689, n19167);
  and g30761 (n19168, n_11688, n_11689);
  not g30762 (n_11690, n19168);
  and g30763 (n19169, n19157, n_11690);
  and g30764 (n19170, n7101, n12540);
  and g30765 (n19171, n6402, n12546);
  and g30766 (n19172, n6951, n12543);
  and g30772 (n19175, n6397, n_8936);
  not g30775 (n_11695, n19176);
  and g30776 (n19177, \a[14] , n_11695);
  not g30777 (n_11696, n19177);
  and g30778 (n19178, n_11695, n_11696);
  and g30779 (n19179, \a[14] , n_11696);
  not g30780 (n_11697, n19178);
  not g30781 (n_11698, n19179);
  and g30782 (n19180, n_11697, n_11698);
  not g30783 (n_11699, n18838);
  and g30784 (n19181, n18836, n_11699);
  not g30785 (n_11700, n19181);
  and g30786 (n19182, n_11413, n_11700);
  not g30787 (n_11701, n19180);
  and g30788 (n19183, n_11701, n19182);
  not g30789 (n_11702, n19183);
  and g30790 (n19184, n_11701, n_11702);
  and g30791 (n19185, n19182, n_11702);
  not g30792 (n_11703, n19184);
  not g30793 (n_11704, n19185);
  and g30794 (n19186, n_11703, n_11704);
  and g30795 (n19187, n7101, n12543);
  and g30796 (n19188, n6402, n12549);
  and g30797 (n19189, n6951, n12546);
  and g30803 (n19192, n6397, n15724);
  not g30806 (n_11709, n19193);
  and g30807 (n19194, \a[14] , n_11709);
  not g30808 (n_11710, n19194);
  and g30809 (n19195, n_11709, n_11710);
  and g30810 (n19196, \a[14] , n_11710);
  not g30811 (n_11711, n19195);
  not g30812 (n_11712, n19196);
  and g30813 (n19197, n_11711, n_11712);
  and g30814 (n19198, n_11406, n_11408);
  and g30815 (n19199, n_11407, n_11408);
  not g30816 (n_11713, n19198);
  not g30817 (n_11714, n19199);
  and g30818 (n19200, n_11713, n_11714);
  not g30819 (n_11715, n19197);
  not g30820 (n_11716, n19200);
  and g30821 (n19201, n_11715, n_11716);
  not g30822 (n_11717, n19201);
  and g30823 (n19202, n_11715, n_11717);
  and g30824 (n19203, n_11716, n_11717);
  not g30825 (n_11718, n19202);
  not g30826 (n_11719, n19203);
  and g30827 (n19204, n_11718, n_11719);
  and g30828 (n19205, n7101, n12546);
  and g30829 (n19206, n6402, n12552);
  and g30830 (n19207, n6951, n12549);
  and g30836 (n19210, n6397, n_8634);
  not g30839 (n_11724, n19211);
  and g30840 (n19212, \a[14] , n_11724);
  not g30841 (n_11725, n19212);
  and g30842 (n19213, n_11724, n_11725);
  and g30843 (n19214, \a[14] , n_11725);
  not g30844 (n_11726, n19213);
  not g30845 (n_11727, n19214);
  and g30846 (n19215, n_11726, n_11727);
  and g30847 (n19216, n_11400, n_11402);
  and g30848 (n19217, n_11401, n_11402);
  not g30849 (n_11728, n19216);
  not g30850 (n_11729, n19217);
  and g30851 (n19218, n_11728, n_11729);
  not g30852 (n_11730, n19215);
  not g30853 (n_11731, n19218);
  and g30854 (n19219, n_11730, n_11731);
  not g30855 (n_11732, n19219);
  and g30856 (n19220, n_11730, n_11732);
  and g30857 (n19221, n_11731, n_11732);
  not g30858 (n_11733, n19220);
  not g30859 (n_11734, n19221);
  and g30860 (n19222, n_11733, n_11734);
  and g30861 (n19223, n18727, n18824);
  not g30862 (n_11735, n19223);
  and g30863 (n19224, n_11396, n_11735);
  and g30864 (n19225, n7101, n12549);
  and g30865 (n19226, n6402, n12555);
  and g30866 (n19227, n6951, n12552);
  not g30867 (n_11736, n19226);
  not g30868 (n_11737, n19227);
  and g30869 (n19228, n_11736, n_11737);
  not g30870 (n_11738, n19225);
  and g30871 (n19229, n_11738, n19228);
  and g30872 (n19230, n_1885, n19229);
  and g30873 (n19231, n_9580, n19229);
  not g30874 (n_11739, n19230);
  not g30875 (n_11740, n19231);
  and g30876 (n19232, n_11739, n_11740);
  not g30877 (n_11741, n19232);
  and g30878 (n19233, \a[14] , n_11741);
  and g30879 (n19234, n_652, n19232);
  not g30880 (n_11742, n19233);
  not g30881 (n_11743, n19234);
  and g30882 (n19235, n_11742, n_11743);
  not g30883 (n_11744, n19235);
  and g30884 (n19236, n19224, n_11744);
  not g30885 (n_11745, n18822);
  and g30886 (n19237, n18820, n_11745);
  not g30887 (n_11746, n19237);
  and g30888 (n19238, n_11393, n_11746);
  and g30889 (n19239, n7101, n12552);
  and g30890 (n19240, n6402, n12558);
  and g30891 (n19241, n6951, n12555);
  not g30892 (n_11747, n19240);
  not g30893 (n_11748, n19241);
  and g30894 (n19242, n_11747, n_11748);
  not g30895 (n_11749, n19239);
  and g30896 (n19243, n_11749, n19242);
  and g30897 (n19244, n_1885, n19243);
  and g30898 (n19245, n15791, n19243);
  not g30899 (n_11750, n19244);
  not g30900 (n_11751, n19245);
  and g30901 (n19246, n_11750, n_11751);
  not g30902 (n_11752, n19246);
  and g30903 (n19247, \a[14] , n_11752);
  and g30904 (n19248, n_652, n19246);
  not g30905 (n_11753, n19247);
  not g30906 (n_11754, n19248);
  and g30907 (n19249, n_11753, n_11754);
  not g30908 (n_11755, n19249);
  and g30909 (n19250, n19238, n_11755);
  and g30910 (n19251, n18759, n18818);
  not g30911 (n_11756, n19251);
  and g30912 (n19252, n_11389, n_11756);
  and g30913 (n19253, n7101, n12555);
  and g30914 (n19254, n6402, n12561);
  and g30915 (n19255, n6951, n12558);
  not g30916 (n_11757, n19254);
  not g30917 (n_11758, n19255);
  and g30918 (n19256, n_11757, n_11758);
  not g30919 (n_11759, n19253);
  and g30920 (n19257, n_11759, n19256);
  and g30921 (n19258, n_1885, n19257);
  and g30922 (n19259, n15816, n19257);
  not g30923 (n_11760, n19258);
  not g30924 (n_11761, n19259);
  and g30925 (n19260, n_11760, n_11761);
  not g30926 (n_11762, n19260);
  and g30927 (n19261, \a[14] , n_11762);
  and g30928 (n19262, n_652, n19260);
  not g30929 (n_11763, n19261);
  not g30930 (n_11764, n19262);
  and g30931 (n19263, n_11763, n_11764);
  not g30932 (n_11765, n19263);
  and g30933 (n19264, n19252, n_11765);
  and g30934 (n19265, n7101, n12558);
  and g30935 (n19266, n6402, n12564);
  and g30936 (n19267, n6951, n12561);
  and g30942 (n19270, n6397, n15847);
  not g30945 (n_11770, n19271);
  and g30946 (n19272, \a[14] , n_11770);
  not g30947 (n_11771, n19272);
  and g30948 (n19273, n_11770, n_11771);
  and g30949 (n19274, \a[14] , n_11771);
  not g30950 (n_11772, n19273);
  not g30951 (n_11773, n19274);
  and g30952 (n19275, n_11772, n_11773);
  not g30953 (n_11774, n18816);
  and g30954 (n19276, n18814, n_11774);
  not g30955 (n_11775, n19276);
  and g30956 (n19277, n_11386, n_11775);
  not g30957 (n_11776, n19275);
  and g30958 (n19278, n_11776, n19277);
  not g30959 (n_11777, n19278);
  and g30960 (n19279, n_11776, n_11777);
  and g30961 (n19280, n19277, n_11777);
  not g30962 (n_11778, n19279);
  not g30963 (n_11779, n19280);
  and g30964 (n19281, n_11778, n_11779);
  and g30965 (n19282, n_11379, n_11381);
  and g30966 (n19283, n_11380, n_11381);
  not g30967 (n_11780, n19282);
  not g30968 (n_11781, n19283);
  and g30969 (n19284, n_11780, n_11781);
  and g30970 (n19285, n7101, n12561);
  and g30971 (n19286, n6402, n12567);
  and g30972 (n19287, n6951, n12564);
  not g30973 (n_11782, n19286);
  not g30974 (n_11783, n19287);
  and g30975 (n19288, n_11782, n_11783);
  not g30976 (n_11784, n19285);
  and g30977 (n19289, n_11784, n19288);
  and g30978 (n19290, n_1885, n19289);
  and g30979 (n19291, n15905, n19289);
  not g30980 (n_11785, n19290);
  not g30981 (n_11786, n19291);
  and g30982 (n19292, n_11785, n_11786);
  not g30983 (n_11787, n19292);
  and g30984 (n19293, \a[14] , n_11787);
  and g30985 (n19294, n_652, n19292);
  not g30986 (n_11788, n19293);
  not g30987 (n_11789, n19294);
  and g30988 (n19295, n_11788, n_11789);
  not g30989 (n_11790, n19284);
  not g30990 (n_11791, n19295);
  and g30991 (n19296, n_11790, n_11791);
  and g30992 (n19297, n7101, n12564);
  and g30993 (n19298, n6402, n12571);
  and g30994 (n19299, n6951, n12567);
  and g31000 (n19302, n6397, n_9006);
  not g31003 (n_11796, n19303);
  and g31004 (n19304, \a[14] , n_11796);
  not g31005 (n_11797, n19304);
  and g31006 (n19305, n_11796, n_11797);
  and g31007 (n19306, \a[14] , n_11797);
  not g31008 (n_11798, n19305);
  not g31009 (n_11799, n19306);
  and g31010 (n19307, n_11798, n_11799);
  not g31011 (n_11800, n18785);
  and g31012 (n19308, n_11800, n18796);
  not g31013 (n_11801, n18797);
  not g31014 (n_11802, n19308);
  and g31015 (n19309, n_11801, n_11802);
  not g31016 (n_11803, n19307);
  and g31017 (n19310, n_11803, n19309);
  not g31018 (n_11804, n19310);
  and g31019 (n19311, n_11803, n_11804);
  and g31020 (n19312, n19309, n_11804);
  not g31021 (n_11805, n19311);
  not g31022 (n_11806, n19312);
  and g31023 (n19313, n_11805, n_11806);
  not g31024 (n_11807, n18784);
  and g31025 (n19314, n18782, n_11807);
  not g31026 (n_11808, n19314);
  and g31027 (n19315, n_11800, n_11808);
  and g31028 (n19316, n7101, n12567);
  and g31029 (n19317, n6402, n12574);
  and g31030 (n19318, n6951, n12571);
  not g31031 (n_11809, n19317);
  not g31032 (n_11810, n19318);
  and g31033 (n19319, n_11809, n_11810);
  not g31034 (n_11811, n19316);
  and g31035 (n19320, n_11811, n19319);
  and g31036 (n19321, n_1885, n19320);
  and g31037 (n19322, n_10006, n19320);
  not g31038 (n_11812, n19321);
  not g31039 (n_11813, n19322);
  and g31040 (n19323, n_11812, n_11813);
  not g31041 (n_11814, n19323);
  and g31042 (n19324, \a[14] , n_11814);
  and g31043 (n19325, n_652, n19323);
  not g31044 (n_11815, n19324);
  not g31045 (n_11816, n19325);
  and g31046 (n19326, n_11815, n_11816);
  not g31047 (n_11817, n19326);
  and g31048 (n19327, n19315, n_11817);
  and g31049 (n19328, n6951, n_6977);
  and g31050 (n19329, n7101, n12577);
  not g31051 (n_11818, n19328);
  not g31052 (n_11819, n19329);
  and g31053 (n19330, n_11818, n_11819);
  and g31054 (n19331, n6397, n_9032);
  not g31055 (n_11820, n19331);
  and g31056 (n19332, n19330, n_11820);
  not g31057 (n_11821, n19332);
  and g31058 (n19333, \a[14] , n_11821);
  not g31059 (n_11822, n19333);
  and g31060 (n19334, \a[14] , n_11822);
  and g31061 (n19335, n_11821, n_11822);
  not g31062 (n_11823, n19334);
  not g31063 (n_11824, n19335);
  and g31064 (n19336, n_11823, n_11824);
  and g31065 (n19337, n_1881, n_6977);
  not g31066 (n_11825, n19337);
  and g31067 (n19338, \a[14] , n_11825);
  not g31068 (n_11826, n19336);
  and g31069 (n19339, n_11826, n19338);
  and g31070 (n19340, n7101, n12574);
  and g31071 (n19341, n6402, n_6977);
  and g31072 (n19342, n6951, n12577);
  not g31073 (n_11827, n19341);
  not g31074 (n_11828, n19342);
  and g31075 (n19343, n_11827, n_11828);
  not g31076 (n_11829, n19340);
  and g31077 (n19344, n_11829, n19343);
  and g31078 (n19345, n_1885, n19344);
  and g31079 (n19346, n16094, n19344);
  not g31080 (n_11830, n19345);
  not g31081 (n_11831, n19346);
  and g31082 (n19347, n_11830, n_11831);
  not g31083 (n_11832, n19347);
  and g31084 (n19348, \a[14] , n_11832);
  and g31085 (n19349, n_652, n19347);
  not g31086 (n_11833, n19348);
  not g31087 (n_11834, n19349);
  and g31088 (n19350, n_11833, n_11834);
  not g31089 (n_11835, n19350);
  and g31090 (n19351, n19339, n_11835);
  and g31091 (n19352, n18783, n19351);
  not g31092 (n_11836, n19352);
  and g31093 (n19353, n19351, n_11836);
  and g31094 (n19354, n18783, n_11836);
  not g31095 (n_11837, n19353);
  not g31096 (n_11838, n19354);
  and g31097 (n19355, n_11837, n_11838);
  and g31098 (n19356, n7101, n12571);
  and g31099 (n19357, n6402, n12577);
  and g31100 (n19358, n6951, n12574);
  and g31106 (n19361, n6397, n16013);
  not g31109 (n_11843, n19362);
  and g31110 (n19363, \a[14] , n_11843);
  not g31111 (n_11844, n19363);
  and g31112 (n19364, \a[14] , n_11844);
  and g31113 (n19365, n_11843, n_11844);
  not g31114 (n_11845, n19364);
  not g31115 (n_11846, n19365);
  and g31116 (n19366, n_11845, n_11846);
  not g31117 (n_11847, n19355);
  not g31118 (n_11848, n19366);
  and g31119 (n19367, n_11847, n_11848);
  not g31120 (n_11849, n19367);
  and g31121 (n19368, n_11836, n_11849);
  not g31122 (n_11850, n19315);
  and g31123 (n19369, n_11850, n19326);
  not g31124 (n_11851, n19327);
  not g31125 (n_11852, n19369);
  and g31126 (n19370, n_11851, n_11852);
  not g31127 (n_11853, n19368);
  and g31128 (n19371, n_11853, n19370);
  not g31129 (n_11854, n19371);
  and g31130 (n19372, n_11851, n_11854);
  not g31131 (n_11855, n19313);
  not g31132 (n_11856, n19372);
  and g31133 (n19373, n_11855, n_11856);
  not g31134 (n_11857, n19373);
  and g31135 (n19374, n_11804, n_11857);
  and g31136 (n19375, n19284, n19295);
  not g31137 (n_11858, n19296);
  not g31138 (n_11859, n19375);
  and g31139 (n19376, n_11858, n_11859);
  not g31140 (n_11860, n19374);
  and g31141 (n19377, n_11860, n19376);
  not g31142 (n_11861, n19377);
  and g31143 (n19378, n_11858, n_11861);
  not g31144 (n_11862, n19281);
  not g31145 (n_11863, n19378);
  and g31146 (n19379, n_11862, n_11863);
  not g31147 (n_11864, n19379);
  and g31148 (n19380, n_11777, n_11864);
  not g31149 (n_11865, n19264);
  and g31150 (n19381, n19252, n_11865);
  and g31151 (n19382, n_11765, n_11865);
  not g31152 (n_11866, n19381);
  not g31153 (n_11867, n19382);
  and g31154 (n19383, n_11866, n_11867);
  not g31155 (n_11868, n19380);
  not g31156 (n_11869, n19383);
  and g31157 (n19384, n_11868, n_11869);
  not g31158 (n_11870, n19384);
  and g31159 (n19385, n_11865, n_11870);
  not g31160 (n_11871, n19250);
  and g31161 (n19386, n19238, n_11871);
  and g31162 (n19387, n_11755, n_11871);
  not g31163 (n_11872, n19386);
  not g31164 (n_11873, n19387);
  and g31165 (n19388, n_11872, n_11873);
  not g31166 (n_11874, n19385);
  not g31167 (n_11875, n19388);
  and g31168 (n19389, n_11874, n_11875);
  not g31169 (n_11876, n19389);
  and g31170 (n19390, n_11871, n_11876);
  not g31171 (n_11877, n19224);
  and g31172 (n19391, n_11877, n19235);
  not g31173 (n_11878, n19236);
  not g31174 (n_11879, n19391);
  and g31175 (n19392, n_11878, n_11879);
  not g31176 (n_11880, n19390);
  and g31177 (n19393, n_11880, n19392);
  not g31178 (n_11881, n19393);
  and g31179 (n19394, n_11878, n_11881);
  not g31180 (n_11882, n19222);
  not g31181 (n_11883, n19394);
  and g31182 (n19395, n_11882, n_11883);
  not g31183 (n_11884, n19395);
  and g31184 (n19396, n_11732, n_11884);
  not g31185 (n_11885, n19204);
  not g31186 (n_11886, n19396);
  and g31187 (n19397, n_11885, n_11886);
  not g31188 (n_11887, n19397);
  and g31189 (n19398, n_11717, n_11887);
  not g31190 (n_11888, n19186);
  not g31191 (n_11889, n19398);
  and g31192 (n19399, n_11888, n_11889);
  not g31193 (n_11890, n19399);
  and g31194 (n19400, n_11702, n_11890);
  not g31195 (n_11891, n19169);
  and g31196 (n19401, n19157, n_11891);
  and g31197 (n19402, n_11690, n_11891);
  not g31198 (n_11892, n19401);
  not g31199 (n_11893, n19402);
  and g31200 (n19403, n_11892, n_11893);
  not g31201 (n_11894, n19400);
  not g31202 (n_11895, n19403);
  and g31203 (n19404, n_11894, n_11895);
  not g31204 (n_11896, n19404);
  and g31205 (n19405, n_11891, n_11896);
  not g31206 (n_11897, n19155);
  and g31207 (n19406, n19143, n_11897);
  and g31208 (n19407, n_11680, n_11897);
  not g31209 (n_11898, n19406);
  not g31210 (n_11899, n19407);
  and g31211 (n19408, n_11898, n_11899);
  not g31212 (n_11900, n19405);
  not g31213 (n_11901, n19408);
  and g31214 (n19409, n_11900, n_11901);
  not g31215 (n_11902, n19409);
  and g31216 (n19410, n_11897, n_11902);
  not g31217 (n_11903, n19129);
  and g31218 (n19411, n_11903, n19140);
  not g31219 (n_11904, n19141);
  not g31220 (n_11905, n19411);
  and g31221 (n19412, n_11904, n_11905);
  not g31222 (n_11906, n19410);
  and g31223 (n19413, n_11906, n19412);
  not g31224 (n_11907, n19413);
  and g31225 (n19414, n_11904, n_11907);
  not g31226 (n_11908, n19127);
  not g31227 (n_11909, n19414);
  and g31228 (n19415, n_11908, n_11909);
  not g31229 (n_11910, n19415);
  and g31230 (n19416, n_11658, n_11910);
  not g31231 (n_11911, n19109);
  not g31232 (n_11912, n19416);
  and g31233 (n19417, n_11911, n_11912);
  not g31234 (n_11913, n19417);
  and g31235 (n19418, n_11643, n_11913);
  not g31236 (n_11914, n19092);
  and g31237 (n19419, n19080, n_11914);
  and g31238 (n19420, n_11631, n_11914);
  not g31239 (n_11915, n19419);
  not g31240 (n_11916, n19420);
  and g31241 (n19421, n_11915, n_11916);
  not g31242 (n_11917, n19418);
  not g31243 (n_11918, n19421);
  and g31244 (n19422, n_11917, n_11918);
  not g31245 (n_11919, n19422);
  and g31246 (n19423, n_11914, n_11919);
  not g31247 (n_11920, n19078);
  and g31248 (n19424, n19066, n_11920);
  and g31249 (n19425, n_11621, n_11920);
  not g31250 (n_11921, n19424);
  not g31251 (n_11922, n19425);
  and g31252 (n19426, n_11921, n_11922);
  not g31253 (n_11923, n19423);
  not g31254 (n_11924, n19426);
  and g31255 (n19427, n_11923, n_11924);
  not g31256 (n_11925, n19427);
  and g31257 (n19428, n_11920, n_11925);
  not g31258 (n_11926, n19064);
  and g31259 (n19429, n19052, n_11926);
  and g31260 (n19430, n_11611, n_11926);
  not g31261 (n_11927, n19429);
  not g31262 (n_11928, n19430);
  and g31263 (n19431, n_11927, n_11928);
  not g31264 (n_11929, n19428);
  not g31265 (n_11930, n19431);
  and g31266 (n19432, n_11929, n_11930);
  not g31267 (n_11931, n19432);
  and g31268 (n19433, n_11926, n_11931);
  not g31269 (n_11932, n19050);
  and g31270 (n19434, n19038, n_11932);
  and g31271 (n19435, n_11601, n_11932);
  not g31272 (n_11933, n19434);
  not g31273 (n_11934, n19435);
  and g31274 (n19436, n_11933, n_11934);
  not g31275 (n_11935, n19433);
  not g31276 (n_11936, n19436);
  and g31277 (n19437, n_11935, n_11936);
  not g31278 (n_11937, n19437);
  and g31279 (n19438, n_11932, n_11937);
  not g31280 (n_11938, n19036);
  and g31281 (n19439, n19024, n_11938);
  and g31282 (n19440, n_11591, n_11938);
  not g31283 (n_11939, n19439);
  not g31284 (n_11940, n19440);
  and g31285 (n19441, n_11939, n_11940);
  not g31286 (n_11941, n19438);
  not g31287 (n_11942, n19441);
  and g31288 (n19442, n_11941, n_11942);
  not g31289 (n_11943, n19442);
  and g31290 (n19443, n_11938, n_11943);
  not g31291 (n_11944, n19022);
  and g31292 (n19444, n19010, n_11944);
  and g31293 (n19445, n_11580, n_11944);
  not g31294 (n_11945, n19444);
  not g31295 (n_11946, n19445);
  and g31296 (n19446, n_11945, n_11946);
  not g31297 (n_11947, n19443);
  not g31298 (n_11948, n19446);
  and g31299 (n19447, n_11947, n_11948);
  not g31300 (n_11949, n19447);
  and g31301 (n19448, n_11944, n_11949);
  not g31302 (n_11950, n19008);
  and g31303 (n19449, n18996, n_11950);
  and g31304 (n19450, n_11570, n_11950);
  not g31305 (n_11951, n19449);
  not g31306 (n_11952, n19450);
  and g31307 (n19451, n_11951, n_11952);
  not g31308 (n_11953, n19448);
  not g31309 (n_11954, n19451);
  and g31310 (n19452, n_11953, n_11954);
  not g31311 (n_11955, n19452);
  and g31312 (n19453, n_11950, n_11955);
  not g31313 (n_11956, n18994);
  and g31314 (n19454, n18982, n_11956);
  and g31315 (n19455, n_11560, n_11956);
  not g31316 (n_11957, n19454);
  not g31317 (n_11958, n19455);
  and g31318 (n19456, n_11957, n_11958);
  not g31319 (n_11959, n19453);
  not g31320 (n_11960, n19456);
  and g31321 (n19457, n_11959, n_11960);
  not g31322 (n_11961, n19457);
  and g31323 (n19458, n_11956, n_11961);
  not g31324 (n_11962, n18980);
  and g31325 (n19459, n18968, n_11962);
  and g31326 (n19460, n_11550, n_11962);
  not g31327 (n_11963, n19459);
  not g31328 (n_11964, n19460);
  and g31329 (n19461, n_11963, n_11964);
  not g31330 (n_11965, n19458);
  not g31331 (n_11966, n19461);
  and g31332 (n19462, n_11965, n_11966);
  not g31333 (n_11967, n19462);
  and g31334 (n19463, n_11962, n_11967);
  not g31335 (n_11968, n18954);
  and g31336 (n19464, n_11968, n18965);
  not g31337 (n_11969, n18966);
  not g31338 (n_11970, n19464);
  and g31339 (n19465, n_11969, n_11970);
  not g31340 (n_11971, n19463);
  and g31341 (n19466, n_11971, n19465);
  not g31342 (n_11972, n19466);
  and g31343 (n19467, n_11969, n_11972);
  not g31344 (n_11973, n18952);
  not g31345 (n_11974, n19467);
  and g31346 (n19468, n_11973, n_11974);
  and g31347 (n19469, n18952, n19467);
  not g31348 (n_11975, n19468);
  not g31349 (n_11976, n19469);
  and g31350 (n19470, n_11975, n_11976);
  and g31351 (n19471, n7983, n13521);
  and g31352 (n19472, n7291, n13491);
  and g31353 (n19473, n7632, n13518);
  and g31359 (n19476, n7294, n_7677);
  not g31362 (n_11981, n19477);
  and g31363 (n19478, \a[11] , n_11981);
  not g31364 (n_11982, n19478);
  and g31365 (n19479, \a[11] , n_11982);
  and g31366 (n19480, n_11981, n_11982);
  not g31367 (n_11983, n19479);
  not g31368 (n_11984, n19480);
  and g31369 (n19481, n_11983, n_11984);
  not g31370 (n_11985, n19481);
  and g31371 (n19482, n19470, n_11985);
  not g31372 (n_11986, n19482);
  and g31373 (n19483, n_11975, n_11986);
  not g31374 (n_11987, n18949);
  not g31375 (n_11988, n19483);
  and g31376 (n19484, n_11987, n_11988);
  and g31377 (n19485, n18949, n19483);
  not g31378 (n_11989, n19484);
  not g31379 (n_11990, n19485);
  and g31380 (n19486, n_11989, n_11990);
  and g31381 (n19487, n9331, n13633);
  and g31382 (n19488, n8418, n13597);
  and g31383 (n19489, n8860, n13630);
  and g31389 (n19492, n8421, n13929);
  not g31392 (n_11995, n19493);
  and g31393 (n19494, \a[8] , n_11995);
  not g31394 (n_11996, n19494);
  and g31395 (n19495, \a[8] , n_11996);
  and g31396 (n19496, n_11995, n_11996);
  not g31397 (n_11997, n19495);
  not g31398 (n_11998, n19496);
  and g31399 (n19497, n_11997, n_11998);
  not g31400 (n_11999, n19497);
  and g31401 (n19498, n19486, n_11999);
  not g31402 (n_12000, n19498);
  and g31403 (n19499, n_11989, n_12000);
  not g31404 (n_12001, n15076);
  and g31405 (n19500, n_7417, n_12001);
  and g31406 (n19501, n9867, n13941);
  not g31407 (n_12002, n19500);
  not g31408 (n_12003, n19501);
  and g31409 (n19502, n_12002, n_12003);
  and g31410 (n19503, n_4684, n19502);
  and g31411 (n19504, n13951, n19502);
  not g31412 (n_12004, n19503);
  not g31413 (n_12005, n19504);
  and g31414 (n19505, n_12004, n_12005);
  not g31415 (n_12006, n19505);
  and g31416 (n19506, \a[5] , n_12006);
  and g31417 (n19507, n_3, n19505);
  not g31418 (n_12007, n19506);
  not g31419 (n_12008, n19507);
  and g31420 (n19508, n_12007, n_12008);
  not g31421 (n_12009, n19499);
  not g31422 (n_12010, n19508);
  and g31423 (n19509, n_12009, n_12010);
  and g31424 (n19510, n18910, n_11505);
  and g31425 (n19511, n_11504, n_11505);
  not g31426 (n_12011, n19510);
  not g31427 (n_12012, n19511);
  and g31428 (n19512, n_12011, n_12012);
  and g31429 (n19513, n19499, n19508);
  not g31430 (n_12013, n19509);
  not g31431 (n_12014, n19513);
  and g31432 (n19514, n_12013, n_12014);
  not g31433 (n_12015, n19512);
  and g31434 (n19515, n_12015, n19514);
  not g31435 (n_12016, n19515);
  and g31436 (n19516, n_12013, n_12016);
  not g31437 (n_12017, n18940);
  and g31438 (n19517, n18938, n_12017);
  not g31439 (n_12018, n19517);
  and g31440 (n19518, n_11521, n_12018);
  not g31441 (n_12019, n19516);
  and g31442 (n19519, n_12019, n19518);
  and g31443 (n19520, n_12015, n_12016);
  and g31444 (n19521, n19514, n_12016);
  not g31445 (n_12020, n19520);
  not g31446 (n_12021, n19521);
  and g31447 (n19522, n_12020, n_12021);
  and g31448 (n19523, n19486, n_12000);
  and g31449 (n19524, n_11999, n_12000);
  not g31450 (n_12022, n19523);
  not g31451 (n_12023, n19524);
  and g31452 (n19525, n_12022, n_12023);
  and g31453 (n19526, n19470, n_11986);
  and g31454 (n19527, n_11985, n_11986);
  not g31455 (n_12024, n19526);
  not g31456 (n_12025, n19527);
  and g31457 (n19528, n_12024, n_12025);
  and g31458 (n19529, n7983, n13518);
  and g31459 (n19530, n7291, n12889);
  and g31460 (n19531, n7632, n13491);
  and g31466 (n19534, n7294, n13584);
  not g31469 (n_12030, n19535);
  and g31470 (n19536, \a[11] , n_12030);
  not g31471 (n_12031, n19536);
  and g31472 (n19537, n_12030, n_12031);
  and g31473 (n19538, \a[11] , n_12031);
  not g31474 (n_12032, n19537);
  not g31475 (n_12033, n19538);
  and g31476 (n19539, n_12032, n_12033);
  not g31477 (n_12034, n19465);
  and g31478 (n19540, n19463, n_12034);
  not g31479 (n_12035, n19540);
  and g31480 (n19541, n_11972, n_12035);
  not g31481 (n_12036, n19539);
  and g31482 (n19542, n_12036, n19541);
  not g31483 (n_12037, n19542);
  and g31484 (n19543, n_12036, n_12037);
  and g31485 (n19544, n19541, n_12037);
  not g31486 (n_12038, n19543);
  not g31487 (n_12039, n19544);
  and g31488 (n19545, n_12038, n_12039);
  and g31489 (n19546, n7983, n13491);
  and g31490 (n19547, n7291, n12769);
  and g31491 (n19548, n7632, n12889);
  and g31497 (n19551, n7294, n_7447);
  not g31500 (n_12044, n19552);
  and g31501 (n19553, \a[11] , n_12044);
  not g31502 (n_12045, n19553);
  and g31503 (n19554, n_12044, n_12045);
  and g31504 (n19555, \a[11] , n_12045);
  not g31505 (n_12046, n19554);
  not g31506 (n_12047, n19555);
  and g31507 (n19556, n_12046, n_12047);
  and g31508 (n19557, n_11965, n_11967);
  and g31509 (n19558, n_11966, n_11967);
  not g31510 (n_12048, n19557);
  not g31511 (n_12049, n19558);
  and g31512 (n19559, n_12048, n_12049);
  not g31513 (n_12050, n19556);
  not g31514 (n_12051, n19559);
  and g31515 (n19560, n_12050, n_12051);
  not g31516 (n_12052, n19560);
  and g31517 (n19561, n_12050, n_12052);
  and g31518 (n19562, n_12051, n_12052);
  not g31519 (n_12053, n19561);
  not g31520 (n_12054, n19562);
  and g31521 (n19563, n_12053, n_12054);
  and g31522 (n19564, n7983, n12889);
  and g31523 (n19565, n7291, n12502);
  and g31524 (n19566, n7632, n12769);
  and g31530 (n19569, n7294, n12895);
  not g31533 (n_12059, n19570);
  and g31534 (n19571, \a[11] , n_12059);
  not g31535 (n_12060, n19571);
  and g31536 (n19572, n_12059, n_12060);
  and g31537 (n19573, \a[11] , n_12060);
  not g31538 (n_12061, n19572);
  not g31539 (n_12062, n19573);
  and g31540 (n19574, n_12061, n_12062);
  and g31541 (n19575, n_11959, n_11961);
  and g31542 (n19576, n_11960, n_11961);
  not g31543 (n_12063, n19575);
  not g31544 (n_12064, n19576);
  and g31545 (n19577, n_12063, n_12064);
  not g31546 (n_12065, n19574);
  not g31547 (n_12066, n19577);
  and g31548 (n19578, n_12065, n_12066);
  not g31549 (n_12067, n19578);
  and g31550 (n19579, n_12065, n_12067);
  and g31551 (n19580, n_12066, n_12067);
  not g31552 (n_12068, n19579);
  not g31553 (n_12069, n19580);
  and g31554 (n19581, n_12068, n_12069);
  and g31555 (n19582, n7983, n12769);
  and g31556 (n19583, n7291, n12370);
  and g31557 (n19584, n7632, n12502);
  and g31563 (n19587, n7294, n12999);
  not g31566 (n_12074, n19588);
  and g31567 (n19589, \a[11] , n_12074);
  not g31568 (n_12075, n19589);
  and g31569 (n19590, n_12074, n_12075);
  and g31570 (n19591, \a[11] , n_12075);
  not g31571 (n_12076, n19590);
  not g31572 (n_12077, n19591);
  and g31573 (n19592, n_12076, n_12077);
  and g31574 (n19593, n_11953, n_11955);
  and g31575 (n19594, n_11954, n_11955);
  not g31576 (n_12078, n19593);
  not g31577 (n_12079, n19594);
  and g31578 (n19595, n_12078, n_12079);
  not g31579 (n_12080, n19592);
  not g31580 (n_12081, n19595);
  and g31581 (n19596, n_12080, n_12081);
  not g31582 (n_12082, n19596);
  and g31583 (n19597, n_12080, n_12082);
  and g31584 (n19598, n_12081, n_12082);
  not g31585 (n_12083, n19597);
  not g31586 (n_12084, n19598);
  and g31587 (n19599, n_12083, n_12084);
  and g31588 (n19600, n7983, n12502);
  and g31589 (n19601, n7291, n12505);
  and g31590 (n19602, n7632, n12370);
  and g31596 (n19605, n7294, n_7594);
  not g31599 (n_12089, n19606);
  and g31600 (n19607, \a[11] , n_12089);
  not g31601 (n_12090, n19607);
  and g31602 (n19608, n_12089, n_12090);
  and g31603 (n19609, \a[11] , n_12090);
  not g31604 (n_12091, n19608);
  not g31605 (n_12092, n19609);
  and g31606 (n19610, n_12091, n_12092);
  and g31607 (n19611, n_11947, n_11949);
  and g31608 (n19612, n_11948, n_11949);
  not g31609 (n_12093, n19611);
  not g31610 (n_12094, n19612);
  and g31611 (n19613, n_12093, n_12094);
  not g31612 (n_12095, n19610);
  not g31613 (n_12096, n19613);
  and g31614 (n19614, n_12095, n_12096);
  not g31615 (n_12097, n19614);
  and g31616 (n19615, n_12095, n_12097);
  and g31617 (n19616, n_12096, n_12097);
  not g31618 (n_12098, n19615);
  not g31619 (n_12099, n19616);
  and g31620 (n19617, n_12098, n_12099);
  and g31621 (n19618, n7983, n12370);
  and g31622 (n19619, n7291, n12508);
  and g31623 (n19620, n7632, n12505);
  and g31629 (n19623, n7294, n_7607);
  not g31632 (n_12104, n19624);
  and g31633 (n19625, \a[11] , n_12104);
  not g31634 (n_12105, n19625);
  and g31635 (n19626, n_12104, n_12105);
  and g31636 (n19627, \a[11] , n_12105);
  not g31637 (n_12106, n19626);
  not g31638 (n_12107, n19627);
  and g31639 (n19628, n_12106, n_12107);
  and g31640 (n19629, n_11941, n_11943);
  and g31641 (n19630, n_11942, n_11943);
  not g31642 (n_12108, n19629);
  not g31643 (n_12109, n19630);
  and g31644 (n19631, n_12108, n_12109);
  not g31645 (n_12110, n19628);
  not g31646 (n_12111, n19631);
  and g31647 (n19632, n_12110, n_12111);
  not g31648 (n_12112, n19632);
  and g31649 (n19633, n_12110, n_12112);
  and g31650 (n19634, n_12111, n_12112);
  not g31651 (n_12113, n19633);
  not g31652 (n_12114, n19634);
  and g31653 (n19635, n_12113, n_12114);
  and g31654 (n19636, n7983, n12505);
  and g31655 (n19637, n7291, n12513);
  and g31656 (n19638, n7632, n12508);
  and g31662 (n19641, n7294, n_7804);
  not g31665 (n_12119, n19642);
  and g31666 (n19643, \a[11] , n_12119);
  not g31667 (n_12120, n19643);
  and g31668 (n19644, n_12119, n_12120);
  and g31669 (n19645, \a[11] , n_12120);
  not g31670 (n_12121, n19644);
  not g31671 (n_12122, n19645);
  and g31672 (n19646, n_12121, n_12122);
  and g31673 (n19647, n_11935, n_11937);
  and g31674 (n19648, n_11936, n_11937);
  not g31675 (n_12123, n19647);
  not g31676 (n_12124, n19648);
  and g31677 (n19649, n_12123, n_12124);
  not g31678 (n_12125, n19646);
  not g31679 (n_12126, n19649);
  and g31680 (n19650, n_12125, n_12126);
  not g31681 (n_12127, n19650);
  and g31682 (n19651, n_12125, n_12127);
  and g31683 (n19652, n_12126, n_12127);
  not g31684 (n_12128, n19651);
  not g31685 (n_12129, n19652);
  and g31686 (n19653, n_12128, n_12129);
  and g31687 (n19654, n7983, n12508);
  and g31688 (n19655, n7291, n12511);
  and g31689 (n19656, n7632, n12513);
  and g31695 (n19659, n7294, n13863);
  not g31698 (n_12134, n19660);
  and g31699 (n19661, \a[11] , n_12134);
  not g31700 (n_12135, n19661);
  and g31701 (n19662, n_12134, n_12135);
  and g31702 (n19663, \a[11] , n_12135);
  not g31703 (n_12136, n19662);
  not g31704 (n_12137, n19663);
  and g31705 (n19664, n_12136, n_12137);
  and g31706 (n19665, n_11929, n_11931);
  and g31707 (n19666, n_11930, n_11931);
  not g31708 (n_12138, n19665);
  not g31709 (n_12139, n19666);
  and g31710 (n19667, n_12138, n_12139);
  not g31711 (n_12140, n19664);
  not g31712 (n_12141, n19667);
  and g31713 (n19668, n_12140, n_12141);
  not g31714 (n_12142, n19668);
  and g31715 (n19669, n_12140, n_12142);
  and g31716 (n19670, n_12141, n_12142);
  not g31717 (n_12143, n19669);
  not g31718 (n_12144, n19670);
  and g31719 (n19671, n_12143, n_12144);
  and g31720 (n19672, n7983, n12513);
  and g31721 (n19673, n7291, n12516);
  and g31722 (n19674, n7632, n12511);
  and g31728 (n19677, n7294, n14177);
  not g31731 (n_12149, n19678);
  and g31732 (n19679, \a[11] , n_12149);
  not g31733 (n_12150, n19679);
  and g31734 (n19680, n_12149, n_12150);
  and g31735 (n19681, \a[11] , n_12150);
  not g31736 (n_12151, n19680);
  not g31737 (n_12152, n19681);
  and g31738 (n19682, n_12151, n_12152);
  and g31739 (n19683, n_11923, n_11925);
  and g31740 (n19684, n_11924, n_11925);
  not g31741 (n_12153, n19683);
  not g31742 (n_12154, n19684);
  and g31743 (n19685, n_12153, n_12154);
  not g31744 (n_12155, n19682);
  not g31745 (n_12156, n19685);
  and g31746 (n19686, n_12155, n_12156);
  not g31747 (n_12157, n19686);
  and g31748 (n19687, n_12155, n_12157);
  and g31749 (n19688, n_12156, n_12157);
  not g31750 (n_12158, n19687);
  not g31751 (n_12159, n19688);
  and g31752 (n19689, n_12158, n_12159);
  and g31753 (n19690, n7983, n12511);
  and g31754 (n19691, n7291, n12519);
  and g31755 (n19692, n7632, n12516);
  and g31761 (n19695, n7294, n_7923);
  not g31764 (n_12164, n19696);
  and g31765 (n19697, \a[11] , n_12164);
  not g31766 (n_12165, n19697);
  and g31767 (n19698, n_12164, n_12165);
  and g31768 (n19699, \a[11] , n_12165);
  not g31769 (n_12166, n19698);
  not g31770 (n_12167, n19699);
  and g31771 (n19700, n_12166, n_12167);
  and g31772 (n19701, n_11917, n_11919);
  and g31773 (n19702, n_11918, n_11919);
  not g31774 (n_12168, n19701);
  not g31775 (n_12169, n19702);
  and g31776 (n19703, n_12168, n_12169);
  not g31777 (n_12170, n19700);
  not g31778 (n_12171, n19703);
  and g31779 (n19704, n_12170, n_12171);
  not g31780 (n_12172, n19704);
  and g31781 (n19705, n_12170, n_12172);
  and g31782 (n19706, n_12171, n_12172);
  not g31783 (n_12173, n19705);
  not g31784 (n_12174, n19706);
  and g31785 (n19707, n_12173, n_12174);
  and g31786 (n19708, n19109, n19416);
  not g31787 (n_12175, n19708);
  and g31788 (n19709, n_11913, n_12175);
  and g31789 (n19710, n7983, n12516);
  and g31790 (n19711, n7291, n12522);
  and g31791 (n19712, n7632, n12519);
  not g31792 (n_12176, n19711);
  not g31793 (n_12177, n19712);
  and g31794 (n19713, n_12176, n_12177);
  not g31795 (n_12178, n19710);
  and g31796 (n19714, n_12178, n19713);
  and g31797 (n19715, n_2446, n19714);
  and g31798 (n19716, n14443, n19714);
  not g31799 (n_12179, n19715);
  not g31800 (n_12180, n19716);
  and g31801 (n19717, n_12179, n_12180);
  not g31802 (n_12181, n19717);
  and g31803 (n19718, \a[11] , n_12181);
  and g31804 (n19719, n_1071, n19717);
  not g31805 (n_12182, n19718);
  not g31806 (n_12183, n19719);
  and g31807 (n19720, n_12182, n_12183);
  not g31808 (n_12184, n19720);
  and g31809 (n19721, n19709, n_12184);
  and g31810 (n19722, n19127, n19414);
  not g31811 (n_12185, n19722);
  and g31812 (n19723, n_11910, n_12185);
  and g31813 (n19724, n7983, n12519);
  and g31814 (n19725, n7291, n12525);
  and g31815 (n19726, n7632, n12522);
  not g31816 (n_12186, n19725);
  not g31817 (n_12187, n19726);
  and g31818 (n19727, n_12186, n_12187);
  not g31819 (n_12188, n19724);
  and g31820 (n19728, n_12188, n19727);
  and g31821 (n19729, n_2446, n19728);
  and g31822 (n19730, n_10664, n19728);
  not g31823 (n_12189, n19729);
  not g31824 (n_12190, n19730);
  and g31825 (n19731, n_12189, n_12190);
  not g31826 (n_12191, n19731);
  and g31827 (n19732, \a[11] , n_12191);
  and g31828 (n19733, n_1071, n19731);
  not g31829 (n_12192, n19732);
  not g31830 (n_12193, n19733);
  and g31831 (n19734, n_12192, n_12193);
  not g31832 (n_12194, n19734);
  and g31833 (n19735, n19723, n_12194);
  and g31834 (n19736, n7983, n12522);
  and g31835 (n19737, n7291, n12528);
  and g31836 (n19738, n7632, n12525);
  and g31842 (n19741, n7294, n14837);
  not g31845 (n_12199, n19742);
  and g31846 (n19743, \a[11] , n_12199);
  not g31847 (n_12200, n19743);
  and g31848 (n19744, n_12199, n_12200);
  and g31849 (n19745, \a[11] , n_12200);
  not g31850 (n_12201, n19744);
  not g31851 (n_12202, n19745);
  and g31852 (n19746, n_12201, n_12202);
  not g31853 (n_12203, n19412);
  and g31854 (n19747, n19410, n_12203);
  not g31855 (n_12204, n19747);
  and g31856 (n19748, n_11907, n_12204);
  not g31857 (n_12205, n19746);
  and g31858 (n19749, n_12205, n19748);
  not g31859 (n_12206, n19749);
  and g31860 (n19750, n_12205, n_12206);
  and g31861 (n19751, n19748, n_12206);
  not g31862 (n_12207, n19750);
  not g31863 (n_12208, n19751);
  and g31864 (n19752, n_12207, n_12208);
  and g31865 (n19753, n7983, n12525);
  and g31866 (n19754, n7291, n12531);
  and g31867 (n19755, n7632, n12528);
  and g31873 (n19758, n7294, n14608);
  not g31876 (n_12213, n19759);
  and g31877 (n19760, \a[11] , n_12213);
  not g31878 (n_12214, n19760);
  and g31879 (n19761, n_12213, n_12214);
  and g31880 (n19762, \a[11] , n_12214);
  not g31881 (n_12215, n19761);
  not g31882 (n_12216, n19762);
  and g31883 (n19763, n_12215, n_12216);
  and g31884 (n19764, n_11900, n_11902);
  and g31885 (n19765, n_11901, n_11902);
  not g31886 (n_12217, n19764);
  not g31887 (n_12218, n19765);
  and g31888 (n19766, n_12217, n_12218);
  not g31889 (n_12219, n19763);
  not g31890 (n_12220, n19766);
  and g31891 (n19767, n_12219, n_12220);
  not g31892 (n_12221, n19767);
  and g31893 (n19768, n_12219, n_12221);
  and g31894 (n19769, n_12220, n_12221);
  not g31895 (n_12222, n19768);
  not g31896 (n_12223, n19769);
  and g31897 (n19770, n_12222, n_12223);
  and g31898 (n19771, n7983, n12528);
  and g31899 (n19772, n7291, n12534);
  and g31900 (n19773, n7632, n12531);
  and g31906 (n19776, n7294, n_8448);
  not g31909 (n_12228, n19777);
  and g31910 (n19778, \a[11] , n_12228);
  not g31911 (n_12229, n19778);
  and g31912 (n19779, n_12228, n_12229);
  and g31913 (n19780, \a[11] , n_12229);
  not g31914 (n_12230, n19779);
  not g31915 (n_12231, n19780);
  and g31916 (n19781, n_12230, n_12231);
  and g31917 (n19782, n_11894, n_11896);
  and g31918 (n19783, n_11895, n_11896);
  not g31919 (n_12232, n19782);
  not g31920 (n_12233, n19783);
  and g31921 (n19784, n_12232, n_12233);
  not g31922 (n_12234, n19781);
  not g31923 (n_12235, n19784);
  and g31924 (n19785, n_12234, n_12235);
  not g31925 (n_12236, n19785);
  and g31926 (n19786, n_12234, n_12236);
  and g31927 (n19787, n_12235, n_12236);
  not g31928 (n_12237, n19786);
  not g31929 (n_12238, n19787);
  and g31930 (n19788, n_12237, n_12238);
  and g31931 (n19789, n19186, n19398);
  not g31932 (n_12239, n19789);
  and g31933 (n19790, n_11890, n_12239);
  and g31934 (n19791, n7983, n12531);
  and g31935 (n19792, n7291, n12537);
  and g31936 (n19793, n7632, n12534);
  not g31937 (n_12240, n19792);
  not g31938 (n_12241, n19793);
  and g31939 (n19794, n_12240, n_12241);
  not g31940 (n_12242, n19791);
  and g31941 (n19795, n_12242, n19794);
  and g31942 (n19796, n_2446, n19795);
  and g31943 (n19797, n_9870, n19795);
  not g31944 (n_12243, n19796);
  not g31945 (n_12244, n19797);
  and g31946 (n19798, n_12243, n_12244);
  not g31947 (n_12245, n19798);
  and g31948 (n19799, \a[11] , n_12245);
  and g31949 (n19800, n_1071, n19798);
  not g31950 (n_12246, n19799);
  not g31951 (n_12247, n19800);
  and g31952 (n19801, n_12246, n_12247);
  not g31953 (n_12248, n19801);
  and g31954 (n19802, n19790, n_12248);
  and g31955 (n19803, n19204, n19396);
  not g31956 (n_12249, n19803);
  and g31957 (n19804, n_11887, n_12249);
  and g31958 (n19805, n7983, n12534);
  and g31959 (n19806, n7291, n12540);
  and g31960 (n19807, n7632, n12537);
  not g31961 (n_12250, n19806);
  not g31962 (n_12251, n19807);
  and g31963 (n19808, n_12250, n_12251);
  not g31964 (n_12252, n19805);
  and g31965 (n19809, n_12252, n19808);
  and g31966 (n19810, n_2446, n19809);
  and g31967 (n19811, n15096, n19809);
  not g31968 (n_12253, n19810);
  not g31969 (n_12254, n19811);
  and g31970 (n19812, n_12253, n_12254);
  not g31971 (n_12255, n19812);
  and g31972 (n19813, \a[11] , n_12255);
  and g31973 (n19814, n_1071, n19812);
  not g31974 (n_12256, n19813);
  not g31975 (n_12257, n19814);
  and g31976 (n19815, n_12256, n_12257);
  not g31977 (n_12258, n19815);
  and g31978 (n19816, n19804, n_12258);
  and g31979 (n19817, n19222, n19394);
  not g31980 (n_12259, n19817);
  and g31981 (n19818, n_11884, n_12259);
  and g31982 (n19819, n7983, n12537);
  and g31983 (n19820, n7291, n12543);
  and g31984 (n19821, n7632, n12540);
  not g31985 (n_12260, n19820);
  not g31986 (n_12261, n19821);
  and g31987 (n19822, n_12260, n_12261);
  not g31988 (n_12262, n19819);
  and g31989 (n19823, n_12262, n19822);
  and g31990 (n19824, n_2446, n19823);
  and g31991 (n19825, n15385, n19823);
  not g31992 (n_12263, n19824);
  not g31993 (n_12264, n19825);
  and g31994 (n19826, n_12263, n_12264);
  not g31995 (n_12265, n19826);
  and g31996 (n19827, \a[11] , n_12265);
  and g31997 (n19828, n_1071, n19826);
  not g31998 (n_12266, n19827);
  not g31999 (n_12267, n19828);
  and g32000 (n19829, n_12266, n_12267);
  not g32001 (n_12268, n19829);
  and g32002 (n19830, n19818, n_12268);
  and g32003 (n19831, n7983, n12540);
  and g32004 (n19832, n7291, n12546);
  and g32005 (n19833, n7632, n12543);
  and g32011 (n19836, n7294, n_8936);
  not g32014 (n_12273, n19837);
  and g32015 (n19838, \a[11] , n_12273);
  not g32016 (n_12274, n19838);
  and g32017 (n19839, n_12273, n_12274);
  and g32018 (n19840, \a[11] , n_12274);
  not g32019 (n_12275, n19839);
  not g32020 (n_12276, n19840);
  and g32021 (n19841, n_12275, n_12276);
  not g32022 (n_12277, n19392);
  and g32023 (n19842, n19390, n_12277);
  not g32024 (n_12278, n19842);
  and g32025 (n19843, n_11881, n_12278);
  not g32026 (n_12279, n19841);
  and g32027 (n19844, n_12279, n19843);
  not g32028 (n_12280, n19844);
  and g32029 (n19845, n_12279, n_12280);
  and g32030 (n19846, n19843, n_12280);
  not g32031 (n_12281, n19845);
  not g32032 (n_12282, n19846);
  and g32033 (n19847, n_12281, n_12282);
  and g32034 (n19848, n7983, n12543);
  and g32035 (n19849, n7291, n12549);
  and g32036 (n19850, n7632, n12546);
  and g32042 (n19853, n7294, n15724);
  not g32045 (n_12287, n19854);
  and g32046 (n19855, \a[11] , n_12287);
  not g32047 (n_12288, n19855);
  and g32048 (n19856, n_12287, n_12288);
  and g32049 (n19857, \a[11] , n_12288);
  not g32050 (n_12289, n19856);
  not g32051 (n_12290, n19857);
  and g32052 (n19858, n_12289, n_12290);
  and g32053 (n19859, n_11874, n_11876);
  and g32054 (n19860, n_11875, n_11876);
  not g32055 (n_12291, n19859);
  not g32056 (n_12292, n19860);
  and g32057 (n19861, n_12291, n_12292);
  not g32058 (n_12293, n19858);
  not g32059 (n_12294, n19861);
  and g32060 (n19862, n_12293, n_12294);
  not g32061 (n_12295, n19862);
  and g32062 (n19863, n_12293, n_12295);
  and g32063 (n19864, n_12294, n_12295);
  not g32064 (n_12296, n19863);
  not g32065 (n_12297, n19864);
  and g32066 (n19865, n_12296, n_12297);
  and g32067 (n19866, n7983, n12546);
  and g32068 (n19867, n7291, n12552);
  and g32069 (n19868, n7632, n12549);
  and g32075 (n19871, n7294, n_8634);
  not g32078 (n_12302, n19872);
  and g32079 (n19873, \a[11] , n_12302);
  not g32080 (n_12303, n19873);
  and g32081 (n19874, n_12302, n_12303);
  and g32082 (n19875, \a[11] , n_12303);
  not g32083 (n_12304, n19874);
  not g32084 (n_12305, n19875);
  and g32085 (n19876, n_12304, n_12305);
  and g32086 (n19877, n_11868, n_11870);
  and g32087 (n19878, n_11869, n_11870);
  not g32088 (n_12306, n19877);
  not g32089 (n_12307, n19878);
  and g32090 (n19879, n_12306, n_12307);
  not g32091 (n_12308, n19876);
  not g32092 (n_12309, n19879);
  and g32093 (n19880, n_12308, n_12309);
  not g32094 (n_12310, n19880);
  and g32095 (n19881, n_12308, n_12310);
  and g32096 (n19882, n_12309, n_12310);
  not g32097 (n_12311, n19881);
  not g32098 (n_12312, n19882);
  and g32099 (n19883, n_12311, n_12312);
  and g32100 (n19884, n19281, n19378);
  not g32101 (n_12313, n19884);
  and g32102 (n19885, n_11864, n_12313);
  and g32103 (n19886, n7983, n12549);
  and g32104 (n19887, n7291, n12555);
  and g32105 (n19888, n7632, n12552);
  not g32106 (n_12314, n19887);
  not g32107 (n_12315, n19888);
  and g32108 (n19889, n_12314, n_12315);
  not g32109 (n_12316, n19886);
  and g32110 (n19890, n_12316, n19889);
  and g32111 (n19891, n_2446, n19890);
  and g32112 (n19892, n_9580, n19890);
  not g32113 (n_12317, n19891);
  not g32114 (n_12318, n19892);
  and g32115 (n19893, n_12317, n_12318);
  not g32116 (n_12319, n19893);
  and g32117 (n19894, \a[11] , n_12319);
  and g32118 (n19895, n_1071, n19893);
  not g32119 (n_12320, n19894);
  not g32120 (n_12321, n19895);
  and g32121 (n19896, n_12320, n_12321);
  not g32122 (n_12322, n19896);
  and g32123 (n19897, n19885, n_12322);
  not g32124 (n_12323, n19376);
  and g32125 (n19898, n19374, n_12323);
  not g32126 (n_12324, n19898);
  and g32127 (n19899, n_11861, n_12324);
  and g32128 (n19900, n7983, n12552);
  and g32129 (n19901, n7291, n12558);
  and g32130 (n19902, n7632, n12555);
  not g32131 (n_12325, n19901);
  not g32132 (n_12326, n19902);
  and g32133 (n19903, n_12325, n_12326);
  not g32134 (n_12327, n19900);
  and g32135 (n19904, n_12327, n19903);
  and g32136 (n19905, n_2446, n19904);
  and g32137 (n19906, n15791, n19904);
  not g32138 (n_12328, n19905);
  not g32139 (n_12329, n19906);
  and g32140 (n19907, n_12328, n_12329);
  not g32141 (n_12330, n19907);
  and g32142 (n19908, \a[11] , n_12330);
  and g32143 (n19909, n_1071, n19907);
  not g32144 (n_12331, n19908);
  not g32145 (n_12332, n19909);
  and g32146 (n19910, n_12331, n_12332);
  not g32147 (n_12333, n19910);
  and g32148 (n19911, n19899, n_12333);
  and g32149 (n19912, n19313, n19372);
  not g32150 (n_12334, n19912);
  and g32151 (n19913, n_11857, n_12334);
  and g32152 (n19914, n7983, n12555);
  and g32153 (n19915, n7291, n12561);
  and g32154 (n19916, n7632, n12558);
  not g32155 (n_12335, n19915);
  not g32156 (n_12336, n19916);
  and g32157 (n19917, n_12335, n_12336);
  not g32158 (n_12337, n19914);
  and g32159 (n19918, n_12337, n19917);
  and g32160 (n19919, n_2446, n19918);
  and g32161 (n19920, n15816, n19918);
  not g32162 (n_12338, n19919);
  not g32163 (n_12339, n19920);
  and g32164 (n19921, n_12338, n_12339);
  not g32165 (n_12340, n19921);
  and g32166 (n19922, \a[11] , n_12340);
  and g32167 (n19923, n_1071, n19921);
  not g32168 (n_12341, n19922);
  not g32169 (n_12342, n19923);
  and g32170 (n19924, n_12341, n_12342);
  not g32171 (n_12343, n19924);
  and g32172 (n19925, n19913, n_12343);
  and g32173 (n19926, n7983, n12558);
  and g32174 (n19927, n7291, n12564);
  and g32175 (n19928, n7632, n12561);
  and g32181 (n19931, n7294, n15847);
  not g32184 (n_12348, n19932);
  and g32185 (n19933, \a[11] , n_12348);
  not g32186 (n_12349, n19933);
  and g32187 (n19934, n_12348, n_12349);
  and g32188 (n19935, \a[11] , n_12349);
  not g32189 (n_12350, n19934);
  not g32190 (n_12351, n19935);
  and g32191 (n19936, n_12350, n_12351);
  not g32192 (n_12352, n19370);
  and g32193 (n19937, n19368, n_12352);
  not g32194 (n_12353, n19937);
  and g32195 (n19938, n_11854, n_12353);
  not g32196 (n_12354, n19936);
  and g32197 (n19939, n_12354, n19938);
  not g32198 (n_12355, n19939);
  and g32199 (n19940, n_12354, n_12355);
  and g32200 (n19941, n19938, n_12355);
  not g32201 (n_12356, n19940);
  not g32202 (n_12357, n19941);
  and g32203 (n19942, n_12356, n_12357);
  and g32204 (n19943, n_11847, n_11849);
  and g32205 (n19944, n_11848, n_11849);
  not g32206 (n_12358, n19943);
  not g32207 (n_12359, n19944);
  and g32208 (n19945, n_12358, n_12359);
  and g32209 (n19946, n7983, n12561);
  and g32210 (n19947, n7291, n12567);
  and g32211 (n19948, n7632, n12564);
  not g32212 (n_12360, n19947);
  not g32213 (n_12361, n19948);
  and g32214 (n19949, n_12360, n_12361);
  not g32215 (n_12362, n19946);
  and g32216 (n19950, n_12362, n19949);
  and g32217 (n19951, n_2446, n19950);
  and g32218 (n19952, n15905, n19950);
  not g32219 (n_12363, n19951);
  not g32220 (n_12364, n19952);
  and g32221 (n19953, n_12363, n_12364);
  not g32222 (n_12365, n19953);
  and g32223 (n19954, \a[11] , n_12365);
  and g32224 (n19955, n_1071, n19953);
  not g32225 (n_12366, n19954);
  not g32226 (n_12367, n19955);
  and g32227 (n19956, n_12366, n_12367);
  not g32228 (n_12368, n19945);
  not g32229 (n_12369, n19956);
  and g32230 (n19957, n_12368, n_12369);
  and g32231 (n19958, n7983, n12564);
  and g32232 (n19959, n7291, n12571);
  and g32233 (n19960, n7632, n12567);
  and g32239 (n19963, n7294, n_9006);
  not g32242 (n_12374, n19964);
  and g32243 (n19965, \a[11] , n_12374);
  not g32244 (n_12375, n19965);
  and g32245 (n19966, n_12374, n_12375);
  and g32246 (n19967, \a[11] , n_12375);
  not g32247 (n_12376, n19966);
  not g32248 (n_12377, n19967);
  and g32249 (n19968, n_12376, n_12377);
  not g32250 (n_12378, n19339);
  and g32251 (n19969, n_12378, n19350);
  not g32252 (n_12379, n19351);
  not g32253 (n_12380, n19969);
  and g32254 (n19970, n_12379, n_12380);
  not g32255 (n_12381, n19968);
  and g32256 (n19971, n_12381, n19970);
  not g32257 (n_12382, n19971);
  and g32258 (n19972, n_12381, n_12382);
  and g32259 (n19973, n19970, n_12382);
  not g32260 (n_12383, n19972);
  not g32261 (n_12384, n19973);
  and g32262 (n19974, n_12383, n_12384);
  not g32263 (n_12385, n19338);
  and g32264 (n19975, n19336, n_12385);
  not g32265 (n_12386, n19975);
  and g32266 (n19976, n_12378, n_12386);
  and g32267 (n19977, n7983, n12567);
  and g32268 (n19978, n7291, n12574);
  and g32269 (n19979, n7632, n12571);
  not g32270 (n_12387, n19978);
  not g32271 (n_12388, n19979);
  and g32272 (n19980, n_12387, n_12388);
  not g32273 (n_12389, n19977);
  and g32274 (n19981, n_12389, n19980);
  and g32275 (n19982, n_2446, n19981);
  and g32276 (n19983, n_10006, n19981);
  not g32277 (n_12390, n19982);
  not g32278 (n_12391, n19983);
  and g32279 (n19984, n_12390, n_12391);
  not g32280 (n_12392, n19984);
  and g32281 (n19985, \a[11] , n_12392);
  and g32282 (n19986, n_1071, n19984);
  not g32283 (n_12393, n19985);
  not g32284 (n_12394, n19986);
  and g32285 (n19987, n_12393, n_12394);
  not g32286 (n_12395, n19987);
  and g32287 (n19988, n19976, n_12395);
  and g32288 (n19989, n7632, n_6977);
  and g32289 (n19990, n7983, n12577);
  not g32290 (n_12396, n19989);
  not g32291 (n_12397, n19990);
  and g32292 (n19991, n_12396, n_12397);
  and g32293 (n19992, n7294, n_9032);
  not g32294 (n_12398, n19992);
  and g32295 (n19993, n19991, n_12398);
  not g32296 (n_12399, n19993);
  and g32297 (n19994, \a[11] , n_12399);
  not g32298 (n_12400, n19994);
  and g32299 (n19995, \a[11] , n_12400);
  and g32300 (n19996, n_12399, n_12400);
  not g32301 (n_12401, n19995);
  not g32302 (n_12402, n19996);
  and g32303 (n19997, n_12401, n_12402);
  and g32304 (n19998, n_2445, n_6977);
  not g32305 (n_12403, n19998);
  and g32306 (n19999, \a[11] , n_12403);
  not g32307 (n_12404, n19997);
  and g32308 (n20000, n_12404, n19999);
  and g32309 (n20001, n7983, n12574);
  and g32310 (n20002, n7291, n_6977);
  and g32311 (n20003, n7632, n12577);
  not g32312 (n_12405, n20002);
  not g32313 (n_12406, n20003);
  and g32314 (n20004, n_12405, n_12406);
  not g32315 (n_12407, n20001);
  and g32316 (n20005, n_12407, n20004);
  and g32317 (n20006, n_2446, n20005);
  and g32318 (n20007, n16094, n20005);
  not g32319 (n_12408, n20006);
  not g32320 (n_12409, n20007);
  and g32321 (n20008, n_12408, n_12409);
  not g32322 (n_12410, n20008);
  and g32323 (n20009, \a[11] , n_12410);
  and g32324 (n20010, n_1071, n20008);
  not g32325 (n_12411, n20009);
  not g32326 (n_12412, n20010);
  and g32327 (n20011, n_12411, n_12412);
  not g32328 (n_12413, n20011);
  and g32329 (n20012, n20000, n_12413);
  and g32330 (n20013, n19337, n20012);
  not g32331 (n_12414, n20013);
  and g32332 (n20014, n20012, n_12414);
  and g32333 (n20015, n19337, n_12414);
  not g32334 (n_12415, n20014);
  not g32335 (n_12416, n20015);
  and g32336 (n20016, n_12415, n_12416);
  and g32337 (n20017, n7983, n12571);
  and g32338 (n20018, n7291, n12577);
  and g32339 (n20019, n7632, n12574);
  and g32345 (n20022, n7294, n16013);
  not g32348 (n_12421, n20023);
  and g32349 (n20024, \a[11] , n_12421);
  not g32350 (n_12422, n20024);
  and g32351 (n20025, \a[11] , n_12422);
  and g32352 (n20026, n_12421, n_12422);
  not g32353 (n_12423, n20025);
  not g32354 (n_12424, n20026);
  and g32355 (n20027, n_12423, n_12424);
  not g32356 (n_12425, n20016);
  not g32357 (n_12426, n20027);
  and g32358 (n20028, n_12425, n_12426);
  not g32359 (n_12427, n20028);
  and g32360 (n20029, n_12414, n_12427);
  not g32361 (n_12428, n19976);
  and g32362 (n20030, n_12428, n19987);
  not g32363 (n_12429, n19988);
  not g32364 (n_12430, n20030);
  and g32365 (n20031, n_12429, n_12430);
  not g32366 (n_12431, n20029);
  and g32367 (n20032, n_12431, n20031);
  not g32368 (n_12432, n20032);
  and g32369 (n20033, n_12429, n_12432);
  not g32370 (n_12433, n19974);
  not g32371 (n_12434, n20033);
  and g32372 (n20034, n_12433, n_12434);
  not g32373 (n_12435, n20034);
  and g32374 (n20035, n_12382, n_12435);
  and g32375 (n20036, n19945, n19956);
  not g32376 (n_12436, n19957);
  not g32377 (n_12437, n20036);
  and g32378 (n20037, n_12436, n_12437);
  not g32379 (n_12438, n20035);
  and g32380 (n20038, n_12438, n20037);
  not g32381 (n_12439, n20038);
  and g32382 (n20039, n_12436, n_12439);
  not g32383 (n_12440, n19942);
  not g32384 (n_12441, n20039);
  and g32385 (n20040, n_12440, n_12441);
  not g32386 (n_12442, n20040);
  and g32387 (n20041, n_12355, n_12442);
  not g32388 (n_12443, n19925);
  and g32389 (n20042, n19913, n_12443);
  and g32390 (n20043, n_12343, n_12443);
  not g32391 (n_12444, n20042);
  not g32392 (n_12445, n20043);
  and g32393 (n20044, n_12444, n_12445);
  not g32394 (n_12446, n20041);
  not g32395 (n_12447, n20044);
  and g32396 (n20045, n_12446, n_12447);
  not g32397 (n_12448, n20045);
  and g32398 (n20046, n_12443, n_12448);
  not g32399 (n_12449, n19911);
  and g32400 (n20047, n19899, n_12449);
  and g32401 (n20048, n_12333, n_12449);
  not g32402 (n_12450, n20047);
  not g32403 (n_12451, n20048);
  and g32404 (n20049, n_12450, n_12451);
  not g32405 (n_12452, n20046);
  not g32406 (n_12453, n20049);
  and g32407 (n20050, n_12452, n_12453);
  not g32408 (n_12454, n20050);
  and g32409 (n20051, n_12449, n_12454);
  not g32410 (n_12455, n19885);
  and g32411 (n20052, n_12455, n19896);
  not g32412 (n_12456, n19897);
  not g32413 (n_12457, n20052);
  and g32414 (n20053, n_12456, n_12457);
  not g32415 (n_12458, n20051);
  and g32416 (n20054, n_12458, n20053);
  not g32417 (n_12459, n20054);
  and g32418 (n20055, n_12456, n_12459);
  not g32419 (n_12460, n19883);
  not g32420 (n_12461, n20055);
  and g32421 (n20056, n_12460, n_12461);
  not g32422 (n_12462, n20056);
  and g32423 (n20057, n_12310, n_12462);
  not g32424 (n_12463, n19865);
  not g32425 (n_12464, n20057);
  and g32426 (n20058, n_12463, n_12464);
  not g32427 (n_12465, n20058);
  and g32428 (n20059, n_12295, n_12465);
  not g32429 (n_12466, n19847);
  not g32430 (n_12467, n20059);
  and g32431 (n20060, n_12466, n_12467);
  not g32432 (n_12468, n20060);
  and g32433 (n20061, n_12280, n_12468);
  not g32434 (n_12469, n19830);
  and g32435 (n20062, n19818, n_12469);
  and g32436 (n20063, n_12268, n_12469);
  not g32437 (n_12470, n20062);
  not g32438 (n_12471, n20063);
  and g32439 (n20064, n_12470, n_12471);
  not g32440 (n_12472, n20061);
  not g32441 (n_12473, n20064);
  and g32442 (n20065, n_12472, n_12473);
  not g32443 (n_12474, n20065);
  and g32444 (n20066, n_12469, n_12474);
  not g32445 (n_12475, n19816);
  and g32446 (n20067, n19804, n_12475);
  and g32447 (n20068, n_12258, n_12475);
  not g32448 (n_12476, n20067);
  not g32449 (n_12477, n20068);
  and g32450 (n20069, n_12476, n_12477);
  not g32451 (n_12478, n20066);
  not g32452 (n_12479, n20069);
  and g32453 (n20070, n_12478, n_12479);
  not g32454 (n_12480, n20070);
  and g32455 (n20071, n_12475, n_12480);
  not g32456 (n_12481, n19790);
  and g32457 (n20072, n_12481, n19801);
  not g32458 (n_12482, n19802);
  not g32459 (n_12483, n20072);
  and g32460 (n20073, n_12482, n_12483);
  not g32461 (n_12484, n20071);
  and g32462 (n20074, n_12484, n20073);
  not g32463 (n_12485, n20074);
  and g32464 (n20075, n_12482, n_12485);
  not g32465 (n_12486, n19788);
  not g32466 (n_12487, n20075);
  and g32467 (n20076, n_12486, n_12487);
  not g32468 (n_12488, n20076);
  and g32469 (n20077, n_12236, n_12488);
  not g32470 (n_12489, n19770);
  not g32471 (n_12490, n20077);
  and g32472 (n20078, n_12489, n_12490);
  not g32473 (n_12491, n20078);
  and g32474 (n20079, n_12221, n_12491);
  not g32475 (n_12492, n19752);
  not g32476 (n_12493, n20079);
  and g32477 (n20080, n_12492, n_12493);
  not g32478 (n_12494, n20080);
  and g32479 (n20081, n_12206, n_12494);
  not g32480 (n_12495, n19735);
  and g32481 (n20082, n19723, n_12495);
  and g32482 (n20083, n_12194, n_12495);
  not g32483 (n_12496, n20082);
  not g32484 (n_12497, n20083);
  and g32485 (n20084, n_12496, n_12497);
  not g32486 (n_12498, n20081);
  not g32487 (n_12499, n20084);
  and g32488 (n20085, n_12498, n_12499);
  not g32489 (n_12500, n20085);
  and g32490 (n20086, n_12495, n_12500);
  not g32491 (n_12501, n19709);
  and g32492 (n20087, n_12501, n19720);
  not g32493 (n_12502, n19721);
  not g32494 (n_12503, n20087);
  and g32495 (n20088, n_12502, n_12503);
  not g32496 (n_12504, n20086);
  and g32497 (n20089, n_12504, n20088);
  not g32498 (n_12505, n20089);
  and g32499 (n20090, n_12502, n_12505);
  not g32500 (n_12506, n19707);
  not g32501 (n_12507, n20090);
  and g32502 (n20091, n_12506, n_12507);
  not g32503 (n_12508, n20091);
  and g32504 (n20092, n_12172, n_12508);
  not g32505 (n_12509, n19689);
  not g32506 (n_12510, n20092);
  and g32507 (n20093, n_12509, n_12510);
  not g32508 (n_12511, n20093);
  and g32509 (n20094, n_12157, n_12511);
  not g32510 (n_12512, n19671);
  not g32511 (n_12513, n20094);
  and g32512 (n20095, n_12512, n_12513);
  not g32513 (n_12514, n20095);
  and g32514 (n20096, n_12142, n_12514);
  not g32515 (n_12515, n19653);
  not g32516 (n_12516, n20096);
  and g32517 (n20097, n_12515, n_12516);
  not g32518 (n_12517, n20097);
  and g32519 (n20098, n_12127, n_12517);
  not g32520 (n_12518, n19635);
  not g32521 (n_12519, n20098);
  and g32522 (n20099, n_12518, n_12519);
  not g32523 (n_12520, n20099);
  and g32524 (n20100, n_12112, n_12520);
  not g32525 (n_12521, n19617);
  not g32526 (n_12522, n20100);
  and g32527 (n20101, n_12521, n_12522);
  not g32528 (n_12523, n20101);
  and g32529 (n20102, n_12097, n_12523);
  not g32530 (n_12524, n19599);
  not g32531 (n_12525, n20102);
  and g32532 (n20103, n_12524, n_12525);
  not g32533 (n_12526, n20103);
  and g32534 (n20104, n_12082, n_12526);
  not g32535 (n_12527, n19581);
  not g32536 (n_12528, n20104);
  and g32537 (n20105, n_12527, n_12528);
  not g32538 (n_12529, n20105);
  and g32539 (n20106, n_12067, n_12529);
  not g32540 (n_12530, n19563);
  not g32541 (n_12531, n20106);
  and g32542 (n20107, n_12530, n_12531);
  not g32543 (n_12532, n20107);
  and g32544 (n20108, n_12052, n_12532);
  not g32545 (n_12533, n19545);
  not g32546 (n_12534, n20108);
  and g32547 (n20109, n_12533, n_12534);
  not g32548 (n_12535, n20109);
  and g32549 (n20110, n_12037, n_12535);
  not g32550 (n_12536, n19528);
  not g32551 (n_12537, n20110);
  and g32552 (n20111, n_12536, n_12537);
  and g32553 (n20112, n19528, n20110);
  not g32554 (n_12538, n20111);
  not g32555 (n_12539, n20112);
  and g32556 (n20113, n_12538, n_12539);
  and g32557 (n20114, n9331, n13630);
  and g32558 (n20115, n8418, n13515);
  and g32559 (n20116, n8860, n13597);
  and g32565 (n20119, n8421, n13976);
  not g32568 (n_12544, n20120);
  and g32569 (n20121, \a[8] , n_12544);
  not g32570 (n_12545, n20121);
  and g32571 (n20122, \a[8] , n_12545);
  and g32572 (n20123, n_12544, n_12545);
  not g32573 (n_12546, n20122);
  not g32574 (n_12547, n20123);
  and g32575 (n20124, n_12546, n_12547);
  not g32576 (n_12548, n20124);
  and g32577 (n20125, n20113, n_12548);
  not g32578 (n_12549, n20125);
  and g32579 (n20126, n_12538, n_12549);
  not g32580 (n_12550, n19525);
  not g32581 (n_12551, n20126);
  and g32582 (n20127, n_12550, n_12551);
  and g32583 (n20128, n19525, n20126);
  not g32584 (n_12552, n20127);
  not g32585 (n_12553, n20128);
  and g32586 (n20129, n_12552, n_12553);
  and g32587 (n20130, n71, n_7417);
  and g32588 (n20131, n9867, n_7540);
  and g32589 (n20132, n10434, n13941);
  and g32595 (n20135, n9870, n14028);
  not g32598 (n_12558, n20136);
  and g32599 (n20137, \a[5] , n_12558);
  not g32600 (n_12559, n20137);
  and g32601 (n20138, \a[5] , n_12559);
  and g32602 (n20139, n_12558, n_12559);
  not g32603 (n_12560, n20138);
  not g32604 (n_12561, n20139);
  and g32605 (n20140, n_12560, n_12561);
  not g32606 (n_12562, n20140);
  and g32607 (n20141, n20129, n_12562);
  not g32608 (n_12563, n20141);
  and g32609 (n20142, n_12552, n_12563);
  not g32610 (n_12564, n19522);
  not g32611 (n_12565, n20142);
  and g32612 (n20143, n_12564, n_12565);
  and g32613 (n20144, n19522, n20142);
  not g32614 (n_12566, n20143);
  not g32615 (n_12567, n20144);
  and g32616 (n20145, n_12566, n_12567);
  and g32617 (n20146, n20129, n_12563);
  and g32618 (n20147, n_12562, n_12563);
  not g32619 (n_12568, n20146);
  not g32620 (n_12569, n20147);
  and g32621 (n20148, n_12568, n_12569);
  and g32622 (n20149, n20113, n_12549);
  and g32623 (n20150, n_12548, n_12549);
  not g32624 (n_12570, n20149);
  not g32625 (n_12571, n20150);
  and g32626 (n20151, n_12570, n_12571);
  and g32627 (n20152, n19545, n20108);
  not g32628 (n_12572, n20152);
  and g32629 (n20153, n_12535, n_12572);
  and g32630 (n20154, n9331, n13597);
  and g32631 (n20155, n8418, n13521);
  and g32632 (n20156, n8860, n13515);
  not g32633 (n_12573, n20155);
  not g32634 (n_12574, n20156);
  and g32635 (n20157, n_12573, n_12574);
  not g32636 (n_12575, n20154);
  and g32637 (n20158, n_12575, n20157);
  and g32638 (n20159, n_3428, n20158);
  and g32639 (n20160, n13612, n20158);
  not g32640 (n_12576, n20159);
  not g32641 (n_12577, n20160);
  and g32642 (n20161, n_12576, n_12577);
  not g32643 (n_12578, n20161);
  and g32644 (n20162, \a[8] , n_12578);
  and g32645 (n20163, n_1106, n20161);
  not g32646 (n_12579, n20162);
  not g32647 (n_12580, n20163);
  and g32648 (n20164, n_12579, n_12580);
  not g32649 (n_12581, n20164);
  and g32650 (n20165, n20153, n_12581);
  and g32651 (n20166, n19563, n20106);
  not g32652 (n_12582, n20166);
  and g32653 (n20167, n_12532, n_12582);
  and g32654 (n20168, n9331, n13515);
  and g32655 (n20169, n8418, n13518);
  and g32656 (n20170, n8860, n13521);
  not g32657 (n_12583, n20169);
  not g32658 (n_12584, n20170);
  and g32659 (n20171, n_12583, n_12584);
  not g32660 (n_12585, n20168);
  and g32661 (n20172, n_12585, n20171);
  and g32662 (n20173, n_3428, n20172);
  and g32663 (n20174, n_7486, n20172);
  not g32664 (n_12586, n20173);
  not g32665 (n_12587, n20174);
  and g32666 (n20175, n_12586, n_12587);
  not g32667 (n_12588, n20175);
  and g32668 (n20176, \a[8] , n_12588);
  and g32669 (n20177, n_1106, n20175);
  not g32670 (n_12589, n20176);
  not g32671 (n_12590, n20177);
  and g32672 (n20178, n_12589, n_12590);
  not g32673 (n_12591, n20178);
  and g32674 (n20179, n20167, n_12591);
  and g32675 (n20180, n19581, n20104);
  not g32676 (n_12592, n20180);
  and g32677 (n20181, n_12529, n_12592);
  and g32678 (n20182, n9331, n13521);
  and g32679 (n20183, n8418, n13491);
  and g32680 (n20184, n8860, n13518);
  not g32681 (n_12593, n20183);
  not g32682 (n_12594, n20184);
  and g32683 (n20185, n_12593, n_12594);
  not g32684 (n_12595, n20182);
  and g32685 (n20186, n_12595, n20185);
  and g32686 (n20187, n_3428, n20186);
  and g32687 (n20188, n13909, n20186);
  not g32688 (n_12596, n20187);
  not g32689 (n_12597, n20188);
  and g32690 (n20189, n_12596, n_12597);
  not g32691 (n_12598, n20189);
  and g32692 (n20190, \a[8] , n_12598);
  and g32693 (n20191, n_1106, n20189);
  not g32694 (n_12599, n20190);
  not g32695 (n_12600, n20191);
  and g32696 (n20192, n_12599, n_12600);
  not g32697 (n_12601, n20192);
  and g32698 (n20193, n20181, n_12601);
  and g32699 (n20194, n19599, n20102);
  not g32700 (n_12602, n20194);
  and g32701 (n20195, n_12526, n_12602);
  and g32702 (n20196, n9331, n13518);
  and g32703 (n20197, n8418, n12889);
  and g32704 (n20198, n8860, n13491);
  not g32705 (n_12603, n20197);
  not g32706 (n_12604, n20198);
  and g32707 (n20199, n_12603, n_12604);
  not g32708 (n_12605, n20196);
  and g32709 (n20200, n_12605, n20199);
  and g32710 (n20201, n_3428, n20200);
  not g32711 (n_12606, n13584);
  and g32712 (n20202, n_12606, n20200);
  not g32713 (n_12607, n20201);
  not g32714 (n_12608, n20202);
  and g32715 (n20203, n_12607, n_12608);
  not g32716 (n_12609, n20203);
  and g32717 (n20204, \a[8] , n_12609);
  and g32718 (n20205, n_1106, n20203);
  not g32719 (n_12610, n20204);
  not g32720 (n_12611, n20205);
  and g32721 (n20206, n_12610, n_12611);
  not g32722 (n_12612, n20206);
  and g32723 (n20207, n20195, n_12612);
  and g32724 (n20208, n19617, n20100);
  not g32725 (n_12613, n20208);
  and g32726 (n20209, n_12523, n_12613);
  and g32727 (n20210, n9331, n13491);
  and g32728 (n20211, n8418, n12769);
  and g32729 (n20212, n8860, n12889);
  not g32730 (n_12614, n20211);
  not g32731 (n_12615, n20212);
  and g32732 (n20213, n_12614, n_12615);
  not g32733 (n_12616, n20210);
  and g32734 (n20214, n_12616, n20213);
  and g32735 (n20215, n_3428, n20214);
  and g32736 (n20216, n13503, n20214);
  not g32737 (n_12617, n20215);
  not g32738 (n_12618, n20216);
  and g32739 (n20217, n_12617, n_12618);
  not g32740 (n_12619, n20217);
  and g32741 (n20218, \a[8] , n_12619);
  and g32742 (n20219, n_1106, n20217);
  not g32743 (n_12620, n20218);
  not g32744 (n_12621, n20219);
  and g32745 (n20220, n_12620, n_12621);
  not g32746 (n_12622, n20220);
  and g32747 (n20221, n20209, n_12622);
  and g32748 (n20222, n19635, n20098);
  not g32749 (n_12623, n20222);
  and g32750 (n20223, n_12520, n_12623);
  and g32751 (n20224, n9331, n12889);
  and g32752 (n20225, n8418, n12502);
  and g32753 (n20226, n8860, n12769);
  not g32754 (n_12624, n20225);
  not g32755 (n_12625, n20226);
  and g32756 (n20227, n_12624, n_12625);
  not g32757 (n_12626, n20224);
  and g32758 (n20228, n_12626, n20227);
  and g32759 (n20229, n_3428, n20228);
  not g32760 (n_12627, n12895);
  and g32761 (n20230, n_12627, n20228);
  not g32762 (n_12628, n20229);
  not g32763 (n_12629, n20230);
  and g32764 (n20231, n_12628, n_12629);
  not g32765 (n_12630, n20231);
  and g32766 (n20232, \a[8] , n_12630);
  and g32767 (n20233, n_1106, n20231);
  not g32768 (n_12631, n20232);
  not g32769 (n_12632, n20233);
  and g32770 (n20234, n_12631, n_12632);
  not g32771 (n_12633, n20234);
  and g32772 (n20235, n20223, n_12633);
  and g32773 (n20236, n19653, n20096);
  not g32774 (n_12634, n20236);
  and g32775 (n20237, n_12517, n_12634);
  and g32776 (n20238, n9331, n12769);
  and g32777 (n20239, n8418, n12370);
  and g32778 (n20240, n8860, n12502);
  not g32779 (n_12635, n20239);
  not g32780 (n_12636, n20240);
  and g32781 (n20241, n_12635, n_12636);
  not g32782 (n_12637, n20238);
  and g32783 (n20242, n_12637, n20241);
  and g32784 (n20243, n_3428, n20242);
  and g32785 (n20244, n_7817, n20242);
  not g32786 (n_12638, n20243);
  not g32787 (n_12639, n20244);
  and g32788 (n20245, n_12638, n_12639);
  not g32789 (n_12640, n20245);
  and g32790 (n20246, \a[8] , n_12640);
  and g32791 (n20247, n_1106, n20245);
  not g32792 (n_12641, n20246);
  not g32793 (n_12642, n20247);
  and g32794 (n20248, n_12641, n_12642);
  not g32795 (n_12643, n20248);
  and g32796 (n20249, n20237, n_12643);
  and g32797 (n20250, n19671, n20094);
  not g32798 (n_12644, n20250);
  and g32799 (n20251, n_12514, n_12644);
  and g32800 (n20252, n9331, n12502);
  and g32801 (n20253, n8418, n12505);
  and g32802 (n20254, n8860, n12370);
  not g32803 (n_12645, n20253);
  not g32804 (n_12646, n20254);
  and g32805 (n20255, n_12645, n_12646);
  not g32806 (n_12647, n20252);
  and g32807 (n20256, n_12647, n20255);
  and g32808 (n20257, n_3428, n20256);
  and g32809 (n20258, n13736, n20256);
  not g32810 (n_12648, n20257);
  not g32811 (n_12649, n20258);
  and g32812 (n20259, n_12648, n_12649);
  not g32813 (n_12650, n20259);
  and g32814 (n20260, \a[8] , n_12650);
  and g32815 (n20261, n_1106, n20259);
  not g32816 (n_12651, n20260);
  not g32817 (n_12652, n20261);
  and g32818 (n20262, n_12651, n_12652);
  not g32819 (n_12653, n20262);
  and g32820 (n20263, n20251, n_12653);
  and g32821 (n20264, n19689, n20092);
  not g32822 (n_12654, n20264);
  and g32823 (n20265, n_12511, n_12654);
  and g32824 (n20266, n9331, n12370);
  and g32825 (n20267, n8418, n12508);
  and g32826 (n20268, n8860, n12505);
  not g32827 (n_12655, n20267);
  not g32828 (n_12656, n20268);
  and g32829 (n20269, n_12655, n_12656);
  not g32830 (n_12657, n20266);
  and g32831 (n20270, n_12657, n20269);
  and g32832 (n20271, n_3428, n20270);
  and g32833 (n20272, n13748, n20270);
  not g32834 (n_12658, n20271);
  not g32835 (n_12659, n20272);
  and g32836 (n20273, n_12658, n_12659);
  not g32837 (n_12660, n20273);
  and g32838 (n20274, \a[8] , n_12660);
  and g32839 (n20275, n_1106, n20273);
  not g32840 (n_12661, n20274);
  not g32841 (n_12662, n20275);
  and g32842 (n20276, n_12661, n_12662);
  not g32843 (n_12663, n20276);
  and g32844 (n20277, n20265, n_12663);
  and g32845 (n20278, n19707, n20090);
  not g32846 (n_12664, n20278);
  and g32847 (n20279, n_12508, n_12664);
  and g32848 (n20280, n9331, n12505);
  and g32849 (n20281, n8418, n12513);
  and g32850 (n20282, n8860, n12508);
  not g32851 (n_12665, n20281);
  not g32852 (n_12666, n20282);
  and g32853 (n20283, n_12665, n_12666);
  not g32854 (n_12667, n20280);
  and g32855 (n20284, n_12667, n20283);
  and g32856 (n20285, n_3428, n20284);
  and g32857 (n20286, n14051, n20284);
  not g32858 (n_12668, n20285);
  not g32859 (n_12669, n20286);
  and g32860 (n20287, n_12668, n_12669);
  not g32861 (n_12670, n20287);
  and g32862 (n20288, \a[8] , n_12670);
  and g32863 (n20289, n_1106, n20287);
  not g32864 (n_12671, n20288);
  not g32865 (n_12672, n20289);
  and g32866 (n20290, n_12671, n_12672);
  not g32867 (n_12673, n20290);
  and g32868 (n20291, n20279, n_12673);
  and g32869 (n20292, n9331, n12508);
  and g32870 (n20293, n8418, n12511);
  and g32871 (n20294, n8860, n12513);
  and g32877 (n20297, n8421, n13863);
  not g32880 (n_12678, n20298);
  and g32881 (n20299, \a[8] , n_12678);
  not g32882 (n_12679, n20299);
  and g32883 (n20300, n_12678, n_12679);
  and g32884 (n20301, \a[8] , n_12679);
  not g32885 (n_12680, n20300);
  not g32886 (n_12681, n20301);
  and g32887 (n20302, n_12680, n_12681);
  not g32888 (n_12682, n20088);
  and g32889 (n20303, n20086, n_12682);
  not g32890 (n_12683, n20303);
  and g32891 (n20304, n_12505, n_12683);
  not g32892 (n_12684, n20302);
  and g32893 (n20305, n_12684, n20304);
  not g32894 (n_12685, n20305);
  and g32895 (n20306, n_12684, n_12685);
  and g32896 (n20307, n20304, n_12685);
  not g32897 (n_12686, n20306);
  not g32898 (n_12687, n20307);
  and g32899 (n20308, n_12686, n_12687);
  and g32900 (n20309, n9331, n12513);
  and g32901 (n20310, n8418, n12516);
  and g32902 (n20311, n8860, n12511);
  and g32908 (n20314, n8421, n14177);
  not g32911 (n_12692, n20315);
  and g32912 (n20316, \a[8] , n_12692);
  not g32913 (n_12693, n20316);
  and g32914 (n20317, n_12692, n_12693);
  and g32915 (n20318, \a[8] , n_12693);
  not g32916 (n_12694, n20317);
  not g32917 (n_12695, n20318);
  and g32918 (n20319, n_12694, n_12695);
  and g32919 (n20320, n_12498, n_12500);
  and g32920 (n20321, n_12499, n_12500);
  not g32921 (n_12696, n20320);
  not g32922 (n_12697, n20321);
  and g32923 (n20322, n_12696, n_12697);
  not g32924 (n_12698, n20319);
  not g32925 (n_12699, n20322);
  and g32926 (n20323, n_12698, n_12699);
  not g32927 (n_12700, n20323);
  and g32928 (n20324, n_12698, n_12700);
  and g32929 (n20325, n_12699, n_12700);
  not g32930 (n_12701, n20324);
  not g32931 (n_12702, n20325);
  and g32932 (n20326, n_12701, n_12702);
  and g32933 (n20327, n19752, n20079);
  not g32934 (n_12703, n20327);
  and g32935 (n20328, n_12494, n_12703);
  and g32936 (n20329, n9331, n12511);
  and g32937 (n20330, n8418, n12519);
  and g32938 (n20331, n8860, n12516);
  not g32939 (n_12704, n20330);
  not g32940 (n_12705, n20331);
  and g32941 (n20332, n_12704, n_12705);
  not g32942 (n_12706, n20329);
  and g32943 (n20333, n_12706, n20332);
  and g32944 (n20334, n_3428, n20333);
  and g32945 (n20335, n14233, n20333);
  not g32946 (n_12707, n20334);
  not g32947 (n_12708, n20335);
  and g32948 (n20336, n_12707, n_12708);
  not g32949 (n_12709, n20336);
  and g32950 (n20337, \a[8] , n_12709);
  and g32951 (n20338, n_1106, n20336);
  not g32952 (n_12710, n20337);
  not g32953 (n_12711, n20338);
  and g32954 (n20339, n_12710, n_12711);
  not g32955 (n_12712, n20339);
  and g32956 (n20340, n20328, n_12712);
  and g32957 (n20341, n19770, n20077);
  not g32958 (n_12713, n20341);
  and g32959 (n20342, n_12491, n_12713);
  and g32960 (n20343, n9331, n12516);
  and g32961 (n20344, n8418, n12522);
  and g32962 (n20345, n8860, n12519);
  not g32963 (n_12714, n20344);
  not g32964 (n_12715, n20345);
  and g32965 (n20346, n_12714, n_12715);
  not g32966 (n_12716, n20343);
  and g32967 (n20347, n_12716, n20346);
  and g32968 (n20348, n_3428, n20347);
  and g32969 (n20349, n14443, n20347);
  not g32970 (n_12717, n20348);
  not g32971 (n_12718, n20349);
  and g32972 (n20350, n_12717, n_12718);
  not g32973 (n_12719, n20350);
  and g32974 (n20351, \a[8] , n_12719);
  and g32975 (n20352, n_1106, n20350);
  not g32976 (n_12720, n20351);
  not g32977 (n_12721, n20352);
  and g32978 (n20353, n_12720, n_12721);
  not g32979 (n_12722, n20353);
  and g32980 (n20354, n20342, n_12722);
  and g32981 (n20355, n19788, n20075);
  not g32982 (n_12723, n20355);
  and g32983 (n20356, n_12488, n_12723);
  and g32984 (n20357, n9331, n12519);
  and g32985 (n20358, n8418, n12525);
  and g32986 (n20359, n8860, n12522);
  not g32987 (n_12724, n20358);
  not g32988 (n_12725, n20359);
  and g32989 (n20360, n_12724, n_12725);
  not g32990 (n_12726, n20357);
  and g32991 (n20361, n_12726, n20360);
  and g32992 (n20362, n_3428, n20361);
  and g32993 (n20363, n_10664, n20361);
  not g32994 (n_12727, n20362);
  not g32995 (n_12728, n20363);
  and g32996 (n20364, n_12727, n_12728);
  not g32997 (n_12729, n20364);
  and g32998 (n20365, \a[8] , n_12729);
  and g32999 (n20366, n_1106, n20364);
  not g33000 (n_12730, n20365);
  not g33001 (n_12731, n20366);
  and g33002 (n20367, n_12730, n_12731);
  not g33003 (n_12732, n20367);
  and g33004 (n20368, n20356, n_12732);
  and g33005 (n20369, n9331, n12522);
  and g33006 (n20370, n8418, n12528);
  and g33007 (n20371, n8860, n12525);
  and g33013 (n20374, n8421, n14837);
  not g33016 (n_12737, n20375);
  and g33017 (n20376, \a[8] , n_12737);
  not g33018 (n_12738, n20376);
  and g33019 (n20377, n_12737, n_12738);
  and g33020 (n20378, \a[8] , n_12738);
  not g33021 (n_12739, n20377);
  not g33022 (n_12740, n20378);
  and g33023 (n20379, n_12739, n_12740);
  not g33024 (n_12741, n20073);
  and g33025 (n20380, n20071, n_12741);
  not g33026 (n_12742, n20380);
  and g33027 (n20381, n_12485, n_12742);
  not g33028 (n_12743, n20379);
  and g33029 (n20382, n_12743, n20381);
  not g33030 (n_12744, n20382);
  and g33031 (n20383, n_12743, n_12744);
  and g33032 (n20384, n20381, n_12744);
  not g33033 (n_12745, n20383);
  not g33034 (n_12746, n20384);
  and g33035 (n20385, n_12745, n_12746);
  and g33036 (n20386, n9331, n12525);
  and g33037 (n20387, n8418, n12531);
  and g33038 (n20388, n8860, n12528);
  and g33044 (n20391, n8421, n14608);
  not g33047 (n_12751, n20392);
  and g33048 (n20393, \a[8] , n_12751);
  not g33049 (n_12752, n20393);
  and g33050 (n20394, n_12751, n_12752);
  and g33051 (n20395, \a[8] , n_12752);
  not g33052 (n_12753, n20394);
  not g33053 (n_12754, n20395);
  and g33054 (n20396, n_12753, n_12754);
  and g33055 (n20397, n_12478, n_12480);
  and g33056 (n20398, n_12479, n_12480);
  not g33057 (n_12755, n20397);
  not g33058 (n_12756, n20398);
  and g33059 (n20399, n_12755, n_12756);
  not g33060 (n_12757, n20396);
  not g33061 (n_12758, n20399);
  and g33062 (n20400, n_12757, n_12758);
  not g33063 (n_12759, n20400);
  and g33064 (n20401, n_12757, n_12759);
  and g33065 (n20402, n_12758, n_12759);
  not g33066 (n_12760, n20401);
  not g33067 (n_12761, n20402);
  and g33068 (n20403, n_12760, n_12761);
  and g33069 (n20404, n9331, n12528);
  and g33070 (n20405, n8418, n12534);
  and g33071 (n20406, n8860, n12531);
  and g33077 (n20409, n8421, n_8448);
  not g33080 (n_12766, n20410);
  and g33081 (n20411, \a[8] , n_12766);
  not g33082 (n_12767, n20411);
  and g33083 (n20412, n_12766, n_12767);
  and g33084 (n20413, \a[8] , n_12767);
  not g33085 (n_12768, n20412);
  not g33086 (n_12769, n20413);
  and g33087 (n20414, n_12768, n_12769);
  and g33088 (n20415, n_12472, n_12474);
  and g33089 (n20416, n_12473, n_12474);
  not g33090 (n_12770, n20415);
  not g33091 (n_12771, n20416);
  and g33092 (n20417, n_12770, n_12771);
  not g33093 (n_12772, n20414);
  not g33094 (n_12773, n20417);
  and g33095 (n20418, n_12772, n_12773);
  not g33096 (n_12774, n20418);
  and g33097 (n20419, n_12772, n_12774);
  and g33098 (n20420, n_12773, n_12774);
  not g33099 (n_12775, n20419);
  not g33100 (n_12776, n20420);
  and g33101 (n20421, n_12775, n_12776);
  and g33102 (n20422, n19847, n20059);
  not g33103 (n_12777, n20422);
  and g33104 (n20423, n_12468, n_12777);
  and g33105 (n20424, n9331, n12531);
  and g33106 (n20425, n8418, n12537);
  and g33107 (n20426, n8860, n12534);
  not g33108 (n_12778, n20425);
  not g33109 (n_12779, n20426);
  and g33110 (n20427, n_12778, n_12779);
  not g33111 (n_12780, n20424);
  and g33112 (n20428, n_12780, n20427);
  and g33113 (n20429, n_3428, n20428);
  and g33114 (n20430, n_9870, n20428);
  not g33115 (n_12781, n20429);
  not g33116 (n_12782, n20430);
  and g33117 (n20431, n_12781, n_12782);
  not g33118 (n_12783, n20431);
  and g33119 (n20432, \a[8] , n_12783);
  and g33120 (n20433, n_1106, n20431);
  not g33121 (n_12784, n20432);
  not g33122 (n_12785, n20433);
  and g33123 (n20434, n_12784, n_12785);
  not g33124 (n_12786, n20434);
  and g33125 (n20435, n20423, n_12786);
  and g33126 (n20436, n19865, n20057);
  not g33127 (n_12787, n20436);
  and g33128 (n20437, n_12465, n_12787);
  and g33129 (n20438, n9331, n12534);
  and g33130 (n20439, n8418, n12540);
  and g33131 (n20440, n8860, n12537);
  not g33132 (n_12788, n20439);
  not g33133 (n_12789, n20440);
  and g33134 (n20441, n_12788, n_12789);
  not g33135 (n_12790, n20438);
  and g33136 (n20442, n_12790, n20441);
  and g33137 (n20443, n_3428, n20442);
  and g33138 (n20444, n15096, n20442);
  not g33139 (n_12791, n20443);
  not g33140 (n_12792, n20444);
  and g33141 (n20445, n_12791, n_12792);
  not g33142 (n_12793, n20445);
  and g33143 (n20446, \a[8] , n_12793);
  and g33144 (n20447, n_1106, n20445);
  not g33145 (n_12794, n20446);
  not g33146 (n_12795, n20447);
  and g33147 (n20448, n_12794, n_12795);
  not g33148 (n_12796, n20448);
  and g33149 (n20449, n20437, n_12796);
  and g33150 (n20450, n19883, n20055);
  not g33151 (n_12797, n20450);
  and g33152 (n20451, n_12462, n_12797);
  and g33153 (n20452, n9331, n12537);
  and g33154 (n20453, n8418, n12543);
  and g33155 (n20454, n8860, n12540);
  not g33156 (n_12798, n20453);
  not g33157 (n_12799, n20454);
  and g33158 (n20455, n_12798, n_12799);
  not g33159 (n_12800, n20452);
  and g33160 (n20456, n_12800, n20455);
  and g33161 (n20457, n_3428, n20456);
  and g33162 (n20458, n15385, n20456);
  not g33163 (n_12801, n20457);
  not g33164 (n_12802, n20458);
  and g33165 (n20459, n_12801, n_12802);
  not g33166 (n_12803, n20459);
  and g33167 (n20460, \a[8] , n_12803);
  and g33168 (n20461, n_1106, n20459);
  not g33169 (n_12804, n20460);
  not g33170 (n_12805, n20461);
  and g33171 (n20462, n_12804, n_12805);
  not g33172 (n_12806, n20462);
  and g33173 (n20463, n20451, n_12806);
  and g33174 (n20464, n9331, n12540);
  and g33175 (n20465, n8418, n12546);
  and g33176 (n20466, n8860, n12543);
  and g33182 (n20469, n8421, n_8936);
  not g33185 (n_12811, n20470);
  and g33186 (n20471, \a[8] , n_12811);
  not g33187 (n_12812, n20471);
  and g33188 (n20472, n_12811, n_12812);
  and g33189 (n20473, \a[8] , n_12812);
  not g33190 (n_12813, n20472);
  not g33191 (n_12814, n20473);
  and g33192 (n20474, n_12813, n_12814);
  not g33193 (n_12815, n20053);
  and g33194 (n20475, n20051, n_12815);
  not g33195 (n_12816, n20475);
  and g33196 (n20476, n_12459, n_12816);
  not g33197 (n_12817, n20474);
  and g33198 (n20477, n_12817, n20476);
  not g33199 (n_12818, n20477);
  and g33200 (n20478, n_12817, n_12818);
  and g33201 (n20479, n20476, n_12818);
  not g33202 (n_12819, n20478);
  not g33203 (n_12820, n20479);
  and g33204 (n20480, n_12819, n_12820);
  and g33205 (n20481, n9331, n12543);
  and g33206 (n20482, n8418, n12549);
  and g33207 (n20483, n8860, n12546);
  and g33213 (n20486, n8421, n15724);
  not g33216 (n_12825, n20487);
  and g33217 (n20488, \a[8] , n_12825);
  not g33218 (n_12826, n20488);
  and g33219 (n20489, n_12825, n_12826);
  and g33220 (n20490, \a[8] , n_12826);
  not g33221 (n_12827, n20489);
  not g33222 (n_12828, n20490);
  and g33223 (n20491, n_12827, n_12828);
  and g33224 (n20492, n_12452, n_12454);
  and g33225 (n20493, n_12453, n_12454);
  not g33226 (n_12829, n20492);
  not g33227 (n_12830, n20493);
  and g33228 (n20494, n_12829, n_12830);
  not g33229 (n_12831, n20491);
  not g33230 (n_12832, n20494);
  and g33231 (n20495, n_12831, n_12832);
  not g33232 (n_12833, n20495);
  and g33233 (n20496, n_12831, n_12833);
  and g33234 (n20497, n_12832, n_12833);
  not g33235 (n_12834, n20496);
  not g33236 (n_12835, n20497);
  and g33237 (n20498, n_12834, n_12835);
  and g33238 (n20499, n9331, n12546);
  and g33239 (n20500, n8418, n12552);
  and g33240 (n20501, n8860, n12549);
  and g33246 (n20504, n8421, n_8634);
  not g33249 (n_12840, n20505);
  and g33250 (n20506, \a[8] , n_12840);
  not g33251 (n_12841, n20506);
  and g33252 (n20507, n_12840, n_12841);
  and g33253 (n20508, \a[8] , n_12841);
  not g33254 (n_12842, n20507);
  not g33255 (n_12843, n20508);
  and g33256 (n20509, n_12842, n_12843);
  and g33257 (n20510, n_12446, n_12448);
  and g33258 (n20511, n_12447, n_12448);
  not g33259 (n_12844, n20510);
  not g33260 (n_12845, n20511);
  and g33261 (n20512, n_12844, n_12845);
  not g33262 (n_12846, n20509);
  not g33263 (n_12847, n20512);
  and g33264 (n20513, n_12846, n_12847);
  not g33265 (n_12848, n20513);
  and g33266 (n20514, n_12846, n_12848);
  and g33267 (n20515, n_12847, n_12848);
  not g33268 (n_12849, n20514);
  not g33269 (n_12850, n20515);
  and g33270 (n20516, n_12849, n_12850);
  and g33271 (n20517, n19942, n20039);
  not g33272 (n_12851, n20517);
  and g33273 (n20518, n_12442, n_12851);
  and g33274 (n20519, n9331, n12549);
  and g33275 (n20520, n8418, n12555);
  and g33276 (n20521, n8860, n12552);
  not g33277 (n_12852, n20520);
  not g33278 (n_12853, n20521);
  and g33279 (n20522, n_12852, n_12853);
  not g33280 (n_12854, n20519);
  and g33281 (n20523, n_12854, n20522);
  and g33282 (n20524, n_3428, n20523);
  and g33283 (n20525, n_9580, n20523);
  not g33284 (n_12855, n20524);
  not g33285 (n_12856, n20525);
  and g33286 (n20526, n_12855, n_12856);
  not g33287 (n_12857, n20526);
  and g33288 (n20527, \a[8] , n_12857);
  and g33289 (n20528, n_1106, n20526);
  not g33290 (n_12858, n20527);
  not g33291 (n_12859, n20528);
  and g33292 (n20529, n_12858, n_12859);
  not g33293 (n_12860, n20529);
  and g33294 (n20530, n20518, n_12860);
  not g33295 (n_12861, n20037);
  and g33296 (n20531, n20035, n_12861);
  not g33297 (n_12862, n20531);
  and g33298 (n20532, n_12439, n_12862);
  and g33299 (n20533, n9331, n12552);
  and g33300 (n20534, n8418, n12558);
  and g33301 (n20535, n8860, n12555);
  not g33302 (n_12863, n20534);
  not g33303 (n_12864, n20535);
  and g33304 (n20536, n_12863, n_12864);
  not g33305 (n_12865, n20533);
  and g33306 (n20537, n_12865, n20536);
  and g33307 (n20538, n_3428, n20537);
  and g33308 (n20539, n15791, n20537);
  not g33309 (n_12866, n20538);
  not g33310 (n_12867, n20539);
  and g33311 (n20540, n_12866, n_12867);
  not g33312 (n_12868, n20540);
  and g33313 (n20541, \a[8] , n_12868);
  and g33314 (n20542, n_1106, n20540);
  not g33315 (n_12869, n20541);
  not g33316 (n_12870, n20542);
  and g33317 (n20543, n_12869, n_12870);
  not g33318 (n_12871, n20543);
  and g33319 (n20544, n20532, n_12871);
  and g33320 (n20545, n19974, n20033);
  not g33321 (n_12872, n20545);
  and g33322 (n20546, n_12435, n_12872);
  and g33323 (n20547, n9331, n12555);
  and g33324 (n20548, n8418, n12561);
  and g33325 (n20549, n8860, n12558);
  not g33326 (n_12873, n20548);
  not g33327 (n_12874, n20549);
  and g33328 (n20550, n_12873, n_12874);
  not g33329 (n_12875, n20547);
  and g33330 (n20551, n_12875, n20550);
  and g33331 (n20552, n_3428, n20551);
  and g33332 (n20553, n15816, n20551);
  not g33333 (n_12876, n20552);
  not g33334 (n_12877, n20553);
  and g33335 (n20554, n_12876, n_12877);
  not g33336 (n_12878, n20554);
  and g33337 (n20555, \a[8] , n_12878);
  and g33338 (n20556, n_1106, n20554);
  not g33339 (n_12879, n20555);
  not g33340 (n_12880, n20556);
  and g33341 (n20557, n_12879, n_12880);
  not g33342 (n_12881, n20557);
  and g33343 (n20558, n20546, n_12881);
  and g33344 (n20559, n9331, n12558);
  and g33345 (n20560, n8418, n12564);
  and g33346 (n20561, n8860, n12561);
  and g33352 (n20564, n8421, n15847);
  not g33355 (n_12886, n20565);
  and g33356 (n20566, \a[8] , n_12886);
  not g33357 (n_12887, n20566);
  and g33358 (n20567, n_12886, n_12887);
  and g33359 (n20568, \a[8] , n_12887);
  not g33360 (n_12888, n20567);
  not g33361 (n_12889, n20568);
  and g33362 (n20569, n_12888, n_12889);
  not g33363 (n_12890, n20031);
  and g33364 (n20570, n20029, n_12890);
  not g33365 (n_12891, n20570);
  and g33366 (n20571, n_12432, n_12891);
  not g33367 (n_12892, n20569);
  and g33368 (n20572, n_12892, n20571);
  not g33369 (n_12893, n20572);
  and g33370 (n20573, n_12892, n_12893);
  and g33371 (n20574, n20571, n_12893);
  not g33372 (n_12894, n20573);
  not g33373 (n_12895, n20574);
  and g33374 (n20575, n_12894, n_12895);
  and g33375 (n20576, n_12425, n_12427);
  and g33376 (n20577, n_12426, n_12427);
  not g33377 (n_12896, n20576);
  not g33378 (n_12897, n20577);
  and g33379 (n20578, n_12896, n_12897);
  and g33380 (n20579, n9331, n12561);
  and g33381 (n20580, n8418, n12567);
  and g33382 (n20581, n8860, n12564);
  not g33383 (n_12898, n20580);
  not g33384 (n_12899, n20581);
  and g33385 (n20582, n_12898, n_12899);
  not g33386 (n_12900, n20579);
  and g33387 (n20583, n_12900, n20582);
  and g33388 (n20584, n_3428, n20583);
  and g33389 (n20585, n15905, n20583);
  not g33390 (n_12901, n20584);
  not g33391 (n_12902, n20585);
  and g33392 (n20586, n_12901, n_12902);
  not g33393 (n_12903, n20586);
  and g33394 (n20587, \a[8] , n_12903);
  and g33395 (n20588, n_1106, n20586);
  not g33396 (n_12904, n20587);
  not g33397 (n_12905, n20588);
  and g33398 (n20589, n_12904, n_12905);
  not g33399 (n_12906, n20578);
  not g33400 (n_12907, n20589);
  and g33401 (n20590, n_12906, n_12907);
  and g33402 (n20591, n9331, n12564);
  and g33403 (n20592, n8418, n12571);
  and g33404 (n20593, n8860, n12567);
  and g33410 (n20596, n8421, n_9006);
  not g33413 (n_12912, n20597);
  and g33414 (n20598, \a[8] , n_12912);
  not g33415 (n_12913, n20598);
  and g33416 (n20599, n_12912, n_12913);
  and g33417 (n20600, \a[8] , n_12913);
  not g33418 (n_12914, n20599);
  not g33419 (n_12915, n20600);
  and g33420 (n20601, n_12914, n_12915);
  not g33421 (n_12916, n20000);
  and g33422 (n20602, n_12916, n20011);
  not g33423 (n_12917, n20012);
  not g33424 (n_12918, n20602);
  and g33425 (n20603, n_12917, n_12918);
  not g33426 (n_12919, n20601);
  and g33427 (n20604, n_12919, n20603);
  not g33428 (n_12920, n20604);
  and g33429 (n20605, n_12919, n_12920);
  and g33430 (n20606, n20603, n_12920);
  not g33431 (n_12921, n20605);
  not g33432 (n_12922, n20606);
  and g33433 (n20607, n_12921, n_12922);
  not g33434 (n_12923, n19999);
  and g33435 (n20608, n19997, n_12923);
  not g33436 (n_12924, n20608);
  and g33437 (n20609, n_12916, n_12924);
  and g33438 (n20610, n9331, n12567);
  and g33439 (n20611, n8418, n12574);
  and g33440 (n20612, n8860, n12571);
  not g33441 (n_12925, n20611);
  not g33442 (n_12926, n20612);
  and g33443 (n20613, n_12925, n_12926);
  not g33444 (n_12927, n20610);
  and g33445 (n20614, n_12927, n20613);
  and g33446 (n20615, n_3428, n20614);
  and g33447 (n20616, n_10006, n20614);
  not g33448 (n_12928, n20615);
  not g33449 (n_12929, n20616);
  and g33450 (n20617, n_12928, n_12929);
  not g33451 (n_12930, n20617);
  and g33452 (n20618, \a[8] , n_12930);
  and g33453 (n20619, n_1106, n20617);
  not g33454 (n_12931, n20618);
  not g33455 (n_12932, n20619);
  and g33456 (n20620, n_12931, n_12932);
  not g33457 (n_12933, n20620);
  and g33458 (n20621, n20609, n_12933);
  and g33459 (n20622, n8860, n_6977);
  and g33460 (n20623, n9331, n12577);
  not g33461 (n_12934, n20622);
  not g33462 (n_12935, n20623);
  and g33463 (n20624, n_12934, n_12935);
  and g33464 (n20625, n8421, n_9032);
  not g33465 (n_12936, n20625);
  and g33466 (n20626, n20624, n_12936);
  not g33467 (n_12937, n20626);
  and g33468 (n20627, \a[8] , n_12937);
  not g33469 (n_12938, n20627);
  and g33470 (n20628, \a[8] , n_12938);
  and g33471 (n20629, n_12937, n_12938);
  not g33472 (n_12939, n20628);
  not g33473 (n_12940, n20629);
  and g33474 (n20630, n_12939, n_12940);
  and g33475 (n20631, n_3427, n_6977);
  not g33476 (n_12941, n20631);
  and g33477 (n20632, \a[8] , n_12941);
  not g33478 (n_12942, n20630);
  and g33479 (n20633, n_12942, n20632);
  and g33480 (n20634, n9331, n12574);
  and g33481 (n20635, n8418, n_6977);
  and g33482 (n20636, n8860, n12577);
  not g33483 (n_12943, n20635);
  not g33484 (n_12944, n20636);
  and g33485 (n20637, n_12943, n_12944);
  not g33486 (n_12945, n20634);
  and g33487 (n20638, n_12945, n20637);
  and g33488 (n20639, n_3428, n20638);
  and g33489 (n20640, n16094, n20638);
  not g33490 (n_12946, n20639);
  not g33491 (n_12947, n20640);
  and g33492 (n20641, n_12946, n_12947);
  not g33493 (n_12948, n20641);
  and g33494 (n20642, \a[8] , n_12948);
  and g33495 (n20643, n_1106, n20641);
  not g33496 (n_12949, n20642);
  not g33497 (n_12950, n20643);
  and g33498 (n20644, n_12949, n_12950);
  not g33499 (n_12951, n20644);
  and g33500 (n20645, n20633, n_12951);
  and g33501 (n20646, n19998, n20645);
  not g33502 (n_12952, n20646);
  and g33503 (n20647, n20645, n_12952);
  and g33504 (n20648, n19998, n_12952);
  not g33505 (n_12953, n20647);
  not g33506 (n_12954, n20648);
  and g33507 (n20649, n_12953, n_12954);
  and g33508 (n20650, n9331, n12571);
  and g33509 (n20651, n8418, n12577);
  and g33510 (n20652, n8860, n12574);
  and g33516 (n20655, n8421, n16013);
  not g33519 (n_12959, n20656);
  and g33520 (n20657, \a[8] , n_12959);
  not g33521 (n_12960, n20657);
  and g33522 (n20658, \a[8] , n_12960);
  and g33523 (n20659, n_12959, n_12960);
  not g33524 (n_12961, n20658);
  not g33525 (n_12962, n20659);
  and g33526 (n20660, n_12961, n_12962);
  not g33527 (n_12963, n20649);
  not g33528 (n_12964, n20660);
  and g33529 (n20661, n_12963, n_12964);
  not g33530 (n_12965, n20661);
  and g33531 (n20662, n_12952, n_12965);
  not g33532 (n_12966, n20609);
  and g33533 (n20663, n_12966, n20620);
  not g33534 (n_12967, n20621);
  not g33535 (n_12968, n20663);
  and g33536 (n20664, n_12967, n_12968);
  not g33537 (n_12969, n20662);
  and g33538 (n20665, n_12969, n20664);
  not g33539 (n_12970, n20665);
  and g33540 (n20666, n_12967, n_12970);
  not g33541 (n_12971, n20607);
  not g33542 (n_12972, n20666);
  and g33543 (n20667, n_12971, n_12972);
  not g33544 (n_12973, n20667);
  and g33545 (n20668, n_12920, n_12973);
  and g33546 (n20669, n20578, n20589);
  not g33547 (n_12974, n20590);
  not g33548 (n_12975, n20669);
  and g33549 (n20670, n_12974, n_12975);
  not g33550 (n_12976, n20668);
  and g33551 (n20671, n_12976, n20670);
  not g33552 (n_12977, n20671);
  and g33553 (n20672, n_12974, n_12977);
  not g33554 (n_12978, n20575);
  not g33555 (n_12979, n20672);
  and g33556 (n20673, n_12978, n_12979);
  not g33557 (n_12980, n20673);
  and g33558 (n20674, n_12893, n_12980);
  not g33559 (n_12981, n20558);
  and g33560 (n20675, n20546, n_12981);
  and g33561 (n20676, n_12881, n_12981);
  not g33562 (n_12982, n20675);
  not g33563 (n_12983, n20676);
  and g33564 (n20677, n_12982, n_12983);
  not g33565 (n_12984, n20674);
  not g33566 (n_12985, n20677);
  and g33567 (n20678, n_12984, n_12985);
  not g33568 (n_12986, n20678);
  and g33569 (n20679, n_12981, n_12986);
  not g33570 (n_12987, n20544);
  and g33571 (n20680, n20532, n_12987);
  and g33572 (n20681, n_12871, n_12987);
  not g33573 (n_12988, n20680);
  not g33574 (n_12989, n20681);
  and g33575 (n20682, n_12988, n_12989);
  not g33576 (n_12990, n20679);
  not g33577 (n_12991, n20682);
  and g33578 (n20683, n_12990, n_12991);
  not g33579 (n_12992, n20683);
  and g33580 (n20684, n_12987, n_12992);
  not g33581 (n_12993, n20518);
  and g33582 (n20685, n_12993, n20529);
  not g33583 (n_12994, n20530);
  not g33584 (n_12995, n20685);
  and g33585 (n20686, n_12994, n_12995);
  not g33586 (n_12996, n20684);
  and g33587 (n20687, n_12996, n20686);
  not g33588 (n_12997, n20687);
  and g33589 (n20688, n_12994, n_12997);
  not g33590 (n_12998, n20516);
  not g33591 (n_12999, n20688);
  and g33592 (n20689, n_12998, n_12999);
  not g33593 (n_13000, n20689);
  and g33594 (n20690, n_12848, n_13000);
  not g33595 (n_13001, n20498);
  not g33596 (n_13002, n20690);
  and g33597 (n20691, n_13001, n_13002);
  not g33598 (n_13003, n20691);
  and g33599 (n20692, n_12833, n_13003);
  not g33600 (n_13004, n20480);
  not g33601 (n_13005, n20692);
  and g33602 (n20693, n_13004, n_13005);
  not g33603 (n_13006, n20693);
  and g33604 (n20694, n_12818, n_13006);
  not g33605 (n_13007, n20463);
  and g33606 (n20695, n20451, n_13007);
  and g33607 (n20696, n_12806, n_13007);
  not g33608 (n_13008, n20695);
  not g33609 (n_13009, n20696);
  and g33610 (n20697, n_13008, n_13009);
  not g33611 (n_13010, n20694);
  not g33612 (n_13011, n20697);
  and g33613 (n20698, n_13010, n_13011);
  not g33614 (n_13012, n20698);
  and g33615 (n20699, n_13007, n_13012);
  not g33616 (n_13013, n20449);
  and g33617 (n20700, n20437, n_13013);
  and g33618 (n20701, n_12796, n_13013);
  not g33619 (n_13014, n20700);
  not g33620 (n_13015, n20701);
  and g33621 (n20702, n_13014, n_13015);
  not g33622 (n_13016, n20699);
  not g33623 (n_13017, n20702);
  and g33624 (n20703, n_13016, n_13017);
  not g33625 (n_13018, n20703);
  and g33626 (n20704, n_13013, n_13018);
  not g33627 (n_13019, n20423);
  and g33628 (n20705, n_13019, n20434);
  not g33629 (n_13020, n20435);
  not g33630 (n_13021, n20705);
  and g33631 (n20706, n_13020, n_13021);
  not g33632 (n_13022, n20704);
  and g33633 (n20707, n_13022, n20706);
  not g33634 (n_13023, n20707);
  and g33635 (n20708, n_13020, n_13023);
  not g33636 (n_13024, n20421);
  not g33637 (n_13025, n20708);
  and g33638 (n20709, n_13024, n_13025);
  not g33639 (n_13026, n20709);
  and g33640 (n20710, n_12774, n_13026);
  not g33641 (n_13027, n20403);
  not g33642 (n_13028, n20710);
  and g33643 (n20711, n_13027, n_13028);
  not g33644 (n_13029, n20711);
  and g33645 (n20712, n_12759, n_13029);
  not g33646 (n_13030, n20385);
  not g33647 (n_13031, n20712);
  and g33648 (n20713, n_13030, n_13031);
  not g33649 (n_13032, n20713);
  and g33650 (n20714, n_12744, n_13032);
  not g33651 (n_13033, n20368);
  and g33652 (n20715, n20356, n_13033);
  and g33653 (n20716, n_12732, n_13033);
  not g33654 (n_13034, n20715);
  not g33655 (n_13035, n20716);
  and g33656 (n20717, n_13034, n_13035);
  not g33657 (n_13036, n20714);
  not g33658 (n_13037, n20717);
  and g33659 (n20718, n_13036, n_13037);
  not g33660 (n_13038, n20718);
  and g33661 (n20719, n_13033, n_13038);
  not g33662 (n_13039, n20354);
  and g33663 (n20720, n20342, n_13039);
  and g33664 (n20721, n_12722, n_13039);
  not g33665 (n_13040, n20720);
  not g33666 (n_13041, n20721);
  and g33667 (n20722, n_13040, n_13041);
  not g33668 (n_13042, n20719);
  not g33669 (n_13043, n20722);
  and g33670 (n20723, n_13042, n_13043);
  not g33671 (n_13044, n20723);
  and g33672 (n20724, n_13039, n_13044);
  not g33673 (n_13045, n20328);
  and g33674 (n20725, n_13045, n20339);
  not g33675 (n_13046, n20340);
  not g33676 (n_13047, n20725);
  and g33677 (n20726, n_13046, n_13047);
  not g33678 (n_13048, n20724);
  and g33679 (n20727, n_13048, n20726);
  not g33680 (n_13049, n20727);
  and g33681 (n20728, n_13046, n_13049);
  not g33682 (n_13050, n20326);
  not g33683 (n_13051, n20728);
  and g33684 (n20729, n_13050, n_13051);
  not g33685 (n_13052, n20729);
  and g33686 (n20730, n_12700, n_13052);
  not g33687 (n_13053, n20308);
  not g33688 (n_13054, n20730);
  and g33689 (n20731, n_13053, n_13054);
  not g33690 (n_13055, n20731);
  and g33691 (n20732, n_12685, n_13055);
  not g33692 (n_13056, n20291);
  and g33693 (n20733, n20279, n_13056);
  and g33694 (n20734, n_12673, n_13056);
  not g33695 (n_13057, n20733);
  not g33696 (n_13058, n20734);
  and g33697 (n20735, n_13057, n_13058);
  not g33698 (n_13059, n20732);
  not g33699 (n_13060, n20735);
  and g33700 (n20736, n_13059, n_13060);
  not g33701 (n_13061, n20736);
  and g33702 (n20737, n_13056, n_13061);
  not g33703 (n_13062, n20277);
  and g33704 (n20738, n20265, n_13062);
  and g33705 (n20739, n_12663, n_13062);
  not g33706 (n_13063, n20738);
  not g33707 (n_13064, n20739);
  and g33708 (n20740, n_13063, n_13064);
  not g33709 (n_13065, n20737);
  not g33710 (n_13066, n20740);
  and g33711 (n20741, n_13065, n_13066);
  not g33712 (n_13067, n20741);
  and g33713 (n20742, n_13062, n_13067);
  not g33714 (n_13068, n20263);
  and g33715 (n20743, n20251, n_13068);
  and g33716 (n20744, n_12653, n_13068);
  not g33717 (n_13069, n20743);
  not g33718 (n_13070, n20744);
  and g33719 (n20745, n_13069, n_13070);
  not g33720 (n_13071, n20742);
  not g33721 (n_13072, n20745);
  and g33722 (n20746, n_13071, n_13072);
  not g33723 (n_13073, n20746);
  and g33724 (n20747, n_13068, n_13073);
  not g33725 (n_13074, n20249);
  and g33726 (n20748, n20237, n_13074);
  and g33727 (n20749, n_12643, n_13074);
  not g33728 (n_13075, n20748);
  not g33729 (n_13076, n20749);
  and g33730 (n20750, n_13075, n_13076);
  not g33731 (n_13077, n20747);
  not g33732 (n_13078, n20750);
  and g33733 (n20751, n_13077, n_13078);
  not g33734 (n_13079, n20751);
  and g33735 (n20752, n_13074, n_13079);
  not g33736 (n_13080, n20235);
  and g33737 (n20753, n20223, n_13080);
  and g33738 (n20754, n_12633, n_13080);
  not g33739 (n_13081, n20753);
  not g33740 (n_13082, n20754);
  and g33741 (n20755, n_13081, n_13082);
  not g33742 (n_13083, n20752);
  not g33743 (n_13084, n20755);
  and g33744 (n20756, n_13083, n_13084);
  not g33745 (n_13085, n20756);
  and g33746 (n20757, n_13080, n_13085);
  not g33747 (n_13086, n20221);
  and g33748 (n20758, n20209, n_13086);
  and g33749 (n20759, n_12622, n_13086);
  not g33750 (n_13087, n20758);
  not g33751 (n_13088, n20759);
  and g33752 (n20760, n_13087, n_13088);
  not g33753 (n_13089, n20757);
  not g33754 (n_13090, n20760);
  and g33755 (n20761, n_13089, n_13090);
  not g33756 (n_13091, n20761);
  and g33757 (n20762, n_13086, n_13091);
  not g33758 (n_13092, n20207);
  and g33759 (n20763, n20195, n_13092);
  and g33760 (n20764, n_12612, n_13092);
  not g33761 (n_13093, n20763);
  not g33762 (n_13094, n20764);
  and g33763 (n20765, n_13093, n_13094);
  not g33764 (n_13095, n20762);
  not g33765 (n_13096, n20765);
  and g33766 (n20766, n_13095, n_13096);
  not g33767 (n_13097, n20766);
  and g33768 (n20767, n_13092, n_13097);
  not g33769 (n_13098, n20193);
  and g33770 (n20768, n20181, n_13098);
  and g33771 (n20769, n_12601, n_13098);
  not g33772 (n_13099, n20768);
  not g33773 (n_13100, n20769);
  and g33774 (n20770, n_13099, n_13100);
  not g33775 (n_13101, n20767);
  not g33776 (n_13102, n20770);
  and g33777 (n20771, n_13101, n_13102);
  not g33778 (n_13103, n20771);
  and g33779 (n20772, n_13098, n_13103);
  not g33780 (n_13104, n20179);
  and g33781 (n20773, n20167, n_13104);
  and g33782 (n20774, n_12591, n_13104);
  not g33783 (n_13105, n20773);
  not g33784 (n_13106, n20774);
  and g33785 (n20775, n_13105, n_13106);
  not g33786 (n_13107, n20772);
  not g33787 (n_13108, n20775);
  and g33788 (n20776, n_13107, n_13108);
  not g33789 (n_13109, n20776);
  and g33790 (n20777, n_13104, n_13109);
  not g33791 (n_13110, n20153);
  and g33792 (n20778, n_13110, n20164);
  not g33793 (n_13111, n20165);
  not g33794 (n_13112, n20778);
  and g33795 (n20779, n_13111, n_13112);
  not g33796 (n_13113, n20777);
  and g33797 (n20780, n_13113, n20779);
  not g33798 (n_13114, n20780);
  and g33799 (n20781, n_13111, n_13114);
  not g33800 (n_13115, n20151);
  not g33801 (n_13116, n20781);
  and g33802 (n20782, n_13115, n_13116);
  and g33803 (n20783, n20151, n20781);
  not g33804 (n_13117, n20782);
  not g33805 (n_13118, n20783);
  and g33806 (n20784, n_13117, n_13118);
  and g33807 (n20785, n71, n13941);
  and g33808 (n20786, n9867, n13633);
  and g33809 (n20787, n10434, n_7540);
  and g33815 (n20790, n9870, n14136);
  not g33818 (n_13123, n20791);
  and g33819 (n20792, \a[5] , n_13123);
  not g33820 (n_13124, n20792);
  and g33821 (n20793, \a[5] , n_13124);
  and g33822 (n20794, n_13123, n_13124);
  not g33823 (n_13125, n20793);
  not g33824 (n_13126, n20794);
  and g33825 (n20795, n_13125, n_13126);
  not g33826 (n_13127, n20795);
  and g33827 (n20796, n20784, n_13127);
  not g33828 (n_13128, n20796);
  and g33829 (n20797, n_13117, n_13128);
  not g33830 (n_13129, n20148);
  not g33831 (n_13130, n20797);
  and g33832 (n20798, n_13129, n_13130);
  and g33833 (n20799, n20148, n20797);
  not g33834 (n_13131, n20798);
  not g33835 (n_13132, n20799);
  and g33836 (n20800, n_13131, n_13132);
  and g33837 (n20801, n20784, n_13128);
  and g33838 (n20802, n_13127, n_13128);
  not g33839 (n_13133, n20801);
  not g33840 (n_13134, n20802);
  and g33841 (n20803, n_13133, n_13134);
  and g33842 (n20804, n71, n_7540);
  and g33843 (n20805, n9867, n13630);
  and g33844 (n20806, n10434, n13633);
  and g33850 (n20809, n9870, n_7563);
  not g33853 (n_13139, n20810);
  and g33854 (n20811, \a[5] , n_13139);
  not g33855 (n_13140, n20811);
  and g33856 (n20812, n_13139, n_13140);
  and g33857 (n20813, \a[5] , n_13140);
  not g33858 (n_13141, n20812);
  not g33859 (n_13142, n20813);
  and g33860 (n20814, n_13141, n_13142);
  not g33861 (n_13143, n20779);
  and g33862 (n20815, n20777, n_13143);
  not g33863 (n_13144, n20815);
  and g33864 (n20816, n_13114, n_13144);
  not g33865 (n_13145, n20814);
  and g33866 (n20817, n_13145, n20816);
  not g33867 (n_13146, n20817);
  and g33868 (n20818, n_13145, n_13146);
  and g33869 (n20819, n20816, n_13146);
  not g33870 (n_13147, n20818);
  not g33871 (n_13148, n20819);
  and g33872 (n20820, n_13147, n_13148);
  not g33873 (n_13149, n11715);
  and g33874 (n20821, n_13149, n_6353);
  not g33875 (n_13150, n20821);
  and g33876 (n20822, n_7417, n_13150);
  and g33877 (n20823, n11055, n13941);
  not g33878 (n_13151, n20822);
  not g33879 (n_13152, n20823);
  and g33880 (n20824, n_13151, n_13152);
  not g33881 (n_13153, n13951);
  and g33882 (n20825, n11057, n_13153);
  not g33883 (n_13154, n20825);
  and g33884 (n20826, n20824, n_13154);
  not g33885 (n_13155, n20826);
  and g33886 (n20827, \a[2] , n_13155);
  not g33887 (n_13156, n20827);
  and g33888 (n20828, \a[2] , n_13156);
  and g33889 (n20829, n_13155, n_13156);
  not g33890 (n_13157, n20828);
  not g33891 (n_13158, n20829);
  and g33892 (n20830, n_13157, n_13158);
  not g33893 (n_13159, n20820);
  not g33894 (n_13160, n20830);
  and g33895 (n20831, n_13159, n_13160);
  not g33896 (n_13161, n20831);
  and g33897 (n20832, n_13146, n_13161);
  not g33898 (n_13162, n20803);
  not g33899 (n_13163, n20832);
  and g33900 (n20833, n_13162, n_13163);
  and g33901 (n20834, n20803, n20832);
  not g33902 (n_13164, n20833);
  not g33903 (n_13165, n20834);
  and g33904 (n20835, n_13164, n_13165);
  and g33905 (n20836, n_13159, n_13161);
  and g33906 (n20837, n_13160, n_13161);
  not g33907 (n_13166, n20836);
  not g33908 (n_13167, n20837);
  and g33909 (n20838, n_13166, n_13167);
  and g33910 (n20839, n71, n13633);
  and g33911 (n20840, n9867, n13597);
  and g33912 (n20841, n10434, n13630);
  and g33918 (n20844, n9870, n13929);
  not g33921 (n_13172, n20845);
  and g33922 (n20846, \a[5] , n_13172);
  not g33923 (n_13173, n20846);
  and g33924 (n20847, n_13172, n_13173);
  and g33925 (n20848, \a[5] , n_13173);
  not g33926 (n_13174, n20847);
  not g33927 (n_13175, n20848);
  and g33928 (n20849, n_13174, n_13175);
  and g33929 (n20850, n_13107, n_13109);
  and g33930 (n20851, n_13108, n_13109);
  not g33931 (n_13176, n20850);
  not g33932 (n_13177, n20851);
  and g33933 (n20852, n_13176, n_13177);
  not g33934 (n_13178, n20849);
  not g33935 (n_13179, n20852);
  and g33936 (n20853, n_13178, n_13179);
  not g33937 (n_13180, n20853);
  and g33938 (n20854, n_13178, n_13180);
  and g33939 (n20855, n_13179, n_13180);
  not g33940 (n_13181, n20854);
  not g33941 (n_13182, n20855);
  and g33942 (n20856, n_13181, n_13182);
  and g33943 (n20857, n71, n13630);
  and g33944 (n20858, n9867, n13515);
  and g33945 (n20859, n10434, n13597);
  and g33951 (n20862, n9870, n13976);
  not g33954 (n_13187, n20863);
  and g33955 (n20864, \a[5] , n_13187);
  not g33956 (n_13188, n20864);
  and g33957 (n20865, n_13187, n_13188);
  and g33958 (n20866, \a[5] , n_13188);
  not g33959 (n_13189, n20865);
  not g33960 (n_13190, n20866);
  and g33961 (n20867, n_13189, n_13190);
  and g33962 (n20868, n_13101, n_13103);
  and g33963 (n20869, n_13102, n_13103);
  not g33964 (n_13191, n20868);
  not g33965 (n_13192, n20869);
  and g33966 (n20870, n_13191, n_13192);
  not g33967 (n_13193, n20867);
  not g33968 (n_13194, n20870);
  and g33969 (n20871, n_13193, n_13194);
  not g33970 (n_13195, n20871);
  and g33971 (n20872, n_13193, n_13195);
  and g33972 (n20873, n_13194, n_13195);
  not g33973 (n_13196, n20872);
  not g33974 (n_13197, n20873);
  and g33975 (n20874, n_13196, n_13197);
  and g33976 (n20875, n71, n13597);
  and g33977 (n20876, n9867, n13521);
  and g33978 (n20877, n10434, n13515);
  and g33984 (n20880, n9870, n_7765);
  not g33987 (n_13202, n20881);
  and g33988 (n20882, \a[5] , n_13202);
  not g33989 (n_13203, n20882);
  and g33990 (n20883, n_13202, n_13203);
  and g33991 (n20884, \a[5] , n_13203);
  not g33992 (n_13204, n20883);
  not g33993 (n_13205, n20884);
  and g33994 (n20885, n_13204, n_13205);
  and g33995 (n20886, n_13095, n_13097);
  and g33996 (n20887, n_13096, n_13097);
  not g33997 (n_13206, n20886);
  not g33998 (n_13207, n20887);
  and g33999 (n20888, n_13206, n_13207);
  not g34000 (n_13208, n20885);
  not g34001 (n_13209, n20888);
  and g34002 (n20889, n_13208, n_13209);
  not g34003 (n_13210, n20889);
  and g34004 (n20890, n_13208, n_13210);
  and g34005 (n20891, n_13209, n_13210);
  not g34006 (n_13211, n20890);
  not g34007 (n_13212, n20891);
  and g34008 (n20892, n_13211, n_13212);
  and g34009 (n20893, n71, n13515);
  and g34010 (n20894, n9867, n13518);
  and g34011 (n20895, n10434, n13521);
  and g34017 (n20898, n9870, n13541);
  not g34020 (n_13217, n20899);
  and g34021 (n20900, \a[5] , n_13217);
  not g34022 (n_13218, n20900);
  and g34023 (n20901, n_13217, n_13218);
  and g34024 (n20902, \a[5] , n_13218);
  not g34025 (n_13219, n20901);
  not g34026 (n_13220, n20902);
  and g34027 (n20903, n_13219, n_13220);
  and g34028 (n20904, n_13089, n_13091);
  and g34029 (n20905, n_13090, n_13091);
  not g34030 (n_13221, n20904);
  not g34031 (n_13222, n20905);
  and g34032 (n20906, n_13221, n_13222);
  not g34033 (n_13223, n20903);
  not g34034 (n_13224, n20906);
  and g34035 (n20907, n_13223, n_13224);
  not g34036 (n_13225, n20907);
  and g34037 (n20908, n_13223, n_13225);
  and g34038 (n20909, n_13224, n_13225);
  not g34039 (n_13226, n20908);
  not g34040 (n_13227, n20909);
  and g34041 (n20910, n_13226, n_13227);
  and g34042 (n20911, n71, n13521);
  and g34043 (n20912, n9867, n13491);
  and g34044 (n20913, n10434, n13518);
  and g34050 (n20916, n9870, n_7677);
  not g34053 (n_13232, n20917);
  and g34054 (n20918, \a[5] , n_13232);
  not g34055 (n_13233, n20918);
  and g34056 (n20919, n_13232, n_13233);
  and g34057 (n20920, \a[5] , n_13233);
  not g34058 (n_13234, n20919);
  not g34059 (n_13235, n20920);
  and g34060 (n20921, n_13234, n_13235);
  and g34061 (n20922, n_13083, n_13085);
  and g34062 (n20923, n_13084, n_13085);
  not g34063 (n_13236, n20922);
  not g34064 (n_13237, n20923);
  and g34065 (n20924, n_13236, n_13237);
  not g34066 (n_13238, n20921);
  not g34067 (n_13239, n20924);
  and g34068 (n20925, n_13238, n_13239);
  not g34069 (n_13240, n20925);
  and g34070 (n20926, n_13238, n_13240);
  and g34071 (n20927, n_13239, n_13240);
  not g34072 (n_13241, n20926);
  not g34073 (n_13242, n20927);
  and g34074 (n20928, n_13241, n_13242);
  and g34075 (n20929, n71, n13518);
  and g34076 (n20930, n9867, n12889);
  and g34077 (n20931, n10434, n13491);
  and g34083 (n20934, n9870, n13584);
  not g34086 (n_13247, n20935);
  and g34087 (n20936, \a[5] , n_13247);
  not g34088 (n_13248, n20936);
  and g34089 (n20937, n_13247, n_13248);
  and g34090 (n20938, \a[5] , n_13248);
  not g34091 (n_13249, n20937);
  not g34092 (n_13250, n20938);
  and g34093 (n20939, n_13249, n_13250);
  and g34094 (n20940, n_13077, n_13079);
  and g34095 (n20941, n_13078, n_13079);
  not g34096 (n_13251, n20940);
  not g34097 (n_13252, n20941);
  and g34098 (n20942, n_13251, n_13252);
  not g34099 (n_13253, n20939);
  not g34100 (n_13254, n20942);
  and g34101 (n20943, n_13253, n_13254);
  not g34102 (n_13255, n20943);
  and g34103 (n20944, n_13253, n_13255);
  and g34104 (n20945, n_13254, n_13255);
  not g34105 (n_13256, n20944);
  not g34106 (n_13257, n20945);
  and g34107 (n20946, n_13256, n_13257);
  and g34108 (n20947, n71, n13491);
  and g34109 (n20948, n9867, n12769);
  and g34110 (n20949, n10434, n12889);
  and g34116 (n20952, n9870, n_7447);
  not g34119 (n_13262, n20953);
  and g34120 (n20954, \a[5] , n_13262);
  not g34121 (n_13263, n20954);
  and g34122 (n20955, n_13262, n_13263);
  and g34123 (n20956, \a[5] , n_13263);
  not g34124 (n_13264, n20955);
  not g34125 (n_13265, n20956);
  and g34126 (n20957, n_13264, n_13265);
  and g34127 (n20958, n_13071, n_13073);
  and g34128 (n20959, n_13072, n_13073);
  not g34129 (n_13266, n20958);
  not g34130 (n_13267, n20959);
  and g34131 (n20960, n_13266, n_13267);
  not g34132 (n_13268, n20957);
  not g34133 (n_13269, n20960);
  and g34134 (n20961, n_13268, n_13269);
  not g34135 (n_13270, n20961);
  and g34136 (n20962, n_13268, n_13270);
  and g34137 (n20963, n_13269, n_13270);
  not g34138 (n_13271, n20962);
  not g34139 (n_13272, n20963);
  and g34140 (n20964, n_13271, n_13272);
  and g34141 (n20965, n71, n12889);
  and g34142 (n20966, n9867, n12502);
  and g34143 (n20967, n10434, n12769);
  and g34149 (n20970, n9870, n12895);
  not g34152 (n_13277, n20971);
  and g34153 (n20972, \a[5] , n_13277);
  not g34154 (n_13278, n20972);
  and g34155 (n20973, n_13277, n_13278);
  and g34156 (n20974, \a[5] , n_13278);
  not g34157 (n_13279, n20973);
  not g34158 (n_13280, n20974);
  and g34159 (n20975, n_13279, n_13280);
  and g34160 (n20976, n_13065, n_13067);
  and g34161 (n20977, n_13066, n_13067);
  not g34162 (n_13281, n20976);
  not g34163 (n_13282, n20977);
  and g34164 (n20978, n_13281, n_13282);
  not g34165 (n_13283, n20975);
  not g34166 (n_13284, n20978);
  and g34167 (n20979, n_13283, n_13284);
  not g34168 (n_13285, n20979);
  and g34169 (n20980, n_13283, n_13285);
  and g34170 (n20981, n_13284, n_13285);
  not g34171 (n_13286, n20980);
  not g34172 (n_13287, n20981);
  and g34173 (n20982, n_13286, n_13287);
  and g34174 (n20983, n71, n12769);
  and g34175 (n20984, n9867, n12370);
  and g34176 (n20985, n10434, n12502);
  and g34182 (n20988, n9870, n12999);
  not g34185 (n_13292, n20989);
  and g34186 (n20990, \a[5] , n_13292);
  not g34187 (n_13293, n20990);
  and g34188 (n20991, n_13292, n_13293);
  and g34189 (n20992, \a[5] , n_13293);
  not g34190 (n_13294, n20991);
  not g34191 (n_13295, n20992);
  and g34192 (n20993, n_13294, n_13295);
  and g34193 (n20994, n_13059, n_13061);
  and g34194 (n20995, n_13060, n_13061);
  not g34195 (n_13296, n20994);
  not g34196 (n_13297, n20995);
  and g34197 (n20996, n_13296, n_13297);
  not g34198 (n_13298, n20993);
  not g34199 (n_13299, n20996);
  and g34200 (n20997, n_13298, n_13299);
  not g34201 (n_13300, n20997);
  and g34202 (n20998, n_13298, n_13300);
  and g34203 (n20999, n_13299, n_13300);
  not g34204 (n_13301, n20998);
  not g34205 (n_13302, n20999);
  and g34206 (n21000, n_13301, n_13302);
  and g34207 (n21001, n20308, n20730);
  not g34208 (n_13303, n21001);
  and g34209 (n21002, n_13055, n_13303);
  and g34210 (n21003, n71, n12502);
  and g34211 (n21004, n9867, n12505);
  and g34212 (n21005, n10434, n12370);
  not g34213 (n_13304, n21004);
  not g34214 (n_13305, n21005);
  and g34215 (n21006, n_13304, n_13305);
  not g34216 (n_13306, n21003);
  and g34217 (n21007, n_13306, n21006);
  and g34218 (n21008, n_4684, n21007);
  and g34219 (n21009, n13736, n21007);
  not g34220 (n_13307, n21008);
  not g34221 (n_13308, n21009);
  and g34222 (n21010, n_13307, n_13308);
  not g34223 (n_13309, n21010);
  and g34224 (n21011, \a[5] , n_13309);
  and g34225 (n21012, n_3, n21010);
  not g34226 (n_13310, n21011);
  not g34227 (n_13311, n21012);
  and g34228 (n21013, n_13310, n_13311);
  not g34229 (n_13312, n21013);
  and g34230 (n21014, n21002, n_13312);
  and g34231 (n21015, n20326, n20728);
  not g34232 (n_13313, n21015);
  and g34233 (n21016, n_13052, n_13313);
  and g34234 (n21017, n71, n12370);
  and g34235 (n21018, n9867, n12508);
  and g34236 (n21019, n10434, n12505);
  not g34237 (n_13314, n21018);
  not g34238 (n_13315, n21019);
  and g34239 (n21020, n_13314, n_13315);
  not g34240 (n_13316, n21017);
  and g34241 (n21021, n_13316, n21020);
  and g34242 (n21022, n_4684, n21021);
  and g34243 (n21023, n13748, n21021);
  not g34244 (n_13317, n21022);
  not g34245 (n_13318, n21023);
  and g34246 (n21024, n_13317, n_13318);
  not g34247 (n_13319, n21024);
  and g34248 (n21025, \a[5] , n_13319);
  and g34249 (n21026, n_3, n21024);
  not g34250 (n_13320, n21025);
  not g34251 (n_13321, n21026);
  and g34252 (n21027, n_13320, n_13321);
  not g34253 (n_13322, n21027);
  and g34254 (n21028, n21016, n_13322);
  and g34255 (n21029, n71, n12505);
  and g34256 (n21030, n9867, n12513);
  and g34257 (n21031, n10434, n12508);
  and g34263 (n21034, n9870, n_7804);
  not g34266 (n_13327, n21035);
  and g34267 (n21036, \a[5] , n_13327);
  not g34268 (n_13328, n21036);
  and g34269 (n21037, n_13327, n_13328);
  and g34270 (n21038, \a[5] , n_13328);
  not g34271 (n_13329, n21037);
  not g34272 (n_13330, n21038);
  and g34273 (n21039, n_13329, n_13330);
  not g34274 (n_13331, n20726);
  and g34275 (n21040, n20724, n_13331);
  not g34276 (n_13332, n21040);
  and g34277 (n21041, n_13049, n_13332);
  not g34278 (n_13333, n21039);
  and g34279 (n21042, n_13333, n21041);
  not g34280 (n_13334, n21042);
  and g34281 (n21043, n_13333, n_13334);
  and g34282 (n21044, n21041, n_13334);
  not g34283 (n_13335, n21043);
  not g34284 (n_13336, n21044);
  and g34285 (n21045, n_13335, n_13336);
  and g34286 (n21046, n71, n12508);
  and g34287 (n21047, n9867, n12511);
  and g34288 (n21048, n10434, n12513);
  and g34294 (n21051, n9870, n13863);
  not g34297 (n_13341, n21052);
  and g34298 (n21053, \a[5] , n_13341);
  not g34299 (n_13342, n21053);
  and g34300 (n21054, n_13341, n_13342);
  and g34301 (n21055, \a[5] , n_13342);
  not g34302 (n_13343, n21054);
  not g34303 (n_13344, n21055);
  and g34304 (n21056, n_13343, n_13344);
  and g34305 (n21057, n_13042, n_13044);
  and g34306 (n21058, n_13043, n_13044);
  not g34307 (n_13345, n21057);
  not g34308 (n_13346, n21058);
  and g34309 (n21059, n_13345, n_13346);
  not g34310 (n_13347, n21056);
  not g34311 (n_13348, n21059);
  and g34312 (n21060, n_13347, n_13348);
  not g34313 (n_13349, n21060);
  and g34314 (n21061, n_13347, n_13349);
  and g34315 (n21062, n_13348, n_13349);
  not g34316 (n_13350, n21061);
  not g34317 (n_13351, n21062);
  and g34318 (n21063, n_13350, n_13351);
  and g34319 (n21064, n71, n12513);
  and g34320 (n21065, n9867, n12516);
  and g34321 (n21066, n10434, n12511);
  and g34327 (n21069, n9870, n14177);
  not g34330 (n_13356, n21070);
  and g34331 (n21071, \a[5] , n_13356);
  not g34332 (n_13357, n21071);
  and g34333 (n21072, n_13356, n_13357);
  and g34334 (n21073, \a[5] , n_13357);
  not g34335 (n_13358, n21072);
  not g34336 (n_13359, n21073);
  and g34337 (n21074, n_13358, n_13359);
  and g34338 (n21075, n_13036, n_13038);
  and g34339 (n21076, n_13037, n_13038);
  not g34340 (n_13360, n21075);
  not g34341 (n_13361, n21076);
  and g34342 (n21077, n_13360, n_13361);
  not g34343 (n_13362, n21074);
  not g34344 (n_13363, n21077);
  and g34345 (n21078, n_13362, n_13363);
  not g34346 (n_13364, n21078);
  and g34347 (n21079, n_13362, n_13364);
  and g34348 (n21080, n_13363, n_13364);
  not g34349 (n_13365, n21079);
  not g34350 (n_13366, n21080);
  and g34351 (n21081, n_13365, n_13366);
  and g34352 (n21082, n20385, n20712);
  not g34353 (n_13367, n21082);
  and g34354 (n21083, n_13032, n_13367);
  and g34355 (n21084, n71, n12511);
  and g34356 (n21085, n9867, n12519);
  and g34357 (n21086, n10434, n12516);
  not g34358 (n_13368, n21085);
  not g34359 (n_13369, n21086);
  and g34360 (n21087, n_13368, n_13369);
  not g34361 (n_13370, n21084);
  and g34362 (n21088, n_13370, n21087);
  and g34363 (n21089, n_4684, n21088);
  and g34364 (n21090, n14233, n21088);
  not g34365 (n_13371, n21089);
  not g34366 (n_13372, n21090);
  and g34367 (n21091, n_13371, n_13372);
  not g34368 (n_13373, n21091);
  and g34369 (n21092, \a[5] , n_13373);
  and g34370 (n21093, n_3, n21091);
  not g34371 (n_13374, n21092);
  not g34372 (n_13375, n21093);
  and g34373 (n21094, n_13374, n_13375);
  not g34374 (n_13376, n21094);
  and g34375 (n21095, n21083, n_13376);
  and g34376 (n21096, n20403, n20710);
  not g34377 (n_13377, n21096);
  and g34378 (n21097, n_13029, n_13377);
  and g34379 (n21098, n71, n12516);
  and g34380 (n21099, n9867, n12522);
  and g34381 (n21100, n10434, n12519);
  not g34382 (n_13378, n21099);
  not g34383 (n_13379, n21100);
  and g34384 (n21101, n_13378, n_13379);
  not g34385 (n_13380, n21098);
  and g34386 (n21102, n_13380, n21101);
  and g34387 (n21103, n_4684, n21102);
  and g34388 (n21104, n14443, n21102);
  not g34389 (n_13381, n21103);
  not g34390 (n_13382, n21104);
  and g34391 (n21105, n_13381, n_13382);
  not g34392 (n_13383, n21105);
  and g34393 (n21106, \a[5] , n_13383);
  and g34394 (n21107, n_3, n21105);
  not g34395 (n_13384, n21106);
  not g34396 (n_13385, n21107);
  and g34397 (n21108, n_13384, n_13385);
  not g34398 (n_13386, n21108);
  and g34399 (n21109, n21097, n_13386);
  and g34400 (n21110, n20421, n20708);
  not g34401 (n_13387, n21110);
  and g34402 (n21111, n_13026, n_13387);
  and g34403 (n21112, n71, n12519);
  and g34404 (n21113, n9867, n12525);
  and g34405 (n21114, n10434, n12522);
  not g34406 (n_13388, n21113);
  not g34407 (n_13389, n21114);
  and g34408 (n21115, n_13388, n_13389);
  not g34409 (n_13390, n21112);
  and g34410 (n21116, n_13390, n21115);
  and g34411 (n21117, n_4684, n21116);
  and g34412 (n21118, n_10664, n21116);
  not g34413 (n_13391, n21117);
  not g34414 (n_13392, n21118);
  and g34415 (n21119, n_13391, n_13392);
  not g34416 (n_13393, n21119);
  and g34417 (n21120, \a[5] , n_13393);
  and g34418 (n21121, n_3, n21119);
  not g34419 (n_13394, n21120);
  not g34420 (n_13395, n21121);
  and g34421 (n21122, n_13394, n_13395);
  not g34422 (n_13396, n21122);
  and g34423 (n21123, n21111, n_13396);
  and g34424 (n21124, n71, n12522);
  and g34425 (n21125, n9867, n12528);
  and g34426 (n21126, n10434, n12525);
  and g34432 (n21129, n9870, n14837);
  not g34435 (n_13401, n21130);
  and g34436 (n21131, \a[5] , n_13401);
  not g34437 (n_13402, n21131);
  and g34438 (n21132, n_13401, n_13402);
  and g34439 (n21133, \a[5] , n_13402);
  not g34440 (n_13403, n21132);
  not g34441 (n_13404, n21133);
  and g34442 (n21134, n_13403, n_13404);
  not g34443 (n_13405, n20706);
  and g34444 (n21135, n20704, n_13405);
  not g34445 (n_13406, n21135);
  and g34446 (n21136, n_13023, n_13406);
  not g34447 (n_13407, n21134);
  and g34448 (n21137, n_13407, n21136);
  not g34449 (n_13408, n21137);
  and g34450 (n21138, n_13407, n_13408);
  and g34451 (n21139, n21136, n_13408);
  not g34452 (n_13409, n21138);
  not g34453 (n_13410, n21139);
  and g34454 (n21140, n_13409, n_13410);
  and g34455 (n21141, n71, n12525);
  and g34456 (n21142, n9867, n12531);
  and g34457 (n21143, n10434, n12528);
  and g34463 (n21146, n9870, n14608);
  not g34466 (n_13415, n21147);
  and g34467 (n21148, \a[5] , n_13415);
  not g34468 (n_13416, n21148);
  and g34469 (n21149, n_13415, n_13416);
  and g34470 (n21150, \a[5] , n_13416);
  not g34471 (n_13417, n21149);
  not g34472 (n_13418, n21150);
  and g34473 (n21151, n_13417, n_13418);
  and g34474 (n21152, n_13016, n_13018);
  and g34475 (n21153, n_13017, n_13018);
  not g34476 (n_13419, n21152);
  not g34477 (n_13420, n21153);
  and g34478 (n21154, n_13419, n_13420);
  not g34479 (n_13421, n21151);
  not g34480 (n_13422, n21154);
  and g34481 (n21155, n_13421, n_13422);
  not g34482 (n_13423, n21155);
  and g34483 (n21156, n_13421, n_13423);
  and g34484 (n21157, n_13422, n_13423);
  not g34485 (n_13424, n21156);
  not g34486 (n_13425, n21157);
  and g34487 (n21158, n_13424, n_13425);
  and g34488 (n21159, n71, n12528);
  and g34489 (n21160, n9867, n12534);
  and g34490 (n21161, n10434, n12531);
  and g34496 (n21164, n9870, n_8448);
  not g34499 (n_13430, n21165);
  and g34500 (n21166, \a[5] , n_13430);
  not g34501 (n_13431, n21166);
  and g34502 (n21167, n_13430, n_13431);
  and g34503 (n21168, \a[5] , n_13431);
  not g34504 (n_13432, n21167);
  not g34505 (n_13433, n21168);
  and g34506 (n21169, n_13432, n_13433);
  and g34507 (n21170, n_13010, n_13012);
  and g34508 (n21171, n_13011, n_13012);
  not g34509 (n_13434, n21170);
  not g34510 (n_13435, n21171);
  and g34511 (n21172, n_13434, n_13435);
  not g34512 (n_13436, n21169);
  not g34513 (n_13437, n21172);
  and g34514 (n21173, n_13436, n_13437);
  not g34515 (n_13438, n21173);
  and g34516 (n21174, n_13436, n_13438);
  and g34517 (n21175, n_13437, n_13438);
  not g34518 (n_13439, n21174);
  not g34519 (n_13440, n21175);
  and g34520 (n21176, n_13439, n_13440);
  and g34521 (n21177, n20480, n20692);
  not g34522 (n_13441, n21177);
  and g34523 (n21178, n_13006, n_13441);
  and g34524 (n21179, n71, n12531);
  and g34525 (n21180, n9867, n12537);
  and g34526 (n21181, n10434, n12534);
  not g34527 (n_13442, n21180);
  not g34528 (n_13443, n21181);
  and g34529 (n21182, n_13442, n_13443);
  not g34530 (n_13444, n21179);
  and g34531 (n21183, n_13444, n21182);
  and g34532 (n21184, n_4684, n21183);
  and g34533 (n21185, n_9870, n21183);
  not g34534 (n_13445, n21184);
  not g34535 (n_13446, n21185);
  and g34536 (n21186, n_13445, n_13446);
  not g34537 (n_13447, n21186);
  and g34538 (n21187, \a[5] , n_13447);
  and g34539 (n21188, n_3, n21186);
  not g34540 (n_13448, n21187);
  not g34541 (n_13449, n21188);
  and g34542 (n21189, n_13448, n_13449);
  not g34543 (n_13450, n21189);
  and g34544 (n21190, n21178, n_13450);
  and g34545 (n21191, n20498, n20690);
  not g34546 (n_13451, n21191);
  and g34547 (n21192, n_13003, n_13451);
  and g34548 (n21193, n71, n12534);
  and g34549 (n21194, n9867, n12540);
  and g34550 (n21195, n10434, n12537);
  not g34551 (n_13452, n21194);
  not g34552 (n_13453, n21195);
  and g34553 (n21196, n_13452, n_13453);
  not g34554 (n_13454, n21193);
  and g34555 (n21197, n_13454, n21196);
  and g34556 (n21198, n_4684, n21197);
  and g34557 (n21199, n15096, n21197);
  not g34558 (n_13455, n21198);
  not g34559 (n_13456, n21199);
  and g34560 (n21200, n_13455, n_13456);
  not g34561 (n_13457, n21200);
  and g34562 (n21201, \a[5] , n_13457);
  and g34563 (n21202, n_3, n21200);
  not g34564 (n_13458, n21201);
  not g34565 (n_13459, n21202);
  and g34566 (n21203, n_13458, n_13459);
  not g34567 (n_13460, n21203);
  and g34568 (n21204, n21192, n_13460);
  and g34569 (n21205, n20516, n20688);
  not g34570 (n_13461, n21205);
  and g34571 (n21206, n_13000, n_13461);
  and g34572 (n21207, n71, n12537);
  and g34573 (n21208, n9867, n12543);
  and g34574 (n21209, n10434, n12540);
  not g34575 (n_13462, n21208);
  not g34576 (n_13463, n21209);
  and g34577 (n21210, n_13462, n_13463);
  not g34578 (n_13464, n21207);
  and g34579 (n21211, n_13464, n21210);
  and g34580 (n21212, n_4684, n21211);
  and g34581 (n21213, n15385, n21211);
  not g34582 (n_13465, n21212);
  not g34583 (n_13466, n21213);
  and g34584 (n21214, n_13465, n_13466);
  not g34585 (n_13467, n21214);
  and g34586 (n21215, \a[5] , n_13467);
  and g34587 (n21216, n_3, n21214);
  not g34588 (n_13468, n21215);
  not g34589 (n_13469, n21216);
  and g34590 (n21217, n_13468, n_13469);
  not g34591 (n_13470, n21217);
  and g34592 (n21218, n21206, n_13470);
  and g34593 (n21219, n71, n12540);
  and g34594 (n21220, n9867, n12546);
  and g34595 (n21221, n10434, n12543);
  and g34601 (n21224, n9870, n_8936);
  not g34604 (n_13475, n21225);
  and g34605 (n21226, \a[5] , n_13475);
  not g34606 (n_13476, n21226);
  and g34607 (n21227, n_13475, n_13476);
  and g34608 (n21228, \a[5] , n_13476);
  not g34609 (n_13477, n21227);
  not g34610 (n_13478, n21228);
  and g34611 (n21229, n_13477, n_13478);
  not g34612 (n_13479, n20686);
  and g34613 (n21230, n20684, n_13479);
  not g34614 (n_13480, n21230);
  and g34615 (n21231, n_12997, n_13480);
  not g34616 (n_13481, n21229);
  and g34617 (n21232, n_13481, n21231);
  not g34618 (n_13482, n21232);
  and g34619 (n21233, n_13481, n_13482);
  and g34620 (n21234, n21231, n_13482);
  not g34621 (n_13483, n21233);
  not g34622 (n_13484, n21234);
  and g34623 (n21235, n_13483, n_13484);
  and g34624 (n21236, n71, n12543);
  and g34625 (n21237, n9867, n12549);
  and g34626 (n21238, n10434, n12546);
  and g34632 (n21241, n9870, n15724);
  not g34635 (n_13489, n21242);
  and g34636 (n21243, \a[5] , n_13489);
  not g34637 (n_13490, n21243);
  and g34638 (n21244, n_13489, n_13490);
  and g34639 (n21245, \a[5] , n_13490);
  not g34640 (n_13491, n21244);
  not g34641 (n_13492, n21245);
  and g34642 (n21246, n_13491, n_13492);
  and g34643 (n21247, n_12990, n_12992);
  and g34644 (n21248, n_12991, n_12992);
  not g34645 (n_13493, n21247);
  not g34646 (n_13494, n21248);
  and g34647 (n21249, n_13493, n_13494);
  not g34648 (n_13495, n21246);
  not g34649 (n_13496, n21249);
  and g34650 (n21250, n_13495, n_13496);
  not g34651 (n_13497, n21250);
  and g34652 (n21251, n_13495, n_13497);
  and g34653 (n21252, n_13496, n_13497);
  not g34654 (n_13498, n21251);
  not g34655 (n_13499, n21252);
  and g34656 (n21253, n_13498, n_13499);
  and g34657 (n21254, n71, n12546);
  and g34658 (n21255, n9867, n12552);
  and g34659 (n21256, n10434, n12549);
  and g34665 (n21259, n9870, n_8634);
  not g34668 (n_13504, n21260);
  and g34669 (n21261, \a[5] , n_13504);
  not g34670 (n_13505, n21261);
  and g34671 (n21262, n_13504, n_13505);
  and g34672 (n21263, \a[5] , n_13505);
  not g34673 (n_13506, n21262);
  not g34674 (n_13507, n21263);
  and g34675 (n21264, n_13506, n_13507);
  and g34676 (n21265, n_12984, n_12986);
  and g34677 (n21266, n_12985, n_12986);
  not g34678 (n_13508, n21265);
  not g34679 (n_13509, n21266);
  and g34680 (n21267, n_13508, n_13509);
  not g34681 (n_13510, n21264);
  not g34682 (n_13511, n21267);
  and g34683 (n21268, n_13510, n_13511);
  not g34684 (n_13512, n21268);
  and g34685 (n21269, n_13510, n_13512);
  and g34686 (n21270, n_13511, n_13512);
  not g34687 (n_13513, n21269);
  not g34688 (n_13514, n21270);
  and g34689 (n21271, n_13513, n_13514);
  and g34690 (n21272, n20575, n20672);
  not g34691 (n_13515, n21272);
  and g34692 (n21273, n_12980, n_13515);
  and g34693 (n21274, n71, n12549);
  and g34694 (n21275, n9867, n12555);
  and g34695 (n21276, n10434, n12552);
  not g34696 (n_13516, n21275);
  not g34697 (n_13517, n21276);
  and g34698 (n21277, n_13516, n_13517);
  not g34699 (n_13518, n21274);
  and g34700 (n21278, n_13518, n21277);
  and g34701 (n21279, n_4684, n21278);
  and g34702 (n21280, n_9580, n21278);
  not g34703 (n_13519, n21279);
  not g34704 (n_13520, n21280);
  and g34705 (n21281, n_13519, n_13520);
  not g34706 (n_13521, n21281);
  and g34707 (n21282, \a[5] , n_13521);
  and g34708 (n21283, n_3, n21281);
  not g34709 (n_13522, n21282);
  not g34710 (n_13523, n21283);
  and g34711 (n21284, n_13522, n_13523);
  not g34712 (n_13524, n21284);
  and g34713 (n21285, n21273, n_13524);
  not g34714 (n_13525, n20670);
  and g34715 (n21286, n20668, n_13525);
  not g34716 (n_13526, n21286);
  and g34717 (n21287, n_12977, n_13526);
  and g34718 (n21288, n71, n12552);
  and g34719 (n21289, n9867, n12558);
  and g34720 (n21290, n10434, n12555);
  not g34721 (n_13527, n21289);
  not g34722 (n_13528, n21290);
  and g34723 (n21291, n_13527, n_13528);
  not g34724 (n_13529, n21288);
  and g34725 (n21292, n_13529, n21291);
  and g34726 (n21293, n_4684, n21292);
  and g34727 (n21294, n15791, n21292);
  not g34728 (n_13530, n21293);
  not g34729 (n_13531, n21294);
  and g34730 (n21295, n_13530, n_13531);
  not g34731 (n_13532, n21295);
  and g34732 (n21296, \a[5] , n_13532);
  and g34733 (n21297, n_3, n21295);
  not g34734 (n_13533, n21296);
  not g34735 (n_13534, n21297);
  and g34736 (n21298, n_13533, n_13534);
  not g34737 (n_13535, n21298);
  and g34738 (n21299, n21287, n_13535);
  and g34739 (n21300, n20607, n20666);
  not g34740 (n_13536, n21300);
  and g34741 (n21301, n_12973, n_13536);
  and g34742 (n21302, n71, n12555);
  and g34743 (n21303, n9867, n12561);
  and g34744 (n21304, n10434, n12558);
  not g34745 (n_13537, n21303);
  not g34746 (n_13538, n21304);
  and g34747 (n21305, n_13537, n_13538);
  not g34748 (n_13539, n21302);
  and g34749 (n21306, n_13539, n21305);
  and g34750 (n21307, n_4684, n21306);
  and g34751 (n21308, n15816, n21306);
  not g34752 (n_13540, n21307);
  not g34753 (n_13541, n21308);
  and g34754 (n21309, n_13540, n_13541);
  not g34755 (n_13542, n21309);
  and g34756 (n21310, \a[5] , n_13542);
  and g34757 (n21311, n_3, n21309);
  not g34758 (n_13543, n21310);
  not g34759 (n_13544, n21311);
  and g34760 (n21312, n_13543, n_13544);
  not g34761 (n_13545, n21312);
  and g34762 (n21313, n21301, n_13545);
  and g34763 (n21314, n71, n12558);
  and g34764 (n21315, n9867, n12564);
  and g34765 (n21316, n10434, n12561);
  and g34771 (n21319, n9870, n15847);
  not g34774 (n_13550, n21320);
  and g34775 (n21321, \a[5] , n_13550);
  not g34776 (n_13551, n21321);
  and g34777 (n21322, n_13550, n_13551);
  and g34778 (n21323, \a[5] , n_13551);
  not g34779 (n_13552, n21322);
  not g34780 (n_13553, n21323);
  and g34781 (n21324, n_13552, n_13553);
  not g34782 (n_13554, n20664);
  and g34783 (n21325, n20662, n_13554);
  not g34784 (n_13555, n21325);
  and g34785 (n21326, n_12970, n_13555);
  not g34786 (n_13556, n21324);
  and g34787 (n21327, n_13556, n21326);
  not g34788 (n_13557, n21327);
  and g34789 (n21328, n_13556, n_13557);
  and g34790 (n21329, n21326, n_13557);
  not g34791 (n_13558, n21328);
  not g34792 (n_13559, n21329);
  and g34793 (n21330, n_13558, n_13559);
  and g34794 (n21331, n_12963, n_12965);
  and g34795 (n21332, n_12964, n_12965);
  not g34796 (n_13560, n21331);
  not g34797 (n_13561, n21332);
  and g34798 (n21333, n_13560, n_13561);
  and g34799 (n21334, n71, n12561);
  and g34800 (n21335, n9867, n12567);
  and g34801 (n21336, n10434, n12564);
  not g34802 (n_13562, n21335);
  not g34803 (n_13563, n21336);
  and g34804 (n21337, n_13562, n_13563);
  not g34805 (n_13564, n21334);
  and g34806 (n21338, n_13564, n21337);
  and g34807 (n21339, n_4684, n21338);
  and g34808 (n21340, n15905, n21338);
  not g34809 (n_13565, n21339);
  not g34810 (n_13566, n21340);
  and g34811 (n21341, n_13565, n_13566);
  not g34812 (n_13567, n21341);
  and g34813 (n21342, \a[5] , n_13567);
  and g34814 (n21343, n_3, n21341);
  not g34815 (n_13568, n21342);
  not g34816 (n_13569, n21343);
  and g34817 (n21344, n_13568, n_13569);
  not g34818 (n_13570, n21333);
  not g34819 (n_13571, n21344);
  and g34820 (n21345, n_13570, n_13571);
  and g34821 (n21346, n71, n12564);
  and g34822 (n21347, n9867, n12571);
  and g34823 (n21348, n10434, n12567);
  and g34829 (n21351, n9870, n_9006);
  not g34832 (n_13576, n21352);
  and g34833 (n21353, \a[5] , n_13576);
  not g34834 (n_13577, n21353);
  and g34835 (n21354, n_13576, n_13577);
  and g34836 (n21355, \a[5] , n_13577);
  not g34837 (n_13578, n21354);
  not g34838 (n_13579, n21355);
  and g34839 (n21356, n_13578, n_13579);
  not g34840 (n_13580, n20633);
  and g34841 (n21357, n_13580, n20644);
  not g34842 (n_13581, n20645);
  not g34843 (n_13582, n21357);
  and g34844 (n21358, n_13581, n_13582);
  not g34845 (n_13583, n21356);
  and g34846 (n21359, n_13583, n21358);
  not g34847 (n_13584, n21359);
  and g34848 (n21360, n_13583, n_13584);
  and g34849 (n21361, n21358, n_13584);
  not g34850 (n_13585, n21360);
  not g34851 (n_13586, n21361);
  and g34852 (n21362, n_13585, n_13586);
  not g34853 (n_13587, n20632);
  and g34854 (n21363, n20630, n_13587);
  not g34855 (n_13588, n21363);
  and g34856 (n21364, n_13580, n_13588);
  and g34857 (n21365, n71, n12567);
  and g34858 (n21366, n9867, n12574);
  and g34859 (n21367, n10434, n12571);
  not g34860 (n_13589, n21366);
  not g34861 (n_13590, n21367);
  and g34862 (n21368, n_13589, n_13590);
  not g34863 (n_13591, n21365);
  and g34864 (n21369, n_13591, n21368);
  and g34865 (n21370, n_4684, n21369);
  and g34866 (n21371, n_10006, n21369);
  not g34867 (n_13592, n21370);
  not g34868 (n_13593, n21371);
  and g34869 (n21372, n_13592, n_13593);
  not g34870 (n_13594, n21372);
  and g34871 (n21373, \a[5] , n_13594);
  and g34872 (n21374, n_3, n21372);
  not g34873 (n_13595, n21373);
  not g34874 (n_13596, n21374);
  and g34875 (n21375, n_13595, n_13596);
  not g34876 (n_13597, n21375);
  and g34877 (n21376, n21364, n_13597);
  and g34878 (n21377, n10434, n_6977);
  and g34879 (n21378, n71, n12577);
  not g34880 (n_13598, n21377);
  not g34881 (n_13599, n21378);
  and g34882 (n21379, n_13598, n_13599);
  and g34883 (n21380, n9870, n_9032);
  not g34884 (n_13600, n21380);
  and g34885 (n21381, n21379, n_13600);
  not g34886 (n_13601, n21381);
  and g34887 (n21382, \a[5] , n_13601);
  not g34888 (n_13602, n21382);
  and g34889 (n21383, \a[5] , n_13602);
  and g34890 (n21384, n_13601, n_13602);
  not g34891 (n_13603, n21383);
  not g34892 (n_13604, n21384);
  and g34893 (n21385, n_13603, n_13604);
  and g34894 (n21386, n_13, n_6977);
  not g34895 (n_13605, n21386);
  and g34896 (n21387, \a[5] , n_13605);
  not g34897 (n_13606, n21385);
  and g34898 (n21388, n_13606, n21387);
  and g34899 (n21389, n71, n12574);
  and g34900 (n21390, n9867, n_6977);
  and g34901 (n21391, n10434, n12577);
  not g34902 (n_13607, n21390);
  not g34903 (n_13608, n21391);
  and g34904 (n21392, n_13607, n_13608);
  not g34905 (n_13609, n21389);
  and g34906 (n21393, n_13609, n21392);
  and g34907 (n21394, n_4684, n21393);
  and g34908 (n21395, n16094, n21393);
  not g34909 (n_13610, n21394);
  not g34910 (n_13611, n21395);
  and g34911 (n21396, n_13610, n_13611);
  not g34912 (n_13612, n21396);
  and g34913 (n21397, \a[5] , n_13612);
  and g34914 (n21398, n_3, n21396);
  not g34915 (n_13613, n21397);
  not g34916 (n_13614, n21398);
  and g34917 (n21399, n_13613, n_13614);
  not g34918 (n_13615, n21399);
  and g34919 (n21400, n21388, n_13615);
  and g34920 (n21401, n20631, n21400);
  not g34921 (n_13616, n21401);
  and g34922 (n21402, n21400, n_13616);
  and g34923 (n21403, n20631, n_13616);
  not g34924 (n_13617, n21402);
  not g34925 (n_13618, n21403);
  and g34926 (n21404, n_13617, n_13618);
  and g34927 (n21405, n71, n12571);
  and g34928 (n21406, n9867, n12577);
  and g34929 (n21407, n10434, n12574);
  and g34935 (n21410, n9870, n16013);
  not g34938 (n_13623, n21411);
  and g34939 (n21412, \a[5] , n_13623);
  not g34940 (n_13624, n21412);
  and g34941 (n21413, \a[5] , n_13624);
  and g34942 (n21414, n_13623, n_13624);
  not g34943 (n_13625, n21413);
  not g34944 (n_13626, n21414);
  and g34945 (n21415, n_13625, n_13626);
  not g34946 (n_13627, n21404);
  not g34947 (n_13628, n21415);
  and g34948 (n21416, n_13627, n_13628);
  not g34949 (n_13629, n21416);
  and g34950 (n21417, n_13616, n_13629);
  not g34951 (n_13630, n21364);
  and g34952 (n21418, n_13630, n21375);
  not g34953 (n_13631, n21376);
  not g34954 (n_13632, n21418);
  and g34955 (n21419, n_13631, n_13632);
  not g34956 (n_13633, n21417);
  and g34957 (n21420, n_13633, n21419);
  not g34958 (n_13634, n21420);
  and g34959 (n21421, n_13631, n_13634);
  not g34960 (n_13635, n21362);
  not g34961 (n_13636, n21421);
  and g34962 (n21422, n_13635, n_13636);
  not g34963 (n_13637, n21422);
  and g34964 (n21423, n_13584, n_13637);
  and g34965 (n21424, n21333, n21344);
  not g34966 (n_13638, n21345);
  not g34967 (n_13639, n21424);
  and g34968 (n21425, n_13638, n_13639);
  not g34969 (n_13640, n21423);
  and g34970 (n21426, n_13640, n21425);
  not g34971 (n_13641, n21426);
  and g34972 (n21427, n_13638, n_13641);
  not g34973 (n_13642, n21330);
  not g34974 (n_13643, n21427);
  and g34975 (n21428, n_13642, n_13643);
  not g34976 (n_13644, n21428);
  and g34977 (n21429, n_13557, n_13644);
  not g34978 (n_13645, n21313);
  and g34979 (n21430, n21301, n_13645);
  and g34980 (n21431, n_13545, n_13645);
  not g34981 (n_13646, n21430);
  not g34982 (n_13647, n21431);
  and g34983 (n21432, n_13646, n_13647);
  not g34984 (n_13648, n21429);
  not g34985 (n_13649, n21432);
  and g34986 (n21433, n_13648, n_13649);
  not g34987 (n_13650, n21433);
  and g34988 (n21434, n_13645, n_13650);
  not g34989 (n_13651, n21299);
  and g34990 (n21435, n21287, n_13651);
  and g34991 (n21436, n_13535, n_13651);
  not g34992 (n_13652, n21435);
  not g34993 (n_13653, n21436);
  and g34994 (n21437, n_13652, n_13653);
  not g34995 (n_13654, n21434);
  not g34996 (n_13655, n21437);
  and g34997 (n21438, n_13654, n_13655);
  not g34998 (n_13656, n21438);
  and g34999 (n21439, n_13651, n_13656);
  not g35000 (n_13657, n21273);
  and g35001 (n21440, n_13657, n21284);
  not g35002 (n_13658, n21285);
  not g35003 (n_13659, n21440);
  and g35004 (n21441, n_13658, n_13659);
  not g35005 (n_13660, n21439);
  and g35006 (n21442, n_13660, n21441);
  not g35007 (n_13661, n21442);
  and g35008 (n21443, n_13658, n_13661);
  not g35009 (n_13662, n21271);
  not g35010 (n_13663, n21443);
  and g35011 (n21444, n_13662, n_13663);
  not g35012 (n_13664, n21444);
  and g35013 (n21445, n_13512, n_13664);
  not g35014 (n_13665, n21253);
  not g35015 (n_13666, n21445);
  and g35016 (n21446, n_13665, n_13666);
  not g35017 (n_13667, n21446);
  and g35018 (n21447, n_13497, n_13667);
  not g35019 (n_13668, n21235);
  not g35020 (n_13669, n21447);
  and g35021 (n21448, n_13668, n_13669);
  not g35022 (n_13670, n21448);
  and g35023 (n21449, n_13482, n_13670);
  not g35024 (n_13671, n21218);
  and g35025 (n21450, n21206, n_13671);
  and g35026 (n21451, n_13470, n_13671);
  not g35027 (n_13672, n21450);
  not g35028 (n_13673, n21451);
  and g35029 (n21452, n_13672, n_13673);
  not g35030 (n_13674, n21449);
  not g35031 (n_13675, n21452);
  and g35032 (n21453, n_13674, n_13675);
  not g35033 (n_13676, n21453);
  and g35034 (n21454, n_13671, n_13676);
  not g35035 (n_13677, n21204);
  and g35036 (n21455, n21192, n_13677);
  and g35037 (n21456, n_13460, n_13677);
  not g35038 (n_13678, n21455);
  not g35039 (n_13679, n21456);
  and g35040 (n21457, n_13678, n_13679);
  not g35041 (n_13680, n21454);
  not g35042 (n_13681, n21457);
  and g35043 (n21458, n_13680, n_13681);
  not g35044 (n_13682, n21458);
  and g35045 (n21459, n_13677, n_13682);
  not g35046 (n_13683, n21178);
  and g35047 (n21460, n_13683, n21189);
  not g35048 (n_13684, n21190);
  not g35049 (n_13685, n21460);
  and g35050 (n21461, n_13684, n_13685);
  not g35051 (n_13686, n21459);
  and g35052 (n21462, n_13686, n21461);
  not g35053 (n_13687, n21462);
  and g35054 (n21463, n_13684, n_13687);
  not g35055 (n_13688, n21176);
  not g35056 (n_13689, n21463);
  and g35057 (n21464, n_13688, n_13689);
  not g35058 (n_13690, n21464);
  and g35059 (n21465, n_13438, n_13690);
  not g35060 (n_13691, n21158);
  not g35061 (n_13692, n21465);
  and g35062 (n21466, n_13691, n_13692);
  not g35063 (n_13693, n21466);
  and g35064 (n21467, n_13423, n_13693);
  not g35065 (n_13694, n21140);
  not g35066 (n_13695, n21467);
  and g35067 (n21468, n_13694, n_13695);
  not g35068 (n_13696, n21468);
  and g35069 (n21469, n_13408, n_13696);
  not g35070 (n_13697, n21123);
  and g35071 (n21470, n21111, n_13697);
  and g35072 (n21471, n_13396, n_13697);
  not g35073 (n_13698, n21470);
  not g35074 (n_13699, n21471);
  and g35075 (n21472, n_13698, n_13699);
  not g35076 (n_13700, n21469);
  not g35077 (n_13701, n21472);
  and g35078 (n21473, n_13700, n_13701);
  not g35079 (n_13702, n21473);
  and g35080 (n21474, n_13697, n_13702);
  not g35081 (n_13703, n21109);
  and g35082 (n21475, n21097, n_13703);
  and g35083 (n21476, n_13386, n_13703);
  not g35084 (n_13704, n21475);
  not g35085 (n_13705, n21476);
  and g35086 (n21477, n_13704, n_13705);
  not g35087 (n_13706, n21474);
  not g35088 (n_13707, n21477);
  and g35089 (n21478, n_13706, n_13707);
  not g35090 (n_13708, n21478);
  and g35091 (n21479, n_13703, n_13708);
  not g35092 (n_13709, n21083);
  and g35093 (n21480, n_13709, n21094);
  not g35094 (n_13710, n21095);
  not g35095 (n_13711, n21480);
  and g35096 (n21481, n_13710, n_13711);
  not g35097 (n_13712, n21479);
  and g35098 (n21482, n_13712, n21481);
  not g35099 (n_13713, n21482);
  and g35100 (n21483, n_13710, n_13713);
  not g35101 (n_13714, n21081);
  not g35102 (n_13715, n21483);
  and g35103 (n21484, n_13714, n_13715);
  not g35104 (n_13716, n21484);
  and g35105 (n21485, n_13364, n_13716);
  not g35106 (n_13717, n21063);
  not g35107 (n_13718, n21485);
  and g35108 (n21486, n_13717, n_13718);
  not g35109 (n_13719, n21486);
  and g35110 (n21487, n_13349, n_13719);
  not g35111 (n_13720, n21045);
  not g35112 (n_13721, n21487);
  and g35113 (n21488, n_13720, n_13721);
  not g35114 (n_13722, n21488);
  and g35115 (n21489, n_13334, n_13722);
  not g35116 (n_13723, n21028);
  and g35117 (n21490, n21016, n_13723);
  and g35118 (n21491, n_13322, n_13723);
  not g35119 (n_13724, n21490);
  not g35120 (n_13725, n21491);
  and g35121 (n21492, n_13724, n_13725);
  not g35122 (n_13726, n21489);
  not g35123 (n_13727, n21492);
  and g35124 (n21493, n_13726, n_13727);
  not g35125 (n_13728, n21493);
  and g35126 (n21494, n_13723, n_13728);
  not g35127 (n_13729, n21002);
  and g35128 (n21495, n_13729, n21013);
  not g35129 (n_13730, n21014);
  not g35130 (n_13731, n21495);
  and g35131 (n21496, n_13730, n_13731);
  not g35132 (n_13732, n21494);
  and g35133 (n21497, n_13732, n21496);
  not g35134 (n_13733, n21497);
  and g35135 (n21498, n_13730, n_13733);
  not g35136 (n_13734, n21000);
  not g35137 (n_13735, n21498);
  and g35138 (n21499, n_13734, n_13735);
  not g35139 (n_13736, n21499);
  and g35140 (n21500, n_13300, n_13736);
  not g35141 (n_13737, n20982);
  not g35142 (n_13738, n21500);
  and g35143 (n21501, n_13737, n_13738);
  not g35144 (n_13739, n21501);
  and g35145 (n21502, n_13285, n_13739);
  not g35146 (n_13740, n20964);
  not g35147 (n_13741, n21502);
  and g35148 (n21503, n_13740, n_13741);
  not g35149 (n_13742, n21503);
  and g35150 (n21504, n_13270, n_13742);
  not g35151 (n_13743, n20946);
  not g35152 (n_13744, n21504);
  and g35153 (n21505, n_13743, n_13744);
  not g35154 (n_13745, n21505);
  and g35155 (n21506, n_13255, n_13745);
  not g35156 (n_13746, n20928);
  not g35157 (n_13747, n21506);
  and g35158 (n21507, n_13746, n_13747);
  not g35159 (n_13748, n21507);
  and g35160 (n21508, n_13240, n_13748);
  not g35161 (n_13749, n20910);
  not g35162 (n_13750, n21508);
  and g35163 (n21509, n_13749, n_13750);
  not g35164 (n_13751, n21509);
  and g35165 (n21510, n_13225, n_13751);
  not g35166 (n_13752, n20892);
  not g35167 (n_13753, n21510);
  and g35168 (n21511, n_13752, n_13753);
  not g35169 (n_13754, n21511);
  and g35170 (n21512, n_13210, n_13754);
  not g35171 (n_13755, n20874);
  not g35172 (n_13756, n21512);
  and g35173 (n21513, n_13755, n_13756);
  not g35174 (n_13757, n21513);
  and g35175 (n21514, n_13195, n_13757);
  not g35176 (n_13758, n20856);
  not g35177 (n_13759, n21514);
  and g35178 (n21515, n_13758, n_13759);
  not g35179 (n_13760, n21515);
  and g35180 (n21516, n_13180, n_13760);
  not g35181 (n_13761, n20838);
  not g35182 (n_13762, n21516);
  and g35183 (n21517, n_13761, n_13762);
  and g35184 (n21518, n20838, n21516);
  not g35185 (n_13763, n21517);
  not g35186 (n_13764, n21518);
  and g35187 (n21519, n_13763, n_13764);
  and g35188 (n21520, n20856, n21514);
  not g35189 (n_13765, n21520);
  and g35190 (n21521, n_13760, n_13765);
  and g35191 (n21522, n11727, n_7417);
  and g35192 (n21523, n11055, n_7540);
  and g35193 (n21524, n11715, n13941);
  not g35194 (n_13766, n21523);
  not g35195 (n_13767, n21524);
  and g35196 (n21525, n_13766, n_13767);
  not g35197 (n_13768, n21522);
  and g35198 (n21526, n_13768, n21525);
  and g35199 (n21527, n_6291, n21526);
  not g35200 (n_13769, n14028);
  and g35201 (n21528, n_13769, n21526);
  not g35202 (n_13770, n21527);
  not g35203 (n_13771, n21528);
  and g35204 (n21529, n_13770, n_13771);
  not g35205 (n_13772, n21529);
  and g35206 (n21530, \a[2] , n_13772);
  and g35207 (n21531, n_10, n21529);
  not g35208 (n_13773, n21530);
  not g35209 (n_13774, n21531);
  and g35210 (n21532, n_13773, n_13774);
  not g35211 (n_13775, n21532);
  and g35212 (n21533, n21521, n_13775);
  and g35213 (n21534, n20874, n21512);
  not g35214 (n_13776, n21534);
  and g35215 (n21535, n_13757, n_13776);
  and g35216 (n21536, n11727, n13941);
  and g35217 (n21537, n11055, n13633);
  and g35218 (n21538, n11715, n_7540);
  not g35219 (n_13777, n21537);
  not g35220 (n_13778, n21538);
  and g35221 (n21539, n_13777, n_13778);
  not g35222 (n_13779, n21536);
  and g35223 (n21540, n_13779, n21539);
  and g35224 (n21541, n_6291, n21540);
  not g35225 (n_13780, n14136);
  and g35226 (n21542, n_13780, n21540);
  not g35227 (n_13781, n21541);
  not g35228 (n_13782, n21542);
  and g35229 (n21543, n_13781, n_13782);
  not g35230 (n_13783, n21543);
  and g35231 (n21544, \a[2] , n_13783);
  and g35232 (n21545, n_10, n21543);
  not g35233 (n_13784, n21544);
  not g35234 (n_13785, n21545);
  and g35235 (n21546, n_13784, n_13785);
  not g35236 (n_13786, n21546);
  and g35237 (n21547, n21535, n_13786);
  and g35238 (n21548, n20892, n21510);
  not g35239 (n_13787, n21548);
  and g35240 (n21549, n_13754, n_13787);
  and g35241 (n21550, n11727, n_7540);
  and g35242 (n21551, n11055, n13630);
  and g35243 (n21552, n11715, n13633);
  not g35244 (n_13788, n21551);
  not g35245 (n_13789, n21552);
  and g35246 (n21553, n_13788, n_13789);
  not g35247 (n_13790, n21550);
  and g35248 (n21554, n_13790, n21553);
  and g35249 (n21555, n_6291, n21554);
  and g35250 (n21556, n13654, n21554);
  not g35251 (n_13791, n21555);
  not g35252 (n_13792, n21556);
  and g35253 (n21557, n_13791, n_13792);
  not g35254 (n_13793, n21557);
  and g35255 (n21558, \a[2] , n_13793);
  and g35256 (n21559, n_10, n21557);
  not g35257 (n_13794, n21558);
  not g35258 (n_13795, n21559);
  and g35259 (n21560, n_13794, n_13795);
  not g35260 (n_13796, n21560);
  and g35261 (n21561, n21549, n_13796);
  and g35262 (n21562, n20910, n21508);
  not g35263 (n_13797, n21562);
  and g35264 (n21563, n_13751, n_13797);
  and g35265 (n21564, n11727, n13633);
  and g35266 (n21565, n11055, n13597);
  and g35267 (n21566, n11715, n13630);
  not g35268 (n_13798, n21565);
  not g35269 (n_13799, n21566);
  and g35270 (n21567, n_13798, n_13799);
  not g35271 (n_13800, n21564);
  and g35272 (n21568, n_13800, n21567);
  and g35273 (n21569, n_6291, n21568);
  not g35274 (n_13801, n13929);
  and g35275 (n21570, n_13801, n21568);
  not g35276 (n_13802, n21569);
  not g35277 (n_13803, n21570);
  and g35278 (n21571, n_13802, n_13803);
  not g35279 (n_13804, n21571);
  and g35280 (n21572, \a[2] , n_13804);
  and g35281 (n21573, n_10, n21571);
  not g35282 (n_13805, n21572);
  not g35283 (n_13806, n21573);
  and g35284 (n21574, n_13805, n_13806);
  not g35285 (n_13807, n21574);
  and g35286 (n21575, n21563, n_13807);
  and g35287 (n21576, n20928, n21506);
  not g35288 (n_13808, n21576);
  and g35289 (n21577, n_13748, n_13808);
  and g35290 (n21578, n11727, n13630);
  and g35291 (n21579, n11055, n13515);
  and g35292 (n21580, n11715, n13597);
  not g35293 (n_13809, n21579);
  not g35294 (n_13810, n21580);
  and g35295 (n21581, n_13809, n_13810);
  not g35296 (n_13811, n21578);
  and g35297 (n21582, n_13811, n21581);
  and g35298 (n21583, n_6291, n21582);
  not g35299 (n_13812, n13976);
  and g35300 (n21584, n_13812, n21582);
  not g35301 (n_13813, n21583);
  not g35302 (n_13814, n21584);
  and g35303 (n21585, n_13813, n_13814);
  not g35304 (n_13815, n21585);
  and g35305 (n21586, \a[2] , n_13815);
  and g35306 (n21587, n_10, n21585);
  not g35307 (n_13816, n21586);
  not g35308 (n_13817, n21587);
  and g35309 (n21588, n_13816, n_13817);
  not g35310 (n_13818, n21588);
  and g35311 (n21589, n21577, n_13818);
  and g35312 (n21590, n20946, n21504);
  not g35313 (n_13819, n21590);
  and g35314 (n21591, n_13745, n_13819);
  and g35315 (n21592, n11727, n13597);
  and g35316 (n21593, n11055, n13521);
  and g35317 (n21594, n11715, n13515);
  not g35318 (n_13820, n21593);
  not g35319 (n_13821, n21594);
  and g35320 (n21595, n_13820, n_13821);
  not g35321 (n_13822, n21592);
  and g35322 (n21596, n_13822, n21595);
  and g35323 (n21597, n_6291, n21596);
  and g35324 (n21598, n13612, n21596);
  not g35325 (n_13823, n21597);
  not g35326 (n_13824, n21598);
  and g35327 (n21599, n_13823, n_13824);
  not g35328 (n_13825, n21599);
  and g35329 (n21600, \a[2] , n_13825);
  and g35330 (n21601, n_10, n21599);
  not g35331 (n_13826, n21600);
  not g35332 (n_13827, n21601);
  and g35333 (n21602, n_13826, n_13827);
  not g35334 (n_13828, n21602);
  and g35335 (n21603, n21591, n_13828);
  and g35336 (n21604, n20964, n21502);
  not g35337 (n_13829, n21604);
  and g35338 (n21605, n_13742, n_13829);
  and g35339 (n21606, n11727, n13515);
  and g35340 (n21607, n11055, n13518);
  and g35341 (n21608, n11715, n13521);
  not g35342 (n_13830, n21607);
  not g35343 (n_13831, n21608);
  and g35344 (n21609, n_13830, n_13831);
  not g35345 (n_13832, n21606);
  and g35346 (n21610, n_13832, n21609);
  and g35347 (n21611, n_6291, n21610);
  and g35348 (n21612, n_7486, n21610);
  not g35349 (n_13833, n21611);
  not g35350 (n_13834, n21612);
  and g35351 (n21613, n_13833, n_13834);
  not g35352 (n_13835, n21613);
  and g35353 (n21614, \a[2] , n_13835);
  and g35354 (n21615, n_10, n21613);
  not g35355 (n_13836, n21614);
  not g35356 (n_13837, n21615);
  and g35357 (n21616, n_13836, n_13837);
  not g35358 (n_13838, n21616);
  and g35359 (n21617, n21605, n_13838);
  and g35360 (n21618, n20982, n21500);
  not g35361 (n_13839, n21618);
  and g35362 (n21619, n_13739, n_13839);
  and g35363 (n21620, n11727, n13521);
  and g35364 (n21621, n11055, n13491);
  and g35365 (n21622, n11715, n13518);
  not g35366 (n_13840, n21621);
  not g35367 (n_13841, n21622);
  and g35368 (n21623, n_13840, n_13841);
  not g35369 (n_13842, n21620);
  and g35370 (n21624, n_13842, n21623);
  and g35371 (n21625, n_6291, n21624);
  and g35372 (n21626, n13909, n21624);
  not g35373 (n_13843, n21625);
  not g35374 (n_13844, n21626);
  and g35375 (n21627, n_13843, n_13844);
  not g35376 (n_13845, n21627);
  and g35377 (n21628, \a[2] , n_13845);
  and g35378 (n21629, n_10, n21627);
  not g35379 (n_13846, n21628);
  not g35380 (n_13847, n21629);
  and g35381 (n21630, n_13846, n_13847);
  not g35382 (n_13848, n21630);
  and g35383 (n21631, n21619, n_13848);
  and g35384 (n21632, n21000, n21498);
  not g35385 (n_13849, n21632);
  and g35386 (n21633, n_13736, n_13849);
  and g35387 (n21634, n11727, n13518);
  and g35388 (n21635, n11055, n12889);
  and g35389 (n21636, n11715, n13491);
  not g35390 (n_13850, n21635);
  not g35391 (n_13851, n21636);
  and g35392 (n21637, n_13850, n_13851);
  not g35393 (n_13852, n21634);
  and g35394 (n21638, n_13852, n21637);
  and g35395 (n21639, n_6291, n21638);
  and g35396 (n21640, n_12606, n21638);
  not g35397 (n_13853, n21639);
  not g35398 (n_13854, n21640);
  and g35399 (n21641, n_13853, n_13854);
  not g35400 (n_13855, n21641);
  and g35401 (n21642, \a[2] , n_13855);
  and g35402 (n21643, n_10, n21641);
  not g35403 (n_13856, n21642);
  not g35404 (n_13857, n21643);
  and g35405 (n21644, n_13856, n_13857);
  not g35406 (n_13858, n21644);
  and g35407 (n21645, n21633, n_13858);
  not g35408 (n_13859, n21496);
  and g35409 (n21646, n21494, n_13859);
  not g35410 (n_13860, n21646);
  and g35411 (n21647, n_13733, n_13860);
  not g35412 (n_13861, n21481);
  and g35413 (n21648, n21479, n_13861);
  not g35414 (n_13862, n21648);
  and g35415 (n21649, n_13713, n_13862);
  not g35416 (n_13863, n21461);
  and g35417 (n21650, n21459, n_13863);
  not g35418 (n_13864, n21650);
  and g35419 (n21651, n_13687, n_13864);
  not g35420 (n_13865, n21441);
  and g35421 (n21652, n21439, n_13865);
  not g35422 (n_13866, n21652);
  and g35423 (n21653, n_13661, n_13866);
  not g35424 (n_13867, n21419);
  and g35425 (n21654, n21417, n_13867);
  not g35426 (n_13868, n21654);
  and g35427 (n21655, n_13634, n_13868);
  not g35428 (n_13869, n21388);
  and g35429 (n21656, n_13869, n21399);
  not g35430 (n_13870, n21400);
  not g35431 (n_13871, n21656);
  and g35432 (n21657, n_13870, n_13871);
  and g35433 (n21658, n_6354, n_6977);
  and g35434 (n21659, n11796, n_9041);
  and g35435 (n21660, n11727, n12574);
  and g35436 (n21661, n11055, n_6977);
  and g35437 (n21662, n11715, n12577);
  not g35438 (n_13872, n21661);
  not g35439 (n_13873, n21662);
  and g35440 (n21663, n_13872, n_13873);
  not g35441 (n_13874, n21660);
  and g35442 (n21664, n_13874, n21663);
  not g35443 (n_13875, n21664);
  and g35444 (n21665, \a[2] , n_13875);
  and g35445 (n21666, n11796, n_9032);
  and g35446 (n21667, n11805, n_6977);
  and g35447 (n21668, n11807, n12577);
  and g35460 (n21675, n21386, n21674);
  not g35461 (n_13882, n21674);
  and g35462 (n21676, n_13605, n_13882);
  and g35463 (n21677, n11727, n12571);
  and g35464 (n21678, n11055, n12577);
  and g35465 (n21679, n11715, n12574);
  and g35471 (n21682, n11057, n16013);
  not g35474 (n_13887, n21683);
  and g35475 (n21684, n_10, n_13887);
  and g35476 (n21685, \a[2] , n21683);
  not g35477 (n_13888, n21684);
  not g35478 (n_13889, n21685);
  and g35479 (n21686, n_13888, n_13889);
  not g35480 (n_13890, n21676);
  not g35481 (n_13891, n21686);
  and g35482 (n21687, n_13890, n_13891);
  not g35483 (n_13892, n21675);
  not g35484 (n_13893, n21687);
  and g35485 (n21688, n_13892, n_13893);
  and g35486 (n21689, n11727, n12567);
  and g35487 (n21690, n11055, n12574);
  and g35488 (n21691, n11715, n12571);
  not g35489 (n_13894, n21690);
  not g35490 (n_13895, n21691);
  and g35491 (n21692, n_13894, n_13895);
  not g35492 (n_13896, n21689);
  and g35493 (n21693, n_13896, n21692);
  and g35494 (n21694, n_6291, n21693);
  and g35495 (n21695, n_10006, n21693);
  not g35496 (n_13897, n21694);
  not g35497 (n_13898, n21695);
  and g35498 (n21696, n_13897, n_13898);
  not g35499 (n_13899, n21696);
  and g35500 (n21697, \a[2] , n_13899);
  and g35501 (n21698, n_10, n21696);
  not g35502 (n_13900, n21697);
  not g35503 (n_13901, n21698);
  and g35504 (n21699, n_13900, n_13901);
  and g35505 (n21700, n21688, n21699);
  not g35506 (n_13902, n21387);
  and g35507 (n21701, n21385, n_13902);
  not g35508 (n_13903, n21701);
  and g35509 (n21702, n_13869, n_13903);
  not g35510 (n_13904, n21700);
  and g35511 (n21703, n_13904, n21702);
  not g35512 (n_13905, n21688);
  not g35513 (n_13906, n21699);
  and g35514 (n21704, n_13905, n_13906);
  not g35515 (n_13907, n21703);
  not g35516 (n_13908, n21704);
  and g35517 (n21705, n_13907, n_13908);
  not g35518 (n_13909, n21705);
  and g35519 (n21706, n21657, n_13909);
  not g35520 (n_13910, n21657);
  and g35521 (n21707, n_13910, n21705);
  and g35522 (n21708, n11727, n12564);
  and g35523 (n21709, n11055, n12571);
  and g35524 (n21710, n11715, n12567);
  and g35530 (n21713, n11057, n_9006);
  not g35533 (n_13915, n21714);
  and g35534 (n21715, n_10, n_13915);
  and g35535 (n21716, \a[2] , n21714);
  not g35536 (n_13916, n21715);
  not g35537 (n_13917, n21716);
  and g35538 (n21717, n_13916, n_13917);
  not g35539 (n_13918, n21707);
  not g35540 (n_13919, n21717);
  and g35541 (n21718, n_13918, n_13919);
  not g35542 (n_13920, n21706);
  not g35543 (n_13921, n21718);
  and g35544 (n21719, n_13920, n_13921);
  and g35545 (n21720, n11727, n12561);
  and g35546 (n21721, n11055, n12567);
  and g35547 (n21722, n11715, n12564);
  not g35548 (n_13922, n21721);
  not g35549 (n_13923, n21722);
  and g35550 (n21723, n_13922, n_13923);
  not g35551 (n_13924, n21720);
  and g35552 (n21724, n_13924, n21723);
  and g35553 (n21725, n_6291, n21724);
  and g35554 (n21726, n15905, n21724);
  not g35555 (n_13925, n21725);
  not g35556 (n_13926, n21726);
  and g35557 (n21727, n_13925, n_13926);
  not g35558 (n_13927, n21727);
  and g35559 (n21728, \a[2] , n_13927);
  and g35560 (n21729, n_10, n21727);
  not g35561 (n_13928, n21728);
  not g35562 (n_13929, n21729);
  and g35563 (n21730, n_13928, n_13929);
  not g35564 (n_13930, n21719);
  not g35565 (n_13931, n21730);
  and g35566 (n21731, n_13930, n_13931);
  and g35567 (n21732, n21719, n21730);
  and g35568 (n21733, n21404, n21415);
  not g35569 (n_13932, n21733);
  and g35570 (n21734, n_13629, n_13932);
  not g35571 (n_13933, n21732);
  and g35572 (n21735, n_13933, n21734);
  not g35573 (n_13934, n21731);
  not g35574 (n_13935, n21735);
  and g35575 (n21736, n_13934, n_13935);
  not g35576 (n_13936, n21736);
  and g35577 (n21737, n21655, n_13936);
  not g35578 (n_13937, n21655);
  and g35579 (n21738, n_13937, n21736);
  and g35580 (n21739, n11727, n12558);
  and g35581 (n21740, n11055, n12564);
  and g35582 (n21741, n11715, n12561);
  and g35588 (n21744, n11057, n15847);
  not g35591 (n_13942, n21745);
  and g35592 (n21746, n_10, n_13942);
  and g35593 (n21747, \a[2] , n21745);
  not g35594 (n_13943, n21746);
  not g35595 (n_13944, n21747);
  and g35596 (n21748, n_13943, n_13944);
  not g35597 (n_13945, n21738);
  not g35598 (n_13946, n21748);
  and g35599 (n21749, n_13945, n_13946);
  not g35600 (n_13947, n21737);
  not g35601 (n_13948, n21749);
  and g35602 (n21750, n_13947, n_13948);
  and g35603 (n21751, n11727, n12555);
  and g35604 (n21752, n11055, n12561);
  and g35605 (n21753, n11715, n12558);
  not g35606 (n_13949, n21752);
  not g35607 (n_13950, n21753);
  and g35608 (n21754, n_13949, n_13950);
  not g35609 (n_13951, n21751);
  and g35610 (n21755, n_13951, n21754);
  and g35611 (n21756, n_6291, n21755);
  and g35612 (n21757, n15816, n21755);
  not g35613 (n_13952, n21756);
  not g35614 (n_13953, n21757);
  and g35615 (n21758, n_13952, n_13953);
  not g35616 (n_13954, n21758);
  and g35617 (n21759, \a[2] , n_13954);
  and g35618 (n21760, n_10, n21758);
  not g35619 (n_13955, n21759);
  not g35620 (n_13956, n21760);
  and g35621 (n21761, n_13955, n_13956);
  and g35622 (n21762, n21750, n21761);
  and g35623 (n21763, n21362, n21421);
  not g35624 (n_13957, n21763);
  and g35625 (n21764, n_13637, n_13957);
  not g35626 (n_13958, n21762);
  and g35627 (n21765, n_13958, n21764);
  not g35628 (n_13959, n21750);
  not g35629 (n_13960, n21761);
  and g35630 (n21766, n_13959, n_13960);
  not g35631 (n_13961, n21765);
  not g35632 (n_13962, n21766);
  and g35633 (n21767, n_13961, n_13962);
  and g35634 (n21768, n11727, n12552);
  and g35635 (n21769, n11055, n12558);
  and g35636 (n21770, n11715, n12555);
  not g35637 (n_13963, n21769);
  not g35638 (n_13964, n21770);
  and g35639 (n21771, n_13963, n_13964);
  not g35640 (n_13965, n21768);
  and g35641 (n21772, n_13965, n21771);
  and g35642 (n21773, n_6291, n21772);
  and g35643 (n21774, n15791, n21772);
  not g35644 (n_13966, n21773);
  not g35645 (n_13967, n21774);
  and g35646 (n21775, n_13966, n_13967);
  not g35647 (n_13968, n21775);
  and g35648 (n21776, \a[2] , n_13968);
  and g35649 (n21777, n_10, n21775);
  not g35650 (n_13969, n21776);
  not g35651 (n_13970, n21777);
  and g35652 (n21778, n_13969, n_13970);
  and g35653 (n21779, n21767, n21778);
  not g35654 (n_13971, n21425);
  and g35655 (n21780, n21423, n_13971);
  not g35656 (n_13972, n21780);
  and g35657 (n21781, n_13641, n_13972);
  not g35658 (n_13973, n21779);
  and g35659 (n21782, n_13973, n21781);
  not g35660 (n_13974, n21767);
  not g35661 (n_13975, n21778);
  and g35662 (n21783, n_13974, n_13975);
  not g35663 (n_13976, n21782);
  not g35664 (n_13977, n21783);
  and g35665 (n21784, n_13976, n_13977);
  and g35666 (n21785, n11727, n12549);
  and g35667 (n21786, n11055, n12555);
  and g35668 (n21787, n11715, n12552);
  not g35669 (n_13978, n21786);
  not g35670 (n_13979, n21787);
  and g35671 (n21788, n_13978, n_13979);
  not g35672 (n_13980, n21785);
  and g35673 (n21789, n_13980, n21788);
  and g35674 (n21790, n_6291, n21789);
  and g35675 (n21791, n_9580, n21789);
  not g35676 (n_13981, n21790);
  not g35677 (n_13982, n21791);
  and g35678 (n21792, n_13981, n_13982);
  not g35679 (n_13983, n21792);
  and g35680 (n21793, \a[2] , n_13983);
  and g35681 (n21794, n_10, n21792);
  not g35682 (n_13984, n21793);
  not g35683 (n_13985, n21794);
  and g35684 (n21795, n_13984, n_13985);
  and g35685 (n21796, n21784, n21795);
  and g35686 (n21797, n21330, n21427);
  not g35687 (n_13986, n21797);
  and g35688 (n21798, n_13644, n_13986);
  not g35689 (n_13987, n21796);
  and g35690 (n21799, n_13987, n21798);
  not g35691 (n_13988, n21784);
  not g35692 (n_13989, n21795);
  and g35693 (n21800, n_13988, n_13989);
  not g35694 (n_13990, n21799);
  not g35695 (n_13991, n21800);
  and g35696 (n21801, n_13990, n_13991);
  and g35697 (n21802, n21429, n_13647);
  and g35698 (n21803, n_13646, n21802);
  not g35699 (n_13992, n21803);
  and g35700 (n21804, n_13650, n_13992);
  not g35701 (n_13993, n21801);
  and g35702 (n21805, n_13993, n21804);
  not g35703 (n_13994, n21804);
  and g35704 (n21806, n21801, n_13994);
  and g35705 (n21807, n11727, n12546);
  and g35706 (n21808, n11055, n12552);
  and g35707 (n21809, n11715, n12549);
  and g35713 (n21812, n11057, n_8634);
  not g35716 (n_13999, n21813);
  and g35717 (n21814, n_10, n_13999);
  and g35718 (n21815, \a[2] , n21813);
  not g35719 (n_14000, n21814);
  not g35720 (n_14001, n21815);
  and g35721 (n21816, n_14000, n_14001);
  not g35722 (n_14002, n21806);
  not g35723 (n_14003, n21816);
  and g35724 (n21817, n_14002, n_14003);
  not g35725 (n_14004, n21805);
  not g35726 (n_14005, n21817);
  and g35727 (n21818, n_14004, n_14005);
  and g35728 (n21819, n21434, n_13653);
  and g35729 (n21820, n_13652, n21819);
  not g35730 (n_14006, n21820);
  and g35731 (n21821, n_13656, n_14006);
  not g35732 (n_14007, n21818);
  and g35733 (n21822, n_14007, n21821);
  not g35734 (n_14008, n21821);
  and g35735 (n21823, n21818, n_14008);
  and g35736 (n21824, n11727, n12543);
  and g35737 (n21825, n11055, n12549);
  and g35738 (n21826, n11715, n12546);
  and g35744 (n21829, n11057, n15724);
  not g35747 (n_14013, n21830);
  and g35748 (n21831, n_10, n_14013);
  and g35749 (n21832, \a[2] , n21830);
  not g35750 (n_14014, n21831);
  not g35751 (n_14015, n21832);
  and g35752 (n21833, n_14014, n_14015);
  not g35753 (n_14016, n21823);
  not g35754 (n_14017, n21833);
  and g35755 (n21834, n_14016, n_14017);
  not g35756 (n_14018, n21822);
  not g35757 (n_14019, n21834);
  and g35758 (n21835, n_14018, n_14019);
  not g35759 (n_14020, n21835);
  and g35760 (n21836, n21653, n_14020);
  not g35761 (n_14021, n21653);
  and g35762 (n21837, n_14021, n21835);
  and g35763 (n21838, n11727, n12540);
  and g35764 (n21839, n11055, n12546);
  and g35765 (n21840, n11715, n12543);
  and g35771 (n21843, n11057, n_8936);
  not g35774 (n_14026, n21844);
  and g35775 (n21845, n_10, n_14026);
  and g35776 (n21846, \a[2] , n21844);
  not g35777 (n_14027, n21845);
  not g35778 (n_14028, n21846);
  and g35779 (n21847, n_14027, n_14028);
  not g35780 (n_14029, n21837);
  not g35781 (n_14030, n21847);
  and g35782 (n21848, n_14029, n_14030);
  not g35783 (n_14031, n21836);
  not g35784 (n_14032, n21848);
  and g35785 (n21849, n_14031, n_14032);
  and g35786 (n21850, n11727, n12537);
  and g35787 (n21851, n11055, n12543);
  and g35788 (n21852, n11715, n12540);
  not g35789 (n_14033, n21851);
  not g35790 (n_14034, n21852);
  and g35791 (n21853, n_14033, n_14034);
  not g35792 (n_14035, n21850);
  and g35793 (n21854, n_14035, n21853);
  and g35794 (n21855, n_6291, n21854);
  and g35795 (n21856, n15385, n21854);
  not g35796 (n_14036, n21855);
  not g35797 (n_14037, n21856);
  and g35798 (n21857, n_14036, n_14037);
  not g35799 (n_14038, n21857);
  and g35800 (n21858, \a[2] , n_14038);
  and g35801 (n21859, n_10, n21857);
  not g35802 (n_14039, n21858);
  not g35803 (n_14040, n21859);
  and g35804 (n21860, n_14039, n_14040);
  and g35805 (n21861, n21849, n21860);
  and g35806 (n21862, n21271, n21443);
  not g35807 (n_14041, n21862);
  and g35808 (n21863, n_13664, n_14041);
  not g35809 (n_14042, n21861);
  and g35810 (n21864, n_14042, n21863);
  not g35811 (n_14043, n21849);
  not g35812 (n_14044, n21860);
  and g35813 (n21865, n_14043, n_14044);
  not g35814 (n_14045, n21864);
  not g35815 (n_14046, n21865);
  and g35816 (n21866, n_14045, n_14046);
  and g35817 (n21867, n11727, n12534);
  and g35818 (n21868, n11055, n12540);
  and g35819 (n21869, n11715, n12537);
  not g35820 (n_14047, n21868);
  not g35821 (n_14048, n21869);
  and g35822 (n21870, n_14047, n_14048);
  not g35823 (n_14049, n21867);
  and g35824 (n21871, n_14049, n21870);
  and g35825 (n21872, n_6291, n21871);
  and g35826 (n21873, n15096, n21871);
  not g35827 (n_14050, n21872);
  not g35828 (n_14051, n21873);
  and g35829 (n21874, n_14050, n_14051);
  not g35830 (n_14052, n21874);
  and g35831 (n21875, \a[2] , n_14052);
  and g35832 (n21876, n_10, n21874);
  not g35833 (n_14053, n21875);
  not g35834 (n_14054, n21876);
  and g35835 (n21877, n_14053, n_14054);
  and g35836 (n21878, n21866, n21877);
  and g35837 (n21879, n21253, n21445);
  not g35838 (n_14055, n21879);
  and g35839 (n21880, n_13667, n_14055);
  not g35840 (n_14056, n21878);
  and g35841 (n21881, n_14056, n21880);
  not g35842 (n_14057, n21866);
  not g35843 (n_14058, n21877);
  and g35844 (n21882, n_14057, n_14058);
  not g35845 (n_14059, n21881);
  not g35846 (n_14060, n21882);
  and g35847 (n21883, n_14059, n_14060);
  and g35848 (n21884, n11727, n12531);
  and g35849 (n21885, n11055, n12537);
  and g35850 (n21886, n11715, n12534);
  not g35851 (n_14061, n21885);
  not g35852 (n_14062, n21886);
  and g35853 (n21887, n_14061, n_14062);
  not g35854 (n_14063, n21884);
  and g35855 (n21888, n_14063, n21887);
  and g35856 (n21889, n_6291, n21888);
  and g35857 (n21890, n_9870, n21888);
  not g35858 (n_14064, n21889);
  not g35859 (n_14065, n21890);
  and g35860 (n21891, n_14064, n_14065);
  not g35861 (n_14066, n21891);
  and g35862 (n21892, \a[2] , n_14066);
  and g35863 (n21893, n_10, n21891);
  not g35864 (n_14067, n21892);
  not g35865 (n_14068, n21893);
  and g35866 (n21894, n_14067, n_14068);
  and g35867 (n21895, n21883, n21894);
  and g35868 (n21896, n21235, n21447);
  not g35869 (n_14069, n21896);
  and g35870 (n21897, n_13670, n_14069);
  not g35871 (n_14070, n21895);
  and g35872 (n21898, n_14070, n21897);
  not g35873 (n_14071, n21883);
  not g35874 (n_14072, n21894);
  and g35875 (n21899, n_14071, n_14072);
  not g35876 (n_14073, n21898);
  not g35877 (n_14074, n21899);
  and g35878 (n21900, n_14073, n_14074);
  and g35879 (n21901, n21449, n_13673);
  and g35880 (n21902, n_13672, n21901);
  not g35881 (n_14075, n21902);
  and g35882 (n21903, n_13676, n_14075);
  not g35883 (n_14076, n21900);
  and g35884 (n21904, n_14076, n21903);
  not g35885 (n_14077, n21903);
  and g35886 (n21905, n21900, n_14077);
  and g35887 (n21906, n11727, n12528);
  and g35888 (n21907, n11055, n12534);
  and g35889 (n21908, n11715, n12531);
  and g35895 (n21911, n11057, n_8448);
  not g35898 (n_14082, n21912);
  and g35899 (n21913, n_10, n_14082);
  and g35900 (n21914, \a[2] , n21912);
  not g35901 (n_14083, n21913);
  not g35902 (n_14084, n21914);
  and g35903 (n21915, n_14083, n_14084);
  not g35904 (n_14085, n21905);
  not g35905 (n_14086, n21915);
  and g35906 (n21916, n_14085, n_14086);
  not g35907 (n_14087, n21904);
  not g35908 (n_14088, n21916);
  and g35909 (n21917, n_14087, n_14088);
  and g35910 (n21918, n21454, n_13679);
  and g35911 (n21919, n_13678, n21918);
  not g35912 (n_14089, n21919);
  and g35913 (n21920, n_13682, n_14089);
  not g35914 (n_14090, n21917);
  and g35915 (n21921, n_14090, n21920);
  not g35916 (n_14091, n21920);
  and g35917 (n21922, n21917, n_14091);
  and g35918 (n21923, n11727, n12525);
  and g35919 (n21924, n11055, n12531);
  and g35920 (n21925, n11715, n12528);
  and g35926 (n21928, n11057, n14608);
  not g35929 (n_14096, n21929);
  and g35930 (n21930, n_10, n_14096);
  and g35931 (n21931, \a[2] , n21929);
  not g35932 (n_14097, n21930);
  not g35933 (n_14098, n21931);
  and g35934 (n21932, n_14097, n_14098);
  not g35935 (n_14099, n21922);
  not g35936 (n_14100, n21932);
  and g35937 (n21933, n_14099, n_14100);
  not g35938 (n_14101, n21921);
  not g35939 (n_14102, n21933);
  and g35940 (n21934, n_14101, n_14102);
  not g35941 (n_14103, n21934);
  and g35942 (n21935, n21651, n_14103);
  not g35943 (n_14104, n21651);
  and g35944 (n21936, n_14104, n21934);
  and g35945 (n21937, n11727, n12522);
  and g35946 (n21938, n11055, n12528);
  and g35947 (n21939, n11715, n12525);
  and g35953 (n21942, n11057, n14837);
  not g35956 (n_14109, n21943);
  and g35957 (n21944, n_10, n_14109);
  and g35958 (n21945, \a[2] , n21943);
  not g35959 (n_14110, n21944);
  not g35960 (n_14111, n21945);
  and g35961 (n21946, n_14110, n_14111);
  not g35962 (n_14112, n21936);
  not g35963 (n_14113, n21946);
  and g35964 (n21947, n_14112, n_14113);
  not g35965 (n_14114, n21935);
  not g35966 (n_14115, n21947);
  and g35967 (n21948, n_14114, n_14115);
  and g35968 (n21949, n11727, n12519);
  and g35969 (n21950, n11055, n12525);
  and g35970 (n21951, n11715, n12522);
  not g35971 (n_14116, n21950);
  not g35972 (n_14117, n21951);
  and g35973 (n21952, n_14116, n_14117);
  not g35974 (n_14118, n21949);
  and g35975 (n21953, n_14118, n21952);
  and g35976 (n21954, n_6291, n21953);
  and g35977 (n21955, n_10664, n21953);
  not g35978 (n_14119, n21954);
  not g35979 (n_14120, n21955);
  and g35980 (n21956, n_14119, n_14120);
  not g35981 (n_14121, n21956);
  and g35982 (n21957, \a[2] , n_14121);
  and g35983 (n21958, n_10, n21956);
  not g35984 (n_14122, n21957);
  not g35985 (n_14123, n21958);
  and g35986 (n21959, n_14122, n_14123);
  and g35987 (n21960, n21948, n21959);
  and g35988 (n21961, n21176, n21463);
  not g35989 (n_14124, n21961);
  and g35990 (n21962, n_13690, n_14124);
  not g35991 (n_14125, n21960);
  and g35992 (n21963, n_14125, n21962);
  not g35993 (n_14126, n21948);
  not g35994 (n_14127, n21959);
  and g35995 (n21964, n_14126, n_14127);
  not g35996 (n_14128, n21963);
  not g35997 (n_14129, n21964);
  and g35998 (n21965, n_14128, n_14129);
  and g35999 (n21966, n11727, n12516);
  and g36000 (n21967, n11055, n12522);
  and g36001 (n21968, n11715, n12519);
  not g36002 (n_14130, n21967);
  not g36003 (n_14131, n21968);
  and g36004 (n21969, n_14130, n_14131);
  not g36005 (n_14132, n21966);
  and g36006 (n21970, n_14132, n21969);
  and g36007 (n21971, n_6291, n21970);
  and g36008 (n21972, n14443, n21970);
  not g36009 (n_14133, n21971);
  not g36010 (n_14134, n21972);
  and g36011 (n21973, n_14133, n_14134);
  not g36012 (n_14135, n21973);
  and g36013 (n21974, \a[2] , n_14135);
  and g36014 (n21975, n_10, n21973);
  not g36015 (n_14136, n21974);
  not g36016 (n_14137, n21975);
  and g36017 (n21976, n_14136, n_14137);
  and g36018 (n21977, n21965, n21976);
  and g36019 (n21978, n21158, n21465);
  not g36020 (n_14138, n21978);
  and g36021 (n21979, n_13693, n_14138);
  not g36022 (n_14139, n21977);
  and g36023 (n21980, n_14139, n21979);
  not g36024 (n_14140, n21965);
  not g36025 (n_14141, n21976);
  and g36026 (n21981, n_14140, n_14141);
  not g36027 (n_14142, n21980);
  not g36028 (n_14143, n21981);
  and g36029 (n21982, n_14142, n_14143);
  and g36030 (n21983, n11727, n12511);
  and g36031 (n21984, n11055, n12519);
  and g36032 (n21985, n11715, n12516);
  not g36033 (n_14144, n21984);
  not g36034 (n_14145, n21985);
  and g36035 (n21986, n_14144, n_14145);
  not g36036 (n_14146, n21983);
  and g36037 (n21987, n_14146, n21986);
  and g36038 (n21988, n_6291, n21987);
  and g36039 (n21989, n14233, n21987);
  not g36040 (n_14147, n21988);
  not g36041 (n_14148, n21989);
  and g36042 (n21990, n_14147, n_14148);
  not g36043 (n_14149, n21990);
  and g36044 (n21991, \a[2] , n_14149);
  and g36045 (n21992, n_10, n21990);
  not g36046 (n_14150, n21991);
  not g36047 (n_14151, n21992);
  and g36048 (n21993, n_14150, n_14151);
  and g36049 (n21994, n21982, n21993);
  and g36050 (n21995, n21140, n21467);
  not g36051 (n_14152, n21995);
  and g36052 (n21996, n_13696, n_14152);
  not g36053 (n_14153, n21994);
  and g36054 (n21997, n_14153, n21996);
  not g36055 (n_14154, n21982);
  not g36056 (n_14155, n21993);
  and g36057 (n21998, n_14154, n_14155);
  not g36058 (n_14156, n21997);
  not g36059 (n_14157, n21998);
  and g36060 (n21999, n_14156, n_14157);
  and g36061 (n22000, n21469, n_13699);
  and g36062 (n22001, n_13698, n22000);
  not g36063 (n_14158, n22001);
  and g36064 (n22002, n_13702, n_14158);
  not g36065 (n_14159, n21999);
  and g36066 (n22003, n_14159, n22002);
  not g36067 (n_14160, n22002);
  and g36068 (n22004, n21999, n_14160);
  and g36069 (n22005, n11727, n12513);
  and g36070 (n22006, n11055, n12516);
  and g36071 (n22007, n11715, n12511);
  and g36077 (n22010, n11057, n14177);
  not g36080 (n_14165, n22011);
  and g36081 (n22012, n_10, n_14165);
  and g36082 (n22013, \a[2] , n22011);
  not g36083 (n_14166, n22012);
  not g36084 (n_14167, n22013);
  and g36085 (n22014, n_14166, n_14167);
  not g36086 (n_14168, n22004);
  not g36087 (n_14169, n22014);
  and g36088 (n22015, n_14168, n_14169);
  not g36089 (n_14170, n22003);
  not g36090 (n_14171, n22015);
  and g36091 (n22016, n_14170, n_14171);
  and g36092 (n22017, n21474, n_13705);
  and g36093 (n22018, n_13704, n22017);
  not g36094 (n_14172, n22018);
  and g36095 (n22019, n_13708, n_14172);
  not g36096 (n_14173, n22016);
  and g36097 (n22020, n_14173, n22019);
  not g36098 (n_14174, n22019);
  and g36099 (n22021, n22016, n_14174);
  and g36100 (n22022, n11727, n12508);
  and g36101 (n22023, n11055, n12511);
  and g36102 (n22024, n11715, n12513);
  and g36108 (n22027, n11057, n13863);
  not g36111 (n_14179, n22028);
  and g36112 (n22029, n_10, n_14179);
  and g36113 (n22030, \a[2] , n22028);
  not g36114 (n_14180, n22029);
  not g36115 (n_14181, n22030);
  and g36116 (n22031, n_14180, n_14181);
  not g36117 (n_14182, n22021);
  not g36118 (n_14183, n22031);
  and g36119 (n22032, n_14182, n_14183);
  not g36120 (n_14184, n22020);
  not g36121 (n_14185, n22032);
  and g36122 (n22033, n_14184, n_14185);
  not g36123 (n_14186, n22033);
  and g36124 (n22034, n21649, n_14186);
  not g36125 (n_14187, n21649);
  and g36126 (n22035, n_14187, n22033);
  and g36127 (n22036, n11727, n12505);
  and g36128 (n22037, n11055, n12513);
  and g36129 (n22038, n11715, n12508);
  and g36135 (n22041, n11057, n_7804);
  not g36138 (n_14192, n22042);
  and g36139 (n22043, n_10, n_14192);
  and g36140 (n22044, \a[2] , n22042);
  not g36141 (n_14193, n22043);
  not g36142 (n_14194, n22044);
  and g36143 (n22045, n_14193, n_14194);
  not g36144 (n_14195, n22035);
  not g36145 (n_14196, n22045);
  and g36146 (n22046, n_14195, n_14196);
  not g36147 (n_14197, n22034);
  not g36148 (n_14198, n22046);
  and g36149 (n22047, n_14197, n_14198);
  and g36150 (n22048, n11727, n12370);
  and g36151 (n22049, n11055, n12508);
  and g36152 (n22050, n11715, n12505);
  not g36153 (n_14199, n22049);
  not g36154 (n_14200, n22050);
  and g36155 (n22051, n_14199, n_14200);
  not g36156 (n_14201, n22048);
  and g36157 (n22052, n_14201, n22051);
  and g36158 (n22053, n_6291, n22052);
  and g36159 (n22054, n13748, n22052);
  not g36160 (n_14202, n22053);
  not g36161 (n_14203, n22054);
  and g36162 (n22055, n_14202, n_14203);
  not g36163 (n_14204, n22055);
  and g36164 (n22056, \a[2] , n_14204);
  and g36165 (n22057, n_10, n22055);
  not g36166 (n_14205, n22056);
  not g36167 (n_14206, n22057);
  and g36168 (n22058, n_14205, n_14206);
  and g36169 (n22059, n22047, n22058);
  and g36170 (n22060, n21081, n21483);
  not g36171 (n_14207, n22060);
  and g36172 (n22061, n_13716, n_14207);
  not g36173 (n_14208, n22059);
  and g36174 (n22062, n_14208, n22061);
  not g36175 (n_14209, n22047);
  not g36176 (n_14210, n22058);
  and g36177 (n22063, n_14209, n_14210);
  not g36178 (n_14211, n22062);
  not g36179 (n_14212, n22063);
  and g36180 (n22064, n_14211, n_14212);
  and g36181 (n22065, n11727, n12502);
  and g36182 (n22066, n11055, n12505);
  and g36183 (n22067, n11715, n12370);
  not g36184 (n_14213, n22066);
  not g36185 (n_14214, n22067);
  and g36186 (n22068, n_14213, n_14214);
  not g36187 (n_14215, n22065);
  and g36188 (n22069, n_14215, n22068);
  and g36189 (n22070, n_6291, n22069);
  and g36190 (n22071, n13736, n22069);
  not g36191 (n_14216, n22070);
  not g36192 (n_14217, n22071);
  and g36193 (n22072, n_14216, n_14217);
  not g36194 (n_14218, n22072);
  and g36195 (n22073, \a[2] , n_14218);
  and g36196 (n22074, n_10, n22072);
  not g36197 (n_14219, n22073);
  not g36198 (n_14220, n22074);
  and g36199 (n22075, n_14219, n_14220);
  and g36200 (n22076, n22064, n22075);
  and g36201 (n22077, n21063, n21485);
  not g36202 (n_14221, n22077);
  and g36203 (n22078, n_13719, n_14221);
  not g36204 (n_14222, n22076);
  and g36205 (n22079, n_14222, n22078);
  not g36206 (n_14223, n22064);
  not g36207 (n_14224, n22075);
  and g36208 (n22080, n_14223, n_14224);
  not g36209 (n_14225, n22079);
  not g36210 (n_14226, n22080);
  and g36211 (n22081, n_14225, n_14226);
  and g36212 (n22082, n11727, n12769);
  and g36213 (n22083, n11055, n12370);
  and g36214 (n22084, n11715, n12502);
  not g36215 (n_14227, n22083);
  not g36216 (n_14228, n22084);
  and g36217 (n22085, n_14227, n_14228);
  not g36218 (n_14229, n22082);
  and g36219 (n22086, n_14229, n22085);
  and g36220 (n22087, n_6291, n22086);
  and g36221 (n22088, n_7817, n22086);
  not g36222 (n_14230, n22087);
  not g36223 (n_14231, n22088);
  and g36224 (n22089, n_14230, n_14231);
  not g36225 (n_14232, n22089);
  and g36226 (n22090, \a[2] , n_14232);
  and g36227 (n22091, n_10, n22089);
  not g36228 (n_14233, n22090);
  not g36229 (n_14234, n22091);
  and g36230 (n22092, n_14233, n_14234);
  and g36231 (n22093, n22081, n22092);
  and g36232 (n22094, n21045, n21487);
  not g36233 (n_14235, n22094);
  and g36234 (n22095, n_13722, n_14235);
  not g36235 (n_14236, n22093);
  and g36236 (n22096, n_14236, n22095);
  not g36237 (n_14237, n22081);
  not g36238 (n_14238, n22092);
  and g36239 (n22097, n_14237, n_14238);
  not g36240 (n_14239, n22096);
  not g36241 (n_14240, n22097);
  and g36242 (n22098, n_14239, n_14240);
  and g36243 (n22099, n21489, n_13725);
  and g36244 (n22100, n_13724, n22099);
  not g36245 (n_14241, n22100);
  and g36246 (n22101, n_13728, n_14241);
  not g36247 (n_14242, n22098);
  and g36248 (n22102, n_14242, n22101);
  not g36249 (n_14243, n22101);
  and g36250 (n22103, n22098, n_14243);
  and g36251 (n22104, n11727, n12889);
  and g36252 (n22105, n11055, n12502);
  and g36253 (n22106, n11715, n12769);
  and g36259 (n22109, n11057, n12895);
  not g36262 (n_14248, n22110);
  and g36263 (n22111, n_10, n_14248);
  and g36264 (n22112, \a[2] , n22110);
  not g36265 (n_14249, n22111);
  not g36266 (n_14250, n22112);
  and g36267 (n22113, n_14249, n_14250);
  not g36268 (n_14251, n22103);
  not g36269 (n_14252, n22113);
  and g36270 (n22114, n_14251, n_14252);
  not g36271 (n_14253, n22102);
  not g36272 (n_14254, n22114);
  and g36273 (n22115, n_14253, n_14254);
  not g36274 (n_14255, n22115);
  and g36275 (n22116, n21647, n_14255);
  not g36276 (n_14256, n21647);
  and g36277 (n22117, n_14256, n22115);
  and g36278 (n22118, n11727, n13491);
  and g36279 (n22119, n11055, n12769);
  and g36280 (n22120, n11715, n12889);
  and g36286 (n22123, n11057, n_7447);
  not g36289 (n_14261, n22124);
  and g36290 (n22125, n_10, n_14261);
  and g36291 (n22126, \a[2] , n22124);
  not g36292 (n_14262, n22125);
  not g36293 (n_14263, n22126);
  and g36294 (n22127, n_14262, n_14263);
  not g36295 (n_14264, n22117);
  not g36296 (n_14265, n22127);
  and g36297 (n22128, n_14264, n_14265);
  not g36298 (n_14266, n22116);
  not g36299 (n_14267, n22128);
  and g36300 (n22129, n_14266, n_14267);
  not g36301 (n_14268, n21645);
  and g36302 (n22130, n21633, n_14268);
  and g36303 (n22131, n_13858, n_14268);
  not g36304 (n_14269, n22130);
  not g36305 (n_14270, n22131);
  and g36306 (n22132, n_14269, n_14270);
  not g36307 (n_14271, n22129);
  not g36308 (n_14272, n22132);
  and g36309 (n22133, n_14271, n_14272);
  not g36310 (n_14273, n22133);
  and g36311 (n22134, n_14268, n_14273);
  not g36312 (n_14274, n21619);
  and g36313 (n22135, n_14274, n21630);
  not g36314 (n_14275, n21631);
  not g36315 (n_14276, n22135);
  and g36316 (n22136, n_14275, n_14276);
  not g36317 (n_14277, n22134);
  and g36318 (n22137, n_14277, n22136);
  not g36319 (n_14278, n22137);
  and g36320 (n22138, n_14275, n_14278);
  not g36321 (n_14279, n21605);
  and g36322 (n22139, n_14279, n21616);
  not g36323 (n_14280, n21617);
  not g36324 (n_14281, n22139);
  and g36325 (n22140, n_14280, n_14281);
  not g36326 (n_14282, n22138);
  and g36327 (n22141, n_14282, n22140);
  not g36328 (n_14283, n22141);
  and g36329 (n22142, n_14280, n_14283);
  not g36330 (n_14284, n21591);
  and g36331 (n22143, n_14284, n21602);
  not g36332 (n_14285, n21603);
  not g36333 (n_14286, n22143);
  and g36334 (n22144, n_14285, n_14286);
  not g36335 (n_14287, n22142);
  and g36336 (n22145, n_14287, n22144);
  not g36337 (n_14288, n22145);
  and g36338 (n22146, n_14285, n_14288);
  not g36339 (n_14289, n21577);
  and g36340 (n22147, n_14289, n21588);
  not g36341 (n_14290, n21589);
  not g36342 (n_14291, n22147);
  and g36343 (n22148, n_14290, n_14291);
  not g36344 (n_14292, n22146);
  and g36345 (n22149, n_14292, n22148);
  not g36346 (n_14293, n22149);
  and g36347 (n22150, n_14290, n_14293);
  not g36348 (n_14294, n21563);
  and g36349 (n22151, n_14294, n21574);
  not g36350 (n_14295, n21575);
  not g36351 (n_14296, n22151);
  and g36352 (n22152, n_14295, n_14296);
  not g36353 (n_14297, n22150);
  and g36354 (n22153, n_14297, n22152);
  not g36355 (n_14298, n22153);
  and g36356 (n22154, n_14295, n_14298);
  not g36357 (n_14299, n21549);
  and g36358 (n22155, n_14299, n21560);
  not g36359 (n_14300, n21561);
  not g36360 (n_14301, n22155);
  and g36361 (n22156, n_14300, n_14301);
  not g36362 (n_14302, n22154);
  and g36363 (n22157, n_14302, n22156);
  not g36364 (n_14303, n22157);
  and g36365 (n22158, n_14300, n_14303);
  not g36366 (n_14304, n21535);
  and g36367 (n22159, n_14304, n21546);
  not g36368 (n_14305, n21547);
  not g36369 (n_14306, n22159);
  and g36370 (n22160, n_14305, n_14306);
  not g36371 (n_14307, n22158);
  and g36372 (n22161, n_14307, n22160);
  not g36373 (n_14308, n22161);
  and g36374 (n22162, n_14305, n_14308);
  not g36375 (n_14309, n21521);
  and g36376 (n22163, n_14309, n21532);
  not g36377 (n_14310, n21533);
  not g36378 (n_14311, n22163);
  and g36379 (n22164, n_14310, n_14311);
  not g36380 (n_14312, n22162);
  and g36381 (n22165, n_14312, n22164);
  not g36382 (n_14313, n22165);
  and g36383 (n22166, n_14310, n_14313);
  not g36384 (n_14314, n22166);
  and g36385 (n22167, n21519, n_14314);
  not g36386 (n_14315, n22167);
  and g36387 (n22168, n_13763, n_14315);
  not g36388 (n_14316, n22168);
  and g36389 (n22169, n20835, n_14316);
  not g36390 (n_14317, n22169);
  and g36391 (n22170, n_13164, n_14317);
  not g36392 (n_14318, n22170);
  and g36393 (n22171, n20800, n_14318);
  not g36394 (n_14319, n22171);
  and g36395 (n22172, n_13131, n_14319);
  not g36396 (n_14320, n22172);
  and g36397 (n22173, n20145, n_14320);
  not g36398 (n_14321, n22173);
  and g36399 (n22174, n_12566, n_14321);
  not g36400 (n_14322, n19518);
  and g36401 (n22175, n19516, n_14322);
  not g36402 (n_14323, n19519);
  not g36403 (n_14324, n22175);
  and g36404 (n22176, n_14323, n_14324);
  not g36405 (n_14325, n22174);
  and g36406 (n22177, n_14325, n22176);
  not g36407 (n_14326, n22177);
  and g36408 (n22178, n_14323, n_14326);
  not g36409 (n_14327, n18946);
  not g36410 (n_14328, n22178);
  and g36411 (n22179, n_14327, n_14328);
  not g36412 (n_14329, n22179);
  and g36413 (n22180, n_11524, n_14329);
  not g36414 (n_14330, n22180);
  and g36415 (n22181, n18396, n_14330);
  not g36416 (n_14331, n22181);
  and g36417 (n22182, n_11044, n_14331);
  not g36418 (n_14332, n17894);
  and g36419 (n22183, n17892, n_14332);
  not g36420 (n_14333, n17895);
  not g36421 (n_14334, n22183);
  and g36422 (n22184, n_14333, n_14334);
  not g36423 (n_14335, n22182);
  and g36424 (n22185, n_14335, n22184);
  not g36425 (n_14336, n22185);
  and g36426 (n22186, n_14333, n_14336);
  not g36427 (n_14337, n17428);
  not g36428 (n_14338, n22186);
  and g36429 (n22187, n_14337, n_14338);
  not g36430 (n_14339, n22187);
  and g36431 (n22188, n_10206, n_14339);
  not g36432 (n_14340, n22188);
  and g36433 (n22189, n17001, n_14340);
  not g36434 (n_14341, n22189);
  and g36435 (n22190, n_9838, n_14341);
  not g36436 (n_14342, n16606);
  and g36437 (n22191, n16604, n_14342);
  not g36438 (n_14343, n16607);
  not g36439 (n_14344, n22191);
  and g36440 (n22192, n_14343, n_14344);
  not g36441 (n_14345, n22190);
  and g36442 (n22193, n_14345, n22192);
  not g36443 (n_14346, n22193);
  and g36444 (n22194, n_14343, n_14346);
  not g36445 (n_14347, n16443);
  not g36446 (n_14348, n22194);
  and g36447 (n22195, n_14347, n_14348);
  not g36448 (n_14349, n22195);
  and g36449 (n22196, n_9358, n_14349);
  not g36450 (n_14350, n22196);
  and g36451 (n22197, n16272, n_14350);
  not g36452 (n_14351, n22197);
  and g36453 (n22198, n_9214, n_14351);
  not g36454 (n_14352, n15652);
  and g36455 (n22199, n15650, n_14352);
  not g36456 (n_14353, n15653);
  not g36457 (n_14354, n22199);
  and g36458 (n22200, n_14353, n_14354);
  not g36459 (n_14355, n22198);
  and g36460 (n22201, n_14355, n22200);
  not g36461 (n_14356, n22201);
  and g36462 (n22202, n_14353, n_14356);
  not g36463 (n_14357, n15508);
  not g36464 (n_14358, n22202);
  and g36465 (n22203, n_14357, n_14358);
  not g36466 (n_14359, n22203);
  and g36467 (n22204, n_8770, n_14359);
  not g36468 (n_14360, n22204);
  and g36469 (n22205, n15203, n_14360);
  not g36470 (n_14361, n22205);
  and g36471 (n22206, n_8578, n_14361);
  not g36472 (n_14362, n14952);
  and g36473 (n22207, n14950, n_14362);
  not g36474 (n_14363, n14953);
  not g36475 (n_14364, n22207);
  and g36476 (n22208, n_14363, n_14364);
  not g36477 (n_14365, n22206);
  and g36478 (n22209, n_14365, n22208);
  not g36479 (n_14366, n22209);
  and g36480 (n22210, n_14363, n_14366);
  not g36481 (n_14367, n14809);
  not g36482 (n_14368, n22210);
  and g36483 (n22211, n_14367, n_14368);
  not g36484 (n_14369, n22211);
  and g36485 (n22212, n_8282, n_14369);
  not g36486 (n_14370, n22212);
  and g36487 (n22213, n14696, n_14370);
  not g36488 (n_14371, n22213);
  and g36489 (n22214, n_8187, n_14371);
  not g36490 (n_14372, n14323);
  and g36491 (n22215, n14321, n_14372);
  not g36492 (n_14373, n14324);
  not g36493 (n_14374, n22215);
  and g36494 (n22216, n_14373, n_14374);
  not g36495 (n_14375, n22214);
  and g36496 (n22217, n_14375, n22216);
  not g36497 (n_14376, n22217);
  and g36498 (n22218, n_14373, n_14376);
  not g36499 (n_14377, n14154);
  not g36500 (n_14378, n22218);
  and g36501 (n22219, n_14377, n_14378);
  not g36502 (n_14379, n22219);
  and g36503 (n22220, n_7894, n_14379);
  not g36504 (n_14380, n22220);
  and g36505 (n22221, n14039, n_14380);
  not g36506 (n_14381, n22221);
  and g36507 (n22222, n_7794, n_14381);
  and g36508 (n22223, n_7723, n_7726);
  and g36509 (n22224, n_7535, n_7570);
  and g36510 (n22225, n3884, n13941);
  and g36511 (n22226, n3967, n13633);
  and g36512 (n22227, n4046, n_7540);
  and g36518 (n22230, n4050, n14136);
  not g36521 (n_14386, n22231);
  and g36522 (n22232, \a[26] , n_14386);
  not g36523 (n_14387, n22232);
  and g36524 (n22233, \a[26] , n_14387);
  and g36525 (n22234, n_14386, n_14387);
  not g36526 (n_14388, n22233);
  not g36527 (n_14389, n22234);
  and g36528 (n22235, n_14388, n_14389);
  not g36529 (n_14390, n22224);
  not g36530 (n_14391, n22235);
  and g36531 (n22236, n_14390, n_14391);
  not g36532 (n_14392, n22236);
  and g36533 (n22237, n_14390, n_14392);
  and g36534 (n22238, n_14391, n_14392);
  not g36535 (n_14393, n22237);
  not g36536 (n_14394, n22238);
  and g36537 (n22239, n_14393, n_14394);
  and g36538 (n22240, n75, n_7677);
  and g36539 (n22241, n3020, n13521);
  and g36540 (n22242, n3023, n13491);
  and g36541 (n22243, n3028, n13518);
  not g36549 (n_14399, n4533);
  and g36550 (n22247, n_14399, n13938);
  and g36551 (n22248, n_732, n22247);
  not g36552 (n_14400, n22248);
  and g36553 (n22249, n_7417, n_14400);
  not g36554 (n_14401, n22249);
  and g36555 (n22250, \a[23] , n_14401);
  and g36556 (n22251, n_27, n22249);
  not g36557 (n_14402, n22250);
  not g36558 (n_14403, n22251);
  and g36559 (n22252, n_14402, n_14403);
  and g36576 (n22269, n13574, n22268);
  not g36577 (n_14404, n22268);
  and g36578 (n22270, n_7494, n_14404);
  not g36579 (n_14405, n22269);
  not g36580 (n_14406, n22270);
  and g36581 (n22271, n_14405, n_14406);
  and g36582 (n22272, n22252, n22271);
  not g36583 (n_14407, n22252);
  not g36584 (n_14408, n22271);
  and g36585 (n22273, n_14407, n_14408);
  not g36586 (n_14409, n22272);
  not g36587 (n_14410, n22273);
  and g36588 (n22274, n_14409, n_14410);
  not g36589 (n_14411, n13580);
  and g36590 (n22275, n_14411, n22274);
  not g36591 (n_14412, n22274);
  and g36592 (n22276, n13580, n_14412);
  not g36593 (n_14413, n22275);
  not g36594 (n_14414, n22276);
  and g36595 (n22277, n_14413, n_14414);
  not g36596 (n_14415, n22246);
  and g36597 (n22278, n_14415, n22277);
  not g36598 (n_14416, n22278);
  and g36599 (n22279, n22277, n_14416);
  and g36600 (n22280, n_14415, n_14416);
  not g36601 (n_14417, n22279);
  not g36602 (n_14418, n22280);
  and g36603 (n22281, n_14417, n_14418);
  and g36604 (n22282, n_7509, n_7531);
  and g36605 (n22283, n22281, n22282);
  not g36606 (n_14419, n22281);
  not g36607 (n_14420, n22282);
  and g36608 (n22284, n_14419, n_14420);
  not g36609 (n_14421, n22283);
  not g36610 (n_14422, n22284);
  and g36611 (n22285, n_14421, n_14422);
  and g36612 (n22286, n3457, n13630);
  and g36613 (n22287, n3542, n13515);
  and g36614 (n22288, n3606, n13597);
  and g36620 (n22291, n3368, n13976);
  not g36623 (n_14427, n22292);
  and g36624 (n22293, \a[29] , n_14427);
  not g36625 (n_14428, n22293);
  and g36626 (n22294, \a[29] , n_14428);
  and g36627 (n22295, n_14427, n_14428);
  not g36628 (n_14429, n22294);
  not g36629 (n_14430, n22295);
  and g36630 (n22296, n_14429, n_14430);
  not g36631 (n_14431, n22296);
  and g36632 (n22297, n22285, n_14431);
  not g36633 (n_14432, n22297);
  and g36634 (n22298, n22285, n_14432);
  and g36635 (n22299, n_14431, n_14432);
  not g36636 (n_14433, n22298);
  not g36637 (n_14434, n22299);
  and g36638 (n22300, n_14433, n_14434);
  not g36639 (n_14435, n22239);
  and g36640 (n22301, n_14435, n22300);
  not g36641 (n_14436, n22300);
  and g36642 (n22302, n22239, n_14436);
  not g36643 (n_14437, n22301);
  not g36644 (n_14438, n22302);
  and g36645 (n22303, n_14437, n_14438);
  not g36646 (n_14439, n22223);
  not g36647 (n_14440, n22303);
  and g36648 (n22304, n_14439, n_14440);
  and g36649 (n22305, n22223, n22303);
  not g36650 (n_14441, n22304);
  not g36651 (n_14442, n22305);
  and g36652 (n22306, n_14441, n_14442);
  not g36653 (n_14443, n22222);
  and g36654 (n22307, n_14443, n22306);
  not g36655 (n_14444, n22306);
  and g36656 (n22308, n22222, n_14444);
  not g36657 (n_14445, n22307);
  not g36658 (n_14446, n22308);
  and g36659 (n22309, n_14445, n_14446);
  and g36660 (n22310, n71, n22309);
  and g36661 (n22311, n14154, n22218);
  not g36662 (n_14447, n22311);
  and g36663 (n22312, n_14379, n_14447);
  and g36664 (n22313, n9867, n22312);
  not g36665 (n_14448, n14039);
  and g36666 (n22314, n_14448, n22220);
  not g36667 (n_14449, n22314);
  and g36668 (n22315, n_14381, n_14449);
  and g36669 (n22316, n10434, n22315);
  not g36675 (n_14453, n22216);
  and g36676 (n22319, n22214, n_14453);
  not g36677 (n_14454, n22319);
  and g36678 (n22320, n_14376, n_14454);
  and g36679 (n22321, n22312, n22320);
  not g36680 (n_14455, n14696);
  and g36681 (n22322, n_14455, n22212);
  not g36682 (n_14456, n22322);
  and g36683 (n22323, n_14371, n_14456);
  and g36684 (n22324, n22320, n22323);
  and g36685 (n22325, n14809, n22210);
  not g36686 (n_14457, n22325);
  and g36687 (n22326, n_14369, n_14457);
  and g36688 (n22327, n22323, n22326);
  not g36689 (n_14458, n22208);
  and g36690 (n22328, n22206, n_14458);
  not g36691 (n_14459, n22328);
  and g36692 (n22329, n_14366, n_14459);
  and g36693 (n22330, n22326, n22329);
  not g36694 (n_14460, n15203);
  and g36695 (n22331, n_14460, n22204);
  not g36696 (n_14461, n22331);
  and g36697 (n22332, n_14361, n_14461);
  and g36698 (n22333, n22329, n22332);
  and g36699 (n22334, n15508, n22202);
  not g36700 (n_14462, n22334);
  and g36701 (n22335, n_14359, n_14462);
  and g36702 (n22336, n22332, n22335);
  not g36703 (n_14463, n22200);
  and g36704 (n22337, n22198, n_14463);
  not g36705 (n_14464, n22337);
  and g36706 (n22338, n_14356, n_14464);
  and g36707 (n22339, n22335, n22338);
  not g36708 (n_14465, n16272);
  and g36709 (n22340, n_14465, n22196);
  not g36710 (n_14466, n22340);
  and g36711 (n22341, n_14351, n_14466);
  and g36712 (n22342, n22338, n22341);
  and g36713 (n22343, n16443, n22194);
  not g36714 (n_14467, n22343);
  and g36715 (n22344, n_14349, n_14467);
  and g36716 (n22345, n22341, n22344);
  not g36717 (n_14468, n22192);
  and g36718 (n22346, n22190, n_14468);
  not g36719 (n_14469, n22346);
  and g36720 (n22347, n_14346, n_14469);
  and g36721 (n22348, n22344, n22347);
  not g36722 (n_14470, n17001);
  and g36723 (n22349, n_14470, n22188);
  not g36724 (n_14471, n22349);
  and g36725 (n22350, n_14341, n_14471);
  and g36726 (n22351, n22347, n22350);
  and g36727 (n22352, n17428, n22186);
  not g36728 (n_14472, n22352);
  and g36729 (n22353, n_14339, n_14472);
  and g36730 (n22354, n22350, n22353);
  not g36731 (n_14473, n22184);
  and g36732 (n22355, n22182, n_14473);
  not g36733 (n_14474, n22355);
  and g36734 (n22356, n_14336, n_14474);
  and g36735 (n22357, n22353, n22356);
  not g36736 (n_14475, n18396);
  and g36737 (n22358, n_14475, n22180);
  not g36738 (n_14476, n22358);
  and g36739 (n22359, n_14331, n_14476);
  and g36740 (n22360, n22356, n22359);
  and g36741 (n22361, n18946, n22178);
  not g36742 (n_14477, n22361);
  and g36743 (n22362, n_14329, n_14477);
  and g36744 (n22363, n22359, n22362);
  not g36745 (n_14478, n22176);
  and g36746 (n22364, n22174, n_14478);
  not g36747 (n_14479, n22364);
  and g36748 (n22365, n_14326, n_14479);
  and g36749 (n22366, n22362, n22365);
  not g36750 (n_14480, n20145);
  and g36751 (n22367, n_14480, n22172);
  not g36752 (n_14481, n22367);
  and g36753 (n22368, n_14321, n_14481);
  and g36754 (n22369, n22365, n22368);
  not g36755 (n_14482, n20800);
  and g36756 (n22370, n_14482, n22170);
  not g36757 (n_14483, n22370);
  and g36758 (n22371, n_14319, n_14483);
  and g36759 (n22372, n22368, n22371);
  not g36760 (n_14484, n20835);
  and g36761 (n22373, n_14484, n22168);
  not g36762 (n_14485, n22373);
  and g36763 (n22374, n_14317, n_14485);
  and g36764 (n22375, n22371, n22374);
  not g36765 (n_14486, n21519);
  and g36766 (n22376, n_14486, n22166);
  not g36767 (n_14487, n22376);
  and g36768 (n22377, n_14315, n_14487);
  and g36769 (n22378, n22374, n22377);
  not g36770 (n_14488, n22164);
  and g36771 (n22379, n22162, n_14488);
  not g36772 (n_14489, n22379);
  and g36773 (n22380, n_14313, n_14489);
  and g36774 (n22381, n22377, n22380);
  not g36775 (n_14490, n22377);
  not g36776 (n_14491, n22380);
  and g36777 (n22382, n_14490, n_14491);
  not g36778 (n_14492, n22160);
  and g36779 (n22383, n22158, n_14492);
  not g36780 (n_14493, n22383);
  and g36781 (n22384, n_14308, n_14493);
  and g36782 (n22385, n22380, n22384);
  not g36783 (n_14494, n22156);
  and g36784 (n22386, n22154, n_14494);
  not g36785 (n_14495, n22386);
  and g36786 (n22387, n_14303, n_14495);
  and g36787 (n22388, n22384, n22387);
  not g36788 (n_14496, n22152);
  and g36789 (n22389, n22150, n_14496);
  not g36790 (n_14497, n22389);
  and g36791 (n22390, n_14298, n_14497);
  and g36792 (n22391, n22387, n22390);
  not g36793 (n_14498, n22148);
  and g36794 (n22392, n22146, n_14498);
  not g36795 (n_14499, n22392);
  and g36796 (n22393, n_14293, n_14499);
  and g36797 (n22394, n22390, n22393);
  not g36798 (n_14500, n22144);
  and g36799 (n22395, n22142, n_14500);
  not g36800 (n_14501, n22395);
  and g36801 (n22396, n_14288, n_14501);
  and g36802 (n22397, n22393, n22396);
  not g36803 (n_14502, n22140);
  and g36804 (n22398, n22138, n_14502);
  not g36805 (n_14503, n22398);
  and g36806 (n22399, n_14283, n_14503);
  and g36807 (n22400, n22396, n22399);
  not g36808 (n_14504, n22136);
  and g36809 (n22401, n22134, n_14504);
  not g36810 (n_14505, n22401);
  and g36811 (n22402, n_14278, n_14505);
  and g36812 (n22403, n22399, n22402);
  and g36813 (n22404, n_14271, n_14273);
  and g36814 (n22405, n_14272, n_14273);
  not g36815 (n_14506, n22404);
  not g36816 (n_14507, n22405);
  and g36817 (n22406, n_14506, n_14507);
  not g36818 (n_14508, n22406);
  and g36819 (n22407, n22402, n_14508);
  not g36820 (n_14509, n22399);
  and g36821 (n22408, n_14509, n22407);
  not g36822 (n_14510, n22403);
  not g36823 (n_14511, n22408);
  and g36824 (n22409, n_14510, n_14511);
  not g36825 (n_14512, n22396);
  and g36826 (n22410, n_14512, n_14509);
  not g36827 (n_14513, n22400);
  not g36828 (n_14514, n22410);
  and g36829 (n22411, n_14513, n_14514);
  not g36830 (n_14515, n22409);
  and g36831 (n22412, n_14515, n22411);
  not g36832 (n_14516, n22412);
  and g36833 (n22413, n_14513, n_14516);
  not g36834 (n_14517, n22393);
  and g36835 (n22414, n_14517, n_14512);
  not g36836 (n_14518, n22397);
  not g36837 (n_14519, n22414);
  and g36838 (n22415, n_14518, n_14519);
  not g36839 (n_14520, n22413);
  and g36840 (n22416, n_14520, n22415);
  not g36841 (n_14521, n22416);
  and g36842 (n22417, n_14518, n_14521);
  not g36843 (n_14522, n22390);
  and g36844 (n22418, n_14522, n_14517);
  not g36845 (n_14523, n22394);
  not g36846 (n_14524, n22418);
  and g36847 (n22419, n_14523, n_14524);
  not g36848 (n_14525, n22417);
  and g36849 (n22420, n_14525, n22419);
  not g36850 (n_14526, n22420);
  and g36851 (n22421, n_14523, n_14526);
  not g36852 (n_14527, n22387);
  and g36853 (n22422, n_14527, n_14522);
  not g36854 (n_14528, n22391);
  not g36855 (n_14529, n22422);
  and g36856 (n22423, n_14528, n_14529);
  not g36857 (n_14530, n22421);
  and g36858 (n22424, n_14530, n22423);
  not g36859 (n_14531, n22424);
  and g36860 (n22425, n_14528, n_14531);
  not g36861 (n_14532, n22384);
  and g36862 (n22426, n_14532, n_14527);
  not g36863 (n_14533, n22388);
  not g36864 (n_14534, n22426);
  and g36865 (n22427, n_14533, n_14534);
  not g36866 (n_14535, n22425);
  and g36867 (n22428, n_14535, n22427);
  not g36868 (n_14536, n22428);
  and g36869 (n22429, n_14533, n_14536);
  and g36870 (n22430, n_14491, n_14532);
  not g36871 (n_14537, n22385);
  not g36872 (n_14538, n22430);
  and g36873 (n22431, n_14537, n_14538);
  not g36874 (n_14539, n22429);
  and g36875 (n22432, n_14539, n22431);
  not g36876 (n_14540, n22432);
  and g36877 (n22433, n_14537, n_14540);
  not g36878 (n_14541, n22381);
  not g36879 (n_14542, n22433);
  and g36880 (n22434, n_14541, n_14542);
  not g36881 (n_14543, n22382);
  and g36882 (n22435, n_14543, n22434);
  not g36883 (n_14544, n22435);
  and g36884 (n22436, n_14541, n_14544);
  not g36885 (n_14545, n22374);
  and g36886 (n22437, n_14545, n_14490);
  not g36887 (n_14546, n22378);
  not g36888 (n_14547, n22437);
  and g36889 (n22438, n_14546, n_14547);
  not g36890 (n_14548, n22436);
  and g36891 (n22439, n_14548, n22438);
  not g36892 (n_14549, n22439);
  and g36893 (n22440, n_14546, n_14549);
  not g36894 (n_14550, n22371);
  and g36895 (n22441, n_14550, n_14545);
  not g36896 (n_14551, n22375);
  not g36897 (n_14552, n22441);
  and g36898 (n22442, n_14551, n_14552);
  not g36899 (n_14553, n22440);
  and g36900 (n22443, n_14553, n22442);
  not g36901 (n_14554, n22443);
  and g36902 (n22444, n_14551, n_14554);
  not g36903 (n_14555, n22368);
  and g36904 (n22445, n_14555, n_14550);
  not g36905 (n_14556, n22372);
  not g36906 (n_14557, n22445);
  and g36907 (n22446, n_14556, n_14557);
  not g36908 (n_14558, n22444);
  and g36909 (n22447, n_14558, n22446);
  not g36910 (n_14559, n22447);
  and g36911 (n22448, n_14556, n_14559);
  not g36912 (n_14560, n22365);
  and g36913 (n22449, n_14560, n_14555);
  not g36914 (n_14561, n22448);
  not g36915 (n_14562, n22449);
  and g36916 (n22450, n_14561, n_14562);
  not g36917 (n_14563, n22369);
  and g36918 (n22451, n_14563, n22450);
  not g36919 (n_14564, n22451);
  and g36920 (n22452, n_14563, n_14564);
  not g36921 (n_14565, n22362);
  and g36922 (n22453, n_14565, n_14560);
  not g36923 (n_14566, n22452);
  not g36924 (n_14567, n22453);
  and g36925 (n22454, n_14566, n_14567);
  not g36926 (n_14568, n22366);
  and g36927 (n22455, n_14568, n22454);
  not g36928 (n_14569, n22455);
  and g36929 (n22456, n_14568, n_14569);
  not g36930 (n_14570, n22359);
  and g36931 (n22457, n_14570, n_14565);
  not g36932 (n_14571, n22363);
  not g36933 (n_14572, n22457);
  and g36934 (n22458, n_14571, n_14572);
  not g36935 (n_14573, n22456);
  and g36936 (n22459, n_14573, n22458);
  not g36937 (n_14574, n22459);
  and g36938 (n22460, n_14571, n_14574);
  not g36939 (n_14575, n22356);
  and g36940 (n22461, n_14575, n_14570);
  not g36941 (n_14576, n22460);
  not g36942 (n_14577, n22461);
  and g36943 (n22462, n_14576, n_14577);
  not g36944 (n_14578, n22360);
  and g36945 (n22463, n_14578, n22462);
  not g36946 (n_14579, n22463);
  and g36947 (n22464, n_14578, n_14579);
  not g36948 (n_14580, n22353);
  and g36949 (n22465, n_14580, n_14575);
  not g36950 (n_14581, n22464);
  not g36951 (n_14582, n22465);
  and g36952 (n22466, n_14581, n_14582);
  not g36953 (n_14583, n22357);
  and g36954 (n22467, n_14583, n22466);
  not g36955 (n_14584, n22467);
  and g36956 (n22468, n_14583, n_14584);
  not g36957 (n_14585, n22350);
  and g36958 (n22469, n_14585, n_14580);
  not g36959 (n_14586, n22354);
  not g36960 (n_14587, n22469);
  and g36961 (n22470, n_14586, n_14587);
  not g36962 (n_14588, n22468);
  and g36963 (n22471, n_14588, n22470);
  not g36964 (n_14589, n22471);
  and g36965 (n22472, n_14586, n_14589);
  not g36966 (n_14590, n22347);
  and g36967 (n22473, n_14590, n_14585);
  not g36968 (n_14591, n22472);
  not g36969 (n_14592, n22473);
  and g36970 (n22474, n_14591, n_14592);
  not g36971 (n_14593, n22351);
  and g36972 (n22475, n_14593, n22474);
  not g36973 (n_14594, n22475);
  and g36974 (n22476, n_14593, n_14594);
  not g36975 (n_14595, n22344);
  and g36976 (n22477, n_14595, n_14590);
  not g36977 (n_14596, n22476);
  not g36978 (n_14597, n22477);
  and g36979 (n22478, n_14596, n_14597);
  not g36980 (n_14598, n22348);
  and g36981 (n22479, n_14598, n22478);
  not g36982 (n_14599, n22479);
  and g36983 (n22480, n_14598, n_14599);
  not g36984 (n_14600, n22341);
  and g36985 (n22481, n_14600, n_14595);
  not g36986 (n_14601, n22345);
  not g36987 (n_14602, n22481);
  and g36988 (n22482, n_14601, n_14602);
  not g36989 (n_14603, n22480);
  and g36990 (n22483, n_14603, n22482);
  not g36991 (n_14604, n22483);
  and g36992 (n22484, n_14601, n_14604);
  not g36993 (n_14605, n22338);
  and g36994 (n22485, n_14605, n_14600);
  not g36995 (n_14606, n22484);
  not g36996 (n_14607, n22485);
  and g36997 (n22486, n_14606, n_14607);
  not g36998 (n_14608, n22342);
  and g36999 (n22487, n_14608, n22486);
  not g37000 (n_14609, n22487);
  and g37001 (n22488, n_14608, n_14609);
  not g37002 (n_14610, n22335);
  and g37003 (n22489, n_14610, n_14605);
  not g37004 (n_14611, n22488);
  not g37005 (n_14612, n22489);
  and g37006 (n22490, n_14611, n_14612);
  not g37007 (n_14613, n22339);
  and g37008 (n22491, n_14613, n22490);
  not g37009 (n_14614, n22491);
  and g37010 (n22492, n_14613, n_14614);
  not g37011 (n_14615, n22332);
  and g37012 (n22493, n_14615, n_14610);
  not g37013 (n_14616, n22336);
  not g37014 (n_14617, n22493);
  and g37015 (n22494, n_14616, n_14617);
  not g37016 (n_14618, n22492);
  and g37017 (n22495, n_14618, n22494);
  not g37018 (n_14619, n22495);
  and g37019 (n22496, n_14616, n_14619);
  not g37020 (n_14620, n22329);
  and g37021 (n22497, n_14620, n_14615);
  not g37022 (n_14621, n22496);
  not g37023 (n_14622, n22497);
  and g37024 (n22498, n_14621, n_14622);
  not g37025 (n_14623, n22333);
  and g37026 (n22499, n_14623, n22498);
  not g37027 (n_14624, n22499);
  and g37028 (n22500, n_14623, n_14624);
  not g37029 (n_14625, n22326);
  and g37030 (n22501, n_14625, n_14620);
  not g37031 (n_14626, n22500);
  not g37032 (n_14627, n22501);
  and g37033 (n22502, n_14626, n_14627);
  not g37034 (n_14628, n22330);
  and g37035 (n22503, n_14628, n22502);
  not g37036 (n_14629, n22503);
  and g37037 (n22504, n_14628, n_14629);
  not g37038 (n_14630, n22323);
  and g37039 (n22505, n_14630, n_14625);
  not g37040 (n_14631, n22327);
  not g37041 (n_14632, n22505);
  and g37042 (n22506, n_14631, n_14632);
  not g37043 (n_14633, n22504);
  and g37044 (n22507, n_14633, n22506);
  not g37045 (n_14634, n22507);
  and g37046 (n22508, n_14631, n_14634);
  not g37047 (n_14635, n22320);
  and g37048 (n22509, n_14635, n_14630);
  not g37049 (n_14636, n22508);
  not g37050 (n_14637, n22509);
  and g37051 (n22510, n_14636, n_14637);
  not g37052 (n_14638, n22324);
  and g37053 (n22511, n_14638, n22510);
  not g37054 (n_14639, n22511);
  and g37055 (n22512, n_14638, n_14639);
  not g37056 (n_14640, n22312);
  and g37057 (n22513, n_14640, n_14635);
  not g37058 (n_14641, n22512);
  not g37059 (n_14642, n22513);
  and g37060 (n22514, n_14641, n_14642);
  not g37061 (n_14643, n22321);
  and g37062 (n22515, n_14643, n22514);
  not g37063 (n_14644, n22515);
  and g37064 (n22516, n_14643, n_14644);
  not g37065 (n_14645, n22315);
  and g37066 (n22517, n_14640, n_14645);
  and g37067 (n22518, n22312, n22315);
  not g37068 (n_14646, n22517);
  not g37069 (n_14647, n22518);
  and g37070 (n22519, n_14646, n_14647);
  not g37071 (n_14648, n22516);
  and g37072 (n22520, n_14648, n22519);
  not g37073 (n_14649, n22520);
  and g37074 (n22521, n_14647, n_14649);
  and g37075 (n22522, n22309, n22315);
  not g37076 (n_14650, n22309);
  and g37077 (n22523, n_14650, n_14645);
  not g37078 (n_14651, n22521);
  not g37079 (n_14652, n22523);
  and g37080 (n22524, n_14651, n_14652);
  not g37081 (n_14653, n22522);
  and g37082 (n22525, n_14653, n22524);
  not g37083 (n_14654, n22525);
  and g37084 (n22526, n_14651, n_14654);
  and g37085 (n22527, n_14653, n_14654);
  and g37086 (n22528, n_14652, n22527);
  not g37087 (n_14655, n22526);
  not g37088 (n_14656, n22528);
  and g37089 (n22529, n_14655, n_14656);
  not g37090 (n_14657, n22529);
  and g37091 (n22530, n9870, n_14657);
  not g37094 (n_14659, n22531);
  and g37095 (n22532, \a[5] , n_14659);
  not g37096 (n_14660, n22532);
  and g37097 (n22533, n_14659, n_14660);
  and g37098 (n22534, \a[5] , n_14660);
  not g37099 (n_14661, n22533);
  not g37100 (n_14662, n22534);
  and g37101 (n22535, n_14661, n_14662);
  and g37102 (n22536, n7983, n22332);
  and g37103 (n22537, n7291, n22338);
  and g37104 (n22538, n7632, n22335);
  not g37110 (n_14666, n22494);
  and g37111 (n22541, n22492, n_14666);
  not g37112 (n_14667, n22541);
  and g37113 (n22542, n_14619, n_14667);
  and g37114 (n22543, n7294, n22542);
  not g37117 (n_14669, n22544);
  and g37118 (n22545, \a[11] , n_14669);
  not g37119 (n_14670, n22545);
  and g37120 (n22546, n_14669, n_14670);
  and g37121 (n22547, \a[11] , n_14670);
  not g37122 (n_14671, n22546);
  not g37123 (n_14672, n22547);
  and g37124 (n22548, n_14671, n_14672);
  and g37125 (n22549, n6233, n22353);
  and g37126 (n22550, n5663, n22359);
  and g37127 (n22551, n5939, n22356);
  and g37133 (n22554, n_14581, n_14584);
  and g37134 (n22555, n_14582, n22468);
  not g37135 (n_14676, n22554);
  not g37136 (n_14677, n22555);
  and g37137 (n22556, n_14676, n_14677);
  not g37138 (n_14678, n22556);
  and g37139 (n22557, n5666, n_14678);
  not g37142 (n_14680, n22558);
  and g37143 (n22559, \a[17] , n_14680);
  not g37144 (n_14681, n22559);
  and g37145 (n22560, n_14680, n_14681);
  and g37146 (n22561, \a[17] , n_14681);
  not g37147 (n_14682, n22560);
  not g37148 (n_14683, n22561);
  and g37149 (n22562, n_14682, n_14683);
  and g37150 (n22563, n4694, n22374);
  and g37151 (n22564, n4533, n22380);
  and g37152 (n22565, n4604, n22377);
  not g37158 (n_14687, n22438);
  and g37159 (n22568, n22436, n_14687);
  not g37160 (n_14688, n22568);
  and g37161 (n22569, n_14549, n_14688);
  and g37162 (n22570, n4536, n22569);
  not g37165 (n_14690, n22571);
  and g37166 (n22572, \a[23] , n_14690);
  not g37167 (n_14691, n22572);
  and g37168 (n22573, n_14690, n_14691);
  and g37169 (n22574, \a[23] , n_14691);
  not g37170 (n_14692, n22573);
  not g37171 (n_14693, n22574);
  and g37172 (n22575, n_14692, n_14693);
  and g37173 (n22576, n3884, n22387);
  and g37174 (n22577, n3967, n22393);
  and g37175 (n22578, n4046, n22390);
  not g37181 (n_14697, n22423);
  and g37182 (n22581, n22421, n_14697);
  not g37183 (n_14698, n22581);
  and g37184 (n22582, n_14531, n_14698);
  and g37185 (n22583, n4050, n22582);
  not g37188 (n_14700, n22584);
  and g37189 (n22585, \a[26] , n_14700);
  not g37190 (n_14701, n22585);
  and g37191 (n22586, n_14700, n_14701);
  and g37192 (n22587, \a[26] , n_14701);
  not g37193 (n_14702, n22586);
  not g37194 (n_14703, n22587);
  and g37195 (n22588, n_14702, n_14703);
  and g37196 (n22589, n3457, n22396);
  and g37197 (n22590, n3542, n22402);
  and g37198 (n22591, n3606, n22399);
  not g37204 (n_14707, n22411);
  and g37205 (n22594, n22409, n_14707);
  not g37206 (n_14708, n22594);
  and g37207 (n22595, n_14516, n_14708);
  and g37208 (n22596, n3368, n22595);
  not g37211 (n_14710, n22597);
  and g37212 (n22598, \a[29] , n_14710);
  not g37213 (n_14711, n22598);
  and g37214 (n22599, n_14710, n_14711);
  and g37215 (n22600, \a[29] , n_14711);
  not g37216 (n_14712, n22599);
  not g37217 (n_14713, n22600);
  and g37218 (n22601, n_14712, n_14713);
  and g37219 (n22602, n_479, n_14508);
  not g37220 (n_14714, n22602);
  and g37221 (n22603, \a[29] , n_14714);
  and g37222 (n22604, n3606, n_14508);
  and g37223 (n22605, n3457, n22402);
  not g37224 (n_14715, n22604);
  not g37225 (n_14716, n22605);
  and g37226 (n22606, n_14715, n_14716);
  and g37227 (n22607, n22402, n22406);
  not g37228 (n_14717, n22402);
  and g37229 (n22608, n_14717, n_14508);
  not g37230 (n_14718, n22607);
  not g37231 (n_14719, n22608);
  and g37232 (n22609, n_14718, n_14719);
  not g37233 (n_14720, n22609);
  and g37234 (n22610, n3368, n_14720);
  not g37235 (n_14721, n22610);
  and g37236 (n22611, n22606, n_14721);
  not g37237 (n_14722, n22611);
  and g37238 (n22612, \a[29] , n_14722);
  not g37239 (n_14723, n22612);
  and g37240 (n22613, \a[29] , n_14723);
  and g37241 (n22614, n_14722, n_14723);
  not g37242 (n_14724, n22613);
  not g37243 (n_14725, n22614);
  and g37244 (n22615, n_14724, n_14725);
  not g37245 (n_14726, n22615);
  and g37246 (n22616, n22603, n_14726);
  and g37247 (n22617, n3457, n22399);
  and g37248 (n22618, n3542, n_14508);
  and g37249 (n22619, n3606, n22402);
  not g37250 (n_14727, n22618);
  not g37251 (n_14728, n22619);
  and g37252 (n22620, n_14727, n_14728);
  not g37253 (n_14729, n22617);
  and g37254 (n22621, n_14729, n22620);
  and g37255 (n22622, n_489, n22621);
  and g37256 (n22623, n_14509, n22607);
  and g37257 (n22624, n22399, n_14718);
  not g37258 (n_14730, n22623);
  not g37259 (n_14731, n22624);
  and g37260 (n22625, n_14730, n_14731);
  and g37261 (n22626, n22621, n22625);
  not g37262 (n_14732, n22622);
  not g37263 (n_14733, n22626);
  and g37264 (n22627, n_14732, n_14733);
  not g37265 (n_14734, n22627);
  and g37266 (n22628, \a[29] , n_14734);
  and g37267 (n22629, n_15, n22627);
  not g37268 (n_14735, n22628);
  not g37269 (n_14736, n22629);
  and g37270 (n22630, n_14735, n_14736);
  not g37271 (n_14737, n22630);
  and g37272 (n22631, n22616, n_14737);
  and g37273 (n22632, n_2599, n_14508);
  not g37274 (n_14738, n22632);
  and g37275 (n22633, n22631, n_14738);
  not g37276 (n_14739, n22631);
  and g37277 (n22634, n_14739, n22632);
  not g37278 (n_14740, n22633);
  not g37279 (n_14741, n22634);
  and g37280 (n22635, n_14740, n_14741);
  not g37281 (n_14742, n22601);
  not g37282 (n_14743, n22635);
  and g37283 (n22636, n_14742, n_14743);
  and g37284 (n22637, n22601, n22635);
  not g37285 (n_14744, n22636);
  not g37286 (n_14745, n22637);
  and g37287 (n22638, n_14744, n_14745);
  not g37288 (n_14746, n22588);
  and g37289 (n22639, n_14746, n22638);
  not g37290 (n_14747, n22639);
  and g37291 (n22640, n_14746, n_14747);
  and g37292 (n22641, n22638, n_14747);
  not g37293 (n_14748, n22640);
  not g37294 (n_14749, n22641);
  and g37295 (n22642, n_14748, n_14749);
  and g37296 (n22643, n3884, n22390);
  and g37297 (n22644, n3967, n22396);
  and g37298 (n22645, n4046, n22393);
  not g37304 (n_14753, n22419);
  and g37305 (n22648, n22417, n_14753);
  not g37306 (n_14754, n22648);
  and g37307 (n22649, n_14526, n_14754);
  and g37308 (n22650, n4050, n22649);
  not g37311 (n_14756, n22651);
  and g37312 (n22652, \a[26] , n_14756);
  not g37313 (n_14757, n22652);
  and g37314 (n22653, n_14756, n_14757);
  and g37315 (n22654, \a[26] , n_14757);
  not g37316 (n_14758, n22653);
  not g37317 (n_14759, n22654);
  and g37318 (n22655, n_14758, n_14759);
  not g37319 (n_14760, n22616);
  and g37320 (n22656, n_14760, n22630);
  not g37321 (n_14761, n22656);
  and g37322 (n22657, n_14739, n_14761);
  not g37323 (n_14762, n22655);
  and g37324 (n22658, n_14762, n22657);
  not g37325 (n_14763, n22658);
  and g37326 (n22659, n_14762, n_14763);
  and g37327 (n22660, n22657, n_14763);
  not g37328 (n_14764, n22659);
  not g37329 (n_14765, n22660);
  and g37330 (n22661, n_14764, n_14765);
  not g37331 (n_14766, n22603);
  and g37332 (n22662, n_14766, n22615);
  not g37333 (n_14767, n22662);
  and g37334 (n22663, n_14760, n_14767);
  and g37335 (n22664, n3884, n22393);
  and g37336 (n22665, n3967, n22399);
  and g37337 (n22666, n4046, n22396);
  not g37338 (n_14768, n22665);
  not g37339 (n_14769, n22666);
  and g37340 (n22667, n_14768, n_14769);
  not g37341 (n_14770, n22664);
  and g37342 (n22668, n_14770, n22667);
  and g37343 (n22669, n_750, n22668);
  not g37344 (n_14771, n22415);
  and g37345 (n22670, n22413, n_14771);
  not g37346 (n_14772, n22670);
  and g37347 (n22671, n_14521, n_14772);
  not g37348 (n_14773, n22671);
  and g37349 (n22672, n22668, n_14773);
  not g37350 (n_14774, n22669);
  not g37351 (n_14775, n22672);
  and g37352 (n22673, n_14774, n_14775);
  not g37353 (n_14776, n22673);
  and g37354 (n22674, \a[26] , n_14776);
  and g37355 (n22675, n_33, n22673);
  not g37356 (n_14777, n22674);
  not g37357 (n_14778, n22675);
  and g37358 (n22676, n_14777, n_14778);
  not g37359 (n_14779, n22676);
  and g37360 (n22677, n22663, n_14779);
  and g37361 (n22678, n_559, n_14508);
  not g37362 (n_14780, n22678);
  and g37363 (n22679, \a[26] , n_14780);
  and g37364 (n22680, n4046, n_14508);
  and g37365 (n22681, n3884, n22402);
  not g37366 (n_14781, n22680);
  not g37367 (n_14782, n22681);
  and g37368 (n22682, n_14781, n_14782);
  and g37369 (n22683, n4050, n_14720);
  not g37370 (n_14783, n22683);
  and g37371 (n22684, n22682, n_14783);
  not g37372 (n_14784, n22684);
  and g37373 (n22685, \a[26] , n_14784);
  not g37374 (n_14785, n22685);
  and g37375 (n22686, \a[26] , n_14785);
  and g37376 (n22687, n_14784, n_14785);
  not g37377 (n_14786, n22686);
  not g37378 (n_14787, n22687);
  and g37379 (n22688, n_14786, n_14787);
  not g37380 (n_14788, n22688);
  and g37381 (n22689, n22679, n_14788);
  and g37382 (n22690, n3884, n22399);
  and g37383 (n22691, n3967, n_14508);
  and g37384 (n22692, n4046, n22402);
  not g37385 (n_14789, n22691);
  not g37386 (n_14790, n22692);
  and g37387 (n22693, n_14789, n_14790);
  not g37388 (n_14791, n22690);
  and g37389 (n22694, n_14791, n22693);
  and g37390 (n22695, n_750, n22694);
  and g37391 (n22696, n22625, n22694);
  not g37392 (n_14792, n22695);
  not g37393 (n_14793, n22696);
  and g37394 (n22697, n_14792, n_14793);
  not g37395 (n_14794, n22697);
  and g37396 (n22698, \a[26] , n_14794);
  and g37397 (n22699, n_33, n22697);
  not g37398 (n_14795, n22698);
  not g37399 (n_14796, n22699);
  and g37400 (n22700, n_14795, n_14796);
  not g37401 (n_14797, n22700);
  and g37402 (n22701, n22689, n_14797);
  and g37403 (n22702, n22602, n22701);
  not g37404 (n_14798, n22702);
  and g37405 (n22703, n22701, n_14798);
  and g37406 (n22704, n22602, n_14798);
  not g37407 (n_14799, n22703);
  not g37408 (n_14800, n22704);
  and g37409 (n22705, n_14799, n_14800);
  and g37410 (n22706, n3884, n22396);
  and g37411 (n22707, n3967, n22402);
  and g37412 (n22708, n4046, n22399);
  and g37418 (n22711, n4050, n22595);
  not g37421 (n_14805, n22712);
  and g37422 (n22713, \a[26] , n_14805);
  not g37423 (n_14806, n22713);
  and g37424 (n22714, \a[26] , n_14806);
  and g37425 (n22715, n_14805, n_14806);
  not g37426 (n_14807, n22714);
  not g37427 (n_14808, n22715);
  and g37428 (n22716, n_14807, n_14808);
  not g37429 (n_14809, n22705);
  not g37430 (n_14810, n22716);
  and g37431 (n22717, n_14809, n_14810);
  not g37432 (n_14811, n22717);
  and g37433 (n22718, n_14798, n_14811);
  not g37434 (n_14812, n22663);
  and g37435 (n22719, n_14812, n22676);
  not g37436 (n_14813, n22677);
  not g37437 (n_14814, n22719);
  and g37438 (n22720, n_14813, n_14814);
  not g37439 (n_14815, n22718);
  and g37440 (n22721, n_14815, n22720);
  not g37441 (n_14816, n22721);
  and g37442 (n22722, n_14813, n_14816);
  not g37443 (n_14817, n22661);
  not g37444 (n_14818, n22722);
  and g37445 (n22723, n_14817, n_14818);
  not g37446 (n_14819, n22723);
  and g37447 (n22724, n_14763, n_14819);
  not g37448 (n_14820, n22642);
  not g37449 (n_14821, n22724);
  and g37450 (n22725, n_14820, n_14821);
  not g37451 (n_14822, n22725);
  and g37452 (n22726, n_14747, n_14822);
  and g37453 (n22727, n3457, n22393);
  and g37454 (n22728, n3542, n22399);
  and g37455 (n22729, n3606, n22396);
  and g37461 (n22732, n3368, n22671);
  not g37464 (n_14827, n22733);
  and g37465 (n22734, \a[29] , n_14827);
  not g37466 (n_14828, n22734);
  and g37467 (n22735, n_14827, n_14828);
  and g37468 (n22736, \a[29] , n_14828);
  not g37469 (n_14829, n22735);
  not g37470 (n_14830, n22736);
  and g37471 (n22737, n_14829, n_14830);
  and g37514 (n22780, n3020, n22402);
  and g37515 (n22781, n75, n_14720);
  and g37516 (n22782, n3028, n_14508);
  not g37517 (n_14831, n22781);
  not g37518 (n_14832, n22782);
  and g37519 (n22783, n_14831, n_14832);
  not g37520 (n_14833, n22780);
  and g37521 (n22784, n_14833, n22783);
  not g37522 (n_14834, n22779);
  not g37523 (n_14835, n22784);
  and g37524 (n22785, n_14834, n_14835);
  not g37525 (n_14836, n22785);
  and g37526 (n22786, n_14834, n_14836);
  and g37527 (n22787, n_14835, n_14836);
  not g37528 (n_14837, n22786);
  not g37529 (n_14838, n22787);
  and g37530 (n22788, n_14837, n_14838);
  not g37531 (n_14839, n22737);
  not g37532 (n_14840, n22788);
  and g37533 (n22789, n_14839, n_14840);
  not g37534 (n_14841, n22789);
  and g37535 (n22790, n_14839, n_14841);
  and g37536 (n22791, n_14840, n_14841);
  not g37537 (n_14842, n22790);
  not g37538 (n_14843, n22791);
  and g37539 (n22792, n_14842, n_14843);
  and g37540 (n22793, n22631, n22632);
  not g37541 (n_14844, n22793);
  and g37542 (n22794, n_14744, n_14844);
  not g37543 (n_14845, n22792);
  not g37544 (n_14846, n22794);
  and g37545 (n22795, n_14845, n_14846);
  not g37546 (n_14847, n22795);
  and g37547 (n22796, n_14845, n_14847);
  and g37548 (n22797, n_14846, n_14847);
  not g37549 (n_14848, n22796);
  not g37550 (n_14849, n22797);
  and g37551 (n22798, n_14848, n_14849);
  and g37552 (n22799, n3884, n22384);
  and g37553 (n22800, n3967, n22390);
  and g37554 (n22801, n4046, n22387);
  not g37555 (n_14850, n22800);
  not g37556 (n_14851, n22801);
  and g37557 (n22802, n_14850, n_14851);
  not g37558 (n_14852, n22799);
  and g37559 (n22803, n_14852, n22802);
  and g37560 (n22804, n_750, n22803);
  not g37561 (n_14853, n22427);
  and g37562 (n22805, n22425, n_14853);
  not g37563 (n_14854, n22805);
  and g37564 (n22806, n_14536, n_14854);
  not g37565 (n_14855, n22806);
  and g37566 (n22807, n22803, n_14855);
  not g37567 (n_14856, n22804);
  not g37568 (n_14857, n22807);
  and g37569 (n22808, n_14856, n_14857);
  not g37570 (n_14858, n22808);
  and g37571 (n22809, \a[26] , n_14858);
  and g37572 (n22810, n_33, n22808);
  not g37573 (n_14859, n22809);
  not g37574 (n_14860, n22810);
  and g37575 (n22811, n_14859, n_14860);
  not g37576 (n_14861, n22798);
  not g37577 (n_14862, n22811);
  and g37578 (n22812, n_14861, n_14862);
  not g37579 (n_14863, n22812);
  and g37580 (n22813, n_14861, n_14863);
  and g37581 (n22814, n_14862, n_14863);
  not g37582 (n_14864, n22813);
  not g37583 (n_14865, n22814);
  and g37584 (n22815, n_14864, n_14865);
  not g37585 (n_14866, n22726);
  not g37586 (n_14867, n22815);
  and g37587 (n22816, n_14866, n_14867);
  not g37588 (n_14868, n22816);
  and g37589 (n22817, n_14866, n_14868);
  and g37590 (n22818, n_14867, n_14868);
  not g37591 (n_14869, n22817);
  not g37592 (n_14870, n22818);
  and g37593 (n22819, n_14869, n_14870);
  not g37594 (n_14871, n22575);
  not g37595 (n_14872, n22819);
  and g37596 (n22820, n_14871, n_14872);
  not g37597 (n_14873, n22820);
  and g37598 (n22821, n_14871, n_14873);
  and g37599 (n22822, n_14872, n_14873);
  not g37600 (n_14874, n22821);
  not g37601 (n_14875, n22822);
  and g37602 (n22823, n_14874, n_14875);
  and g37603 (n22824, n22642, n22724);
  not g37604 (n_14876, n22824);
  and g37605 (n22825, n_14822, n_14876);
  and g37606 (n22826, n4694, n22377);
  and g37607 (n22827, n4533, n22384);
  and g37608 (n22828, n4604, n22380);
  not g37609 (n_14877, n22827);
  not g37610 (n_14878, n22828);
  and g37611 (n22829, n_14877, n_14878);
  not g37612 (n_14879, n22826);
  and g37613 (n22830, n_14879, n22829);
  and g37614 (n22831, n_732, n22830);
  and g37615 (n22832, n_14542, n_14544);
  and g37616 (n22833, n_14543, n22436);
  not g37617 (n_14880, n22832);
  not g37618 (n_14881, n22833);
  and g37619 (n22834, n_14880, n_14881);
  and g37620 (n22835, n22830, n22834);
  not g37621 (n_14882, n22831);
  not g37622 (n_14883, n22835);
  and g37623 (n22836, n_14882, n_14883);
  not g37624 (n_14884, n22836);
  and g37625 (n22837, \a[23] , n_14884);
  and g37626 (n22838, n_27, n22836);
  not g37627 (n_14885, n22837);
  not g37628 (n_14886, n22838);
  and g37629 (n22839, n_14885, n_14886);
  not g37630 (n_14887, n22839);
  and g37631 (n22840, n22825, n_14887);
  and g37632 (n22841, n22661, n22722);
  not g37633 (n_14888, n22841);
  and g37634 (n22842, n_14819, n_14888);
  and g37635 (n22843, n4694, n22380);
  and g37636 (n22844, n4533, n22387);
  and g37637 (n22845, n4604, n22384);
  not g37638 (n_14889, n22844);
  not g37639 (n_14890, n22845);
  and g37640 (n22846, n_14889, n_14890);
  not g37641 (n_14891, n22843);
  and g37642 (n22847, n_14891, n22846);
  and g37643 (n22848, n_732, n22847);
  not g37644 (n_14892, n22431);
  and g37645 (n22849, n22429, n_14892);
  not g37646 (n_14893, n22849);
  and g37647 (n22850, n_14540, n_14893);
  not g37648 (n_14894, n22850);
  and g37649 (n22851, n22847, n_14894);
  not g37650 (n_14895, n22848);
  not g37651 (n_14896, n22851);
  and g37652 (n22852, n_14895, n_14896);
  not g37653 (n_14897, n22852);
  and g37654 (n22853, \a[23] , n_14897);
  and g37655 (n22854, n_27, n22852);
  not g37656 (n_14898, n22853);
  not g37657 (n_14899, n22854);
  and g37658 (n22855, n_14898, n_14899);
  not g37659 (n_14900, n22855);
  and g37660 (n22856, n22842, n_14900);
  and g37661 (n22857, n4694, n22384);
  and g37662 (n22858, n4533, n22390);
  and g37663 (n22859, n4604, n22387);
  and g37669 (n22862, n4536, n22806);
  not g37672 (n_14905, n22863);
  and g37673 (n22864, \a[23] , n_14905);
  not g37674 (n_14906, n22864);
  and g37675 (n22865, n_14905, n_14906);
  and g37676 (n22866, \a[23] , n_14906);
  not g37677 (n_14907, n22865);
  not g37678 (n_14908, n22866);
  and g37679 (n22867, n_14907, n_14908);
  not g37680 (n_14909, n22720);
  and g37681 (n22868, n22718, n_14909);
  not g37682 (n_14910, n22868);
  and g37683 (n22869, n_14816, n_14910);
  not g37684 (n_14911, n22867);
  and g37685 (n22870, n_14911, n22869);
  not g37686 (n_14912, n22870);
  and g37687 (n22871, n_14911, n_14912);
  and g37688 (n22872, n22869, n_14912);
  not g37689 (n_14913, n22871);
  not g37690 (n_14914, n22872);
  and g37691 (n22873, n_14913, n_14914);
  and g37692 (n22874, n_14809, n_14811);
  and g37693 (n22875, n_14810, n_14811);
  not g37694 (n_14915, n22874);
  not g37695 (n_14916, n22875);
  and g37696 (n22876, n_14915, n_14916);
  and g37697 (n22877, n4694, n22387);
  and g37698 (n22878, n4533, n22393);
  and g37699 (n22879, n4604, n22390);
  not g37700 (n_14917, n22878);
  not g37701 (n_14918, n22879);
  and g37702 (n22880, n_14917, n_14918);
  not g37703 (n_14919, n22877);
  and g37704 (n22881, n_14919, n22880);
  and g37705 (n22882, n_732, n22881);
  not g37706 (n_14920, n22582);
  and g37707 (n22883, n_14920, n22881);
  not g37708 (n_14921, n22882);
  not g37709 (n_14922, n22883);
  and g37710 (n22884, n_14921, n_14922);
  not g37711 (n_14923, n22884);
  and g37712 (n22885, \a[23] , n_14923);
  and g37713 (n22886, n_27, n22884);
  not g37714 (n_14924, n22885);
  not g37715 (n_14925, n22886);
  and g37716 (n22887, n_14924, n_14925);
  not g37717 (n_14926, n22876);
  not g37718 (n_14927, n22887);
  and g37719 (n22888, n_14926, n_14927);
  and g37720 (n22889, n4694, n22390);
  and g37721 (n22890, n4533, n22396);
  and g37722 (n22891, n4604, n22393);
  and g37728 (n22894, n4536, n22649);
  not g37731 (n_14932, n22895);
  and g37732 (n22896, \a[23] , n_14932);
  not g37733 (n_14933, n22896);
  and g37734 (n22897, n_14932, n_14933);
  and g37735 (n22898, \a[23] , n_14933);
  not g37736 (n_14934, n22897);
  not g37737 (n_14935, n22898);
  and g37738 (n22899, n_14934, n_14935);
  not g37739 (n_14936, n22689);
  and g37740 (n22900, n_14936, n22700);
  not g37741 (n_14937, n22701);
  not g37742 (n_14938, n22900);
  and g37743 (n22901, n_14937, n_14938);
  not g37744 (n_14939, n22899);
  and g37745 (n22902, n_14939, n22901);
  not g37746 (n_14940, n22902);
  and g37747 (n22903, n_14939, n_14940);
  and g37748 (n22904, n22901, n_14940);
  not g37749 (n_14941, n22903);
  not g37750 (n_14942, n22904);
  and g37751 (n22905, n_14941, n_14942);
  not g37752 (n_14943, n22679);
  and g37753 (n22906, n_14943, n22688);
  not g37754 (n_14944, n22906);
  and g37755 (n22907, n_14936, n_14944);
  and g37756 (n22908, n4694, n22393);
  and g37757 (n22909, n4533, n22399);
  and g37758 (n22910, n4604, n22396);
  not g37759 (n_14945, n22909);
  not g37760 (n_14946, n22910);
  and g37761 (n22911, n_14945, n_14946);
  not g37762 (n_14947, n22908);
  and g37763 (n22912, n_14947, n22911);
  and g37764 (n22913, n_732, n22912);
  and g37765 (n22914, n_14773, n22912);
  not g37766 (n_14948, n22913);
  not g37767 (n_14949, n22914);
  and g37768 (n22915, n_14948, n_14949);
  not g37769 (n_14950, n22915);
  and g37770 (n22916, \a[23] , n_14950);
  and g37771 (n22917, n_27, n22915);
  not g37772 (n_14951, n22916);
  not g37773 (n_14952, n22917);
  and g37774 (n22918, n_14951, n_14952);
  not g37775 (n_14953, n22918);
  and g37776 (n22919, n22907, n_14953);
  and g37777 (n22920, n_731, n_14508);
  not g37778 (n_14954, n22920);
  and g37779 (n22921, \a[23] , n_14954);
  and g37780 (n22922, n4604, n_14508);
  and g37781 (n22923, n4694, n22402);
  not g37782 (n_14955, n22922);
  not g37783 (n_14956, n22923);
  and g37784 (n22924, n_14955, n_14956);
  and g37785 (n22925, n4536, n_14720);
  not g37786 (n_14957, n22925);
  and g37787 (n22926, n22924, n_14957);
  not g37788 (n_14958, n22926);
  and g37789 (n22927, \a[23] , n_14958);
  not g37790 (n_14959, n22927);
  and g37791 (n22928, \a[23] , n_14959);
  and g37792 (n22929, n_14958, n_14959);
  not g37793 (n_14960, n22928);
  not g37794 (n_14961, n22929);
  and g37795 (n22930, n_14960, n_14961);
  not g37796 (n_14962, n22930);
  and g37797 (n22931, n22921, n_14962);
  and g37798 (n22932, n4694, n22399);
  and g37799 (n22933, n4533, n_14508);
  and g37800 (n22934, n4604, n22402);
  not g37801 (n_14963, n22933);
  not g37802 (n_14964, n22934);
  and g37803 (n22935, n_14963, n_14964);
  not g37804 (n_14965, n22932);
  and g37805 (n22936, n_14965, n22935);
  and g37806 (n22937, n_732, n22936);
  and g37807 (n22938, n22625, n22936);
  not g37808 (n_14966, n22937);
  not g37809 (n_14967, n22938);
  and g37810 (n22939, n_14966, n_14967);
  not g37811 (n_14968, n22939);
  and g37812 (n22940, \a[23] , n_14968);
  and g37813 (n22941, n_27, n22939);
  not g37814 (n_14969, n22940);
  not g37815 (n_14970, n22941);
  and g37816 (n22942, n_14969, n_14970);
  not g37817 (n_14971, n22942);
  and g37818 (n22943, n22931, n_14971);
  and g37819 (n22944, n22678, n22943);
  not g37820 (n_14972, n22944);
  and g37821 (n22945, n22943, n_14972);
  and g37822 (n22946, n22678, n_14972);
  not g37823 (n_14973, n22945);
  not g37824 (n_14974, n22946);
  and g37825 (n22947, n_14973, n_14974);
  and g37826 (n22948, n4694, n22396);
  and g37827 (n22949, n4533, n22402);
  and g37828 (n22950, n4604, n22399);
  and g37834 (n22953, n4536, n22595);
  not g37837 (n_14979, n22954);
  and g37838 (n22955, \a[23] , n_14979);
  not g37839 (n_14980, n22955);
  and g37840 (n22956, \a[23] , n_14980);
  and g37841 (n22957, n_14979, n_14980);
  not g37842 (n_14981, n22956);
  not g37843 (n_14982, n22957);
  and g37844 (n22958, n_14981, n_14982);
  not g37845 (n_14983, n22947);
  not g37846 (n_14984, n22958);
  and g37847 (n22959, n_14983, n_14984);
  not g37848 (n_14985, n22959);
  and g37849 (n22960, n_14972, n_14985);
  not g37850 (n_14986, n22907);
  and g37851 (n22961, n_14986, n22918);
  not g37852 (n_14987, n22919);
  not g37853 (n_14988, n22961);
  and g37854 (n22962, n_14987, n_14988);
  not g37855 (n_14989, n22960);
  and g37856 (n22963, n_14989, n22962);
  not g37857 (n_14990, n22963);
  and g37858 (n22964, n_14987, n_14990);
  not g37859 (n_14991, n22905);
  not g37860 (n_14992, n22964);
  and g37861 (n22965, n_14991, n_14992);
  not g37862 (n_14993, n22965);
  and g37863 (n22966, n_14940, n_14993);
  and g37864 (n22967, n22876, n22887);
  not g37865 (n_14994, n22888);
  not g37866 (n_14995, n22967);
  and g37867 (n22968, n_14994, n_14995);
  not g37868 (n_14996, n22966);
  and g37869 (n22969, n_14996, n22968);
  not g37870 (n_14997, n22969);
  and g37871 (n22970, n_14994, n_14997);
  not g37872 (n_14998, n22873);
  not g37873 (n_14999, n22970);
  and g37874 (n22971, n_14998, n_14999);
  not g37875 (n_15000, n22971);
  and g37876 (n22972, n_14912, n_15000);
  not g37877 (n_15001, n22856);
  and g37878 (n22973, n22842, n_15001);
  and g37879 (n22974, n_14900, n_15001);
  not g37880 (n_15002, n22973);
  not g37881 (n_15003, n22974);
  and g37882 (n22975, n_15002, n_15003);
  not g37883 (n_15004, n22972);
  not g37884 (n_15005, n22975);
  and g37885 (n22976, n_15004, n_15005);
  not g37886 (n_15006, n22976);
  and g37887 (n22977, n_15001, n_15006);
  not g37888 (n_15007, n22825);
  and g37889 (n22978, n_15007, n22839);
  not g37890 (n_15008, n22840);
  not g37891 (n_15009, n22978);
  and g37892 (n22979, n_15008, n_15009);
  not g37893 (n_15010, n22977);
  and g37894 (n22980, n_15010, n22979);
  not g37895 (n_15011, n22980);
  and g37896 (n22981, n_15008, n_15011);
  and g37897 (n22982, n22823, n22981);
  not g37898 (n_15012, n22823);
  not g37899 (n_15013, n22981);
  and g37900 (n22983, n_15012, n_15013);
  not g37901 (n_15014, n22982);
  not g37902 (n_15015, n22983);
  and g37903 (n22984, n_15014, n_15015);
  and g37904 (n22985, n5496, n22365);
  and g37905 (n22986, n4935, n22371);
  and g37906 (n22987, n5407, n22368);
  not g37907 (n_15016, n22986);
  not g37908 (n_15017, n22987);
  and g37909 (n22988, n_15016, n_15017);
  not g37910 (n_15018, n22985);
  and g37911 (n22989, n_15018, n22988);
  and g37912 (n22990, n_1011, n22989);
  and g37913 (n22991, n_14561, n_14564);
  and g37914 (n22992, n_14562, n22452);
  not g37915 (n_15019, n22991);
  not g37916 (n_15020, n22992);
  and g37917 (n22993, n_15019, n_15020);
  and g37918 (n22994, n22989, n22993);
  not g37919 (n_15021, n22990);
  not g37920 (n_15022, n22994);
  and g37921 (n22995, n_15021, n_15022);
  not g37922 (n_15023, n22995);
  and g37923 (n22996, \a[20] , n_15023);
  and g37924 (n22997, n_435, n22995);
  not g37925 (n_15024, n22996);
  not g37926 (n_15025, n22997);
  and g37927 (n22998, n_15024, n_15025);
  not g37928 (n_15026, n22998);
  and g37929 (n22999, n22984, n_15026);
  and g37930 (n23000, n5496, n22368);
  and g37931 (n23001, n4935, n22374);
  and g37932 (n23002, n5407, n22371);
  not g37938 (n_15030, n22446);
  and g37939 (n23005, n22444, n_15030);
  not g37940 (n_15031, n23005);
  and g37941 (n23006, n_14559, n_15031);
  and g37942 (n23007, n4938, n23006);
  not g37945 (n_15033, n23008);
  and g37946 (n23009, \a[20] , n_15033);
  not g37947 (n_15034, n23009);
  and g37948 (n23010, n_15033, n_15034);
  and g37949 (n23011, \a[20] , n_15034);
  not g37950 (n_15035, n23010);
  not g37951 (n_15036, n23011);
  and g37952 (n23012, n_15035, n_15036);
  not g37953 (n_15037, n22979);
  and g37954 (n23013, n22977, n_15037);
  not g37955 (n_15038, n23013);
  and g37956 (n23014, n_15011, n_15038);
  not g37957 (n_15039, n23012);
  and g37958 (n23015, n_15039, n23014);
  not g37959 (n_15040, n23015);
  and g37960 (n23016, n_15039, n_15040);
  and g37961 (n23017, n23014, n_15040);
  not g37962 (n_15041, n23016);
  not g37963 (n_15042, n23017);
  and g37964 (n23018, n_15041, n_15042);
  and g37965 (n23019, n5496, n22371);
  and g37966 (n23020, n4935, n22377);
  and g37967 (n23021, n5407, n22374);
  not g37973 (n_15046, n22442);
  and g37974 (n23024, n22440, n_15046);
  not g37975 (n_15047, n23024);
  and g37976 (n23025, n_14554, n_15047);
  and g37977 (n23026, n4938, n23025);
  not g37980 (n_15049, n23027);
  and g37981 (n23028, \a[20] , n_15049);
  not g37982 (n_15050, n23028);
  and g37983 (n23029, n_15049, n_15050);
  and g37984 (n23030, \a[20] , n_15050);
  not g37985 (n_15051, n23029);
  not g37986 (n_15052, n23030);
  and g37987 (n23031, n_15051, n_15052);
  and g37988 (n23032, n_15004, n_15006);
  and g37989 (n23033, n_15005, n_15006);
  not g37990 (n_15053, n23032);
  not g37991 (n_15054, n23033);
  and g37992 (n23034, n_15053, n_15054);
  not g37993 (n_15055, n23031);
  not g37994 (n_15056, n23034);
  and g37995 (n23035, n_15055, n_15056);
  not g37996 (n_15057, n23035);
  and g37997 (n23036, n_15055, n_15057);
  and g37998 (n23037, n_15056, n_15057);
  not g37999 (n_15058, n23036);
  not g38000 (n_15059, n23037);
  and g38001 (n23038, n_15058, n_15059);
  and g38002 (n23039, n22873, n22970);
  not g38003 (n_15060, n23039);
  and g38004 (n23040, n_15000, n_15060);
  and g38005 (n23041, n5496, n22374);
  and g38006 (n23042, n4935, n22380);
  and g38007 (n23043, n5407, n22377);
  not g38008 (n_15061, n23042);
  not g38009 (n_15062, n23043);
  and g38010 (n23044, n_15061, n_15062);
  not g38011 (n_15063, n23041);
  and g38012 (n23045, n_15063, n23044);
  and g38013 (n23046, n_1011, n23045);
  not g38014 (n_15064, n22569);
  and g38015 (n23047, n_15064, n23045);
  not g38016 (n_15065, n23046);
  not g38017 (n_15066, n23047);
  and g38018 (n23048, n_15065, n_15066);
  not g38019 (n_15067, n23048);
  and g38020 (n23049, \a[20] , n_15067);
  and g38021 (n23050, n_435, n23048);
  not g38022 (n_15068, n23049);
  not g38023 (n_15069, n23050);
  and g38024 (n23051, n_15068, n_15069);
  not g38025 (n_15070, n23051);
  and g38026 (n23052, n23040, n_15070);
  not g38027 (n_15071, n22968);
  and g38028 (n23053, n22966, n_15071);
  not g38029 (n_15072, n23053);
  and g38030 (n23054, n_14997, n_15072);
  and g38031 (n23055, n5496, n22377);
  and g38032 (n23056, n4935, n22384);
  and g38033 (n23057, n5407, n22380);
  not g38034 (n_15073, n23056);
  not g38035 (n_15074, n23057);
  and g38036 (n23058, n_15073, n_15074);
  not g38037 (n_15075, n23055);
  and g38038 (n23059, n_15075, n23058);
  and g38039 (n23060, n_1011, n23059);
  and g38040 (n23061, n22834, n23059);
  not g38041 (n_15076, n23060);
  not g38042 (n_15077, n23061);
  and g38043 (n23062, n_15076, n_15077);
  not g38044 (n_15078, n23062);
  and g38045 (n23063, \a[20] , n_15078);
  and g38046 (n23064, n_435, n23062);
  not g38047 (n_15079, n23063);
  not g38048 (n_15080, n23064);
  and g38049 (n23065, n_15079, n_15080);
  not g38050 (n_15081, n23065);
  and g38051 (n23066, n23054, n_15081);
  and g38052 (n23067, n22905, n22964);
  not g38053 (n_15082, n23067);
  and g38054 (n23068, n_14993, n_15082);
  and g38055 (n23069, n5496, n22380);
  and g38056 (n23070, n4935, n22387);
  and g38057 (n23071, n5407, n22384);
  not g38058 (n_15083, n23070);
  not g38059 (n_15084, n23071);
  and g38060 (n23072, n_15083, n_15084);
  not g38061 (n_15085, n23069);
  and g38062 (n23073, n_15085, n23072);
  and g38063 (n23074, n_1011, n23073);
  and g38064 (n23075, n_14894, n23073);
  not g38065 (n_15086, n23074);
  not g38066 (n_15087, n23075);
  and g38067 (n23076, n_15086, n_15087);
  not g38068 (n_15088, n23076);
  and g38069 (n23077, \a[20] , n_15088);
  and g38070 (n23078, n_435, n23076);
  not g38071 (n_15089, n23077);
  not g38072 (n_15090, n23078);
  and g38073 (n23079, n_15089, n_15090);
  not g38074 (n_15091, n23079);
  and g38075 (n23080, n23068, n_15091);
  and g38076 (n23081, n5496, n22384);
  and g38077 (n23082, n4935, n22390);
  and g38078 (n23083, n5407, n22387);
  and g38084 (n23086, n4938, n22806);
  not g38087 (n_15096, n23087);
  and g38088 (n23088, \a[20] , n_15096);
  not g38089 (n_15097, n23088);
  and g38090 (n23089, n_15096, n_15097);
  and g38091 (n23090, \a[20] , n_15097);
  not g38092 (n_15098, n23089);
  not g38093 (n_15099, n23090);
  and g38094 (n23091, n_15098, n_15099);
  not g38095 (n_15100, n22962);
  and g38096 (n23092, n22960, n_15100);
  not g38097 (n_15101, n23092);
  and g38098 (n23093, n_14990, n_15101);
  not g38099 (n_15102, n23091);
  and g38100 (n23094, n_15102, n23093);
  not g38101 (n_15103, n23094);
  and g38102 (n23095, n_15102, n_15103);
  and g38103 (n23096, n23093, n_15103);
  not g38104 (n_15104, n23095);
  not g38105 (n_15105, n23096);
  and g38106 (n23097, n_15104, n_15105);
  and g38107 (n23098, n_14983, n_14985);
  and g38108 (n23099, n_14984, n_14985);
  not g38109 (n_15106, n23098);
  not g38110 (n_15107, n23099);
  and g38111 (n23100, n_15106, n_15107);
  and g38112 (n23101, n5496, n22387);
  and g38113 (n23102, n4935, n22393);
  and g38114 (n23103, n5407, n22390);
  not g38115 (n_15108, n23102);
  not g38116 (n_15109, n23103);
  and g38117 (n23104, n_15108, n_15109);
  not g38118 (n_15110, n23101);
  and g38119 (n23105, n_15110, n23104);
  and g38120 (n23106, n_1011, n23105);
  and g38121 (n23107, n_14920, n23105);
  not g38122 (n_15111, n23106);
  not g38123 (n_15112, n23107);
  and g38124 (n23108, n_15111, n_15112);
  not g38125 (n_15113, n23108);
  and g38126 (n23109, \a[20] , n_15113);
  and g38127 (n23110, n_435, n23108);
  not g38128 (n_15114, n23109);
  not g38129 (n_15115, n23110);
  and g38130 (n23111, n_15114, n_15115);
  not g38131 (n_15116, n23100);
  not g38132 (n_15117, n23111);
  and g38133 (n23112, n_15116, n_15117);
  and g38134 (n23113, n5496, n22390);
  and g38135 (n23114, n4935, n22396);
  and g38136 (n23115, n5407, n22393);
  and g38142 (n23118, n4938, n22649);
  not g38145 (n_15122, n23119);
  and g38146 (n23120, \a[20] , n_15122);
  not g38147 (n_15123, n23120);
  and g38148 (n23121, n_15122, n_15123);
  and g38149 (n23122, \a[20] , n_15123);
  not g38150 (n_15124, n23121);
  not g38151 (n_15125, n23122);
  and g38152 (n23123, n_15124, n_15125);
  not g38153 (n_15126, n22931);
  and g38154 (n23124, n_15126, n22942);
  not g38155 (n_15127, n22943);
  not g38156 (n_15128, n23124);
  and g38157 (n23125, n_15127, n_15128);
  not g38158 (n_15129, n23123);
  and g38159 (n23126, n_15129, n23125);
  not g38160 (n_15130, n23126);
  and g38161 (n23127, n_15129, n_15130);
  and g38162 (n23128, n23125, n_15130);
  not g38163 (n_15131, n23127);
  not g38164 (n_15132, n23128);
  and g38165 (n23129, n_15131, n_15132);
  not g38166 (n_15133, n22921);
  and g38167 (n23130, n_15133, n22930);
  not g38168 (n_15134, n23130);
  and g38169 (n23131, n_15126, n_15134);
  and g38170 (n23132, n5496, n22393);
  and g38171 (n23133, n4935, n22399);
  and g38172 (n23134, n5407, n22396);
  not g38173 (n_15135, n23133);
  not g38174 (n_15136, n23134);
  and g38175 (n23135, n_15135, n_15136);
  not g38176 (n_15137, n23132);
  and g38177 (n23136, n_15137, n23135);
  and g38178 (n23137, n_1011, n23136);
  and g38179 (n23138, n_14773, n23136);
  not g38180 (n_15138, n23137);
  not g38181 (n_15139, n23138);
  and g38182 (n23139, n_15138, n_15139);
  not g38183 (n_15140, n23139);
  and g38184 (n23140, \a[20] , n_15140);
  and g38185 (n23141, n_435, n23139);
  not g38186 (n_15141, n23140);
  not g38187 (n_15142, n23141);
  and g38188 (n23142, n_15141, n_15142);
  not g38189 (n_15143, n23142);
  and g38190 (n23143, n23131, n_15143);
  and g38191 (n23144, n5407, n_14508);
  and g38192 (n23145, n5496, n22402);
  not g38193 (n_15144, n23144);
  not g38194 (n_15145, n23145);
  and g38195 (n23146, n_15144, n_15145);
  and g38196 (n23147, n4938, n_14720);
  not g38197 (n_15146, n23147);
  and g38198 (n23148, n23146, n_15146);
  not g38199 (n_15147, n23148);
  and g38200 (n23149, \a[20] , n_15147);
  not g38201 (n_15148, n23149);
  and g38202 (n23150, \a[20] , n_15148);
  and g38203 (n23151, n_15147, n_15148);
  not g38204 (n_15149, n23150);
  not g38205 (n_15150, n23151);
  and g38206 (n23152, n_15149, n_15150);
  and g38207 (n23153, n_1010, n_14508);
  not g38208 (n_15151, n23153);
  and g38209 (n23154, \a[20] , n_15151);
  not g38210 (n_15152, n23152);
  and g38211 (n23155, n_15152, n23154);
  and g38212 (n23156, n5496, n22399);
  and g38213 (n23157, n4935, n_14508);
  and g38214 (n23158, n5407, n22402);
  not g38215 (n_15153, n23157);
  not g38216 (n_15154, n23158);
  and g38217 (n23159, n_15153, n_15154);
  not g38218 (n_15155, n23156);
  and g38219 (n23160, n_15155, n23159);
  and g38220 (n23161, n_1011, n23160);
  and g38221 (n23162, n22625, n23160);
  not g38222 (n_15156, n23161);
  not g38223 (n_15157, n23162);
  and g38224 (n23163, n_15156, n_15157);
  not g38225 (n_15158, n23163);
  and g38226 (n23164, \a[20] , n_15158);
  and g38227 (n23165, n_435, n23163);
  not g38228 (n_15159, n23164);
  not g38229 (n_15160, n23165);
  and g38230 (n23166, n_15159, n_15160);
  not g38231 (n_15161, n23166);
  and g38232 (n23167, n23155, n_15161);
  and g38233 (n23168, n22920, n23167);
  not g38234 (n_15162, n23168);
  and g38235 (n23169, n23167, n_15162);
  and g38236 (n23170, n22920, n_15162);
  not g38237 (n_15163, n23169);
  not g38238 (n_15164, n23170);
  and g38239 (n23171, n_15163, n_15164);
  and g38240 (n23172, n5496, n22396);
  and g38241 (n23173, n4935, n22402);
  and g38242 (n23174, n5407, n22399);
  and g38248 (n23177, n4938, n22595);
  not g38251 (n_15169, n23178);
  and g38252 (n23179, \a[20] , n_15169);
  not g38253 (n_15170, n23179);
  and g38254 (n23180, \a[20] , n_15170);
  and g38255 (n23181, n_15169, n_15170);
  not g38256 (n_15171, n23180);
  not g38257 (n_15172, n23181);
  and g38258 (n23182, n_15171, n_15172);
  not g38259 (n_15173, n23171);
  not g38260 (n_15174, n23182);
  and g38261 (n23183, n_15173, n_15174);
  not g38262 (n_15175, n23183);
  and g38263 (n23184, n_15162, n_15175);
  not g38264 (n_15176, n23131);
  and g38265 (n23185, n_15176, n23142);
  not g38266 (n_15177, n23143);
  not g38267 (n_15178, n23185);
  and g38268 (n23186, n_15177, n_15178);
  not g38269 (n_15179, n23184);
  and g38270 (n23187, n_15179, n23186);
  not g38271 (n_15180, n23187);
  and g38272 (n23188, n_15177, n_15180);
  not g38273 (n_15181, n23129);
  not g38274 (n_15182, n23188);
  and g38275 (n23189, n_15181, n_15182);
  not g38276 (n_15183, n23189);
  and g38277 (n23190, n_15130, n_15183);
  and g38278 (n23191, n23100, n23111);
  not g38279 (n_15184, n23112);
  not g38280 (n_15185, n23191);
  and g38281 (n23192, n_15184, n_15185);
  not g38282 (n_15186, n23190);
  and g38283 (n23193, n_15186, n23192);
  not g38284 (n_15187, n23193);
  and g38285 (n23194, n_15184, n_15187);
  not g38286 (n_15188, n23097);
  not g38287 (n_15189, n23194);
  and g38288 (n23195, n_15188, n_15189);
  not g38289 (n_15190, n23195);
  and g38290 (n23196, n_15103, n_15190);
  not g38291 (n_15191, n23080);
  and g38292 (n23197, n23068, n_15191);
  and g38293 (n23198, n_15091, n_15191);
  not g38294 (n_15192, n23197);
  not g38295 (n_15193, n23198);
  and g38296 (n23199, n_15192, n_15193);
  not g38297 (n_15194, n23196);
  not g38298 (n_15195, n23199);
  and g38299 (n23200, n_15194, n_15195);
  not g38300 (n_15196, n23200);
  and g38301 (n23201, n_15191, n_15196);
  not g38302 (n_15197, n23066);
  and g38303 (n23202, n23054, n_15197);
  and g38304 (n23203, n_15081, n_15197);
  not g38305 (n_15198, n23202);
  not g38306 (n_15199, n23203);
  and g38307 (n23204, n_15198, n_15199);
  not g38308 (n_15200, n23201);
  not g38309 (n_15201, n23204);
  and g38310 (n23205, n_15200, n_15201);
  not g38311 (n_15202, n23205);
  and g38312 (n23206, n_15197, n_15202);
  not g38313 (n_15203, n23040);
  and g38314 (n23207, n_15203, n23051);
  not g38315 (n_15204, n23052);
  not g38316 (n_15205, n23207);
  and g38317 (n23208, n_15204, n_15205);
  not g38318 (n_15206, n23206);
  and g38319 (n23209, n_15206, n23208);
  not g38320 (n_15207, n23209);
  and g38321 (n23210, n_15204, n_15207);
  not g38322 (n_15208, n23038);
  not g38323 (n_15209, n23210);
  and g38324 (n23211, n_15208, n_15209);
  not g38325 (n_15210, n23211);
  and g38326 (n23212, n_15057, n_15210);
  not g38327 (n_15211, n23018);
  not g38328 (n_15212, n23212);
  and g38329 (n23213, n_15211, n_15212);
  not g38330 (n_15213, n23213);
  and g38331 (n23214, n_15040, n_15213);
  not g38332 (n_15214, n22999);
  and g38333 (n23215, n22984, n_15214);
  and g38334 (n23216, n_15026, n_15214);
  not g38335 (n_15215, n23215);
  not g38336 (n_15216, n23216);
  and g38337 (n23217, n_15215, n_15216);
  not g38338 (n_15217, n23214);
  not g38339 (n_15218, n23217);
  and g38340 (n23218, n_15217, n_15218);
  not g38341 (n_15219, n23218);
  and g38342 (n23219, n_15214, n_15219);
  and g38343 (n23220, n4694, n22371);
  and g38344 (n23221, n4533, n22377);
  and g38345 (n23222, n4604, n22374);
  and g38351 (n23225, n4536, n23025);
  not g38354 (n_15224, n23226);
  and g38355 (n23227, \a[23] , n_15224);
  not g38356 (n_15225, n23227);
  and g38357 (n23228, n_15224, n_15225);
  and g38358 (n23229, \a[23] , n_15225);
  not g38359 (n_15226, n23228);
  not g38360 (n_15227, n23229);
  and g38361 (n23230, n_15226, n_15227);
  and g38362 (n23231, n_14863, n_14868);
  and g38363 (n23232, n3457, n22390);
  and g38364 (n23233, n3542, n22396);
  and g38365 (n23234, n3606, n22393);
  and g38371 (n23237, n3368, n22649);
  not g38374 (n_15232, n23238);
  and g38375 (n23239, \a[29] , n_15232);
  not g38376 (n_15233, n23239);
  and g38377 (n23240, n_15232, n_15233);
  and g38378 (n23241, \a[29] , n_15233);
  not g38379 (n_15234, n23240);
  not g38380 (n_15235, n23241);
  and g38381 (n23242, n_15234, n_15235);
  not g38382 (n_15236, n22625);
  and g38383 (n23243, n75, n_15236);
  and g38384 (n23244, n3020, n22399);
  and g38385 (n23245, n3023, n_14508);
  and g38386 (n23246, n3028, n22402);
  and g38394 (n23250, n_91, n_139);
  and g38395 (n23251, n_168, n23250);
  not g38414 (n_15241, n23269);
  and g38415 (n23270, n22785, n_15241);
  and g38416 (n23271, n_14836, n23269);
  not g38417 (n_15242, n23270);
  not g38418 (n_15243, n23271);
  and g38419 (n23272, n_15242, n_15243);
  not g38420 (n_15244, n23249);
  and g38421 (n23273, n_15244, n23272);
  not g38422 (n_15245, n23273);
  and g38423 (n23274, n_15244, n_15245);
  and g38424 (n23275, n23272, n_15245);
  not g38425 (n_15246, n23274);
  not g38426 (n_15247, n23275);
  and g38427 (n23276, n_15246, n_15247);
  not g38428 (n_15248, n23242);
  not g38429 (n_15249, n23276);
  and g38430 (n23277, n_15248, n_15249);
  not g38431 (n_15250, n23277);
  and g38432 (n23278, n_15248, n_15250);
  and g38433 (n23279, n_15249, n_15250);
  not g38434 (n_15251, n23278);
  not g38435 (n_15252, n23279);
  and g38436 (n23280, n_15251, n_15252);
  and g38437 (n23281, n_14841, n_14847);
  and g38438 (n23282, n23280, n23281);
  not g38439 (n_15253, n23280);
  not g38440 (n_15254, n23281);
  and g38441 (n23283, n_15253, n_15254);
  not g38442 (n_15255, n23282);
  not g38443 (n_15256, n23283);
  and g38444 (n23284, n_15255, n_15256);
  and g38445 (n23285, n3884, n22380);
  and g38446 (n23286, n3967, n22387);
  and g38447 (n23287, n4046, n22384);
  not g38448 (n_15257, n23286);
  not g38449 (n_15258, n23287);
  and g38450 (n23288, n_15257, n_15258);
  not g38451 (n_15259, n23285);
  and g38452 (n23289, n_15259, n23288);
  and g38453 (n23290, n_750, n23289);
  and g38454 (n23291, n_14894, n23289);
  not g38455 (n_15260, n23290);
  not g38456 (n_15261, n23291);
  and g38457 (n23292, n_15260, n_15261);
  not g38458 (n_15262, n23292);
  and g38459 (n23293, \a[26] , n_15262);
  and g38460 (n23294, n_33, n23292);
  not g38461 (n_15263, n23293);
  not g38462 (n_15264, n23294);
  and g38463 (n23295, n_15263, n_15264);
  not g38464 (n_15265, n23295);
  and g38465 (n23296, n23284, n_15265);
  not g38466 (n_15266, n23296);
  and g38467 (n23297, n23284, n_15266);
  and g38468 (n23298, n_15265, n_15266);
  not g38469 (n_15267, n23297);
  not g38470 (n_15268, n23298);
  and g38471 (n23299, n_15267, n_15268);
  not g38472 (n_15269, n23231);
  not g38473 (n_15270, n23299);
  and g38474 (n23300, n_15269, n_15270);
  not g38475 (n_15271, n23300);
  and g38476 (n23301, n_15269, n_15271);
  and g38477 (n23302, n_15270, n_15271);
  not g38478 (n_15272, n23301);
  not g38479 (n_15273, n23302);
  and g38480 (n23303, n_15272, n_15273);
  not g38481 (n_15274, n23230);
  not g38482 (n_15275, n23303);
  and g38483 (n23304, n_15274, n_15275);
  not g38484 (n_15276, n23304);
  and g38485 (n23305, n_15274, n_15276);
  and g38486 (n23306, n_15275, n_15276);
  not g38487 (n_15277, n23305);
  not g38488 (n_15278, n23306);
  and g38489 (n23307, n_15277, n_15278);
  and g38490 (n23308, n_14873, n_15015);
  and g38491 (n23309, n23307, n23308);
  not g38492 (n_15279, n23307);
  not g38493 (n_15280, n23308);
  and g38494 (n23310, n_15279, n_15280);
  not g38495 (n_15281, n23309);
  not g38496 (n_15282, n23310);
  and g38497 (n23311, n_15281, n_15282);
  and g38498 (n23312, n5496, n22362);
  and g38499 (n23313, n4935, n22368);
  and g38500 (n23314, n5407, n22365);
  not g38501 (n_15283, n23313);
  not g38502 (n_15284, n23314);
  and g38503 (n23315, n_15283, n_15284);
  not g38504 (n_15285, n23312);
  and g38505 (n23316, n_15285, n23315);
  and g38506 (n23317, n_1011, n23316);
  and g38507 (n23318, n_14566, n_14569);
  and g38508 (n23319, n_14567, n22456);
  not g38509 (n_15286, n23318);
  not g38510 (n_15287, n23319);
  and g38511 (n23320, n_15286, n_15287);
  and g38512 (n23321, n23316, n23320);
  not g38513 (n_15288, n23317);
  not g38514 (n_15289, n23321);
  and g38515 (n23322, n_15288, n_15289);
  not g38516 (n_15290, n23322);
  and g38517 (n23323, \a[20] , n_15290);
  and g38518 (n23324, n_435, n23322);
  not g38519 (n_15291, n23323);
  not g38520 (n_15292, n23324);
  and g38521 (n23325, n_15291, n_15292);
  not g38522 (n_15293, n23325);
  and g38523 (n23326, n23311, n_15293);
  not g38524 (n_15294, n23326);
  and g38525 (n23327, n23311, n_15294);
  and g38526 (n23328, n_15293, n_15294);
  not g38527 (n_15295, n23327);
  not g38528 (n_15296, n23328);
  and g38529 (n23329, n_15295, n_15296);
  not g38530 (n_15297, n23219);
  not g38531 (n_15298, n23329);
  and g38532 (n23330, n_15297, n_15298);
  not g38533 (n_15299, n23330);
  and g38534 (n23331, n_15297, n_15299);
  and g38535 (n23332, n_15298, n_15299);
  not g38536 (n_15300, n23331);
  not g38537 (n_15301, n23332);
  and g38538 (n23333, n_15300, n_15301);
  not g38539 (n_15302, n22562);
  not g38540 (n_15303, n23333);
  and g38541 (n23334, n_15302, n_15303);
  not g38542 (n_15304, n23334);
  and g38543 (n23335, n_15302, n_15304);
  and g38544 (n23336, n_15303, n_15304);
  not g38545 (n_15305, n23335);
  not g38546 (n_15306, n23336);
  and g38547 (n23337, n_15305, n_15306);
  and g38548 (n23338, n6233, n22356);
  and g38549 (n23339, n5663, n22362);
  and g38550 (n23340, n5939, n22359);
  and g38556 (n23343, n_14576, n_14579);
  and g38557 (n23344, n_14577, n22464);
  not g38558 (n_15310, n23343);
  not g38559 (n_15311, n23344);
  and g38560 (n23345, n_15310, n_15311);
  not g38561 (n_15312, n23345);
  and g38562 (n23346, n5666, n_15312);
  not g38565 (n_15314, n23347);
  and g38566 (n23348, \a[17] , n_15314);
  not g38567 (n_15315, n23348);
  and g38568 (n23349, n_15314, n_15315);
  and g38569 (n23350, \a[17] , n_15315);
  not g38570 (n_15316, n23349);
  not g38571 (n_15317, n23350);
  and g38572 (n23351, n_15316, n_15317);
  and g38573 (n23352, n_15217, n_15219);
  and g38574 (n23353, n_15218, n_15219);
  not g38575 (n_15318, n23352);
  not g38576 (n_15319, n23353);
  and g38577 (n23354, n_15318, n_15319);
  not g38578 (n_15320, n23351);
  not g38579 (n_15321, n23354);
  and g38580 (n23355, n_15320, n_15321);
  not g38581 (n_15322, n23355);
  and g38582 (n23356, n_15320, n_15322);
  and g38583 (n23357, n_15321, n_15322);
  not g38584 (n_15323, n23356);
  not g38585 (n_15324, n23357);
  and g38586 (n23358, n_15323, n_15324);
  and g38587 (n23359, n23018, n23212);
  not g38588 (n_15325, n23359);
  and g38589 (n23360, n_15213, n_15325);
  and g38590 (n23361, n6233, n22359);
  and g38591 (n23362, n5663, n22365);
  and g38592 (n23363, n5939, n22362);
  not g38593 (n_15326, n23362);
  not g38594 (n_15327, n23363);
  and g38595 (n23364, n_15326, n_15327);
  not g38596 (n_15328, n23361);
  and g38597 (n23365, n_15328, n23364);
  and g38598 (n23366, n_1409, n23365);
  not g38599 (n_15329, n22458);
  and g38600 (n23367, n22456, n_15329);
  not g38601 (n_15330, n23367);
  and g38602 (n23368, n_14574, n_15330);
  not g38603 (n_15331, n23368);
  and g38604 (n23369, n23365, n_15331);
  not g38605 (n_15332, n23366);
  not g38606 (n_15333, n23369);
  and g38607 (n23370, n_15332, n_15333);
  not g38608 (n_15334, n23370);
  and g38609 (n23371, \a[17] , n_15334);
  and g38610 (n23372, n_617, n23370);
  not g38611 (n_15335, n23371);
  not g38612 (n_15336, n23372);
  and g38613 (n23373, n_15335, n_15336);
  not g38614 (n_15337, n23373);
  and g38615 (n23374, n23360, n_15337);
  and g38616 (n23375, n23038, n23210);
  not g38617 (n_15338, n23375);
  and g38618 (n23376, n_15210, n_15338);
  and g38619 (n23377, n6233, n22362);
  and g38620 (n23378, n5663, n22368);
  and g38621 (n23379, n5939, n22365);
  not g38622 (n_15339, n23378);
  not g38623 (n_15340, n23379);
  and g38624 (n23380, n_15339, n_15340);
  not g38625 (n_15341, n23377);
  and g38626 (n23381, n_15341, n23380);
  and g38627 (n23382, n_1409, n23381);
  and g38628 (n23383, n23320, n23381);
  not g38629 (n_15342, n23382);
  not g38630 (n_15343, n23383);
  and g38631 (n23384, n_15342, n_15343);
  not g38632 (n_15344, n23384);
  and g38633 (n23385, \a[17] , n_15344);
  and g38634 (n23386, n_617, n23384);
  not g38635 (n_15345, n23385);
  not g38636 (n_15346, n23386);
  and g38637 (n23387, n_15345, n_15346);
  not g38638 (n_15347, n23387);
  and g38639 (n23388, n23376, n_15347);
  and g38640 (n23389, n6233, n22365);
  and g38641 (n23390, n5663, n22371);
  and g38642 (n23391, n5939, n22368);
  not g38648 (n_15351, n22993);
  and g38649 (n23394, n5666, n_15351);
  not g38652 (n_15353, n23395);
  and g38653 (n23396, \a[17] , n_15353);
  not g38654 (n_15354, n23396);
  and g38655 (n23397, n_15353, n_15354);
  and g38656 (n23398, \a[17] , n_15354);
  not g38657 (n_15355, n23397);
  not g38658 (n_15356, n23398);
  and g38659 (n23399, n_15355, n_15356);
  not g38660 (n_15357, n23208);
  and g38661 (n23400, n23206, n_15357);
  not g38662 (n_15358, n23400);
  and g38663 (n23401, n_15207, n_15358);
  not g38664 (n_15359, n23399);
  and g38665 (n23402, n_15359, n23401);
  not g38666 (n_15360, n23402);
  and g38667 (n23403, n_15359, n_15360);
  and g38668 (n23404, n23401, n_15360);
  not g38669 (n_15361, n23403);
  not g38670 (n_15362, n23404);
  and g38671 (n23405, n_15361, n_15362);
  and g38672 (n23406, n6233, n22368);
  and g38673 (n23407, n5663, n22374);
  and g38674 (n23408, n5939, n22371);
  and g38680 (n23411, n5666, n23006);
  not g38683 (n_15367, n23412);
  and g38684 (n23413, \a[17] , n_15367);
  not g38685 (n_15368, n23413);
  and g38686 (n23414, n_15367, n_15368);
  and g38687 (n23415, \a[17] , n_15368);
  not g38688 (n_15369, n23414);
  not g38689 (n_15370, n23415);
  and g38690 (n23416, n_15369, n_15370);
  and g38691 (n23417, n_15200, n_15202);
  and g38692 (n23418, n_15201, n_15202);
  not g38693 (n_15371, n23417);
  not g38694 (n_15372, n23418);
  and g38695 (n23419, n_15371, n_15372);
  not g38696 (n_15373, n23416);
  not g38697 (n_15374, n23419);
  and g38698 (n23420, n_15373, n_15374);
  not g38699 (n_15375, n23420);
  and g38700 (n23421, n_15373, n_15375);
  and g38701 (n23422, n_15374, n_15375);
  not g38702 (n_15376, n23421);
  not g38703 (n_15377, n23422);
  and g38704 (n23423, n_15376, n_15377);
  and g38705 (n23424, n6233, n22371);
  and g38706 (n23425, n5663, n22377);
  and g38707 (n23426, n5939, n22374);
  and g38713 (n23429, n5666, n23025);
  not g38716 (n_15382, n23430);
  and g38717 (n23431, \a[17] , n_15382);
  not g38718 (n_15383, n23431);
  and g38719 (n23432, n_15382, n_15383);
  and g38720 (n23433, \a[17] , n_15383);
  not g38721 (n_15384, n23432);
  not g38722 (n_15385, n23433);
  and g38723 (n23434, n_15384, n_15385);
  and g38724 (n23435, n_15194, n_15196);
  and g38725 (n23436, n_15195, n_15196);
  not g38726 (n_15386, n23435);
  not g38727 (n_15387, n23436);
  and g38728 (n23437, n_15386, n_15387);
  not g38729 (n_15388, n23434);
  not g38730 (n_15389, n23437);
  and g38731 (n23438, n_15388, n_15389);
  not g38732 (n_15390, n23438);
  and g38733 (n23439, n_15388, n_15390);
  and g38734 (n23440, n_15389, n_15390);
  not g38735 (n_15391, n23439);
  not g38736 (n_15392, n23440);
  and g38737 (n23441, n_15391, n_15392);
  and g38738 (n23442, n23097, n23194);
  not g38739 (n_15393, n23442);
  and g38740 (n23443, n_15190, n_15393);
  and g38741 (n23444, n6233, n22374);
  and g38742 (n23445, n5663, n22380);
  and g38743 (n23446, n5939, n22377);
  not g38744 (n_15394, n23445);
  not g38745 (n_15395, n23446);
  and g38746 (n23447, n_15394, n_15395);
  not g38747 (n_15396, n23444);
  and g38748 (n23448, n_15396, n23447);
  and g38749 (n23449, n_1409, n23448);
  and g38750 (n23450, n_15064, n23448);
  not g38751 (n_15397, n23449);
  not g38752 (n_15398, n23450);
  and g38753 (n23451, n_15397, n_15398);
  not g38754 (n_15399, n23451);
  and g38755 (n23452, \a[17] , n_15399);
  and g38756 (n23453, n_617, n23451);
  not g38757 (n_15400, n23452);
  not g38758 (n_15401, n23453);
  and g38759 (n23454, n_15400, n_15401);
  not g38760 (n_15402, n23454);
  and g38761 (n23455, n23443, n_15402);
  not g38762 (n_15403, n23192);
  and g38763 (n23456, n23190, n_15403);
  not g38764 (n_15404, n23456);
  and g38765 (n23457, n_15187, n_15404);
  and g38766 (n23458, n6233, n22377);
  and g38767 (n23459, n5663, n22384);
  and g38768 (n23460, n5939, n22380);
  not g38769 (n_15405, n23459);
  not g38770 (n_15406, n23460);
  and g38771 (n23461, n_15405, n_15406);
  not g38772 (n_15407, n23458);
  and g38773 (n23462, n_15407, n23461);
  and g38774 (n23463, n_1409, n23462);
  and g38775 (n23464, n22834, n23462);
  not g38776 (n_15408, n23463);
  not g38777 (n_15409, n23464);
  and g38778 (n23465, n_15408, n_15409);
  not g38779 (n_15410, n23465);
  and g38780 (n23466, \a[17] , n_15410);
  and g38781 (n23467, n_617, n23465);
  not g38782 (n_15411, n23466);
  not g38783 (n_15412, n23467);
  and g38784 (n23468, n_15411, n_15412);
  not g38785 (n_15413, n23468);
  and g38786 (n23469, n23457, n_15413);
  and g38787 (n23470, n23129, n23188);
  not g38788 (n_15414, n23470);
  and g38789 (n23471, n_15183, n_15414);
  and g38790 (n23472, n6233, n22380);
  and g38791 (n23473, n5663, n22387);
  and g38792 (n23474, n5939, n22384);
  not g38793 (n_15415, n23473);
  not g38794 (n_15416, n23474);
  and g38795 (n23475, n_15415, n_15416);
  not g38796 (n_15417, n23472);
  and g38797 (n23476, n_15417, n23475);
  and g38798 (n23477, n_1409, n23476);
  and g38799 (n23478, n_14894, n23476);
  not g38800 (n_15418, n23477);
  not g38801 (n_15419, n23478);
  and g38802 (n23479, n_15418, n_15419);
  not g38803 (n_15420, n23479);
  and g38804 (n23480, \a[17] , n_15420);
  and g38805 (n23481, n_617, n23479);
  not g38806 (n_15421, n23480);
  not g38807 (n_15422, n23481);
  and g38808 (n23482, n_15421, n_15422);
  not g38809 (n_15423, n23482);
  and g38810 (n23483, n23471, n_15423);
  and g38811 (n23484, n6233, n22384);
  and g38812 (n23485, n5663, n22390);
  and g38813 (n23486, n5939, n22387);
  and g38819 (n23489, n5666, n22806);
  not g38822 (n_15428, n23490);
  and g38823 (n23491, \a[17] , n_15428);
  not g38824 (n_15429, n23491);
  and g38825 (n23492, n_15428, n_15429);
  and g38826 (n23493, \a[17] , n_15429);
  not g38827 (n_15430, n23492);
  not g38828 (n_15431, n23493);
  and g38829 (n23494, n_15430, n_15431);
  not g38830 (n_15432, n23186);
  and g38831 (n23495, n23184, n_15432);
  not g38832 (n_15433, n23495);
  and g38833 (n23496, n_15180, n_15433);
  not g38834 (n_15434, n23494);
  and g38835 (n23497, n_15434, n23496);
  not g38836 (n_15435, n23497);
  and g38837 (n23498, n_15434, n_15435);
  and g38838 (n23499, n23496, n_15435);
  not g38839 (n_15436, n23498);
  not g38840 (n_15437, n23499);
  and g38841 (n23500, n_15436, n_15437);
  and g38842 (n23501, n_15173, n_15175);
  and g38843 (n23502, n_15174, n_15175);
  not g38844 (n_15438, n23501);
  not g38845 (n_15439, n23502);
  and g38846 (n23503, n_15438, n_15439);
  and g38847 (n23504, n6233, n22387);
  and g38848 (n23505, n5663, n22393);
  and g38849 (n23506, n5939, n22390);
  not g38850 (n_15440, n23505);
  not g38851 (n_15441, n23506);
  and g38852 (n23507, n_15440, n_15441);
  not g38853 (n_15442, n23504);
  and g38854 (n23508, n_15442, n23507);
  and g38855 (n23509, n_1409, n23508);
  and g38856 (n23510, n_14920, n23508);
  not g38857 (n_15443, n23509);
  not g38858 (n_15444, n23510);
  and g38859 (n23511, n_15443, n_15444);
  not g38860 (n_15445, n23511);
  and g38861 (n23512, \a[17] , n_15445);
  and g38862 (n23513, n_617, n23511);
  not g38863 (n_15446, n23512);
  not g38864 (n_15447, n23513);
  and g38865 (n23514, n_15446, n_15447);
  not g38866 (n_15448, n23503);
  not g38867 (n_15449, n23514);
  and g38868 (n23515, n_15448, n_15449);
  and g38869 (n23516, n6233, n22390);
  and g38870 (n23517, n5663, n22396);
  and g38871 (n23518, n5939, n22393);
  and g38877 (n23521, n5666, n22649);
  not g38880 (n_15454, n23522);
  and g38881 (n23523, \a[17] , n_15454);
  not g38882 (n_15455, n23523);
  and g38883 (n23524, n_15454, n_15455);
  and g38884 (n23525, \a[17] , n_15455);
  not g38885 (n_15456, n23524);
  not g38886 (n_15457, n23525);
  and g38887 (n23526, n_15456, n_15457);
  not g38888 (n_15458, n23155);
  and g38889 (n23527, n_15458, n23166);
  not g38890 (n_15459, n23167);
  not g38891 (n_15460, n23527);
  and g38892 (n23528, n_15459, n_15460);
  not g38893 (n_15461, n23526);
  and g38894 (n23529, n_15461, n23528);
  not g38895 (n_15462, n23529);
  and g38896 (n23530, n_15461, n_15462);
  and g38897 (n23531, n23528, n_15462);
  not g38898 (n_15463, n23530);
  not g38899 (n_15464, n23531);
  and g38900 (n23532, n_15463, n_15464);
  not g38901 (n_15465, n23154);
  and g38902 (n23533, n23152, n_15465);
  not g38903 (n_15466, n23533);
  and g38904 (n23534, n_15458, n_15466);
  and g38905 (n23535, n6233, n22393);
  and g38906 (n23536, n5663, n22399);
  and g38907 (n23537, n5939, n22396);
  not g38908 (n_15467, n23536);
  not g38909 (n_15468, n23537);
  and g38910 (n23538, n_15467, n_15468);
  not g38911 (n_15469, n23535);
  and g38912 (n23539, n_15469, n23538);
  and g38913 (n23540, n_1409, n23539);
  and g38914 (n23541, n_14773, n23539);
  not g38915 (n_15470, n23540);
  not g38916 (n_15471, n23541);
  and g38917 (n23542, n_15470, n_15471);
  not g38918 (n_15472, n23542);
  and g38919 (n23543, \a[17] , n_15472);
  and g38920 (n23544, n_617, n23542);
  not g38921 (n_15473, n23543);
  not g38922 (n_15474, n23544);
  and g38923 (n23545, n_15473, n_15474);
  not g38924 (n_15475, n23545);
  and g38925 (n23546, n23534, n_15475);
  and g38926 (n23547, n5939, n_14508);
  and g38927 (n23548, n6233, n22402);
  not g38928 (n_15476, n23547);
  not g38929 (n_15477, n23548);
  and g38930 (n23549, n_15476, n_15477);
  and g38931 (n23550, n5666, n_14720);
  not g38932 (n_15478, n23550);
  and g38933 (n23551, n23549, n_15478);
  not g38934 (n_15479, n23551);
  and g38935 (n23552, \a[17] , n_15479);
  not g38936 (n_15480, n23552);
  and g38937 (n23553, \a[17] , n_15480);
  and g38938 (n23554, n_15479, n_15480);
  not g38939 (n_15481, n23553);
  not g38940 (n_15482, n23554);
  and g38941 (n23555, n_15481, n_15482);
  and g38942 (n23556, n_1408, n_14508);
  not g38943 (n_15483, n23556);
  and g38944 (n23557, \a[17] , n_15483);
  not g38945 (n_15484, n23555);
  and g38946 (n23558, n_15484, n23557);
  and g38947 (n23559, n6233, n22399);
  and g38948 (n23560, n5663, n_14508);
  and g38949 (n23561, n5939, n22402);
  not g38950 (n_15485, n23560);
  not g38951 (n_15486, n23561);
  and g38952 (n23562, n_15485, n_15486);
  not g38953 (n_15487, n23559);
  and g38954 (n23563, n_15487, n23562);
  and g38955 (n23564, n_1409, n23563);
  and g38956 (n23565, n22625, n23563);
  not g38957 (n_15488, n23564);
  not g38958 (n_15489, n23565);
  and g38959 (n23566, n_15488, n_15489);
  not g38960 (n_15490, n23566);
  and g38961 (n23567, \a[17] , n_15490);
  and g38962 (n23568, n_617, n23566);
  not g38963 (n_15491, n23567);
  not g38964 (n_15492, n23568);
  and g38965 (n23569, n_15491, n_15492);
  not g38966 (n_15493, n23569);
  and g38967 (n23570, n23558, n_15493);
  and g38968 (n23571, n23153, n23570);
  not g38969 (n_15494, n23571);
  and g38970 (n23572, n23570, n_15494);
  and g38971 (n23573, n23153, n_15494);
  not g38972 (n_15495, n23572);
  not g38973 (n_15496, n23573);
  and g38974 (n23574, n_15495, n_15496);
  and g38975 (n23575, n6233, n22396);
  and g38976 (n23576, n5663, n22402);
  and g38977 (n23577, n5939, n22399);
  and g38983 (n23580, n5666, n22595);
  not g38986 (n_15501, n23581);
  and g38987 (n23582, \a[17] , n_15501);
  not g38988 (n_15502, n23582);
  and g38989 (n23583, \a[17] , n_15502);
  and g38990 (n23584, n_15501, n_15502);
  not g38991 (n_15503, n23583);
  not g38992 (n_15504, n23584);
  and g38993 (n23585, n_15503, n_15504);
  not g38994 (n_15505, n23574);
  not g38995 (n_15506, n23585);
  and g38996 (n23586, n_15505, n_15506);
  not g38997 (n_15507, n23586);
  and g38998 (n23587, n_15494, n_15507);
  not g38999 (n_15508, n23534);
  and g39000 (n23588, n_15508, n23545);
  not g39001 (n_15509, n23546);
  not g39002 (n_15510, n23588);
  and g39003 (n23589, n_15509, n_15510);
  not g39004 (n_15511, n23587);
  and g39005 (n23590, n_15511, n23589);
  not g39006 (n_15512, n23590);
  and g39007 (n23591, n_15509, n_15512);
  not g39008 (n_15513, n23532);
  not g39009 (n_15514, n23591);
  and g39010 (n23592, n_15513, n_15514);
  not g39011 (n_15515, n23592);
  and g39012 (n23593, n_15462, n_15515);
  and g39013 (n23594, n23503, n23514);
  not g39014 (n_15516, n23515);
  not g39015 (n_15517, n23594);
  and g39016 (n23595, n_15516, n_15517);
  not g39017 (n_15518, n23593);
  and g39018 (n23596, n_15518, n23595);
  not g39019 (n_15519, n23596);
  and g39020 (n23597, n_15516, n_15519);
  not g39021 (n_15520, n23500);
  not g39022 (n_15521, n23597);
  and g39023 (n23598, n_15520, n_15521);
  not g39024 (n_15522, n23598);
  and g39025 (n23599, n_15435, n_15522);
  not g39026 (n_15523, n23483);
  and g39027 (n23600, n23471, n_15523);
  and g39028 (n23601, n_15423, n_15523);
  not g39029 (n_15524, n23600);
  not g39030 (n_15525, n23601);
  and g39031 (n23602, n_15524, n_15525);
  not g39032 (n_15526, n23599);
  not g39033 (n_15527, n23602);
  and g39034 (n23603, n_15526, n_15527);
  not g39035 (n_15528, n23603);
  and g39036 (n23604, n_15523, n_15528);
  not g39037 (n_15529, n23469);
  and g39038 (n23605, n23457, n_15529);
  and g39039 (n23606, n_15413, n_15529);
  not g39040 (n_15530, n23605);
  not g39041 (n_15531, n23606);
  and g39042 (n23607, n_15530, n_15531);
  not g39043 (n_15532, n23604);
  not g39044 (n_15533, n23607);
  and g39045 (n23608, n_15532, n_15533);
  not g39046 (n_15534, n23608);
  and g39047 (n23609, n_15529, n_15534);
  not g39048 (n_15535, n23443);
  and g39049 (n23610, n_15535, n23454);
  not g39050 (n_15536, n23455);
  not g39051 (n_15537, n23610);
  and g39052 (n23611, n_15536, n_15537);
  not g39053 (n_15538, n23609);
  and g39054 (n23612, n_15538, n23611);
  not g39055 (n_15539, n23612);
  and g39056 (n23613, n_15536, n_15539);
  not g39057 (n_15540, n23441);
  not g39058 (n_15541, n23613);
  and g39059 (n23614, n_15540, n_15541);
  not g39060 (n_15542, n23614);
  and g39061 (n23615, n_15390, n_15542);
  not g39062 (n_15543, n23423);
  not g39063 (n_15544, n23615);
  and g39064 (n23616, n_15543, n_15544);
  not g39065 (n_15545, n23616);
  and g39066 (n23617, n_15375, n_15545);
  not g39067 (n_15546, n23405);
  not g39068 (n_15547, n23617);
  and g39069 (n23618, n_15546, n_15547);
  not g39070 (n_15548, n23618);
  and g39071 (n23619, n_15360, n_15548);
  not g39072 (n_15549, n23388);
  and g39073 (n23620, n23376, n_15549);
  and g39074 (n23621, n_15347, n_15549);
  not g39075 (n_15550, n23620);
  not g39076 (n_15551, n23621);
  and g39077 (n23622, n_15550, n_15551);
  not g39078 (n_15552, n23619);
  not g39079 (n_15553, n23622);
  and g39080 (n23623, n_15552, n_15553);
  not g39081 (n_15554, n23623);
  and g39082 (n23624, n_15549, n_15554);
  not g39083 (n_15555, n23360);
  and g39084 (n23625, n_15555, n23373);
  not g39085 (n_15556, n23374);
  not g39086 (n_15557, n23625);
  and g39087 (n23626, n_15556, n_15557);
  not g39088 (n_15558, n23624);
  and g39089 (n23627, n_15558, n23626);
  not g39090 (n_15559, n23627);
  and g39091 (n23628, n_15556, n_15559);
  not g39092 (n_15560, n23358);
  not g39093 (n_15561, n23628);
  and g39094 (n23629, n_15560, n_15561);
  not g39095 (n_15562, n23629);
  and g39096 (n23630, n_15322, n_15562);
  and g39097 (n23631, n23337, n23630);
  not g39098 (n_15563, n23337);
  not g39099 (n_15564, n23630);
  and g39100 (n23632, n_15563, n_15564);
  not g39101 (n_15565, n23631);
  not g39102 (n_15566, n23632);
  and g39103 (n23633, n_15565, n_15566);
  and g39104 (n23634, n7101, n22344);
  and g39105 (n23635, n6402, n22350);
  and g39106 (n23636, n6951, n22347);
  not g39107 (n_15567, n23635);
  not g39108 (n_15568, n23636);
  and g39109 (n23637, n_15567, n_15568);
  not g39110 (n_15569, n23634);
  and g39111 (n23638, n_15569, n23637);
  and g39112 (n23639, n_1885, n23638);
  and g39113 (n23640, n_14596, n_14599);
  and g39114 (n23641, n_14597, n22480);
  not g39115 (n_15570, n23640);
  not g39116 (n_15571, n23641);
  and g39117 (n23642, n_15570, n_15571);
  and g39118 (n23643, n23638, n23642);
  not g39119 (n_15572, n23639);
  not g39120 (n_15573, n23643);
  and g39121 (n23644, n_15572, n_15573);
  not g39122 (n_15574, n23644);
  and g39123 (n23645, \a[14] , n_15574);
  and g39124 (n23646, n_652, n23644);
  not g39125 (n_15575, n23645);
  not g39126 (n_15576, n23646);
  and g39127 (n23647, n_15575, n_15576);
  not g39128 (n_15577, n23647);
  and g39129 (n23648, n23633, n_15577);
  and g39130 (n23649, n23358, n23628);
  not g39131 (n_15578, n23649);
  and g39132 (n23650, n_15562, n_15578);
  and g39133 (n23651, n7101, n22347);
  and g39134 (n23652, n6402, n22353);
  and g39135 (n23653, n6951, n22350);
  not g39136 (n_15579, n23652);
  not g39137 (n_15580, n23653);
  and g39138 (n23654, n_15579, n_15580);
  not g39139 (n_15581, n23651);
  and g39140 (n23655, n_15581, n23654);
  and g39141 (n23656, n_1885, n23655);
  and g39142 (n23657, n_14591, n_14594);
  and g39143 (n23658, n_14592, n22476);
  not g39144 (n_15582, n23657);
  not g39145 (n_15583, n23658);
  and g39146 (n23659, n_15582, n_15583);
  and g39147 (n23660, n23655, n23659);
  not g39148 (n_15584, n23656);
  not g39149 (n_15585, n23660);
  and g39150 (n23661, n_15584, n_15585);
  not g39151 (n_15586, n23661);
  and g39152 (n23662, \a[14] , n_15586);
  and g39153 (n23663, n_652, n23661);
  not g39154 (n_15587, n23662);
  not g39155 (n_15588, n23663);
  and g39156 (n23664, n_15587, n_15588);
  not g39157 (n_15589, n23664);
  and g39158 (n23665, n23650, n_15589);
  and g39159 (n23666, n7101, n22350);
  and g39160 (n23667, n6402, n22356);
  and g39161 (n23668, n6951, n22353);
  not g39167 (n_15593, n22470);
  and g39168 (n23671, n22468, n_15593);
  not g39169 (n_15594, n23671);
  and g39170 (n23672, n_14589, n_15594);
  and g39171 (n23673, n6397, n23672);
  not g39174 (n_15596, n23674);
  and g39175 (n23675, \a[14] , n_15596);
  not g39176 (n_15597, n23675);
  and g39177 (n23676, n_15596, n_15597);
  and g39178 (n23677, \a[14] , n_15597);
  not g39179 (n_15598, n23676);
  not g39180 (n_15599, n23677);
  and g39181 (n23678, n_15598, n_15599);
  not g39182 (n_15600, n23626);
  and g39183 (n23679, n23624, n_15600);
  not g39184 (n_15601, n23679);
  and g39185 (n23680, n_15559, n_15601);
  not g39186 (n_15602, n23678);
  and g39187 (n23681, n_15602, n23680);
  not g39188 (n_15603, n23681);
  and g39189 (n23682, n_15602, n_15603);
  and g39190 (n23683, n23680, n_15603);
  not g39191 (n_15604, n23682);
  not g39192 (n_15605, n23683);
  and g39193 (n23684, n_15604, n_15605);
  and g39194 (n23685, n7101, n22353);
  and g39195 (n23686, n6402, n22359);
  and g39196 (n23687, n6951, n22356);
  and g39202 (n23690, n6397, n_14678);
  not g39205 (n_15610, n23691);
  and g39206 (n23692, \a[14] , n_15610);
  not g39207 (n_15611, n23692);
  and g39208 (n23693, n_15610, n_15611);
  and g39209 (n23694, \a[14] , n_15611);
  not g39210 (n_15612, n23693);
  not g39211 (n_15613, n23694);
  and g39212 (n23695, n_15612, n_15613);
  and g39213 (n23696, n_15552, n_15554);
  and g39214 (n23697, n_15553, n_15554);
  not g39215 (n_15614, n23696);
  not g39216 (n_15615, n23697);
  and g39217 (n23698, n_15614, n_15615);
  not g39218 (n_15616, n23695);
  not g39219 (n_15617, n23698);
  and g39220 (n23699, n_15616, n_15617);
  not g39221 (n_15618, n23699);
  and g39222 (n23700, n_15616, n_15618);
  and g39223 (n23701, n_15617, n_15618);
  not g39224 (n_15619, n23700);
  not g39225 (n_15620, n23701);
  and g39226 (n23702, n_15619, n_15620);
  and g39227 (n23703, n23405, n23617);
  not g39228 (n_15621, n23703);
  and g39229 (n23704, n_15548, n_15621);
  and g39230 (n23705, n7101, n22356);
  and g39231 (n23706, n6402, n22362);
  and g39232 (n23707, n6951, n22359);
  not g39233 (n_15622, n23706);
  not g39234 (n_15623, n23707);
  and g39235 (n23708, n_15622, n_15623);
  not g39236 (n_15624, n23705);
  and g39237 (n23709, n_15624, n23708);
  and g39238 (n23710, n_1885, n23709);
  and g39239 (n23711, n23345, n23709);
  not g39240 (n_15625, n23710);
  not g39241 (n_15626, n23711);
  and g39242 (n23712, n_15625, n_15626);
  not g39243 (n_15627, n23712);
  and g39244 (n23713, \a[14] , n_15627);
  and g39245 (n23714, n_652, n23712);
  not g39246 (n_15628, n23713);
  not g39247 (n_15629, n23714);
  and g39248 (n23715, n_15628, n_15629);
  not g39249 (n_15630, n23715);
  and g39250 (n23716, n23704, n_15630);
  and g39251 (n23717, n23423, n23615);
  not g39252 (n_15631, n23717);
  and g39253 (n23718, n_15545, n_15631);
  and g39254 (n23719, n7101, n22359);
  and g39255 (n23720, n6402, n22365);
  and g39256 (n23721, n6951, n22362);
  not g39257 (n_15632, n23720);
  not g39258 (n_15633, n23721);
  and g39259 (n23722, n_15632, n_15633);
  not g39260 (n_15634, n23719);
  and g39261 (n23723, n_15634, n23722);
  and g39262 (n23724, n_1885, n23723);
  and g39263 (n23725, n_15331, n23723);
  not g39264 (n_15635, n23724);
  not g39265 (n_15636, n23725);
  and g39266 (n23726, n_15635, n_15636);
  not g39267 (n_15637, n23726);
  and g39268 (n23727, \a[14] , n_15637);
  and g39269 (n23728, n_652, n23726);
  not g39270 (n_15638, n23727);
  not g39271 (n_15639, n23728);
  and g39272 (n23729, n_15638, n_15639);
  not g39273 (n_15640, n23729);
  and g39274 (n23730, n23718, n_15640);
  and g39275 (n23731, n23441, n23613);
  not g39276 (n_15641, n23731);
  and g39277 (n23732, n_15542, n_15641);
  and g39278 (n23733, n7101, n22362);
  and g39279 (n23734, n6402, n22368);
  and g39280 (n23735, n6951, n22365);
  not g39281 (n_15642, n23734);
  not g39282 (n_15643, n23735);
  and g39283 (n23736, n_15642, n_15643);
  not g39284 (n_15644, n23733);
  and g39285 (n23737, n_15644, n23736);
  and g39286 (n23738, n_1885, n23737);
  and g39287 (n23739, n23320, n23737);
  not g39288 (n_15645, n23738);
  not g39289 (n_15646, n23739);
  and g39290 (n23740, n_15645, n_15646);
  not g39291 (n_15647, n23740);
  and g39292 (n23741, \a[14] , n_15647);
  and g39293 (n23742, n_652, n23740);
  not g39294 (n_15648, n23741);
  not g39295 (n_15649, n23742);
  and g39296 (n23743, n_15648, n_15649);
  not g39297 (n_15650, n23743);
  and g39298 (n23744, n23732, n_15650);
  and g39299 (n23745, n7101, n22365);
  and g39300 (n23746, n6402, n22371);
  and g39301 (n23747, n6951, n22368);
  and g39307 (n23750, n6397, n_15351);
  not g39310 (n_15655, n23751);
  and g39311 (n23752, \a[14] , n_15655);
  not g39312 (n_15656, n23752);
  and g39313 (n23753, n_15655, n_15656);
  and g39314 (n23754, \a[14] , n_15656);
  not g39315 (n_15657, n23753);
  not g39316 (n_15658, n23754);
  and g39317 (n23755, n_15657, n_15658);
  not g39318 (n_15659, n23611);
  and g39319 (n23756, n23609, n_15659);
  not g39320 (n_15660, n23756);
  and g39321 (n23757, n_15539, n_15660);
  not g39322 (n_15661, n23755);
  and g39323 (n23758, n_15661, n23757);
  not g39324 (n_15662, n23758);
  and g39325 (n23759, n_15661, n_15662);
  and g39326 (n23760, n23757, n_15662);
  not g39327 (n_15663, n23759);
  not g39328 (n_15664, n23760);
  and g39329 (n23761, n_15663, n_15664);
  and g39330 (n23762, n7101, n22368);
  and g39331 (n23763, n6402, n22374);
  and g39332 (n23764, n6951, n22371);
  and g39338 (n23767, n6397, n23006);
  not g39341 (n_15669, n23768);
  and g39342 (n23769, \a[14] , n_15669);
  not g39343 (n_15670, n23769);
  and g39344 (n23770, n_15669, n_15670);
  and g39345 (n23771, \a[14] , n_15670);
  not g39346 (n_15671, n23770);
  not g39347 (n_15672, n23771);
  and g39348 (n23772, n_15671, n_15672);
  and g39349 (n23773, n_15532, n_15534);
  and g39350 (n23774, n_15533, n_15534);
  not g39351 (n_15673, n23773);
  not g39352 (n_15674, n23774);
  and g39353 (n23775, n_15673, n_15674);
  not g39354 (n_15675, n23772);
  not g39355 (n_15676, n23775);
  and g39356 (n23776, n_15675, n_15676);
  not g39357 (n_15677, n23776);
  and g39358 (n23777, n_15675, n_15677);
  and g39359 (n23778, n_15676, n_15677);
  not g39360 (n_15678, n23777);
  not g39361 (n_15679, n23778);
  and g39362 (n23779, n_15678, n_15679);
  and g39363 (n23780, n7101, n22371);
  and g39364 (n23781, n6402, n22377);
  and g39365 (n23782, n6951, n22374);
  and g39371 (n23785, n6397, n23025);
  not g39374 (n_15684, n23786);
  and g39375 (n23787, \a[14] , n_15684);
  not g39376 (n_15685, n23787);
  and g39377 (n23788, n_15684, n_15685);
  and g39378 (n23789, \a[14] , n_15685);
  not g39379 (n_15686, n23788);
  not g39380 (n_15687, n23789);
  and g39381 (n23790, n_15686, n_15687);
  and g39382 (n23791, n_15526, n_15528);
  and g39383 (n23792, n_15527, n_15528);
  not g39384 (n_15688, n23791);
  not g39385 (n_15689, n23792);
  and g39386 (n23793, n_15688, n_15689);
  not g39387 (n_15690, n23790);
  not g39388 (n_15691, n23793);
  and g39389 (n23794, n_15690, n_15691);
  not g39390 (n_15692, n23794);
  and g39391 (n23795, n_15690, n_15692);
  and g39392 (n23796, n_15691, n_15692);
  not g39393 (n_15693, n23795);
  not g39394 (n_15694, n23796);
  and g39395 (n23797, n_15693, n_15694);
  and g39396 (n23798, n23500, n23597);
  not g39397 (n_15695, n23798);
  and g39398 (n23799, n_15522, n_15695);
  and g39399 (n23800, n7101, n22374);
  and g39400 (n23801, n6402, n22380);
  and g39401 (n23802, n6951, n22377);
  not g39402 (n_15696, n23801);
  not g39403 (n_15697, n23802);
  and g39404 (n23803, n_15696, n_15697);
  not g39405 (n_15698, n23800);
  and g39406 (n23804, n_15698, n23803);
  and g39407 (n23805, n_1885, n23804);
  and g39408 (n23806, n_15064, n23804);
  not g39409 (n_15699, n23805);
  not g39410 (n_15700, n23806);
  and g39411 (n23807, n_15699, n_15700);
  not g39412 (n_15701, n23807);
  and g39413 (n23808, \a[14] , n_15701);
  and g39414 (n23809, n_652, n23807);
  not g39415 (n_15702, n23808);
  not g39416 (n_15703, n23809);
  and g39417 (n23810, n_15702, n_15703);
  not g39418 (n_15704, n23810);
  and g39419 (n23811, n23799, n_15704);
  not g39420 (n_15705, n23595);
  and g39421 (n23812, n23593, n_15705);
  not g39422 (n_15706, n23812);
  and g39423 (n23813, n_15519, n_15706);
  and g39424 (n23814, n7101, n22377);
  and g39425 (n23815, n6402, n22384);
  and g39426 (n23816, n6951, n22380);
  not g39427 (n_15707, n23815);
  not g39428 (n_15708, n23816);
  and g39429 (n23817, n_15707, n_15708);
  not g39430 (n_15709, n23814);
  and g39431 (n23818, n_15709, n23817);
  and g39432 (n23819, n_1885, n23818);
  and g39433 (n23820, n22834, n23818);
  not g39434 (n_15710, n23819);
  not g39435 (n_15711, n23820);
  and g39436 (n23821, n_15710, n_15711);
  not g39437 (n_15712, n23821);
  and g39438 (n23822, \a[14] , n_15712);
  and g39439 (n23823, n_652, n23821);
  not g39440 (n_15713, n23822);
  not g39441 (n_15714, n23823);
  and g39442 (n23824, n_15713, n_15714);
  not g39443 (n_15715, n23824);
  and g39444 (n23825, n23813, n_15715);
  and g39445 (n23826, n23532, n23591);
  not g39446 (n_15716, n23826);
  and g39447 (n23827, n_15515, n_15716);
  and g39448 (n23828, n7101, n22380);
  and g39449 (n23829, n6402, n22387);
  and g39450 (n23830, n6951, n22384);
  not g39451 (n_15717, n23829);
  not g39452 (n_15718, n23830);
  and g39453 (n23831, n_15717, n_15718);
  not g39454 (n_15719, n23828);
  and g39455 (n23832, n_15719, n23831);
  and g39456 (n23833, n_1885, n23832);
  and g39457 (n23834, n_14894, n23832);
  not g39458 (n_15720, n23833);
  not g39459 (n_15721, n23834);
  and g39460 (n23835, n_15720, n_15721);
  not g39461 (n_15722, n23835);
  and g39462 (n23836, \a[14] , n_15722);
  and g39463 (n23837, n_652, n23835);
  not g39464 (n_15723, n23836);
  not g39465 (n_15724, n23837);
  and g39466 (n23838, n_15723, n_15724);
  not g39467 (n_15725, n23838);
  and g39468 (n23839, n23827, n_15725);
  and g39469 (n23840, n7101, n22384);
  and g39470 (n23841, n6402, n22390);
  and g39471 (n23842, n6951, n22387);
  and g39477 (n23845, n6397, n22806);
  not g39480 (n_15730, n23846);
  and g39481 (n23847, \a[14] , n_15730);
  not g39482 (n_15731, n23847);
  and g39483 (n23848, n_15730, n_15731);
  and g39484 (n23849, \a[14] , n_15731);
  not g39485 (n_15732, n23848);
  not g39486 (n_15733, n23849);
  and g39487 (n23850, n_15732, n_15733);
  not g39488 (n_15734, n23589);
  and g39489 (n23851, n23587, n_15734);
  not g39490 (n_15735, n23851);
  and g39491 (n23852, n_15512, n_15735);
  not g39492 (n_15736, n23850);
  and g39493 (n23853, n_15736, n23852);
  not g39494 (n_15737, n23853);
  and g39495 (n23854, n_15736, n_15737);
  and g39496 (n23855, n23852, n_15737);
  not g39497 (n_15738, n23854);
  not g39498 (n_15739, n23855);
  and g39499 (n23856, n_15738, n_15739);
  and g39500 (n23857, n_15505, n_15507);
  and g39501 (n23858, n_15506, n_15507);
  not g39502 (n_15740, n23857);
  not g39503 (n_15741, n23858);
  and g39504 (n23859, n_15740, n_15741);
  and g39505 (n23860, n7101, n22387);
  and g39506 (n23861, n6402, n22393);
  and g39507 (n23862, n6951, n22390);
  not g39508 (n_15742, n23861);
  not g39509 (n_15743, n23862);
  and g39510 (n23863, n_15742, n_15743);
  not g39511 (n_15744, n23860);
  and g39512 (n23864, n_15744, n23863);
  and g39513 (n23865, n_1885, n23864);
  and g39514 (n23866, n_14920, n23864);
  not g39515 (n_15745, n23865);
  not g39516 (n_15746, n23866);
  and g39517 (n23867, n_15745, n_15746);
  not g39518 (n_15747, n23867);
  and g39519 (n23868, \a[14] , n_15747);
  and g39520 (n23869, n_652, n23867);
  not g39521 (n_15748, n23868);
  not g39522 (n_15749, n23869);
  and g39523 (n23870, n_15748, n_15749);
  not g39524 (n_15750, n23859);
  not g39525 (n_15751, n23870);
  and g39526 (n23871, n_15750, n_15751);
  and g39527 (n23872, n7101, n22390);
  and g39528 (n23873, n6402, n22396);
  and g39529 (n23874, n6951, n22393);
  and g39535 (n23877, n6397, n22649);
  not g39538 (n_15756, n23878);
  and g39539 (n23879, \a[14] , n_15756);
  not g39540 (n_15757, n23879);
  and g39541 (n23880, n_15756, n_15757);
  and g39542 (n23881, \a[14] , n_15757);
  not g39543 (n_15758, n23880);
  not g39544 (n_15759, n23881);
  and g39545 (n23882, n_15758, n_15759);
  not g39546 (n_15760, n23558);
  and g39547 (n23883, n_15760, n23569);
  not g39548 (n_15761, n23570);
  not g39549 (n_15762, n23883);
  and g39550 (n23884, n_15761, n_15762);
  not g39551 (n_15763, n23882);
  and g39552 (n23885, n_15763, n23884);
  not g39553 (n_15764, n23885);
  and g39554 (n23886, n_15763, n_15764);
  and g39555 (n23887, n23884, n_15764);
  not g39556 (n_15765, n23886);
  not g39557 (n_15766, n23887);
  and g39558 (n23888, n_15765, n_15766);
  not g39559 (n_15767, n23557);
  and g39560 (n23889, n23555, n_15767);
  not g39561 (n_15768, n23889);
  and g39562 (n23890, n_15760, n_15768);
  and g39563 (n23891, n7101, n22393);
  and g39564 (n23892, n6402, n22399);
  and g39565 (n23893, n6951, n22396);
  not g39566 (n_15769, n23892);
  not g39567 (n_15770, n23893);
  and g39568 (n23894, n_15769, n_15770);
  not g39569 (n_15771, n23891);
  and g39570 (n23895, n_15771, n23894);
  and g39571 (n23896, n_1885, n23895);
  and g39572 (n23897, n_14773, n23895);
  not g39573 (n_15772, n23896);
  not g39574 (n_15773, n23897);
  and g39575 (n23898, n_15772, n_15773);
  not g39576 (n_15774, n23898);
  and g39577 (n23899, \a[14] , n_15774);
  and g39578 (n23900, n_652, n23898);
  not g39579 (n_15775, n23899);
  not g39580 (n_15776, n23900);
  and g39581 (n23901, n_15775, n_15776);
  not g39582 (n_15777, n23901);
  and g39583 (n23902, n23890, n_15777);
  and g39584 (n23903, n6951, n_14508);
  and g39585 (n23904, n7101, n22402);
  not g39586 (n_15778, n23903);
  not g39587 (n_15779, n23904);
  and g39588 (n23905, n_15778, n_15779);
  and g39589 (n23906, n6397, n_14720);
  not g39590 (n_15780, n23906);
  and g39591 (n23907, n23905, n_15780);
  not g39592 (n_15781, n23907);
  and g39593 (n23908, \a[14] , n_15781);
  not g39594 (n_15782, n23908);
  and g39595 (n23909, \a[14] , n_15782);
  and g39596 (n23910, n_15781, n_15782);
  not g39597 (n_15783, n23909);
  not g39598 (n_15784, n23910);
  and g39599 (n23911, n_15783, n_15784);
  and g39600 (n23912, n_1881, n_14508);
  not g39601 (n_15785, n23912);
  and g39602 (n23913, \a[14] , n_15785);
  not g39603 (n_15786, n23911);
  and g39604 (n23914, n_15786, n23913);
  and g39605 (n23915, n7101, n22399);
  and g39606 (n23916, n6402, n_14508);
  and g39607 (n23917, n6951, n22402);
  not g39608 (n_15787, n23916);
  not g39609 (n_15788, n23917);
  and g39610 (n23918, n_15787, n_15788);
  not g39611 (n_15789, n23915);
  and g39612 (n23919, n_15789, n23918);
  and g39613 (n23920, n_1885, n23919);
  and g39614 (n23921, n22625, n23919);
  not g39615 (n_15790, n23920);
  not g39616 (n_15791, n23921);
  and g39617 (n23922, n_15790, n_15791);
  not g39618 (n_15792, n23922);
  and g39619 (n23923, \a[14] , n_15792);
  and g39620 (n23924, n_652, n23922);
  not g39621 (n_15793, n23923);
  not g39622 (n_15794, n23924);
  and g39623 (n23925, n_15793, n_15794);
  not g39624 (n_15795, n23925);
  and g39625 (n23926, n23914, n_15795);
  and g39626 (n23927, n23556, n23926);
  not g39627 (n_15796, n23927);
  and g39628 (n23928, n23926, n_15796);
  and g39629 (n23929, n23556, n_15796);
  not g39630 (n_15797, n23928);
  not g39631 (n_15798, n23929);
  and g39632 (n23930, n_15797, n_15798);
  and g39633 (n23931, n7101, n22396);
  and g39634 (n23932, n6402, n22402);
  and g39635 (n23933, n6951, n22399);
  and g39641 (n23936, n6397, n22595);
  not g39644 (n_15803, n23937);
  and g39645 (n23938, \a[14] , n_15803);
  not g39646 (n_15804, n23938);
  and g39647 (n23939, \a[14] , n_15804);
  and g39648 (n23940, n_15803, n_15804);
  not g39649 (n_15805, n23939);
  not g39650 (n_15806, n23940);
  and g39651 (n23941, n_15805, n_15806);
  not g39652 (n_15807, n23930);
  not g39653 (n_15808, n23941);
  and g39654 (n23942, n_15807, n_15808);
  not g39655 (n_15809, n23942);
  and g39656 (n23943, n_15796, n_15809);
  not g39657 (n_15810, n23890);
  and g39658 (n23944, n_15810, n23901);
  not g39659 (n_15811, n23902);
  not g39660 (n_15812, n23944);
  and g39661 (n23945, n_15811, n_15812);
  not g39662 (n_15813, n23943);
  and g39663 (n23946, n_15813, n23945);
  not g39664 (n_15814, n23946);
  and g39665 (n23947, n_15811, n_15814);
  not g39666 (n_15815, n23888);
  not g39667 (n_15816, n23947);
  and g39668 (n23948, n_15815, n_15816);
  not g39669 (n_15817, n23948);
  and g39670 (n23949, n_15764, n_15817);
  and g39671 (n23950, n23859, n23870);
  not g39672 (n_15818, n23871);
  not g39673 (n_15819, n23950);
  and g39674 (n23951, n_15818, n_15819);
  not g39675 (n_15820, n23949);
  and g39676 (n23952, n_15820, n23951);
  not g39677 (n_15821, n23952);
  and g39678 (n23953, n_15818, n_15821);
  not g39679 (n_15822, n23856);
  not g39680 (n_15823, n23953);
  and g39681 (n23954, n_15822, n_15823);
  not g39682 (n_15824, n23954);
  and g39683 (n23955, n_15737, n_15824);
  not g39684 (n_15825, n23839);
  and g39685 (n23956, n23827, n_15825);
  and g39686 (n23957, n_15725, n_15825);
  not g39687 (n_15826, n23956);
  not g39688 (n_15827, n23957);
  and g39689 (n23958, n_15826, n_15827);
  not g39690 (n_15828, n23955);
  not g39691 (n_15829, n23958);
  and g39692 (n23959, n_15828, n_15829);
  not g39693 (n_15830, n23959);
  and g39694 (n23960, n_15825, n_15830);
  not g39695 (n_15831, n23825);
  and g39696 (n23961, n23813, n_15831);
  and g39697 (n23962, n_15715, n_15831);
  not g39698 (n_15832, n23961);
  not g39699 (n_15833, n23962);
  and g39700 (n23963, n_15832, n_15833);
  not g39701 (n_15834, n23960);
  not g39702 (n_15835, n23963);
  and g39703 (n23964, n_15834, n_15835);
  not g39704 (n_15836, n23964);
  and g39705 (n23965, n_15831, n_15836);
  not g39706 (n_15837, n23799);
  and g39707 (n23966, n_15837, n23810);
  not g39708 (n_15838, n23811);
  not g39709 (n_15839, n23966);
  and g39710 (n23967, n_15838, n_15839);
  not g39711 (n_15840, n23965);
  and g39712 (n23968, n_15840, n23967);
  not g39713 (n_15841, n23968);
  and g39714 (n23969, n_15838, n_15841);
  not g39715 (n_15842, n23797);
  not g39716 (n_15843, n23969);
  and g39717 (n23970, n_15842, n_15843);
  not g39718 (n_15844, n23970);
  and g39719 (n23971, n_15692, n_15844);
  not g39720 (n_15845, n23779);
  not g39721 (n_15846, n23971);
  and g39722 (n23972, n_15845, n_15846);
  not g39723 (n_15847, n23972);
  and g39724 (n23973, n_15677, n_15847);
  not g39725 (n_15848, n23761);
  not g39726 (n_15849, n23973);
  and g39727 (n23974, n_15848, n_15849);
  not g39728 (n_15850, n23974);
  and g39729 (n23975, n_15662, n_15850);
  not g39730 (n_15851, n23744);
  and g39731 (n23976, n23732, n_15851);
  and g39732 (n23977, n_15650, n_15851);
  not g39733 (n_15852, n23976);
  not g39734 (n_15853, n23977);
  and g39735 (n23978, n_15852, n_15853);
  not g39736 (n_15854, n23975);
  not g39737 (n_15855, n23978);
  and g39738 (n23979, n_15854, n_15855);
  not g39739 (n_15856, n23979);
  and g39740 (n23980, n_15851, n_15856);
  not g39741 (n_15857, n23730);
  and g39742 (n23981, n23718, n_15857);
  and g39743 (n23982, n_15640, n_15857);
  not g39744 (n_15858, n23981);
  not g39745 (n_15859, n23982);
  and g39746 (n23983, n_15858, n_15859);
  not g39747 (n_15860, n23980);
  not g39748 (n_15861, n23983);
  and g39749 (n23984, n_15860, n_15861);
  not g39750 (n_15862, n23984);
  and g39751 (n23985, n_15857, n_15862);
  not g39752 (n_15863, n23704);
  and g39753 (n23986, n_15863, n23715);
  not g39754 (n_15864, n23716);
  not g39755 (n_15865, n23986);
  and g39756 (n23987, n_15864, n_15865);
  not g39757 (n_15866, n23985);
  and g39758 (n23988, n_15866, n23987);
  not g39759 (n_15867, n23988);
  and g39760 (n23989, n_15864, n_15867);
  not g39761 (n_15868, n23702);
  not g39762 (n_15869, n23989);
  and g39763 (n23990, n_15868, n_15869);
  not g39764 (n_15870, n23990);
  and g39765 (n23991, n_15618, n_15870);
  not g39766 (n_15871, n23684);
  not g39767 (n_15872, n23991);
  and g39768 (n23992, n_15871, n_15872);
  not g39769 (n_15873, n23992);
  and g39770 (n23993, n_15603, n_15873);
  not g39771 (n_15874, n23665);
  and g39772 (n23994, n23650, n_15874);
  and g39773 (n23995, n_15589, n_15874);
  not g39774 (n_15875, n23994);
  not g39775 (n_15876, n23995);
  and g39776 (n23996, n_15875, n_15876);
  not g39777 (n_15877, n23993);
  not g39778 (n_15878, n23996);
  and g39779 (n23997, n_15877, n_15878);
  not g39780 (n_15879, n23997);
  and g39781 (n23998, n_15874, n_15879);
  not g39782 (n_15880, n23648);
  and g39783 (n23999, n23633, n_15880);
  and g39784 (n24000, n_15577, n_15880);
  not g39785 (n_15881, n23999);
  not g39786 (n_15882, n24000);
  and g39787 (n24001, n_15881, n_15882);
  not g39788 (n_15883, n23998);
  not g39789 (n_15884, n24001);
  and g39790 (n24002, n_15883, n_15884);
  not g39791 (n_15885, n24002);
  and g39792 (n24003, n_15880, n_15885);
  and g39793 (n24004, n6233, n22350);
  and g39794 (n24005, n5663, n22356);
  and g39795 (n24006, n5939, n22353);
  and g39801 (n24009, n5666, n23672);
  not g39804 (n_15890, n24010);
  and g39805 (n24011, \a[17] , n_15890);
  not g39806 (n_15891, n24011);
  and g39807 (n24012, n_15890, n_15891);
  and g39808 (n24013, \a[17] , n_15891);
  not g39809 (n_15892, n24012);
  not g39810 (n_15893, n24013);
  and g39811 (n24014, n_15892, n_15893);
  and g39812 (n24015, n_15294, n_15299);
  and g39813 (n24016, n4694, n22368);
  and g39814 (n24017, n4533, n22374);
  and g39815 (n24018, n4604, n22371);
  and g39821 (n24021, n4536, n23006);
  not g39824 (n_15898, n24022);
  and g39825 (n24023, \a[23] , n_15898);
  not g39826 (n_15899, n24023);
  and g39827 (n24024, n_15898, n_15899);
  and g39828 (n24025, \a[23] , n_15899);
  not g39829 (n_15900, n24024);
  not g39830 (n_15901, n24025);
  and g39831 (n24026, n_15900, n_15901);
  and g39832 (n24027, n_15266, n_15271);
  and g39833 (n24028, n3457, n22387);
  and g39834 (n24029, n3542, n22393);
  and g39835 (n24030, n3606, n22390);
  and g39841 (n24033, n3368, n22582);
  not g39844 (n_15906, n24034);
  and g39845 (n24035, \a[29] , n_15906);
  not g39846 (n_15907, n24035);
  and g39847 (n24036, n_15906, n_15907);
  and g39848 (n24037, \a[29] , n_15907);
  not g39849 (n_15908, n24036);
  not g39850 (n_15909, n24037);
  and g39851 (n24038, n_15908, n_15909);
  and g39852 (n24039, n_15242, n_15245);
  and g39853 (n24040, n116, n_212);
  and g39854 (n24041, n_215, n24040);
  and g39871 (n24058, n3020, n22396);
  and g39872 (n24059, n3028, n22399);
  and g39873 (n24060, n3023, n22402);
  and g39874 (n24061, n75, n22595);
  not g39882 (n_15914, n24057);
  not g39883 (n_15915, n24064);
  and g39884 (n24065, n_15914, n_15915);
  not g39885 (n_15916, n24065);
  and g39886 (n24066, n_15914, n_15916);
  and g39887 (n24067, n_15915, n_15916);
  not g39888 (n_15917, n24066);
  not g39889 (n_15918, n24067);
  and g39890 (n24068, n_15917, n_15918);
  not g39891 (n_15919, n24039);
  not g39892 (n_15920, n24068);
  and g39893 (n24069, n_15919, n_15920);
  not g39894 (n_15921, n24069);
  and g39895 (n24070, n_15919, n_15921);
  and g39896 (n24071, n_15920, n_15921);
  not g39897 (n_15922, n24070);
  not g39898 (n_15923, n24071);
  and g39899 (n24072, n_15922, n_15923);
  not g39900 (n_15924, n24038);
  not g39901 (n_15925, n24072);
  and g39902 (n24073, n_15924, n_15925);
  not g39903 (n_15926, n24073);
  and g39904 (n24074, n_15924, n_15926);
  and g39905 (n24075, n_15925, n_15926);
  not g39906 (n_15927, n24074);
  not g39907 (n_15928, n24075);
  and g39908 (n24076, n_15927, n_15928);
  and g39909 (n24077, n_15250, n_15256);
  and g39910 (n24078, n24076, n24077);
  not g39911 (n_15929, n24076);
  not g39912 (n_15930, n24077);
  and g39913 (n24079, n_15929, n_15930);
  not g39914 (n_15931, n24078);
  not g39915 (n_15932, n24079);
  and g39916 (n24080, n_15931, n_15932);
  and g39917 (n24081, n3884, n22377);
  and g39918 (n24082, n3967, n22384);
  and g39919 (n24083, n4046, n22380);
  not g39920 (n_15933, n24082);
  not g39921 (n_15934, n24083);
  and g39922 (n24084, n_15933, n_15934);
  not g39923 (n_15935, n24081);
  and g39924 (n24085, n_15935, n24084);
  and g39925 (n24086, n_750, n24085);
  and g39926 (n24087, n22834, n24085);
  not g39927 (n_15936, n24086);
  not g39928 (n_15937, n24087);
  and g39929 (n24088, n_15936, n_15937);
  not g39930 (n_15938, n24088);
  and g39931 (n24089, \a[26] , n_15938);
  and g39932 (n24090, n_33, n24088);
  not g39933 (n_15939, n24089);
  not g39934 (n_15940, n24090);
  and g39935 (n24091, n_15939, n_15940);
  not g39936 (n_15941, n24091);
  and g39937 (n24092, n24080, n_15941);
  not g39938 (n_15942, n24092);
  and g39939 (n24093, n24080, n_15942);
  and g39940 (n24094, n_15941, n_15942);
  not g39941 (n_15943, n24093);
  not g39942 (n_15944, n24094);
  and g39943 (n24095, n_15943, n_15944);
  not g39944 (n_15945, n24027);
  not g39945 (n_15946, n24095);
  and g39946 (n24096, n_15945, n_15946);
  not g39947 (n_15947, n24096);
  and g39948 (n24097, n_15945, n_15947);
  and g39949 (n24098, n_15946, n_15947);
  not g39950 (n_15948, n24097);
  not g39951 (n_15949, n24098);
  and g39952 (n24099, n_15948, n_15949);
  not g39953 (n_15950, n24026);
  not g39954 (n_15951, n24099);
  and g39955 (n24100, n_15950, n_15951);
  not g39956 (n_15952, n24100);
  and g39957 (n24101, n_15950, n_15952);
  and g39958 (n24102, n_15951, n_15952);
  not g39959 (n_15953, n24101);
  not g39960 (n_15954, n24102);
  and g39961 (n24103, n_15953, n_15954);
  and g39962 (n24104, n_15276, n_15282);
  and g39963 (n24105, n24103, n24104);
  not g39964 (n_15955, n24103);
  not g39965 (n_15956, n24104);
  and g39966 (n24106, n_15955, n_15956);
  not g39967 (n_15957, n24105);
  not g39968 (n_15958, n24106);
  and g39969 (n24107, n_15957, n_15958);
  and g39970 (n24108, n5496, n22359);
  and g39971 (n24109, n4935, n22365);
  and g39972 (n24110, n5407, n22362);
  not g39973 (n_15959, n24109);
  not g39974 (n_15960, n24110);
  and g39975 (n24111, n_15959, n_15960);
  not g39976 (n_15961, n24108);
  and g39977 (n24112, n_15961, n24111);
  and g39978 (n24113, n_1011, n24112);
  and g39979 (n24114, n_15331, n24112);
  not g39980 (n_15962, n24113);
  not g39981 (n_15963, n24114);
  and g39982 (n24115, n_15962, n_15963);
  not g39983 (n_15964, n24115);
  and g39984 (n24116, \a[20] , n_15964);
  and g39985 (n24117, n_435, n24115);
  not g39986 (n_15965, n24116);
  not g39987 (n_15966, n24117);
  and g39988 (n24118, n_15965, n_15966);
  not g39989 (n_15967, n24118);
  and g39990 (n24119, n24107, n_15967);
  not g39991 (n_15968, n24119);
  and g39992 (n24120, n24107, n_15968);
  and g39993 (n24121, n_15967, n_15968);
  not g39994 (n_15969, n24120);
  not g39995 (n_15970, n24121);
  and g39996 (n24122, n_15969, n_15970);
  not g39997 (n_15971, n24015);
  not g39998 (n_15972, n24122);
  and g39999 (n24123, n_15971, n_15972);
  not g40000 (n_15973, n24123);
  and g40001 (n24124, n_15971, n_15973);
  and g40002 (n24125, n_15972, n_15973);
  not g40003 (n_15974, n24124);
  not g40004 (n_15975, n24125);
  and g40005 (n24126, n_15974, n_15975);
  not g40006 (n_15976, n24014);
  not g40007 (n_15977, n24126);
  and g40008 (n24127, n_15976, n_15977);
  not g40009 (n_15978, n24127);
  and g40010 (n24128, n_15976, n_15978);
  and g40011 (n24129, n_15977, n_15978);
  not g40012 (n_15979, n24128);
  not g40013 (n_15980, n24129);
  and g40014 (n24130, n_15979, n_15980);
  and g40015 (n24131, n_15304, n_15566);
  and g40016 (n24132, n24130, n24131);
  not g40017 (n_15981, n24130);
  not g40018 (n_15982, n24131);
  and g40019 (n24133, n_15981, n_15982);
  not g40020 (n_15983, n24132);
  not g40021 (n_15984, n24133);
  and g40022 (n24134, n_15983, n_15984);
  and g40023 (n24135, n7101, n22341);
  and g40024 (n24136, n6402, n22347);
  and g40025 (n24137, n6951, n22344);
  not g40026 (n_15985, n24136);
  not g40027 (n_15986, n24137);
  and g40028 (n24138, n_15985, n_15986);
  not g40029 (n_15987, n24135);
  and g40030 (n24139, n_15987, n24138);
  and g40031 (n24140, n_1885, n24139);
  not g40032 (n_15988, n22482);
  and g40033 (n24141, n22480, n_15988);
  not g40034 (n_15989, n24141);
  and g40035 (n24142, n_14604, n_15989);
  not g40036 (n_15990, n24142);
  and g40037 (n24143, n24139, n_15990);
  not g40038 (n_15991, n24140);
  not g40039 (n_15992, n24143);
  and g40040 (n24144, n_15991, n_15992);
  not g40041 (n_15993, n24144);
  and g40042 (n24145, \a[14] , n_15993);
  and g40043 (n24146, n_652, n24144);
  not g40044 (n_15994, n24145);
  not g40045 (n_15995, n24146);
  and g40046 (n24147, n_15994, n_15995);
  not g40047 (n_15996, n24147);
  and g40048 (n24148, n24134, n_15996);
  not g40049 (n_15997, n24148);
  and g40050 (n24149, n24134, n_15997);
  and g40051 (n24150, n_15996, n_15997);
  not g40052 (n_15998, n24149);
  not g40053 (n_15999, n24150);
  and g40054 (n24151, n_15998, n_15999);
  not g40055 (n_16000, n24003);
  not g40056 (n_16001, n24151);
  and g40057 (n24152, n_16000, n_16001);
  not g40058 (n_16002, n24152);
  and g40059 (n24153, n_16000, n_16002);
  and g40060 (n24154, n_16001, n_16002);
  not g40061 (n_16003, n24153);
  not g40062 (n_16004, n24154);
  and g40063 (n24155, n_16003, n_16004);
  not g40064 (n_16005, n22548);
  not g40065 (n_16006, n24155);
  and g40066 (n24156, n_16005, n_16006);
  not g40067 (n_16007, n24156);
  and g40068 (n24157, n_16005, n_16007);
  and g40069 (n24158, n_16006, n_16007);
  not g40070 (n_16008, n24157);
  not g40071 (n_16009, n24158);
  and g40072 (n24159, n_16008, n_16009);
  and g40073 (n24160, n7983, n22335);
  and g40074 (n24161, n7291, n22341);
  and g40075 (n24162, n7632, n22338);
  and g40081 (n24165, n_14611, n_14614);
  and g40082 (n24166, n_14612, n22492);
  not g40083 (n_16013, n24165);
  not g40084 (n_16014, n24166);
  and g40085 (n24167, n_16013, n_16014);
  not g40086 (n_16015, n24167);
  and g40087 (n24168, n7294, n_16015);
  not g40090 (n_16017, n24169);
  and g40091 (n24170, \a[11] , n_16017);
  not g40092 (n_16018, n24170);
  and g40093 (n24171, n_16017, n_16018);
  and g40094 (n24172, \a[11] , n_16018);
  not g40095 (n_16019, n24171);
  not g40096 (n_16020, n24172);
  and g40097 (n24173, n_16019, n_16020);
  and g40098 (n24174, n_15883, n_15885);
  and g40099 (n24175, n_15884, n_15885);
  not g40100 (n_16021, n24174);
  not g40101 (n_16022, n24175);
  and g40102 (n24176, n_16021, n_16022);
  not g40103 (n_16023, n24173);
  not g40104 (n_16024, n24176);
  and g40105 (n24177, n_16023, n_16024);
  not g40106 (n_16025, n24177);
  and g40107 (n24178, n_16023, n_16025);
  and g40108 (n24179, n_16024, n_16025);
  not g40109 (n_16026, n24178);
  not g40110 (n_16027, n24179);
  and g40111 (n24180, n_16026, n_16027);
  and g40112 (n24181, n7983, n22338);
  and g40113 (n24182, n7291, n22344);
  and g40114 (n24183, n7632, n22341);
  and g40120 (n24186, n_14606, n_14609);
  and g40121 (n24187, n_14607, n22488);
  not g40122 (n_16031, n24186);
  not g40123 (n_16032, n24187);
  and g40124 (n24188, n_16031, n_16032);
  not g40125 (n_16033, n24188);
  and g40126 (n24189, n7294, n_16033);
  not g40129 (n_16035, n24190);
  and g40130 (n24191, \a[11] , n_16035);
  not g40131 (n_16036, n24191);
  and g40132 (n24192, n_16035, n_16036);
  and g40133 (n24193, \a[11] , n_16036);
  not g40134 (n_16037, n24192);
  not g40135 (n_16038, n24193);
  and g40136 (n24194, n_16037, n_16038);
  and g40137 (n24195, n_15877, n_15879);
  and g40138 (n24196, n_15878, n_15879);
  not g40139 (n_16039, n24195);
  not g40140 (n_16040, n24196);
  and g40141 (n24197, n_16039, n_16040);
  not g40142 (n_16041, n24194);
  not g40143 (n_16042, n24197);
  and g40144 (n24198, n_16041, n_16042);
  not g40145 (n_16043, n24198);
  and g40146 (n24199, n_16041, n_16043);
  and g40147 (n24200, n_16042, n_16043);
  not g40148 (n_16044, n24199);
  not g40149 (n_16045, n24200);
  and g40150 (n24201, n_16044, n_16045);
  and g40151 (n24202, n23684, n23991);
  not g40152 (n_16046, n24202);
  and g40153 (n24203, n_15873, n_16046);
  and g40154 (n24204, n7983, n22341);
  and g40155 (n24205, n7291, n22347);
  and g40156 (n24206, n7632, n22344);
  not g40157 (n_16047, n24205);
  not g40158 (n_16048, n24206);
  and g40159 (n24207, n_16047, n_16048);
  not g40160 (n_16049, n24204);
  and g40161 (n24208, n_16049, n24207);
  and g40162 (n24209, n_2446, n24208);
  and g40163 (n24210, n_15990, n24208);
  not g40164 (n_16050, n24209);
  not g40165 (n_16051, n24210);
  and g40166 (n24211, n_16050, n_16051);
  not g40167 (n_16052, n24211);
  and g40168 (n24212, \a[11] , n_16052);
  and g40169 (n24213, n_1071, n24211);
  not g40170 (n_16053, n24212);
  not g40171 (n_16054, n24213);
  and g40172 (n24214, n_16053, n_16054);
  not g40173 (n_16055, n24214);
  and g40174 (n24215, n24203, n_16055);
  and g40175 (n24216, n23702, n23989);
  not g40176 (n_16056, n24216);
  and g40177 (n24217, n_15870, n_16056);
  and g40178 (n24218, n7983, n22344);
  and g40179 (n24219, n7291, n22350);
  and g40180 (n24220, n7632, n22347);
  not g40181 (n_16057, n24219);
  not g40182 (n_16058, n24220);
  and g40183 (n24221, n_16057, n_16058);
  not g40184 (n_16059, n24218);
  and g40185 (n24222, n_16059, n24221);
  and g40186 (n24223, n_2446, n24222);
  and g40187 (n24224, n23642, n24222);
  not g40188 (n_16060, n24223);
  not g40189 (n_16061, n24224);
  and g40190 (n24225, n_16060, n_16061);
  not g40191 (n_16062, n24225);
  and g40192 (n24226, \a[11] , n_16062);
  and g40193 (n24227, n_1071, n24225);
  not g40194 (n_16063, n24226);
  not g40195 (n_16064, n24227);
  and g40196 (n24228, n_16063, n_16064);
  not g40197 (n_16065, n24228);
  and g40198 (n24229, n24217, n_16065);
  and g40199 (n24230, n7983, n22347);
  and g40200 (n24231, n7291, n22353);
  and g40201 (n24232, n7632, n22350);
  not g40207 (n_16069, n23659);
  and g40208 (n24235, n7294, n_16069);
  not g40211 (n_16071, n24236);
  and g40212 (n24237, \a[11] , n_16071);
  not g40213 (n_16072, n24237);
  and g40214 (n24238, n_16071, n_16072);
  and g40215 (n24239, \a[11] , n_16072);
  not g40216 (n_16073, n24238);
  not g40217 (n_16074, n24239);
  and g40218 (n24240, n_16073, n_16074);
  not g40219 (n_16075, n23987);
  and g40220 (n24241, n23985, n_16075);
  not g40221 (n_16076, n24241);
  and g40222 (n24242, n_15867, n_16076);
  not g40223 (n_16077, n24240);
  and g40224 (n24243, n_16077, n24242);
  not g40225 (n_16078, n24243);
  and g40226 (n24244, n_16077, n_16078);
  and g40227 (n24245, n24242, n_16078);
  not g40228 (n_16079, n24244);
  not g40229 (n_16080, n24245);
  and g40230 (n24246, n_16079, n_16080);
  and g40231 (n24247, n7983, n22350);
  and g40232 (n24248, n7291, n22356);
  and g40233 (n24249, n7632, n22353);
  and g40239 (n24252, n7294, n23672);
  not g40242 (n_16085, n24253);
  and g40243 (n24254, \a[11] , n_16085);
  not g40244 (n_16086, n24254);
  and g40245 (n24255, n_16085, n_16086);
  and g40246 (n24256, \a[11] , n_16086);
  not g40247 (n_16087, n24255);
  not g40248 (n_16088, n24256);
  and g40249 (n24257, n_16087, n_16088);
  and g40250 (n24258, n_15860, n_15862);
  and g40251 (n24259, n_15861, n_15862);
  not g40252 (n_16089, n24258);
  not g40253 (n_16090, n24259);
  and g40254 (n24260, n_16089, n_16090);
  not g40255 (n_16091, n24257);
  not g40256 (n_16092, n24260);
  and g40257 (n24261, n_16091, n_16092);
  not g40258 (n_16093, n24261);
  and g40259 (n24262, n_16091, n_16093);
  and g40260 (n24263, n_16092, n_16093);
  not g40261 (n_16094, n24262);
  not g40262 (n_16095, n24263);
  and g40263 (n24264, n_16094, n_16095);
  and g40264 (n24265, n7983, n22353);
  and g40265 (n24266, n7291, n22359);
  and g40266 (n24267, n7632, n22356);
  and g40272 (n24270, n7294, n_14678);
  not g40275 (n_16100, n24271);
  and g40276 (n24272, \a[11] , n_16100);
  not g40277 (n_16101, n24272);
  and g40278 (n24273, n_16100, n_16101);
  and g40279 (n24274, \a[11] , n_16101);
  not g40280 (n_16102, n24273);
  not g40281 (n_16103, n24274);
  and g40282 (n24275, n_16102, n_16103);
  and g40283 (n24276, n_15854, n_15856);
  and g40284 (n24277, n_15855, n_15856);
  not g40285 (n_16104, n24276);
  not g40286 (n_16105, n24277);
  and g40287 (n24278, n_16104, n_16105);
  not g40288 (n_16106, n24275);
  not g40289 (n_16107, n24278);
  and g40290 (n24279, n_16106, n_16107);
  not g40291 (n_16108, n24279);
  and g40292 (n24280, n_16106, n_16108);
  and g40293 (n24281, n_16107, n_16108);
  not g40294 (n_16109, n24280);
  not g40295 (n_16110, n24281);
  and g40296 (n24282, n_16109, n_16110);
  and g40297 (n24283, n23761, n23973);
  not g40298 (n_16111, n24283);
  and g40299 (n24284, n_15850, n_16111);
  and g40300 (n24285, n7983, n22356);
  and g40301 (n24286, n7291, n22362);
  and g40302 (n24287, n7632, n22359);
  not g40303 (n_16112, n24286);
  not g40304 (n_16113, n24287);
  and g40305 (n24288, n_16112, n_16113);
  not g40306 (n_16114, n24285);
  and g40307 (n24289, n_16114, n24288);
  and g40308 (n24290, n_2446, n24289);
  and g40309 (n24291, n23345, n24289);
  not g40310 (n_16115, n24290);
  not g40311 (n_16116, n24291);
  and g40312 (n24292, n_16115, n_16116);
  not g40313 (n_16117, n24292);
  and g40314 (n24293, \a[11] , n_16117);
  and g40315 (n24294, n_1071, n24292);
  not g40316 (n_16118, n24293);
  not g40317 (n_16119, n24294);
  and g40318 (n24295, n_16118, n_16119);
  not g40319 (n_16120, n24295);
  and g40320 (n24296, n24284, n_16120);
  and g40321 (n24297, n23779, n23971);
  not g40322 (n_16121, n24297);
  and g40323 (n24298, n_15847, n_16121);
  and g40324 (n24299, n7983, n22359);
  and g40325 (n24300, n7291, n22365);
  and g40326 (n24301, n7632, n22362);
  not g40327 (n_16122, n24300);
  not g40328 (n_16123, n24301);
  and g40329 (n24302, n_16122, n_16123);
  not g40330 (n_16124, n24299);
  and g40331 (n24303, n_16124, n24302);
  and g40332 (n24304, n_2446, n24303);
  and g40333 (n24305, n_15331, n24303);
  not g40334 (n_16125, n24304);
  not g40335 (n_16126, n24305);
  and g40336 (n24306, n_16125, n_16126);
  not g40337 (n_16127, n24306);
  and g40338 (n24307, \a[11] , n_16127);
  and g40339 (n24308, n_1071, n24306);
  not g40340 (n_16128, n24307);
  not g40341 (n_16129, n24308);
  and g40342 (n24309, n_16128, n_16129);
  not g40343 (n_16130, n24309);
  and g40344 (n24310, n24298, n_16130);
  and g40345 (n24311, n23797, n23969);
  not g40346 (n_16131, n24311);
  and g40347 (n24312, n_15844, n_16131);
  and g40348 (n24313, n7983, n22362);
  and g40349 (n24314, n7291, n22368);
  and g40350 (n24315, n7632, n22365);
  not g40351 (n_16132, n24314);
  not g40352 (n_16133, n24315);
  and g40353 (n24316, n_16132, n_16133);
  not g40354 (n_16134, n24313);
  and g40355 (n24317, n_16134, n24316);
  and g40356 (n24318, n_2446, n24317);
  and g40357 (n24319, n23320, n24317);
  not g40358 (n_16135, n24318);
  not g40359 (n_16136, n24319);
  and g40360 (n24320, n_16135, n_16136);
  not g40361 (n_16137, n24320);
  and g40362 (n24321, \a[11] , n_16137);
  and g40363 (n24322, n_1071, n24320);
  not g40364 (n_16138, n24321);
  not g40365 (n_16139, n24322);
  and g40366 (n24323, n_16138, n_16139);
  not g40367 (n_16140, n24323);
  and g40368 (n24324, n24312, n_16140);
  and g40369 (n24325, n7983, n22365);
  and g40370 (n24326, n7291, n22371);
  and g40371 (n24327, n7632, n22368);
  and g40377 (n24330, n7294, n_15351);
  not g40380 (n_16145, n24331);
  and g40381 (n24332, \a[11] , n_16145);
  not g40382 (n_16146, n24332);
  and g40383 (n24333, n_16145, n_16146);
  and g40384 (n24334, \a[11] , n_16146);
  not g40385 (n_16147, n24333);
  not g40386 (n_16148, n24334);
  and g40387 (n24335, n_16147, n_16148);
  not g40388 (n_16149, n23967);
  and g40389 (n24336, n23965, n_16149);
  not g40390 (n_16150, n24336);
  and g40391 (n24337, n_15841, n_16150);
  not g40392 (n_16151, n24335);
  and g40393 (n24338, n_16151, n24337);
  not g40394 (n_16152, n24338);
  and g40395 (n24339, n_16151, n_16152);
  and g40396 (n24340, n24337, n_16152);
  not g40397 (n_16153, n24339);
  not g40398 (n_16154, n24340);
  and g40399 (n24341, n_16153, n_16154);
  and g40400 (n24342, n7983, n22368);
  and g40401 (n24343, n7291, n22374);
  and g40402 (n24344, n7632, n22371);
  and g40408 (n24347, n7294, n23006);
  not g40411 (n_16159, n24348);
  and g40412 (n24349, \a[11] , n_16159);
  not g40413 (n_16160, n24349);
  and g40414 (n24350, n_16159, n_16160);
  and g40415 (n24351, \a[11] , n_16160);
  not g40416 (n_16161, n24350);
  not g40417 (n_16162, n24351);
  and g40418 (n24352, n_16161, n_16162);
  and g40419 (n24353, n_15834, n_15836);
  and g40420 (n24354, n_15835, n_15836);
  not g40421 (n_16163, n24353);
  not g40422 (n_16164, n24354);
  and g40423 (n24355, n_16163, n_16164);
  not g40424 (n_16165, n24352);
  not g40425 (n_16166, n24355);
  and g40426 (n24356, n_16165, n_16166);
  not g40427 (n_16167, n24356);
  and g40428 (n24357, n_16165, n_16167);
  and g40429 (n24358, n_16166, n_16167);
  not g40430 (n_16168, n24357);
  not g40431 (n_16169, n24358);
  and g40432 (n24359, n_16168, n_16169);
  and g40433 (n24360, n7983, n22371);
  and g40434 (n24361, n7291, n22377);
  and g40435 (n24362, n7632, n22374);
  and g40441 (n24365, n7294, n23025);
  not g40444 (n_16174, n24366);
  and g40445 (n24367, \a[11] , n_16174);
  not g40446 (n_16175, n24367);
  and g40447 (n24368, n_16174, n_16175);
  and g40448 (n24369, \a[11] , n_16175);
  not g40449 (n_16176, n24368);
  not g40450 (n_16177, n24369);
  and g40451 (n24370, n_16176, n_16177);
  and g40452 (n24371, n_15828, n_15830);
  and g40453 (n24372, n_15829, n_15830);
  not g40454 (n_16178, n24371);
  not g40455 (n_16179, n24372);
  and g40456 (n24373, n_16178, n_16179);
  not g40457 (n_16180, n24370);
  not g40458 (n_16181, n24373);
  and g40459 (n24374, n_16180, n_16181);
  not g40460 (n_16182, n24374);
  and g40461 (n24375, n_16180, n_16182);
  and g40462 (n24376, n_16181, n_16182);
  not g40463 (n_16183, n24375);
  not g40464 (n_16184, n24376);
  and g40465 (n24377, n_16183, n_16184);
  and g40466 (n24378, n23856, n23953);
  not g40467 (n_16185, n24378);
  and g40468 (n24379, n_15824, n_16185);
  and g40469 (n24380, n7983, n22374);
  and g40470 (n24381, n7291, n22380);
  and g40471 (n24382, n7632, n22377);
  not g40472 (n_16186, n24381);
  not g40473 (n_16187, n24382);
  and g40474 (n24383, n_16186, n_16187);
  not g40475 (n_16188, n24380);
  and g40476 (n24384, n_16188, n24383);
  and g40477 (n24385, n_2446, n24384);
  and g40478 (n24386, n_15064, n24384);
  not g40479 (n_16189, n24385);
  not g40480 (n_16190, n24386);
  and g40481 (n24387, n_16189, n_16190);
  not g40482 (n_16191, n24387);
  and g40483 (n24388, \a[11] , n_16191);
  and g40484 (n24389, n_1071, n24387);
  not g40485 (n_16192, n24388);
  not g40486 (n_16193, n24389);
  and g40487 (n24390, n_16192, n_16193);
  not g40488 (n_16194, n24390);
  and g40489 (n24391, n24379, n_16194);
  not g40490 (n_16195, n23951);
  and g40491 (n24392, n23949, n_16195);
  not g40492 (n_16196, n24392);
  and g40493 (n24393, n_15821, n_16196);
  and g40494 (n24394, n7983, n22377);
  and g40495 (n24395, n7291, n22384);
  and g40496 (n24396, n7632, n22380);
  not g40497 (n_16197, n24395);
  not g40498 (n_16198, n24396);
  and g40499 (n24397, n_16197, n_16198);
  not g40500 (n_16199, n24394);
  and g40501 (n24398, n_16199, n24397);
  and g40502 (n24399, n_2446, n24398);
  and g40503 (n24400, n22834, n24398);
  not g40504 (n_16200, n24399);
  not g40505 (n_16201, n24400);
  and g40506 (n24401, n_16200, n_16201);
  not g40507 (n_16202, n24401);
  and g40508 (n24402, \a[11] , n_16202);
  and g40509 (n24403, n_1071, n24401);
  not g40510 (n_16203, n24402);
  not g40511 (n_16204, n24403);
  and g40512 (n24404, n_16203, n_16204);
  not g40513 (n_16205, n24404);
  and g40514 (n24405, n24393, n_16205);
  and g40515 (n24406, n23888, n23947);
  not g40516 (n_16206, n24406);
  and g40517 (n24407, n_15817, n_16206);
  and g40518 (n24408, n7983, n22380);
  and g40519 (n24409, n7291, n22387);
  and g40520 (n24410, n7632, n22384);
  not g40521 (n_16207, n24409);
  not g40522 (n_16208, n24410);
  and g40523 (n24411, n_16207, n_16208);
  not g40524 (n_16209, n24408);
  and g40525 (n24412, n_16209, n24411);
  and g40526 (n24413, n_2446, n24412);
  and g40527 (n24414, n_14894, n24412);
  not g40528 (n_16210, n24413);
  not g40529 (n_16211, n24414);
  and g40530 (n24415, n_16210, n_16211);
  not g40531 (n_16212, n24415);
  and g40532 (n24416, \a[11] , n_16212);
  and g40533 (n24417, n_1071, n24415);
  not g40534 (n_16213, n24416);
  not g40535 (n_16214, n24417);
  and g40536 (n24418, n_16213, n_16214);
  not g40537 (n_16215, n24418);
  and g40538 (n24419, n24407, n_16215);
  and g40539 (n24420, n7983, n22384);
  and g40540 (n24421, n7291, n22390);
  and g40541 (n24422, n7632, n22387);
  and g40547 (n24425, n7294, n22806);
  not g40550 (n_16220, n24426);
  and g40551 (n24427, \a[11] , n_16220);
  not g40552 (n_16221, n24427);
  and g40553 (n24428, n_16220, n_16221);
  and g40554 (n24429, \a[11] , n_16221);
  not g40555 (n_16222, n24428);
  not g40556 (n_16223, n24429);
  and g40557 (n24430, n_16222, n_16223);
  not g40558 (n_16224, n23945);
  and g40559 (n24431, n23943, n_16224);
  not g40560 (n_16225, n24431);
  and g40561 (n24432, n_15814, n_16225);
  not g40562 (n_16226, n24430);
  and g40563 (n24433, n_16226, n24432);
  not g40564 (n_16227, n24433);
  and g40565 (n24434, n_16226, n_16227);
  and g40566 (n24435, n24432, n_16227);
  not g40567 (n_16228, n24434);
  not g40568 (n_16229, n24435);
  and g40569 (n24436, n_16228, n_16229);
  and g40570 (n24437, n_15807, n_15809);
  and g40571 (n24438, n_15808, n_15809);
  not g40572 (n_16230, n24437);
  not g40573 (n_16231, n24438);
  and g40574 (n24439, n_16230, n_16231);
  and g40575 (n24440, n7983, n22387);
  and g40576 (n24441, n7291, n22393);
  and g40577 (n24442, n7632, n22390);
  not g40578 (n_16232, n24441);
  not g40579 (n_16233, n24442);
  and g40580 (n24443, n_16232, n_16233);
  not g40581 (n_16234, n24440);
  and g40582 (n24444, n_16234, n24443);
  and g40583 (n24445, n_2446, n24444);
  and g40584 (n24446, n_14920, n24444);
  not g40585 (n_16235, n24445);
  not g40586 (n_16236, n24446);
  and g40587 (n24447, n_16235, n_16236);
  not g40588 (n_16237, n24447);
  and g40589 (n24448, \a[11] , n_16237);
  and g40590 (n24449, n_1071, n24447);
  not g40591 (n_16238, n24448);
  not g40592 (n_16239, n24449);
  and g40593 (n24450, n_16238, n_16239);
  not g40594 (n_16240, n24439);
  not g40595 (n_16241, n24450);
  and g40596 (n24451, n_16240, n_16241);
  and g40597 (n24452, n7983, n22390);
  and g40598 (n24453, n7291, n22396);
  and g40599 (n24454, n7632, n22393);
  and g40605 (n24457, n7294, n22649);
  not g40608 (n_16246, n24458);
  and g40609 (n24459, \a[11] , n_16246);
  not g40610 (n_16247, n24459);
  and g40611 (n24460, n_16246, n_16247);
  and g40612 (n24461, \a[11] , n_16247);
  not g40613 (n_16248, n24460);
  not g40614 (n_16249, n24461);
  and g40615 (n24462, n_16248, n_16249);
  not g40616 (n_16250, n23914);
  and g40617 (n24463, n_16250, n23925);
  not g40618 (n_16251, n23926);
  not g40619 (n_16252, n24463);
  and g40620 (n24464, n_16251, n_16252);
  not g40621 (n_16253, n24462);
  and g40622 (n24465, n_16253, n24464);
  not g40623 (n_16254, n24465);
  and g40624 (n24466, n_16253, n_16254);
  and g40625 (n24467, n24464, n_16254);
  not g40626 (n_16255, n24466);
  not g40627 (n_16256, n24467);
  and g40628 (n24468, n_16255, n_16256);
  not g40629 (n_16257, n23913);
  and g40630 (n24469, n23911, n_16257);
  not g40631 (n_16258, n24469);
  and g40632 (n24470, n_16250, n_16258);
  and g40633 (n24471, n7983, n22393);
  and g40634 (n24472, n7291, n22399);
  and g40635 (n24473, n7632, n22396);
  not g40636 (n_16259, n24472);
  not g40637 (n_16260, n24473);
  and g40638 (n24474, n_16259, n_16260);
  not g40639 (n_16261, n24471);
  and g40640 (n24475, n_16261, n24474);
  and g40641 (n24476, n_2446, n24475);
  and g40642 (n24477, n_14773, n24475);
  not g40643 (n_16262, n24476);
  not g40644 (n_16263, n24477);
  and g40645 (n24478, n_16262, n_16263);
  not g40646 (n_16264, n24478);
  and g40647 (n24479, \a[11] , n_16264);
  and g40648 (n24480, n_1071, n24478);
  not g40649 (n_16265, n24479);
  not g40650 (n_16266, n24480);
  and g40651 (n24481, n_16265, n_16266);
  not g40652 (n_16267, n24481);
  and g40653 (n24482, n24470, n_16267);
  and g40654 (n24483, n7632, n_14508);
  and g40655 (n24484, n7983, n22402);
  not g40656 (n_16268, n24483);
  not g40657 (n_16269, n24484);
  and g40658 (n24485, n_16268, n_16269);
  and g40659 (n24486, n7294, n_14720);
  not g40660 (n_16270, n24486);
  and g40661 (n24487, n24485, n_16270);
  not g40662 (n_16271, n24487);
  and g40663 (n24488, \a[11] , n_16271);
  not g40664 (n_16272, n24488);
  and g40665 (n24489, \a[11] , n_16272);
  and g40666 (n24490, n_16271, n_16272);
  not g40667 (n_16273, n24489);
  not g40668 (n_16274, n24490);
  and g40669 (n24491, n_16273, n_16274);
  and g40670 (n24492, n_2445, n_14508);
  not g40671 (n_16275, n24492);
  and g40672 (n24493, \a[11] , n_16275);
  not g40673 (n_16276, n24491);
  and g40674 (n24494, n_16276, n24493);
  and g40675 (n24495, n7983, n22399);
  and g40676 (n24496, n7291, n_14508);
  and g40677 (n24497, n7632, n22402);
  not g40678 (n_16277, n24496);
  not g40679 (n_16278, n24497);
  and g40680 (n24498, n_16277, n_16278);
  not g40681 (n_16279, n24495);
  and g40682 (n24499, n_16279, n24498);
  and g40683 (n24500, n_2446, n24499);
  and g40684 (n24501, n22625, n24499);
  not g40685 (n_16280, n24500);
  not g40686 (n_16281, n24501);
  and g40687 (n24502, n_16280, n_16281);
  not g40688 (n_16282, n24502);
  and g40689 (n24503, \a[11] , n_16282);
  and g40690 (n24504, n_1071, n24502);
  not g40691 (n_16283, n24503);
  not g40692 (n_16284, n24504);
  and g40693 (n24505, n_16283, n_16284);
  not g40694 (n_16285, n24505);
  and g40695 (n24506, n24494, n_16285);
  and g40696 (n24507, n23912, n24506);
  not g40697 (n_16286, n24507);
  and g40698 (n24508, n24506, n_16286);
  and g40699 (n24509, n23912, n_16286);
  not g40700 (n_16287, n24508);
  not g40701 (n_16288, n24509);
  and g40702 (n24510, n_16287, n_16288);
  and g40703 (n24511, n7983, n22396);
  and g40704 (n24512, n7291, n22402);
  and g40705 (n24513, n7632, n22399);
  and g40711 (n24516, n7294, n22595);
  not g40714 (n_16293, n24517);
  and g40715 (n24518, \a[11] , n_16293);
  not g40716 (n_16294, n24518);
  and g40717 (n24519, \a[11] , n_16294);
  and g40718 (n24520, n_16293, n_16294);
  not g40719 (n_16295, n24519);
  not g40720 (n_16296, n24520);
  and g40721 (n24521, n_16295, n_16296);
  not g40722 (n_16297, n24510);
  not g40723 (n_16298, n24521);
  and g40724 (n24522, n_16297, n_16298);
  not g40725 (n_16299, n24522);
  and g40726 (n24523, n_16286, n_16299);
  not g40727 (n_16300, n24470);
  and g40728 (n24524, n_16300, n24481);
  not g40729 (n_16301, n24482);
  not g40730 (n_16302, n24524);
  and g40731 (n24525, n_16301, n_16302);
  not g40732 (n_16303, n24523);
  and g40733 (n24526, n_16303, n24525);
  not g40734 (n_16304, n24526);
  and g40735 (n24527, n_16301, n_16304);
  not g40736 (n_16305, n24468);
  not g40737 (n_16306, n24527);
  and g40738 (n24528, n_16305, n_16306);
  not g40739 (n_16307, n24528);
  and g40740 (n24529, n_16254, n_16307);
  and g40741 (n24530, n24439, n24450);
  not g40742 (n_16308, n24451);
  not g40743 (n_16309, n24530);
  and g40744 (n24531, n_16308, n_16309);
  not g40745 (n_16310, n24529);
  and g40746 (n24532, n_16310, n24531);
  not g40747 (n_16311, n24532);
  and g40748 (n24533, n_16308, n_16311);
  not g40749 (n_16312, n24436);
  not g40750 (n_16313, n24533);
  and g40751 (n24534, n_16312, n_16313);
  not g40752 (n_16314, n24534);
  and g40753 (n24535, n_16227, n_16314);
  not g40754 (n_16315, n24419);
  and g40755 (n24536, n24407, n_16315);
  and g40756 (n24537, n_16215, n_16315);
  not g40757 (n_16316, n24536);
  not g40758 (n_16317, n24537);
  and g40759 (n24538, n_16316, n_16317);
  not g40760 (n_16318, n24535);
  not g40761 (n_16319, n24538);
  and g40762 (n24539, n_16318, n_16319);
  not g40763 (n_16320, n24539);
  and g40764 (n24540, n_16315, n_16320);
  not g40765 (n_16321, n24405);
  and g40766 (n24541, n24393, n_16321);
  and g40767 (n24542, n_16205, n_16321);
  not g40768 (n_16322, n24541);
  not g40769 (n_16323, n24542);
  and g40770 (n24543, n_16322, n_16323);
  not g40771 (n_16324, n24540);
  not g40772 (n_16325, n24543);
  and g40773 (n24544, n_16324, n_16325);
  not g40774 (n_16326, n24544);
  and g40775 (n24545, n_16321, n_16326);
  not g40776 (n_16327, n24379);
  and g40777 (n24546, n_16327, n24390);
  not g40778 (n_16328, n24391);
  not g40779 (n_16329, n24546);
  and g40780 (n24547, n_16328, n_16329);
  not g40781 (n_16330, n24545);
  and g40782 (n24548, n_16330, n24547);
  not g40783 (n_16331, n24548);
  and g40784 (n24549, n_16328, n_16331);
  not g40785 (n_16332, n24377);
  not g40786 (n_16333, n24549);
  and g40787 (n24550, n_16332, n_16333);
  not g40788 (n_16334, n24550);
  and g40789 (n24551, n_16182, n_16334);
  not g40790 (n_16335, n24359);
  not g40791 (n_16336, n24551);
  and g40792 (n24552, n_16335, n_16336);
  not g40793 (n_16337, n24552);
  and g40794 (n24553, n_16167, n_16337);
  not g40795 (n_16338, n24341);
  not g40796 (n_16339, n24553);
  and g40797 (n24554, n_16338, n_16339);
  not g40798 (n_16340, n24554);
  and g40799 (n24555, n_16152, n_16340);
  not g40800 (n_16341, n24324);
  and g40801 (n24556, n24312, n_16341);
  and g40802 (n24557, n_16140, n_16341);
  not g40803 (n_16342, n24556);
  not g40804 (n_16343, n24557);
  and g40805 (n24558, n_16342, n_16343);
  not g40806 (n_16344, n24555);
  not g40807 (n_16345, n24558);
  and g40808 (n24559, n_16344, n_16345);
  not g40809 (n_16346, n24559);
  and g40810 (n24560, n_16341, n_16346);
  not g40811 (n_16347, n24310);
  and g40812 (n24561, n24298, n_16347);
  and g40813 (n24562, n_16130, n_16347);
  not g40814 (n_16348, n24561);
  not g40815 (n_16349, n24562);
  and g40816 (n24563, n_16348, n_16349);
  not g40817 (n_16350, n24560);
  not g40818 (n_16351, n24563);
  and g40819 (n24564, n_16350, n_16351);
  not g40820 (n_16352, n24564);
  and g40821 (n24565, n_16347, n_16352);
  not g40822 (n_16353, n24284);
  and g40823 (n24566, n_16353, n24295);
  not g40824 (n_16354, n24296);
  not g40825 (n_16355, n24566);
  and g40826 (n24567, n_16354, n_16355);
  not g40827 (n_16356, n24565);
  and g40828 (n24568, n_16356, n24567);
  not g40829 (n_16357, n24568);
  and g40830 (n24569, n_16354, n_16357);
  not g40831 (n_16358, n24282);
  not g40832 (n_16359, n24569);
  and g40833 (n24570, n_16358, n_16359);
  not g40834 (n_16360, n24570);
  and g40835 (n24571, n_16108, n_16360);
  not g40836 (n_16361, n24264);
  not g40837 (n_16362, n24571);
  and g40838 (n24572, n_16361, n_16362);
  not g40839 (n_16363, n24572);
  and g40840 (n24573, n_16093, n_16363);
  not g40841 (n_16364, n24246);
  not g40842 (n_16365, n24573);
  and g40843 (n24574, n_16364, n_16365);
  not g40844 (n_16366, n24574);
  and g40845 (n24575, n_16078, n_16366);
  not g40846 (n_16367, n24229);
  and g40847 (n24576, n24217, n_16367);
  and g40848 (n24577, n_16065, n_16367);
  not g40849 (n_16368, n24576);
  not g40850 (n_16369, n24577);
  and g40851 (n24578, n_16368, n_16369);
  not g40852 (n_16370, n24575);
  not g40853 (n_16371, n24578);
  and g40854 (n24579, n_16370, n_16371);
  not g40855 (n_16372, n24579);
  and g40856 (n24580, n_16367, n_16372);
  not g40857 (n_16373, n24203);
  and g40858 (n24581, n_16373, n24214);
  not g40859 (n_16374, n24215);
  not g40860 (n_16375, n24581);
  and g40861 (n24582, n_16374, n_16375);
  not g40862 (n_16376, n24580);
  and g40863 (n24583, n_16376, n24582);
  not g40864 (n_16377, n24583);
  and g40865 (n24584, n_16374, n_16377);
  not g40866 (n_16378, n24201);
  not g40867 (n_16379, n24584);
  and g40868 (n24585, n_16378, n_16379);
  not g40869 (n_16380, n24585);
  and g40870 (n24586, n_16043, n_16380);
  not g40871 (n_16381, n24180);
  not g40872 (n_16382, n24586);
  and g40873 (n24587, n_16381, n_16382);
  not g40874 (n_16383, n24587);
  and g40875 (n24588, n_16025, n_16383);
  and g40876 (n24589, n24159, n24588);
  not g40877 (n_16384, n24159);
  not g40878 (n_16385, n24588);
  and g40879 (n24590, n_16384, n_16385);
  not g40880 (n_16386, n24589);
  not g40881 (n_16387, n24590);
  and g40882 (n24591, n_16386, n_16387);
  and g40883 (n24592, n9331, n22323);
  and g40884 (n24593, n8418, n22329);
  and g40885 (n24594, n8860, n22326);
  not g40886 (n_16388, n24593);
  not g40887 (n_16389, n24594);
  and g40888 (n24595, n_16388, n_16389);
  not g40889 (n_16390, n24592);
  and g40890 (n24596, n_16390, n24595);
  and g40891 (n24597, n_3428, n24596);
  not g40892 (n_16391, n22506);
  and g40893 (n24598, n22504, n_16391);
  not g40894 (n_16392, n24598);
  and g40895 (n24599, n_14634, n_16392);
  not g40896 (n_16393, n24599);
  and g40897 (n24600, n24596, n_16393);
  not g40898 (n_16394, n24597);
  not g40899 (n_16395, n24600);
  and g40900 (n24601, n_16394, n_16395);
  not g40901 (n_16396, n24601);
  and g40902 (n24602, \a[8] , n_16396);
  and g40903 (n24603, n_1106, n24601);
  not g40904 (n_16397, n24602);
  not g40905 (n_16398, n24603);
  and g40906 (n24604, n_16397, n_16398);
  not g40907 (n_16399, n24604);
  and g40908 (n24605, n24591, n_16399);
  and g40909 (n24606, n24180, n24586);
  not g40910 (n_16400, n24606);
  and g40911 (n24607, n_16383, n_16400);
  and g40912 (n24608, n9331, n22326);
  and g40913 (n24609, n8418, n22332);
  and g40914 (n24610, n8860, n22329);
  not g40915 (n_16401, n24609);
  not g40916 (n_16402, n24610);
  and g40917 (n24611, n_16401, n_16402);
  not g40918 (n_16403, n24608);
  and g40919 (n24612, n_16403, n24611);
  and g40920 (n24613, n_3428, n24612);
  and g40921 (n24614, n_14626, n_14629);
  and g40922 (n24615, n_14627, n22504);
  not g40923 (n_16404, n24614);
  not g40924 (n_16405, n24615);
  and g40925 (n24616, n_16404, n_16405);
  and g40926 (n24617, n24612, n24616);
  not g40927 (n_16406, n24613);
  not g40928 (n_16407, n24617);
  and g40929 (n24618, n_16406, n_16407);
  not g40930 (n_16408, n24618);
  and g40931 (n24619, \a[8] , n_16408);
  and g40932 (n24620, n_1106, n24618);
  not g40933 (n_16409, n24619);
  not g40934 (n_16410, n24620);
  and g40935 (n24621, n_16409, n_16410);
  not g40936 (n_16411, n24621);
  and g40937 (n24622, n24607, n_16411);
  and g40938 (n24623, n24201, n24584);
  not g40939 (n_16412, n24623);
  and g40940 (n24624, n_16380, n_16412);
  and g40941 (n24625, n9331, n22329);
  and g40942 (n24626, n8418, n22335);
  and g40943 (n24627, n8860, n22332);
  not g40944 (n_16413, n24626);
  not g40945 (n_16414, n24627);
  and g40946 (n24628, n_16413, n_16414);
  not g40947 (n_16415, n24625);
  and g40948 (n24629, n_16415, n24628);
  and g40949 (n24630, n_3428, n24629);
  and g40950 (n24631, n_14621, n_14624);
  and g40951 (n24632, n_14622, n22500);
  not g40952 (n_16416, n24631);
  not g40953 (n_16417, n24632);
  and g40954 (n24633, n_16416, n_16417);
  and g40955 (n24634, n24629, n24633);
  not g40956 (n_16418, n24630);
  not g40957 (n_16419, n24634);
  and g40958 (n24635, n_16418, n_16419);
  not g40959 (n_16420, n24635);
  and g40960 (n24636, \a[8] , n_16420);
  and g40961 (n24637, n_1106, n24635);
  not g40962 (n_16421, n24636);
  not g40963 (n_16422, n24637);
  and g40964 (n24638, n_16421, n_16422);
  not g40965 (n_16423, n24638);
  and g40966 (n24639, n24624, n_16423);
  and g40967 (n24640, n9331, n22332);
  and g40968 (n24641, n8418, n22338);
  and g40969 (n24642, n8860, n22335);
  and g40975 (n24645, n8421, n22542);
  not g40978 (n_16428, n24646);
  and g40979 (n24647, \a[8] , n_16428);
  not g40980 (n_16429, n24647);
  and g40981 (n24648, n_16428, n_16429);
  and g40982 (n24649, \a[8] , n_16429);
  not g40983 (n_16430, n24648);
  not g40984 (n_16431, n24649);
  and g40985 (n24650, n_16430, n_16431);
  not g40986 (n_16432, n24582);
  and g40987 (n24651, n24580, n_16432);
  not g40988 (n_16433, n24651);
  and g40989 (n24652, n_16377, n_16433);
  not g40990 (n_16434, n24650);
  and g40991 (n24653, n_16434, n24652);
  not g40992 (n_16435, n24653);
  and g40993 (n24654, n_16434, n_16435);
  and g40994 (n24655, n24652, n_16435);
  not g40995 (n_16436, n24654);
  not g40996 (n_16437, n24655);
  and g40997 (n24656, n_16436, n_16437);
  and g40998 (n24657, n9331, n22335);
  and g40999 (n24658, n8418, n22341);
  and g41000 (n24659, n8860, n22338);
  and g41006 (n24662, n8421, n_16015);
  not g41009 (n_16442, n24663);
  and g41010 (n24664, \a[8] , n_16442);
  not g41011 (n_16443, n24664);
  and g41012 (n24665, n_16442, n_16443);
  and g41013 (n24666, \a[8] , n_16443);
  not g41014 (n_16444, n24665);
  not g41015 (n_16445, n24666);
  and g41016 (n24667, n_16444, n_16445);
  and g41017 (n24668, n_16370, n_16372);
  and g41018 (n24669, n_16371, n_16372);
  not g41019 (n_16446, n24668);
  not g41020 (n_16447, n24669);
  and g41021 (n24670, n_16446, n_16447);
  not g41022 (n_16448, n24667);
  not g41023 (n_16449, n24670);
  and g41024 (n24671, n_16448, n_16449);
  not g41025 (n_16450, n24671);
  and g41026 (n24672, n_16448, n_16450);
  and g41027 (n24673, n_16449, n_16450);
  not g41028 (n_16451, n24672);
  not g41029 (n_16452, n24673);
  and g41030 (n24674, n_16451, n_16452);
  and g41031 (n24675, n24246, n24573);
  not g41032 (n_16453, n24675);
  and g41033 (n24676, n_16366, n_16453);
  and g41034 (n24677, n9331, n22338);
  and g41035 (n24678, n8418, n22344);
  and g41036 (n24679, n8860, n22341);
  not g41037 (n_16454, n24678);
  not g41038 (n_16455, n24679);
  and g41039 (n24680, n_16454, n_16455);
  not g41040 (n_16456, n24677);
  and g41041 (n24681, n_16456, n24680);
  and g41042 (n24682, n_3428, n24681);
  and g41043 (n24683, n24188, n24681);
  not g41044 (n_16457, n24682);
  not g41045 (n_16458, n24683);
  and g41046 (n24684, n_16457, n_16458);
  not g41047 (n_16459, n24684);
  and g41048 (n24685, \a[8] , n_16459);
  and g41049 (n24686, n_1106, n24684);
  not g41050 (n_16460, n24685);
  not g41051 (n_16461, n24686);
  and g41052 (n24687, n_16460, n_16461);
  not g41053 (n_16462, n24687);
  and g41054 (n24688, n24676, n_16462);
  and g41055 (n24689, n24264, n24571);
  not g41056 (n_16463, n24689);
  and g41057 (n24690, n_16363, n_16463);
  and g41058 (n24691, n9331, n22341);
  and g41059 (n24692, n8418, n22347);
  and g41060 (n24693, n8860, n22344);
  not g41061 (n_16464, n24692);
  not g41062 (n_16465, n24693);
  and g41063 (n24694, n_16464, n_16465);
  not g41064 (n_16466, n24691);
  and g41065 (n24695, n_16466, n24694);
  and g41066 (n24696, n_3428, n24695);
  and g41067 (n24697, n_15990, n24695);
  not g41068 (n_16467, n24696);
  not g41069 (n_16468, n24697);
  and g41070 (n24698, n_16467, n_16468);
  not g41071 (n_16469, n24698);
  and g41072 (n24699, \a[8] , n_16469);
  and g41073 (n24700, n_1106, n24698);
  not g41074 (n_16470, n24699);
  not g41075 (n_16471, n24700);
  and g41076 (n24701, n_16470, n_16471);
  not g41077 (n_16472, n24701);
  and g41078 (n24702, n24690, n_16472);
  and g41079 (n24703, n24282, n24569);
  not g41080 (n_16473, n24703);
  and g41081 (n24704, n_16360, n_16473);
  and g41082 (n24705, n9331, n22344);
  and g41083 (n24706, n8418, n22350);
  and g41084 (n24707, n8860, n22347);
  not g41085 (n_16474, n24706);
  not g41086 (n_16475, n24707);
  and g41087 (n24708, n_16474, n_16475);
  not g41088 (n_16476, n24705);
  and g41089 (n24709, n_16476, n24708);
  and g41090 (n24710, n_3428, n24709);
  and g41091 (n24711, n23642, n24709);
  not g41092 (n_16477, n24710);
  not g41093 (n_16478, n24711);
  and g41094 (n24712, n_16477, n_16478);
  not g41095 (n_16479, n24712);
  and g41096 (n24713, \a[8] , n_16479);
  and g41097 (n24714, n_1106, n24712);
  not g41098 (n_16480, n24713);
  not g41099 (n_16481, n24714);
  and g41100 (n24715, n_16480, n_16481);
  not g41101 (n_16482, n24715);
  and g41102 (n24716, n24704, n_16482);
  and g41103 (n24717, n9331, n22347);
  and g41104 (n24718, n8418, n22353);
  and g41105 (n24719, n8860, n22350);
  and g41111 (n24722, n8421, n_16069);
  not g41114 (n_16487, n24723);
  and g41115 (n24724, \a[8] , n_16487);
  not g41116 (n_16488, n24724);
  and g41117 (n24725, n_16487, n_16488);
  and g41118 (n24726, \a[8] , n_16488);
  not g41119 (n_16489, n24725);
  not g41120 (n_16490, n24726);
  and g41121 (n24727, n_16489, n_16490);
  not g41122 (n_16491, n24567);
  and g41123 (n24728, n24565, n_16491);
  not g41124 (n_16492, n24728);
  and g41125 (n24729, n_16357, n_16492);
  not g41126 (n_16493, n24727);
  and g41127 (n24730, n_16493, n24729);
  not g41128 (n_16494, n24730);
  and g41129 (n24731, n_16493, n_16494);
  and g41130 (n24732, n24729, n_16494);
  not g41131 (n_16495, n24731);
  not g41132 (n_16496, n24732);
  and g41133 (n24733, n_16495, n_16496);
  and g41134 (n24734, n9331, n22350);
  and g41135 (n24735, n8418, n22356);
  and g41136 (n24736, n8860, n22353);
  and g41142 (n24739, n8421, n23672);
  not g41145 (n_16501, n24740);
  and g41146 (n24741, \a[8] , n_16501);
  not g41147 (n_16502, n24741);
  and g41148 (n24742, n_16501, n_16502);
  and g41149 (n24743, \a[8] , n_16502);
  not g41150 (n_16503, n24742);
  not g41151 (n_16504, n24743);
  and g41152 (n24744, n_16503, n_16504);
  and g41153 (n24745, n_16350, n_16352);
  and g41154 (n24746, n_16351, n_16352);
  not g41155 (n_16505, n24745);
  not g41156 (n_16506, n24746);
  and g41157 (n24747, n_16505, n_16506);
  not g41158 (n_16507, n24744);
  not g41159 (n_16508, n24747);
  and g41160 (n24748, n_16507, n_16508);
  not g41161 (n_16509, n24748);
  and g41162 (n24749, n_16507, n_16509);
  and g41163 (n24750, n_16508, n_16509);
  not g41164 (n_16510, n24749);
  not g41165 (n_16511, n24750);
  and g41166 (n24751, n_16510, n_16511);
  and g41167 (n24752, n9331, n22353);
  and g41168 (n24753, n8418, n22359);
  and g41169 (n24754, n8860, n22356);
  and g41175 (n24757, n8421, n_14678);
  not g41178 (n_16516, n24758);
  and g41179 (n24759, \a[8] , n_16516);
  not g41180 (n_16517, n24759);
  and g41181 (n24760, n_16516, n_16517);
  and g41182 (n24761, \a[8] , n_16517);
  not g41183 (n_16518, n24760);
  not g41184 (n_16519, n24761);
  and g41185 (n24762, n_16518, n_16519);
  and g41186 (n24763, n_16344, n_16346);
  and g41187 (n24764, n_16345, n_16346);
  not g41188 (n_16520, n24763);
  not g41189 (n_16521, n24764);
  and g41190 (n24765, n_16520, n_16521);
  not g41191 (n_16522, n24762);
  not g41192 (n_16523, n24765);
  and g41193 (n24766, n_16522, n_16523);
  not g41194 (n_16524, n24766);
  and g41195 (n24767, n_16522, n_16524);
  and g41196 (n24768, n_16523, n_16524);
  not g41197 (n_16525, n24767);
  not g41198 (n_16526, n24768);
  and g41199 (n24769, n_16525, n_16526);
  and g41200 (n24770, n24341, n24553);
  not g41201 (n_16527, n24770);
  and g41202 (n24771, n_16340, n_16527);
  and g41203 (n24772, n9331, n22356);
  and g41204 (n24773, n8418, n22362);
  and g41205 (n24774, n8860, n22359);
  not g41206 (n_16528, n24773);
  not g41207 (n_16529, n24774);
  and g41208 (n24775, n_16528, n_16529);
  not g41209 (n_16530, n24772);
  and g41210 (n24776, n_16530, n24775);
  and g41211 (n24777, n_3428, n24776);
  and g41212 (n24778, n23345, n24776);
  not g41213 (n_16531, n24777);
  not g41214 (n_16532, n24778);
  and g41215 (n24779, n_16531, n_16532);
  not g41216 (n_16533, n24779);
  and g41217 (n24780, \a[8] , n_16533);
  and g41218 (n24781, n_1106, n24779);
  not g41219 (n_16534, n24780);
  not g41220 (n_16535, n24781);
  and g41221 (n24782, n_16534, n_16535);
  not g41222 (n_16536, n24782);
  and g41223 (n24783, n24771, n_16536);
  and g41224 (n24784, n24359, n24551);
  not g41225 (n_16537, n24784);
  and g41226 (n24785, n_16337, n_16537);
  and g41227 (n24786, n9331, n22359);
  and g41228 (n24787, n8418, n22365);
  and g41229 (n24788, n8860, n22362);
  not g41230 (n_16538, n24787);
  not g41231 (n_16539, n24788);
  and g41232 (n24789, n_16538, n_16539);
  not g41233 (n_16540, n24786);
  and g41234 (n24790, n_16540, n24789);
  and g41235 (n24791, n_3428, n24790);
  and g41236 (n24792, n_15331, n24790);
  not g41237 (n_16541, n24791);
  not g41238 (n_16542, n24792);
  and g41239 (n24793, n_16541, n_16542);
  not g41240 (n_16543, n24793);
  and g41241 (n24794, \a[8] , n_16543);
  and g41242 (n24795, n_1106, n24793);
  not g41243 (n_16544, n24794);
  not g41244 (n_16545, n24795);
  and g41245 (n24796, n_16544, n_16545);
  not g41246 (n_16546, n24796);
  and g41247 (n24797, n24785, n_16546);
  and g41248 (n24798, n24377, n24549);
  not g41249 (n_16547, n24798);
  and g41250 (n24799, n_16334, n_16547);
  and g41251 (n24800, n9331, n22362);
  and g41252 (n24801, n8418, n22368);
  and g41253 (n24802, n8860, n22365);
  not g41254 (n_16548, n24801);
  not g41255 (n_16549, n24802);
  and g41256 (n24803, n_16548, n_16549);
  not g41257 (n_16550, n24800);
  and g41258 (n24804, n_16550, n24803);
  and g41259 (n24805, n_3428, n24804);
  and g41260 (n24806, n23320, n24804);
  not g41261 (n_16551, n24805);
  not g41262 (n_16552, n24806);
  and g41263 (n24807, n_16551, n_16552);
  not g41264 (n_16553, n24807);
  and g41265 (n24808, \a[8] , n_16553);
  and g41266 (n24809, n_1106, n24807);
  not g41267 (n_16554, n24808);
  not g41268 (n_16555, n24809);
  and g41269 (n24810, n_16554, n_16555);
  not g41270 (n_16556, n24810);
  and g41271 (n24811, n24799, n_16556);
  and g41272 (n24812, n9331, n22365);
  and g41273 (n24813, n8418, n22371);
  and g41274 (n24814, n8860, n22368);
  and g41280 (n24817, n8421, n_15351);
  not g41283 (n_16561, n24818);
  and g41284 (n24819, \a[8] , n_16561);
  not g41285 (n_16562, n24819);
  and g41286 (n24820, n_16561, n_16562);
  and g41287 (n24821, \a[8] , n_16562);
  not g41288 (n_16563, n24820);
  not g41289 (n_16564, n24821);
  and g41290 (n24822, n_16563, n_16564);
  not g41291 (n_16565, n24547);
  and g41292 (n24823, n24545, n_16565);
  not g41293 (n_16566, n24823);
  and g41294 (n24824, n_16331, n_16566);
  not g41295 (n_16567, n24822);
  and g41296 (n24825, n_16567, n24824);
  not g41297 (n_16568, n24825);
  and g41298 (n24826, n_16567, n_16568);
  and g41299 (n24827, n24824, n_16568);
  not g41300 (n_16569, n24826);
  not g41301 (n_16570, n24827);
  and g41302 (n24828, n_16569, n_16570);
  and g41303 (n24829, n9331, n22368);
  and g41304 (n24830, n8418, n22374);
  and g41305 (n24831, n8860, n22371);
  and g41311 (n24834, n8421, n23006);
  not g41314 (n_16575, n24835);
  and g41315 (n24836, \a[8] , n_16575);
  not g41316 (n_16576, n24836);
  and g41317 (n24837, n_16575, n_16576);
  and g41318 (n24838, \a[8] , n_16576);
  not g41319 (n_16577, n24837);
  not g41320 (n_16578, n24838);
  and g41321 (n24839, n_16577, n_16578);
  and g41322 (n24840, n_16324, n_16326);
  and g41323 (n24841, n_16325, n_16326);
  not g41324 (n_16579, n24840);
  not g41325 (n_16580, n24841);
  and g41326 (n24842, n_16579, n_16580);
  not g41327 (n_16581, n24839);
  not g41328 (n_16582, n24842);
  and g41329 (n24843, n_16581, n_16582);
  not g41330 (n_16583, n24843);
  and g41331 (n24844, n_16581, n_16583);
  and g41332 (n24845, n_16582, n_16583);
  not g41333 (n_16584, n24844);
  not g41334 (n_16585, n24845);
  and g41335 (n24846, n_16584, n_16585);
  and g41336 (n24847, n9331, n22371);
  and g41337 (n24848, n8418, n22377);
  and g41338 (n24849, n8860, n22374);
  and g41344 (n24852, n8421, n23025);
  not g41347 (n_16590, n24853);
  and g41348 (n24854, \a[8] , n_16590);
  not g41349 (n_16591, n24854);
  and g41350 (n24855, n_16590, n_16591);
  and g41351 (n24856, \a[8] , n_16591);
  not g41352 (n_16592, n24855);
  not g41353 (n_16593, n24856);
  and g41354 (n24857, n_16592, n_16593);
  and g41355 (n24858, n_16318, n_16320);
  and g41356 (n24859, n_16319, n_16320);
  not g41357 (n_16594, n24858);
  not g41358 (n_16595, n24859);
  and g41359 (n24860, n_16594, n_16595);
  not g41360 (n_16596, n24857);
  not g41361 (n_16597, n24860);
  and g41362 (n24861, n_16596, n_16597);
  not g41363 (n_16598, n24861);
  and g41364 (n24862, n_16596, n_16598);
  and g41365 (n24863, n_16597, n_16598);
  not g41366 (n_16599, n24862);
  not g41367 (n_16600, n24863);
  and g41368 (n24864, n_16599, n_16600);
  and g41369 (n24865, n24436, n24533);
  not g41370 (n_16601, n24865);
  and g41371 (n24866, n_16314, n_16601);
  and g41372 (n24867, n9331, n22374);
  and g41373 (n24868, n8418, n22380);
  and g41374 (n24869, n8860, n22377);
  not g41375 (n_16602, n24868);
  not g41376 (n_16603, n24869);
  and g41377 (n24870, n_16602, n_16603);
  not g41378 (n_16604, n24867);
  and g41379 (n24871, n_16604, n24870);
  and g41380 (n24872, n_3428, n24871);
  and g41381 (n24873, n_15064, n24871);
  not g41382 (n_16605, n24872);
  not g41383 (n_16606, n24873);
  and g41384 (n24874, n_16605, n_16606);
  not g41385 (n_16607, n24874);
  and g41386 (n24875, \a[8] , n_16607);
  and g41387 (n24876, n_1106, n24874);
  not g41388 (n_16608, n24875);
  not g41389 (n_16609, n24876);
  and g41390 (n24877, n_16608, n_16609);
  not g41391 (n_16610, n24877);
  and g41392 (n24878, n24866, n_16610);
  not g41393 (n_16611, n24531);
  and g41394 (n24879, n24529, n_16611);
  not g41395 (n_16612, n24879);
  and g41396 (n24880, n_16311, n_16612);
  and g41397 (n24881, n9331, n22377);
  and g41398 (n24882, n8418, n22384);
  and g41399 (n24883, n8860, n22380);
  not g41400 (n_16613, n24882);
  not g41401 (n_16614, n24883);
  and g41402 (n24884, n_16613, n_16614);
  not g41403 (n_16615, n24881);
  and g41404 (n24885, n_16615, n24884);
  and g41405 (n24886, n_3428, n24885);
  and g41406 (n24887, n22834, n24885);
  not g41407 (n_16616, n24886);
  not g41408 (n_16617, n24887);
  and g41409 (n24888, n_16616, n_16617);
  not g41410 (n_16618, n24888);
  and g41411 (n24889, \a[8] , n_16618);
  and g41412 (n24890, n_1106, n24888);
  not g41413 (n_16619, n24889);
  not g41414 (n_16620, n24890);
  and g41415 (n24891, n_16619, n_16620);
  not g41416 (n_16621, n24891);
  and g41417 (n24892, n24880, n_16621);
  and g41418 (n24893, n24468, n24527);
  not g41419 (n_16622, n24893);
  and g41420 (n24894, n_16307, n_16622);
  and g41421 (n24895, n9331, n22380);
  and g41422 (n24896, n8418, n22387);
  and g41423 (n24897, n8860, n22384);
  not g41424 (n_16623, n24896);
  not g41425 (n_16624, n24897);
  and g41426 (n24898, n_16623, n_16624);
  not g41427 (n_16625, n24895);
  and g41428 (n24899, n_16625, n24898);
  and g41429 (n24900, n_3428, n24899);
  and g41430 (n24901, n_14894, n24899);
  not g41431 (n_16626, n24900);
  not g41432 (n_16627, n24901);
  and g41433 (n24902, n_16626, n_16627);
  not g41434 (n_16628, n24902);
  and g41435 (n24903, \a[8] , n_16628);
  and g41436 (n24904, n_1106, n24902);
  not g41437 (n_16629, n24903);
  not g41438 (n_16630, n24904);
  and g41439 (n24905, n_16629, n_16630);
  not g41440 (n_16631, n24905);
  and g41441 (n24906, n24894, n_16631);
  and g41442 (n24907, n9331, n22384);
  and g41443 (n24908, n8418, n22390);
  and g41444 (n24909, n8860, n22387);
  and g41450 (n24912, n8421, n22806);
  not g41453 (n_16636, n24913);
  and g41454 (n24914, \a[8] , n_16636);
  not g41455 (n_16637, n24914);
  and g41456 (n24915, n_16636, n_16637);
  and g41457 (n24916, \a[8] , n_16637);
  not g41458 (n_16638, n24915);
  not g41459 (n_16639, n24916);
  and g41460 (n24917, n_16638, n_16639);
  not g41461 (n_16640, n24525);
  and g41462 (n24918, n24523, n_16640);
  not g41463 (n_16641, n24918);
  and g41464 (n24919, n_16304, n_16641);
  not g41465 (n_16642, n24917);
  and g41466 (n24920, n_16642, n24919);
  not g41467 (n_16643, n24920);
  and g41468 (n24921, n_16642, n_16643);
  and g41469 (n24922, n24919, n_16643);
  not g41470 (n_16644, n24921);
  not g41471 (n_16645, n24922);
  and g41472 (n24923, n_16644, n_16645);
  and g41473 (n24924, n_16297, n_16299);
  and g41474 (n24925, n_16298, n_16299);
  not g41475 (n_16646, n24924);
  not g41476 (n_16647, n24925);
  and g41477 (n24926, n_16646, n_16647);
  and g41478 (n24927, n9331, n22387);
  and g41479 (n24928, n8418, n22393);
  and g41480 (n24929, n8860, n22390);
  not g41481 (n_16648, n24928);
  not g41482 (n_16649, n24929);
  and g41483 (n24930, n_16648, n_16649);
  not g41484 (n_16650, n24927);
  and g41485 (n24931, n_16650, n24930);
  and g41486 (n24932, n_3428, n24931);
  and g41487 (n24933, n_14920, n24931);
  not g41488 (n_16651, n24932);
  not g41489 (n_16652, n24933);
  and g41490 (n24934, n_16651, n_16652);
  not g41491 (n_16653, n24934);
  and g41492 (n24935, \a[8] , n_16653);
  and g41493 (n24936, n_1106, n24934);
  not g41494 (n_16654, n24935);
  not g41495 (n_16655, n24936);
  and g41496 (n24937, n_16654, n_16655);
  not g41497 (n_16656, n24926);
  not g41498 (n_16657, n24937);
  and g41499 (n24938, n_16656, n_16657);
  and g41500 (n24939, n9331, n22390);
  and g41501 (n24940, n8418, n22396);
  and g41502 (n24941, n8860, n22393);
  and g41508 (n24944, n8421, n22649);
  not g41511 (n_16662, n24945);
  and g41512 (n24946, \a[8] , n_16662);
  not g41513 (n_16663, n24946);
  and g41514 (n24947, n_16662, n_16663);
  and g41515 (n24948, \a[8] , n_16663);
  not g41516 (n_16664, n24947);
  not g41517 (n_16665, n24948);
  and g41518 (n24949, n_16664, n_16665);
  not g41519 (n_16666, n24494);
  and g41520 (n24950, n_16666, n24505);
  not g41521 (n_16667, n24506);
  not g41522 (n_16668, n24950);
  and g41523 (n24951, n_16667, n_16668);
  not g41524 (n_16669, n24949);
  and g41525 (n24952, n_16669, n24951);
  not g41526 (n_16670, n24952);
  and g41527 (n24953, n_16669, n_16670);
  and g41528 (n24954, n24951, n_16670);
  not g41529 (n_16671, n24953);
  not g41530 (n_16672, n24954);
  and g41531 (n24955, n_16671, n_16672);
  not g41532 (n_16673, n24493);
  and g41533 (n24956, n24491, n_16673);
  not g41534 (n_16674, n24956);
  and g41535 (n24957, n_16666, n_16674);
  and g41536 (n24958, n9331, n22393);
  and g41537 (n24959, n8418, n22399);
  and g41538 (n24960, n8860, n22396);
  not g41539 (n_16675, n24959);
  not g41540 (n_16676, n24960);
  and g41541 (n24961, n_16675, n_16676);
  not g41542 (n_16677, n24958);
  and g41543 (n24962, n_16677, n24961);
  and g41544 (n24963, n_3428, n24962);
  and g41545 (n24964, n_14773, n24962);
  not g41546 (n_16678, n24963);
  not g41547 (n_16679, n24964);
  and g41548 (n24965, n_16678, n_16679);
  not g41549 (n_16680, n24965);
  and g41550 (n24966, \a[8] , n_16680);
  and g41551 (n24967, n_1106, n24965);
  not g41552 (n_16681, n24966);
  not g41553 (n_16682, n24967);
  and g41554 (n24968, n_16681, n_16682);
  not g41555 (n_16683, n24968);
  and g41556 (n24969, n24957, n_16683);
  and g41557 (n24970, n8860, n_14508);
  and g41558 (n24971, n9331, n22402);
  not g41559 (n_16684, n24970);
  not g41560 (n_16685, n24971);
  and g41561 (n24972, n_16684, n_16685);
  and g41562 (n24973, n8421, n_14720);
  not g41563 (n_16686, n24973);
  and g41564 (n24974, n24972, n_16686);
  not g41565 (n_16687, n24974);
  and g41566 (n24975, \a[8] , n_16687);
  not g41567 (n_16688, n24975);
  and g41568 (n24976, \a[8] , n_16688);
  and g41569 (n24977, n_16687, n_16688);
  not g41570 (n_16689, n24976);
  not g41571 (n_16690, n24977);
  and g41572 (n24978, n_16689, n_16690);
  and g41573 (n24979, n_3427, n_14508);
  not g41574 (n_16691, n24979);
  and g41575 (n24980, \a[8] , n_16691);
  not g41576 (n_16692, n24978);
  and g41577 (n24981, n_16692, n24980);
  and g41578 (n24982, n9331, n22399);
  and g41579 (n24983, n8418, n_14508);
  and g41580 (n24984, n8860, n22402);
  not g41581 (n_16693, n24983);
  not g41582 (n_16694, n24984);
  and g41583 (n24985, n_16693, n_16694);
  not g41584 (n_16695, n24982);
  and g41585 (n24986, n_16695, n24985);
  and g41586 (n24987, n_3428, n24986);
  and g41587 (n24988, n22625, n24986);
  not g41588 (n_16696, n24987);
  not g41589 (n_16697, n24988);
  and g41590 (n24989, n_16696, n_16697);
  not g41591 (n_16698, n24989);
  and g41592 (n24990, \a[8] , n_16698);
  and g41593 (n24991, n_1106, n24989);
  not g41594 (n_16699, n24990);
  not g41595 (n_16700, n24991);
  and g41596 (n24992, n_16699, n_16700);
  not g41597 (n_16701, n24992);
  and g41598 (n24993, n24981, n_16701);
  and g41599 (n24994, n24492, n24993);
  not g41600 (n_16702, n24994);
  and g41601 (n24995, n24993, n_16702);
  and g41602 (n24996, n24492, n_16702);
  not g41603 (n_16703, n24995);
  not g41604 (n_16704, n24996);
  and g41605 (n24997, n_16703, n_16704);
  and g41606 (n24998, n9331, n22396);
  and g41607 (n24999, n8418, n22402);
  and g41608 (n25000, n8860, n22399);
  and g41614 (n25003, n8421, n22595);
  not g41617 (n_16709, n25004);
  and g41618 (n25005, \a[8] , n_16709);
  not g41619 (n_16710, n25005);
  and g41620 (n25006, \a[8] , n_16710);
  and g41621 (n25007, n_16709, n_16710);
  not g41622 (n_16711, n25006);
  not g41623 (n_16712, n25007);
  and g41624 (n25008, n_16711, n_16712);
  not g41625 (n_16713, n24997);
  not g41626 (n_16714, n25008);
  and g41627 (n25009, n_16713, n_16714);
  not g41628 (n_16715, n25009);
  and g41629 (n25010, n_16702, n_16715);
  not g41630 (n_16716, n24957);
  and g41631 (n25011, n_16716, n24968);
  not g41632 (n_16717, n24969);
  not g41633 (n_16718, n25011);
  and g41634 (n25012, n_16717, n_16718);
  not g41635 (n_16719, n25010);
  and g41636 (n25013, n_16719, n25012);
  not g41637 (n_16720, n25013);
  and g41638 (n25014, n_16717, n_16720);
  not g41639 (n_16721, n24955);
  not g41640 (n_16722, n25014);
  and g41641 (n25015, n_16721, n_16722);
  not g41642 (n_16723, n25015);
  and g41643 (n25016, n_16670, n_16723);
  and g41644 (n25017, n24926, n24937);
  not g41645 (n_16724, n24938);
  not g41646 (n_16725, n25017);
  and g41647 (n25018, n_16724, n_16725);
  not g41648 (n_16726, n25016);
  and g41649 (n25019, n_16726, n25018);
  not g41650 (n_16727, n25019);
  and g41651 (n25020, n_16724, n_16727);
  not g41652 (n_16728, n24923);
  not g41653 (n_16729, n25020);
  and g41654 (n25021, n_16728, n_16729);
  not g41655 (n_16730, n25021);
  and g41656 (n25022, n_16643, n_16730);
  not g41657 (n_16731, n24906);
  and g41658 (n25023, n24894, n_16731);
  and g41659 (n25024, n_16631, n_16731);
  not g41660 (n_16732, n25023);
  not g41661 (n_16733, n25024);
  and g41662 (n25025, n_16732, n_16733);
  not g41663 (n_16734, n25022);
  not g41664 (n_16735, n25025);
  and g41665 (n25026, n_16734, n_16735);
  not g41666 (n_16736, n25026);
  and g41667 (n25027, n_16731, n_16736);
  not g41668 (n_16737, n24892);
  and g41669 (n25028, n24880, n_16737);
  and g41670 (n25029, n_16621, n_16737);
  not g41671 (n_16738, n25028);
  not g41672 (n_16739, n25029);
  and g41673 (n25030, n_16738, n_16739);
  not g41674 (n_16740, n25027);
  not g41675 (n_16741, n25030);
  and g41676 (n25031, n_16740, n_16741);
  not g41677 (n_16742, n25031);
  and g41678 (n25032, n_16737, n_16742);
  not g41679 (n_16743, n24866);
  and g41680 (n25033, n_16743, n24877);
  not g41681 (n_16744, n24878);
  not g41682 (n_16745, n25033);
  and g41683 (n25034, n_16744, n_16745);
  not g41684 (n_16746, n25032);
  and g41685 (n25035, n_16746, n25034);
  not g41686 (n_16747, n25035);
  and g41687 (n25036, n_16744, n_16747);
  not g41688 (n_16748, n24864);
  not g41689 (n_16749, n25036);
  and g41690 (n25037, n_16748, n_16749);
  not g41691 (n_16750, n25037);
  and g41692 (n25038, n_16598, n_16750);
  not g41693 (n_16751, n24846);
  not g41694 (n_16752, n25038);
  and g41695 (n25039, n_16751, n_16752);
  not g41696 (n_16753, n25039);
  and g41697 (n25040, n_16583, n_16753);
  not g41698 (n_16754, n24828);
  not g41699 (n_16755, n25040);
  and g41700 (n25041, n_16754, n_16755);
  not g41701 (n_16756, n25041);
  and g41702 (n25042, n_16568, n_16756);
  not g41703 (n_16757, n24811);
  and g41704 (n25043, n24799, n_16757);
  and g41705 (n25044, n_16556, n_16757);
  not g41706 (n_16758, n25043);
  not g41707 (n_16759, n25044);
  and g41708 (n25045, n_16758, n_16759);
  not g41709 (n_16760, n25042);
  not g41710 (n_16761, n25045);
  and g41711 (n25046, n_16760, n_16761);
  not g41712 (n_16762, n25046);
  and g41713 (n25047, n_16757, n_16762);
  not g41714 (n_16763, n24797);
  and g41715 (n25048, n24785, n_16763);
  and g41716 (n25049, n_16546, n_16763);
  not g41717 (n_16764, n25048);
  not g41718 (n_16765, n25049);
  and g41719 (n25050, n_16764, n_16765);
  not g41720 (n_16766, n25047);
  not g41721 (n_16767, n25050);
  and g41722 (n25051, n_16766, n_16767);
  not g41723 (n_16768, n25051);
  and g41724 (n25052, n_16763, n_16768);
  not g41725 (n_16769, n24771);
  and g41726 (n25053, n_16769, n24782);
  not g41727 (n_16770, n24783);
  not g41728 (n_16771, n25053);
  and g41729 (n25054, n_16770, n_16771);
  not g41730 (n_16772, n25052);
  and g41731 (n25055, n_16772, n25054);
  not g41732 (n_16773, n25055);
  and g41733 (n25056, n_16770, n_16773);
  not g41734 (n_16774, n24769);
  not g41735 (n_16775, n25056);
  and g41736 (n25057, n_16774, n_16775);
  not g41737 (n_16776, n25057);
  and g41738 (n25058, n_16524, n_16776);
  not g41739 (n_16777, n24751);
  not g41740 (n_16778, n25058);
  and g41741 (n25059, n_16777, n_16778);
  not g41742 (n_16779, n25059);
  and g41743 (n25060, n_16509, n_16779);
  not g41744 (n_16780, n24733);
  not g41745 (n_16781, n25060);
  and g41746 (n25061, n_16780, n_16781);
  not g41747 (n_16782, n25061);
  and g41748 (n25062, n_16494, n_16782);
  not g41749 (n_16783, n24716);
  and g41750 (n25063, n24704, n_16783);
  and g41751 (n25064, n_16482, n_16783);
  not g41752 (n_16784, n25063);
  not g41753 (n_16785, n25064);
  and g41754 (n25065, n_16784, n_16785);
  not g41755 (n_16786, n25062);
  not g41756 (n_16787, n25065);
  and g41757 (n25066, n_16786, n_16787);
  not g41758 (n_16788, n25066);
  and g41759 (n25067, n_16783, n_16788);
  not g41760 (n_16789, n24702);
  and g41761 (n25068, n24690, n_16789);
  and g41762 (n25069, n_16472, n_16789);
  not g41763 (n_16790, n25068);
  not g41764 (n_16791, n25069);
  and g41765 (n25070, n_16790, n_16791);
  not g41766 (n_16792, n25067);
  not g41767 (n_16793, n25070);
  and g41768 (n25071, n_16792, n_16793);
  not g41769 (n_16794, n25071);
  and g41770 (n25072, n_16789, n_16794);
  not g41771 (n_16795, n24676);
  and g41772 (n25073, n_16795, n24687);
  not g41773 (n_16796, n24688);
  not g41774 (n_16797, n25073);
  and g41775 (n25074, n_16796, n_16797);
  not g41776 (n_16798, n25072);
  and g41777 (n25075, n_16798, n25074);
  not g41778 (n_16799, n25075);
  and g41779 (n25076, n_16796, n_16799);
  not g41780 (n_16800, n24674);
  not g41781 (n_16801, n25076);
  and g41782 (n25077, n_16800, n_16801);
  not g41783 (n_16802, n25077);
  and g41784 (n25078, n_16450, n_16802);
  not g41785 (n_16803, n24656);
  not g41786 (n_16804, n25078);
  and g41787 (n25079, n_16803, n_16804);
  not g41788 (n_16805, n25079);
  and g41789 (n25080, n_16435, n_16805);
  not g41790 (n_16806, n24639);
  and g41791 (n25081, n24624, n_16806);
  and g41792 (n25082, n_16423, n_16806);
  not g41793 (n_16807, n25081);
  not g41794 (n_16808, n25082);
  and g41795 (n25083, n_16807, n_16808);
  not g41796 (n_16809, n25080);
  not g41797 (n_16810, n25083);
  and g41798 (n25084, n_16809, n_16810);
  not g41799 (n_16811, n25084);
  and g41800 (n25085, n_16806, n_16811);
  not g41801 (n_16812, n24622);
  and g41802 (n25086, n24607, n_16812);
  and g41803 (n25087, n_16411, n_16812);
  not g41804 (n_16813, n25086);
  not g41805 (n_16814, n25087);
  and g41806 (n25088, n_16813, n_16814);
  not g41807 (n_16815, n25085);
  not g41808 (n_16816, n25088);
  and g41809 (n25089, n_16815, n_16816);
  not g41810 (n_16817, n25089);
  and g41811 (n25090, n_16812, n_16817);
  not g41812 (n_16818, n24605);
  and g41813 (n25091, n24591, n_16818);
  and g41814 (n25092, n_16399, n_16818);
  not g41815 (n_16819, n25091);
  not g41816 (n_16820, n25092);
  and g41817 (n25093, n_16819, n_16820);
  not g41818 (n_16821, n25090);
  not g41819 (n_16822, n25093);
  and g41820 (n25094, n_16821, n_16822);
  not g41821 (n_16823, n25094);
  and g41822 (n25095, n_16818, n_16823);
  and g41823 (n25096, n7983, n22329);
  and g41824 (n25097, n7291, n22335);
  and g41825 (n25098, n7632, n22332);
  not g41831 (n_16827, n24633);
  and g41832 (n25101, n7294, n_16827);
  not g41835 (n_16829, n25102);
  and g41836 (n25103, \a[11] , n_16829);
  not g41837 (n_16830, n25103);
  and g41838 (n25104, n_16829, n_16830);
  and g41839 (n25105, \a[11] , n_16830);
  not g41840 (n_16831, n25104);
  not g41841 (n_16832, n25105);
  and g41842 (n25106, n_16831, n_16832);
  and g41843 (n25107, n_15997, n_16002);
  and g41844 (n25108, n6233, n22347);
  and g41845 (n25109, n5663, n22353);
  and g41846 (n25110, n5939, n22350);
  and g41852 (n25113, n5666, n_16069);
  not g41855 (n_16837, n25114);
  and g41856 (n25115, \a[17] , n_16837);
  not g41857 (n_16838, n25115);
  and g41858 (n25116, n_16837, n_16838);
  and g41859 (n25117, \a[17] , n_16838);
  not g41860 (n_16839, n25116);
  not g41861 (n_16840, n25117);
  and g41862 (n25118, n_16839, n_16840);
  and g41863 (n25119, n_15968, n_15973);
  and g41864 (n25120, n4694, n22365);
  and g41865 (n25121, n4533, n22371);
  and g41866 (n25122, n4604, n22368);
  and g41872 (n25125, n4536, n_15351);
  not g41875 (n_16845, n25126);
  and g41876 (n25127, \a[23] , n_16845);
  not g41877 (n_16846, n25127);
  and g41878 (n25128, n_16845, n_16846);
  and g41879 (n25129, \a[23] , n_16846);
  not g41880 (n_16847, n25128);
  not g41881 (n_16848, n25129);
  and g41882 (n25130, n_16847, n_16848);
  and g41883 (n25131, n_15942, n_15947);
  and g41884 (n25132, n3457, n22384);
  and g41885 (n25133, n3542, n22390);
  and g41886 (n25134, n3606, n22387);
  and g41892 (n25137, n3368, n22806);
  not g41895 (n_16853, n25138);
  and g41896 (n25139, \a[29] , n_16853);
  not g41897 (n_16854, n25139);
  and g41898 (n25140, n_16853, n_16854);
  and g41899 (n25141, \a[29] , n_16854);
  not g41900 (n_16855, n25140);
  not g41901 (n_16856, n25141);
  and g41902 (n25142, n_16855, n_16856);
  and g41903 (n25143, n_15916, n_15921);
  and g41918 (n25158, n3020, n22393);
  and g41919 (n25159, n3028, n22396);
  and g41920 (n25160, n3023, n22399);
  and g41921 (n25161, n75, n22671);
  not g41929 (n_16861, n25157);
  not g41930 (n_16862, n25164);
  and g41931 (n25165, n_16861, n_16862);
  not g41932 (n_16863, n25165);
  and g41933 (n25166, n_16861, n_16863);
  and g41934 (n25167, n_16862, n_16863);
  not g41935 (n_16864, n25166);
  not g41936 (n_16865, n25167);
  and g41937 (n25168, n_16864, n_16865);
  not g41938 (n_16866, n25143);
  not g41939 (n_16867, n25168);
  and g41940 (n25169, n_16866, n_16867);
  not g41941 (n_16868, n25169);
  and g41942 (n25170, n_16866, n_16868);
  and g41943 (n25171, n_16867, n_16868);
  not g41944 (n_16869, n25170);
  not g41945 (n_16870, n25171);
  and g41946 (n25172, n_16869, n_16870);
  not g41947 (n_16871, n25142);
  not g41948 (n_16872, n25172);
  and g41949 (n25173, n_16871, n_16872);
  not g41950 (n_16873, n25173);
  and g41951 (n25174, n_16871, n_16873);
  and g41952 (n25175, n_16872, n_16873);
  not g41953 (n_16874, n25174);
  not g41954 (n_16875, n25175);
  and g41955 (n25176, n_16874, n_16875);
  and g41956 (n25177, n_15926, n_15932);
  and g41957 (n25178, n25176, n25177);
  not g41958 (n_16876, n25176);
  not g41959 (n_16877, n25177);
  and g41960 (n25179, n_16876, n_16877);
  not g41961 (n_16878, n25178);
  not g41962 (n_16879, n25179);
  and g41963 (n25180, n_16878, n_16879);
  and g41964 (n25181, n3884, n22374);
  and g41965 (n25182, n3967, n22380);
  and g41966 (n25183, n4046, n22377);
  not g41967 (n_16880, n25182);
  not g41968 (n_16881, n25183);
  and g41969 (n25184, n_16880, n_16881);
  not g41970 (n_16882, n25181);
  and g41971 (n25185, n_16882, n25184);
  and g41972 (n25186, n_750, n25185);
  and g41973 (n25187, n_15064, n25185);
  not g41974 (n_16883, n25186);
  not g41975 (n_16884, n25187);
  and g41976 (n25188, n_16883, n_16884);
  not g41977 (n_16885, n25188);
  and g41978 (n25189, \a[26] , n_16885);
  and g41979 (n25190, n_33, n25188);
  not g41980 (n_16886, n25189);
  not g41981 (n_16887, n25190);
  and g41982 (n25191, n_16886, n_16887);
  not g41983 (n_16888, n25191);
  and g41984 (n25192, n25180, n_16888);
  not g41985 (n_16889, n25192);
  and g41986 (n25193, n25180, n_16889);
  and g41987 (n25194, n_16888, n_16889);
  not g41988 (n_16890, n25193);
  not g41989 (n_16891, n25194);
  and g41990 (n25195, n_16890, n_16891);
  not g41991 (n_16892, n25131);
  not g41992 (n_16893, n25195);
  and g41993 (n25196, n_16892, n_16893);
  not g41994 (n_16894, n25196);
  and g41995 (n25197, n_16892, n_16894);
  and g41996 (n25198, n_16893, n_16894);
  not g41997 (n_16895, n25197);
  not g41998 (n_16896, n25198);
  and g41999 (n25199, n_16895, n_16896);
  not g42000 (n_16897, n25130);
  not g42001 (n_16898, n25199);
  and g42002 (n25200, n_16897, n_16898);
  not g42003 (n_16899, n25200);
  and g42004 (n25201, n_16897, n_16899);
  and g42005 (n25202, n_16898, n_16899);
  not g42006 (n_16900, n25201);
  not g42007 (n_16901, n25202);
  and g42008 (n25203, n_16900, n_16901);
  and g42009 (n25204, n_15952, n_15958);
  and g42010 (n25205, n25203, n25204);
  not g42011 (n_16902, n25203);
  not g42012 (n_16903, n25204);
  and g42013 (n25206, n_16902, n_16903);
  not g42014 (n_16904, n25205);
  not g42015 (n_16905, n25206);
  and g42016 (n25207, n_16904, n_16905);
  and g42017 (n25208, n5496, n22356);
  and g42018 (n25209, n4935, n22362);
  and g42019 (n25210, n5407, n22359);
  not g42020 (n_16906, n25209);
  not g42021 (n_16907, n25210);
  and g42022 (n25211, n_16906, n_16907);
  not g42023 (n_16908, n25208);
  and g42024 (n25212, n_16908, n25211);
  and g42025 (n25213, n_1011, n25212);
  and g42026 (n25214, n23345, n25212);
  not g42027 (n_16909, n25213);
  not g42028 (n_16910, n25214);
  and g42029 (n25215, n_16909, n_16910);
  not g42030 (n_16911, n25215);
  and g42031 (n25216, \a[20] , n_16911);
  and g42032 (n25217, n_435, n25215);
  not g42033 (n_16912, n25216);
  not g42034 (n_16913, n25217);
  and g42035 (n25218, n_16912, n_16913);
  not g42036 (n_16914, n25218);
  and g42037 (n25219, n25207, n_16914);
  not g42038 (n_16915, n25219);
  and g42039 (n25220, n25207, n_16915);
  and g42040 (n25221, n_16914, n_16915);
  not g42041 (n_16916, n25220);
  not g42042 (n_16917, n25221);
  and g42043 (n25222, n_16916, n_16917);
  not g42044 (n_16918, n25119);
  not g42045 (n_16919, n25222);
  and g42046 (n25223, n_16918, n_16919);
  not g42047 (n_16920, n25223);
  and g42048 (n25224, n_16918, n_16920);
  and g42049 (n25225, n_16919, n_16920);
  not g42050 (n_16921, n25224);
  not g42051 (n_16922, n25225);
  and g42052 (n25226, n_16921, n_16922);
  not g42053 (n_16923, n25118);
  not g42054 (n_16924, n25226);
  and g42055 (n25227, n_16923, n_16924);
  not g42056 (n_16925, n25227);
  and g42057 (n25228, n_16923, n_16925);
  and g42058 (n25229, n_16924, n_16925);
  not g42059 (n_16926, n25228);
  not g42060 (n_16927, n25229);
  and g42061 (n25230, n_16926, n_16927);
  and g42062 (n25231, n_15978, n_15984);
  and g42063 (n25232, n25230, n25231);
  not g42064 (n_16928, n25230);
  not g42065 (n_16929, n25231);
  and g42066 (n25233, n_16928, n_16929);
  not g42067 (n_16930, n25232);
  not g42068 (n_16931, n25233);
  and g42069 (n25234, n_16930, n_16931);
  and g42070 (n25235, n7101, n22338);
  and g42071 (n25236, n6402, n22344);
  and g42072 (n25237, n6951, n22341);
  not g42073 (n_16932, n25236);
  not g42074 (n_16933, n25237);
  and g42075 (n25238, n_16932, n_16933);
  not g42076 (n_16934, n25235);
  and g42077 (n25239, n_16934, n25238);
  and g42078 (n25240, n_1885, n25239);
  and g42079 (n25241, n24188, n25239);
  not g42080 (n_16935, n25240);
  not g42081 (n_16936, n25241);
  and g42082 (n25242, n_16935, n_16936);
  not g42083 (n_16937, n25242);
  and g42084 (n25243, \a[14] , n_16937);
  and g42085 (n25244, n_652, n25242);
  not g42086 (n_16938, n25243);
  not g42087 (n_16939, n25244);
  and g42088 (n25245, n_16938, n_16939);
  not g42089 (n_16940, n25245);
  and g42090 (n25246, n25234, n_16940);
  not g42091 (n_16941, n25246);
  and g42092 (n25247, n25234, n_16941);
  and g42093 (n25248, n_16940, n_16941);
  not g42094 (n_16942, n25247);
  not g42095 (n_16943, n25248);
  and g42096 (n25249, n_16942, n_16943);
  not g42097 (n_16944, n25107);
  not g42098 (n_16945, n25249);
  and g42099 (n25250, n_16944, n_16945);
  not g42100 (n_16946, n25250);
  and g42101 (n25251, n_16944, n_16946);
  and g42102 (n25252, n_16945, n_16946);
  not g42103 (n_16947, n25251);
  not g42104 (n_16948, n25252);
  and g42105 (n25253, n_16947, n_16948);
  not g42106 (n_16949, n25106);
  not g42107 (n_16950, n25253);
  and g42108 (n25254, n_16949, n_16950);
  not g42109 (n_16951, n25254);
  and g42110 (n25255, n_16949, n_16951);
  and g42111 (n25256, n_16950, n_16951);
  not g42112 (n_16952, n25255);
  not g42113 (n_16953, n25256);
  and g42114 (n25257, n_16952, n_16953);
  and g42115 (n25258, n_16007, n_16387);
  and g42116 (n25259, n25257, n25258);
  not g42117 (n_16954, n25257);
  not g42118 (n_16955, n25258);
  and g42119 (n25260, n_16954, n_16955);
  not g42120 (n_16956, n25259);
  not g42121 (n_16957, n25260);
  and g42122 (n25261, n_16956, n_16957);
  and g42123 (n25262, n9331, n22320);
  and g42124 (n25263, n8418, n22326);
  and g42125 (n25264, n8860, n22323);
  not g42126 (n_16958, n25263);
  not g42127 (n_16959, n25264);
  and g42128 (n25265, n_16958, n_16959);
  not g42129 (n_16960, n25262);
  and g42130 (n25266, n_16960, n25265);
  and g42131 (n25267, n_3428, n25266);
  and g42132 (n25268, n_14636, n_14639);
  and g42133 (n25269, n_14637, n22512);
  not g42134 (n_16961, n25268);
  not g42135 (n_16962, n25269);
  and g42136 (n25270, n_16961, n_16962);
  and g42137 (n25271, n25266, n25270);
  not g42138 (n_16963, n25267);
  not g42139 (n_16964, n25271);
  and g42140 (n25272, n_16963, n_16964);
  not g42141 (n_16965, n25272);
  and g42142 (n25273, \a[8] , n_16965);
  and g42143 (n25274, n_1106, n25272);
  not g42144 (n_16966, n25273);
  not g42145 (n_16967, n25274);
  and g42146 (n25275, n_16966, n_16967);
  not g42147 (n_16968, n25275);
  and g42148 (n25276, n25261, n_16968);
  not g42149 (n_16969, n25276);
  and g42150 (n25277, n25261, n_16969);
  and g42151 (n25278, n_16968, n_16969);
  not g42152 (n_16970, n25277);
  not g42153 (n_16971, n25278);
  and g42154 (n25279, n_16970, n_16971);
  not g42155 (n_16972, n25095);
  not g42156 (n_16973, n25279);
  and g42157 (n25280, n_16972, n_16973);
  not g42158 (n_16974, n25280);
  and g42159 (n25281, n_16972, n_16974);
  and g42160 (n25282, n_16973, n_16974);
  not g42161 (n_16975, n25281);
  not g42162 (n_16976, n25282);
  and g42163 (n25283, n_16975, n_16976);
  not g42164 (n_16977, n22535);
  not g42165 (n_16978, n25283);
  and g42166 (n25284, n_16977, n_16978);
  not g42167 (n_16979, n25284);
  and g42168 (n25285, n_16977, n_16979);
  and g42169 (n25286, n_16978, n_16979);
  not g42170 (n_16980, n25285);
  not g42171 (n_16981, n25286);
  and g42172 (n25287, n_16980, n_16981);
  and g42173 (n25288, n71, n22315);
  and g42174 (n25289, n9867, n22320);
  and g42175 (n25290, n10434, n22312);
  not g42181 (n_16985, n22519);
  and g42182 (n25293, n22516, n_16985);
  not g42183 (n_16986, n25293);
  and g42184 (n25294, n_14649, n_16986);
  and g42185 (n25295, n9870, n25294);
  not g42188 (n_16988, n25296);
  and g42189 (n25297, \a[5] , n_16988);
  not g42190 (n_16989, n25297);
  and g42191 (n25298, n_16988, n_16989);
  and g42192 (n25299, \a[5] , n_16989);
  not g42193 (n_16990, n25298);
  not g42194 (n_16991, n25299);
  and g42195 (n25300, n_16990, n_16991);
  and g42196 (n25301, n_16821, n_16823);
  and g42197 (n25302, n_16822, n_16823);
  not g42198 (n_16992, n25301);
  not g42199 (n_16993, n25302);
  and g42200 (n25303, n_16992, n_16993);
  not g42201 (n_16994, n25300);
  not g42202 (n_16995, n25303);
  and g42203 (n25304, n_16994, n_16995);
  not g42204 (n_16996, n25304);
  and g42205 (n25305, n_16994, n_16996);
  and g42206 (n25306, n_16995, n_16996);
  not g42207 (n_16997, n25305);
  not g42208 (n_16998, n25306);
  and g42209 (n25307, n_16997, n_16998);
  and g42210 (n25308, n71, n22312);
  and g42211 (n25309, n9867, n22323);
  and g42212 (n25310, n10434, n22320);
  and g42218 (n25313, n_14641, n_14644);
  and g42219 (n25314, n_14642, n22516);
  not g42220 (n_17002, n25313);
  not g42221 (n_17003, n25314);
  and g42222 (n25315, n_17002, n_17003);
  not g42223 (n_17004, n25315);
  and g42224 (n25316, n9870, n_17004);
  not g42227 (n_17006, n25317);
  and g42228 (n25318, \a[5] , n_17006);
  not g42229 (n_17007, n25318);
  and g42230 (n25319, n_17006, n_17007);
  and g42231 (n25320, \a[5] , n_17007);
  not g42232 (n_17008, n25319);
  not g42233 (n_17009, n25320);
  and g42234 (n25321, n_17008, n_17009);
  and g42235 (n25322, n_16815, n_16817);
  and g42236 (n25323, n_16816, n_16817);
  not g42237 (n_17010, n25322);
  not g42238 (n_17011, n25323);
  and g42239 (n25324, n_17010, n_17011);
  not g42240 (n_17012, n25321);
  not g42241 (n_17013, n25324);
  and g42242 (n25325, n_17012, n_17013);
  not g42243 (n_17014, n25325);
  and g42244 (n25326, n_17012, n_17014);
  and g42245 (n25327, n_17013, n_17014);
  not g42246 (n_17015, n25326);
  not g42247 (n_17016, n25327);
  and g42248 (n25328, n_17015, n_17016);
  and g42249 (n25329, n71, n22320);
  and g42250 (n25330, n9867, n22326);
  and g42251 (n25331, n10434, n22323);
  not g42257 (n_17020, n25270);
  and g42258 (n25334, n9870, n_17020);
  not g42261 (n_17022, n25335);
  and g42262 (n25336, \a[5] , n_17022);
  not g42263 (n_17023, n25336);
  and g42264 (n25337, n_17022, n_17023);
  and g42265 (n25338, \a[5] , n_17023);
  not g42266 (n_17024, n25337);
  not g42267 (n_17025, n25338);
  and g42268 (n25339, n_17024, n_17025);
  and g42269 (n25340, n_16809, n_16811);
  and g42270 (n25341, n_16810, n_16811);
  not g42271 (n_17026, n25340);
  not g42272 (n_17027, n25341);
  and g42273 (n25342, n_17026, n_17027);
  not g42274 (n_17028, n25339);
  not g42275 (n_17029, n25342);
  and g42276 (n25343, n_17028, n_17029);
  not g42277 (n_17030, n25343);
  and g42278 (n25344, n_17028, n_17030);
  and g42279 (n25345, n_17029, n_17030);
  not g42280 (n_17031, n25344);
  not g42281 (n_17032, n25345);
  and g42282 (n25346, n_17031, n_17032);
  and g42283 (n25347, n24656, n25078);
  not g42284 (n_17033, n25347);
  and g42285 (n25348, n_16805, n_17033);
  and g42286 (n25349, n71, n22323);
  and g42287 (n25350, n9867, n22329);
  and g42288 (n25351, n10434, n22326);
  not g42289 (n_17034, n25350);
  not g42290 (n_17035, n25351);
  and g42291 (n25352, n_17034, n_17035);
  not g42292 (n_17036, n25349);
  and g42293 (n25353, n_17036, n25352);
  and g42294 (n25354, n_4684, n25353);
  and g42295 (n25355, n_16393, n25353);
  not g42296 (n_17037, n25354);
  not g42297 (n_17038, n25355);
  and g42298 (n25356, n_17037, n_17038);
  not g42299 (n_17039, n25356);
  and g42300 (n25357, \a[5] , n_17039);
  and g42301 (n25358, n_3, n25356);
  not g42302 (n_17040, n25357);
  not g42303 (n_17041, n25358);
  and g42304 (n25359, n_17040, n_17041);
  not g42305 (n_17042, n25359);
  and g42306 (n25360, n25348, n_17042);
  and g42307 (n25361, n24674, n25076);
  not g42308 (n_17043, n25361);
  and g42309 (n25362, n_16802, n_17043);
  and g42310 (n25363, n71, n22326);
  and g42311 (n25364, n9867, n22332);
  and g42312 (n25365, n10434, n22329);
  not g42313 (n_17044, n25364);
  not g42314 (n_17045, n25365);
  and g42315 (n25366, n_17044, n_17045);
  not g42316 (n_17046, n25363);
  and g42317 (n25367, n_17046, n25366);
  and g42318 (n25368, n_4684, n25367);
  and g42319 (n25369, n24616, n25367);
  not g42320 (n_17047, n25368);
  not g42321 (n_17048, n25369);
  and g42322 (n25370, n_17047, n_17048);
  not g42323 (n_17049, n25370);
  and g42324 (n25371, \a[5] , n_17049);
  and g42325 (n25372, n_3, n25370);
  not g42326 (n_17050, n25371);
  not g42327 (n_17051, n25372);
  and g42328 (n25373, n_17050, n_17051);
  not g42329 (n_17052, n25373);
  and g42330 (n25374, n25362, n_17052);
  and g42331 (n25375, n71, n22329);
  and g42332 (n25376, n9867, n22335);
  and g42333 (n25377, n10434, n22332);
  and g42339 (n25380, n9870, n_16827);
  not g42342 (n_17057, n25381);
  and g42343 (n25382, \a[5] , n_17057);
  not g42344 (n_17058, n25382);
  and g42345 (n25383, n_17057, n_17058);
  and g42346 (n25384, \a[5] , n_17058);
  not g42347 (n_17059, n25383);
  not g42348 (n_17060, n25384);
  and g42349 (n25385, n_17059, n_17060);
  not g42350 (n_17061, n25074);
  and g42351 (n25386, n25072, n_17061);
  not g42352 (n_17062, n25386);
  and g42353 (n25387, n_16799, n_17062);
  not g42354 (n_17063, n25385);
  and g42355 (n25388, n_17063, n25387);
  not g42356 (n_17064, n25388);
  and g42357 (n25389, n_17063, n_17064);
  and g42358 (n25390, n25387, n_17064);
  not g42359 (n_17065, n25389);
  not g42360 (n_17066, n25390);
  and g42361 (n25391, n_17065, n_17066);
  and g42362 (n25392, n71, n22332);
  and g42363 (n25393, n9867, n22338);
  and g42364 (n25394, n10434, n22335);
  and g42370 (n25397, n9870, n22542);
  not g42373 (n_17071, n25398);
  and g42374 (n25399, \a[5] , n_17071);
  not g42375 (n_17072, n25399);
  and g42376 (n25400, n_17071, n_17072);
  and g42377 (n25401, \a[5] , n_17072);
  not g42378 (n_17073, n25400);
  not g42379 (n_17074, n25401);
  and g42380 (n25402, n_17073, n_17074);
  and g42381 (n25403, n_16792, n_16794);
  and g42382 (n25404, n_16793, n_16794);
  not g42383 (n_17075, n25403);
  not g42384 (n_17076, n25404);
  and g42385 (n25405, n_17075, n_17076);
  not g42386 (n_17077, n25402);
  not g42387 (n_17078, n25405);
  and g42388 (n25406, n_17077, n_17078);
  not g42389 (n_17079, n25406);
  and g42390 (n25407, n_17077, n_17079);
  and g42391 (n25408, n_17078, n_17079);
  not g42392 (n_17080, n25407);
  not g42393 (n_17081, n25408);
  and g42394 (n25409, n_17080, n_17081);
  and g42395 (n25410, n71, n22335);
  and g42396 (n25411, n9867, n22341);
  and g42397 (n25412, n10434, n22338);
  and g42403 (n25415, n9870, n_16015);
  not g42406 (n_17086, n25416);
  and g42407 (n25417, \a[5] , n_17086);
  not g42408 (n_17087, n25417);
  and g42409 (n25418, n_17086, n_17087);
  and g42410 (n25419, \a[5] , n_17087);
  not g42411 (n_17088, n25418);
  not g42412 (n_17089, n25419);
  and g42413 (n25420, n_17088, n_17089);
  and g42414 (n25421, n_16786, n_16788);
  and g42415 (n25422, n_16787, n_16788);
  not g42416 (n_17090, n25421);
  not g42417 (n_17091, n25422);
  and g42418 (n25423, n_17090, n_17091);
  not g42419 (n_17092, n25420);
  not g42420 (n_17093, n25423);
  and g42421 (n25424, n_17092, n_17093);
  not g42422 (n_17094, n25424);
  and g42423 (n25425, n_17092, n_17094);
  and g42424 (n25426, n_17093, n_17094);
  not g42425 (n_17095, n25425);
  not g42426 (n_17096, n25426);
  and g42427 (n25427, n_17095, n_17096);
  and g42428 (n25428, n24733, n25060);
  not g42429 (n_17097, n25428);
  and g42430 (n25429, n_16782, n_17097);
  and g42431 (n25430, n71, n22338);
  and g42432 (n25431, n9867, n22344);
  and g42433 (n25432, n10434, n22341);
  not g42434 (n_17098, n25431);
  not g42435 (n_17099, n25432);
  and g42436 (n25433, n_17098, n_17099);
  not g42437 (n_17100, n25430);
  and g42438 (n25434, n_17100, n25433);
  and g42439 (n25435, n_4684, n25434);
  and g42440 (n25436, n24188, n25434);
  not g42441 (n_17101, n25435);
  not g42442 (n_17102, n25436);
  and g42443 (n25437, n_17101, n_17102);
  not g42444 (n_17103, n25437);
  and g42445 (n25438, \a[5] , n_17103);
  and g42446 (n25439, n_3, n25437);
  not g42447 (n_17104, n25438);
  not g42448 (n_17105, n25439);
  and g42449 (n25440, n_17104, n_17105);
  not g42450 (n_17106, n25440);
  and g42451 (n25441, n25429, n_17106);
  and g42452 (n25442, n24751, n25058);
  not g42453 (n_17107, n25442);
  and g42454 (n25443, n_16779, n_17107);
  and g42455 (n25444, n71, n22341);
  and g42456 (n25445, n9867, n22347);
  and g42457 (n25446, n10434, n22344);
  not g42458 (n_17108, n25445);
  not g42459 (n_17109, n25446);
  and g42460 (n25447, n_17108, n_17109);
  not g42461 (n_17110, n25444);
  and g42462 (n25448, n_17110, n25447);
  and g42463 (n25449, n_4684, n25448);
  and g42464 (n25450, n_15990, n25448);
  not g42465 (n_17111, n25449);
  not g42466 (n_17112, n25450);
  and g42467 (n25451, n_17111, n_17112);
  not g42468 (n_17113, n25451);
  and g42469 (n25452, \a[5] , n_17113);
  and g42470 (n25453, n_3, n25451);
  not g42471 (n_17114, n25452);
  not g42472 (n_17115, n25453);
  and g42473 (n25454, n_17114, n_17115);
  not g42474 (n_17116, n25454);
  and g42475 (n25455, n25443, n_17116);
  and g42476 (n25456, n24769, n25056);
  not g42477 (n_17117, n25456);
  and g42478 (n25457, n_16776, n_17117);
  and g42479 (n25458, n71, n22344);
  and g42480 (n25459, n9867, n22350);
  and g42481 (n25460, n10434, n22347);
  not g42482 (n_17118, n25459);
  not g42483 (n_17119, n25460);
  and g42484 (n25461, n_17118, n_17119);
  not g42485 (n_17120, n25458);
  and g42486 (n25462, n_17120, n25461);
  and g42487 (n25463, n_4684, n25462);
  and g42488 (n25464, n23642, n25462);
  not g42489 (n_17121, n25463);
  not g42490 (n_17122, n25464);
  and g42491 (n25465, n_17121, n_17122);
  not g42492 (n_17123, n25465);
  and g42493 (n25466, \a[5] , n_17123);
  and g42494 (n25467, n_3, n25465);
  not g42495 (n_17124, n25466);
  not g42496 (n_17125, n25467);
  and g42497 (n25468, n_17124, n_17125);
  not g42498 (n_17126, n25468);
  and g42499 (n25469, n25457, n_17126);
  and g42500 (n25470, n71, n22347);
  and g42501 (n25471, n9867, n22353);
  and g42502 (n25472, n10434, n22350);
  and g42508 (n25475, n9870, n_16069);
  not g42511 (n_17131, n25476);
  and g42512 (n25477, \a[5] , n_17131);
  not g42513 (n_17132, n25477);
  and g42514 (n25478, n_17131, n_17132);
  and g42515 (n25479, \a[5] , n_17132);
  not g42516 (n_17133, n25478);
  not g42517 (n_17134, n25479);
  and g42518 (n25480, n_17133, n_17134);
  not g42519 (n_17135, n25054);
  and g42520 (n25481, n25052, n_17135);
  not g42521 (n_17136, n25481);
  and g42522 (n25482, n_16773, n_17136);
  not g42523 (n_17137, n25480);
  and g42524 (n25483, n_17137, n25482);
  not g42525 (n_17138, n25483);
  and g42526 (n25484, n_17137, n_17138);
  and g42527 (n25485, n25482, n_17138);
  not g42528 (n_17139, n25484);
  not g42529 (n_17140, n25485);
  and g42530 (n25486, n_17139, n_17140);
  and g42531 (n25487, n71, n22350);
  and g42532 (n25488, n9867, n22356);
  and g42533 (n25489, n10434, n22353);
  and g42539 (n25492, n9870, n23672);
  not g42542 (n_17145, n25493);
  and g42543 (n25494, \a[5] , n_17145);
  not g42544 (n_17146, n25494);
  and g42545 (n25495, n_17145, n_17146);
  and g42546 (n25496, \a[5] , n_17146);
  not g42547 (n_17147, n25495);
  not g42548 (n_17148, n25496);
  and g42549 (n25497, n_17147, n_17148);
  and g42550 (n25498, n_16766, n_16768);
  and g42551 (n25499, n_16767, n_16768);
  not g42552 (n_17149, n25498);
  not g42553 (n_17150, n25499);
  and g42554 (n25500, n_17149, n_17150);
  not g42555 (n_17151, n25497);
  not g42556 (n_17152, n25500);
  and g42557 (n25501, n_17151, n_17152);
  not g42558 (n_17153, n25501);
  and g42559 (n25502, n_17151, n_17153);
  and g42560 (n25503, n_17152, n_17153);
  not g42561 (n_17154, n25502);
  not g42562 (n_17155, n25503);
  and g42563 (n25504, n_17154, n_17155);
  and g42564 (n25505, n71, n22353);
  and g42565 (n25506, n9867, n22359);
  and g42566 (n25507, n10434, n22356);
  and g42572 (n25510, n9870, n_14678);
  not g42575 (n_17160, n25511);
  and g42576 (n25512, \a[5] , n_17160);
  not g42577 (n_17161, n25512);
  and g42578 (n25513, n_17160, n_17161);
  and g42579 (n25514, \a[5] , n_17161);
  not g42580 (n_17162, n25513);
  not g42581 (n_17163, n25514);
  and g42582 (n25515, n_17162, n_17163);
  and g42583 (n25516, n_16760, n_16762);
  and g42584 (n25517, n_16761, n_16762);
  not g42585 (n_17164, n25516);
  not g42586 (n_17165, n25517);
  and g42587 (n25518, n_17164, n_17165);
  not g42588 (n_17166, n25515);
  not g42589 (n_17167, n25518);
  and g42590 (n25519, n_17166, n_17167);
  not g42591 (n_17168, n25519);
  and g42592 (n25520, n_17166, n_17168);
  and g42593 (n25521, n_17167, n_17168);
  not g42594 (n_17169, n25520);
  not g42595 (n_17170, n25521);
  and g42596 (n25522, n_17169, n_17170);
  and g42597 (n25523, n24828, n25040);
  not g42598 (n_17171, n25523);
  and g42599 (n25524, n_16756, n_17171);
  and g42600 (n25525, n71, n22356);
  and g42601 (n25526, n9867, n22362);
  and g42602 (n25527, n10434, n22359);
  not g42603 (n_17172, n25526);
  not g42604 (n_17173, n25527);
  and g42605 (n25528, n_17172, n_17173);
  not g42606 (n_17174, n25525);
  and g42607 (n25529, n_17174, n25528);
  and g42608 (n25530, n_4684, n25529);
  and g42609 (n25531, n23345, n25529);
  not g42610 (n_17175, n25530);
  not g42611 (n_17176, n25531);
  and g42612 (n25532, n_17175, n_17176);
  not g42613 (n_17177, n25532);
  and g42614 (n25533, \a[5] , n_17177);
  and g42615 (n25534, n_3, n25532);
  not g42616 (n_17178, n25533);
  not g42617 (n_17179, n25534);
  and g42618 (n25535, n_17178, n_17179);
  not g42619 (n_17180, n25535);
  and g42620 (n25536, n25524, n_17180);
  and g42621 (n25537, n24846, n25038);
  not g42622 (n_17181, n25537);
  and g42623 (n25538, n_16753, n_17181);
  and g42624 (n25539, n71, n22359);
  and g42625 (n25540, n9867, n22365);
  and g42626 (n25541, n10434, n22362);
  not g42627 (n_17182, n25540);
  not g42628 (n_17183, n25541);
  and g42629 (n25542, n_17182, n_17183);
  not g42630 (n_17184, n25539);
  and g42631 (n25543, n_17184, n25542);
  and g42632 (n25544, n_4684, n25543);
  and g42633 (n25545, n_15331, n25543);
  not g42634 (n_17185, n25544);
  not g42635 (n_17186, n25545);
  and g42636 (n25546, n_17185, n_17186);
  not g42637 (n_17187, n25546);
  and g42638 (n25547, \a[5] , n_17187);
  and g42639 (n25548, n_3, n25546);
  not g42640 (n_17188, n25547);
  not g42641 (n_17189, n25548);
  and g42642 (n25549, n_17188, n_17189);
  not g42643 (n_17190, n25549);
  and g42644 (n25550, n25538, n_17190);
  and g42645 (n25551, n24864, n25036);
  not g42646 (n_17191, n25551);
  and g42647 (n25552, n_16750, n_17191);
  and g42648 (n25553, n71, n22362);
  and g42649 (n25554, n9867, n22368);
  and g42650 (n25555, n10434, n22365);
  not g42651 (n_17192, n25554);
  not g42652 (n_17193, n25555);
  and g42653 (n25556, n_17192, n_17193);
  not g42654 (n_17194, n25553);
  and g42655 (n25557, n_17194, n25556);
  and g42656 (n25558, n_4684, n25557);
  and g42657 (n25559, n23320, n25557);
  not g42658 (n_17195, n25558);
  not g42659 (n_17196, n25559);
  and g42660 (n25560, n_17195, n_17196);
  not g42661 (n_17197, n25560);
  and g42662 (n25561, \a[5] , n_17197);
  and g42663 (n25562, n_3, n25560);
  not g42664 (n_17198, n25561);
  not g42665 (n_17199, n25562);
  and g42666 (n25563, n_17198, n_17199);
  not g42667 (n_17200, n25563);
  and g42668 (n25564, n25552, n_17200);
  and g42669 (n25565, n71, n22365);
  and g42670 (n25566, n9867, n22371);
  and g42671 (n25567, n10434, n22368);
  and g42677 (n25570, n9870, n_15351);
  not g42680 (n_17205, n25571);
  and g42681 (n25572, \a[5] , n_17205);
  not g42682 (n_17206, n25572);
  and g42683 (n25573, n_17205, n_17206);
  and g42684 (n25574, \a[5] , n_17206);
  not g42685 (n_17207, n25573);
  not g42686 (n_17208, n25574);
  and g42687 (n25575, n_17207, n_17208);
  not g42688 (n_17209, n25034);
  and g42689 (n25576, n25032, n_17209);
  not g42690 (n_17210, n25576);
  and g42691 (n25577, n_16747, n_17210);
  not g42692 (n_17211, n25575);
  and g42693 (n25578, n_17211, n25577);
  not g42694 (n_17212, n25578);
  and g42695 (n25579, n_17211, n_17212);
  and g42696 (n25580, n25577, n_17212);
  not g42697 (n_17213, n25579);
  not g42698 (n_17214, n25580);
  and g42699 (n25581, n_17213, n_17214);
  and g42700 (n25582, n71, n22368);
  and g42701 (n25583, n9867, n22374);
  and g42702 (n25584, n10434, n22371);
  and g42708 (n25587, n9870, n23006);
  not g42711 (n_17219, n25588);
  and g42712 (n25589, \a[5] , n_17219);
  not g42713 (n_17220, n25589);
  and g42714 (n25590, n_17219, n_17220);
  and g42715 (n25591, \a[5] , n_17220);
  not g42716 (n_17221, n25590);
  not g42717 (n_17222, n25591);
  and g42718 (n25592, n_17221, n_17222);
  and g42719 (n25593, n_16740, n_16742);
  and g42720 (n25594, n_16741, n_16742);
  not g42721 (n_17223, n25593);
  not g42722 (n_17224, n25594);
  and g42723 (n25595, n_17223, n_17224);
  not g42724 (n_17225, n25592);
  not g42725 (n_17226, n25595);
  and g42726 (n25596, n_17225, n_17226);
  not g42727 (n_17227, n25596);
  and g42728 (n25597, n_17225, n_17227);
  and g42729 (n25598, n_17226, n_17227);
  not g42730 (n_17228, n25597);
  not g42731 (n_17229, n25598);
  and g42732 (n25599, n_17228, n_17229);
  and g42733 (n25600, n71, n22371);
  and g42734 (n25601, n9867, n22377);
  and g42735 (n25602, n10434, n22374);
  and g42741 (n25605, n9870, n23025);
  not g42744 (n_17234, n25606);
  and g42745 (n25607, \a[5] , n_17234);
  not g42746 (n_17235, n25607);
  and g42747 (n25608, n_17234, n_17235);
  and g42748 (n25609, \a[5] , n_17235);
  not g42749 (n_17236, n25608);
  not g42750 (n_17237, n25609);
  and g42751 (n25610, n_17236, n_17237);
  and g42752 (n25611, n_16734, n_16736);
  and g42753 (n25612, n_16735, n_16736);
  not g42754 (n_17238, n25611);
  not g42755 (n_17239, n25612);
  and g42756 (n25613, n_17238, n_17239);
  not g42757 (n_17240, n25610);
  not g42758 (n_17241, n25613);
  and g42759 (n25614, n_17240, n_17241);
  not g42760 (n_17242, n25614);
  and g42761 (n25615, n_17240, n_17242);
  and g42762 (n25616, n_17241, n_17242);
  not g42763 (n_17243, n25615);
  not g42764 (n_17244, n25616);
  and g42765 (n25617, n_17243, n_17244);
  and g42766 (n25618, n24923, n25020);
  not g42767 (n_17245, n25618);
  and g42768 (n25619, n_16730, n_17245);
  and g42769 (n25620, n71, n22374);
  and g42770 (n25621, n9867, n22380);
  and g42771 (n25622, n10434, n22377);
  not g42772 (n_17246, n25621);
  not g42773 (n_17247, n25622);
  and g42774 (n25623, n_17246, n_17247);
  not g42775 (n_17248, n25620);
  and g42776 (n25624, n_17248, n25623);
  and g42777 (n25625, n_4684, n25624);
  and g42778 (n25626, n_15064, n25624);
  not g42779 (n_17249, n25625);
  not g42780 (n_17250, n25626);
  and g42781 (n25627, n_17249, n_17250);
  not g42782 (n_17251, n25627);
  and g42783 (n25628, \a[5] , n_17251);
  and g42784 (n25629, n_3, n25627);
  not g42785 (n_17252, n25628);
  not g42786 (n_17253, n25629);
  and g42787 (n25630, n_17252, n_17253);
  not g42788 (n_17254, n25630);
  and g42789 (n25631, n25619, n_17254);
  not g42790 (n_17255, n25018);
  and g42791 (n25632, n25016, n_17255);
  not g42792 (n_17256, n25632);
  and g42793 (n25633, n_16727, n_17256);
  and g42794 (n25634, n71, n22377);
  and g42795 (n25635, n9867, n22384);
  and g42796 (n25636, n10434, n22380);
  not g42797 (n_17257, n25635);
  not g42798 (n_17258, n25636);
  and g42799 (n25637, n_17257, n_17258);
  not g42800 (n_17259, n25634);
  and g42801 (n25638, n_17259, n25637);
  and g42802 (n25639, n_4684, n25638);
  and g42803 (n25640, n22834, n25638);
  not g42804 (n_17260, n25639);
  not g42805 (n_17261, n25640);
  and g42806 (n25641, n_17260, n_17261);
  not g42807 (n_17262, n25641);
  and g42808 (n25642, \a[5] , n_17262);
  and g42809 (n25643, n_3, n25641);
  not g42810 (n_17263, n25642);
  not g42811 (n_17264, n25643);
  and g42812 (n25644, n_17263, n_17264);
  not g42813 (n_17265, n25644);
  and g42814 (n25645, n25633, n_17265);
  and g42815 (n25646, n24955, n25014);
  not g42816 (n_17266, n25646);
  and g42817 (n25647, n_16723, n_17266);
  and g42818 (n25648, n71, n22380);
  and g42819 (n25649, n9867, n22387);
  and g42820 (n25650, n10434, n22384);
  not g42821 (n_17267, n25649);
  not g42822 (n_17268, n25650);
  and g42823 (n25651, n_17267, n_17268);
  not g42824 (n_17269, n25648);
  and g42825 (n25652, n_17269, n25651);
  and g42826 (n25653, n_4684, n25652);
  and g42827 (n25654, n_14894, n25652);
  not g42828 (n_17270, n25653);
  not g42829 (n_17271, n25654);
  and g42830 (n25655, n_17270, n_17271);
  not g42831 (n_17272, n25655);
  and g42832 (n25656, \a[5] , n_17272);
  and g42833 (n25657, n_3, n25655);
  not g42834 (n_17273, n25656);
  not g42835 (n_17274, n25657);
  and g42836 (n25658, n_17273, n_17274);
  not g42837 (n_17275, n25658);
  and g42838 (n25659, n25647, n_17275);
  and g42839 (n25660, n71, n22384);
  and g42840 (n25661, n9867, n22390);
  and g42841 (n25662, n10434, n22387);
  and g42847 (n25665, n9870, n22806);
  not g42850 (n_17280, n25666);
  and g42851 (n25667, \a[5] , n_17280);
  not g42852 (n_17281, n25667);
  and g42853 (n25668, n_17280, n_17281);
  and g42854 (n25669, \a[5] , n_17281);
  not g42855 (n_17282, n25668);
  not g42856 (n_17283, n25669);
  and g42857 (n25670, n_17282, n_17283);
  not g42858 (n_17284, n25012);
  and g42859 (n25671, n25010, n_17284);
  not g42860 (n_17285, n25671);
  and g42861 (n25672, n_16720, n_17285);
  not g42862 (n_17286, n25670);
  and g42863 (n25673, n_17286, n25672);
  not g42864 (n_17287, n25673);
  and g42865 (n25674, n_17286, n_17287);
  and g42866 (n25675, n25672, n_17287);
  not g42867 (n_17288, n25674);
  not g42868 (n_17289, n25675);
  and g42869 (n25676, n_17288, n_17289);
  and g42870 (n25677, n_16713, n_16715);
  and g42871 (n25678, n_16714, n_16715);
  not g42872 (n_17290, n25677);
  not g42873 (n_17291, n25678);
  and g42874 (n25679, n_17290, n_17291);
  and g42875 (n25680, n71, n22387);
  and g42876 (n25681, n9867, n22393);
  and g42877 (n25682, n10434, n22390);
  not g42878 (n_17292, n25681);
  not g42879 (n_17293, n25682);
  and g42880 (n25683, n_17292, n_17293);
  not g42881 (n_17294, n25680);
  and g42882 (n25684, n_17294, n25683);
  and g42883 (n25685, n_4684, n25684);
  and g42884 (n25686, n_14920, n25684);
  not g42885 (n_17295, n25685);
  not g42886 (n_17296, n25686);
  and g42887 (n25687, n_17295, n_17296);
  not g42888 (n_17297, n25687);
  and g42889 (n25688, \a[5] , n_17297);
  and g42890 (n25689, n_3, n25687);
  not g42891 (n_17298, n25688);
  not g42892 (n_17299, n25689);
  and g42893 (n25690, n_17298, n_17299);
  not g42894 (n_17300, n25679);
  not g42895 (n_17301, n25690);
  and g42896 (n25691, n_17300, n_17301);
  and g42897 (n25692, n71, n22390);
  and g42898 (n25693, n9867, n22396);
  and g42899 (n25694, n10434, n22393);
  and g42905 (n25697, n9870, n22649);
  not g42908 (n_17306, n25698);
  and g42909 (n25699, \a[5] , n_17306);
  not g42910 (n_17307, n25699);
  and g42911 (n25700, n_17306, n_17307);
  and g42912 (n25701, \a[5] , n_17307);
  not g42913 (n_17308, n25700);
  not g42914 (n_17309, n25701);
  and g42915 (n25702, n_17308, n_17309);
  not g42916 (n_17310, n24981);
  and g42917 (n25703, n_17310, n24992);
  not g42918 (n_17311, n24993);
  not g42919 (n_17312, n25703);
  and g42920 (n25704, n_17311, n_17312);
  not g42921 (n_17313, n25702);
  and g42922 (n25705, n_17313, n25704);
  not g42923 (n_17314, n25705);
  and g42924 (n25706, n_17313, n_17314);
  and g42925 (n25707, n25704, n_17314);
  not g42926 (n_17315, n25706);
  not g42927 (n_17316, n25707);
  and g42928 (n25708, n_17315, n_17316);
  not g42929 (n_17317, n24980);
  and g42930 (n25709, n24978, n_17317);
  not g42931 (n_17318, n25709);
  and g42932 (n25710, n_17310, n_17318);
  and g42933 (n25711, n71, n22393);
  and g42934 (n25712, n9867, n22399);
  and g42935 (n25713, n10434, n22396);
  not g42936 (n_17319, n25712);
  not g42937 (n_17320, n25713);
  and g42938 (n25714, n_17319, n_17320);
  not g42939 (n_17321, n25711);
  and g42940 (n25715, n_17321, n25714);
  and g42941 (n25716, n_4684, n25715);
  and g42942 (n25717, n_14773, n25715);
  not g42943 (n_17322, n25716);
  not g42944 (n_17323, n25717);
  and g42945 (n25718, n_17322, n_17323);
  not g42946 (n_17324, n25718);
  and g42947 (n25719, \a[5] , n_17324);
  and g42948 (n25720, n_3, n25718);
  not g42949 (n_17325, n25719);
  not g42950 (n_17326, n25720);
  and g42951 (n25721, n_17325, n_17326);
  not g42952 (n_17327, n25721);
  and g42953 (n25722, n25710, n_17327);
  and g42954 (n25723, n10434, n_14508);
  and g42955 (n25724, n71, n22402);
  not g42956 (n_17328, n25723);
  not g42957 (n_17329, n25724);
  and g42958 (n25725, n_17328, n_17329);
  and g42959 (n25726, n9870, n_14720);
  not g42960 (n_17330, n25726);
  and g42961 (n25727, n25725, n_17330);
  not g42962 (n_17331, n25727);
  and g42963 (n25728, \a[5] , n_17331);
  not g42964 (n_17332, n25728);
  and g42965 (n25729, \a[5] , n_17332);
  and g42966 (n25730, n_17331, n_17332);
  not g42967 (n_17333, n25729);
  not g42968 (n_17334, n25730);
  and g42969 (n25731, n_17333, n_17334);
  and g42970 (n25732, n_13, n_14508);
  not g42971 (n_17335, n25732);
  and g42972 (n25733, \a[5] , n_17335);
  not g42973 (n_17336, n25731);
  and g42974 (n25734, n_17336, n25733);
  and g42975 (n25735, n71, n22399);
  and g42976 (n25736, n9867, n_14508);
  and g42977 (n25737, n10434, n22402);
  not g42978 (n_17337, n25736);
  not g42979 (n_17338, n25737);
  and g42980 (n25738, n_17337, n_17338);
  not g42981 (n_17339, n25735);
  and g42982 (n25739, n_17339, n25738);
  and g42983 (n25740, n_4684, n25739);
  and g42984 (n25741, n22625, n25739);
  not g42985 (n_17340, n25740);
  not g42986 (n_17341, n25741);
  and g42987 (n25742, n_17340, n_17341);
  not g42988 (n_17342, n25742);
  and g42989 (n25743, \a[5] , n_17342);
  and g42990 (n25744, n_3, n25742);
  not g42991 (n_17343, n25743);
  not g42992 (n_17344, n25744);
  and g42993 (n25745, n_17343, n_17344);
  not g42994 (n_17345, n25745);
  and g42995 (n25746, n25734, n_17345);
  and g42996 (n25747, n24979, n25746);
  not g42997 (n_17346, n25747);
  and g42998 (n25748, n25746, n_17346);
  and g42999 (n25749, n24979, n_17346);
  not g43000 (n_17347, n25748);
  not g43001 (n_17348, n25749);
  and g43002 (n25750, n_17347, n_17348);
  and g43003 (n25751, n71, n22396);
  and g43004 (n25752, n9867, n22402);
  and g43005 (n25753, n10434, n22399);
  and g43011 (n25756, n9870, n22595);
  not g43014 (n_17353, n25757);
  and g43015 (n25758, \a[5] , n_17353);
  not g43016 (n_17354, n25758);
  and g43017 (n25759, \a[5] , n_17354);
  and g43018 (n25760, n_17353, n_17354);
  not g43019 (n_17355, n25759);
  not g43020 (n_17356, n25760);
  and g43021 (n25761, n_17355, n_17356);
  not g43022 (n_17357, n25750);
  not g43023 (n_17358, n25761);
  and g43024 (n25762, n_17357, n_17358);
  not g43025 (n_17359, n25762);
  and g43026 (n25763, n_17346, n_17359);
  not g43027 (n_17360, n25710);
  and g43028 (n25764, n_17360, n25721);
  not g43029 (n_17361, n25722);
  not g43030 (n_17362, n25764);
  and g43031 (n25765, n_17361, n_17362);
  not g43032 (n_17363, n25763);
  and g43033 (n25766, n_17363, n25765);
  not g43034 (n_17364, n25766);
  and g43035 (n25767, n_17361, n_17364);
  not g43036 (n_17365, n25708);
  not g43037 (n_17366, n25767);
  and g43038 (n25768, n_17365, n_17366);
  not g43039 (n_17367, n25768);
  and g43040 (n25769, n_17314, n_17367);
  and g43041 (n25770, n25679, n25690);
  not g43042 (n_17368, n25691);
  not g43043 (n_17369, n25770);
  and g43044 (n25771, n_17368, n_17369);
  not g43045 (n_17370, n25769);
  and g43046 (n25772, n_17370, n25771);
  not g43047 (n_17371, n25772);
  and g43048 (n25773, n_17368, n_17371);
  not g43049 (n_17372, n25676);
  not g43050 (n_17373, n25773);
  and g43051 (n25774, n_17372, n_17373);
  not g43052 (n_17374, n25774);
  and g43053 (n25775, n_17287, n_17374);
  not g43054 (n_17375, n25659);
  and g43055 (n25776, n25647, n_17375);
  and g43056 (n25777, n_17275, n_17375);
  not g43057 (n_17376, n25776);
  not g43058 (n_17377, n25777);
  and g43059 (n25778, n_17376, n_17377);
  not g43060 (n_17378, n25775);
  not g43061 (n_17379, n25778);
  and g43062 (n25779, n_17378, n_17379);
  not g43063 (n_17380, n25779);
  and g43064 (n25780, n_17375, n_17380);
  not g43065 (n_17381, n25645);
  and g43066 (n25781, n25633, n_17381);
  and g43067 (n25782, n_17265, n_17381);
  not g43068 (n_17382, n25781);
  not g43069 (n_17383, n25782);
  and g43070 (n25783, n_17382, n_17383);
  not g43071 (n_17384, n25780);
  not g43072 (n_17385, n25783);
  and g43073 (n25784, n_17384, n_17385);
  not g43074 (n_17386, n25784);
  and g43075 (n25785, n_17381, n_17386);
  not g43076 (n_17387, n25619);
  and g43077 (n25786, n_17387, n25630);
  not g43078 (n_17388, n25631);
  not g43079 (n_17389, n25786);
  and g43080 (n25787, n_17388, n_17389);
  not g43081 (n_17390, n25785);
  and g43082 (n25788, n_17390, n25787);
  not g43083 (n_17391, n25788);
  and g43084 (n25789, n_17388, n_17391);
  not g43085 (n_17392, n25617);
  not g43086 (n_17393, n25789);
  and g43087 (n25790, n_17392, n_17393);
  not g43088 (n_17394, n25790);
  and g43089 (n25791, n_17242, n_17394);
  not g43090 (n_17395, n25599);
  not g43091 (n_17396, n25791);
  and g43092 (n25792, n_17395, n_17396);
  not g43093 (n_17397, n25792);
  and g43094 (n25793, n_17227, n_17397);
  not g43095 (n_17398, n25581);
  not g43096 (n_17399, n25793);
  and g43097 (n25794, n_17398, n_17399);
  not g43098 (n_17400, n25794);
  and g43099 (n25795, n_17212, n_17400);
  not g43100 (n_17401, n25564);
  and g43101 (n25796, n25552, n_17401);
  and g43102 (n25797, n_17200, n_17401);
  not g43103 (n_17402, n25796);
  not g43104 (n_17403, n25797);
  and g43105 (n25798, n_17402, n_17403);
  not g43106 (n_17404, n25795);
  not g43107 (n_17405, n25798);
  and g43108 (n25799, n_17404, n_17405);
  not g43109 (n_17406, n25799);
  and g43110 (n25800, n_17401, n_17406);
  not g43111 (n_17407, n25550);
  and g43112 (n25801, n25538, n_17407);
  and g43113 (n25802, n_17190, n_17407);
  not g43114 (n_17408, n25801);
  not g43115 (n_17409, n25802);
  and g43116 (n25803, n_17408, n_17409);
  not g43117 (n_17410, n25800);
  not g43118 (n_17411, n25803);
  and g43119 (n25804, n_17410, n_17411);
  not g43120 (n_17412, n25804);
  and g43121 (n25805, n_17407, n_17412);
  not g43122 (n_17413, n25524);
  and g43123 (n25806, n_17413, n25535);
  not g43124 (n_17414, n25536);
  not g43125 (n_17415, n25806);
  and g43126 (n25807, n_17414, n_17415);
  not g43127 (n_17416, n25805);
  and g43128 (n25808, n_17416, n25807);
  not g43129 (n_17417, n25808);
  and g43130 (n25809, n_17414, n_17417);
  not g43131 (n_17418, n25522);
  not g43132 (n_17419, n25809);
  and g43133 (n25810, n_17418, n_17419);
  not g43134 (n_17420, n25810);
  and g43135 (n25811, n_17168, n_17420);
  not g43136 (n_17421, n25504);
  not g43137 (n_17422, n25811);
  and g43138 (n25812, n_17421, n_17422);
  not g43139 (n_17423, n25812);
  and g43140 (n25813, n_17153, n_17423);
  not g43141 (n_17424, n25486);
  not g43142 (n_17425, n25813);
  and g43143 (n25814, n_17424, n_17425);
  not g43144 (n_17426, n25814);
  and g43145 (n25815, n_17138, n_17426);
  not g43146 (n_17427, n25469);
  and g43147 (n25816, n25457, n_17427);
  and g43148 (n25817, n_17126, n_17427);
  not g43149 (n_17428, n25816);
  not g43150 (n_17429, n25817);
  and g43151 (n25818, n_17428, n_17429);
  not g43152 (n_17430, n25815);
  not g43153 (n_17431, n25818);
  and g43154 (n25819, n_17430, n_17431);
  not g43155 (n_17432, n25819);
  and g43156 (n25820, n_17427, n_17432);
  not g43157 (n_17433, n25455);
  and g43158 (n25821, n25443, n_17433);
  and g43159 (n25822, n_17116, n_17433);
  not g43160 (n_17434, n25821);
  not g43161 (n_17435, n25822);
  and g43162 (n25823, n_17434, n_17435);
  not g43163 (n_17436, n25820);
  not g43164 (n_17437, n25823);
  and g43165 (n25824, n_17436, n_17437);
  not g43166 (n_17438, n25824);
  and g43167 (n25825, n_17433, n_17438);
  not g43168 (n_17439, n25429);
  and g43169 (n25826, n_17439, n25440);
  not g43170 (n_17440, n25441);
  not g43171 (n_17441, n25826);
  and g43172 (n25827, n_17440, n_17441);
  not g43173 (n_17442, n25825);
  and g43174 (n25828, n_17442, n25827);
  not g43175 (n_17443, n25828);
  and g43176 (n25829, n_17440, n_17443);
  not g43177 (n_17444, n25427);
  not g43178 (n_17445, n25829);
  and g43179 (n25830, n_17444, n_17445);
  not g43180 (n_17446, n25830);
  and g43181 (n25831, n_17094, n_17446);
  not g43182 (n_17447, n25409);
  not g43183 (n_17448, n25831);
  and g43184 (n25832, n_17447, n_17448);
  not g43185 (n_17449, n25832);
  and g43186 (n25833, n_17079, n_17449);
  not g43187 (n_17450, n25391);
  not g43188 (n_17451, n25833);
  and g43189 (n25834, n_17450, n_17451);
  not g43190 (n_17452, n25834);
  and g43191 (n25835, n_17064, n_17452);
  not g43192 (n_17453, n25374);
  and g43193 (n25836, n25362, n_17453);
  and g43194 (n25837, n_17052, n_17453);
  not g43195 (n_17454, n25836);
  not g43196 (n_17455, n25837);
  and g43197 (n25838, n_17454, n_17455);
  not g43198 (n_17456, n25835);
  not g43199 (n_17457, n25838);
  and g43200 (n25839, n_17456, n_17457);
  not g43201 (n_17458, n25839);
  and g43202 (n25840, n_17453, n_17458);
  not g43203 (n_17459, n25348);
  and g43204 (n25841, n_17459, n25359);
  not g43205 (n_17460, n25360);
  not g43206 (n_17461, n25841);
  and g43207 (n25842, n_17460, n_17461);
  not g43208 (n_17462, n25840);
  and g43209 (n25843, n_17462, n25842);
  not g43210 (n_17463, n25843);
  and g43211 (n25844, n_17460, n_17463);
  not g43212 (n_17464, n25346);
  not g43213 (n_17465, n25844);
  and g43214 (n25845, n_17464, n_17465);
  not g43215 (n_17466, n25845);
  and g43216 (n25846, n_17030, n_17466);
  not g43217 (n_17467, n25328);
  not g43218 (n_17468, n25846);
  and g43219 (n25847, n_17467, n_17468);
  not g43220 (n_17469, n25847);
  and g43221 (n25848, n_17014, n_17469);
  not g43222 (n_17470, n25307);
  not g43223 (n_17471, n25848);
  and g43224 (n25849, n_17470, n_17471);
  not g43225 (n_17472, n25849);
  and g43226 (n25850, n_16996, n_17472);
  and g43227 (n25851, n25287, n25850);
  not g43228 (n_17473, n25287);
  not g43229 (n_17474, n25850);
  and g43230 (n25852, n_17473, n_17474);
  not g43231 (n_17475, n25851);
  not g43232 (n_17476, n25852);
  and g43233 (n25853, n_17475, n_17476);
  and g43234 (n25854, n_14422, n_14432);
  and g43235 (n25855, n_14413, n_14416);
  and g43236 (n25856, n_14406, n_14409);
  not g43255 (n_17477, n25856);
  and g43256 (n25875, n_17477, n25874);
  not g43257 (n_17478, n25874);
  and g43258 (n25876, n25856, n_17478);
  not g43259 (n_17479, n25875);
  not g43260 (n_17480, n25876);
  and g43261 (n25877, n_17479, n_17480);
  and g43262 (n25878, n3020, n13515);
  and g43263 (n25879, n3028, n13521);
  and g43264 (n25880, n3023, n13518);
  and g43265 (n25881, n75, n13541);
  not g43273 (n_17485, n25884);
  and g43274 (n25885, n25877, n_17485);
  not g43275 (n_17486, n25877);
  and g43276 (n25886, n_17486, n25884);
  not g43277 (n_17487, n25885);
  not g43278 (n_17488, n25886);
  and g43279 (n25887, n_17487, n_17488);
  not g43280 (n_17489, n25855);
  and g43281 (n25888, n_17489, n25887);
  not g43282 (n_17490, n25887);
  and g43283 (n25889, n25855, n_17490);
  not g43284 (n_17491, n25888);
  not g43285 (n_17492, n25889);
  and g43286 (n25890, n_17491, n_17492);
  and g43287 (n25891, n3457, n13633);
  and g43288 (n25892, n3542, n13597);
  and g43289 (n25893, n3606, n13630);
  not g43290 (n_17493, n25892);
  not g43291 (n_17494, n25893);
  and g43292 (n25894, n_17493, n_17494);
  not g43293 (n_17495, n25891);
  and g43294 (n25895, n_17495, n25894);
  and g43295 (n25896, n_489, n25895);
  and g43296 (n25897, n_13801, n25895);
  not g43297 (n_17496, n25896);
  not g43298 (n_17497, n25897);
  and g43299 (n25898, n_17496, n_17497);
  not g43300 (n_17498, n25898);
  and g43301 (n25899, \a[29] , n_17498);
  and g43302 (n25900, n_15, n25898);
  not g43303 (n_17499, n25899);
  not g43304 (n_17500, n25900);
  and g43305 (n25901, n_17499, n_17500);
  not g43306 (n_17501, n25901);
  and g43307 (n25902, n25890, n_17501);
  not g43308 (n_17502, n25890);
  and g43309 (n25903, n_17502, n25901);
  not g43310 (n_17503, n25902);
  not g43311 (n_17504, n25903);
  and g43312 (n25904, n_17503, n_17504);
  not g43313 (n_17505, n25854);
  and g43314 (n25905, n_17505, n25904);
  not g43315 (n_17506, n25904);
  and g43316 (n25906, n25854, n_17506);
  not g43317 (n_17507, n25905);
  not g43318 (n_17508, n25906);
  and g43319 (n25907, n_17507, n_17508);
  and g43320 (n25908, n3884, n_7417);
  and g43321 (n25909, n3967, n_7540);
  and g43322 (n25910, n4046, n13941);
  and g43328 (n25913, n4050, n14028);
  not g43331 (n_17513, n25914);
  and g43332 (n25915, \a[26] , n_17513);
  not g43333 (n_17514, n25915);
  and g43334 (n25916, \a[26] , n_17514);
  and g43335 (n25917, n_17513, n_17514);
  not g43336 (n_17515, n25916);
  not g43337 (n_17516, n25917);
  and g43338 (n25918, n_17515, n_17516);
  not g43339 (n_17517, n25918);
  and g43340 (n25919, n25907, n_17517);
  not g43341 (n_17518, n25919);
  and g43342 (n25920, n_17507, n_17518);
  and g43343 (n25921, n75, n_7765);
  and g43344 (n25922, n3020, n13597);
  and g43345 (n25923, n3023, n13521);
  and g43346 (n25924, n3028, n13515);
  and g43367 (n25941, n_17478, n25940);
  not g43368 (n_17523, n25940);
  and g43369 (n25942, n25874, n_17523);
  not g43370 (n_17524, n25927);
  not g43371 (n_17525, n25942);
  and g43372 (n25943, n_17524, n_17525);
  not g43373 (n_17526, n25941);
  and g43374 (n25944, n_17526, n25943);
  not g43375 (n_17527, n25944);
  and g43376 (n25945, n_17524, n_17527);
  and g43377 (n25946, n_17525, n_17527);
  and g43378 (n25947, n_17526, n25946);
  not g43379 (n_17528, n25945);
  not g43380 (n_17529, n25947);
  and g43381 (n25948, n_17528, n_17529);
  and g43382 (n25949, n_17479, n_17487);
  and g43383 (n25950, n25948, n25949);
  not g43384 (n_17530, n25948);
  not g43385 (n_17531, n25949);
  and g43386 (n25951, n_17530, n_17531);
  not g43387 (n_17532, n25950);
  not g43388 (n_17533, n25951);
  and g43389 (n25952, n_17532, n_17533);
  and g43390 (n25953, n_17491, n_17503);
  not g43391 (n_17534, n25952);
  and g43392 (n25954, n_17534, n25953);
  not g43393 (n_17535, n25953);
  and g43394 (n25955, n25952, n_17535);
  not g43395 (n_17536, n25954);
  not g43396 (n_17537, n25955);
  and g43397 (n25956, n_17536, n_17537);
  not g43398 (n_17538, n3884);
  not g43399 (n_17539, n4046);
  and g43400 (n25957, n_17538, n_17539);
  not g43401 (n_17540, n25957);
  and g43402 (n25958, n_7417, n_17540);
  and g43403 (n25959, n3967, n13941);
  not g43404 (n_17541, n25958);
  not g43405 (n_17542, n25959);
  and g43406 (n25960, n_17541, n_17542);
  and g43407 (n25961, n4050, n_13153);
  not g43408 (n_17543, n25961);
  and g43409 (n25962, n25960, n_17543);
  not g43410 (n_17544, n25962);
  and g43411 (n25963, \a[26] , n_17544);
  not g43412 (n_17545, n25963);
  and g43413 (n25964, n_17544, n_17545);
  and g43414 (n25965, \a[26] , n_17545);
  not g43415 (n_17546, n25964);
  not g43416 (n_17547, n25965);
  and g43417 (n25966, n_17546, n_17547);
  and g43418 (n25967, n3457, n_7540);
  and g43419 (n25968, n3542, n13630);
  and g43420 (n25969, n3606, n13633);
  and g43426 (n25972, n3368, n_7563);
  not g43429 (n_17552, n25973);
  and g43430 (n25974, \a[29] , n_17552);
  not g43431 (n_17553, n25974);
  and g43432 (n25975, \a[29] , n_17553);
  and g43433 (n25976, n_17552, n_17553);
  not g43434 (n_17554, n25975);
  not g43435 (n_17555, n25976);
  and g43436 (n25977, n_17554, n_17555);
  not g43437 (n_17556, n25966);
  not g43438 (n_17557, n25977);
  and g43439 (n25978, n_17556, n_17557);
  not g43440 (n_17558, n25978);
  and g43441 (n25979, n_17556, n_17558);
  and g43442 (n25980, n_17557, n_17558);
  not g43443 (n_17559, n25979);
  not g43444 (n_17560, n25980);
  and g43445 (n25981, n_17559, n_17560);
  not g43446 (n_17561, n25956);
  and g43447 (n25982, n_17561, n25981);
  not g43448 (n_17562, n25981);
  and g43449 (n25983, n25956, n_17562);
  not g43450 (n_17563, n25982);
  not g43451 (n_17564, n25983);
  and g43452 (n25984, n_17563, n_17564);
  not g43453 (n_17565, n25920);
  and g43454 (n25985, n_17565, n25984);
  and g43455 (n25986, n25907, n_17518);
  and g43456 (n25987, n_17517, n_17518);
  not g43457 (n_17566, n25986);
  not g43458 (n_17567, n25987);
  and g43459 (n25988, n_17566, n_17567);
  and g43460 (n25989, n_14435, n_14436);
  not g43461 (n_17568, n25989);
  and g43462 (n25990, n_14392, n_17568);
  not g43463 (n_17569, n25988);
  not g43464 (n_17570, n25990);
  and g43465 (n25991, n_17569, n_17570);
  not g43466 (n_17571, n25991);
  and g43467 (n25992, n_17569, n_17571);
  and g43468 (n25993, n_17570, n_17571);
  not g43469 (n_17572, n25992);
  not g43470 (n_17573, n25993);
  and g43471 (n25994, n_17572, n_17573);
  and g43472 (n25995, n_14441, n_14445);
  not g43473 (n_17574, n25994);
  not g43474 (n_17575, n25995);
  and g43475 (n25996, n_17574, n_17575);
  not g43476 (n_17576, n25996);
  and g43477 (n25997, n_17571, n_17576);
  not g43478 (n_17577, n25984);
  and g43479 (n25998, n25920, n_17577);
  not g43480 (n_17578, n25985);
  not g43481 (n_17579, n25998);
  and g43482 (n25999, n_17578, n_17579);
  not g43483 (n_17580, n25997);
  and g43484 (n26000, n_17580, n25999);
  not g43485 (n_17581, n26000);
  and g43486 (n26001, n_17578, n_17581);
  and g43487 (n26002, n75, n13976);
  and g43488 (n26003, n3020, n13630);
  and g43489 (n26004, n3023, n13515);
  and g43490 (n26005, n3028, n13597);
  not g43498 (n_17586, n3967);
  and g43499 (n26009, n_17586, n25957);
  and g43500 (n26010, n_750, n26009);
  not g43501 (n_17587, n26010);
  and g43502 (n26011, n_7417, n_17587);
  not g43503 (n_17588, n26011);
  and g43504 (n26012, \a[26] , n_17588);
  and g43505 (n26013, n_33, n26011);
  not g43506 (n_17589, n26012);
  not g43507 (n_17590, n26013);
  and g43508 (n26014, n_17589, n_17590);
  and g43509 (n26015, n3873, n3972);
  and g43510 (n26016, n_123, n26015);
  and g43516 (n26022, n25874, n26021);
  not g43517 (n_17591, n26021);
  and g43518 (n26023, n_17478, n_17591);
  not g43519 (n_17592, n26022);
  not g43520 (n_17593, n26023);
  and g43521 (n26024, n_17592, n_17593);
  and g43522 (n26025, n26014, n26024);
  not g43523 (n_17594, n26014);
  not g43524 (n_17595, n26024);
  and g43525 (n26026, n_17594, n_17595);
  not g43526 (n_17596, n26025);
  not g43527 (n_17597, n26026);
  and g43528 (n26027, n_17596, n_17597);
  not g43529 (n_17598, n25946);
  and g43530 (n26028, n_17598, n26027);
  not g43531 (n_17599, n26027);
  and g43532 (n26029, n25946, n_17599);
  not g43533 (n_17600, n26028);
  not g43534 (n_17601, n26029);
  and g43535 (n26030, n_17600, n_17601);
  not g43536 (n_17602, n26008);
  and g43537 (n26031, n_17602, n26030);
  not g43538 (n_17603, n26031);
  and g43539 (n26032, n26030, n_17603);
  and g43540 (n26033, n_17602, n_17603);
  not g43541 (n_17604, n26032);
  not g43542 (n_17605, n26033);
  and g43543 (n26034, n_17604, n_17605);
  and g43544 (n26035, n3457, n13941);
  and g43545 (n26036, n3542, n13633);
  and g43546 (n26037, n3606, n_7540);
  and g43552 (n26040, n3368, n14136);
  not g43555 (n_17610, n26041);
  and g43556 (n26042, \a[29] , n_17610);
  not g43557 (n_17611, n26042);
  and g43558 (n26043, \a[29] , n_17611);
  and g43559 (n26044, n_17610, n_17611);
  not g43560 (n_17612, n26043);
  not g43561 (n_17613, n26044);
  and g43562 (n26045, n_17612, n_17613);
  not g43563 (n_17614, n26034);
  not g43564 (n_17615, n26045);
  and g43565 (n26046, n_17614, n_17615);
  not g43566 (n_17616, n26046);
  and g43567 (n26047, n_17614, n_17616);
  and g43568 (n26048, n_17615, n_17616);
  not g43569 (n_17617, n26047);
  not g43570 (n_17618, n26048);
  and g43571 (n26049, n_17617, n_17618);
  and g43572 (n26050, n_17533, n_17537);
  and g43573 (n26051, n26049, n26050);
  not g43574 (n_17619, n26049);
  not g43575 (n_17620, n26050);
  and g43576 (n26052, n_17619, n_17620);
  not g43577 (n_17621, n26051);
  not g43578 (n_17622, n26052);
  and g43579 (n26053, n_17621, n_17622);
  and g43580 (n26054, n_17558, n_17564);
  not g43581 (n_17623, n26054);
  and g43582 (n26055, n26053, n_17623);
  not g43583 (n_17624, n26053);
  and g43584 (n26056, n_17624, n26054);
  not g43585 (n_17625, n26055);
  not g43586 (n_17626, n26056);
  and g43587 (n26057, n_17625, n_17626);
  not g43588 (n_17627, n26057);
  and g43589 (n26058, n26001, n_17627);
  not g43590 (n_17628, n26001);
  and g43591 (n26059, n_17628, n26057);
  not g43592 (n_17629, n26058);
  not g43593 (n_17630, n26059);
  and g43594 (n26060, n_17629, n_17630);
  and g43595 (n26061, n11727, n26060);
  and g43596 (n26062, n25994, n25995);
  not g43597 (n_17631, n26062);
  and g43598 (n26063, n_17576, n_17631);
  and g43599 (n26064, n11055, n26063);
  not g43600 (n_17632, n25999);
  and g43601 (n26065, n25997, n_17632);
  not g43602 (n_17633, n26065);
  and g43603 (n26066, n_17581, n_17633);
  and g43604 (n26067, n11715, n26066);
  not g43605 (n_17634, n26064);
  not g43606 (n_17635, n26067);
  and g43607 (n26068, n_17634, n_17635);
  not g43608 (n_17636, n26061);
  and g43609 (n26069, n_17636, n26068);
  and g43610 (n26070, n_6291, n26069);
  and g43611 (n26071, n26063, n26066);
  and g43612 (n26072, n22309, n26063);
  not g43613 (n_17637, n26063);
  and g43614 (n26073, n_14650, n_17637);
  not g43615 (n_17638, n22527);
  not g43616 (n_17639, n26073);
  and g43617 (n26074, n_17638, n_17639);
  not g43618 (n_17640, n26072);
  and g43619 (n26075, n_17640, n26074);
  not g43620 (n_17641, n26075);
  and g43621 (n26076, n_17640, n_17641);
  not g43622 (n_17642, n26066);
  and g43623 (n26077, n_17637, n_17642);
  not g43624 (n_17643, n26076);
  not g43625 (n_17644, n26077);
  and g43626 (n26078, n_17643, n_17644);
  not g43627 (n_17645, n26071);
  and g43628 (n26079, n_17645, n26078);
  not g43629 (n_17646, n26079);
  and g43630 (n26080, n_17645, n_17646);
  and g43631 (n26081, n26060, n26066);
  not g43632 (n_17647, n26060);
  and g43633 (n26082, n_17647, n_17642);
  not g43634 (n_17648, n26080);
  not g43635 (n_17649, n26082);
  and g43636 (n26083, n_17648, n_17649);
  not g43637 (n_17650, n26081);
  and g43638 (n26084, n_17650, n26083);
  not g43639 (n_17651, n26084);
  and g43640 (n26085, n_17648, n_17651);
  and g43641 (n26086, n_17650, n_17651);
  and g43642 (n26087, n_17649, n26086);
  not g43643 (n_17652, n26085);
  not g43644 (n_17653, n26087);
  and g43645 (n26088, n_17652, n_17653);
  and g43646 (n26089, n26069, n26088);
  not g43647 (n_17654, n26070);
  not g43648 (n_17655, n26089);
  and g43649 (n26090, n_17654, n_17655);
  not g43650 (n_17656, n26090);
  and g43651 (n26091, \a[2] , n_17656);
  and g43652 (n26092, n_10, n26090);
  not g43653 (n_17657, n26091);
  not g43654 (n_17658, n26092);
  and g43655 (n26093, n_17657, n_17658);
  not g43656 (n_17659, n26093);
  and g43657 (n26094, n25853, n_17659);
  not g43658 (n_17660, n25842);
  and g43659 (n26095, n25840, n_17660);
  not g43660 (n_17661, n26095);
  and g43661 (n26096, n_17463, n_17661);
  not g43662 (n_17662, n25827);
  and g43663 (n26097, n25825, n_17662);
  not g43664 (n_17663, n26097);
  and g43665 (n26098, n_17443, n_17663);
  not g43666 (n_17664, n25807);
  and g43667 (n26099, n25805, n_17664);
  not g43668 (n_17665, n26099);
  and g43669 (n26100, n_17417, n_17665);
  not g43670 (n_17666, n25787);
  and g43671 (n26101, n25785, n_17666);
  not g43672 (n_17667, n26101);
  and g43673 (n26102, n_17391, n_17667);
  not g43674 (n_17668, n25765);
  and g43675 (n26103, n25763, n_17668);
  not g43676 (n_17669, n26103);
  and g43677 (n26104, n_17364, n_17669);
  not g43678 (n_17670, n25734);
  and g43679 (n26105, n_17670, n25745);
  not g43680 (n_17671, n25746);
  not g43681 (n_17672, n26105);
  and g43682 (n26106, n_17671, n_17672);
  and g43683 (n26107, n_6354, n_14508);
  and g43684 (n26108, n11796, n_15236);
  and g43685 (n26109, n11727, n22399);
  and g43686 (n26110, n11055, n_14508);
  and g43687 (n26111, n11715, n22402);
  not g43688 (n_17673, n26110);
  not g43689 (n_17674, n26111);
  and g43690 (n26112, n_17673, n_17674);
  not g43691 (n_17675, n26109);
  and g43692 (n26113, n_17675, n26112);
  not g43693 (n_17676, n26113);
  and g43694 (n26114, \a[2] , n_17676);
  and g43695 (n26115, n11796, n_14720);
  and g43696 (n26116, n11805, n_14508);
  and g43697 (n26117, n11807, n22402);
  and g43710 (n26124, n25732, n26123);
  not g43711 (n_17683, n26123);
  and g43712 (n26125, n_17335, n_17683);
  and g43713 (n26126, n11727, n22396);
  and g43714 (n26127, n11055, n22402);
  and g43715 (n26128, n11715, n22399);
  and g43721 (n26131, n11057, n22595);
  not g43724 (n_17688, n26132);
  and g43725 (n26133, n_10, n_17688);
  and g43726 (n26134, \a[2] , n26132);
  not g43727 (n_17689, n26133);
  not g43728 (n_17690, n26134);
  and g43729 (n26135, n_17689, n_17690);
  not g43730 (n_17691, n26125);
  not g43731 (n_17692, n26135);
  and g43732 (n26136, n_17691, n_17692);
  not g43733 (n_17693, n26124);
  not g43734 (n_17694, n26136);
  and g43735 (n26137, n_17693, n_17694);
  and g43736 (n26138, n11727, n22393);
  and g43737 (n26139, n11055, n22399);
  and g43738 (n26140, n11715, n22396);
  not g43739 (n_17695, n26139);
  not g43740 (n_17696, n26140);
  and g43741 (n26141, n_17695, n_17696);
  not g43742 (n_17697, n26138);
  and g43743 (n26142, n_17697, n26141);
  and g43744 (n26143, n_6291, n26142);
  and g43745 (n26144, n_14773, n26142);
  not g43746 (n_17698, n26143);
  not g43747 (n_17699, n26144);
  and g43748 (n26145, n_17698, n_17699);
  not g43749 (n_17700, n26145);
  and g43750 (n26146, \a[2] , n_17700);
  and g43751 (n26147, n_10, n26145);
  not g43752 (n_17701, n26146);
  not g43753 (n_17702, n26147);
  and g43754 (n26148, n_17701, n_17702);
  and g43755 (n26149, n26137, n26148);
  not g43756 (n_17703, n25733);
  and g43757 (n26150, n25731, n_17703);
  not g43758 (n_17704, n26150);
  and g43759 (n26151, n_17670, n_17704);
  not g43760 (n_17705, n26149);
  and g43761 (n26152, n_17705, n26151);
  not g43762 (n_17706, n26137);
  not g43763 (n_17707, n26148);
  and g43764 (n26153, n_17706, n_17707);
  not g43765 (n_17708, n26152);
  not g43766 (n_17709, n26153);
  and g43767 (n26154, n_17708, n_17709);
  not g43768 (n_17710, n26154);
  and g43769 (n26155, n26106, n_17710);
  not g43770 (n_17711, n26106);
  and g43771 (n26156, n_17711, n26154);
  and g43772 (n26157, n11727, n22390);
  and g43773 (n26158, n11055, n22396);
  and g43774 (n26159, n11715, n22393);
  and g43780 (n26162, n11057, n22649);
  not g43783 (n_17716, n26163);
  and g43784 (n26164, n_10, n_17716);
  and g43785 (n26165, \a[2] , n26163);
  not g43786 (n_17717, n26164);
  not g43787 (n_17718, n26165);
  and g43788 (n26166, n_17717, n_17718);
  not g43789 (n_17719, n26156);
  not g43790 (n_17720, n26166);
  and g43791 (n26167, n_17719, n_17720);
  not g43792 (n_17721, n26155);
  not g43793 (n_17722, n26167);
  and g43794 (n26168, n_17721, n_17722);
  and g43795 (n26169, n11727, n22387);
  and g43796 (n26170, n11055, n22393);
  and g43797 (n26171, n11715, n22390);
  not g43798 (n_17723, n26170);
  not g43799 (n_17724, n26171);
  and g43800 (n26172, n_17723, n_17724);
  not g43801 (n_17725, n26169);
  and g43802 (n26173, n_17725, n26172);
  and g43803 (n26174, n_6291, n26173);
  and g43804 (n26175, n_14920, n26173);
  not g43805 (n_17726, n26174);
  not g43806 (n_17727, n26175);
  and g43807 (n26176, n_17726, n_17727);
  not g43808 (n_17728, n26176);
  and g43809 (n26177, \a[2] , n_17728);
  and g43810 (n26178, n_10, n26176);
  not g43811 (n_17729, n26177);
  not g43812 (n_17730, n26178);
  and g43813 (n26179, n_17729, n_17730);
  not g43814 (n_17731, n26168);
  not g43815 (n_17732, n26179);
  and g43816 (n26180, n_17731, n_17732);
  and g43817 (n26181, n26168, n26179);
  and g43818 (n26182, n25750, n25761);
  not g43819 (n_17733, n26182);
  and g43820 (n26183, n_17359, n_17733);
  not g43821 (n_17734, n26181);
  and g43822 (n26184, n_17734, n26183);
  not g43823 (n_17735, n26180);
  not g43824 (n_17736, n26184);
  and g43825 (n26185, n_17735, n_17736);
  not g43826 (n_17737, n26185);
  and g43827 (n26186, n26104, n_17737);
  not g43828 (n_17738, n26104);
  and g43829 (n26187, n_17738, n26185);
  and g43830 (n26188, n11727, n22384);
  and g43831 (n26189, n11055, n22390);
  and g43832 (n26190, n11715, n22387);
  and g43838 (n26193, n11057, n22806);
  not g43841 (n_17743, n26194);
  and g43842 (n26195, n_10, n_17743);
  and g43843 (n26196, \a[2] , n26194);
  not g43844 (n_17744, n26195);
  not g43845 (n_17745, n26196);
  and g43846 (n26197, n_17744, n_17745);
  not g43847 (n_17746, n26187);
  not g43848 (n_17747, n26197);
  and g43849 (n26198, n_17746, n_17747);
  not g43850 (n_17748, n26186);
  not g43851 (n_17749, n26198);
  and g43852 (n26199, n_17748, n_17749);
  and g43853 (n26200, n11727, n22380);
  and g43854 (n26201, n11055, n22387);
  and g43855 (n26202, n11715, n22384);
  not g43856 (n_17750, n26201);
  not g43857 (n_17751, n26202);
  and g43858 (n26203, n_17750, n_17751);
  not g43859 (n_17752, n26200);
  and g43860 (n26204, n_17752, n26203);
  and g43861 (n26205, n_6291, n26204);
  and g43862 (n26206, n_14894, n26204);
  not g43863 (n_17753, n26205);
  not g43864 (n_17754, n26206);
  and g43865 (n26207, n_17753, n_17754);
  not g43866 (n_17755, n26207);
  and g43867 (n26208, \a[2] , n_17755);
  and g43868 (n26209, n_10, n26207);
  not g43869 (n_17756, n26208);
  not g43870 (n_17757, n26209);
  and g43871 (n26210, n_17756, n_17757);
  and g43872 (n26211, n26199, n26210);
  and g43873 (n26212, n25708, n25767);
  not g43874 (n_17758, n26212);
  and g43875 (n26213, n_17367, n_17758);
  not g43876 (n_17759, n26211);
  and g43877 (n26214, n_17759, n26213);
  not g43878 (n_17760, n26199);
  not g43879 (n_17761, n26210);
  and g43880 (n26215, n_17760, n_17761);
  not g43881 (n_17762, n26214);
  not g43882 (n_17763, n26215);
  and g43883 (n26216, n_17762, n_17763);
  and g43884 (n26217, n11727, n22377);
  and g43885 (n26218, n11055, n22384);
  and g43886 (n26219, n11715, n22380);
  not g43887 (n_17764, n26218);
  not g43888 (n_17765, n26219);
  and g43889 (n26220, n_17764, n_17765);
  not g43890 (n_17766, n26217);
  and g43891 (n26221, n_17766, n26220);
  and g43892 (n26222, n_6291, n26221);
  and g43893 (n26223, n22834, n26221);
  not g43894 (n_17767, n26222);
  not g43895 (n_17768, n26223);
  and g43896 (n26224, n_17767, n_17768);
  not g43897 (n_17769, n26224);
  and g43898 (n26225, \a[2] , n_17769);
  and g43899 (n26226, n_10, n26224);
  not g43900 (n_17770, n26225);
  not g43901 (n_17771, n26226);
  and g43902 (n26227, n_17770, n_17771);
  and g43903 (n26228, n26216, n26227);
  not g43904 (n_17772, n25771);
  and g43905 (n26229, n25769, n_17772);
  not g43906 (n_17773, n26229);
  and g43907 (n26230, n_17371, n_17773);
  not g43908 (n_17774, n26228);
  and g43909 (n26231, n_17774, n26230);
  not g43910 (n_17775, n26216);
  not g43911 (n_17776, n26227);
  and g43912 (n26232, n_17775, n_17776);
  not g43913 (n_17777, n26231);
  not g43914 (n_17778, n26232);
  and g43915 (n26233, n_17777, n_17778);
  and g43916 (n26234, n11727, n22374);
  and g43917 (n26235, n11055, n22380);
  and g43918 (n26236, n11715, n22377);
  not g43919 (n_17779, n26235);
  not g43920 (n_17780, n26236);
  and g43921 (n26237, n_17779, n_17780);
  not g43922 (n_17781, n26234);
  and g43923 (n26238, n_17781, n26237);
  and g43924 (n26239, n_6291, n26238);
  and g43925 (n26240, n_15064, n26238);
  not g43926 (n_17782, n26239);
  not g43927 (n_17783, n26240);
  and g43928 (n26241, n_17782, n_17783);
  not g43929 (n_17784, n26241);
  and g43930 (n26242, \a[2] , n_17784);
  and g43931 (n26243, n_10, n26241);
  not g43932 (n_17785, n26242);
  not g43933 (n_17786, n26243);
  and g43934 (n26244, n_17785, n_17786);
  and g43935 (n26245, n26233, n26244);
  and g43936 (n26246, n25676, n25773);
  not g43937 (n_17787, n26246);
  and g43938 (n26247, n_17374, n_17787);
  not g43939 (n_17788, n26245);
  and g43940 (n26248, n_17788, n26247);
  not g43941 (n_17789, n26233);
  not g43942 (n_17790, n26244);
  and g43943 (n26249, n_17789, n_17790);
  not g43944 (n_17791, n26248);
  not g43945 (n_17792, n26249);
  and g43946 (n26250, n_17791, n_17792);
  and g43947 (n26251, n25775, n_17377);
  and g43948 (n26252, n_17376, n26251);
  not g43949 (n_17793, n26252);
  and g43950 (n26253, n_17380, n_17793);
  not g43951 (n_17794, n26250);
  and g43952 (n26254, n_17794, n26253);
  not g43953 (n_17795, n26253);
  and g43954 (n26255, n26250, n_17795);
  and g43955 (n26256, n11727, n22371);
  and g43956 (n26257, n11055, n22377);
  and g43957 (n26258, n11715, n22374);
  and g43963 (n26261, n11057, n23025);
  not g43966 (n_17800, n26262);
  and g43967 (n26263, n_10, n_17800);
  and g43968 (n26264, \a[2] , n26262);
  not g43969 (n_17801, n26263);
  not g43970 (n_17802, n26264);
  and g43971 (n26265, n_17801, n_17802);
  not g43972 (n_17803, n26255);
  not g43973 (n_17804, n26265);
  and g43974 (n26266, n_17803, n_17804);
  not g43975 (n_17805, n26254);
  not g43976 (n_17806, n26266);
  and g43977 (n26267, n_17805, n_17806);
  and g43978 (n26268, n25780, n_17383);
  and g43979 (n26269, n_17382, n26268);
  not g43980 (n_17807, n26269);
  and g43981 (n26270, n_17386, n_17807);
  not g43982 (n_17808, n26267);
  and g43983 (n26271, n_17808, n26270);
  not g43984 (n_17809, n26270);
  and g43985 (n26272, n26267, n_17809);
  and g43986 (n26273, n11727, n22368);
  and g43987 (n26274, n11055, n22374);
  and g43988 (n26275, n11715, n22371);
  and g43994 (n26278, n11057, n23006);
  not g43997 (n_17814, n26279);
  and g43998 (n26280, n_10, n_17814);
  and g43999 (n26281, \a[2] , n26279);
  not g44000 (n_17815, n26280);
  not g44001 (n_17816, n26281);
  and g44002 (n26282, n_17815, n_17816);
  not g44003 (n_17817, n26272);
  not g44004 (n_17818, n26282);
  and g44005 (n26283, n_17817, n_17818);
  not g44006 (n_17819, n26271);
  not g44007 (n_17820, n26283);
  and g44008 (n26284, n_17819, n_17820);
  not g44009 (n_17821, n26284);
  and g44010 (n26285, n26102, n_17821);
  not g44011 (n_17822, n26102);
  and g44012 (n26286, n_17822, n26284);
  and g44013 (n26287, n11727, n22365);
  and g44014 (n26288, n11055, n22371);
  and g44015 (n26289, n11715, n22368);
  and g44021 (n26292, n11057, n_15351);
  not g44024 (n_17827, n26293);
  and g44025 (n26294, n_10, n_17827);
  and g44026 (n26295, \a[2] , n26293);
  not g44027 (n_17828, n26294);
  not g44028 (n_17829, n26295);
  and g44029 (n26296, n_17828, n_17829);
  not g44030 (n_17830, n26286);
  not g44031 (n_17831, n26296);
  and g44032 (n26297, n_17830, n_17831);
  not g44033 (n_17832, n26285);
  not g44034 (n_17833, n26297);
  and g44035 (n26298, n_17832, n_17833);
  and g44036 (n26299, n11727, n22362);
  and g44037 (n26300, n11055, n22368);
  and g44038 (n26301, n11715, n22365);
  not g44039 (n_17834, n26300);
  not g44040 (n_17835, n26301);
  and g44041 (n26302, n_17834, n_17835);
  not g44042 (n_17836, n26299);
  and g44043 (n26303, n_17836, n26302);
  and g44044 (n26304, n_6291, n26303);
  and g44045 (n26305, n23320, n26303);
  not g44046 (n_17837, n26304);
  not g44047 (n_17838, n26305);
  and g44048 (n26306, n_17837, n_17838);
  not g44049 (n_17839, n26306);
  and g44050 (n26307, \a[2] , n_17839);
  and g44051 (n26308, n_10, n26306);
  not g44052 (n_17840, n26307);
  not g44053 (n_17841, n26308);
  and g44054 (n26309, n_17840, n_17841);
  and g44055 (n26310, n26298, n26309);
  and g44056 (n26311, n25617, n25789);
  not g44057 (n_17842, n26311);
  and g44058 (n26312, n_17394, n_17842);
  not g44059 (n_17843, n26310);
  and g44060 (n26313, n_17843, n26312);
  not g44061 (n_17844, n26298);
  not g44062 (n_17845, n26309);
  and g44063 (n26314, n_17844, n_17845);
  not g44064 (n_17846, n26313);
  not g44065 (n_17847, n26314);
  and g44066 (n26315, n_17846, n_17847);
  and g44067 (n26316, n11727, n22359);
  and g44068 (n26317, n11055, n22365);
  and g44069 (n26318, n11715, n22362);
  not g44070 (n_17848, n26317);
  not g44071 (n_17849, n26318);
  and g44072 (n26319, n_17848, n_17849);
  not g44073 (n_17850, n26316);
  and g44074 (n26320, n_17850, n26319);
  and g44075 (n26321, n_6291, n26320);
  and g44076 (n26322, n_15331, n26320);
  not g44077 (n_17851, n26321);
  not g44078 (n_17852, n26322);
  and g44079 (n26323, n_17851, n_17852);
  not g44080 (n_17853, n26323);
  and g44081 (n26324, \a[2] , n_17853);
  and g44082 (n26325, n_10, n26323);
  not g44083 (n_17854, n26324);
  not g44084 (n_17855, n26325);
  and g44085 (n26326, n_17854, n_17855);
  and g44086 (n26327, n26315, n26326);
  and g44087 (n26328, n25599, n25791);
  not g44088 (n_17856, n26328);
  and g44089 (n26329, n_17397, n_17856);
  not g44090 (n_17857, n26327);
  and g44091 (n26330, n_17857, n26329);
  not g44092 (n_17858, n26315);
  not g44093 (n_17859, n26326);
  and g44094 (n26331, n_17858, n_17859);
  not g44095 (n_17860, n26330);
  not g44096 (n_17861, n26331);
  and g44097 (n26332, n_17860, n_17861);
  and g44098 (n26333, n11727, n22356);
  and g44099 (n26334, n11055, n22362);
  and g44100 (n26335, n11715, n22359);
  not g44101 (n_17862, n26334);
  not g44102 (n_17863, n26335);
  and g44103 (n26336, n_17862, n_17863);
  not g44104 (n_17864, n26333);
  and g44105 (n26337, n_17864, n26336);
  and g44106 (n26338, n_6291, n26337);
  and g44107 (n26339, n23345, n26337);
  not g44108 (n_17865, n26338);
  not g44109 (n_17866, n26339);
  and g44110 (n26340, n_17865, n_17866);
  not g44111 (n_17867, n26340);
  and g44112 (n26341, \a[2] , n_17867);
  and g44113 (n26342, n_10, n26340);
  not g44114 (n_17868, n26341);
  not g44115 (n_17869, n26342);
  and g44116 (n26343, n_17868, n_17869);
  and g44117 (n26344, n26332, n26343);
  and g44118 (n26345, n25581, n25793);
  not g44119 (n_17870, n26345);
  and g44120 (n26346, n_17400, n_17870);
  not g44121 (n_17871, n26344);
  and g44122 (n26347, n_17871, n26346);
  not g44123 (n_17872, n26332);
  not g44124 (n_17873, n26343);
  and g44125 (n26348, n_17872, n_17873);
  not g44126 (n_17874, n26347);
  not g44127 (n_17875, n26348);
  and g44128 (n26349, n_17874, n_17875);
  and g44129 (n26350, n25795, n_17403);
  and g44130 (n26351, n_17402, n26350);
  not g44131 (n_17876, n26351);
  and g44132 (n26352, n_17406, n_17876);
  not g44133 (n_17877, n26349);
  and g44134 (n26353, n_17877, n26352);
  not g44135 (n_17878, n26352);
  and g44136 (n26354, n26349, n_17878);
  and g44137 (n26355, n11727, n22353);
  and g44138 (n26356, n11055, n22359);
  and g44139 (n26357, n11715, n22356);
  and g44145 (n26360, n11057, n_14678);
  not g44148 (n_17883, n26361);
  and g44149 (n26362, n_10, n_17883);
  and g44150 (n26363, \a[2] , n26361);
  not g44151 (n_17884, n26362);
  not g44152 (n_17885, n26363);
  and g44153 (n26364, n_17884, n_17885);
  not g44154 (n_17886, n26354);
  not g44155 (n_17887, n26364);
  and g44156 (n26365, n_17886, n_17887);
  not g44157 (n_17888, n26353);
  not g44158 (n_17889, n26365);
  and g44159 (n26366, n_17888, n_17889);
  and g44160 (n26367, n25800, n_17409);
  and g44161 (n26368, n_17408, n26367);
  not g44162 (n_17890, n26368);
  and g44163 (n26369, n_17412, n_17890);
  not g44164 (n_17891, n26366);
  and g44165 (n26370, n_17891, n26369);
  not g44166 (n_17892, n26369);
  and g44167 (n26371, n26366, n_17892);
  and g44168 (n26372, n11727, n22350);
  and g44169 (n26373, n11055, n22356);
  and g44170 (n26374, n11715, n22353);
  and g44176 (n26377, n11057, n23672);
  not g44179 (n_17897, n26378);
  and g44180 (n26379, n_10, n_17897);
  and g44181 (n26380, \a[2] , n26378);
  not g44182 (n_17898, n26379);
  not g44183 (n_17899, n26380);
  and g44184 (n26381, n_17898, n_17899);
  not g44185 (n_17900, n26371);
  not g44186 (n_17901, n26381);
  and g44187 (n26382, n_17900, n_17901);
  not g44188 (n_17902, n26370);
  not g44189 (n_17903, n26382);
  and g44190 (n26383, n_17902, n_17903);
  not g44191 (n_17904, n26383);
  and g44192 (n26384, n26100, n_17904);
  not g44193 (n_17905, n26100);
  and g44194 (n26385, n_17905, n26383);
  and g44195 (n26386, n11727, n22347);
  and g44196 (n26387, n11055, n22353);
  and g44197 (n26388, n11715, n22350);
  and g44203 (n26391, n11057, n_16069);
  not g44206 (n_17910, n26392);
  and g44207 (n26393, n_10, n_17910);
  and g44208 (n26394, \a[2] , n26392);
  not g44209 (n_17911, n26393);
  not g44210 (n_17912, n26394);
  and g44211 (n26395, n_17911, n_17912);
  not g44212 (n_17913, n26385);
  not g44213 (n_17914, n26395);
  and g44214 (n26396, n_17913, n_17914);
  not g44215 (n_17915, n26384);
  not g44216 (n_17916, n26396);
  and g44217 (n26397, n_17915, n_17916);
  and g44218 (n26398, n11727, n22344);
  and g44219 (n26399, n11055, n22350);
  and g44220 (n26400, n11715, n22347);
  not g44221 (n_17917, n26399);
  not g44222 (n_17918, n26400);
  and g44223 (n26401, n_17917, n_17918);
  not g44224 (n_17919, n26398);
  and g44225 (n26402, n_17919, n26401);
  and g44226 (n26403, n_6291, n26402);
  and g44227 (n26404, n23642, n26402);
  not g44228 (n_17920, n26403);
  not g44229 (n_17921, n26404);
  and g44230 (n26405, n_17920, n_17921);
  not g44231 (n_17922, n26405);
  and g44232 (n26406, \a[2] , n_17922);
  and g44233 (n26407, n_10, n26405);
  not g44234 (n_17923, n26406);
  not g44235 (n_17924, n26407);
  and g44236 (n26408, n_17923, n_17924);
  and g44237 (n26409, n26397, n26408);
  and g44238 (n26410, n25522, n25809);
  not g44239 (n_17925, n26410);
  and g44240 (n26411, n_17420, n_17925);
  not g44241 (n_17926, n26409);
  and g44242 (n26412, n_17926, n26411);
  not g44243 (n_17927, n26397);
  not g44244 (n_17928, n26408);
  and g44245 (n26413, n_17927, n_17928);
  not g44246 (n_17929, n26412);
  not g44247 (n_17930, n26413);
  and g44248 (n26414, n_17929, n_17930);
  and g44249 (n26415, n11727, n22341);
  and g44250 (n26416, n11055, n22347);
  and g44251 (n26417, n11715, n22344);
  not g44252 (n_17931, n26416);
  not g44253 (n_17932, n26417);
  and g44254 (n26418, n_17931, n_17932);
  not g44255 (n_17933, n26415);
  and g44256 (n26419, n_17933, n26418);
  and g44257 (n26420, n_6291, n26419);
  and g44258 (n26421, n_15990, n26419);
  not g44259 (n_17934, n26420);
  not g44260 (n_17935, n26421);
  and g44261 (n26422, n_17934, n_17935);
  not g44262 (n_17936, n26422);
  and g44263 (n26423, \a[2] , n_17936);
  and g44264 (n26424, n_10, n26422);
  not g44265 (n_17937, n26423);
  not g44266 (n_17938, n26424);
  and g44267 (n26425, n_17937, n_17938);
  and g44268 (n26426, n26414, n26425);
  and g44269 (n26427, n25504, n25811);
  not g44270 (n_17939, n26427);
  and g44271 (n26428, n_17423, n_17939);
  not g44272 (n_17940, n26426);
  and g44273 (n26429, n_17940, n26428);
  not g44274 (n_17941, n26414);
  not g44275 (n_17942, n26425);
  and g44276 (n26430, n_17941, n_17942);
  not g44277 (n_17943, n26429);
  not g44278 (n_17944, n26430);
  and g44279 (n26431, n_17943, n_17944);
  and g44280 (n26432, n11727, n22338);
  and g44281 (n26433, n11055, n22344);
  and g44282 (n26434, n11715, n22341);
  not g44283 (n_17945, n26433);
  not g44284 (n_17946, n26434);
  and g44285 (n26435, n_17945, n_17946);
  not g44286 (n_17947, n26432);
  and g44287 (n26436, n_17947, n26435);
  and g44288 (n26437, n_6291, n26436);
  and g44289 (n26438, n24188, n26436);
  not g44290 (n_17948, n26437);
  not g44291 (n_17949, n26438);
  and g44292 (n26439, n_17948, n_17949);
  not g44293 (n_17950, n26439);
  and g44294 (n26440, \a[2] , n_17950);
  and g44295 (n26441, n_10, n26439);
  not g44296 (n_17951, n26440);
  not g44297 (n_17952, n26441);
  and g44298 (n26442, n_17951, n_17952);
  and g44299 (n26443, n26431, n26442);
  and g44300 (n26444, n25486, n25813);
  not g44301 (n_17953, n26444);
  and g44302 (n26445, n_17426, n_17953);
  not g44303 (n_17954, n26443);
  and g44304 (n26446, n_17954, n26445);
  not g44305 (n_17955, n26431);
  not g44306 (n_17956, n26442);
  and g44307 (n26447, n_17955, n_17956);
  not g44308 (n_17957, n26446);
  not g44309 (n_17958, n26447);
  and g44310 (n26448, n_17957, n_17958);
  and g44311 (n26449, n25815, n_17429);
  and g44312 (n26450, n_17428, n26449);
  not g44313 (n_17959, n26450);
  and g44314 (n26451, n_17432, n_17959);
  not g44315 (n_17960, n26448);
  and g44316 (n26452, n_17960, n26451);
  not g44317 (n_17961, n26451);
  and g44318 (n26453, n26448, n_17961);
  and g44319 (n26454, n11727, n22335);
  and g44320 (n26455, n11055, n22341);
  and g44321 (n26456, n11715, n22338);
  and g44327 (n26459, n11057, n_16015);
  not g44330 (n_17966, n26460);
  and g44331 (n26461, n_10, n_17966);
  and g44332 (n26462, \a[2] , n26460);
  not g44333 (n_17967, n26461);
  not g44334 (n_17968, n26462);
  and g44335 (n26463, n_17967, n_17968);
  not g44336 (n_17969, n26453);
  not g44337 (n_17970, n26463);
  and g44338 (n26464, n_17969, n_17970);
  not g44339 (n_17971, n26452);
  not g44340 (n_17972, n26464);
  and g44341 (n26465, n_17971, n_17972);
  and g44342 (n26466, n25820, n_17435);
  and g44343 (n26467, n_17434, n26466);
  not g44344 (n_17973, n26467);
  and g44345 (n26468, n_17438, n_17973);
  not g44346 (n_17974, n26465);
  and g44347 (n26469, n_17974, n26468);
  not g44348 (n_17975, n26468);
  and g44349 (n26470, n26465, n_17975);
  and g44350 (n26471, n11727, n22332);
  and g44351 (n26472, n11055, n22338);
  and g44352 (n26473, n11715, n22335);
  and g44358 (n26476, n11057, n22542);
  not g44361 (n_17980, n26477);
  and g44362 (n26478, n_10, n_17980);
  and g44363 (n26479, \a[2] , n26477);
  not g44364 (n_17981, n26478);
  not g44365 (n_17982, n26479);
  and g44366 (n26480, n_17981, n_17982);
  not g44367 (n_17983, n26470);
  not g44368 (n_17984, n26480);
  and g44369 (n26481, n_17983, n_17984);
  not g44370 (n_17985, n26469);
  not g44371 (n_17986, n26481);
  and g44372 (n26482, n_17985, n_17986);
  not g44373 (n_17987, n26482);
  and g44374 (n26483, n26098, n_17987);
  not g44375 (n_17988, n26098);
  and g44376 (n26484, n_17988, n26482);
  and g44377 (n26485, n11727, n22329);
  and g44378 (n26486, n11055, n22335);
  and g44379 (n26487, n11715, n22332);
  and g44385 (n26490, n11057, n_16827);
  not g44388 (n_17993, n26491);
  and g44389 (n26492, n_10, n_17993);
  and g44390 (n26493, \a[2] , n26491);
  not g44391 (n_17994, n26492);
  not g44392 (n_17995, n26493);
  and g44393 (n26494, n_17994, n_17995);
  not g44394 (n_17996, n26484);
  not g44395 (n_17997, n26494);
  and g44396 (n26495, n_17996, n_17997);
  not g44397 (n_17998, n26483);
  not g44398 (n_17999, n26495);
  and g44399 (n26496, n_17998, n_17999);
  and g44400 (n26497, n11727, n22326);
  and g44401 (n26498, n11055, n22332);
  and g44402 (n26499, n11715, n22329);
  not g44403 (n_18000, n26498);
  not g44404 (n_18001, n26499);
  and g44405 (n26500, n_18000, n_18001);
  not g44406 (n_18002, n26497);
  and g44407 (n26501, n_18002, n26500);
  and g44408 (n26502, n_6291, n26501);
  and g44409 (n26503, n24616, n26501);
  not g44410 (n_18003, n26502);
  not g44411 (n_18004, n26503);
  and g44412 (n26504, n_18003, n_18004);
  not g44413 (n_18005, n26504);
  and g44414 (n26505, \a[2] , n_18005);
  and g44415 (n26506, n_10, n26504);
  not g44416 (n_18006, n26505);
  not g44417 (n_18007, n26506);
  and g44418 (n26507, n_18006, n_18007);
  and g44419 (n26508, n26496, n26507);
  and g44420 (n26509, n25427, n25829);
  not g44421 (n_18008, n26509);
  and g44422 (n26510, n_17446, n_18008);
  not g44423 (n_18009, n26508);
  and g44424 (n26511, n_18009, n26510);
  not g44425 (n_18010, n26496);
  not g44426 (n_18011, n26507);
  and g44427 (n26512, n_18010, n_18011);
  not g44428 (n_18012, n26511);
  not g44429 (n_18013, n26512);
  and g44430 (n26513, n_18012, n_18013);
  and g44431 (n26514, n11727, n22323);
  and g44432 (n26515, n11055, n22329);
  and g44433 (n26516, n11715, n22326);
  not g44434 (n_18014, n26515);
  not g44435 (n_18015, n26516);
  and g44436 (n26517, n_18014, n_18015);
  not g44437 (n_18016, n26514);
  and g44438 (n26518, n_18016, n26517);
  and g44439 (n26519, n_6291, n26518);
  and g44440 (n26520, n_16393, n26518);
  not g44441 (n_18017, n26519);
  not g44442 (n_18018, n26520);
  and g44443 (n26521, n_18017, n_18018);
  not g44444 (n_18019, n26521);
  and g44445 (n26522, \a[2] , n_18019);
  and g44446 (n26523, n_10, n26521);
  not g44447 (n_18020, n26522);
  not g44448 (n_18021, n26523);
  and g44449 (n26524, n_18020, n_18021);
  and g44450 (n26525, n26513, n26524);
  and g44451 (n26526, n25409, n25831);
  not g44452 (n_18022, n26526);
  and g44453 (n26527, n_17449, n_18022);
  not g44454 (n_18023, n26525);
  and g44455 (n26528, n_18023, n26527);
  not g44456 (n_18024, n26513);
  not g44457 (n_18025, n26524);
  and g44458 (n26529, n_18024, n_18025);
  not g44459 (n_18026, n26528);
  not g44460 (n_18027, n26529);
  and g44461 (n26530, n_18026, n_18027);
  and g44462 (n26531, n11727, n22320);
  and g44463 (n26532, n11055, n22326);
  and g44464 (n26533, n11715, n22323);
  not g44465 (n_18028, n26532);
  not g44466 (n_18029, n26533);
  and g44467 (n26534, n_18028, n_18029);
  not g44468 (n_18030, n26531);
  and g44469 (n26535, n_18030, n26534);
  and g44470 (n26536, n_6291, n26535);
  and g44471 (n26537, n25270, n26535);
  not g44472 (n_18031, n26536);
  not g44473 (n_18032, n26537);
  and g44474 (n26538, n_18031, n_18032);
  not g44475 (n_18033, n26538);
  and g44476 (n26539, \a[2] , n_18033);
  and g44477 (n26540, n_10, n26538);
  not g44478 (n_18034, n26539);
  not g44479 (n_18035, n26540);
  and g44480 (n26541, n_18034, n_18035);
  and g44481 (n26542, n26530, n26541);
  and g44482 (n26543, n25391, n25833);
  not g44483 (n_18036, n26543);
  and g44484 (n26544, n_17452, n_18036);
  not g44485 (n_18037, n26542);
  and g44486 (n26545, n_18037, n26544);
  not g44487 (n_18038, n26530);
  not g44488 (n_18039, n26541);
  and g44489 (n26546, n_18038, n_18039);
  not g44490 (n_18040, n26545);
  not g44491 (n_18041, n26546);
  and g44492 (n26547, n_18040, n_18041);
  and g44493 (n26548, n25835, n_17455);
  and g44494 (n26549, n_17454, n26548);
  not g44495 (n_18042, n26549);
  and g44496 (n26550, n_17458, n_18042);
  not g44497 (n_18043, n26547);
  and g44498 (n26551, n_18043, n26550);
  not g44499 (n_18044, n26550);
  and g44500 (n26552, n26547, n_18044);
  and g44501 (n26553, n11727, n22312);
  and g44502 (n26554, n11055, n22323);
  and g44503 (n26555, n11715, n22320);
  and g44509 (n26558, n11057, n_17004);
  not g44512 (n_18049, n26559);
  and g44513 (n26560, n_10, n_18049);
  and g44514 (n26561, \a[2] , n26559);
  not g44515 (n_18050, n26560);
  not g44516 (n_18051, n26561);
  and g44517 (n26562, n_18050, n_18051);
  not g44518 (n_18052, n26552);
  not g44519 (n_18053, n26562);
  and g44520 (n26563, n_18052, n_18053);
  not g44521 (n_18054, n26551);
  not g44522 (n_18055, n26563);
  and g44523 (n26564, n_18054, n_18055);
  not g44524 (n_18056, n26564);
  and g44525 (n26565, n26096, n_18056);
  not g44526 (n_18057, n26096);
  and g44527 (n26566, n_18057, n26564);
  and g44528 (n26567, n11727, n22315);
  and g44529 (n26568, n11055, n22320);
  and g44530 (n26569, n11715, n22312);
  and g44536 (n26572, n11057, n25294);
  not g44539 (n_18062, n26573);
  and g44540 (n26574, n_10, n_18062);
  and g44541 (n26575, \a[2] , n26573);
  not g44542 (n_18063, n26574);
  not g44543 (n_18064, n26575);
  and g44544 (n26576, n_18063, n_18064);
  not g44545 (n_18065, n26566);
  not g44546 (n_18066, n26576);
  and g44547 (n26577, n_18065, n_18066);
  not g44548 (n_18067, n26565);
  not g44549 (n_18068, n26577);
  and g44550 (n26578, n_18067, n_18068);
  and g44551 (n26579, n11727, n22309);
  and g44552 (n26580, n11055, n22312);
  and g44553 (n26581, n11715, n22315);
  not g44554 (n_18069, n26580);
  not g44555 (n_18070, n26581);
  and g44556 (n26582, n_18069, n_18070);
  not g44557 (n_18071, n26579);
  and g44558 (n26583, n_18071, n26582);
  and g44559 (n26584, n_6291, n26583);
  and g44560 (n26585, n22529, n26583);
  not g44561 (n_18072, n26584);
  not g44562 (n_18073, n26585);
  and g44563 (n26586, n_18072, n_18073);
  not g44564 (n_18074, n26586);
  and g44565 (n26587, \a[2] , n_18074);
  and g44566 (n26588, n_10, n26586);
  not g44567 (n_18075, n26587);
  not g44568 (n_18076, n26588);
  and g44569 (n26589, n_18075, n_18076);
  and g44570 (n26590, n26578, n26589);
  and g44571 (n26591, n25346, n25844);
  not g44572 (n_18077, n26591);
  and g44573 (n26592, n_17466, n_18077);
  not g44574 (n_18078, n26590);
  and g44575 (n26593, n_18078, n26592);
  not g44576 (n_18079, n26578);
  not g44577 (n_18080, n26589);
  and g44578 (n26594, n_18079, n_18080);
  not g44579 (n_18081, n26593);
  not g44580 (n_18082, n26594);
  and g44581 (n26595, n_18081, n_18082);
  and g44582 (n26596, n11727, n26063);
  and g44583 (n26597, n11055, n22315);
  and g44584 (n26598, n11715, n22309);
  not g44585 (n_18083, n26597);
  not g44586 (n_18084, n26598);
  and g44587 (n26599, n_18083, n_18084);
  not g44588 (n_18085, n26596);
  and g44589 (n26600, n_18085, n26599);
  and g44590 (n26601, n_6291, n26600);
  and g44591 (n26602, n_17638, n_17641);
  and g44592 (n26603, n_17639, n26076);
  not g44593 (n_18086, n26602);
  not g44594 (n_18087, n26603);
  and g44595 (n26604, n_18086, n_18087);
  and g44596 (n26605, n26600, n26604);
  not g44597 (n_18088, n26601);
  not g44598 (n_18089, n26605);
  and g44599 (n26606, n_18088, n_18089);
  not g44600 (n_18090, n26606);
  and g44601 (n26607, \a[2] , n_18090);
  and g44602 (n26608, n_10, n26606);
  not g44603 (n_18091, n26607);
  not g44604 (n_18092, n26608);
  and g44605 (n26609, n_18091, n_18092);
  and g44606 (n26610, n26595, n26609);
  and g44607 (n26611, n25328, n25846);
  not g44608 (n_18093, n26611);
  and g44609 (n26612, n_17469, n_18093);
  not g44610 (n_18094, n26610);
  and g44611 (n26613, n_18094, n26612);
  not g44612 (n_18095, n26595);
  not g44613 (n_18096, n26609);
  and g44614 (n26614, n_18095, n_18096);
  not g44615 (n_18097, n26613);
  not g44616 (n_18098, n26614);
  and g44617 (n26615, n_18097, n_18098);
  and g44618 (n26616, n11727, n26066);
  and g44619 (n26617, n11055, n22309);
  and g44620 (n26618, n11715, n26063);
  not g44621 (n_18099, n26617);
  not g44622 (n_18100, n26618);
  and g44623 (n26619, n_18099, n_18100);
  not g44624 (n_18101, n26616);
  and g44625 (n26620, n_18101, n26619);
  and g44626 (n26621, n_6291, n26620);
  and g44627 (n26622, n_17643, n_17646);
  and g44628 (n26623, n_17644, n26080);
  not g44629 (n_18102, n26622);
  not g44630 (n_18103, n26623);
  and g44631 (n26624, n_18102, n_18103);
  and g44632 (n26625, n26620, n26624);
  not g44633 (n_18104, n26621);
  not g44634 (n_18105, n26625);
  and g44635 (n26626, n_18104, n_18105);
  not g44636 (n_18106, n26626);
  and g44637 (n26627, \a[2] , n_18106);
  and g44638 (n26628, n_10, n26626);
  not g44639 (n_18107, n26627);
  not g44640 (n_18108, n26628);
  and g44641 (n26629, n_18107, n_18108);
  and g44642 (n26630, n26615, n26629);
  and g44643 (n26631, n25307, n25848);
  not g44644 (n_18109, n26631);
  and g44645 (n26632, n_17472, n_18109);
  not g44646 (n_18110, n26630);
  and g44647 (n26633, n_18110, n26632);
  not g44648 (n_18111, n26615);
  not g44649 (n_18112, n26629);
  and g44650 (n26634, n_18111, n_18112);
  not g44651 (n_18113, n26633);
  not g44652 (n_18114, n26634);
  and g44653 (n26635, n_18113, n_18114);
  not g44654 (n_18115, n26094);
  and g44655 (n26636, n25853, n_18115);
  and g44656 (n26637, n_17659, n_18115);
  not g44657 (n_18116, n26636);
  not g44658 (n_18117, n26637);
  and g44659 (n26638, n_18116, n_18117);
  not g44660 (n_18118, n26635);
  not g44661 (n_18119, n26638);
  and g44662 (n26639, n_18118, n_18119);
  not g44663 (n_18120, n26639);
  and g44664 (n26640, n_18115, n_18120);
  and g44665 (n26641, n71, n26063);
  and g44666 (n26642, n9867, n22315);
  and g44667 (n26643, n10434, n22309);
  not g44673 (n_18124, n26604);
  and g44674 (n26646, n9870, n_18124);
  not g44677 (n_18126, n26647);
  and g44678 (n26648, \a[5] , n_18126);
  not g44679 (n_18127, n26648);
  and g44680 (n26649, n_18126, n_18127);
  and g44681 (n26650, \a[5] , n_18127);
  not g44682 (n_18128, n26649);
  not g44683 (n_18129, n26650);
  and g44684 (n26651, n_18128, n_18129);
  and g44685 (n26652, n_16969, n_16974);
  and g44686 (n26653, n7983, n22326);
  and g44687 (n26654, n7291, n22332);
  and g44688 (n26655, n7632, n22329);
  not g44694 (n_18133, n24616);
  and g44695 (n26658, n7294, n_18133);
  not g44698 (n_18135, n26659);
  and g44699 (n26660, \a[11] , n_18135);
  not g44700 (n_18136, n26660);
  and g44701 (n26661, n_18135, n_18136);
  and g44702 (n26662, \a[11] , n_18136);
  not g44703 (n_18137, n26661);
  not g44704 (n_18138, n26662);
  and g44705 (n26663, n_18137, n_18138);
  and g44706 (n26664, n_16941, n_16946);
  and g44707 (n26665, n6233, n22344);
  and g44708 (n26666, n5663, n22350);
  and g44709 (n26667, n5939, n22347);
  not g44715 (n_18142, n23642);
  and g44716 (n26670, n5666, n_18142);
  not g44719 (n_18144, n26671);
  and g44720 (n26672, \a[17] , n_18144);
  not g44721 (n_18145, n26672);
  and g44722 (n26673, n_18144, n_18145);
  and g44723 (n26674, \a[17] , n_18145);
  not g44724 (n_18146, n26673);
  not g44725 (n_18147, n26674);
  and g44726 (n26675, n_18146, n_18147);
  and g44727 (n26676, n_16915, n_16920);
  and g44728 (n26677, n4694, n22362);
  and g44729 (n26678, n4533, n22368);
  and g44730 (n26679, n4604, n22365);
  not g44736 (n_18151, n23320);
  and g44737 (n26682, n4536, n_18151);
  not g44740 (n_18153, n26683);
  and g44741 (n26684, \a[23] , n_18153);
  not g44742 (n_18154, n26684);
  and g44743 (n26685, n_18153, n_18154);
  and g44744 (n26686, \a[23] , n_18154);
  not g44745 (n_18155, n26685);
  not g44746 (n_18156, n26686);
  and g44747 (n26687, n_18155, n_18156);
  and g44748 (n26688, n_16889, n_16894);
  and g44749 (n26689, n3457, n22380);
  and g44750 (n26690, n3542, n22387);
  and g44751 (n26691, n3606, n22384);
  and g44757 (n26694, n3368, n22850);
  not g44760 (n_18161, n26695);
  and g44761 (n26696, \a[29] , n_18161);
  not g44762 (n_18162, n26696);
  and g44763 (n26697, n_18161, n_18162);
  and g44764 (n26698, \a[29] , n_18162);
  not g44765 (n_18163, n26697);
  not g44766 (n_18164, n26698);
  and g44767 (n26699, n_18163, n_18164);
  and g44768 (n26700, n_16863, n_16868);
  and g44784 (n26716, n3020, n22390);
  and g44785 (n26717, n3028, n22393);
  and g44786 (n26718, n3023, n22396);
  and g44787 (n26719, n75, n22649);
  not g44795 (n_18169, n26715);
  not g44796 (n_18170, n26722);
  and g44797 (n26723, n_18169, n_18170);
  not g44798 (n_18171, n26723);
  and g44799 (n26724, n_18169, n_18171);
  and g44800 (n26725, n_18170, n_18171);
  not g44801 (n_18172, n26724);
  not g44802 (n_18173, n26725);
  and g44803 (n26726, n_18172, n_18173);
  not g44804 (n_18174, n26700);
  not g44805 (n_18175, n26726);
  and g44806 (n26727, n_18174, n_18175);
  not g44807 (n_18176, n26727);
  and g44808 (n26728, n_18174, n_18176);
  and g44809 (n26729, n_18175, n_18176);
  not g44810 (n_18177, n26728);
  not g44811 (n_18178, n26729);
  and g44812 (n26730, n_18177, n_18178);
  not g44813 (n_18179, n26699);
  not g44814 (n_18180, n26730);
  and g44815 (n26731, n_18179, n_18180);
  not g44816 (n_18181, n26731);
  and g44817 (n26732, n_18179, n_18181);
  and g44818 (n26733, n_18180, n_18181);
  not g44819 (n_18182, n26732);
  not g44820 (n_18183, n26733);
  and g44821 (n26734, n_18182, n_18183);
  and g44822 (n26735, n_16873, n_16879);
  and g44823 (n26736, n26734, n26735);
  not g44824 (n_18184, n26734);
  not g44825 (n_18185, n26735);
  and g44826 (n26737, n_18184, n_18185);
  not g44827 (n_18186, n26736);
  not g44828 (n_18187, n26737);
  and g44829 (n26738, n_18186, n_18187);
  and g44830 (n26739, n3884, n22371);
  and g44831 (n26740, n3967, n22377);
  and g44832 (n26741, n4046, n22374);
  not g44833 (n_18188, n26740);
  not g44834 (n_18189, n26741);
  and g44835 (n26742, n_18188, n_18189);
  not g44836 (n_18190, n26739);
  and g44837 (n26743, n_18190, n26742);
  and g44838 (n26744, n_750, n26743);
  not g44839 (n_18191, n23025);
  and g44840 (n26745, n_18191, n26743);
  not g44841 (n_18192, n26744);
  not g44842 (n_18193, n26745);
  and g44843 (n26746, n_18192, n_18193);
  not g44844 (n_18194, n26746);
  and g44845 (n26747, \a[26] , n_18194);
  and g44846 (n26748, n_33, n26746);
  not g44847 (n_18195, n26747);
  not g44848 (n_18196, n26748);
  and g44849 (n26749, n_18195, n_18196);
  not g44850 (n_18197, n26749);
  and g44851 (n26750, n26738, n_18197);
  not g44852 (n_18198, n26750);
  and g44853 (n26751, n26738, n_18198);
  and g44854 (n26752, n_18197, n_18198);
  not g44855 (n_18199, n26751);
  not g44856 (n_18200, n26752);
  and g44857 (n26753, n_18199, n_18200);
  not g44858 (n_18201, n26688);
  not g44859 (n_18202, n26753);
  and g44860 (n26754, n_18201, n_18202);
  not g44861 (n_18203, n26754);
  and g44862 (n26755, n_18201, n_18203);
  and g44863 (n26756, n_18202, n_18203);
  not g44864 (n_18204, n26755);
  not g44865 (n_18205, n26756);
  and g44866 (n26757, n_18204, n_18205);
  not g44867 (n_18206, n26687);
  not g44868 (n_18207, n26757);
  and g44869 (n26758, n_18206, n_18207);
  not g44870 (n_18208, n26758);
  and g44871 (n26759, n_18206, n_18208);
  and g44872 (n26760, n_18207, n_18208);
  not g44873 (n_18209, n26759);
  not g44874 (n_18210, n26760);
  and g44875 (n26761, n_18209, n_18210);
  and g44876 (n26762, n_16899, n_16905);
  and g44877 (n26763, n26761, n26762);
  not g44878 (n_18211, n26761);
  not g44879 (n_18212, n26762);
  and g44880 (n26764, n_18211, n_18212);
  not g44881 (n_18213, n26763);
  not g44882 (n_18214, n26764);
  and g44883 (n26765, n_18213, n_18214);
  and g44884 (n26766, n5496, n22353);
  and g44885 (n26767, n4935, n22359);
  and g44886 (n26768, n5407, n22356);
  not g44887 (n_18215, n26767);
  not g44888 (n_18216, n26768);
  and g44889 (n26769, n_18215, n_18216);
  not g44890 (n_18217, n26766);
  and g44891 (n26770, n_18217, n26769);
  and g44892 (n26771, n_1011, n26770);
  and g44893 (n26772, n22556, n26770);
  not g44894 (n_18218, n26771);
  not g44895 (n_18219, n26772);
  and g44896 (n26773, n_18218, n_18219);
  not g44897 (n_18220, n26773);
  and g44898 (n26774, \a[20] , n_18220);
  and g44899 (n26775, n_435, n26773);
  not g44900 (n_18221, n26774);
  not g44901 (n_18222, n26775);
  and g44902 (n26776, n_18221, n_18222);
  not g44903 (n_18223, n26776);
  and g44904 (n26777, n26765, n_18223);
  not g44905 (n_18224, n26777);
  and g44906 (n26778, n26765, n_18224);
  and g44907 (n26779, n_18223, n_18224);
  not g44908 (n_18225, n26778);
  not g44909 (n_18226, n26779);
  and g44910 (n26780, n_18225, n_18226);
  not g44911 (n_18227, n26676);
  not g44912 (n_18228, n26780);
  and g44913 (n26781, n_18227, n_18228);
  not g44914 (n_18229, n26781);
  and g44915 (n26782, n_18227, n_18229);
  and g44916 (n26783, n_18228, n_18229);
  not g44917 (n_18230, n26782);
  not g44918 (n_18231, n26783);
  and g44919 (n26784, n_18230, n_18231);
  not g44920 (n_18232, n26675);
  not g44921 (n_18233, n26784);
  and g44922 (n26785, n_18232, n_18233);
  not g44923 (n_18234, n26785);
  and g44924 (n26786, n_18232, n_18234);
  and g44925 (n26787, n_18233, n_18234);
  not g44926 (n_18235, n26786);
  not g44927 (n_18236, n26787);
  and g44928 (n26788, n_18235, n_18236);
  and g44929 (n26789, n_16925, n_16931);
  and g44930 (n26790, n26788, n26789);
  not g44931 (n_18237, n26788);
  not g44932 (n_18238, n26789);
  and g44933 (n26791, n_18237, n_18238);
  not g44934 (n_18239, n26790);
  not g44935 (n_18240, n26791);
  and g44936 (n26792, n_18239, n_18240);
  and g44937 (n26793, n7101, n22335);
  and g44938 (n26794, n6402, n22341);
  and g44939 (n26795, n6951, n22338);
  not g44940 (n_18241, n26794);
  not g44941 (n_18242, n26795);
  and g44942 (n26796, n_18241, n_18242);
  not g44943 (n_18243, n26793);
  and g44944 (n26797, n_18243, n26796);
  and g44945 (n26798, n_1885, n26797);
  and g44946 (n26799, n24167, n26797);
  not g44947 (n_18244, n26798);
  not g44948 (n_18245, n26799);
  and g44949 (n26800, n_18244, n_18245);
  not g44950 (n_18246, n26800);
  and g44951 (n26801, \a[14] , n_18246);
  and g44952 (n26802, n_652, n26800);
  not g44953 (n_18247, n26801);
  not g44954 (n_18248, n26802);
  and g44955 (n26803, n_18247, n_18248);
  not g44956 (n_18249, n26803);
  and g44957 (n26804, n26792, n_18249);
  not g44958 (n_18250, n26804);
  and g44959 (n26805, n26792, n_18250);
  and g44960 (n26806, n_18249, n_18250);
  not g44961 (n_18251, n26805);
  not g44962 (n_18252, n26806);
  and g44963 (n26807, n_18251, n_18252);
  not g44964 (n_18253, n26664);
  not g44965 (n_18254, n26807);
  and g44966 (n26808, n_18253, n_18254);
  not g44967 (n_18255, n26808);
  and g44968 (n26809, n_18253, n_18255);
  and g44969 (n26810, n_18254, n_18255);
  not g44970 (n_18256, n26809);
  not g44971 (n_18257, n26810);
  and g44972 (n26811, n_18256, n_18257);
  not g44973 (n_18258, n26663);
  not g44974 (n_18259, n26811);
  and g44975 (n26812, n_18258, n_18259);
  not g44976 (n_18260, n26812);
  and g44977 (n26813, n_18258, n_18260);
  and g44978 (n26814, n_18259, n_18260);
  not g44979 (n_18261, n26813);
  not g44980 (n_18262, n26814);
  and g44981 (n26815, n_18261, n_18262);
  and g44982 (n26816, n_16951, n_16957);
  and g44983 (n26817, n26815, n26816);
  not g44984 (n_18263, n26815);
  not g44985 (n_18264, n26816);
  and g44986 (n26818, n_18263, n_18264);
  not g44987 (n_18265, n26817);
  not g44988 (n_18266, n26818);
  and g44989 (n26819, n_18265, n_18266);
  and g44990 (n26820, n9331, n22312);
  and g44991 (n26821, n8418, n22323);
  and g44992 (n26822, n8860, n22320);
  not g44993 (n_18267, n26821);
  not g44994 (n_18268, n26822);
  and g44995 (n26823, n_18267, n_18268);
  not g44996 (n_18269, n26820);
  and g44997 (n26824, n_18269, n26823);
  and g44998 (n26825, n_3428, n26824);
  and g44999 (n26826, n25315, n26824);
  not g45000 (n_18270, n26825);
  not g45001 (n_18271, n26826);
  and g45002 (n26827, n_18270, n_18271);
  not g45003 (n_18272, n26827);
  and g45004 (n26828, \a[8] , n_18272);
  and g45005 (n26829, n_1106, n26827);
  not g45006 (n_18273, n26828);
  not g45007 (n_18274, n26829);
  and g45008 (n26830, n_18273, n_18274);
  not g45009 (n_18275, n26830);
  and g45010 (n26831, n26819, n_18275);
  not g45011 (n_18276, n26831);
  and g45012 (n26832, n26819, n_18276);
  and g45013 (n26833, n_18275, n_18276);
  not g45014 (n_18277, n26832);
  not g45015 (n_18278, n26833);
  and g45016 (n26834, n_18277, n_18278);
  not g45017 (n_18279, n26652);
  not g45018 (n_18280, n26834);
  and g45019 (n26835, n_18279, n_18280);
  not g45020 (n_18281, n26835);
  and g45021 (n26836, n_18279, n_18281);
  and g45022 (n26837, n_18280, n_18281);
  not g45023 (n_18282, n26836);
  not g45024 (n_18283, n26837);
  and g45025 (n26838, n_18282, n_18283);
  not g45026 (n_18284, n26651);
  not g45027 (n_18285, n26838);
  and g45028 (n26839, n_18284, n_18285);
  not g45029 (n_18286, n26839);
  and g45030 (n26840, n_18284, n_18286);
  and g45031 (n26841, n_18285, n_18286);
  not g45032 (n_18287, n26840);
  not g45033 (n_18288, n26841);
  and g45034 (n26842, n_18287, n_18288);
  and g45035 (n26843, n_16979, n_17476);
  and g45036 (n26844, n26842, n26843);
  not g45037 (n_18289, n26842);
  not g45038 (n_18290, n26843);
  and g45039 (n26845, n_18289, n_18290);
  not g45040 (n_18291, n26844);
  not g45041 (n_18292, n26845);
  and g45042 (n26846, n_18291, n_18292);
  and g45043 (n26847, n_17625, n_17630);
  and g45044 (n26848, n_17616, n_17622);
  and g45045 (n26849, n75, n13929);
  and g45046 (n26850, n3020, n13633);
  and g45047 (n26851, n3023, n13597);
  and g45048 (n26852, n3028, n13630);
  and g45056 (n26856, n_17593, n_17596);
  not g45060 (n_18297, n26856);
  and g45061 (n26860, n_18297, n26859);
  not g45062 (n_18298, n26859);
  and g45063 (n26861, n26856, n_18298);
  not g45064 (n_18299, n26860);
  not g45065 (n_18300, n26861);
  and g45066 (n26862, n_18299, n_18300);
  not g45067 (n_18301, n26855);
  and g45068 (n26863, n_18301, n26862);
  not g45069 (n_18302, n26863);
  and g45070 (n26864, n_18301, n_18302);
  and g45071 (n26865, n26862, n_18302);
  not g45072 (n_18303, n26864);
  not g45073 (n_18304, n26865);
  and g45074 (n26866, n_18303, n_18304);
  and g45075 (n26867, n_17600, n_17603);
  and g45076 (n26868, n26866, n26867);
  not g45077 (n_18305, n26866);
  not g45078 (n_18306, n26867);
  and g45079 (n26869, n_18305, n_18306);
  not g45080 (n_18307, n26868);
  not g45081 (n_18308, n26869);
  and g45082 (n26870, n_18307, n_18308);
  and g45083 (n26871, n3457, n_7417);
  and g45084 (n26872, n3542, n_7540);
  and g45085 (n26873, n3606, n13941);
  not g45086 (n_18309, n26872);
  not g45087 (n_18310, n26873);
  and g45088 (n26874, n_18309, n_18310);
  not g45089 (n_18311, n26871);
  and g45090 (n26875, n_18311, n26874);
  and g45091 (n26876, n_489, n26875);
  and g45092 (n26877, n_13769, n26875);
  not g45093 (n_18312, n26876);
  not g45094 (n_18313, n26877);
  and g45095 (n26878, n_18312, n_18313);
  not g45096 (n_18314, n26878);
  and g45097 (n26879, \a[29] , n_18314);
  and g45098 (n26880, n_15, n26878);
  not g45099 (n_18315, n26879);
  not g45100 (n_18316, n26880);
  and g45101 (n26881, n_18315, n_18316);
  not g45102 (n_18317, n26881);
  and g45103 (n26882, n26870, n_18317);
  not g45104 (n_18318, n26870);
  and g45105 (n26883, n_18318, n26881);
  not g45106 (n_18319, n26882);
  not g45107 (n_18320, n26883);
  and g45108 (n26884, n_18319, n_18320);
  not g45109 (n_18321, n26848);
  and g45110 (n26885, n_18321, n26884);
  not g45111 (n_18322, n26884);
  and g45112 (n26886, n26848, n_18322);
  not g45113 (n_18323, n26885);
  not g45114 (n_18324, n26886);
  and g45115 (n26887, n_18323, n_18324);
  not g45116 (n_18325, n26847);
  and g45117 (n26888, n_18325, n26887);
  not g45118 (n_18326, n26887);
  and g45119 (n26889, n26847, n_18326);
  not g45120 (n_18327, n26888);
  not g45121 (n_18328, n26889);
  and g45122 (n26890, n_18327, n_18328);
  and g45123 (n26891, n11727, n26890);
  and g45124 (n26892, n11055, n26066);
  and g45125 (n26893, n11715, n26060);
  not g45126 (n_18329, n26892);
  not g45127 (n_18330, n26893);
  and g45128 (n26894, n_18329, n_18330);
  not g45129 (n_18331, n26891);
  and g45130 (n26895, n_18331, n26894);
  and g45131 (n26896, n_6291, n26895);
  and g45132 (n26897, n26060, n26890);
  not g45133 (n_18332, n26890);
  and g45134 (n26898, n_17647, n_18332);
  not g45135 (n_18333, n26086);
  not g45136 (n_18334, n26898);
  and g45137 (n26899, n_18333, n_18334);
  not g45138 (n_18335, n26897);
  and g45139 (n26900, n_18335, n26899);
  not g45140 (n_18336, n26900);
  and g45141 (n26901, n_18333, n_18336);
  and g45142 (n26902, n_18335, n_18336);
  and g45143 (n26903, n_18334, n26902);
  not g45144 (n_18337, n26901);
  not g45145 (n_18338, n26903);
  and g45146 (n26904, n_18337, n_18338);
  and g45147 (n26905, n26895, n26904);
  not g45148 (n_18339, n26896);
  not g45149 (n_18340, n26905);
  and g45150 (n26906, n_18339, n_18340);
  not g45151 (n_18341, n26906);
  and g45152 (n26907, \a[2] , n_18341);
  and g45153 (n26908, n_10, n26906);
  not g45154 (n_18342, n26907);
  not g45155 (n_18343, n26908);
  and g45156 (n26909, n_18342, n_18343);
  not g45157 (n_18344, n26909);
  and g45158 (n26910, n26846, n_18344);
  not g45159 (n_18345, n26846);
  and g45160 (n26911, n_18345, n26909);
  not g45161 (n_18346, n26910);
  not g45162 (n_18347, n26911);
  and g45163 (n26912, n_18346, n_18347);
  not g45164 (n_18348, n26640);
  and g45165 (n26913, n_18348, n26912);
  not g45166 (n_18349, n26912);
  and g45167 (n26914, n26640, n_18349);
  not g45168 (n_18350, n26913);
  not g45169 (n_18351, n26914);
  and g45170 (n26915, n_18350, n_18351);
  and g45171 (n26916, n_18118, n_18120);
  and g45172 (n26917, n_18119, n_18120);
  not g45173 (n_18352, n26916);
  not g45174 (n_18353, n26917);
  and g45175 (n26918, n_18352, n_18353);
  and g45176 (n26919, n26915, n26918);
  not g45177 (n_18354, n26915);
  not g45178 (n_18355, n26918);
  and g45179 (n26920, n_18354, n_18355);
  or g45180 (\result[0] , n26919, n26920);
  and g45181 (n26922, n26915, n_18355);
  and g45182 (n26923, n_18346, n_18350);
  and g45183 (n26924, n71, n26066);
  and g45184 (n26925, n9867, n22309);
  and g45185 (n26926, n10434, n26063);
  not g45191 (n_18359, n26624);
  and g45192 (n26929, n9870, n_18359);
  not g45195 (n_18361, n26930);
  and g45196 (n26931, \a[5] , n_18361);
  not g45197 (n_18362, n26931);
  and g45198 (n26932, n_18361, n_18362);
  and g45199 (n26933, \a[5] , n_18362);
  not g45200 (n_18363, n26932);
  not g45201 (n_18364, n26933);
  and g45202 (n26934, n_18363, n_18364);
  and g45203 (n26935, n_18276, n_18281);
  and g45204 (n26936, n7983, n22323);
  and g45205 (n26937, n7291, n22329);
  and g45206 (n26938, n7632, n22326);
  and g45212 (n26941, n7294, n24599);
  not g45215 (n_18369, n26942);
  and g45216 (n26943, \a[11] , n_18369);
  not g45217 (n_18370, n26943);
  and g45218 (n26944, n_18369, n_18370);
  and g45219 (n26945, \a[11] , n_18370);
  not g45220 (n_18371, n26944);
  not g45221 (n_18372, n26945);
  and g45222 (n26946, n_18371, n_18372);
  and g45223 (n26947, n_18250, n_18255);
  and g45224 (n26948, n6233, n22341);
  and g45225 (n26949, n5663, n22347);
  and g45226 (n26950, n5939, n22344);
  and g45232 (n26953, n5666, n24142);
  not g45235 (n_18377, n26954);
  and g45236 (n26955, \a[17] , n_18377);
  not g45237 (n_18378, n26955);
  and g45238 (n26956, n_18377, n_18378);
  and g45239 (n26957, \a[17] , n_18378);
  not g45240 (n_18379, n26956);
  not g45241 (n_18380, n26957);
  and g45242 (n26958, n_18379, n_18380);
  and g45243 (n26959, n_18224, n_18229);
  and g45244 (n26960, n4694, n22359);
  and g45245 (n26961, n4533, n22365);
  and g45246 (n26962, n4604, n22362);
  and g45252 (n26965, n4536, n23368);
  not g45255 (n_18385, n26966);
  and g45256 (n26967, \a[23] , n_18385);
  not g45257 (n_18386, n26967);
  and g45258 (n26968, n_18385, n_18386);
  and g45259 (n26969, \a[23] , n_18386);
  not g45260 (n_18387, n26968);
  not g45261 (n_18388, n26969);
  and g45262 (n26970, n_18387, n_18388);
  and g45263 (n26971, n_18198, n_18203);
  and g45264 (n26972, n_18181, n_18187);
  and g45265 (n26973, n_18171, n_18176);
  and g45284 (n26992, n3020, n22387);
  and g45285 (n26993, n3028, n22390);
  and g45286 (n26994, n3023, n22393);
  and g45287 (n26995, n75, n22582);
  not g45295 (n_18393, n26991);
  not g45296 (n_18394, n26998);
  and g45297 (n26999, n_18393, n_18394);
  not g45298 (n_18395, n26999);
  and g45299 (n27000, n_18393, n_18395);
  and g45300 (n27001, n_18394, n_18395);
  not g45301 (n_18396, n27000);
  not g45302 (n_18397, n27001);
  and g45303 (n27002, n_18396, n_18397);
  not g45304 (n_18398, n26973);
  not g45305 (n_18399, n27002);
  and g45306 (n27003, n_18398, n_18399);
  not g45307 (n_18400, n27003);
  and g45308 (n27004, n_18398, n_18400);
  and g45309 (n27005, n_18399, n_18400);
  not g45310 (n_18401, n27004);
  not g45311 (n_18402, n27005);
  and g45312 (n27006, n_18401, n_18402);
  and g45313 (n27007, n3457, n22377);
  and g45314 (n27008, n3542, n22384);
  and g45315 (n27009, n3606, n22380);
  not g45316 (n_18403, n27008);
  not g45317 (n_18404, n27009);
  and g45318 (n27010, n_18403, n_18404);
  not g45319 (n_18405, n27007);
  and g45320 (n27011, n_18405, n27010);
  and g45321 (n27012, n_489, n27011);
  and g45322 (n27013, n22834, n27011);
  not g45323 (n_18406, n27012);
  not g45324 (n_18407, n27013);
  and g45325 (n27014, n_18406, n_18407);
  not g45326 (n_18408, n27014);
  and g45327 (n27015, \a[29] , n_18408);
  and g45328 (n27016, n_15, n27014);
  not g45329 (n_18409, n27015);
  not g45330 (n_18410, n27016);
  and g45331 (n27017, n_18409, n_18410);
  not g45332 (n_18411, n27006);
  not g45333 (n_18412, n27017);
  and g45334 (n27018, n_18411, n_18412);
  and g45335 (n27019, n27006, n27017);
  not g45336 (n_18413, n27018);
  not g45337 (n_18414, n27019);
  and g45338 (n27020, n_18413, n_18414);
  not g45339 (n_18415, n26972);
  and g45340 (n27021, n_18415, n27020);
  not g45341 (n_18416, n27020);
  and g45342 (n27022, n26972, n_18416);
  not g45343 (n_18417, n27021);
  not g45344 (n_18418, n27022);
  and g45345 (n27023, n_18417, n_18418);
  and g45346 (n27024, n3884, n22368);
  and g45347 (n27025, n3967, n22374);
  and g45348 (n27026, n4046, n22371);
  not g45349 (n_18419, n27025);
  not g45350 (n_18420, n27026);
  and g45351 (n27027, n_18419, n_18420);
  not g45352 (n_18421, n27024);
  and g45353 (n27028, n_18421, n27027);
  and g45354 (n27029, n_750, n27028);
  not g45355 (n_18422, n23006);
  and g45356 (n27030, n_18422, n27028);
  not g45357 (n_18423, n27029);
  not g45358 (n_18424, n27030);
  and g45359 (n27031, n_18423, n_18424);
  not g45360 (n_18425, n27031);
  and g45361 (n27032, \a[26] , n_18425);
  and g45362 (n27033, n_33, n27031);
  not g45363 (n_18426, n27032);
  not g45364 (n_18427, n27033);
  and g45365 (n27034, n_18426, n_18427);
  not g45366 (n_18428, n27034);
  and g45367 (n27035, n27023, n_18428);
  not g45368 (n_18429, n27035);
  and g45369 (n27036, n27023, n_18429);
  and g45370 (n27037, n_18428, n_18429);
  not g45371 (n_18430, n27036);
  not g45372 (n_18431, n27037);
  and g45373 (n27038, n_18430, n_18431);
  not g45374 (n_18432, n26971);
  not g45375 (n_18433, n27038);
  and g45376 (n27039, n_18432, n_18433);
  not g45377 (n_18434, n27039);
  and g45378 (n27040, n_18432, n_18434);
  and g45379 (n27041, n_18433, n_18434);
  not g45380 (n_18435, n27040);
  not g45381 (n_18436, n27041);
  and g45382 (n27042, n_18435, n_18436);
  not g45383 (n_18437, n26970);
  not g45384 (n_18438, n27042);
  and g45385 (n27043, n_18437, n_18438);
  not g45386 (n_18439, n27043);
  and g45387 (n27044, n_18437, n_18439);
  and g45388 (n27045, n_18438, n_18439);
  not g45389 (n_18440, n27044);
  not g45390 (n_18441, n27045);
  and g45391 (n27046, n_18440, n_18441);
  and g45392 (n27047, n_18208, n_18214);
  and g45393 (n27048, n27046, n27047);
  not g45394 (n_18442, n27046);
  not g45395 (n_18443, n27047);
  and g45396 (n27049, n_18442, n_18443);
  not g45397 (n_18444, n27048);
  not g45398 (n_18445, n27049);
  and g45399 (n27050, n_18444, n_18445);
  and g45400 (n27051, n5496, n22350);
  and g45401 (n27052, n4935, n22356);
  and g45402 (n27053, n5407, n22353);
  not g45403 (n_18446, n27052);
  not g45404 (n_18447, n27053);
  and g45405 (n27054, n_18446, n_18447);
  not g45406 (n_18448, n27051);
  and g45407 (n27055, n_18448, n27054);
  and g45408 (n27056, n_1011, n27055);
  not g45409 (n_18449, n23672);
  and g45410 (n27057, n_18449, n27055);
  not g45411 (n_18450, n27056);
  not g45412 (n_18451, n27057);
  and g45413 (n27058, n_18450, n_18451);
  not g45414 (n_18452, n27058);
  and g45415 (n27059, \a[20] , n_18452);
  and g45416 (n27060, n_435, n27058);
  not g45417 (n_18453, n27059);
  not g45418 (n_18454, n27060);
  and g45419 (n27061, n_18453, n_18454);
  not g45420 (n_18455, n27061);
  and g45421 (n27062, n27050, n_18455);
  not g45422 (n_18456, n27062);
  and g45423 (n27063, n27050, n_18456);
  and g45424 (n27064, n_18455, n_18456);
  not g45425 (n_18457, n27063);
  not g45426 (n_18458, n27064);
  and g45427 (n27065, n_18457, n_18458);
  not g45428 (n_18459, n26959);
  not g45429 (n_18460, n27065);
  and g45430 (n27066, n_18459, n_18460);
  not g45431 (n_18461, n27066);
  and g45432 (n27067, n_18459, n_18461);
  and g45433 (n27068, n_18460, n_18461);
  not g45434 (n_18462, n27067);
  not g45435 (n_18463, n27068);
  and g45436 (n27069, n_18462, n_18463);
  not g45437 (n_18464, n26958);
  not g45438 (n_18465, n27069);
  and g45439 (n27070, n_18464, n_18465);
  not g45440 (n_18466, n27070);
  and g45441 (n27071, n_18464, n_18466);
  and g45442 (n27072, n_18465, n_18466);
  not g45443 (n_18467, n27071);
  not g45444 (n_18468, n27072);
  and g45445 (n27073, n_18467, n_18468);
  and g45446 (n27074, n_18234, n_18240);
  and g45447 (n27075, n27073, n27074);
  not g45448 (n_18469, n27073);
  not g45449 (n_18470, n27074);
  and g45450 (n27076, n_18469, n_18470);
  not g45451 (n_18471, n27075);
  not g45452 (n_18472, n27076);
  and g45453 (n27077, n_18471, n_18472);
  and g45454 (n27078, n7101, n22332);
  and g45455 (n27079, n6402, n22338);
  and g45456 (n27080, n6951, n22335);
  not g45457 (n_18473, n27079);
  not g45458 (n_18474, n27080);
  and g45459 (n27081, n_18473, n_18474);
  not g45460 (n_18475, n27078);
  and g45461 (n27082, n_18475, n27081);
  and g45462 (n27083, n_1885, n27082);
  not g45463 (n_18476, n22542);
  and g45464 (n27084, n_18476, n27082);
  not g45465 (n_18477, n27083);
  not g45466 (n_18478, n27084);
  and g45467 (n27085, n_18477, n_18478);
  not g45468 (n_18479, n27085);
  and g45469 (n27086, \a[14] , n_18479);
  and g45470 (n27087, n_652, n27085);
  not g45471 (n_18480, n27086);
  not g45472 (n_18481, n27087);
  and g45473 (n27088, n_18480, n_18481);
  not g45474 (n_18482, n27088);
  and g45475 (n27089, n27077, n_18482);
  not g45476 (n_18483, n27089);
  and g45477 (n27090, n27077, n_18483);
  and g45478 (n27091, n_18482, n_18483);
  not g45479 (n_18484, n27090);
  not g45480 (n_18485, n27091);
  and g45481 (n27092, n_18484, n_18485);
  not g45482 (n_18486, n26947);
  not g45483 (n_18487, n27092);
  and g45484 (n27093, n_18486, n_18487);
  not g45485 (n_18488, n27093);
  and g45486 (n27094, n_18486, n_18488);
  and g45487 (n27095, n_18487, n_18488);
  not g45488 (n_18489, n27094);
  not g45489 (n_18490, n27095);
  and g45490 (n27096, n_18489, n_18490);
  not g45491 (n_18491, n26946);
  not g45492 (n_18492, n27096);
  and g45493 (n27097, n_18491, n_18492);
  not g45494 (n_18493, n27097);
  and g45495 (n27098, n_18491, n_18493);
  and g45496 (n27099, n_18492, n_18493);
  not g45497 (n_18494, n27098);
  not g45498 (n_18495, n27099);
  and g45499 (n27100, n_18494, n_18495);
  and g45500 (n27101, n_18260, n_18266);
  and g45501 (n27102, n27100, n27101);
  not g45502 (n_18496, n27100);
  not g45503 (n_18497, n27101);
  and g45504 (n27103, n_18496, n_18497);
  not g45505 (n_18498, n27102);
  not g45506 (n_18499, n27103);
  and g45507 (n27104, n_18498, n_18499);
  and g45508 (n27105, n9331, n22315);
  and g45509 (n27106, n8418, n22320);
  and g45510 (n27107, n8860, n22312);
  not g45511 (n_18500, n27106);
  not g45512 (n_18501, n27107);
  and g45513 (n27108, n_18500, n_18501);
  not g45514 (n_18502, n27105);
  and g45515 (n27109, n_18502, n27108);
  and g45516 (n27110, n_3428, n27109);
  not g45517 (n_18503, n25294);
  and g45518 (n27111, n_18503, n27109);
  not g45519 (n_18504, n27110);
  not g45520 (n_18505, n27111);
  and g45521 (n27112, n_18504, n_18505);
  not g45522 (n_18506, n27112);
  and g45523 (n27113, \a[8] , n_18506);
  and g45524 (n27114, n_1106, n27112);
  not g45525 (n_18507, n27113);
  not g45526 (n_18508, n27114);
  and g45527 (n27115, n_18507, n_18508);
  not g45528 (n_18509, n27115);
  and g45529 (n27116, n27104, n_18509);
  not g45530 (n_18510, n27116);
  and g45531 (n27117, n27104, n_18510);
  and g45532 (n27118, n_18509, n_18510);
  not g45533 (n_18511, n27117);
  not g45534 (n_18512, n27118);
  and g45535 (n27119, n_18511, n_18512);
  not g45536 (n_18513, n26935);
  not g45537 (n_18514, n27119);
  and g45538 (n27120, n_18513, n_18514);
  not g45539 (n_18515, n27120);
  and g45540 (n27121, n_18513, n_18515);
  and g45541 (n27122, n_18514, n_18515);
  not g45542 (n_18516, n27121);
  not g45543 (n_18517, n27122);
  and g45544 (n27123, n_18516, n_18517);
  not g45545 (n_18518, n26934);
  not g45546 (n_18519, n27123);
  and g45547 (n27124, n_18518, n_18519);
  not g45548 (n_18520, n27124);
  and g45549 (n27125, n_18518, n_18520);
  and g45550 (n27126, n_18519, n_18520);
  not g45551 (n_18521, n27125);
  not g45552 (n_18522, n27126);
  and g45553 (n27127, n_18521, n_18522);
  and g45554 (n27128, n_18286, n_18292);
  and g45555 (n27129, n27127, n27128);
  not g45556 (n_18523, n27127);
  not g45557 (n_18524, n27128);
  and g45558 (n27130, n_18523, n_18524);
  not g45559 (n_18525, n27129);
  not g45560 (n_18526, n27130);
  and g45561 (n27131, n_18525, n_18526);
  and g45562 (n27132, n_18323, n_18327);
  and g45563 (n27133, n_18308, n_18319);
  and g45564 (n27134, n_18299, n_18302);
  and g45565 (n27135, n3856, n4514);
  not g45566 (n_18527, n27135);
  and g45567 (n27136, n26859, n_18527);
  and g45568 (n27137, n_18298, n27135);
  not g45569 (n_18528, n27134);
  not g45570 (n_18529, n27137);
  and g45571 (n27138, n_18528, n_18529);
  not g45572 (n_18530, n27136);
  and g45573 (n27139, n_18530, n27138);
  not g45574 (n_18531, n27139);
  and g45575 (n27140, n_18528, n_18531);
  and g45576 (n27141, n_18529, n_18531);
  and g45577 (n27142, n_18530, n27141);
  not g45578 (n_18532, n27140);
  not g45579 (n_18533, n27142);
  and g45580 (n27143, n_18532, n_18533);
  not g45581 (n_18534, n3457);
  not g45582 (n_18535, n3606);
  and g45583 (n27144, n_18534, n_18535);
  not g45584 (n_18536, n27144);
  and g45585 (n27145, n_7417, n_18536);
  and g45586 (n27146, n3542, n13941);
  not g45587 (n_18537, n27145);
  not g45588 (n_18538, n27146);
  and g45589 (n27147, n_18537, n_18538);
  and g45590 (n27148, n3368, n_13153);
  not g45591 (n_18539, n27148);
  and g45592 (n27149, n27147, n_18539);
  not g45593 (n_18540, n27149);
  and g45594 (n27150, \a[29] , n_18540);
  not g45595 (n_18541, n27150);
  and g45596 (n27151, n_18540, n_18541);
  and g45597 (n27152, \a[29] , n_18541);
  not g45598 (n_18542, n27151);
  not g45599 (n_18543, n27152);
  and g45600 (n27153, n_18542, n_18543);
  and g45601 (n27154, n75, n_7563);
  and g45602 (n27155, n3020, n_7540);
  and g45603 (n27156, n3023, n13630);
  and g45604 (n27157, n3028, n13633);
  not g45612 (n_18548, n27153);
  not g45613 (n_18549, n27160);
  and g45614 (n27161, n_18548, n_18549);
  not g45615 (n_18550, n27161);
  and g45616 (n27162, n_18548, n_18550);
  and g45617 (n27163, n_18549, n_18550);
  not g45618 (n_18551, n27162);
  not g45619 (n_18552, n27163);
  and g45620 (n27164, n_18551, n_18552);
  not g45621 (n_18553, n27143);
  and g45622 (n27165, n_18553, n27164);
  not g45623 (n_18554, n27164);
  and g45624 (n27166, n27143, n_18554);
  not g45625 (n_18555, n27165);
  not g45626 (n_18556, n27166);
  and g45627 (n27167, n_18555, n_18556);
  not g45628 (n_18557, n27133);
  not g45629 (n_18558, n27167);
  and g45630 (n27168, n_18557, n_18558);
  and g45631 (n27169, n27133, n27167);
  not g45632 (n_18559, n27168);
  not g45633 (n_18560, n27169);
  and g45634 (n27170, n_18559, n_18560);
  not g45635 (n_18561, n27132);
  and g45636 (n27171, n_18561, n27170);
  not g45637 (n_18562, n27170);
  and g45638 (n27172, n27132, n_18562);
  not g45639 (n_18563, n27171);
  not g45640 (n_18564, n27172);
  and g45641 (n27173, n_18563, n_18564);
  and g45642 (n27174, n11727, n27173);
  and g45643 (n27175, n11055, n26060);
  and g45644 (n27176, n11715, n26890);
  not g45645 (n_18565, n27175);
  not g45646 (n_18566, n27176);
  and g45647 (n27177, n_18565, n_18566);
  not g45648 (n_18567, n27174);
  and g45649 (n27178, n_18567, n27177);
  and g45650 (n27179, n_6291, n27178);
  not g45651 (n_18568, n27173);
  and g45652 (n27180, n_18332, n_18568);
  and g45653 (n27181, n26890, n27173);
  not g45654 (n_18569, n27180);
  not g45655 (n_18570, n27181);
  and g45656 (n27182, n_18569, n_18570);
  not g45657 (n_18571, n26902);
  and g45658 (n27183, n_18571, n27182);
  not g45659 (n_18572, n27182);
  and g45660 (n27184, n26902, n_18572);
  not g45661 (n_18573, n27183);
  not g45662 (n_18574, n27184);
  and g45663 (n27185, n_18573, n_18574);
  not g45664 (n_18575, n27185);
  and g45665 (n27186, n27178, n_18575);
  not g45666 (n_18576, n27179);
  not g45667 (n_18577, n27186);
  and g45668 (n27187, n_18576, n_18577);
  not g45669 (n_18578, n27187);
  and g45670 (n27188, \a[2] , n_18578);
  and g45671 (n27189, n_10, n27187);
  not g45672 (n_18579, n27188);
  not g45673 (n_18580, n27189);
  and g45674 (n27190, n_18579, n_18580);
  not g45675 (n_18581, n27190);
  and g45676 (n27191, n27131, n_18581);
  not g45677 (n_18582, n27131);
  and g45678 (n27192, n_18582, n27190);
  not g45679 (n_18583, n27191);
  not g45680 (n_18584, n27192);
  and g45681 (n27193, n_18583, n_18584);
  not g45682 (n_18585, n26923);
  and g45683 (n27194, n_18585, n27193);
  not g45684 (n_18586, n27193);
  and g45685 (n27195, n26923, n_18586);
  not g45686 (n_18587, n27194);
  not g45687 (n_18588, n27195);
  and g45688 (n27196, n_18587, n_18588);
  and g45689 (n27197, n26922, n27196);
  not g45690 (n_18589, n26922);
  not g45691 (n_18590, n27196);
  and g45692 (n27198, n_18589, n_18590);
  not g45693 (n_18591, n27197);
  not g45694 (n_18592, n27198);
  and g45695 (\result[1] , n_18591, n_18592);
  and g45696 (n27200, n_18583, n_18587);
  and g45697 (n27201, n71, n26060);
  and g45698 (n27202, n9867, n26063);
  and g45699 (n27203, n10434, n26066);
  not g45705 (n_18596, n26088);
  and g45706 (n27206, n9870, n_18596);
  not g45709 (n_18598, n27207);
  and g45710 (n27208, \a[5] , n_18598);
  not g45711 (n_18599, n27208);
  and g45712 (n27209, n_18598, n_18599);
  and g45713 (n27210, \a[5] , n_18599);
  not g45714 (n_18600, n27209);
  not g45715 (n_18601, n27210);
  and g45716 (n27211, n_18600, n_18601);
  and g45717 (n27212, n_18510, n_18515);
  and g45718 (n27213, n7983, n22320);
  and g45719 (n27214, n7291, n22326);
  and g45720 (n27215, n7632, n22323);
  and g45726 (n27218, n7294, n_17020);
  not g45729 (n_18606, n27219);
  and g45730 (n27220, \a[11] , n_18606);
  not g45731 (n_18607, n27220);
  and g45732 (n27221, n_18606, n_18607);
  and g45733 (n27222, \a[11] , n_18607);
  not g45734 (n_18608, n27221);
  not g45735 (n_18609, n27222);
  and g45736 (n27223, n_18608, n_18609);
  and g45737 (n27224, n_18483, n_18488);
  and g45738 (n27225, n6233, n22338);
  and g45739 (n27226, n5663, n22344);
  and g45740 (n27227, n5939, n22341);
  and g45746 (n27230, n5666, n_16033);
  not g45749 (n_18614, n27231);
  and g45750 (n27232, \a[17] , n_18614);
  not g45751 (n_18615, n27232);
  and g45752 (n27233, n_18614, n_18615);
  and g45753 (n27234, \a[17] , n_18615);
  not g45754 (n_18616, n27233);
  not g45755 (n_18617, n27234);
  and g45756 (n27235, n_18616, n_18617);
  and g45757 (n27236, n_18456, n_18461);
  and g45758 (n27237, n4694, n22356);
  and g45759 (n27238, n4533, n22362);
  and g45760 (n27239, n4604, n22359);
  and g45766 (n27242, n4536, n_15312);
  not g45769 (n_18622, n27243);
  and g45770 (n27244, \a[23] , n_18622);
  not g45771 (n_18623, n27244);
  and g45772 (n27245, n_18622, n_18623);
  and g45773 (n27246, \a[23] , n_18623);
  not g45774 (n_18624, n27245);
  not g45775 (n_18625, n27246);
  and g45776 (n27247, n_18624, n_18625);
  and g45777 (n27248, n_18429, n_18434);
  and g45778 (n27249, n_18413, n_18417);
  and g45779 (n27250, n_18395, n_18400);
  and g45797 (n27268, n3020, n22384);
  and g45798 (n27269, n3028, n22387);
  and g45799 (n27270, n3023, n22390);
  and g45800 (n27271, n75, n22806);
  not g45808 (n_18630, n27267);
  not g45809 (n_18631, n27274);
  and g45810 (n27275, n_18630, n_18631);
  not g45811 (n_18632, n27275);
  and g45812 (n27276, n_18630, n_18632);
  and g45813 (n27277, n_18631, n_18632);
  not g45814 (n_18633, n27276);
  not g45815 (n_18634, n27277);
  and g45816 (n27278, n_18633, n_18634);
  not g45817 (n_18635, n27250);
  not g45818 (n_18636, n27278);
  and g45819 (n27279, n_18635, n_18636);
  not g45820 (n_18637, n27279);
  and g45821 (n27280, n_18635, n_18637);
  and g45822 (n27281, n_18636, n_18637);
  not g45823 (n_18638, n27280);
  not g45824 (n_18639, n27281);
  and g45825 (n27282, n_18638, n_18639);
  and g45826 (n27283, n3457, n22374);
  and g45827 (n27284, n3542, n22380);
  and g45828 (n27285, n3606, n22377);
  not g45829 (n_18640, n27284);
  not g45830 (n_18641, n27285);
  and g45831 (n27286, n_18640, n_18641);
  not g45832 (n_18642, n27283);
  and g45833 (n27287, n_18642, n27286);
  and g45834 (n27288, n_489, n27287);
  and g45835 (n27289, n_15064, n27287);
  not g45836 (n_18643, n27288);
  not g45837 (n_18644, n27289);
  and g45838 (n27290, n_18643, n_18644);
  not g45839 (n_18645, n27290);
  and g45840 (n27291, \a[29] , n_18645);
  and g45841 (n27292, n_15, n27290);
  not g45842 (n_18646, n27291);
  not g45843 (n_18647, n27292);
  and g45844 (n27293, n_18646, n_18647);
  not g45845 (n_18648, n27282);
  not g45846 (n_18649, n27293);
  and g45847 (n27294, n_18648, n_18649);
  and g45848 (n27295, n27282, n27293);
  not g45849 (n_18650, n27294);
  not g45850 (n_18651, n27295);
  and g45851 (n27296, n_18650, n_18651);
  not g45852 (n_18652, n27249);
  and g45853 (n27297, n_18652, n27296);
  not g45854 (n_18653, n27296);
  and g45855 (n27298, n27249, n_18653);
  not g45856 (n_18654, n27297);
  not g45857 (n_18655, n27298);
  and g45858 (n27299, n_18654, n_18655);
  and g45859 (n27300, n3884, n22365);
  and g45860 (n27301, n3967, n22371);
  and g45861 (n27302, n4046, n22368);
  not g45862 (n_18656, n27301);
  not g45863 (n_18657, n27302);
  and g45864 (n27303, n_18656, n_18657);
  not g45865 (n_18658, n27300);
  and g45866 (n27304, n_18658, n27303);
  and g45867 (n27305, n_750, n27304);
  and g45868 (n27306, n22993, n27304);
  not g45869 (n_18659, n27305);
  not g45870 (n_18660, n27306);
  and g45871 (n27307, n_18659, n_18660);
  not g45872 (n_18661, n27307);
  and g45873 (n27308, \a[26] , n_18661);
  and g45874 (n27309, n_33, n27307);
  not g45875 (n_18662, n27308);
  not g45876 (n_18663, n27309);
  and g45877 (n27310, n_18662, n_18663);
  not g45878 (n_18664, n27310);
  and g45879 (n27311, n27299, n_18664);
  not g45880 (n_18665, n27311);
  and g45881 (n27312, n27299, n_18665);
  and g45882 (n27313, n_18664, n_18665);
  not g45883 (n_18666, n27312);
  not g45884 (n_18667, n27313);
  and g45885 (n27314, n_18666, n_18667);
  not g45886 (n_18668, n27248);
  not g45887 (n_18669, n27314);
  and g45888 (n27315, n_18668, n_18669);
  not g45889 (n_18670, n27315);
  and g45890 (n27316, n_18668, n_18670);
  and g45891 (n27317, n_18669, n_18670);
  not g45892 (n_18671, n27316);
  not g45893 (n_18672, n27317);
  and g45894 (n27318, n_18671, n_18672);
  not g45895 (n_18673, n27247);
  not g45896 (n_18674, n27318);
  and g45897 (n27319, n_18673, n_18674);
  not g45898 (n_18675, n27319);
  and g45899 (n27320, n_18673, n_18675);
  and g45900 (n27321, n_18674, n_18675);
  not g45901 (n_18676, n27320);
  not g45902 (n_18677, n27321);
  and g45903 (n27322, n_18676, n_18677);
  and g45904 (n27323, n_18439, n_18445);
  and g45905 (n27324, n27322, n27323);
  not g45906 (n_18678, n27322);
  not g45907 (n_18679, n27323);
  and g45908 (n27325, n_18678, n_18679);
  not g45909 (n_18680, n27324);
  not g45910 (n_18681, n27325);
  and g45911 (n27326, n_18680, n_18681);
  and g45912 (n27327, n5496, n22347);
  and g45913 (n27328, n4935, n22353);
  and g45914 (n27329, n5407, n22350);
  not g45915 (n_18682, n27328);
  not g45916 (n_18683, n27329);
  and g45917 (n27330, n_18682, n_18683);
  not g45918 (n_18684, n27327);
  and g45919 (n27331, n_18684, n27330);
  and g45920 (n27332, n_1011, n27331);
  and g45921 (n27333, n23659, n27331);
  not g45922 (n_18685, n27332);
  not g45923 (n_18686, n27333);
  and g45924 (n27334, n_18685, n_18686);
  not g45925 (n_18687, n27334);
  and g45926 (n27335, \a[20] , n_18687);
  and g45927 (n27336, n_435, n27334);
  not g45928 (n_18688, n27335);
  not g45929 (n_18689, n27336);
  and g45930 (n27337, n_18688, n_18689);
  not g45931 (n_18690, n27337);
  and g45932 (n27338, n27326, n_18690);
  not g45933 (n_18691, n27338);
  and g45934 (n27339, n27326, n_18691);
  and g45935 (n27340, n_18690, n_18691);
  not g45936 (n_18692, n27339);
  not g45937 (n_18693, n27340);
  and g45938 (n27341, n_18692, n_18693);
  not g45939 (n_18694, n27236);
  not g45940 (n_18695, n27341);
  and g45941 (n27342, n_18694, n_18695);
  not g45942 (n_18696, n27342);
  and g45943 (n27343, n_18694, n_18696);
  and g45944 (n27344, n_18695, n_18696);
  not g45945 (n_18697, n27343);
  not g45946 (n_18698, n27344);
  and g45947 (n27345, n_18697, n_18698);
  not g45948 (n_18699, n27235);
  not g45949 (n_18700, n27345);
  and g45950 (n27346, n_18699, n_18700);
  not g45951 (n_18701, n27346);
  and g45952 (n27347, n_18699, n_18701);
  and g45953 (n27348, n_18700, n_18701);
  not g45954 (n_18702, n27347);
  not g45955 (n_18703, n27348);
  and g45956 (n27349, n_18702, n_18703);
  and g45957 (n27350, n_18466, n_18472);
  and g45958 (n27351, n27349, n27350);
  not g45959 (n_18704, n27349);
  not g45960 (n_18705, n27350);
  and g45961 (n27352, n_18704, n_18705);
  not g45962 (n_18706, n27351);
  not g45963 (n_18707, n27352);
  and g45964 (n27353, n_18706, n_18707);
  and g45965 (n27354, n7101, n22329);
  and g45966 (n27355, n6402, n22335);
  and g45967 (n27356, n6951, n22332);
  not g45968 (n_18708, n27355);
  not g45969 (n_18709, n27356);
  and g45970 (n27357, n_18708, n_18709);
  not g45971 (n_18710, n27354);
  and g45972 (n27358, n_18710, n27357);
  and g45973 (n27359, n_1885, n27358);
  and g45974 (n27360, n24633, n27358);
  not g45975 (n_18711, n27359);
  not g45976 (n_18712, n27360);
  and g45977 (n27361, n_18711, n_18712);
  not g45978 (n_18713, n27361);
  and g45979 (n27362, \a[14] , n_18713);
  and g45980 (n27363, n_652, n27361);
  not g45981 (n_18714, n27362);
  not g45982 (n_18715, n27363);
  and g45983 (n27364, n_18714, n_18715);
  not g45984 (n_18716, n27364);
  and g45985 (n27365, n27353, n_18716);
  not g45986 (n_18717, n27365);
  and g45987 (n27366, n27353, n_18717);
  and g45988 (n27367, n_18716, n_18717);
  not g45989 (n_18718, n27366);
  not g45990 (n_18719, n27367);
  and g45991 (n27368, n_18718, n_18719);
  not g45992 (n_18720, n27224);
  not g45993 (n_18721, n27368);
  and g45994 (n27369, n_18720, n_18721);
  not g45995 (n_18722, n27369);
  and g45996 (n27370, n_18720, n_18722);
  and g45997 (n27371, n_18721, n_18722);
  not g45998 (n_18723, n27370);
  not g45999 (n_18724, n27371);
  and g46000 (n27372, n_18723, n_18724);
  not g46001 (n_18725, n27223);
  not g46002 (n_18726, n27372);
  and g46003 (n27373, n_18725, n_18726);
  not g46004 (n_18727, n27373);
  and g46005 (n27374, n_18725, n_18727);
  and g46006 (n27375, n_18726, n_18727);
  not g46007 (n_18728, n27374);
  not g46008 (n_18729, n27375);
  and g46009 (n27376, n_18728, n_18729);
  and g46010 (n27377, n_18493, n_18499);
  and g46011 (n27378, n27376, n27377);
  not g46012 (n_18730, n27376);
  not g46013 (n_18731, n27377);
  and g46014 (n27379, n_18730, n_18731);
  not g46015 (n_18732, n27378);
  not g46016 (n_18733, n27379);
  and g46017 (n27380, n_18732, n_18733);
  and g46018 (n27381, n9331, n22309);
  and g46019 (n27382, n8418, n22312);
  and g46020 (n27383, n8860, n22315);
  not g46021 (n_18734, n27382);
  not g46022 (n_18735, n27383);
  and g46023 (n27384, n_18734, n_18735);
  not g46024 (n_18736, n27381);
  and g46025 (n27385, n_18736, n27384);
  and g46026 (n27386, n_3428, n27385);
  and g46027 (n27387, n22529, n27385);
  not g46028 (n_18737, n27386);
  not g46029 (n_18738, n27387);
  and g46030 (n27388, n_18737, n_18738);
  not g46031 (n_18739, n27388);
  and g46032 (n27389, \a[8] , n_18739);
  and g46033 (n27390, n_1106, n27388);
  not g46034 (n_18740, n27389);
  not g46035 (n_18741, n27390);
  and g46036 (n27391, n_18740, n_18741);
  not g46037 (n_18742, n27391);
  and g46038 (n27392, n27380, n_18742);
  not g46039 (n_18743, n27392);
  and g46040 (n27393, n27380, n_18743);
  and g46041 (n27394, n_18742, n_18743);
  not g46042 (n_18744, n27393);
  not g46043 (n_18745, n27394);
  and g46044 (n27395, n_18744, n_18745);
  not g46045 (n_18746, n27212);
  not g46046 (n_18747, n27395);
  and g46047 (n27396, n_18746, n_18747);
  not g46048 (n_18748, n27396);
  and g46049 (n27397, n_18746, n_18748);
  and g46050 (n27398, n_18747, n_18748);
  not g46051 (n_18749, n27397);
  not g46052 (n_18750, n27398);
  and g46053 (n27399, n_18749, n_18750);
  not g46054 (n_18751, n27211);
  not g46055 (n_18752, n27399);
  and g46056 (n27400, n_18751, n_18752);
  not g46057 (n_18753, n27400);
  and g46058 (n27401, n_18751, n_18753);
  and g46059 (n27402, n_18752, n_18753);
  not g46060 (n_18754, n27401);
  not g46061 (n_18755, n27402);
  and g46062 (n27403, n_18754, n_18755);
  and g46063 (n27404, n_18520, n_18526);
  and g46064 (n27405, n27403, n27404);
  not g46065 (n_18756, n27403);
  not g46066 (n_18757, n27404);
  and g46067 (n27406, n_18756, n_18757);
  not g46068 (n_18758, n27405);
  not g46069 (n_18759, n27406);
  and g46070 (n27407, n_18758, n_18759);
  and g46071 (n27408, n_18559, n_18563);
  and g46072 (n27409, n_18553, n_18554);
  not g46073 (n_18760, n27409);
  and g46074 (n27410, n_18550, n_18760);
  and g46075 (n27411, n75, n14136);
  and g46076 (n27412, n3020, n13941);
  and g46077 (n27413, n3023, n13633);
  and g46078 (n27414, n3028, n_7540);
  not g46086 (n_18765, n3542);
  and g46087 (n27418, n_18765, n_18535);
  and g46088 (n27419, n3367, n27418);
  not g46089 (n_18766, n27419);
  and g46090 (n27420, n_7417, n_18766);
  not g46091 (n_18767, n27420);
  and g46092 (n27421, \a[29] , n_18767);
  and g46093 (n27422, n_15, n27420);
  not g46094 (n_18768, n27421);
  not g46095 (n_18769, n27422);
  and g46096 (n27423, n_18768, n_18769);
  and g46097 (n27424, n13056, n27135);
  not g46098 (n_18770, n13056);
  and g46099 (n27425, n_18770, n_18527);
  not g46100 (n_18771, n27424);
  not g46101 (n_18772, n27425);
  and g46102 (n27426, n_18771, n_18772);
  and g46103 (n27427, n27423, n27426);
  not g46104 (n_18773, n27423);
  not g46105 (n_18774, n27426);
  and g46106 (n27428, n_18773, n_18774);
  not g46107 (n_18775, n27427);
  not g46108 (n_18776, n27428);
  and g46109 (n27429, n_18775, n_18776);
  not g46110 (n_18777, n27417);
  and g46111 (n27430, n_18777, n27429);
  not g46112 (n_18778, n27430);
  and g46113 (n27431, n27429, n_18778);
  and g46114 (n27432, n_18777, n_18778);
  not g46115 (n_18779, n27431);
  not g46116 (n_18780, n27432);
  and g46117 (n27433, n_18779, n_18780);
  not g46118 (n_18781, n27141);
  not g46119 (n_18782, n27433);
  and g46120 (n27434, n_18781, n_18782);
  and g46121 (n27435, n27141, n27433);
  not g46122 (n_18783, n27434);
  not g46123 (n_18784, n27435);
  and g46124 (n27436, n_18783, n_18784);
  not g46125 (n_18785, n27410);
  and g46126 (n27437, n_18785, n27436);
  not g46127 (n_18786, n27436);
  and g46128 (n27438, n27410, n_18786);
  not g46129 (n_18787, n27437);
  not g46130 (n_18788, n27438);
  and g46131 (n27439, n_18787, n_18788);
  not g46132 (n_18789, n27408);
  and g46133 (n27440, n_18789, n27439);
  not g46134 (n_18790, n27439);
  and g46135 (n27441, n27408, n_18790);
  not g46136 (n_18791, n27440);
  not g46137 (n_18792, n27441);
  and g46138 (n27442, n_18791, n_18792);
  and g46139 (n27443, n11727, n27442);
  and g46140 (n27444, n11055, n26890);
  and g46141 (n27445, n11715, n27173);
  not g46142 (n_18793, n27444);
  not g46143 (n_18794, n27445);
  and g46144 (n27446, n_18793, n_18794);
  not g46145 (n_18795, n27443);
  and g46146 (n27447, n_18795, n27446);
  and g46147 (n27448, n_6291, n27447);
  and g46148 (n27449, n_18570, n_18573);
  not g46149 (n_18796, n27442);
  and g46150 (n27450, n_18568, n_18796);
  and g46151 (n27451, n27173, n27442);
  not g46152 (n_18797, n27450);
  not g46153 (n_18798, n27451);
  and g46154 (n27452, n_18797, n_18798);
  not g46155 (n_18799, n27449);
  and g46156 (n27453, n_18799, n27452);
  not g46157 (n_18800, n27452);
  and g46158 (n27454, n27449, n_18800);
  not g46159 (n_18801, n27453);
  not g46160 (n_18802, n27454);
  and g46161 (n27455, n_18801, n_18802);
  not g46162 (n_18803, n27455);
  and g46163 (n27456, n27447, n_18803);
  not g46164 (n_18804, n27448);
  not g46165 (n_18805, n27456);
  and g46166 (n27457, n_18804, n_18805);
  not g46167 (n_18806, n27457);
  and g46168 (n27458, \a[2] , n_18806);
  and g46169 (n27459, n_10, n27457);
  not g46170 (n_18807, n27458);
  not g46171 (n_18808, n27459);
  and g46172 (n27460, n_18807, n_18808);
  not g46173 (n_18809, n27460);
  and g46174 (n27461, n27407, n_18809);
  not g46175 (n_18810, n27407);
  and g46176 (n27462, n_18810, n27460);
  not g46177 (n_18811, n27461);
  not g46178 (n_18812, n27462);
  and g46179 (n27463, n_18811, n_18812);
  not g46180 (n_18813, n27200);
  and g46181 (n27464, n_18813, n27463);
  not g46182 (n_18814, n27463);
  and g46183 (n27465, n27200, n_18814);
  not g46184 (n_18815, n27464);
  not g46185 (n_18816, n27465);
  and g46186 (n27466, n_18815, n_18816);
  and g46187 (n27467, n27197, n27466);
  not g46188 (n_18817, n27466);
  and g46189 (n27468, n_18591, n_18817);
  not g46190 (n_18818, n27467);
  not g46191 (n_18819, n27468);
  and g46192 (\result[2] , n_18818, n_18819);
  and g46193 (n27470, n_18811, n_18815);
  and g46194 (n27471, n71, n26890);
  and g46195 (n27472, n9867, n26066);
  and g46196 (n27473, n10434, n26060);
  not g46202 (n_18823, n26904);
  and g46203 (n27476, n9870, n_18823);
  not g46206 (n_18825, n27477);
  and g46207 (n27478, \a[5] , n_18825);
  not g46208 (n_18826, n27478);
  and g46209 (n27479, n_18825, n_18826);
  and g46210 (n27480, \a[5] , n_18826);
  not g46211 (n_18827, n27479);
  not g46212 (n_18828, n27480);
  and g46213 (n27481, n_18827, n_18828);
  and g46214 (n27482, n_18743, n_18748);
  and g46215 (n27483, n7983, n22312);
  and g46216 (n27484, n7291, n22323);
  and g46217 (n27485, n7632, n22320);
  and g46223 (n27488, n7294, n_17004);
  not g46226 (n_18833, n27489);
  and g46227 (n27490, \a[11] , n_18833);
  not g46228 (n_18834, n27490);
  and g46229 (n27491, n_18833, n_18834);
  and g46230 (n27492, \a[11] , n_18834);
  not g46231 (n_18835, n27491);
  not g46232 (n_18836, n27492);
  and g46233 (n27493, n_18835, n_18836);
  and g46234 (n27494, n_18717, n_18722);
  and g46235 (n27495, n6233, n22335);
  and g46236 (n27496, n5663, n22341);
  and g46237 (n27497, n5939, n22338);
  and g46243 (n27500, n5666, n_16015);
  not g46246 (n_18841, n27501);
  and g46247 (n27502, \a[17] , n_18841);
  not g46248 (n_18842, n27502);
  and g46249 (n27503, n_18841, n_18842);
  and g46250 (n27504, \a[17] , n_18842);
  not g46251 (n_18843, n27503);
  not g46252 (n_18844, n27504);
  and g46253 (n27505, n_18843, n_18844);
  and g46254 (n27506, n_18691, n_18696);
  and g46255 (n27507, n4694, n22353);
  and g46256 (n27508, n4533, n22359);
  and g46257 (n27509, n4604, n22356);
  and g46263 (n27512, n4536, n_14678);
  not g46266 (n_18849, n27513);
  and g46267 (n27514, \a[23] , n_18849);
  not g46268 (n_18850, n27514);
  and g46269 (n27515, n_18849, n_18850);
  and g46270 (n27516, \a[23] , n_18850);
  not g46271 (n_18851, n27515);
  not g46272 (n_18852, n27516);
  and g46273 (n27517, n_18851, n_18852);
  and g46274 (n27518, n_18665, n_18670);
  and g46275 (n27519, n_18650, n_18654);
  and g46276 (n27520, n_18632, n_18637);
  and g46277 (n27521, n156, n2466);
  and g46278 (n27522, n2993, n27521);
  and g46292 (n27536, n3020, n22380);
  and g46293 (n27537, n3028, n22384);
  and g46294 (n27538, n3023, n22387);
  and g46295 (n27539, n75, n22850);
  not g46303 (n_18857, n27535);
  not g46304 (n_18858, n27542);
  and g46305 (n27543, n_18857, n_18858);
  not g46306 (n_18859, n27543);
  and g46307 (n27544, n_18857, n_18859);
  and g46308 (n27545, n_18858, n_18859);
  not g46309 (n_18860, n27544);
  not g46310 (n_18861, n27545);
  and g46311 (n27546, n_18860, n_18861);
  not g46312 (n_18862, n27520);
  not g46313 (n_18863, n27546);
  and g46314 (n27547, n_18862, n_18863);
  not g46315 (n_18864, n27547);
  and g46316 (n27548, n_18862, n_18864);
  and g46317 (n27549, n_18863, n_18864);
  not g46318 (n_18865, n27548);
  not g46319 (n_18866, n27549);
  and g46320 (n27550, n_18865, n_18866);
  and g46321 (n27551, n3457, n22371);
  and g46322 (n27552, n3542, n22377);
  and g46323 (n27553, n3606, n22374);
  not g46324 (n_18867, n27552);
  not g46325 (n_18868, n27553);
  and g46326 (n27554, n_18867, n_18868);
  not g46327 (n_18869, n27551);
  and g46328 (n27555, n_18869, n27554);
  and g46329 (n27556, n_489, n27555);
  and g46330 (n27557, n_18191, n27555);
  not g46331 (n_18870, n27556);
  not g46332 (n_18871, n27557);
  and g46333 (n27558, n_18870, n_18871);
  not g46334 (n_18872, n27558);
  and g46335 (n27559, \a[29] , n_18872);
  and g46336 (n27560, n_15, n27558);
  not g46337 (n_18873, n27559);
  not g46338 (n_18874, n27560);
  and g46339 (n27561, n_18873, n_18874);
  not g46340 (n_18875, n27550);
  not g46341 (n_18876, n27561);
  and g46342 (n27562, n_18875, n_18876);
  and g46343 (n27563, n27550, n27561);
  not g46344 (n_18877, n27562);
  not g46345 (n_18878, n27563);
  and g46346 (n27564, n_18877, n_18878);
  not g46347 (n_18879, n27519);
  and g46348 (n27565, n_18879, n27564);
  not g46349 (n_18880, n27564);
  and g46350 (n27566, n27519, n_18880);
  not g46351 (n_18881, n27565);
  not g46352 (n_18882, n27566);
  and g46353 (n27567, n_18881, n_18882);
  and g46354 (n27568, n3884, n22362);
  and g46355 (n27569, n3967, n22368);
  and g46356 (n27570, n4046, n22365);
  not g46357 (n_18883, n27569);
  not g46358 (n_18884, n27570);
  and g46359 (n27571, n_18883, n_18884);
  not g46360 (n_18885, n27568);
  and g46361 (n27572, n_18885, n27571);
  and g46362 (n27573, n_750, n27572);
  and g46363 (n27574, n23320, n27572);
  not g46364 (n_18886, n27573);
  not g46365 (n_18887, n27574);
  and g46366 (n27575, n_18886, n_18887);
  not g46367 (n_18888, n27575);
  and g46368 (n27576, \a[26] , n_18888);
  and g46369 (n27577, n_33, n27575);
  not g46370 (n_18889, n27576);
  not g46371 (n_18890, n27577);
  and g46372 (n27578, n_18889, n_18890);
  not g46373 (n_18891, n27578);
  and g46374 (n27579, n27567, n_18891);
  not g46375 (n_18892, n27579);
  and g46376 (n27580, n27567, n_18892);
  and g46377 (n27581, n_18891, n_18892);
  not g46378 (n_18893, n27580);
  not g46379 (n_18894, n27581);
  and g46380 (n27582, n_18893, n_18894);
  not g46381 (n_18895, n27518);
  not g46382 (n_18896, n27582);
  and g46383 (n27583, n_18895, n_18896);
  not g46384 (n_18897, n27583);
  and g46385 (n27584, n_18895, n_18897);
  and g46386 (n27585, n_18896, n_18897);
  not g46387 (n_18898, n27584);
  not g46388 (n_18899, n27585);
  and g46389 (n27586, n_18898, n_18899);
  not g46390 (n_18900, n27517);
  not g46391 (n_18901, n27586);
  and g46392 (n27587, n_18900, n_18901);
  not g46393 (n_18902, n27587);
  and g46394 (n27588, n_18900, n_18902);
  and g46395 (n27589, n_18901, n_18902);
  not g46396 (n_18903, n27588);
  not g46397 (n_18904, n27589);
  and g46398 (n27590, n_18903, n_18904);
  and g46399 (n27591, n_18675, n_18681);
  and g46400 (n27592, n27590, n27591);
  not g46401 (n_18905, n27590);
  not g46402 (n_18906, n27591);
  and g46403 (n27593, n_18905, n_18906);
  not g46404 (n_18907, n27592);
  not g46405 (n_18908, n27593);
  and g46406 (n27594, n_18907, n_18908);
  and g46407 (n27595, n5496, n22344);
  and g46408 (n27596, n4935, n22350);
  and g46409 (n27597, n5407, n22347);
  not g46410 (n_18909, n27596);
  not g46411 (n_18910, n27597);
  and g46412 (n27598, n_18909, n_18910);
  not g46413 (n_18911, n27595);
  and g46414 (n27599, n_18911, n27598);
  and g46415 (n27600, n_1011, n27599);
  and g46416 (n27601, n23642, n27599);
  not g46417 (n_18912, n27600);
  not g46418 (n_18913, n27601);
  and g46419 (n27602, n_18912, n_18913);
  not g46420 (n_18914, n27602);
  and g46421 (n27603, \a[20] , n_18914);
  and g46422 (n27604, n_435, n27602);
  not g46423 (n_18915, n27603);
  not g46424 (n_18916, n27604);
  and g46425 (n27605, n_18915, n_18916);
  not g46426 (n_18917, n27605);
  and g46427 (n27606, n27594, n_18917);
  not g46428 (n_18918, n27606);
  and g46429 (n27607, n27594, n_18918);
  and g46430 (n27608, n_18917, n_18918);
  not g46431 (n_18919, n27607);
  not g46432 (n_18920, n27608);
  and g46433 (n27609, n_18919, n_18920);
  not g46434 (n_18921, n27506);
  not g46435 (n_18922, n27609);
  and g46436 (n27610, n_18921, n_18922);
  not g46437 (n_18923, n27610);
  and g46438 (n27611, n_18921, n_18923);
  and g46439 (n27612, n_18922, n_18923);
  not g46440 (n_18924, n27611);
  not g46441 (n_18925, n27612);
  and g46442 (n27613, n_18924, n_18925);
  not g46443 (n_18926, n27505);
  not g46444 (n_18927, n27613);
  and g46445 (n27614, n_18926, n_18927);
  not g46446 (n_18928, n27614);
  and g46447 (n27615, n_18926, n_18928);
  and g46448 (n27616, n_18927, n_18928);
  not g46449 (n_18929, n27615);
  not g46450 (n_18930, n27616);
  and g46451 (n27617, n_18929, n_18930);
  and g46452 (n27618, n_18701, n_18707);
  and g46453 (n27619, n27617, n27618);
  not g46454 (n_18931, n27617);
  not g46455 (n_18932, n27618);
  and g46456 (n27620, n_18931, n_18932);
  not g46457 (n_18933, n27619);
  not g46458 (n_18934, n27620);
  and g46459 (n27621, n_18933, n_18934);
  and g46460 (n27622, n7101, n22326);
  and g46461 (n27623, n6402, n22332);
  and g46462 (n27624, n6951, n22329);
  not g46463 (n_18935, n27623);
  not g46464 (n_18936, n27624);
  and g46465 (n27625, n_18935, n_18936);
  not g46466 (n_18937, n27622);
  and g46467 (n27626, n_18937, n27625);
  and g46468 (n27627, n_1885, n27626);
  and g46469 (n27628, n24616, n27626);
  not g46470 (n_18938, n27627);
  not g46471 (n_18939, n27628);
  and g46472 (n27629, n_18938, n_18939);
  not g46473 (n_18940, n27629);
  and g46474 (n27630, \a[14] , n_18940);
  and g46475 (n27631, n_652, n27629);
  not g46476 (n_18941, n27630);
  not g46477 (n_18942, n27631);
  and g46478 (n27632, n_18941, n_18942);
  not g46479 (n_18943, n27632);
  and g46480 (n27633, n27621, n_18943);
  not g46481 (n_18944, n27633);
  and g46482 (n27634, n27621, n_18944);
  and g46483 (n27635, n_18943, n_18944);
  not g46484 (n_18945, n27634);
  not g46485 (n_18946, n27635);
  and g46486 (n27636, n_18945, n_18946);
  not g46487 (n_18947, n27494);
  not g46488 (n_18948, n27636);
  and g46489 (n27637, n_18947, n_18948);
  not g46490 (n_18949, n27637);
  and g46491 (n27638, n_18947, n_18949);
  and g46492 (n27639, n_18948, n_18949);
  not g46493 (n_18950, n27638);
  not g46494 (n_18951, n27639);
  and g46495 (n27640, n_18950, n_18951);
  not g46496 (n_18952, n27493);
  not g46497 (n_18953, n27640);
  and g46498 (n27641, n_18952, n_18953);
  not g46499 (n_18954, n27641);
  and g46500 (n27642, n_18952, n_18954);
  and g46501 (n27643, n_18953, n_18954);
  not g46502 (n_18955, n27642);
  not g46503 (n_18956, n27643);
  and g46504 (n27644, n_18955, n_18956);
  and g46505 (n27645, n_18727, n_18733);
  and g46506 (n27646, n27644, n27645);
  not g46507 (n_18957, n27644);
  not g46508 (n_18958, n27645);
  and g46509 (n27647, n_18957, n_18958);
  not g46510 (n_18959, n27646);
  not g46511 (n_18960, n27647);
  and g46512 (n27648, n_18959, n_18960);
  and g46513 (n27649, n9331, n26063);
  and g46514 (n27650, n8418, n22315);
  and g46515 (n27651, n8860, n22309);
  not g46516 (n_18961, n27650);
  not g46517 (n_18962, n27651);
  and g46518 (n27652, n_18961, n_18962);
  not g46519 (n_18963, n27649);
  and g46520 (n27653, n_18963, n27652);
  and g46521 (n27654, n_3428, n27653);
  and g46522 (n27655, n26604, n27653);
  not g46523 (n_18964, n27654);
  not g46524 (n_18965, n27655);
  and g46525 (n27656, n_18964, n_18965);
  not g46526 (n_18966, n27656);
  and g46527 (n27657, \a[8] , n_18966);
  and g46528 (n27658, n_1106, n27656);
  not g46529 (n_18967, n27657);
  not g46530 (n_18968, n27658);
  and g46531 (n27659, n_18967, n_18968);
  not g46532 (n_18969, n27659);
  and g46533 (n27660, n27648, n_18969);
  not g46534 (n_18970, n27660);
  and g46535 (n27661, n27648, n_18970);
  and g46536 (n27662, n_18969, n_18970);
  not g46537 (n_18971, n27661);
  not g46538 (n_18972, n27662);
  and g46539 (n27663, n_18971, n_18972);
  not g46540 (n_18973, n27482);
  not g46541 (n_18974, n27663);
  and g46542 (n27664, n_18973, n_18974);
  not g46543 (n_18975, n27664);
  and g46544 (n27665, n_18973, n_18975);
  and g46545 (n27666, n_18974, n_18975);
  not g46546 (n_18976, n27665);
  not g46547 (n_18977, n27666);
  and g46548 (n27667, n_18976, n_18977);
  not g46549 (n_18978, n27481);
  not g46550 (n_18979, n27667);
  and g46551 (n27668, n_18978, n_18979);
  not g46552 (n_18980, n27668);
  and g46553 (n27669, n_18978, n_18980);
  and g46554 (n27670, n_18979, n_18980);
  not g46555 (n_18981, n27669);
  not g46556 (n_18982, n27670);
  and g46557 (n27671, n_18981, n_18982);
  and g46558 (n27672, n_18753, n_18759);
  and g46559 (n27673, n27671, n27672);
  not g46560 (n_18983, n27671);
  not g46561 (n_18984, n27672);
  and g46562 (n27674, n_18983, n_18984);
  not g46563 (n_18985, n27673);
  not g46564 (n_18986, n27674);
  and g46565 (n27675, n_18985, n_18986);
  and g46566 (n27676, n75, n14028);
  and g46567 (n27677, n3020, n_7417);
  and g46568 (n27678, n3023, n_7540);
  and g46569 (n27679, n3028, n13941);
  and g46577 (n27683, n_18772, n_18775);
  not g46578 (n_18991, n27683);
  and g46579 (n27684, n3839, n_18991);
  not g46580 (n_18992, n3839);
  and g46581 (n27685, n_18992, n27683);
  not g46582 (n_18993, n27684);
  not g46583 (n_18994, n27685);
  and g46584 (n27686, n_18993, n_18994);
  not g46585 (n_18995, n27682);
  and g46586 (n27687, n_18995, n27686);
  not g46587 (n_18996, n27687);
  and g46588 (n27688, n_18995, n_18996);
  and g46589 (n27689, n27686, n_18996);
  not g46590 (n_18997, n27688);
  not g46591 (n_18998, n27689);
  and g46592 (n27690, n_18997, n_18998);
  and g46593 (n27691, n_18778, n_18783);
  and g46594 (n27692, n27690, n27691);
  not g46595 (n_18999, n27690);
  not g46596 (n_19000, n27691);
  and g46597 (n27693, n_18999, n_19000);
  not g46598 (n_19001, n27692);
  not g46599 (n_19002, n27693);
  and g46600 (n27694, n_19001, n_19002);
  and g46601 (n27695, n_18787, n_18791);
  not g46602 (n_19003, n27694);
  and g46603 (n27696, n_19003, n27695);
  not g46604 (n_19004, n27695);
  and g46605 (n27697, n27694, n_19004);
  not g46606 (n_19005, n27696);
  not g46607 (n_19006, n27697);
  and g46608 (n27698, n_19005, n_19006);
  and g46609 (n27699, n11727, n27698);
  and g46610 (n27700, n11055, n27173);
  and g46611 (n27701, n11715, n27442);
  not g46612 (n_19007, n27700);
  not g46613 (n_19008, n27701);
  and g46614 (n27702, n_19007, n_19008);
  not g46615 (n_19009, n27699);
  and g46616 (n27703, n_19009, n27702);
  and g46617 (n27704, n_6291, n27703);
  and g46618 (n27705, n_18798, n_18801);
  and g46619 (n27706, n27442, n27698);
  not g46620 (n_19010, n27698);
  and g46621 (n27707, n_18796, n_19010);
  not g46622 (n_19011, n27705);
  not g46623 (n_19012, n27707);
  and g46624 (n27708, n_19011, n_19012);
  not g46625 (n_19013, n27706);
  and g46626 (n27709, n_19013, n27708);
  not g46627 (n_19014, n27709);
  and g46628 (n27710, n_19011, n_19014);
  and g46629 (n27711, n_19013, n_19014);
  and g46630 (n27712, n_19012, n27711);
  not g46631 (n_19015, n27710);
  not g46632 (n_19016, n27712);
  and g46633 (n27713, n_19015, n_19016);
  and g46634 (n27714, n27703, n27713);
  not g46635 (n_19017, n27704);
  not g46636 (n_19018, n27714);
  and g46637 (n27715, n_19017, n_19018);
  not g46638 (n_19019, n27715);
  and g46639 (n27716, \a[2] , n_19019);
  and g46640 (n27717, n_10, n27715);
  not g46641 (n_19020, n27716);
  not g46642 (n_19021, n27717);
  and g46643 (n27718, n_19020, n_19021);
  not g46644 (n_19022, n27718);
  and g46645 (n27719, n27675, n_19022);
  not g46646 (n_19023, n27675);
  and g46647 (n27720, n_19023, n27718);
  not g46648 (n_19024, n27719);
  not g46649 (n_19025, n27720);
  and g46650 (n27721, n_19024, n_19025);
  not g46651 (n_19026, n27470);
  and g46652 (n27722, n_19026, n27721);
  not g46653 (n_19027, n27721);
  and g46654 (n27723, n27470, n_19027);
  not g46655 (n_19028, n27722);
  not g46656 (n_19029, n27723);
  and g46657 (n27724, n_19028, n_19029);
  and g46658 (n27725, n27467, n27724);
  not g46659 (n_19030, n27724);
  and g46660 (n27726, n_18818, n_19030);
  not g46661 (n_19031, n27725);
  not g46662 (n_19032, n27726);
  and g46663 (\result[3] , n_19031, n_19032);
  and g46664 (n27728, n_19024, n_19028);
  and g46665 (n27729, n71, n27173);
  and g46666 (n27730, n9867, n26060);
  and g46667 (n27731, n10434, n26890);
  and g46673 (n27734, n9870, n27185);
  not g46676 (n_19037, n27735);
  and g46677 (n27736, \a[5] , n_19037);
  not g46678 (n_19038, n27736);
  and g46679 (n27737, n_19037, n_19038);
  and g46680 (n27738, \a[5] , n_19038);
  not g46681 (n_19039, n27737);
  not g46682 (n_19040, n27738);
  and g46683 (n27739, n_19039, n_19040);
  and g46684 (n27740, n_18970, n_18975);
  and g46685 (n27741, n7983, n22315);
  and g46686 (n27742, n7291, n22320);
  and g46687 (n27743, n7632, n22312);
  and g46693 (n27746, n7294, n25294);
  not g46696 (n_19045, n27747);
  and g46697 (n27748, \a[11] , n_19045);
  not g46698 (n_19046, n27748);
  and g46699 (n27749, n_19045, n_19046);
  and g46700 (n27750, \a[11] , n_19046);
  not g46701 (n_19047, n27749);
  not g46702 (n_19048, n27750);
  and g46703 (n27751, n_19047, n_19048);
  and g46704 (n27752, n_18944, n_18949);
  and g46705 (n27753, n6233, n22332);
  and g46706 (n27754, n5663, n22338);
  and g46707 (n27755, n5939, n22335);
  and g46713 (n27758, n5666, n22542);
  not g46716 (n_19053, n27759);
  and g46717 (n27760, \a[17] , n_19053);
  not g46718 (n_19054, n27760);
  and g46719 (n27761, n_19053, n_19054);
  and g46720 (n27762, \a[17] , n_19054);
  not g46721 (n_19055, n27761);
  not g46722 (n_19056, n27762);
  and g46723 (n27763, n_19055, n_19056);
  and g46724 (n27764, n_18918, n_18923);
  and g46725 (n27765, n4694, n22350);
  and g46726 (n27766, n4533, n22356);
  and g46727 (n27767, n4604, n22353);
  and g46733 (n27770, n4536, n23672);
  not g46736 (n_19061, n27771);
  and g46737 (n27772, \a[23] , n_19061);
  not g46738 (n_19062, n27772);
  and g46739 (n27773, n_19061, n_19062);
  and g46740 (n27774, \a[23] , n_19062);
  not g46741 (n_19063, n27773);
  not g46742 (n_19064, n27774);
  and g46743 (n27775, n_19063, n_19064);
  and g46744 (n27776, n_18892, n_18897);
  and g46745 (n27777, n_18877, n_18881);
  and g46746 (n27778, n_18859, n_18864);
  and g46776 (n27808, n3020, n22377);
  and g46777 (n27809, n3028, n22380);
  and g46778 (n27810, n3023, n22384);
  not g46779 (n_19065, n22834);
  and g46780 (n27811, n75, n_19065);
  not g46788 (n_19070, n27807);
  not g46789 (n_19071, n27814);
  and g46790 (n27815, n_19070, n_19071);
  not g46791 (n_19072, n27815);
  and g46792 (n27816, n_19070, n_19072);
  and g46793 (n27817, n_19071, n_19072);
  not g46794 (n_19073, n27816);
  not g46795 (n_19074, n27817);
  and g46796 (n27818, n_19073, n_19074);
  not g46797 (n_19075, n27778);
  not g46798 (n_19076, n27818);
  and g46799 (n27819, n_19075, n_19076);
  not g46800 (n_19077, n27819);
  and g46801 (n27820, n_19075, n_19077);
  and g46802 (n27821, n_19076, n_19077);
  not g46803 (n_19078, n27820);
  not g46804 (n_19079, n27821);
  and g46805 (n27822, n_19078, n_19079);
  and g46806 (n27823, n3457, n22368);
  and g46807 (n27824, n3542, n22374);
  and g46808 (n27825, n3606, n22371);
  not g46809 (n_19080, n27824);
  not g46810 (n_19081, n27825);
  and g46811 (n27826, n_19080, n_19081);
  not g46812 (n_19082, n27823);
  and g46813 (n27827, n_19082, n27826);
  and g46814 (n27828, n_489, n27827);
  and g46815 (n27829, n_18422, n27827);
  not g46816 (n_19083, n27828);
  not g46817 (n_19084, n27829);
  and g46818 (n27830, n_19083, n_19084);
  not g46819 (n_19085, n27830);
  and g46820 (n27831, \a[29] , n_19085);
  and g46821 (n27832, n_15, n27830);
  not g46822 (n_19086, n27831);
  not g46823 (n_19087, n27832);
  and g46824 (n27833, n_19086, n_19087);
  not g46825 (n_19088, n27822);
  not g46826 (n_19089, n27833);
  and g46827 (n27834, n_19088, n_19089);
  and g46828 (n27835, n27822, n27833);
  not g46829 (n_19090, n27834);
  not g46830 (n_19091, n27835);
  and g46831 (n27836, n_19090, n_19091);
  not g46832 (n_19092, n27777);
  and g46833 (n27837, n_19092, n27836);
  not g46834 (n_19093, n27836);
  and g46835 (n27838, n27777, n_19093);
  not g46836 (n_19094, n27837);
  not g46837 (n_19095, n27838);
  and g46838 (n27839, n_19094, n_19095);
  and g46839 (n27840, n3884, n22359);
  and g46840 (n27841, n3967, n22365);
  and g46841 (n27842, n4046, n22362);
  not g46842 (n_19096, n27841);
  not g46843 (n_19097, n27842);
  and g46844 (n27843, n_19096, n_19097);
  not g46845 (n_19098, n27840);
  and g46846 (n27844, n_19098, n27843);
  and g46847 (n27845, n_750, n27844);
  and g46848 (n27846, n_15331, n27844);
  not g46849 (n_19099, n27845);
  not g46850 (n_19100, n27846);
  and g46851 (n27847, n_19099, n_19100);
  not g46852 (n_19101, n27847);
  and g46853 (n27848, \a[26] , n_19101);
  and g46854 (n27849, n_33, n27847);
  not g46855 (n_19102, n27848);
  not g46856 (n_19103, n27849);
  and g46857 (n27850, n_19102, n_19103);
  not g46858 (n_19104, n27850);
  and g46859 (n27851, n27839, n_19104);
  not g46860 (n_19105, n27851);
  and g46861 (n27852, n27839, n_19105);
  and g46862 (n27853, n_19104, n_19105);
  not g46863 (n_19106, n27852);
  not g46864 (n_19107, n27853);
  and g46865 (n27854, n_19106, n_19107);
  not g46866 (n_19108, n27776);
  not g46867 (n_19109, n27854);
  and g46868 (n27855, n_19108, n_19109);
  not g46869 (n_19110, n27855);
  and g46870 (n27856, n_19108, n_19110);
  and g46871 (n27857, n_19109, n_19110);
  not g46872 (n_19111, n27856);
  not g46873 (n_19112, n27857);
  and g46874 (n27858, n_19111, n_19112);
  not g46875 (n_19113, n27775);
  not g46876 (n_19114, n27858);
  and g46877 (n27859, n_19113, n_19114);
  not g46878 (n_19115, n27859);
  and g46879 (n27860, n_19113, n_19115);
  and g46880 (n27861, n_19114, n_19115);
  not g46881 (n_19116, n27860);
  not g46882 (n_19117, n27861);
  and g46883 (n27862, n_19116, n_19117);
  and g46884 (n27863, n_18902, n_18908);
  and g46885 (n27864, n27862, n27863);
  not g46886 (n_19118, n27862);
  not g46887 (n_19119, n27863);
  and g46888 (n27865, n_19118, n_19119);
  not g46889 (n_19120, n27864);
  not g46890 (n_19121, n27865);
  and g46891 (n27866, n_19120, n_19121);
  and g46892 (n27867, n5496, n22341);
  and g46893 (n27868, n4935, n22347);
  and g46894 (n27869, n5407, n22344);
  not g46895 (n_19122, n27868);
  not g46896 (n_19123, n27869);
  and g46897 (n27870, n_19122, n_19123);
  not g46898 (n_19124, n27867);
  and g46899 (n27871, n_19124, n27870);
  and g46900 (n27872, n_1011, n27871);
  and g46901 (n27873, n_15990, n27871);
  not g46902 (n_19125, n27872);
  not g46903 (n_19126, n27873);
  and g46904 (n27874, n_19125, n_19126);
  not g46905 (n_19127, n27874);
  and g46906 (n27875, \a[20] , n_19127);
  and g46907 (n27876, n_435, n27874);
  not g46908 (n_19128, n27875);
  not g46909 (n_19129, n27876);
  and g46910 (n27877, n_19128, n_19129);
  not g46911 (n_19130, n27877);
  and g46912 (n27878, n27866, n_19130);
  not g46913 (n_19131, n27878);
  and g46914 (n27879, n27866, n_19131);
  and g46915 (n27880, n_19130, n_19131);
  not g46916 (n_19132, n27879);
  not g46917 (n_19133, n27880);
  and g46918 (n27881, n_19132, n_19133);
  not g46919 (n_19134, n27764);
  not g46920 (n_19135, n27881);
  and g46921 (n27882, n_19134, n_19135);
  not g46922 (n_19136, n27882);
  and g46923 (n27883, n_19134, n_19136);
  and g46924 (n27884, n_19135, n_19136);
  not g46925 (n_19137, n27883);
  not g46926 (n_19138, n27884);
  and g46927 (n27885, n_19137, n_19138);
  not g46928 (n_19139, n27763);
  not g46929 (n_19140, n27885);
  and g46930 (n27886, n_19139, n_19140);
  not g46931 (n_19141, n27886);
  and g46932 (n27887, n_19139, n_19141);
  and g46933 (n27888, n_19140, n_19141);
  not g46934 (n_19142, n27887);
  not g46935 (n_19143, n27888);
  and g46936 (n27889, n_19142, n_19143);
  and g46937 (n27890, n_18928, n_18934);
  and g46938 (n27891, n27889, n27890);
  not g46939 (n_19144, n27889);
  not g46940 (n_19145, n27890);
  and g46941 (n27892, n_19144, n_19145);
  not g46942 (n_19146, n27891);
  not g46943 (n_19147, n27892);
  and g46944 (n27893, n_19146, n_19147);
  and g46945 (n27894, n7101, n22323);
  and g46946 (n27895, n6402, n22329);
  and g46947 (n27896, n6951, n22326);
  not g46948 (n_19148, n27895);
  not g46949 (n_19149, n27896);
  and g46950 (n27897, n_19148, n_19149);
  not g46951 (n_19150, n27894);
  and g46952 (n27898, n_19150, n27897);
  and g46953 (n27899, n_1885, n27898);
  and g46954 (n27900, n_16393, n27898);
  not g46955 (n_19151, n27899);
  not g46956 (n_19152, n27900);
  and g46957 (n27901, n_19151, n_19152);
  not g46958 (n_19153, n27901);
  and g46959 (n27902, \a[14] , n_19153);
  and g46960 (n27903, n_652, n27901);
  not g46961 (n_19154, n27902);
  not g46962 (n_19155, n27903);
  and g46963 (n27904, n_19154, n_19155);
  not g46964 (n_19156, n27904);
  and g46965 (n27905, n27893, n_19156);
  not g46966 (n_19157, n27905);
  and g46967 (n27906, n27893, n_19157);
  and g46968 (n27907, n_19156, n_19157);
  not g46969 (n_19158, n27906);
  not g46970 (n_19159, n27907);
  and g46971 (n27908, n_19158, n_19159);
  not g46972 (n_19160, n27752);
  not g46973 (n_19161, n27908);
  and g46974 (n27909, n_19160, n_19161);
  not g46975 (n_19162, n27909);
  and g46976 (n27910, n_19160, n_19162);
  and g46977 (n27911, n_19161, n_19162);
  not g46978 (n_19163, n27910);
  not g46979 (n_19164, n27911);
  and g46980 (n27912, n_19163, n_19164);
  not g46981 (n_19165, n27751);
  not g46982 (n_19166, n27912);
  and g46983 (n27913, n_19165, n_19166);
  not g46984 (n_19167, n27913);
  and g46985 (n27914, n_19165, n_19167);
  and g46986 (n27915, n_19166, n_19167);
  not g46987 (n_19168, n27914);
  not g46988 (n_19169, n27915);
  and g46989 (n27916, n_19168, n_19169);
  and g46990 (n27917, n_18954, n_18960);
  and g46991 (n27918, n27916, n27917);
  not g46992 (n_19170, n27916);
  not g46993 (n_19171, n27917);
  and g46994 (n27919, n_19170, n_19171);
  not g46995 (n_19172, n27918);
  not g46996 (n_19173, n27919);
  and g46997 (n27920, n_19172, n_19173);
  and g46998 (n27921, n9331, n26066);
  and g46999 (n27922, n8418, n22309);
  and g47000 (n27923, n8860, n26063);
  not g47001 (n_19174, n27922);
  not g47002 (n_19175, n27923);
  and g47003 (n27924, n_19174, n_19175);
  not g47004 (n_19176, n27921);
  and g47005 (n27925, n_19176, n27924);
  and g47006 (n27926, n_3428, n27925);
  and g47007 (n27927, n26624, n27925);
  not g47008 (n_19177, n27926);
  not g47009 (n_19178, n27927);
  and g47010 (n27928, n_19177, n_19178);
  not g47011 (n_19179, n27928);
  and g47012 (n27929, \a[8] , n_19179);
  and g47013 (n27930, n_1106, n27928);
  not g47014 (n_19180, n27929);
  not g47015 (n_19181, n27930);
  and g47016 (n27931, n_19180, n_19181);
  not g47017 (n_19182, n27931);
  and g47018 (n27932, n27920, n_19182);
  not g47019 (n_19183, n27932);
  and g47020 (n27933, n27920, n_19183);
  and g47021 (n27934, n_19182, n_19183);
  not g47022 (n_19184, n27933);
  not g47023 (n_19185, n27934);
  and g47024 (n27935, n_19184, n_19185);
  not g47025 (n_19186, n27740);
  not g47026 (n_19187, n27935);
  and g47027 (n27936, n_19186, n_19187);
  not g47028 (n_19188, n27936);
  and g47029 (n27937, n_19186, n_19188);
  and g47030 (n27938, n_19187, n_19188);
  not g47031 (n_19189, n27937);
  not g47032 (n_19190, n27938);
  and g47033 (n27939, n_19189, n_19190);
  not g47034 (n_19191, n27739);
  not g47035 (n_19192, n27939);
  and g47036 (n27940, n_19191, n_19192);
  not g47037 (n_19193, n27940);
  and g47038 (n27941, n_19191, n_19193);
  and g47039 (n27942, n_19192, n_19193);
  not g47040 (n_19194, n27941);
  not g47041 (n_19195, n27942);
  and g47042 (n27943, n_19194, n_19195);
  and g47043 (n27944, n_18980, n_18986);
  and g47044 (n27945, n27943, n27944);
  not g47045 (n_19196, n27943);
  not g47046 (n_19197, n27944);
  and g47047 (n27946, n_19196, n_19197);
  not g47048 (n_19198, n27945);
  not g47049 (n_19199, n27946);
  and g47050 (n27947, n_19198, n_19199);
  and g47051 (n27948, n75, n_13153);
  not g47052 (n_19200, n3028);
  and g47053 (n27949, n_2598, n_19200);
  not g47054 (n_19201, n27949);
  and g47055 (n27950, n_7417, n_19201);
  and g47056 (n27951, n3023, n13941);
  not g47057 (n_19202, n27950);
  not g47058 (n_19203, n27951);
  and g47059 (n27952, n_19202, n_19203);
  not g47060 (n_19204, n27948);
  and g47061 (n27953, n_19204, n27952);
  and g47062 (n27954, n3839, n27953);
  not g47063 (n_19205, n27953);
  and g47064 (n27955, n_18992, n_19205);
  not g47065 (n_19206, n27954);
  not g47066 (n_19207, n27955);
  and g47067 (n27956, n_19206, n_19207);
  and g47068 (n27957, n_18993, n_18996);
  and g47069 (n27958, n27956, n27957);
  not g47070 (n_19208, n27956);
  not g47071 (n_19209, n27957);
  and g47072 (n27959, n_19208, n_19209);
  not g47073 (n_19210, n27958);
  not g47074 (n_19211, n27959);
  and g47075 (n27960, n_19210, n_19211);
  and g47076 (n27961, n_19002, n_19006);
  not g47077 (n_19212, n27960);
  and g47078 (n27962, n_19212, n27961);
  not g47079 (n_19213, n27961);
  and g47080 (n27963, n27960, n_19213);
  not g47081 (n_19214, n27962);
  not g47082 (n_19215, n27963);
  and g47083 (n27964, n_19214, n_19215);
  and g47084 (n27965, n11727, n27964);
  and g47085 (n27966, n11055, n27442);
  and g47086 (n27967, n11715, n27698);
  not g47087 (n_19216, n27966);
  not g47088 (n_19217, n27967);
  and g47089 (n27968, n_19216, n_19217);
  not g47090 (n_19218, n27965);
  and g47091 (n27969, n_19218, n27968);
  and g47092 (n27970, n_6291, n27969);
  not g47093 (n_19219, n27964);
  and g47094 (n27971, n_19010, n_19219);
  and g47095 (n27972, n27698, n27964);
  not g47096 (n_19220, n27971);
  not g47097 (n_19221, n27972);
  and g47098 (n27973, n_19220, n_19221);
  not g47099 (n_19222, n27711);
  and g47100 (n27974, n_19222, n27973);
  not g47101 (n_19223, n27973);
  and g47102 (n27975, n27711, n_19223);
  not g47103 (n_19224, n27974);
  not g47104 (n_19225, n27975);
  and g47105 (n27976, n_19224, n_19225);
  not g47106 (n_19226, n27976);
  and g47107 (n27977, n27969, n_19226);
  not g47108 (n_19227, n27970);
  not g47109 (n_19228, n27977);
  and g47110 (n27978, n_19227, n_19228);
  not g47111 (n_19229, n27978);
  and g47112 (n27979, \a[2] , n_19229);
  and g47113 (n27980, n_10, n27978);
  not g47114 (n_19230, n27979);
  not g47115 (n_19231, n27980);
  and g47116 (n27981, n_19230, n_19231);
  not g47117 (n_19232, n27981);
  and g47118 (n27982, n27947, n_19232);
  not g47119 (n_19233, n27947);
  and g47120 (n27983, n_19233, n27981);
  not g47121 (n_19234, n27982);
  not g47122 (n_19235, n27983);
  and g47123 (n27984, n_19234, n_19235);
  not g47124 (n_19236, n27728);
  and g47125 (n27985, n_19236, n27984);
  not g47126 (n_19237, n27984);
  and g47127 (n27986, n27728, n_19237);
  not g47128 (n_19238, n27985);
  not g47129 (n_19239, n27986);
  and g47130 (n27987, n_19238, n_19239);
  and g47131 (n27988, n27725, n27987);
  not g47132 (n_19240, n27987);
  and g47133 (n27989, n_19031, n_19240);
  not g47134 (n_19241, n27988);
  not g47135 (n_19242, n27989);
  and g47136 (\result[4] , n_19241, n_19242);
  and g47137 (n27991, n_19234, n_19238);
  and g47138 (n27992, n71, n27442);
  and g47139 (n27993, n9867, n26890);
  and g47140 (n27994, n10434, n27173);
  and g47146 (n27997, n9870, n27455);
  not g47149 (n_19247, n27998);
  and g47150 (n27999, \a[5] , n_19247);
  not g47151 (n_19248, n27999);
  and g47152 (n28000, n_19247, n_19248);
  and g47153 (n28001, \a[5] , n_19248);
  not g47154 (n_19249, n28000);
  not g47155 (n_19250, n28001);
  and g47156 (n28002, n_19249, n_19250);
  and g47157 (n28003, n_19183, n_19188);
  and g47158 (n28004, n7983, n22309);
  and g47159 (n28005, n7291, n22312);
  and g47160 (n28006, n7632, n22315);
  and g47166 (n28009, n7294, n_14657);
  not g47169 (n_19255, n28010);
  and g47170 (n28011, \a[11] , n_19255);
  not g47171 (n_19256, n28011);
  and g47172 (n28012, n_19255, n_19256);
  and g47173 (n28013, \a[11] , n_19256);
  not g47174 (n_19257, n28012);
  not g47175 (n_19258, n28013);
  and g47176 (n28014, n_19257, n_19258);
  and g47177 (n28015, n_19157, n_19162);
  and g47178 (n28016, n6233, n22329);
  and g47179 (n28017, n5663, n22335);
  and g47180 (n28018, n5939, n22332);
  and g47186 (n28021, n5666, n_16827);
  not g47189 (n_19263, n28022);
  and g47190 (n28023, \a[17] , n_19263);
  not g47191 (n_19264, n28023);
  and g47192 (n28024, n_19263, n_19264);
  and g47193 (n28025, \a[17] , n_19264);
  not g47194 (n_19265, n28024);
  not g47195 (n_19266, n28025);
  and g47196 (n28026, n_19265, n_19266);
  and g47197 (n28027, n_19131, n_19136);
  and g47198 (n28028, n4694, n22347);
  and g47199 (n28029, n4533, n22353);
  and g47200 (n28030, n4604, n22350);
  and g47206 (n28033, n4536, n_16069);
  not g47209 (n_19271, n28034);
  and g47210 (n28035, \a[23] , n_19271);
  not g47211 (n_19272, n28035);
  and g47212 (n28036, n_19271, n_19272);
  and g47213 (n28037, \a[23] , n_19272);
  not g47214 (n_19273, n28036);
  not g47215 (n_19274, n28037);
  and g47216 (n28038, n_19273, n_19274);
  and g47217 (n28039, n_19105, n_19110);
  and g47218 (n28040, n_19090, n_19094);
  and g47219 (n28041, n_19072, n_19077);
  and g47238 (n28060, n3020, n22374);
  and g47239 (n28061, n3028, n22377);
  and g47240 (n28062, n3023, n22380);
  and g47241 (n28063, n75, n22569);
  not g47249 (n_19279, n28059);
  not g47250 (n_19280, n28066);
  and g47251 (n28067, n_19279, n_19280);
  not g47252 (n_19281, n28067);
  and g47253 (n28068, n_19279, n_19281);
  and g47254 (n28069, n_19280, n_19281);
  not g47255 (n_19282, n28068);
  not g47256 (n_19283, n28069);
  and g47257 (n28070, n_19282, n_19283);
  not g47258 (n_19284, n28041);
  not g47259 (n_19285, n28070);
  and g47260 (n28071, n_19284, n_19285);
  not g47261 (n_19286, n28071);
  and g47262 (n28072, n_19284, n_19286);
  and g47263 (n28073, n_19285, n_19286);
  not g47264 (n_19287, n28072);
  not g47265 (n_19288, n28073);
  and g47266 (n28074, n_19287, n_19288);
  and g47267 (n28075, n3457, n22365);
  and g47268 (n28076, n3542, n22371);
  and g47269 (n28077, n3606, n22368);
  not g47270 (n_19289, n28076);
  not g47271 (n_19290, n28077);
  and g47272 (n28078, n_19289, n_19290);
  not g47273 (n_19291, n28075);
  and g47274 (n28079, n_19291, n28078);
  and g47275 (n28080, n_489, n28079);
  and g47276 (n28081, n22993, n28079);
  not g47277 (n_19292, n28080);
  not g47278 (n_19293, n28081);
  and g47279 (n28082, n_19292, n_19293);
  not g47280 (n_19294, n28082);
  and g47281 (n28083, \a[29] , n_19294);
  and g47282 (n28084, n_15, n28082);
  not g47283 (n_19295, n28083);
  not g47284 (n_19296, n28084);
  and g47285 (n28085, n_19295, n_19296);
  not g47286 (n_19297, n28074);
  not g47287 (n_19298, n28085);
  and g47288 (n28086, n_19297, n_19298);
  and g47289 (n28087, n28074, n28085);
  not g47290 (n_19299, n28086);
  not g47291 (n_19300, n28087);
  and g47292 (n28088, n_19299, n_19300);
  not g47293 (n_19301, n28040);
  and g47294 (n28089, n_19301, n28088);
  not g47295 (n_19302, n28088);
  and g47296 (n28090, n28040, n_19302);
  not g47297 (n_19303, n28089);
  not g47298 (n_19304, n28090);
  and g47299 (n28091, n_19303, n_19304);
  and g47300 (n28092, n3884, n22356);
  and g47301 (n28093, n3967, n22362);
  and g47302 (n28094, n4046, n22359);
  not g47303 (n_19305, n28093);
  not g47304 (n_19306, n28094);
  and g47305 (n28095, n_19305, n_19306);
  not g47306 (n_19307, n28092);
  and g47307 (n28096, n_19307, n28095);
  and g47308 (n28097, n_750, n28096);
  and g47309 (n28098, n23345, n28096);
  not g47310 (n_19308, n28097);
  not g47311 (n_19309, n28098);
  and g47312 (n28099, n_19308, n_19309);
  not g47313 (n_19310, n28099);
  and g47314 (n28100, \a[26] , n_19310);
  and g47315 (n28101, n_33, n28099);
  not g47316 (n_19311, n28100);
  not g47317 (n_19312, n28101);
  and g47318 (n28102, n_19311, n_19312);
  not g47319 (n_19313, n28102);
  and g47320 (n28103, n28091, n_19313);
  not g47321 (n_19314, n28103);
  and g47322 (n28104, n28091, n_19314);
  and g47323 (n28105, n_19313, n_19314);
  not g47324 (n_19315, n28104);
  not g47325 (n_19316, n28105);
  and g47326 (n28106, n_19315, n_19316);
  not g47327 (n_19317, n28039);
  not g47328 (n_19318, n28106);
  and g47329 (n28107, n_19317, n_19318);
  not g47330 (n_19319, n28107);
  and g47331 (n28108, n_19317, n_19319);
  and g47332 (n28109, n_19318, n_19319);
  not g47333 (n_19320, n28108);
  not g47334 (n_19321, n28109);
  and g47335 (n28110, n_19320, n_19321);
  not g47336 (n_19322, n28038);
  not g47337 (n_19323, n28110);
  and g47338 (n28111, n_19322, n_19323);
  not g47339 (n_19324, n28111);
  and g47340 (n28112, n_19322, n_19324);
  and g47341 (n28113, n_19323, n_19324);
  not g47342 (n_19325, n28112);
  not g47343 (n_19326, n28113);
  and g47344 (n28114, n_19325, n_19326);
  and g47345 (n28115, n_19115, n_19121);
  and g47346 (n28116, n28114, n28115);
  not g47347 (n_19327, n28114);
  not g47348 (n_19328, n28115);
  and g47349 (n28117, n_19327, n_19328);
  not g47350 (n_19329, n28116);
  not g47351 (n_19330, n28117);
  and g47352 (n28118, n_19329, n_19330);
  and g47353 (n28119, n5496, n22338);
  and g47354 (n28120, n4935, n22344);
  and g47355 (n28121, n5407, n22341);
  not g47356 (n_19331, n28120);
  not g47357 (n_19332, n28121);
  and g47358 (n28122, n_19331, n_19332);
  not g47359 (n_19333, n28119);
  and g47360 (n28123, n_19333, n28122);
  and g47361 (n28124, n_1011, n28123);
  and g47362 (n28125, n24188, n28123);
  not g47363 (n_19334, n28124);
  not g47364 (n_19335, n28125);
  and g47365 (n28126, n_19334, n_19335);
  not g47366 (n_19336, n28126);
  and g47367 (n28127, \a[20] , n_19336);
  and g47368 (n28128, n_435, n28126);
  not g47369 (n_19337, n28127);
  not g47370 (n_19338, n28128);
  and g47371 (n28129, n_19337, n_19338);
  not g47372 (n_19339, n28129);
  and g47373 (n28130, n28118, n_19339);
  not g47374 (n_19340, n28130);
  and g47375 (n28131, n28118, n_19340);
  and g47376 (n28132, n_19339, n_19340);
  not g47377 (n_19341, n28131);
  not g47378 (n_19342, n28132);
  and g47379 (n28133, n_19341, n_19342);
  not g47380 (n_19343, n28027);
  not g47381 (n_19344, n28133);
  and g47382 (n28134, n_19343, n_19344);
  not g47383 (n_19345, n28134);
  and g47384 (n28135, n_19343, n_19345);
  and g47385 (n28136, n_19344, n_19345);
  not g47386 (n_19346, n28135);
  not g47387 (n_19347, n28136);
  and g47388 (n28137, n_19346, n_19347);
  not g47389 (n_19348, n28026);
  not g47390 (n_19349, n28137);
  and g47391 (n28138, n_19348, n_19349);
  not g47392 (n_19350, n28138);
  and g47393 (n28139, n_19348, n_19350);
  and g47394 (n28140, n_19349, n_19350);
  not g47395 (n_19351, n28139);
  not g47396 (n_19352, n28140);
  and g47397 (n28141, n_19351, n_19352);
  and g47398 (n28142, n_19141, n_19147);
  and g47399 (n28143, n28141, n28142);
  not g47400 (n_19353, n28141);
  not g47401 (n_19354, n28142);
  and g47402 (n28144, n_19353, n_19354);
  not g47403 (n_19355, n28143);
  not g47404 (n_19356, n28144);
  and g47405 (n28145, n_19355, n_19356);
  and g47406 (n28146, n7101, n22320);
  and g47407 (n28147, n6402, n22326);
  and g47408 (n28148, n6951, n22323);
  not g47409 (n_19357, n28147);
  not g47410 (n_19358, n28148);
  and g47411 (n28149, n_19357, n_19358);
  not g47412 (n_19359, n28146);
  and g47413 (n28150, n_19359, n28149);
  and g47414 (n28151, n_1885, n28150);
  and g47415 (n28152, n25270, n28150);
  not g47416 (n_19360, n28151);
  not g47417 (n_19361, n28152);
  and g47418 (n28153, n_19360, n_19361);
  not g47419 (n_19362, n28153);
  and g47420 (n28154, \a[14] , n_19362);
  and g47421 (n28155, n_652, n28153);
  not g47422 (n_19363, n28154);
  not g47423 (n_19364, n28155);
  and g47424 (n28156, n_19363, n_19364);
  not g47425 (n_19365, n28156);
  and g47426 (n28157, n28145, n_19365);
  not g47427 (n_19366, n28157);
  and g47428 (n28158, n28145, n_19366);
  and g47429 (n28159, n_19365, n_19366);
  not g47430 (n_19367, n28158);
  not g47431 (n_19368, n28159);
  and g47432 (n28160, n_19367, n_19368);
  not g47433 (n_19369, n28015);
  not g47434 (n_19370, n28160);
  and g47435 (n28161, n_19369, n_19370);
  not g47436 (n_19371, n28161);
  and g47437 (n28162, n_19369, n_19371);
  and g47438 (n28163, n_19370, n_19371);
  not g47439 (n_19372, n28162);
  not g47440 (n_19373, n28163);
  and g47441 (n28164, n_19372, n_19373);
  not g47442 (n_19374, n28014);
  not g47443 (n_19375, n28164);
  and g47444 (n28165, n_19374, n_19375);
  not g47445 (n_19376, n28165);
  and g47446 (n28166, n_19374, n_19376);
  and g47447 (n28167, n_19375, n_19376);
  not g47448 (n_19377, n28166);
  not g47449 (n_19378, n28167);
  and g47450 (n28168, n_19377, n_19378);
  and g47451 (n28169, n_19167, n_19173);
  and g47452 (n28170, n28168, n28169);
  not g47453 (n_19379, n28168);
  not g47454 (n_19380, n28169);
  and g47455 (n28171, n_19379, n_19380);
  not g47456 (n_19381, n28170);
  not g47457 (n_19382, n28171);
  and g47458 (n28172, n_19381, n_19382);
  and g47459 (n28173, n9331, n26060);
  and g47460 (n28174, n8418, n26063);
  and g47461 (n28175, n8860, n26066);
  not g47462 (n_19383, n28174);
  not g47463 (n_19384, n28175);
  and g47464 (n28176, n_19383, n_19384);
  not g47465 (n_19385, n28173);
  and g47466 (n28177, n_19385, n28176);
  and g47467 (n28178, n_3428, n28177);
  and g47468 (n28179, n26088, n28177);
  not g47469 (n_19386, n28178);
  not g47470 (n_19387, n28179);
  and g47471 (n28180, n_19386, n_19387);
  not g47472 (n_19388, n28180);
  and g47473 (n28181, \a[8] , n_19388);
  and g47474 (n28182, n_1106, n28180);
  not g47475 (n_19389, n28181);
  not g47476 (n_19390, n28182);
  and g47477 (n28183, n_19389, n_19390);
  not g47478 (n_19391, n28183);
  and g47479 (n28184, n28172, n_19391);
  not g47480 (n_19392, n28184);
  and g47481 (n28185, n28172, n_19392);
  and g47482 (n28186, n_19391, n_19392);
  not g47483 (n_19393, n28185);
  not g47484 (n_19394, n28186);
  and g47485 (n28187, n_19393, n_19394);
  not g47486 (n_19395, n28003);
  not g47487 (n_19396, n28187);
  and g47488 (n28188, n_19395, n_19396);
  not g47489 (n_19397, n28188);
  and g47490 (n28189, n_19395, n_19397);
  and g47491 (n28190, n_19396, n_19397);
  not g47492 (n_19398, n28189);
  not g47493 (n_19399, n28190);
  and g47494 (n28191, n_19398, n_19399);
  not g47495 (n_19400, n28002);
  not g47496 (n_19401, n28191);
  and g47497 (n28192, n_19400, n_19401);
  not g47498 (n_19402, n28192);
  and g47499 (n28193, n_19400, n_19402);
  and g47500 (n28194, n_19401, n_19402);
  not g47501 (n_19403, n28193);
  not g47502 (n_19404, n28194);
  and g47503 (n28195, n_19403, n_19404);
  and g47504 (n28196, n_19193, n_19199);
  and g47505 (n28197, n28195, n28196);
  not g47506 (n_19405, n28195);
  not g47507 (n_19406, n28196);
  and g47508 (n28198, n_19405, n_19406);
  not g47509 (n_19407, n28197);
  not g47510 (n_19408, n28198);
  and g47511 (n28199, n_19407, n_19408);
  and g47512 (n28200, n_19211, n_19215);
  and g47513 (n28201, n_422, n97);
  not g47514 (n_19409, n28201);
  and g47515 (n28202, n_7417, n_19409);
  not g47516 (n_19410, n28202);
  and g47517 (n28203, n27954, n_19410);
  and g47518 (n28204, n_19206, n28202);
  not g47519 (n_19411, n28203);
  not g47520 (n_19412, n28204);
  and g47521 (n28205, n_19411, n_19412);
  not g47522 (n_19413, n28205);
  and g47523 (n28206, n28200, n_19413);
  not g47524 (n_19414, n28200);
  and g47525 (n28207, n_19414, n28205);
  not g47526 (n_19415, n28206);
  not g47527 (n_19416, n28207);
  and g47528 (n28208, n_19415, n_19416);
  not g47529 (n_19417, n28208);
  and g47530 (n28209, n11727, n_19417);
  and g47531 (n28210, n11055, n27698);
  and g47532 (n28211, n11715, n27964);
  not g47533 (n_19418, n28210);
  not g47534 (n_19419, n28211);
  and g47535 (n28212, n_19418, n_19419);
  not g47536 (n_19420, n28209);
  and g47537 (n28213, n_19420, n28212);
  and g47538 (n28214, n_6291, n28213);
  and g47539 (n28215, n_19221, n_19224);
  and g47540 (n28216, n27964, n_19417);
  and g47541 (n28217, n_19219, n28208);
  not g47542 (n_19421, n28215);
  not g47543 (n_19422, n28217);
  and g47544 (n28218, n_19421, n_19422);
  not g47545 (n_19423, n28216);
  and g47546 (n28219, n_19423, n28218);
  not g47547 (n_19424, n28219);
  and g47548 (n28220, n_19421, n_19424);
  and g47549 (n28221, n_19423, n_19424);
  and g47550 (n28222, n_19422, n28221);
  not g47551 (n_19425, n28220);
  not g47552 (n_19426, n28222);
  and g47553 (n28223, n_19425, n_19426);
  and g47554 (n28224, n28213, n28223);
  not g47555 (n_19427, n28214);
  not g47556 (n_19428, n28224);
  and g47557 (n28225, n_19427, n_19428);
  not g47558 (n_19429, n28225);
  and g47559 (n28226, \a[2] , n_19429);
  and g47560 (n28227, n_10, n28225);
  not g47561 (n_19430, n28226);
  not g47562 (n_19431, n28227);
  and g47563 (n28228, n_19430, n_19431);
  not g47564 (n_19432, n28228);
  and g47565 (n28229, n28199, n_19432);
  not g47566 (n_19433, n28199);
  and g47567 (n28230, n_19433, n28228);
  not g47568 (n_19434, n28229);
  not g47569 (n_19435, n28230);
  and g47570 (n28231, n_19434, n_19435);
  not g47571 (n_19436, n27991);
  and g47572 (n28232, n_19436, n28231);
  not g47573 (n_19437, n28231);
  and g47574 (n28233, n27991, n_19437);
  not g47575 (n_19438, n28232);
  not g47576 (n_19439, n28233);
  and g47577 (n28234, n_19438, n_19439);
  and g47578 (n28235, n27988, n28234);
  not g47579 (n_19440, n28234);
  and g47580 (n28236, n_19241, n_19440);
  not g47581 (n_19441, n28235);
  not g47582 (n_19442, n28236);
  and g47583 (\result[5] , n_19441, n_19442);
  and g47584 (n28238, n71, n27698);
  and g47585 (n28239, n9867, n27173);
  and g47586 (n28240, n10434, n27442);
  not g47592 (n_19446, n27713);
  and g47593 (n28243, n9870, n_19446);
  not g47596 (n_19448, n28244);
  and g47597 (n28245, \a[5] , n_19448);
  not g47598 (n_19449, n28245);
  and g47599 (n28246, n_19448, n_19449);
  and g47600 (n28247, \a[5] , n_19449);
  not g47601 (n_19450, n28246);
  not g47602 (n_19451, n28247);
  and g47603 (n28248, n_19450, n_19451);
  and g47604 (n28249, n_19392, n_19397);
  and g47605 (n28250, n7983, n26063);
  and g47606 (n28251, n7291, n22315);
  and g47607 (n28252, n7632, n22309);
  and g47613 (n28255, n7294, n_18124);
  not g47616 (n_19456, n28256);
  and g47617 (n28257, \a[11] , n_19456);
  not g47618 (n_19457, n28257);
  and g47619 (n28258, n_19456, n_19457);
  and g47620 (n28259, \a[11] , n_19457);
  not g47621 (n_19458, n28258);
  not g47622 (n_19459, n28259);
  and g47623 (n28260, n_19458, n_19459);
  and g47624 (n28261, n_19366, n_19371);
  and g47625 (n28262, n6233, n22326);
  and g47626 (n28263, n5663, n22332);
  and g47627 (n28264, n5939, n22329);
  and g47633 (n28267, n5666, n_18133);
  not g47636 (n_19464, n28268);
  and g47637 (n28269, \a[17] , n_19464);
  not g47638 (n_19465, n28269);
  and g47639 (n28270, n_19464, n_19465);
  and g47640 (n28271, \a[17] , n_19465);
  not g47641 (n_19466, n28270);
  not g47642 (n_19467, n28271);
  and g47643 (n28272, n_19466, n_19467);
  and g47644 (n28273, n_19340, n_19345);
  and g47645 (n28274, n4694, n22344);
  and g47646 (n28275, n4533, n22350);
  and g47647 (n28276, n4604, n22347);
  and g47653 (n28279, n4536, n_18142);
  not g47656 (n_19472, n28280);
  and g47657 (n28281, \a[23] , n_19472);
  not g47658 (n_19473, n28281);
  and g47659 (n28282, n_19472, n_19473);
  and g47660 (n28283, \a[23] , n_19473);
  not g47661 (n_19474, n28282);
  not g47662 (n_19475, n28283);
  and g47663 (n28284, n_19474, n_19475);
  and g47664 (n28285, n_19314, n_19319);
  and g47665 (n28286, n_19299, n_19303);
  and g47666 (n28287, n_19281, n_19286);
  and g47694 (n28315, n3020, n22371);
  and g47695 (n28316, n3028, n22374);
  and g47696 (n28317, n3023, n22377);
  and g47697 (n28318, n75, n23025);
  not g47705 (n_19480, n28314);
  not g47706 (n_19481, n28321);
  and g47707 (n28322, n_19480, n_19481);
  not g47708 (n_19482, n28322);
  and g47709 (n28323, n_19480, n_19482);
  and g47710 (n28324, n_19481, n_19482);
  not g47711 (n_19483, n28323);
  not g47712 (n_19484, n28324);
  and g47713 (n28325, n_19483, n_19484);
  not g47714 (n_19485, n28287);
  not g47715 (n_19486, n28325);
  and g47716 (n28326, n_19485, n_19486);
  not g47717 (n_19487, n28326);
  and g47718 (n28327, n_19485, n_19487);
  and g47719 (n28328, n_19486, n_19487);
  not g47720 (n_19488, n28327);
  not g47721 (n_19489, n28328);
  and g47722 (n28329, n_19488, n_19489);
  and g47723 (n28330, n3457, n22362);
  and g47724 (n28331, n3542, n22368);
  and g47725 (n28332, n3606, n22365);
  not g47726 (n_19490, n28331);
  not g47727 (n_19491, n28332);
  and g47728 (n28333, n_19490, n_19491);
  not g47729 (n_19492, n28330);
  and g47730 (n28334, n_19492, n28333);
  and g47731 (n28335, n_489, n28334);
  and g47732 (n28336, n23320, n28334);
  not g47733 (n_19493, n28335);
  not g47734 (n_19494, n28336);
  and g47735 (n28337, n_19493, n_19494);
  not g47736 (n_19495, n28337);
  and g47737 (n28338, \a[29] , n_19495);
  and g47738 (n28339, n_15, n28337);
  not g47739 (n_19496, n28338);
  not g47740 (n_19497, n28339);
  and g47741 (n28340, n_19496, n_19497);
  not g47742 (n_19498, n28329);
  not g47743 (n_19499, n28340);
  and g47744 (n28341, n_19498, n_19499);
  and g47745 (n28342, n28329, n28340);
  not g47746 (n_19500, n28341);
  not g47747 (n_19501, n28342);
  and g47748 (n28343, n_19500, n_19501);
  not g47749 (n_19502, n28286);
  and g47750 (n28344, n_19502, n28343);
  not g47751 (n_19503, n28343);
  and g47752 (n28345, n28286, n_19503);
  not g47753 (n_19504, n28344);
  not g47754 (n_19505, n28345);
  and g47755 (n28346, n_19504, n_19505);
  and g47756 (n28347, n3884, n22353);
  and g47757 (n28348, n3967, n22359);
  and g47758 (n28349, n4046, n22356);
  not g47759 (n_19506, n28348);
  not g47760 (n_19507, n28349);
  and g47761 (n28350, n_19506, n_19507);
  not g47762 (n_19508, n28347);
  and g47763 (n28351, n_19508, n28350);
  and g47764 (n28352, n_750, n28351);
  and g47765 (n28353, n22556, n28351);
  not g47766 (n_19509, n28352);
  not g47767 (n_19510, n28353);
  and g47768 (n28354, n_19509, n_19510);
  not g47769 (n_19511, n28354);
  and g47770 (n28355, \a[26] , n_19511);
  and g47771 (n28356, n_33, n28354);
  not g47772 (n_19512, n28355);
  not g47773 (n_19513, n28356);
  and g47774 (n28357, n_19512, n_19513);
  not g47775 (n_19514, n28357);
  and g47776 (n28358, n28346, n_19514);
  not g47777 (n_19515, n28346);
  and g47778 (n28359, n_19515, n28357);
  not g47779 (n_19516, n28358);
  not g47780 (n_19517, n28359);
  and g47781 (n28360, n_19516, n_19517);
  not g47782 (n_19518, n28285);
  and g47783 (n28361, n_19518, n28360);
  not g47784 (n_19519, n28360);
  and g47785 (n28362, n28285, n_19519);
  not g47786 (n_19520, n28361);
  not g47787 (n_19521, n28362);
  and g47788 (n28363, n_19520, n_19521);
  not g47789 (n_19522, n28284);
  and g47790 (n28364, n_19522, n28363);
  not g47791 (n_19523, n28364);
  and g47792 (n28365, n_19522, n_19523);
  and g47793 (n28366, n28363, n_19523);
  not g47794 (n_19524, n28365);
  not g47795 (n_19525, n28366);
  and g47796 (n28367, n_19524, n_19525);
  and g47797 (n28368, n_19324, n_19330);
  and g47798 (n28369, n28367, n28368);
  not g47799 (n_19526, n28367);
  not g47800 (n_19527, n28368);
  and g47801 (n28370, n_19526, n_19527);
  not g47802 (n_19528, n28369);
  not g47803 (n_19529, n28370);
  and g47804 (n28371, n_19528, n_19529);
  and g47805 (n28372, n5496, n22335);
  and g47806 (n28373, n4935, n22341);
  and g47807 (n28374, n5407, n22338);
  not g47808 (n_19530, n28373);
  not g47809 (n_19531, n28374);
  and g47810 (n28375, n_19530, n_19531);
  not g47811 (n_19532, n28372);
  and g47812 (n28376, n_19532, n28375);
  and g47813 (n28377, n_1011, n28376);
  and g47814 (n28378, n24167, n28376);
  not g47815 (n_19533, n28377);
  not g47816 (n_19534, n28378);
  and g47817 (n28379, n_19533, n_19534);
  not g47818 (n_19535, n28379);
  and g47819 (n28380, \a[20] , n_19535);
  and g47820 (n28381, n_435, n28379);
  not g47821 (n_19536, n28380);
  not g47822 (n_19537, n28381);
  and g47823 (n28382, n_19536, n_19537);
  not g47824 (n_19538, n28382);
  and g47825 (n28383, n28371, n_19538);
  not g47826 (n_19539, n28371);
  and g47827 (n28384, n_19539, n28382);
  not g47828 (n_19540, n28383);
  not g47829 (n_19541, n28384);
  and g47830 (n28385, n_19540, n_19541);
  not g47831 (n_19542, n28273);
  and g47832 (n28386, n_19542, n28385);
  not g47833 (n_19543, n28385);
  and g47834 (n28387, n28273, n_19543);
  not g47835 (n_19544, n28386);
  not g47836 (n_19545, n28387);
  and g47837 (n28388, n_19544, n_19545);
  not g47838 (n_19546, n28272);
  and g47839 (n28389, n_19546, n28388);
  not g47840 (n_19547, n28389);
  and g47841 (n28390, n_19546, n_19547);
  and g47842 (n28391, n28388, n_19547);
  not g47843 (n_19548, n28390);
  not g47844 (n_19549, n28391);
  and g47845 (n28392, n_19548, n_19549);
  and g47846 (n28393, n_19350, n_19356);
  and g47847 (n28394, n28392, n28393);
  not g47848 (n_19550, n28392);
  not g47849 (n_19551, n28393);
  and g47850 (n28395, n_19550, n_19551);
  not g47851 (n_19552, n28394);
  not g47852 (n_19553, n28395);
  and g47853 (n28396, n_19552, n_19553);
  and g47854 (n28397, n7101, n22312);
  and g47855 (n28398, n6402, n22323);
  and g47856 (n28399, n6951, n22320);
  not g47857 (n_19554, n28398);
  not g47858 (n_19555, n28399);
  and g47859 (n28400, n_19554, n_19555);
  not g47860 (n_19556, n28397);
  and g47861 (n28401, n_19556, n28400);
  and g47862 (n28402, n_1885, n28401);
  and g47863 (n28403, n25315, n28401);
  not g47864 (n_19557, n28402);
  not g47865 (n_19558, n28403);
  and g47866 (n28404, n_19557, n_19558);
  not g47867 (n_19559, n28404);
  and g47868 (n28405, \a[14] , n_19559);
  and g47869 (n28406, n_652, n28404);
  not g47870 (n_19560, n28405);
  not g47871 (n_19561, n28406);
  and g47872 (n28407, n_19560, n_19561);
  not g47873 (n_19562, n28407);
  and g47874 (n28408, n28396, n_19562);
  not g47875 (n_19563, n28396);
  and g47876 (n28409, n_19563, n28407);
  not g47877 (n_19564, n28408);
  not g47878 (n_19565, n28409);
  and g47879 (n28410, n_19564, n_19565);
  not g47880 (n_19566, n28261);
  and g47881 (n28411, n_19566, n28410);
  not g47882 (n_19567, n28410);
  and g47883 (n28412, n28261, n_19567);
  not g47884 (n_19568, n28411);
  not g47885 (n_19569, n28412);
  and g47886 (n28413, n_19568, n_19569);
  not g47887 (n_19570, n28260);
  and g47888 (n28414, n_19570, n28413);
  not g47889 (n_19571, n28414);
  and g47890 (n28415, n_19570, n_19571);
  and g47891 (n28416, n28413, n_19571);
  not g47892 (n_19572, n28415);
  not g47893 (n_19573, n28416);
  and g47894 (n28417, n_19572, n_19573);
  and g47895 (n28418, n_19376, n_19382);
  and g47896 (n28419, n28417, n28418);
  not g47897 (n_19574, n28417);
  not g47898 (n_19575, n28418);
  and g47899 (n28420, n_19574, n_19575);
  not g47900 (n_19576, n28419);
  not g47901 (n_19577, n28420);
  and g47902 (n28421, n_19576, n_19577);
  and g47903 (n28422, n9331, n26890);
  and g47904 (n28423, n8418, n26066);
  and g47905 (n28424, n8860, n26060);
  not g47906 (n_19578, n28423);
  not g47907 (n_19579, n28424);
  and g47908 (n28425, n_19578, n_19579);
  not g47909 (n_19580, n28422);
  and g47910 (n28426, n_19580, n28425);
  and g47911 (n28427, n_3428, n28426);
  and g47912 (n28428, n26904, n28426);
  not g47913 (n_19581, n28427);
  not g47914 (n_19582, n28428);
  and g47915 (n28429, n_19581, n_19582);
  not g47916 (n_19583, n28429);
  and g47917 (n28430, \a[8] , n_19583);
  and g47918 (n28431, n_1106, n28429);
  not g47919 (n_19584, n28430);
  not g47920 (n_19585, n28431);
  and g47921 (n28432, n_19584, n_19585);
  not g47922 (n_19586, n28432);
  and g47923 (n28433, n28421, n_19586);
  not g47924 (n_19587, n28421);
  and g47925 (n28434, n_19587, n28432);
  not g47926 (n_19588, n28433);
  not g47927 (n_19589, n28434);
  and g47928 (n28435, n_19588, n_19589);
  not g47929 (n_19590, n28249);
  and g47930 (n28436, n_19590, n28435);
  not g47931 (n_19591, n28435);
  and g47932 (n28437, n28249, n_19591);
  not g47933 (n_19592, n28436);
  not g47934 (n_19593, n28437);
  and g47935 (n28438, n_19592, n_19593);
  not g47936 (n_19594, n28248);
  and g47937 (n28439, n_19594, n28438);
  not g47938 (n_19595, n28439);
  and g47939 (n28440, n_19594, n_19595);
  and g47940 (n28441, n28438, n_19595);
  not g47941 (n_19596, n28440);
  not g47942 (n_19597, n28441);
  and g47943 (n28442, n_19596, n_19597);
  and g47944 (n28443, n_13150, n_19417);
  and g47945 (n28444, n11055, n27964);
  not g47946 (n_19598, n28443);
  not g47947 (n_19599, n28444);
  and g47948 (n28445, n_19598, n_19599);
  not g47949 (n_19600, n28221);
  and g47950 (n28446, n11057, n_19600);
  not g47951 (n_19601, n28446);
  and g47952 (n28447, n28445, n_19601);
  not g47953 (n_19602, n28447);
  and g47954 (n28448, \a[2] , n_19602);
  not g47955 (n_19603, n28448);
  and g47956 (n28449, \a[2] , n_19603);
  and g47957 (n28450, n_19602, n_19603);
  not g47958 (n_19604, n28449);
  not g47959 (n_19605, n28450);
  and g47960 (n28451, n_19604, n_19605);
  not g47961 (n_19606, n28442);
  not g47962 (n_19607, n28451);
  and g47963 (n28452, n_19606, n_19607);
  not g47964 (n_19608, n28452);
  and g47965 (n28453, n_19606, n_19608);
  and g47966 (n28454, n_19607, n_19608);
  not g47967 (n_19609, n28453);
  not g47968 (n_19610, n28454);
  and g47969 (n28455, n_19609, n_19610);
  and g47970 (n28456, n_19402, n_19408);
  and g47971 (n28457, n28455, n28456);
  not g47972 (n_19611, n28455);
  not g47973 (n_19612, n28456);
  and g47974 (n28458, n_19611, n_19612);
  not g47975 (n_19613, n28457);
  not g47976 (n_19614, n28458);
  and g47977 (n28459, n_19613, n_19614);
  and g47978 (n28460, n_19434, n_19438);
  not g47979 (n_19615, n28459);
  and g47980 (n28461, n_19615, n28460);
  not g47981 (n_19616, n28460);
  and g47982 (n28462, n28459, n_19616);
  not g47983 (n_19617, n28461);
  not g47984 (n_19618, n28462);
  and g47985 (n28463, n_19617, n_19618);
  and g47986 (n28464, n28235, n28463);
  not g47987 (n_19619, n28463);
  and g47988 (n28465, n_19441, n_19619);
  not g47989 (n_19620, n28464);
  not g47990 (n_19621, n28465);
  and g47991 (\result[6] , n_19620, n_19621);
  and g47992 (n28467, n_19500, n_19504);
  and g47993 (n28468, n75, n23006);
  and g47994 (n28469, n3020, n22368);
  and g47995 (n28470, n3023, n22374);
  and g47996 (n28471, n3028, n22371);
  and g48022 (n28493, n_8454, n_19417);
  not g48023 (n_19626, n28493);
  and g48024 (n28494, \a[2] , n_19626);
  and g48025 (n28495, n_10, n28493);
  not g48026 (n_19627, n28494);
  not g48027 (n_19628, n28495);
  and g48028 (n28496, n_19627, n_19628);
  not g48029 (n_19629, n28492);
  not g48030 (n_19630, n28496);
  and g48031 (n28497, n_19629, n_19630);
  and g48032 (n28498, n28492, n28496);
  not g48033 (n_19631, n28474);
  not g48034 (n_19632, n28498);
  and g48035 (n28499, n_19631, n_19632);
  not g48036 (n_19633, n28497);
  and g48037 (n28500, n_19633, n28499);
  not g48038 (n_19634, n28500);
  and g48039 (n28501, n_19631, n_19634);
  and g48040 (n28502, n_19633, n_19634);
  and g48041 (n28503, n_19632, n28502);
  not g48042 (n_19635, n28501);
  not g48043 (n_19636, n28503);
  and g48044 (n28504, n_19635, n_19636);
  and g48045 (n28505, n_19482, n_19487);
  and g48046 (n28506, n28504, n28505);
  not g48047 (n_19637, n28504);
  not g48048 (n_19638, n28505);
  and g48049 (n28507, n_19637, n_19638);
  not g48050 (n_19639, n28506);
  not g48051 (n_19640, n28507);
  and g48052 (n28508, n_19639, n_19640);
  and g48053 (n28509, n3457, n22359);
  and g48054 (n28510, n3542, n22365);
  and g48055 (n28511, n3606, n22362);
  not g48056 (n_19641, n28510);
  not g48057 (n_19642, n28511);
  and g48058 (n28512, n_19641, n_19642);
  not g48059 (n_19643, n28509);
  and g48060 (n28513, n_19643, n28512);
  and g48061 (n28514, n_489, n28513);
  and g48062 (n28515, n_15331, n28513);
  not g48063 (n_19644, n28514);
  not g48064 (n_19645, n28515);
  and g48065 (n28516, n_19644, n_19645);
  not g48066 (n_19646, n28516);
  and g48067 (n28517, \a[29] , n_19646);
  and g48068 (n28518, n_15, n28516);
  not g48069 (n_19647, n28517);
  not g48070 (n_19648, n28518);
  and g48071 (n28519, n_19647, n_19648);
  not g48072 (n_19649, n28519);
  and g48073 (n28520, n28508, n_19649);
  not g48074 (n_19650, n28508);
  and g48075 (n28521, n_19650, n28519);
  not g48076 (n_19651, n28520);
  not g48077 (n_19652, n28521);
  and g48078 (n28522, n_19651, n_19652);
  not g48079 (n_19653, n28467);
  and g48080 (n28523, n_19653, n28522);
  not g48081 (n_19654, n28522);
  and g48082 (n28524, n28467, n_19654);
  not g48083 (n_19655, n28523);
  not g48084 (n_19656, n28524);
  and g48085 (n28525, n_19655, n_19656);
  and g48086 (n28526, n3884, n22350);
  and g48087 (n28527, n3967, n22356);
  and g48088 (n28528, n4046, n22353);
  and g48094 (n28531, n4050, n23672);
  not g48097 (n_19661, n28532);
  and g48098 (n28533, \a[26] , n_19661);
  not g48099 (n_19662, n28533);
  and g48100 (n28534, \a[26] , n_19662);
  and g48101 (n28535, n_19661, n_19662);
  not g48102 (n_19663, n28534);
  not g48103 (n_19664, n28535);
  and g48104 (n28536, n_19663, n_19664);
  not g48105 (n_19665, n28536);
  and g48106 (n28537, n28525, n_19665);
  not g48107 (n_19666, n28537);
  and g48108 (n28538, n28525, n_19666);
  and g48109 (n28539, n_19665, n_19666);
  not g48110 (n_19667, n28538);
  not g48111 (n_19668, n28539);
  and g48112 (n28540, n_19667, n_19668);
  and g48113 (n28541, n_19516, n_19520);
  and g48114 (n28542, n28540, n28541);
  not g48115 (n_19669, n28540);
  not g48116 (n_19670, n28541);
  and g48117 (n28543, n_19669, n_19670);
  not g48118 (n_19671, n28542);
  not g48119 (n_19672, n28543);
  and g48120 (n28544, n_19671, n_19672);
  and g48121 (n28545, n4694, n22341);
  and g48122 (n28546, n4533, n22347);
  and g48123 (n28547, n4604, n22344);
  and g48129 (n28550, n4536, n24142);
  not g48132 (n_19677, n28551);
  and g48133 (n28552, \a[23] , n_19677);
  not g48134 (n_19678, n28552);
  and g48135 (n28553, \a[23] , n_19678);
  and g48136 (n28554, n_19677, n_19678);
  not g48137 (n_19679, n28553);
  not g48138 (n_19680, n28554);
  and g48139 (n28555, n_19679, n_19680);
  not g48140 (n_19681, n28555);
  and g48141 (n28556, n28544, n_19681);
  not g48142 (n_19682, n28556);
  and g48143 (n28557, n28544, n_19682);
  and g48144 (n28558, n_19681, n_19682);
  not g48145 (n_19683, n28557);
  not g48146 (n_19684, n28558);
  and g48147 (n28559, n_19683, n_19684);
  and g48148 (n28560, n_19523, n_19529);
  and g48149 (n28561, n28559, n28560);
  not g48150 (n_19685, n28559);
  not g48151 (n_19686, n28560);
  and g48152 (n28562, n_19685, n_19686);
  not g48153 (n_19687, n28561);
  not g48154 (n_19688, n28562);
  and g48155 (n28563, n_19687, n_19688);
  and g48156 (n28564, n5496, n22332);
  and g48157 (n28565, n4935, n22338);
  and g48158 (n28566, n5407, n22335);
  and g48164 (n28569, n4938, n22542);
  not g48167 (n_19693, n28570);
  and g48168 (n28571, \a[20] , n_19693);
  not g48169 (n_19694, n28571);
  and g48170 (n28572, \a[20] , n_19694);
  and g48171 (n28573, n_19693, n_19694);
  not g48172 (n_19695, n28572);
  not g48173 (n_19696, n28573);
  and g48174 (n28574, n_19695, n_19696);
  not g48175 (n_19697, n28574);
  and g48176 (n28575, n28563, n_19697);
  not g48177 (n_19698, n28575);
  and g48178 (n28576, n28563, n_19698);
  and g48179 (n28577, n_19697, n_19698);
  not g48180 (n_19699, n28576);
  not g48181 (n_19700, n28577);
  and g48182 (n28578, n_19699, n_19700);
  and g48183 (n28579, n_19540, n_19544);
  and g48184 (n28580, n28578, n28579);
  not g48185 (n_19701, n28578);
  not g48186 (n_19702, n28579);
  and g48187 (n28581, n_19701, n_19702);
  not g48188 (n_19703, n28580);
  not g48189 (n_19704, n28581);
  and g48190 (n28582, n_19703, n_19704);
  and g48191 (n28583, n6233, n22323);
  and g48192 (n28584, n5663, n22329);
  and g48193 (n28585, n5939, n22326);
  and g48199 (n28588, n5666, n24599);
  not g48202 (n_19709, n28589);
  and g48203 (n28590, \a[17] , n_19709);
  not g48204 (n_19710, n28590);
  and g48205 (n28591, \a[17] , n_19710);
  and g48206 (n28592, n_19709, n_19710);
  not g48207 (n_19711, n28591);
  not g48208 (n_19712, n28592);
  and g48209 (n28593, n_19711, n_19712);
  not g48210 (n_19713, n28593);
  and g48211 (n28594, n28582, n_19713);
  not g48212 (n_19714, n28594);
  and g48213 (n28595, n28582, n_19714);
  and g48214 (n28596, n_19713, n_19714);
  not g48215 (n_19715, n28595);
  not g48216 (n_19716, n28596);
  and g48217 (n28597, n_19715, n_19716);
  and g48218 (n28598, n_19547, n_19553);
  and g48219 (n28599, n28597, n28598);
  not g48220 (n_19717, n28597);
  not g48221 (n_19718, n28598);
  and g48222 (n28600, n_19717, n_19718);
  not g48223 (n_19719, n28599);
  not g48224 (n_19720, n28600);
  and g48225 (n28601, n_19719, n_19720);
  and g48226 (n28602, n7101, n22315);
  and g48227 (n28603, n6402, n22320);
  and g48228 (n28604, n6951, n22312);
  and g48234 (n28607, n6397, n25294);
  not g48237 (n_19725, n28608);
  and g48238 (n28609, \a[14] , n_19725);
  not g48239 (n_19726, n28609);
  and g48240 (n28610, \a[14] , n_19726);
  and g48241 (n28611, n_19725, n_19726);
  not g48242 (n_19727, n28610);
  not g48243 (n_19728, n28611);
  and g48244 (n28612, n_19727, n_19728);
  not g48245 (n_19729, n28612);
  and g48246 (n28613, n28601, n_19729);
  not g48247 (n_19730, n28613);
  and g48248 (n28614, n28601, n_19730);
  and g48249 (n28615, n_19729, n_19730);
  not g48250 (n_19731, n28614);
  not g48251 (n_19732, n28615);
  and g48252 (n28616, n_19731, n_19732);
  and g48253 (n28617, n_19564, n_19568);
  and g48254 (n28618, n28616, n28617);
  not g48255 (n_19733, n28616);
  not g48256 (n_19734, n28617);
  and g48257 (n28619, n_19733, n_19734);
  not g48258 (n_19735, n28618);
  not g48259 (n_19736, n28619);
  and g48260 (n28620, n_19735, n_19736);
  and g48261 (n28621, n7983, n26066);
  and g48262 (n28622, n7291, n22309);
  and g48263 (n28623, n7632, n26063);
  and g48269 (n28626, n7294, n_18359);
  not g48272 (n_19741, n28627);
  and g48273 (n28628, \a[11] , n_19741);
  not g48274 (n_19742, n28628);
  and g48275 (n28629, \a[11] , n_19742);
  and g48276 (n28630, n_19741, n_19742);
  not g48277 (n_19743, n28629);
  not g48278 (n_19744, n28630);
  and g48279 (n28631, n_19743, n_19744);
  not g48280 (n_19745, n28631);
  and g48281 (n28632, n28620, n_19745);
  not g48282 (n_19746, n28632);
  and g48283 (n28633, n28620, n_19746);
  and g48284 (n28634, n_19745, n_19746);
  not g48285 (n_19747, n28633);
  not g48286 (n_19748, n28634);
  and g48287 (n28635, n_19747, n_19748);
  and g48288 (n28636, n_19571, n_19577);
  and g48289 (n28637, n28635, n28636);
  not g48290 (n_19749, n28635);
  not g48291 (n_19750, n28636);
  and g48292 (n28638, n_19749, n_19750);
  not g48293 (n_19751, n28637);
  not g48294 (n_19752, n28638);
  and g48295 (n28639, n_19751, n_19752);
  and g48296 (n28640, n9331, n27173);
  and g48297 (n28641, n8418, n26060);
  and g48298 (n28642, n8860, n26890);
  and g48304 (n28645, n8421, n27185);
  not g48307 (n_19757, n28646);
  and g48308 (n28647, \a[8] , n_19757);
  not g48309 (n_19758, n28647);
  and g48310 (n28648, \a[8] , n_19758);
  and g48311 (n28649, n_19757, n_19758);
  not g48312 (n_19759, n28648);
  not g48313 (n_19760, n28649);
  and g48314 (n28650, n_19759, n_19760);
  not g48315 (n_19761, n28650);
  and g48316 (n28651, n28639, n_19761);
  not g48317 (n_19762, n28651);
  and g48318 (n28652, n28639, n_19762);
  and g48319 (n28653, n_19761, n_19762);
  not g48320 (n_19763, n28652);
  not g48321 (n_19764, n28653);
  and g48322 (n28654, n_19763, n_19764);
  and g48323 (n28655, n_19588, n_19592);
  and g48324 (n28656, n28654, n28655);
  not g48325 (n_19765, n28654);
  not g48326 (n_19766, n28655);
  and g48327 (n28657, n_19765, n_19766);
  not g48328 (n_19767, n28656);
  not g48329 (n_19768, n28657);
  and g48330 (n28658, n_19767, n_19768);
  and g48331 (n28659, n71, n27964);
  and g48332 (n28660, n9867, n27442);
  and g48333 (n28661, n10434, n27698);
  and g48339 (n28664, n9870, n27976);
  not g48342 (n_19773, n28665);
  and g48343 (n28666, \a[5] , n_19773);
  not g48344 (n_19774, n28666);
  and g48345 (n28667, \a[5] , n_19774);
  and g48346 (n28668, n_19773, n_19774);
  not g48347 (n_19775, n28667);
  not g48348 (n_19776, n28668);
  and g48349 (n28669, n_19775, n_19776);
  not g48350 (n_19777, n28669);
  and g48351 (n28670, n28658, n_19777);
  not g48352 (n_19778, n28670);
  and g48353 (n28671, n28658, n_19778);
  and g48354 (n28672, n_19777, n_19778);
  not g48355 (n_19779, n28671);
  not g48356 (n_19780, n28672);
  and g48357 (n28673, n_19779, n_19780);
  and g48358 (n28674, n_19595, n_19608);
  and g48359 (n28675, n28673, n28674);
  not g48360 (n_19781, n28673);
  not g48361 (n_19782, n28674);
  and g48362 (n28676, n_19781, n_19782);
  not g48363 (n_19783, n28675);
  not g48364 (n_19784, n28676);
  and g48365 (n28677, n_19783, n_19784);
  and g48366 (n28678, n_19614, n_19618);
  not g48367 (n_19785, n28677);
  and g48368 (n28679, n_19785, n28678);
  not g48369 (n_19786, n28678);
  and g48370 (n28680, n28677, n_19786);
  not g48371 (n_19787, n28679);
  not g48372 (n_19788, n28680);
  and g48373 (n28681, n_19787, n_19788);
  and g48374 (n28682, n28464, n28681);
  not g48375 (n_19789, n28681);
  and g48376 (n28683, n_19620, n_19789);
  not g48377 (n_19790, n28682);
  not g48378 (n_19791, n28683);
  and g48379 (\result[7] , n_19790, n_19791);
  not g48402 (n_19792, n28706);
  and g48403 (n28707, n_19630, n_19792);
  and g48404 (n28708, n28496, n28706);
  not g48405 (n_19793, n28502);
  not g48406 (n_19794, n28708);
  and g48407 (n28709, n_19793, n_19794);
  not g48408 (n_19795, n28707);
  and g48409 (n28710, n_19795, n28709);
  not g48410 (n_19796, n28710);
  and g48411 (n28711, n_19793, n_19796);
  and g48412 (n28712, n_19795, n_19796);
  and g48413 (n28713, n_19794, n28712);
  not g48414 (n_19797, n28711);
  not g48415 (n_19798, n28713);
  and g48416 (n28714, n_19797, n_19798);
  and g48417 (n28715, n75, n_15351);
  and g48418 (n28716, n3020, n22365);
  and g48419 (n28717, n3023, n22371);
  and g48420 (n28718, n3028, n22368);
  not g48428 (n_19803, n28714);
  not g48429 (n_19804, n28721);
  and g48430 (n28722, n_19803, n_19804);
  not g48431 (n_19805, n28722);
  and g48432 (n28723, n_19803, n_19805);
  and g48433 (n28724, n_19804, n_19805);
  not g48434 (n_19806, n28723);
  not g48435 (n_19807, n28724);
  and g48436 (n28725, n_19806, n_19807);
  and g48437 (n28726, n_19640, n_19651);
  and g48438 (n28727, n28725, n28726);
  not g48439 (n_19808, n28725);
  not g48440 (n_19809, n28726);
  and g48441 (n28728, n_19808, n_19809);
  not g48442 (n_19810, n28727);
  not g48443 (n_19811, n28728);
  and g48444 (n28729, n_19810, n_19811);
  and g48445 (n28730, n3457, n22356);
  and g48446 (n28731, n3542, n22362);
  and g48447 (n28732, n3606, n22359);
  and g48453 (n28735, n3368, n_15312);
  not g48456 (n_19816, n28736);
  and g48457 (n28737, \a[29] , n_19816);
  not g48458 (n_19817, n28737);
  and g48459 (n28738, \a[29] , n_19817);
  and g48460 (n28739, n_19816, n_19817);
  not g48461 (n_19818, n28738);
  not g48462 (n_19819, n28739);
  and g48463 (n28740, n_19818, n_19819);
  not g48464 (n_19820, n28740);
  and g48465 (n28741, n28729, n_19820);
  not g48466 (n_19821, n28741);
  and g48467 (n28742, n28729, n_19821);
  and g48468 (n28743, n_19820, n_19821);
  not g48469 (n_19822, n28742);
  not g48470 (n_19823, n28743);
  and g48471 (n28744, n_19822, n_19823);
  and g48472 (n28745, n3884, n22347);
  and g48473 (n28746, n3967, n22353);
  and g48474 (n28747, n4046, n22350);
  and g48480 (n28750, n4050, n_16069);
  not g48483 (n_19828, n28751);
  and g48484 (n28752, \a[26] , n_19828);
  not g48485 (n_19829, n28752);
  and g48486 (n28753, \a[26] , n_19829);
  and g48487 (n28754, n_19828, n_19829);
  not g48488 (n_19830, n28753);
  not g48489 (n_19831, n28754);
  and g48490 (n28755, n_19830, n_19831);
  not g48491 (n_19832, n28744);
  not g48492 (n_19833, n28755);
  and g48493 (n28756, n_19832, n_19833);
  not g48494 (n_19834, n28756);
  and g48495 (n28757, n_19832, n_19834);
  and g48496 (n28758, n_19833, n_19834);
  not g48497 (n_19835, n28757);
  not g48498 (n_19836, n28758);
  and g48499 (n28759, n_19835, n_19836);
  and g48500 (n28760, n_19655, n_19666);
  and g48501 (n28761, n28759, n28760);
  not g48502 (n_19837, n28759);
  not g48503 (n_19838, n28760);
  and g48504 (n28762, n_19837, n_19838);
  not g48505 (n_19839, n28761);
  not g48506 (n_19840, n28762);
  and g48507 (n28763, n_19839, n_19840);
  and g48508 (n28764, n4694, n22338);
  and g48509 (n28765, n4533, n22344);
  and g48510 (n28766, n4604, n22341);
  and g48516 (n28769, n4536, n_16033);
  not g48519 (n_19845, n28770);
  and g48520 (n28771, \a[23] , n_19845);
  not g48521 (n_19846, n28771);
  and g48522 (n28772, \a[23] , n_19846);
  and g48523 (n28773, n_19845, n_19846);
  not g48524 (n_19847, n28772);
  not g48525 (n_19848, n28773);
  and g48526 (n28774, n_19847, n_19848);
  not g48527 (n_19849, n28774);
  and g48528 (n28775, n28763, n_19849);
  not g48529 (n_19850, n28775);
  and g48530 (n28776, n28763, n_19850);
  and g48531 (n28777, n_19849, n_19850);
  not g48532 (n_19851, n28776);
  not g48533 (n_19852, n28777);
  and g48534 (n28778, n_19851, n_19852);
  and g48535 (n28779, n_19672, n_19682);
  and g48536 (n28780, n28778, n28779);
  not g48537 (n_19853, n28778);
  not g48538 (n_19854, n28779);
  and g48539 (n28781, n_19853, n_19854);
  not g48540 (n_19855, n28780);
  not g48541 (n_19856, n28781);
  and g48542 (n28782, n_19855, n_19856);
  and g48543 (n28783, n5496, n22329);
  and g48544 (n28784, n4935, n22335);
  and g48545 (n28785, n5407, n22332);
  and g48551 (n28788, n4938, n_16827);
  not g48554 (n_19861, n28789);
  and g48555 (n28790, \a[20] , n_19861);
  not g48556 (n_19862, n28790);
  and g48557 (n28791, \a[20] , n_19862);
  and g48558 (n28792, n_19861, n_19862);
  not g48559 (n_19863, n28791);
  not g48560 (n_19864, n28792);
  and g48561 (n28793, n_19863, n_19864);
  not g48562 (n_19865, n28793);
  and g48563 (n28794, n28782, n_19865);
  not g48564 (n_19866, n28794);
  and g48565 (n28795, n28782, n_19866);
  and g48566 (n28796, n_19865, n_19866);
  not g48567 (n_19867, n28795);
  not g48568 (n_19868, n28796);
  and g48569 (n28797, n_19867, n_19868);
  and g48570 (n28798, n_19688, n_19698);
  and g48571 (n28799, n28797, n28798);
  not g48572 (n_19869, n28797);
  not g48573 (n_19870, n28798);
  and g48574 (n28800, n_19869, n_19870);
  not g48575 (n_19871, n28799);
  not g48576 (n_19872, n28800);
  and g48577 (n28801, n_19871, n_19872);
  and g48578 (n28802, n6233, n22320);
  and g48579 (n28803, n5663, n22326);
  and g48580 (n28804, n5939, n22323);
  and g48586 (n28807, n5666, n_17020);
  not g48589 (n_19877, n28808);
  and g48590 (n28809, \a[17] , n_19877);
  not g48591 (n_19878, n28809);
  and g48592 (n28810, \a[17] , n_19878);
  and g48593 (n28811, n_19877, n_19878);
  not g48594 (n_19879, n28810);
  not g48595 (n_19880, n28811);
  and g48596 (n28812, n_19879, n_19880);
  not g48597 (n_19881, n28812);
  and g48598 (n28813, n28801, n_19881);
  not g48599 (n_19882, n28813);
  and g48600 (n28814, n28801, n_19882);
  and g48601 (n28815, n_19881, n_19882);
  not g48602 (n_19883, n28814);
  not g48603 (n_19884, n28815);
  and g48604 (n28816, n_19883, n_19884);
  and g48605 (n28817, n_19704, n_19714);
  and g48606 (n28818, n28816, n28817);
  not g48607 (n_19885, n28816);
  not g48608 (n_19886, n28817);
  and g48609 (n28819, n_19885, n_19886);
  not g48610 (n_19887, n28818);
  not g48611 (n_19888, n28819);
  and g48612 (n28820, n_19887, n_19888);
  and g48613 (n28821, n7101, n22309);
  and g48614 (n28822, n6402, n22312);
  and g48615 (n28823, n6951, n22315);
  and g48621 (n28826, n6397, n_14657);
  not g48624 (n_19893, n28827);
  and g48625 (n28828, \a[14] , n_19893);
  not g48626 (n_19894, n28828);
  and g48627 (n28829, \a[14] , n_19894);
  and g48628 (n28830, n_19893, n_19894);
  not g48629 (n_19895, n28829);
  not g48630 (n_19896, n28830);
  and g48631 (n28831, n_19895, n_19896);
  not g48632 (n_19897, n28831);
  and g48633 (n28832, n28820, n_19897);
  not g48634 (n_19898, n28832);
  and g48635 (n28833, n28820, n_19898);
  and g48636 (n28834, n_19897, n_19898);
  not g48637 (n_19899, n28833);
  not g48638 (n_19900, n28834);
  and g48639 (n28835, n_19899, n_19900);
  and g48640 (n28836, n_19720, n_19730);
  and g48641 (n28837, n28835, n28836);
  not g48642 (n_19901, n28835);
  not g48643 (n_19902, n28836);
  and g48644 (n28838, n_19901, n_19902);
  not g48645 (n_19903, n28837);
  not g48646 (n_19904, n28838);
  and g48647 (n28839, n_19903, n_19904);
  and g48648 (n28840, n7983, n26060);
  and g48649 (n28841, n7291, n26063);
  and g48650 (n28842, n7632, n26066);
  and g48656 (n28845, n7294, n_18596);
  not g48659 (n_19909, n28846);
  and g48660 (n28847, \a[11] , n_19909);
  not g48661 (n_19910, n28847);
  and g48662 (n28848, \a[11] , n_19910);
  and g48663 (n28849, n_19909, n_19910);
  not g48664 (n_19911, n28848);
  not g48665 (n_19912, n28849);
  and g48666 (n28850, n_19911, n_19912);
  not g48667 (n_19913, n28850);
  and g48668 (n28851, n28839, n_19913);
  not g48669 (n_19914, n28851);
  and g48670 (n28852, n28839, n_19914);
  and g48671 (n28853, n_19913, n_19914);
  not g48672 (n_19915, n28852);
  not g48673 (n_19916, n28853);
  and g48674 (n28854, n_19915, n_19916);
  and g48675 (n28855, n_19736, n_19746);
  and g48676 (n28856, n28854, n28855);
  not g48677 (n_19917, n28854);
  not g48678 (n_19918, n28855);
  and g48679 (n28857, n_19917, n_19918);
  not g48680 (n_19919, n28856);
  not g48681 (n_19920, n28857);
  and g48682 (n28858, n_19919, n_19920);
  and g48683 (n28859, n9331, n27442);
  and g48684 (n28860, n8418, n26890);
  and g48685 (n28861, n8860, n27173);
  and g48691 (n28864, n8421, n27455);
  not g48694 (n_19925, n28865);
  and g48695 (n28866, \a[8] , n_19925);
  not g48696 (n_19926, n28866);
  and g48697 (n28867, \a[8] , n_19926);
  and g48698 (n28868, n_19925, n_19926);
  not g48699 (n_19927, n28867);
  not g48700 (n_19928, n28868);
  and g48701 (n28869, n_19927, n_19928);
  not g48702 (n_19929, n28869);
  and g48703 (n28870, n28858, n_19929);
  not g48704 (n_19930, n28870);
  and g48705 (n28871, n28858, n_19930);
  and g48706 (n28872, n_19929, n_19930);
  not g48707 (n_19931, n28871);
  not g48708 (n_19932, n28872);
  and g48709 (n28873, n_19931, n_19932);
  and g48710 (n28874, n_19752, n_19762);
  and g48711 (n28875, n28873, n28874);
  not g48712 (n_19933, n28873);
  not g48713 (n_19934, n28874);
  and g48714 (n28876, n_19933, n_19934);
  not g48715 (n_19935, n28875);
  not g48716 (n_19936, n28876);
  and g48717 (n28877, n_19935, n_19936);
  and g48718 (n28878, n71, n_19417);
  and g48719 (n28879, n9867, n27698);
  and g48720 (n28880, n10434, n27964);
  not g48726 (n_19940, n28223);
  and g48727 (n28883, n9870, n_19940);
  not g48730 (n_19942, n28884);
  and g48731 (n28885, \a[5] , n_19942);
  not g48732 (n_19943, n28885);
  and g48733 (n28886, \a[5] , n_19943);
  and g48734 (n28887, n_19942, n_19943);
  not g48735 (n_19944, n28886);
  not g48736 (n_19945, n28887);
  and g48737 (n28888, n_19944, n_19945);
  not g48738 (n_19946, n28888);
  and g48739 (n28889, n28877, n_19946);
  not g48740 (n_19947, n28889);
  and g48741 (n28890, n28877, n_19947);
  and g48742 (n28891, n_19946, n_19947);
  not g48743 (n_19948, n28890);
  not g48744 (n_19949, n28891);
  and g48745 (n28892, n_19948, n_19949);
  and g48746 (n28893, n_19768, n_19778);
  and g48747 (n28894, n28892, n28893);
  not g48748 (n_19950, n28892);
  not g48749 (n_19951, n28893);
  and g48750 (n28895, n_19950, n_19951);
  not g48751 (n_19952, n28894);
  not g48752 (n_19953, n28895);
  and g48753 (n28896, n_19952, n_19953);
  and g48754 (n28897, n_19784, n_19788);
  not g48755 (n_19954, n28896);
  and g48756 (n28898, n_19954, n28897);
  not g48757 (n_19955, n28897);
  and g48758 (n28899, n28896, n_19955);
  not g48759 (n_19956, n28898);
  not g48760 (n_19957, n28899);
  and g48761 (n28900, n_19956, n_19957);
  and g48762 (n28901, n28682, n28900);
  not g48763 (n_19958, n28900);
  and g48764 (n28902, n_19790, n_19958);
  not g48765 (n_19959, n28901);
  not g48766 (n_19960, n28902);
  and g48767 (\result[8] , n_19959, n_19960);
  not g48784 (n_19961, n28919);
  and g48785 (n28920, n_19630, n_19961);
  and g48786 (n28921, n28496, n28919);
  not g48787 (n_19962, n28712);
  not g48788 (n_19963, n28921);
  and g48789 (n28922, n_19962, n_19963);
  not g48790 (n_19964, n28920);
  and g48791 (n28923, n_19964, n28922);
  not g48792 (n_19965, n28923);
  and g48793 (n28924, n_19962, n_19965);
  and g48794 (n28925, n_19964, n_19965);
  and g48795 (n28926, n_19963, n28925);
  not g48796 (n_19966, n28924);
  not g48797 (n_19967, n28926);
  and g48798 (n28927, n_19966, n_19967);
  and g48799 (n28928, n75, n_18151);
  and g48800 (n28929, n3020, n22362);
  and g48801 (n28930, n3023, n22368);
  and g48802 (n28931, n3028, n22365);
  not g48810 (n_19972, n28927);
  not g48811 (n_19973, n28934);
  and g48812 (n28935, n_19972, n_19973);
  not g48813 (n_19974, n28935);
  and g48814 (n28936, n_19972, n_19974);
  and g48815 (n28937, n_19973, n_19974);
  not g48816 (n_19975, n28936);
  not g48817 (n_19976, n28937);
  and g48818 (n28938, n_19975, n_19976);
  and g48819 (n28939, n_19805, n_19811);
  and g48820 (n28940, n28938, n28939);
  not g48821 (n_19977, n28938);
  not g48822 (n_19978, n28939);
  and g48823 (n28941, n_19977, n_19978);
  not g48824 (n_19979, n28940);
  not g48825 (n_19980, n28941);
  and g48826 (n28942, n_19979, n_19980);
  and g48827 (n28943, n3457, n22353);
  and g48828 (n28944, n3542, n22359);
  and g48829 (n28945, n3606, n22356);
  and g48835 (n28948, n3368, n_14678);
  not g48838 (n_19985, n28949);
  and g48839 (n28950, \a[29] , n_19985);
  not g48840 (n_19986, n28950);
  and g48841 (n28951, \a[29] , n_19986);
  and g48842 (n28952, n_19985, n_19986);
  not g48843 (n_19987, n28951);
  not g48844 (n_19988, n28952);
  and g48845 (n28953, n_19987, n_19988);
  not g48846 (n_19989, n28953);
  and g48847 (n28954, n28942, n_19989);
  not g48848 (n_19990, n28954);
  and g48849 (n28955, n28942, n_19990);
  and g48850 (n28956, n_19989, n_19990);
  not g48851 (n_19991, n28955);
  not g48852 (n_19992, n28956);
  and g48853 (n28957, n_19991, n_19992);
  and g48854 (n28958, n3884, n22344);
  and g48855 (n28959, n3967, n22350);
  and g48856 (n28960, n4046, n22347);
  and g48862 (n28963, n4050, n_18142);
  not g48865 (n_19997, n28964);
  and g48866 (n28965, \a[26] , n_19997);
  not g48867 (n_19998, n28965);
  and g48868 (n28966, \a[26] , n_19998);
  and g48869 (n28967, n_19997, n_19998);
  not g48870 (n_19999, n28966);
  not g48871 (n_20000, n28967);
  and g48872 (n28968, n_19999, n_20000);
  not g48873 (n_20001, n28957);
  not g48874 (n_20002, n28968);
  and g48875 (n28969, n_20001, n_20002);
  not g48876 (n_20003, n28969);
  and g48877 (n28970, n_20001, n_20003);
  and g48878 (n28971, n_20002, n_20003);
  not g48879 (n_20004, n28970);
  not g48880 (n_20005, n28971);
  and g48881 (n28972, n_20004, n_20005);
  and g48882 (n28973, n_19821, n_19834);
  and g48883 (n28974, n28972, n28973);
  not g48884 (n_20006, n28972);
  not g48885 (n_20007, n28973);
  and g48886 (n28975, n_20006, n_20007);
  not g48887 (n_20008, n28974);
  not g48888 (n_20009, n28975);
  and g48889 (n28976, n_20008, n_20009);
  and g48890 (n28977, n4694, n22335);
  and g48891 (n28978, n4533, n22341);
  and g48892 (n28979, n4604, n22338);
  and g48898 (n28982, n4536, n_16015);
  not g48901 (n_20014, n28983);
  and g48902 (n28984, \a[23] , n_20014);
  not g48903 (n_20015, n28984);
  and g48904 (n28985, \a[23] , n_20015);
  and g48905 (n28986, n_20014, n_20015);
  not g48906 (n_20016, n28985);
  not g48907 (n_20017, n28986);
  and g48908 (n28987, n_20016, n_20017);
  not g48909 (n_20018, n28987);
  and g48910 (n28988, n28976, n_20018);
  not g48911 (n_20019, n28988);
  and g48912 (n28989, n28976, n_20019);
  and g48913 (n28990, n_20018, n_20019);
  not g48914 (n_20020, n28989);
  not g48915 (n_20021, n28990);
  and g48916 (n28991, n_20020, n_20021);
  and g48917 (n28992, n_19840, n_19850);
  and g48918 (n28993, n28991, n28992);
  not g48919 (n_20022, n28991);
  not g48920 (n_20023, n28992);
  and g48921 (n28994, n_20022, n_20023);
  not g48922 (n_20024, n28993);
  not g48923 (n_20025, n28994);
  and g48924 (n28995, n_20024, n_20025);
  and g48925 (n28996, n5496, n22326);
  and g48926 (n28997, n4935, n22332);
  and g48927 (n28998, n5407, n22329);
  and g48933 (n29001, n4938, n_18133);
  not g48936 (n_20030, n29002);
  and g48937 (n29003, \a[20] , n_20030);
  not g48938 (n_20031, n29003);
  and g48939 (n29004, \a[20] , n_20031);
  and g48940 (n29005, n_20030, n_20031);
  not g48941 (n_20032, n29004);
  not g48942 (n_20033, n29005);
  and g48943 (n29006, n_20032, n_20033);
  not g48944 (n_20034, n29006);
  and g48945 (n29007, n28995, n_20034);
  not g48946 (n_20035, n29007);
  and g48947 (n29008, n28995, n_20035);
  and g48948 (n29009, n_20034, n_20035);
  not g48949 (n_20036, n29008);
  not g48950 (n_20037, n29009);
  and g48951 (n29010, n_20036, n_20037);
  and g48952 (n29011, n_19856, n_19866);
  and g48953 (n29012, n29010, n29011);
  not g48954 (n_20038, n29010);
  not g48955 (n_20039, n29011);
  and g48956 (n29013, n_20038, n_20039);
  not g48957 (n_20040, n29012);
  not g48958 (n_20041, n29013);
  and g48959 (n29014, n_20040, n_20041);
  and g48960 (n29015, n6233, n22312);
  and g48961 (n29016, n5663, n22323);
  and g48962 (n29017, n5939, n22320);
  and g48968 (n29020, n5666, n_17004);
  not g48971 (n_20046, n29021);
  and g48972 (n29022, \a[17] , n_20046);
  not g48973 (n_20047, n29022);
  and g48974 (n29023, \a[17] , n_20047);
  and g48975 (n29024, n_20046, n_20047);
  not g48976 (n_20048, n29023);
  not g48977 (n_20049, n29024);
  and g48978 (n29025, n_20048, n_20049);
  not g48979 (n_20050, n29025);
  and g48980 (n29026, n29014, n_20050);
  not g48981 (n_20051, n29026);
  and g48982 (n29027, n29014, n_20051);
  and g48983 (n29028, n_20050, n_20051);
  not g48984 (n_20052, n29027);
  not g48985 (n_20053, n29028);
  and g48986 (n29029, n_20052, n_20053);
  and g48987 (n29030, n_19872, n_19882);
  and g48988 (n29031, n29029, n29030);
  not g48989 (n_20054, n29029);
  not g48990 (n_20055, n29030);
  and g48991 (n29032, n_20054, n_20055);
  not g48992 (n_20056, n29031);
  not g48993 (n_20057, n29032);
  and g48994 (n29033, n_20056, n_20057);
  and g48995 (n29034, n7101, n26063);
  and g48996 (n29035, n6402, n22315);
  and g48997 (n29036, n6951, n22309);
  and g49003 (n29039, n6397, n_18124);
  not g49006 (n_20062, n29040);
  and g49007 (n29041, \a[14] , n_20062);
  not g49008 (n_20063, n29041);
  and g49009 (n29042, \a[14] , n_20063);
  and g49010 (n29043, n_20062, n_20063);
  not g49011 (n_20064, n29042);
  not g49012 (n_20065, n29043);
  and g49013 (n29044, n_20064, n_20065);
  not g49014 (n_20066, n29044);
  and g49015 (n29045, n29033, n_20066);
  not g49016 (n_20067, n29045);
  and g49017 (n29046, n29033, n_20067);
  and g49018 (n29047, n_20066, n_20067);
  not g49019 (n_20068, n29046);
  not g49020 (n_20069, n29047);
  and g49021 (n29048, n_20068, n_20069);
  and g49022 (n29049, n_19888, n_19898);
  and g49023 (n29050, n29048, n29049);
  not g49024 (n_20070, n29048);
  not g49025 (n_20071, n29049);
  and g49026 (n29051, n_20070, n_20071);
  not g49027 (n_20072, n29050);
  not g49028 (n_20073, n29051);
  and g49029 (n29052, n_20072, n_20073);
  and g49030 (n29053, n7983, n26890);
  and g49031 (n29054, n7291, n26066);
  and g49032 (n29055, n7632, n26060);
  and g49038 (n29058, n7294, n_18823);
  not g49041 (n_20078, n29059);
  and g49042 (n29060, \a[11] , n_20078);
  not g49043 (n_20079, n29060);
  and g49044 (n29061, \a[11] , n_20079);
  and g49045 (n29062, n_20078, n_20079);
  not g49046 (n_20080, n29061);
  not g49047 (n_20081, n29062);
  and g49048 (n29063, n_20080, n_20081);
  not g49049 (n_20082, n29063);
  and g49050 (n29064, n29052, n_20082);
  not g49051 (n_20083, n29064);
  and g49052 (n29065, n29052, n_20083);
  and g49053 (n29066, n_20082, n_20083);
  not g49054 (n_20084, n29065);
  not g49055 (n_20085, n29066);
  and g49056 (n29067, n_20084, n_20085);
  and g49057 (n29068, n_19904, n_19914);
  and g49058 (n29069, n29067, n29068);
  not g49059 (n_20086, n29067);
  not g49060 (n_20087, n29068);
  and g49061 (n29070, n_20086, n_20087);
  not g49062 (n_20088, n29069);
  not g49063 (n_20089, n29070);
  and g49064 (n29071, n_20088, n_20089);
  and g49065 (n29072, n9331, n27698);
  and g49066 (n29073, n8418, n27173);
  and g49067 (n29074, n8860, n27442);
  and g49073 (n29077, n8421, n_19446);
  not g49076 (n_20094, n29078);
  and g49077 (n29079, \a[8] , n_20094);
  not g49078 (n_20095, n29079);
  and g49079 (n29080, \a[8] , n_20095);
  and g49080 (n29081, n_20094, n_20095);
  not g49081 (n_20096, n29080);
  not g49082 (n_20097, n29081);
  and g49083 (n29082, n_20096, n_20097);
  not g49084 (n_20098, n29082);
  and g49085 (n29083, n29071, n_20098);
  not g49086 (n_20099, n29083);
  and g49087 (n29084, n29071, n_20099);
  and g49088 (n29085, n_20098, n_20099);
  not g49089 (n_20100, n29084);
  not g49090 (n_20101, n29085);
  and g49091 (n29086, n_20100, n_20101);
  and g49092 (n29087, n_19920, n_19930);
  and g49093 (n29088, n_12001, n_19417);
  and g49094 (n29089, n9867, n27964);
  not g49095 (n_20102, n29088);
  not g49096 (n_20103, n29089);
  and g49097 (n29090, n_20102, n_20103);
  and g49098 (n29091, n_4684, n29090);
  and g49099 (n29092, n28221, n29090);
  not g49100 (n_20104, n29091);
  not g49101 (n_20105, n29092);
  and g49102 (n29093, n_20104, n_20105);
  not g49103 (n_20106, n29093);
  and g49104 (n29094, \a[5] , n_20106);
  and g49105 (n29095, n_3, n29093);
  not g49106 (n_20107, n29094);
  not g49107 (n_20108, n29095);
  and g49108 (n29096, n_20107, n_20108);
  not g49109 (n_20109, n29087);
  not g49110 (n_20110, n29096);
  and g49111 (n29097, n_20109, n_20110);
  and g49112 (n29098, n29087, n29096);
  not g49113 (n_20111, n29097);
  not g49114 (n_20112, n29098);
  and g49115 (n29099, n_20111, n_20112);
  not g49116 (n_20113, n29086);
  and g49117 (n29100, n_20113, n29099);
  not g49118 (n_20114, n29100);
  and g49119 (n29101, n_20113, n_20114);
  and g49120 (n29102, n29099, n_20114);
  not g49121 (n_20115, n29101);
  not g49122 (n_20116, n29102);
  and g49123 (n29103, n_20115, n_20116);
  and g49124 (n29104, n_19936, n_19947);
  and g49125 (n29105, n29103, n29104);
  not g49126 (n_20117, n29103);
  not g49127 (n_20118, n29104);
  and g49128 (n29106, n_20117, n_20118);
  not g49129 (n_20119, n29105);
  not g49130 (n_20120, n29106);
  and g49131 (n29107, n_20119, n_20120);
  and g49132 (n29108, n_19953, n_19957);
  not g49133 (n_20121, n29107);
  and g49134 (n29109, n_20121, n29108);
  not g49135 (n_20122, n29108);
  and g49136 (n29110, n29107, n_20122);
  not g49137 (n_20123, n29109);
  not g49138 (n_20124, n29110);
  and g49139 (n29111, n_20123, n_20124);
  and g49140 (n29112, n28901, n29111);
  not g49141 (n_20125, n29111);
  and g49142 (n29113, n_19959, n_20125);
  not g49143 (n_20126, n29112);
  not g49144 (n_20127, n29113);
  and g49145 (\result[9] , n_20126, n_20127);
  and g49146 (n29115, n_20120, n_20124);
  and g49147 (n29116, n_20111, n_20114);
  and g49148 (n29117, n_19974, n_19980);
  and g49164 (n29133, n28496, n29132);
  not g49165 (n_20128, n29132);
  and g49166 (n29134, n_19630, n_20128);
  not g49167 (n_20129, n29133);
  not g49168 (n_20130, n29134);
  and g49169 (n29135, n_20129, n_20130);
  and g49170 (n29136, n_8462, n_19417);
  and g49171 (n29137, n_3, n29136);
  not g49172 (n_20131, n29136);
  and g49173 (n29138, \a[5] , n_20131);
  not g49174 (n_20132, n29135);
  not g49175 (n_20133, n29138);
  and g49176 (n29139, n_20132, n_20133);
  not g49177 (n_20134, n29137);
  and g49178 (n29140, n_20134, n29139);
  not g49179 (n_20135, n29140);
  and g49180 (n29141, n_20132, n_20135);
  and g49181 (n29142, n_20133, n_20135);
  and g49182 (n29143, n_20134, n29142);
  not g49183 (n_20136, n29141);
  not g49184 (n_20137, n29143);
  and g49185 (n29144, n_20136, n_20137);
  not g49186 (n_20138, n28925);
  and g49187 (n29145, n_20138, n29144);
  not g49188 (n_20139, n29144);
  and g49189 (n29146, n28925, n_20139);
  not g49190 (n_20140, n29145);
  not g49191 (n_20141, n29146);
  and g49192 (n29147, n_20140, n_20141);
  and g49193 (n29148, n75, n23368);
  and g49194 (n29149, n3020, n22359);
  and g49195 (n29150, n3023, n22365);
  and g49196 (n29151, n3028, n22362);
  not g49204 (n_20146, n29147);
  not g49205 (n_20147, n29154);
  and g49206 (n29155, n_20146, n_20147);
  and g49207 (n29156, n29147, n29154);
  not g49208 (n_20148, n29155);
  not g49209 (n_20149, n29156);
  and g49210 (n29157, n_20148, n_20149);
  not g49211 (n_20150, n29157);
  and g49212 (n29158, n29117, n_20150);
  not g49213 (n_20151, n29117);
  and g49214 (n29159, n_20151, n29157);
  not g49215 (n_20152, n29158);
  not g49216 (n_20153, n29159);
  and g49217 (n29160, n_20152, n_20153);
  and g49218 (n29161, n3457, n22350);
  and g49219 (n29162, n3542, n22356);
  and g49220 (n29163, n3606, n22353);
  and g49226 (n29166, n3368, n23672);
  not g49229 (n_20158, n29167);
  and g49230 (n29168, \a[29] , n_20158);
  not g49231 (n_20159, n29168);
  and g49232 (n29169, \a[29] , n_20159);
  and g49233 (n29170, n_20158, n_20159);
  not g49234 (n_20160, n29169);
  not g49235 (n_20161, n29170);
  and g49236 (n29171, n_20160, n_20161);
  not g49237 (n_20162, n29171);
  and g49238 (n29172, n29160, n_20162);
  not g49239 (n_20163, n29172);
  and g49240 (n29173, n29160, n_20163);
  and g49241 (n29174, n_20162, n_20163);
  not g49242 (n_20164, n29173);
  not g49243 (n_20165, n29174);
  and g49244 (n29175, n_20164, n_20165);
  and g49245 (n29176, n3884, n22341);
  and g49246 (n29177, n3967, n22347);
  and g49247 (n29178, n4046, n22344);
  and g49253 (n29181, n4050, n24142);
  not g49256 (n_20170, n29182);
  and g49257 (n29183, \a[26] , n_20170);
  not g49258 (n_20171, n29183);
  and g49259 (n29184, \a[26] , n_20171);
  and g49260 (n29185, n_20170, n_20171);
  not g49261 (n_20172, n29184);
  not g49262 (n_20173, n29185);
  and g49263 (n29186, n_20172, n_20173);
  not g49264 (n_20174, n29175);
  not g49265 (n_20175, n29186);
  and g49266 (n29187, n_20174, n_20175);
  not g49267 (n_20176, n29187);
  and g49268 (n29188, n_20174, n_20176);
  and g49269 (n29189, n_20175, n_20176);
  not g49270 (n_20177, n29188);
  not g49271 (n_20178, n29189);
  and g49272 (n29190, n_20177, n_20178);
  and g49273 (n29191, n_19990, n_20003);
  and g49274 (n29192, n29190, n29191);
  not g49275 (n_20179, n29190);
  not g49276 (n_20180, n29191);
  and g49277 (n29193, n_20179, n_20180);
  not g49278 (n_20181, n29192);
  not g49279 (n_20182, n29193);
  and g49280 (n29194, n_20181, n_20182);
  and g49281 (n29195, n4694, n22332);
  and g49282 (n29196, n4533, n22338);
  and g49283 (n29197, n4604, n22335);
  and g49289 (n29200, n4536, n22542);
  not g49292 (n_20187, n29201);
  and g49293 (n29202, \a[23] , n_20187);
  not g49294 (n_20188, n29202);
  and g49295 (n29203, \a[23] , n_20188);
  and g49296 (n29204, n_20187, n_20188);
  not g49297 (n_20189, n29203);
  not g49298 (n_20190, n29204);
  and g49299 (n29205, n_20189, n_20190);
  not g49300 (n_20191, n29205);
  and g49301 (n29206, n29194, n_20191);
  not g49302 (n_20192, n29206);
  and g49303 (n29207, n29194, n_20192);
  and g49304 (n29208, n_20191, n_20192);
  not g49305 (n_20193, n29207);
  not g49306 (n_20194, n29208);
  and g49307 (n29209, n_20193, n_20194);
  and g49308 (n29210, n_20009, n_20019);
  and g49309 (n29211, n29209, n29210);
  not g49310 (n_20195, n29209);
  not g49311 (n_20196, n29210);
  and g49312 (n29212, n_20195, n_20196);
  not g49313 (n_20197, n29211);
  not g49314 (n_20198, n29212);
  and g49315 (n29213, n_20197, n_20198);
  and g49316 (n29214, n5496, n22323);
  and g49317 (n29215, n4935, n22329);
  and g49318 (n29216, n5407, n22326);
  and g49324 (n29219, n4938, n24599);
  not g49327 (n_20203, n29220);
  and g49328 (n29221, \a[20] , n_20203);
  not g49329 (n_20204, n29221);
  and g49330 (n29222, \a[20] , n_20204);
  and g49331 (n29223, n_20203, n_20204);
  not g49332 (n_20205, n29222);
  not g49333 (n_20206, n29223);
  and g49334 (n29224, n_20205, n_20206);
  not g49335 (n_20207, n29224);
  and g49336 (n29225, n29213, n_20207);
  not g49337 (n_20208, n29225);
  and g49338 (n29226, n29213, n_20208);
  and g49339 (n29227, n_20207, n_20208);
  not g49340 (n_20209, n29226);
  not g49341 (n_20210, n29227);
  and g49342 (n29228, n_20209, n_20210);
  and g49343 (n29229, n_20025, n_20035);
  and g49344 (n29230, n29228, n29229);
  not g49345 (n_20211, n29228);
  not g49346 (n_20212, n29229);
  and g49347 (n29231, n_20211, n_20212);
  not g49348 (n_20213, n29230);
  not g49349 (n_20214, n29231);
  and g49350 (n29232, n_20213, n_20214);
  and g49351 (n29233, n6233, n22315);
  and g49352 (n29234, n5663, n22320);
  and g49353 (n29235, n5939, n22312);
  and g49359 (n29238, n5666, n25294);
  not g49362 (n_20219, n29239);
  and g49363 (n29240, \a[17] , n_20219);
  not g49364 (n_20220, n29240);
  and g49365 (n29241, \a[17] , n_20220);
  and g49366 (n29242, n_20219, n_20220);
  not g49367 (n_20221, n29241);
  not g49368 (n_20222, n29242);
  and g49369 (n29243, n_20221, n_20222);
  not g49370 (n_20223, n29243);
  and g49371 (n29244, n29232, n_20223);
  not g49372 (n_20224, n29244);
  and g49373 (n29245, n29232, n_20224);
  and g49374 (n29246, n_20223, n_20224);
  not g49375 (n_20225, n29245);
  not g49376 (n_20226, n29246);
  and g49377 (n29247, n_20225, n_20226);
  and g49378 (n29248, n_20041, n_20051);
  and g49379 (n29249, n29247, n29248);
  not g49380 (n_20227, n29247);
  not g49381 (n_20228, n29248);
  and g49382 (n29250, n_20227, n_20228);
  not g49383 (n_20229, n29249);
  not g49384 (n_20230, n29250);
  and g49385 (n29251, n_20229, n_20230);
  and g49386 (n29252, n_20057, n_20067);
  and g49387 (n29253, n7101, n26066);
  and g49388 (n29254, n6402, n22309);
  and g49389 (n29255, n6951, n26063);
  and g49395 (n29258, n6397, n_18359);
  not g49398 (n_20235, n29259);
  and g49399 (n29260, \a[14] , n_20235);
  not g49400 (n_20236, n29260);
  and g49401 (n29261, \a[14] , n_20236);
  and g49402 (n29262, n_20235, n_20236);
  not g49403 (n_20237, n29261);
  not g49404 (n_20238, n29262);
  and g49405 (n29263, n_20237, n_20238);
  not g49406 (n_20239, n29252);
  not g49407 (n_20240, n29263);
  and g49408 (n29264, n_20239, n_20240);
  not g49409 (n_20241, n29264);
  and g49410 (n29265, n_20239, n_20241);
  and g49411 (n29266, n_20240, n_20241);
  not g49412 (n_20242, n29265);
  not g49413 (n_20243, n29266);
  and g49414 (n29267, n_20242, n_20243);
  not g49415 (n_20244, n29251);
  and g49416 (n29268, n_20244, n29267);
  not g49417 (n_20245, n29267);
  and g49418 (n29269, n29251, n_20245);
  not g49419 (n_20246, n29268);
  not g49420 (n_20247, n29269);
  and g49421 (n29270, n_20246, n_20247);
  and g49422 (n29271, n7983, n27173);
  and g49423 (n29272, n7291, n26060);
  and g49424 (n29273, n7632, n26890);
  and g49430 (n29276, n7294, n27185);
  not g49433 (n_20252, n29277);
  and g49434 (n29278, \a[11] , n_20252);
  not g49435 (n_20253, n29278);
  and g49436 (n29279, \a[11] , n_20253);
  and g49437 (n29280, n_20252, n_20253);
  not g49438 (n_20254, n29279);
  not g49439 (n_20255, n29280);
  and g49440 (n29281, n_20254, n_20255);
  not g49441 (n_20256, n29281);
  and g49442 (n29282, n29270, n_20256);
  not g49443 (n_20257, n29282);
  and g49444 (n29283, n29270, n_20257);
  and g49445 (n29284, n_20256, n_20257);
  not g49446 (n_20258, n29283);
  not g49447 (n_20259, n29284);
  and g49448 (n29285, n_20258, n_20259);
  and g49449 (n29286, n_20073, n_20083);
  and g49450 (n29287, n29285, n29286);
  not g49451 (n_20260, n29285);
  not g49452 (n_20261, n29286);
  and g49453 (n29288, n_20260, n_20261);
  not g49454 (n_20262, n29287);
  not g49455 (n_20263, n29288);
  and g49456 (n29289, n_20262, n_20263);
  and g49457 (n29290, n_20089, n_20099);
  and g49458 (n29291, n9331, n27964);
  and g49459 (n29292, n8418, n27442);
  and g49460 (n29293, n8860, n27698);
  and g49466 (n29296, n8421, n27976);
  not g49469 (n_20268, n29297);
  and g49470 (n29298, \a[8] , n_20268);
  not g49471 (n_20269, n29298);
  and g49472 (n29299, \a[8] , n_20269);
  and g49473 (n29300, n_20268, n_20269);
  not g49474 (n_20270, n29299);
  not g49475 (n_20271, n29300);
  and g49476 (n29301, n_20270, n_20271);
  not g49477 (n_20272, n29290);
  not g49478 (n_20273, n29301);
  and g49479 (n29302, n_20272, n_20273);
  not g49480 (n_20274, n29302);
  and g49481 (n29303, n_20272, n_20274);
  and g49482 (n29304, n_20273, n_20274);
  not g49483 (n_20275, n29303);
  not g49484 (n_20276, n29304);
  and g49485 (n29305, n_20275, n_20276);
  not g49486 (n_20277, n29289);
  and g49487 (n29306, n_20277, n29305);
  not g49488 (n_20278, n29305);
  and g49489 (n29307, n29289, n_20278);
  not g49490 (n_20279, n29306);
  not g49491 (n_20280, n29307);
  and g49492 (n29308, n_20279, n_20280);
  not g49493 (n_20281, n29116);
  and g49494 (n29309, n_20281, n29308);
  not g49495 (n_20282, n29308);
  and g49496 (n29310, n29116, n_20282);
  not g49497 (n_20283, n29309);
  not g49498 (n_20284, n29310);
  and g49499 (n29311, n_20283, n_20284);
  not g49500 (n_20285, n29115);
  and g49501 (n29312, n_20285, n29311);
  not g49502 (n_20286, n29311);
  and g49503 (n29313, n29115, n_20286);
  not g49504 (n_20287, n29312);
  not g49505 (n_20288, n29313);
  and g49506 (n29314, n_20287, n_20288);
  not g49507 (n_20289, n29314);
  and g49508 (n29315, n_20126, n_20289);
  and g49509 (n29316, n29112, n29314);
  not g49510 (n_20290, n29315);
  not g49511 (n_20291, n29316);
  and g49512 (\result[10] , n_20290, n_20291);
  and g49513 (n29318, n_20153, n_20163);
  and g49514 (n29319, n75, n_15312);
  and g49515 (n29320, n3020, n22356);
  and g49516 (n29321, n3023, n22362);
  and g49517 (n29322, n3028, n22359);
  and g49555 (n29356, n28496, n_20128);
  not g49556 (n_20296, n29356);
  and g49557 (n29357, n_20135, n_20296);
  not g49558 (n_20297, n29357);
  and g49559 (n29358, n29355, n_20297);
  not g49560 (n_20298, n29355);
  and g49561 (n29359, n_20298, n29357);
  not g49562 (n_20299, n29358);
  not g49563 (n_20300, n29359);
  and g49564 (n29360, n_20299, n_20300);
  not g49565 (n_20301, n29325);
  and g49566 (n29361, n_20301, n29360);
  not g49567 (n_20302, n29361);
  and g49568 (n29362, n_20301, n_20302);
  and g49569 (n29363, n29360, n_20302);
  not g49570 (n_20303, n29362);
  not g49571 (n_20304, n29363);
  and g49572 (n29364, n_20303, n_20304);
  and g49573 (n29365, n_20138, n_20139);
  not g49574 (n_20305, n29365);
  and g49575 (n29366, n_20148, n_20305);
  and g49576 (n29367, n29364, n29366);
  not g49577 (n_20306, n29364);
  not g49578 (n_20307, n29366);
  and g49579 (n29368, n_20306, n_20307);
  not g49580 (n_20308, n29367);
  not g49581 (n_20309, n29368);
  and g49582 (n29369, n_20308, n_20309);
  and g49583 (n29370, n3457, n22347);
  and g49584 (n29371, n3542, n22353);
  and g49585 (n29372, n3606, n22350);
  not g49586 (n_20310, n29371);
  not g49587 (n_20311, n29372);
  and g49588 (n29373, n_20310, n_20311);
  not g49589 (n_20312, n29370);
  and g49590 (n29374, n_20312, n29373);
  and g49591 (n29375, n_489, n29374);
  and g49592 (n29376, n23659, n29374);
  not g49593 (n_20313, n29375);
  not g49594 (n_20314, n29376);
  and g49595 (n29377, n_20313, n_20314);
  not g49596 (n_20315, n29377);
  and g49597 (n29378, \a[29] , n_20315);
  and g49598 (n29379, n_15, n29377);
  not g49599 (n_20316, n29378);
  not g49600 (n_20317, n29379);
  and g49601 (n29380, n_20316, n_20317);
  not g49602 (n_20318, n29380);
  and g49603 (n29381, n29369, n_20318);
  not g49604 (n_20319, n29369);
  and g49605 (n29382, n_20319, n29380);
  not g49606 (n_20320, n29381);
  not g49607 (n_20321, n29382);
  and g49608 (n29383, n_20320, n_20321);
  not g49609 (n_20322, n29318);
  and g49610 (n29384, n_20322, n29383);
  not g49611 (n_20323, n29383);
  and g49612 (n29385, n29318, n_20323);
  not g49613 (n_20324, n29384);
  not g49614 (n_20325, n29385);
  and g49615 (n29386, n_20324, n_20325);
  and g49616 (n29387, n3884, n22338);
  and g49617 (n29388, n3967, n22344);
  and g49618 (n29389, n4046, n22341);
  and g49624 (n29392, n4050, n_16033);
  not g49627 (n_20330, n29393);
  and g49628 (n29394, \a[26] , n_20330);
  not g49629 (n_20331, n29394);
  and g49630 (n29395, \a[26] , n_20331);
  and g49631 (n29396, n_20330, n_20331);
  not g49632 (n_20332, n29395);
  not g49633 (n_20333, n29396);
  and g49634 (n29397, n_20332, n_20333);
  not g49635 (n_20334, n29397);
  and g49636 (n29398, n29386, n_20334);
  not g49637 (n_20335, n29398);
  and g49638 (n29399, n29386, n_20335);
  and g49639 (n29400, n_20334, n_20335);
  not g49640 (n_20336, n29399);
  not g49641 (n_20337, n29400);
  and g49642 (n29401, n_20336, n_20337);
  and g49643 (n29402, n_20176, n_20182);
  and g49644 (n29403, n29401, n29402);
  not g49645 (n_20338, n29401);
  not g49646 (n_20339, n29402);
  and g49647 (n29404, n_20338, n_20339);
  not g49648 (n_20340, n29403);
  not g49649 (n_20341, n29404);
  and g49650 (n29405, n_20340, n_20341);
  and g49651 (n29406, n4694, n22329);
  and g49652 (n29407, n4533, n22335);
  and g49653 (n29408, n4604, n22332);
  and g49659 (n29411, n4536, n_16827);
  not g49662 (n_20346, n29412);
  and g49663 (n29413, \a[23] , n_20346);
  not g49664 (n_20347, n29413);
  and g49665 (n29414, \a[23] , n_20347);
  and g49666 (n29415, n_20346, n_20347);
  not g49667 (n_20348, n29414);
  not g49668 (n_20349, n29415);
  and g49669 (n29416, n_20348, n_20349);
  not g49670 (n_20350, n29416);
  and g49671 (n29417, n29405, n_20350);
  not g49672 (n_20351, n29417);
  and g49673 (n29418, n29405, n_20351);
  and g49674 (n29419, n_20350, n_20351);
  not g49675 (n_20352, n29418);
  not g49676 (n_20353, n29419);
  and g49677 (n29420, n_20352, n_20353);
  and g49678 (n29421, n_20192, n_20198);
  and g49679 (n29422, n29420, n29421);
  not g49680 (n_20354, n29420);
  not g49681 (n_20355, n29421);
  and g49682 (n29423, n_20354, n_20355);
  not g49683 (n_20356, n29422);
  not g49684 (n_20357, n29423);
  and g49685 (n29424, n_20356, n_20357);
  and g49686 (n29425, n5496, n22320);
  and g49687 (n29426, n4935, n22326);
  and g49688 (n29427, n5407, n22323);
  and g49694 (n29430, n4938, n_17020);
  not g49697 (n_20362, n29431);
  and g49698 (n29432, \a[20] , n_20362);
  not g49699 (n_20363, n29432);
  and g49700 (n29433, \a[20] , n_20363);
  and g49701 (n29434, n_20362, n_20363);
  not g49702 (n_20364, n29433);
  not g49703 (n_20365, n29434);
  and g49704 (n29435, n_20364, n_20365);
  not g49705 (n_20366, n29435);
  and g49706 (n29436, n29424, n_20366);
  not g49707 (n_20367, n29436);
  and g49708 (n29437, n29424, n_20367);
  and g49709 (n29438, n_20366, n_20367);
  not g49710 (n_20368, n29437);
  not g49711 (n_20369, n29438);
  and g49712 (n29439, n_20368, n_20369);
  and g49713 (n29440, n_20208, n_20214);
  and g49714 (n29441, n29439, n29440);
  not g49715 (n_20370, n29439);
  not g49716 (n_20371, n29440);
  and g49717 (n29442, n_20370, n_20371);
  not g49718 (n_20372, n29441);
  not g49719 (n_20373, n29442);
  and g49720 (n29443, n_20372, n_20373);
  and g49721 (n29444, n6233, n22309);
  and g49722 (n29445, n5663, n22312);
  and g49723 (n29446, n5939, n22315);
  and g49729 (n29449, n5666, n_14657);
  not g49732 (n_20378, n29450);
  and g49733 (n29451, \a[17] , n_20378);
  not g49734 (n_20379, n29451);
  and g49735 (n29452, \a[17] , n_20379);
  and g49736 (n29453, n_20378, n_20379);
  not g49737 (n_20380, n29452);
  not g49738 (n_20381, n29453);
  and g49739 (n29454, n_20380, n_20381);
  not g49740 (n_20382, n29454);
  and g49741 (n29455, n29443, n_20382);
  not g49742 (n_20383, n29455);
  and g49743 (n29456, n29443, n_20383);
  and g49744 (n29457, n_20382, n_20383);
  not g49745 (n_20384, n29456);
  not g49746 (n_20385, n29457);
  and g49747 (n29458, n_20384, n_20385);
  and g49748 (n29459, n_20224, n_20230);
  and g49749 (n29460, n29458, n29459);
  not g49750 (n_20386, n29458);
  not g49751 (n_20387, n29459);
  and g49752 (n29461, n_20386, n_20387);
  not g49753 (n_20388, n29460);
  not g49754 (n_20389, n29461);
  and g49755 (n29462, n_20388, n_20389);
  and g49756 (n29463, n7101, n26060);
  and g49757 (n29464, n6402, n26063);
  and g49758 (n29465, n6951, n26066);
  and g49764 (n29468, n6397, n_18596);
  not g49767 (n_20394, n29469);
  and g49768 (n29470, \a[14] , n_20394);
  not g49769 (n_20395, n29470);
  and g49770 (n29471, \a[14] , n_20395);
  and g49771 (n29472, n_20394, n_20395);
  not g49772 (n_20396, n29471);
  not g49773 (n_20397, n29472);
  and g49774 (n29473, n_20396, n_20397);
  not g49775 (n_20398, n29473);
  and g49776 (n29474, n29462, n_20398);
  not g49777 (n_20399, n29474);
  and g49778 (n29475, n29462, n_20399);
  and g49779 (n29476, n_20398, n_20399);
  not g49780 (n_20400, n29475);
  not g49781 (n_20401, n29476);
  and g49782 (n29477, n_20400, n_20401);
  and g49783 (n29478, n_20241, n_20247);
  not g49784 (n_20402, n29477);
  not g49785 (n_20403, n29478);
  and g49786 (n29479, n_20402, n_20403);
  not g49787 (n_20404, n29479);
  and g49788 (n29480, n_20402, n_20404);
  and g49789 (n29481, n_20403, n_20404);
  not g49790 (n_20405, n29480);
  not g49791 (n_20406, n29481);
  and g49792 (n29482, n_20405, n_20406);
  and g49793 (n29483, n7983, n27442);
  and g49794 (n29484, n7291, n26890);
  and g49795 (n29485, n7632, n27173);
  and g49801 (n29488, n7294, n27455);
  not g49804 (n_20411, n29489);
  and g49805 (n29490, \a[11] , n_20411);
  not g49806 (n_20412, n29490);
  and g49807 (n29491, \a[11] , n_20412);
  and g49808 (n29492, n_20411, n_20412);
  not g49809 (n_20413, n29491);
  not g49810 (n_20414, n29492);
  and g49811 (n29493, n_20413, n_20414);
  not g49812 (n_20415, n29482);
  not g49813 (n_20416, n29493);
  and g49814 (n29494, n_20415, n_20416);
  not g49815 (n_20417, n29494);
  and g49816 (n29495, n_20415, n_20417);
  and g49817 (n29496, n_20416, n_20417);
  not g49818 (n_20418, n29495);
  not g49819 (n_20419, n29496);
  and g49820 (n29497, n_20418, n_20419);
  and g49821 (n29498, n_20257, n_20263);
  and g49822 (n29499, n29497, n29498);
  not g49823 (n_20420, n29497);
  not g49824 (n_20421, n29498);
  and g49825 (n29500, n_20420, n_20421);
  not g49826 (n_20422, n29499);
  not g49827 (n_20423, n29500);
  and g49828 (n29501, n_20422, n_20423);
  and g49829 (n29502, n9331, n_19417);
  and g49830 (n29503, n8418, n27698);
  and g49831 (n29504, n8860, n27964);
  and g49837 (n29507, n8421, n_19940);
  not g49840 (n_20428, n29508);
  and g49841 (n29509, \a[8] , n_20428);
  not g49842 (n_20429, n29509);
  and g49843 (n29510, \a[8] , n_20429);
  and g49844 (n29511, n_20428, n_20429);
  not g49845 (n_20430, n29510);
  not g49846 (n_20431, n29511);
  and g49847 (n29512, n_20430, n_20431);
  not g49848 (n_20432, n29512);
  and g49849 (n29513, n29501, n_20432);
  not g49850 (n_20433, n29513);
  and g49851 (n29514, n29501, n_20433);
  and g49852 (n29515, n_20432, n_20433);
  not g49853 (n_20434, n29514);
  not g49854 (n_20435, n29515);
  and g49855 (n29516, n_20434, n_20435);
  and g49856 (n29517, n_20274, n_20280);
  not g49857 (n_20436, n29516);
  not g49858 (n_20437, n29517);
  and g49859 (n29518, n_20436, n_20437);
  not g49860 (n_20438, n29518);
  and g49861 (n29519, n_20436, n_20438);
  and g49862 (n29520, n_20437, n_20438);
  not g49863 (n_20439, n29519);
  not g49864 (n_20440, n29520);
  and g49865 (n29521, n_20439, n_20440);
  and g49866 (n29522, n_20283, n_20287);
  and g49867 (n29523, n29521, n29522);
  not g49868 (n_20441, n29521);
  not g49869 (n_20442, n29522);
  and g49870 (n29524, n_20441, n_20442);
  not g49871 (n_20443, n29523);
  not g49872 (n_20444, n29524);
  and g49873 (n29525, n_20443, n_20444);
  and g49874 (n29526, n_20291, n29525);
  not g49875 (n_20445, n29525);
  and g49876 (n29527, n29316, n_20445);
  or g49877 (\result[11] , n29526, n29527);
  and g49878 (n29529, n29316, n29525);
  and g49879 (n29530, n_20299, n_20302);
  and g49914 (n29565, n_20298, n29564);
  not g49915 (n_20446, n29564);
  and g49916 (n29566, n29355, n_20446);
  not g49917 (n_20447, n29530);
  not g49918 (n_20448, n29566);
  and g49919 (n29567, n_20447, n_20448);
  not g49920 (n_20449, n29565);
  and g49921 (n29568, n_20449, n29567);
  not g49922 (n_20450, n29568);
  and g49923 (n29569, n_20447, n_20450);
  and g49924 (n29570, n_20448, n_20450);
  and g49925 (n29571, n_20449, n29570);
  not g49926 (n_20451, n29569);
  not g49927 (n_20452, n29571);
  and g49928 (n29572, n_20451, n_20452);
  and g49929 (n29573, n75, n_14678);
  and g49930 (n29574, n3020, n22353);
  and g49931 (n29575, n3023, n22359);
  and g49932 (n29576, n3028, n22356);
  not g49940 (n_20457, n29572);
  not g49941 (n_20458, n29579);
  and g49942 (n29580, n_20457, n_20458);
  not g49943 (n_20459, n29580);
  and g49944 (n29581, n_20457, n_20459);
  and g49945 (n29582, n_20458, n_20459);
  not g49946 (n_20460, n29581);
  not g49947 (n_20461, n29582);
  and g49948 (n29583, n_20460, n_20461);
  and g49949 (n29584, n_20309, n_20320);
  and g49950 (n29585, n29583, n29584);
  not g49951 (n_20462, n29583);
  not g49952 (n_20463, n29584);
  and g49953 (n29586, n_20462, n_20463);
  not g49954 (n_20464, n29585);
  not g49955 (n_20465, n29586);
  and g49956 (n29587, n_20464, n_20465);
  and g49957 (n29588, n3457, n22344);
  and g49958 (n29589, n3542, n22350);
  and g49959 (n29590, n3606, n22347);
  and g49965 (n29593, n3368, n_18142);
  not g49968 (n_20470, n29594);
  and g49969 (n29595, \a[29] , n_20470);
  not g49970 (n_20471, n29595);
  and g49971 (n29596, \a[29] , n_20471);
  and g49972 (n29597, n_20470, n_20471);
  not g49973 (n_20472, n29596);
  not g49974 (n_20473, n29597);
  and g49975 (n29598, n_20472, n_20473);
  not g49976 (n_20474, n29598);
  and g49977 (n29599, n29587, n_20474);
  not g49978 (n_20475, n29599);
  and g49979 (n29600, n29587, n_20475);
  and g49980 (n29601, n_20474, n_20475);
  not g49981 (n_20476, n29600);
  not g49982 (n_20477, n29601);
  and g49983 (n29602, n_20476, n_20477);
  and g49984 (n29603, n3884, n22335);
  and g49985 (n29604, n3967, n22341);
  and g49986 (n29605, n4046, n22338);
  and g49992 (n29608, n4050, n_16015);
  not g49995 (n_20482, n29609);
  and g49996 (n29610, \a[26] , n_20482);
  not g49997 (n_20483, n29610);
  and g49998 (n29611, \a[26] , n_20483);
  and g49999 (n29612, n_20482, n_20483);
  not g50000 (n_20484, n29611);
  not g50001 (n_20485, n29612);
  and g50002 (n29613, n_20484, n_20485);
  not g50003 (n_20486, n29602);
  not g50004 (n_20487, n29613);
  and g50005 (n29614, n_20486, n_20487);
  not g50006 (n_20488, n29614);
  and g50007 (n29615, n_20486, n_20488);
  and g50008 (n29616, n_20487, n_20488);
  not g50009 (n_20489, n29615);
  not g50010 (n_20490, n29616);
  and g50011 (n29617, n_20489, n_20490);
  and g50012 (n29618, n_20324, n_20335);
  and g50013 (n29619, n29617, n29618);
  not g50014 (n_20491, n29617);
  not g50015 (n_20492, n29618);
  and g50016 (n29620, n_20491, n_20492);
  not g50017 (n_20493, n29619);
  not g50018 (n_20494, n29620);
  and g50019 (n29621, n_20493, n_20494);
  and g50020 (n29622, n4694, n22326);
  and g50021 (n29623, n4533, n22332);
  and g50022 (n29624, n4604, n22329);
  and g50028 (n29627, n4536, n_18133);
  not g50031 (n_20499, n29628);
  and g50032 (n29629, \a[23] , n_20499);
  not g50033 (n_20500, n29629);
  and g50034 (n29630, \a[23] , n_20500);
  and g50035 (n29631, n_20499, n_20500);
  not g50036 (n_20501, n29630);
  not g50037 (n_20502, n29631);
  and g50038 (n29632, n_20501, n_20502);
  not g50039 (n_20503, n29632);
  and g50040 (n29633, n29621, n_20503);
  not g50041 (n_20504, n29633);
  and g50042 (n29634, n29621, n_20504);
  and g50043 (n29635, n_20503, n_20504);
  not g50044 (n_20505, n29634);
  not g50045 (n_20506, n29635);
  and g50046 (n29636, n_20505, n_20506);
  and g50047 (n29637, n_20341, n_20351);
  and g50048 (n29638, n29636, n29637);
  not g50049 (n_20507, n29636);
  not g50050 (n_20508, n29637);
  and g50051 (n29639, n_20507, n_20508);
  not g50052 (n_20509, n29638);
  not g50053 (n_20510, n29639);
  and g50054 (n29640, n_20509, n_20510);
  and g50055 (n29641, n5496, n22312);
  and g50056 (n29642, n4935, n22323);
  and g50057 (n29643, n5407, n22320);
  and g50063 (n29646, n4938, n_17004);
  not g50066 (n_20515, n29647);
  and g50067 (n29648, \a[20] , n_20515);
  not g50068 (n_20516, n29648);
  and g50069 (n29649, \a[20] , n_20516);
  and g50070 (n29650, n_20515, n_20516);
  not g50071 (n_20517, n29649);
  not g50072 (n_20518, n29650);
  and g50073 (n29651, n_20517, n_20518);
  not g50074 (n_20519, n29651);
  and g50075 (n29652, n29640, n_20519);
  not g50076 (n_20520, n29652);
  and g50077 (n29653, n29640, n_20520);
  and g50078 (n29654, n_20519, n_20520);
  not g50079 (n_20521, n29653);
  not g50080 (n_20522, n29654);
  and g50081 (n29655, n_20521, n_20522);
  and g50082 (n29656, n_20357, n_20367);
  and g50083 (n29657, n29655, n29656);
  not g50084 (n_20523, n29655);
  not g50085 (n_20524, n29656);
  and g50086 (n29658, n_20523, n_20524);
  not g50087 (n_20525, n29657);
  not g50088 (n_20526, n29658);
  and g50089 (n29659, n_20525, n_20526);
  and g50090 (n29660, n6233, n26063);
  and g50091 (n29661, n5663, n22315);
  and g50092 (n29662, n5939, n22309);
  and g50098 (n29665, n5666, n_18124);
  not g50101 (n_20531, n29666);
  and g50102 (n29667, \a[17] , n_20531);
  not g50103 (n_20532, n29667);
  and g50104 (n29668, \a[17] , n_20532);
  and g50105 (n29669, n_20531, n_20532);
  not g50106 (n_20533, n29668);
  not g50107 (n_20534, n29669);
  and g50108 (n29670, n_20533, n_20534);
  not g50109 (n_20535, n29670);
  and g50110 (n29671, n29659, n_20535);
  not g50111 (n_20536, n29671);
  and g50112 (n29672, n29659, n_20536);
  and g50113 (n29673, n_20535, n_20536);
  not g50114 (n_20537, n29672);
  not g50115 (n_20538, n29673);
  and g50116 (n29674, n_20537, n_20538);
  and g50117 (n29675, n_20373, n_20383);
  and g50118 (n29676, n29674, n29675);
  not g50119 (n_20539, n29674);
  not g50120 (n_20540, n29675);
  and g50121 (n29677, n_20539, n_20540);
  not g50122 (n_20541, n29676);
  not g50123 (n_20542, n29677);
  and g50124 (n29678, n_20541, n_20542);
  and g50125 (n29679, n7101, n26890);
  and g50126 (n29680, n6402, n26066);
  and g50127 (n29681, n6951, n26060);
  and g50133 (n29684, n6397, n_18823);
  not g50136 (n_20547, n29685);
  and g50137 (n29686, \a[14] , n_20547);
  not g50138 (n_20548, n29686);
  and g50139 (n29687, \a[14] , n_20548);
  and g50140 (n29688, n_20547, n_20548);
  not g50141 (n_20549, n29687);
  not g50142 (n_20550, n29688);
  and g50143 (n29689, n_20549, n_20550);
  not g50144 (n_20551, n29689);
  and g50145 (n29690, n29678, n_20551);
  not g50146 (n_20552, n29690);
  and g50147 (n29691, n29678, n_20552);
  and g50148 (n29692, n_20551, n_20552);
  not g50149 (n_20553, n29691);
  not g50150 (n_20554, n29692);
  and g50151 (n29693, n_20553, n_20554);
  and g50152 (n29694, n_20389, n_20399);
  and g50153 (n29695, n29693, n29694);
  not g50154 (n_20555, n29693);
  not g50155 (n_20556, n29694);
  and g50156 (n29696, n_20555, n_20556);
  not g50157 (n_20557, n29695);
  not g50158 (n_20558, n29696);
  and g50159 (n29697, n_20557, n_20558);
  and g50160 (n29698, n7983, n27698);
  and g50161 (n29699, n7291, n27173);
  and g50162 (n29700, n7632, n27442);
  and g50168 (n29703, n7294, n_19446);
  not g50171 (n_20563, n29704);
  and g50172 (n29705, \a[11] , n_20563);
  not g50173 (n_20564, n29705);
  and g50174 (n29706, \a[11] , n_20564);
  and g50175 (n29707, n_20563, n_20564);
  not g50176 (n_20565, n29706);
  not g50177 (n_20566, n29707);
  and g50178 (n29708, n_20565, n_20566);
  not g50179 (n_20567, n29708);
  and g50180 (n29709, n29697, n_20567);
  not g50181 (n_20568, n29709);
  and g50182 (n29710, n29697, n_20568);
  and g50183 (n29711, n_20567, n_20568);
  not g50184 (n_20569, n29710);
  not g50185 (n_20570, n29711);
  and g50186 (n29712, n_20569, n_20570);
  and g50187 (n29713, n_20404, n_20417);
  and g50188 (n29714, n_10598, n_19417);
  and g50189 (n29715, n8418, n27964);
  not g50190 (n_20571, n29714);
  not g50191 (n_20572, n29715);
  and g50192 (n29716, n_20571, n_20572);
  and g50193 (n29717, n_3428, n29716);
  and g50194 (n29718, n28221, n29716);
  not g50195 (n_20573, n29717);
  not g50196 (n_20574, n29718);
  and g50197 (n29719, n_20573, n_20574);
  not g50198 (n_20575, n29719);
  and g50199 (n29720, \a[8] , n_20575);
  and g50200 (n29721, n_1106, n29719);
  not g50201 (n_20576, n29720);
  not g50202 (n_20577, n29721);
  and g50203 (n29722, n_20576, n_20577);
  not g50204 (n_20578, n29713);
  not g50205 (n_20579, n29722);
  and g50206 (n29723, n_20578, n_20579);
  and g50207 (n29724, n29713, n29722);
  not g50208 (n_20580, n29723);
  not g50209 (n_20581, n29724);
  and g50210 (n29725, n_20580, n_20581);
  not g50211 (n_20582, n29712);
  and g50212 (n29726, n_20582, n29725);
  not g50213 (n_20583, n29726);
  and g50214 (n29727, n_20582, n_20583);
  and g50215 (n29728, n29725, n_20583);
  not g50216 (n_20584, n29727);
  not g50217 (n_20585, n29728);
  and g50218 (n29729, n_20584, n_20585);
  and g50219 (n29730, n_20423, n_20433);
  and g50220 (n29731, n29729, n29730);
  not g50221 (n_20586, n29729);
  not g50222 (n_20587, n29730);
  and g50223 (n29732, n_20586, n_20587);
  not g50224 (n_20588, n29731);
  not g50225 (n_20589, n29732);
  and g50226 (n29733, n_20588, n_20589);
  and g50227 (n29734, n_20438, n_20444);
  not g50228 (n_20590, n29733);
  and g50229 (n29735, n_20590, n29734);
  not g50230 (n_20591, n29734);
  and g50231 (n29736, n29733, n_20591);
  not g50232 (n_20592, n29735);
  not g50233 (n_20593, n29736);
  and g50234 (n29737, n_20592, n_20593);
  and g50235 (n29738, n29529, n29737);
  not g50236 (n_20594, n29529);
  not g50237 (n_20595, n29737);
  and g50238 (n29739, n_20594, n_20595);
  not g50239 (n_20596, n29738);
  not g50240 (n_20597, n29739);
  and g50241 (\result[12] , n_20596, n_20597);
  and g50242 (n29741, n_20589, n_20593);
  and g50243 (n29742, n_20580, n_20583);
  and g50244 (n29743, n75, n23672);
  and g50245 (n29744, n3020, n22350);
  and g50246 (n29745, n3023, n22356);
  and g50247 (n29746, n3028, n22353);
  and g50255 (n29750, n_8091, n_19417);
  not g50256 (n_20602, n29750);
  and g50257 (n29751, \a[8] , n_20602);
  and g50258 (n29752, n_1106, n29750);
  not g50259 (n_20603, n29751);
  not g50260 (n_20604, n29752);
  and g50261 (n29753, n_20603, n_20604);
  and g50276 (n29768, n29355, n29767);
  not g50277 (n_20605, n29767);
  and g50278 (n29769, n_20298, n_20605);
  not g50279 (n_20606, n29768);
  not g50280 (n_20607, n29769);
  and g50281 (n29770, n_20606, n_20607);
  and g50282 (n29771, n29753, n29770);
  not g50283 (n_20608, n29753);
  not g50284 (n_20609, n29770);
  and g50285 (n29772, n_20608, n_20609);
  not g50286 (n_20610, n29771);
  not g50287 (n_20611, n29772);
  and g50288 (n29773, n_20610, n_20611);
  not g50289 (n_20612, n29570);
  and g50290 (n29774, n_20612, n29773);
  not g50291 (n_20613, n29773);
  and g50292 (n29775, n29570, n_20613);
  not g50293 (n_20614, n29774);
  not g50294 (n_20615, n29775);
  and g50295 (n29776, n_20614, n_20615);
  not g50296 (n_20616, n29749);
  and g50297 (n29777, n_20616, n29776);
  not g50298 (n_20617, n29777);
  and g50299 (n29778, n29776, n_20617);
  and g50300 (n29779, n_20616, n_20617);
  not g50301 (n_20618, n29778);
  not g50302 (n_20619, n29779);
  and g50303 (n29780, n_20618, n_20619);
  and g50304 (n29781, n3457, n22341);
  and g50305 (n29782, n3542, n22347);
  and g50306 (n29783, n3606, n22344);
  and g50312 (n29786, n3368, n24142);
  not g50315 (n_20624, n29787);
  and g50316 (n29788, \a[29] , n_20624);
  not g50317 (n_20625, n29788);
  and g50318 (n29789, \a[29] , n_20625);
  and g50319 (n29790, n_20624, n_20625);
  not g50320 (n_20626, n29789);
  not g50321 (n_20627, n29790);
  and g50322 (n29791, n_20626, n_20627);
  not g50323 (n_20628, n29780);
  not g50324 (n_20629, n29791);
  and g50325 (n29792, n_20628, n_20629);
  not g50326 (n_20630, n29792);
  and g50327 (n29793, n_20628, n_20630);
  and g50328 (n29794, n_20629, n_20630);
  not g50329 (n_20631, n29793);
  not g50330 (n_20632, n29794);
  and g50331 (n29795, n_20631, n_20632);
  and g50332 (n29796, n_20459, n_20465);
  and g50333 (n29797, n29795, n29796);
  not g50334 (n_20633, n29795);
  not g50335 (n_20634, n29796);
  and g50336 (n29798, n_20633, n_20634);
  not g50337 (n_20635, n29797);
  not g50338 (n_20636, n29798);
  and g50339 (n29799, n_20635, n_20636);
  and g50340 (n29800, n3884, n22332);
  and g50341 (n29801, n3967, n22338);
  and g50342 (n29802, n4046, n22335);
  and g50348 (n29805, n4050, n22542);
  not g50351 (n_20641, n29806);
  and g50352 (n29807, \a[26] , n_20641);
  not g50353 (n_20642, n29807);
  and g50354 (n29808, \a[26] , n_20642);
  and g50355 (n29809, n_20641, n_20642);
  not g50356 (n_20643, n29808);
  not g50357 (n_20644, n29809);
  and g50358 (n29810, n_20643, n_20644);
  not g50359 (n_20645, n29810);
  and g50360 (n29811, n29799, n_20645);
  not g50361 (n_20646, n29811);
  and g50362 (n29812, n29799, n_20646);
  and g50363 (n29813, n_20645, n_20646);
  not g50364 (n_20647, n29812);
  not g50365 (n_20648, n29813);
  and g50366 (n29814, n_20647, n_20648);
  and g50367 (n29815, n_20475, n_20488);
  and g50368 (n29816, n29814, n29815);
  not g50369 (n_20649, n29814);
  not g50370 (n_20650, n29815);
  and g50371 (n29817, n_20649, n_20650);
  not g50372 (n_20651, n29816);
  not g50373 (n_20652, n29817);
  and g50374 (n29818, n_20651, n_20652);
  and g50375 (n29819, n4694, n22323);
  and g50376 (n29820, n4533, n22329);
  and g50377 (n29821, n4604, n22326);
  and g50383 (n29824, n4536, n24599);
  not g50386 (n_20657, n29825);
  and g50387 (n29826, \a[23] , n_20657);
  not g50388 (n_20658, n29826);
  and g50389 (n29827, \a[23] , n_20658);
  and g50390 (n29828, n_20657, n_20658);
  not g50391 (n_20659, n29827);
  not g50392 (n_20660, n29828);
  and g50393 (n29829, n_20659, n_20660);
  not g50394 (n_20661, n29829);
  and g50395 (n29830, n29818, n_20661);
  not g50396 (n_20662, n29830);
  and g50397 (n29831, n29818, n_20662);
  and g50398 (n29832, n_20661, n_20662);
  not g50399 (n_20663, n29831);
  not g50400 (n_20664, n29832);
  and g50401 (n29833, n_20663, n_20664);
  and g50402 (n29834, n_20494, n_20504);
  and g50403 (n29835, n29833, n29834);
  not g50404 (n_20665, n29833);
  not g50405 (n_20666, n29834);
  and g50406 (n29836, n_20665, n_20666);
  not g50407 (n_20667, n29835);
  not g50408 (n_20668, n29836);
  and g50409 (n29837, n_20667, n_20668);
  and g50410 (n29838, n5496, n22315);
  and g50411 (n29839, n4935, n22320);
  and g50412 (n29840, n5407, n22312);
  and g50418 (n29843, n4938, n25294);
  not g50421 (n_20673, n29844);
  and g50422 (n29845, \a[20] , n_20673);
  not g50423 (n_20674, n29845);
  and g50424 (n29846, \a[20] , n_20674);
  and g50425 (n29847, n_20673, n_20674);
  not g50426 (n_20675, n29846);
  not g50427 (n_20676, n29847);
  and g50428 (n29848, n_20675, n_20676);
  not g50429 (n_20677, n29848);
  and g50430 (n29849, n29837, n_20677);
  not g50431 (n_20678, n29849);
  and g50432 (n29850, n29837, n_20678);
  and g50433 (n29851, n_20677, n_20678);
  not g50434 (n_20679, n29850);
  not g50435 (n_20680, n29851);
  and g50436 (n29852, n_20679, n_20680);
  and g50437 (n29853, n_20510, n_20520);
  and g50438 (n29854, n29852, n29853);
  not g50439 (n_20681, n29852);
  not g50440 (n_20682, n29853);
  and g50441 (n29855, n_20681, n_20682);
  not g50442 (n_20683, n29854);
  not g50443 (n_20684, n29855);
  and g50444 (n29856, n_20683, n_20684);
  and g50445 (n29857, n_20526, n_20536);
  and g50446 (n29858, n6233, n26066);
  and g50447 (n29859, n5663, n22309);
  and g50448 (n29860, n5939, n26063);
  and g50454 (n29863, n5666, n_18359);
  not g50457 (n_20689, n29864);
  and g50458 (n29865, \a[17] , n_20689);
  not g50459 (n_20690, n29865);
  and g50460 (n29866, \a[17] , n_20690);
  and g50461 (n29867, n_20689, n_20690);
  not g50462 (n_20691, n29866);
  not g50463 (n_20692, n29867);
  and g50464 (n29868, n_20691, n_20692);
  not g50465 (n_20693, n29857);
  not g50466 (n_20694, n29868);
  and g50467 (n29869, n_20693, n_20694);
  not g50468 (n_20695, n29869);
  and g50469 (n29870, n_20693, n_20695);
  and g50470 (n29871, n_20694, n_20695);
  not g50471 (n_20696, n29870);
  not g50472 (n_20697, n29871);
  and g50473 (n29872, n_20696, n_20697);
  not g50474 (n_20698, n29856);
  and g50475 (n29873, n_20698, n29872);
  not g50476 (n_20699, n29872);
  and g50477 (n29874, n29856, n_20699);
  not g50478 (n_20700, n29873);
  not g50479 (n_20701, n29874);
  and g50480 (n29875, n_20700, n_20701);
  and g50481 (n29876, n7101, n27173);
  and g50482 (n29877, n6402, n26060);
  and g50483 (n29878, n6951, n26890);
  and g50489 (n29881, n6397, n27185);
  not g50492 (n_20706, n29882);
  and g50493 (n29883, \a[14] , n_20706);
  not g50494 (n_20707, n29883);
  and g50495 (n29884, \a[14] , n_20707);
  and g50496 (n29885, n_20706, n_20707);
  not g50497 (n_20708, n29884);
  not g50498 (n_20709, n29885);
  and g50499 (n29886, n_20708, n_20709);
  not g50500 (n_20710, n29886);
  and g50501 (n29887, n29875, n_20710);
  not g50502 (n_20711, n29887);
  and g50503 (n29888, n29875, n_20711);
  and g50504 (n29889, n_20710, n_20711);
  not g50505 (n_20712, n29888);
  not g50506 (n_20713, n29889);
  and g50507 (n29890, n_20712, n_20713);
  and g50508 (n29891, n_20542, n_20552);
  and g50509 (n29892, n29890, n29891);
  not g50510 (n_20714, n29890);
  not g50511 (n_20715, n29891);
  and g50512 (n29893, n_20714, n_20715);
  not g50513 (n_20716, n29892);
  not g50514 (n_20717, n29893);
  and g50515 (n29894, n_20716, n_20717);
  and g50516 (n29895, n_20558, n_20568);
  and g50517 (n29896, n7983, n27964);
  and g50518 (n29897, n7291, n27442);
  and g50519 (n29898, n7632, n27698);
  and g50525 (n29901, n7294, n27976);
  not g50528 (n_20722, n29902);
  and g50529 (n29903, \a[11] , n_20722);
  not g50530 (n_20723, n29903);
  and g50531 (n29904, \a[11] , n_20723);
  and g50532 (n29905, n_20722, n_20723);
  not g50533 (n_20724, n29904);
  not g50534 (n_20725, n29905);
  and g50535 (n29906, n_20724, n_20725);
  not g50536 (n_20726, n29895);
  not g50537 (n_20727, n29906);
  and g50538 (n29907, n_20726, n_20727);
  not g50539 (n_20728, n29907);
  and g50540 (n29908, n_20726, n_20728);
  and g50541 (n29909, n_20727, n_20728);
  not g50542 (n_20729, n29908);
  not g50543 (n_20730, n29909);
  and g50544 (n29910, n_20729, n_20730);
  not g50545 (n_20731, n29894);
  and g50546 (n29911, n_20731, n29910);
  not g50547 (n_20732, n29910);
  and g50548 (n29912, n29894, n_20732);
  not g50549 (n_20733, n29911);
  not g50550 (n_20734, n29912);
  and g50551 (n29913, n_20733, n_20734);
  not g50552 (n_20735, n29742);
  and g50553 (n29914, n_20735, n29913);
  not g50554 (n_20736, n29913);
  and g50555 (n29915, n29742, n_20736);
  not g50556 (n_20737, n29914);
  not g50557 (n_20738, n29915);
  and g50558 (n29916, n_20737, n_20738);
  not g50559 (n_20739, n29741);
  and g50560 (n29917, n_20739, n29916);
  not g50561 (n_20740, n29916);
  and g50562 (n29918, n29741, n_20740);
  not g50563 (n_20741, n29917);
  not g50564 (n_20742, n29918);
  and g50565 (n29919, n_20741, n_20742);
  not g50566 (n_20743, n29919);
  and g50567 (n29920, n_20596, n_20743);
  and g50568 (n29921, n29738, n29919);
  not g50569 (n_20744, n29920);
  not g50570 (n_20745, n29921);
  and g50571 (\result[13] , n_20744, n_20745);
  and g50572 (n29923, n_20630, n_20636);
  and g50573 (n29924, n75, n_16069);
  and g50574 (n29925, n3020, n22347);
  and g50575 (n29926, n3023, n22353);
  and g50576 (n29927, n3028, n22350);
  and g50584 (n29931, n_20607, n_20610);
  not g50600 (n_20750, n29931);
  and g50601 (n29947, n_20750, n29946);
  not g50602 (n_20751, n29946);
  and g50603 (n29948, n29931, n_20751);
  not g50604 (n_20752, n29947);
  not g50605 (n_20753, n29948);
  and g50606 (n29949, n_20752, n_20753);
  not g50607 (n_20754, n29930);
  and g50608 (n29950, n_20754, n29949);
  not g50609 (n_20755, n29950);
  and g50610 (n29951, n_20754, n_20755);
  and g50611 (n29952, n29949, n_20755);
  not g50612 (n_20756, n29951);
  not g50613 (n_20757, n29952);
  and g50614 (n29953, n_20756, n_20757);
  and g50615 (n29954, n_20614, n_20617);
  and g50616 (n29955, n29953, n29954);
  not g50617 (n_20758, n29953);
  not g50618 (n_20759, n29954);
  and g50619 (n29956, n_20758, n_20759);
  not g50620 (n_20760, n29955);
  not g50621 (n_20761, n29956);
  and g50622 (n29957, n_20760, n_20761);
  and g50623 (n29958, n3457, n22338);
  and g50624 (n29959, n3542, n22344);
  and g50625 (n29960, n3606, n22341);
  not g50626 (n_20762, n29959);
  not g50627 (n_20763, n29960);
  and g50628 (n29961, n_20762, n_20763);
  not g50629 (n_20764, n29958);
  and g50630 (n29962, n_20764, n29961);
  and g50631 (n29963, n_489, n29962);
  and g50632 (n29964, n24188, n29962);
  not g50633 (n_20765, n29963);
  not g50634 (n_20766, n29964);
  and g50635 (n29965, n_20765, n_20766);
  not g50636 (n_20767, n29965);
  and g50637 (n29966, \a[29] , n_20767);
  and g50638 (n29967, n_15, n29965);
  not g50639 (n_20768, n29966);
  not g50640 (n_20769, n29967);
  and g50641 (n29968, n_20768, n_20769);
  not g50642 (n_20770, n29968);
  and g50643 (n29969, n29957, n_20770);
  not g50644 (n_20771, n29957);
  and g50645 (n29970, n_20771, n29968);
  not g50646 (n_20772, n29969);
  not g50647 (n_20773, n29970);
  and g50648 (n29971, n_20772, n_20773);
  not g50649 (n_20774, n29923);
  and g50650 (n29972, n_20774, n29971);
  not g50651 (n_20775, n29971);
  and g50652 (n29973, n29923, n_20775);
  not g50653 (n_20776, n29972);
  not g50654 (n_20777, n29973);
  and g50655 (n29974, n_20776, n_20777);
  and g50656 (n29975, n3884, n22329);
  and g50657 (n29976, n3967, n22335);
  and g50658 (n29977, n4046, n22332);
  and g50664 (n29980, n4050, n_16827);
  not g50667 (n_20782, n29981);
  and g50668 (n29982, \a[26] , n_20782);
  not g50669 (n_20783, n29982);
  and g50670 (n29983, \a[26] , n_20783);
  and g50671 (n29984, n_20782, n_20783);
  not g50672 (n_20784, n29983);
  not g50673 (n_20785, n29984);
  and g50674 (n29985, n_20784, n_20785);
  not g50675 (n_20786, n29985);
  and g50676 (n29986, n29974, n_20786);
  not g50677 (n_20787, n29986);
  and g50678 (n29987, n29974, n_20787);
  and g50679 (n29988, n_20786, n_20787);
  not g50680 (n_20788, n29987);
  not g50681 (n_20789, n29988);
  and g50682 (n29989, n_20788, n_20789);
  and g50683 (n29990, n_20646, n_20652);
  and g50684 (n29991, n29989, n29990);
  not g50685 (n_20790, n29989);
  not g50686 (n_20791, n29990);
  and g50687 (n29992, n_20790, n_20791);
  not g50688 (n_20792, n29991);
  not g50689 (n_20793, n29992);
  and g50690 (n29993, n_20792, n_20793);
  and g50691 (n29994, n4694, n22320);
  and g50692 (n29995, n4533, n22326);
  and g50693 (n29996, n4604, n22323);
  and g50699 (n29999, n4536, n_17020);
  not g50702 (n_20798, n30000);
  and g50703 (n30001, \a[23] , n_20798);
  not g50704 (n_20799, n30001);
  and g50705 (n30002, \a[23] , n_20799);
  and g50706 (n30003, n_20798, n_20799);
  not g50707 (n_20800, n30002);
  not g50708 (n_20801, n30003);
  and g50709 (n30004, n_20800, n_20801);
  not g50710 (n_20802, n30004);
  and g50711 (n30005, n29993, n_20802);
  not g50712 (n_20803, n30005);
  and g50713 (n30006, n29993, n_20803);
  and g50714 (n30007, n_20802, n_20803);
  not g50715 (n_20804, n30006);
  not g50716 (n_20805, n30007);
  and g50717 (n30008, n_20804, n_20805);
  and g50718 (n30009, n_20662, n_20668);
  and g50719 (n30010, n30008, n30009);
  not g50720 (n_20806, n30008);
  not g50721 (n_20807, n30009);
  and g50722 (n30011, n_20806, n_20807);
  not g50723 (n_20808, n30010);
  not g50724 (n_20809, n30011);
  and g50725 (n30012, n_20808, n_20809);
  and g50726 (n30013, n5496, n22309);
  and g50727 (n30014, n4935, n22312);
  and g50728 (n30015, n5407, n22315);
  and g50734 (n30018, n4938, n_14657);
  not g50737 (n_20814, n30019);
  and g50738 (n30020, \a[20] , n_20814);
  not g50739 (n_20815, n30020);
  and g50740 (n30021, \a[20] , n_20815);
  and g50741 (n30022, n_20814, n_20815);
  not g50742 (n_20816, n30021);
  not g50743 (n_20817, n30022);
  and g50744 (n30023, n_20816, n_20817);
  not g50745 (n_20818, n30023);
  and g50746 (n30024, n30012, n_20818);
  not g50747 (n_20819, n30024);
  and g50748 (n30025, n30012, n_20819);
  and g50749 (n30026, n_20818, n_20819);
  not g50750 (n_20820, n30025);
  not g50751 (n_20821, n30026);
  and g50752 (n30027, n_20820, n_20821);
  and g50753 (n30028, n_20678, n_20684);
  and g50754 (n30029, n30027, n30028);
  not g50755 (n_20822, n30027);
  not g50756 (n_20823, n30028);
  and g50757 (n30030, n_20822, n_20823);
  not g50758 (n_20824, n30029);
  not g50759 (n_20825, n30030);
  and g50760 (n30031, n_20824, n_20825);
  and g50761 (n30032, n6233, n26060);
  and g50762 (n30033, n5663, n26063);
  and g50763 (n30034, n5939, n26066);
  and g50769 (n30037, n5666, n_18596);
  not g50772 (n_20830, n30038);
  and g50773 (n30039, \a[17] , n_20830);
  not g50774 (n_20831, n30039);
  and g50775 (n30040, \a[17] , n_20831);
  and g50776 (n30041, n_20830, n_20831);
  not g50777 (n_20832, n30040);
  not g50778 (n_20833, n30041);
  and g50779 (n30042, n_20832, n_20833);
  not g50780 (n_20834, n30042);
  and g50781 (n30043, n30031, n_20834);
  not g50782 (n_20835, n30043);
  and g50783 (n30044, n30031, n_20835);
  and g50784 (n30045, n_20834, n_20835);
  not g50785 (n_20836, n30044);
  not g50786 (n_20837, n30045);
  and g50787 (n30046, n_20836, n_20837);
  and g50788 (n30047, n_20695, n_20701);
  not g50789 (n_20838, n30046);
  not g50790 (n_20839, n30047);
  and g50791 (n30048, n_20838, n_20839);
  not g50792 (n_20840, n30048);
  and g50793 (n30049, n_20838, n_20840);
  and g50794 (n30050, n_20839, n_20840);
  not g50795 (n_20841, n30049);
  not g50796 (n_20842, n30050);
  and g50797 (n30051, n_20841, n_20842);
  and g50798 (n30052, n7101, n27442);
  and g50799 (n30053, n6402, n26890);
  and g50800 (n30054, n6951, n27173);
  and g50806 (n30057, n6397, n27455);
  not g50809 (n_20847, n30058);
  and g50810 (n30059, \a[14] , n_20847);
  not g50811 (n_20848, n30059);
  and g50812 (n30060, \a[14] , n_20848);
  and g50813 (n30061, n_20847, n_20848);
  not g50814 (n_20849, n30060);
  not g50815 (n_20850, n30061);
  and g50816 (n30062, n_20849, n_20850);
  not g50817 (n_20851, n30051);
  not g50818 (n_20852, n30062);
  and g50819 (n30063, n_20851, n_20852);
  not g50820 (n_20853, n30063);
  and g50821 (n30064, n_20851, n_20853);
  and g50822 (n30065, n_20852, n_20853);
  not g50823 (n_20854, n30064);
  not g50824 (n_20855, n30065);
  and g50825 (n30066, n_20854, n_20855);
  and g50826 (n30067, n_20711, n_20717);
  and g50827 (n30068, n30066, n30067);
  not g50828 (n_20856, n30066);
  not g50829 (n_20857, n30067);
  and g50830 (n30069, n_20856, n_20857);
  not g50831 (n_20858, n30068);
  not g50832 (n_20859, n30069);
  and g50833 (n30070, n_20858, n_20859);
  and g50834 (n30071, n7983, n_19417);
  and g50835 (n30072, n7291, n27698);
  and g50836 (n30073, n7632, n27964);
  and g50842 (n30076, n7294, n_19940);
  not g50845 (n_20864, n30077);
  and g50846 (n30078, \a[11] , n_20864);
  not g50847 (n_20865, n30078);
  and g50848 (n30079, \a[11] , n_20865);
  and g50849 (n30080, n_20864, n_20865);
  not g50850 (n_20866, n30079);
  not g50851 (n_20867, n30080);
  and g50852 (n30081, n_20866, n_20867);
  not g50853 (n_20868, n30081);
  and g50854 (n30082, n30070, n_20868);
  not g50855 (n_20869, n30082);
  and g50856 (n30083, n30070, n_20869);
  and g50857 (n30084, n_20868, n_20869);
  not g50858 (n_20870, n30083);
  not g50859 (n_20871, n30084);
  and g50860 (n30085, n_20870, n_20871);
  and g50861 (n30086, n_20728, n_20734);
  not g50862 (n_20872, n30085);
  not g50863 (n_20873, n30086);
  and g50864 (n30087, n_20872, n_20873);
  not g50865 (n_20874, n30087);
  and g50866 (n30088, n_20872, n_20874);
  and g50867 (n30089, n_20873, n_20874);
  not g50868 (n_20875, n30088);
  not g50869 (n_20876, n30089);
  and g50870 (n30090, n_20875, n_20876);
  and g50871 (n30091, n_20737, n_20741);
  and g50872 (n30092, n30090, n30091);
  not g50873 (n_20877, n30090);
  not g50874 (n_20878, n30091);
  and g50875 (n30093, n_20877, n_20878);
  not g50876 (n_20879, n30092);
  not g50877 (n_20880, n30093);
  and g50878 (n30094, n_20879, n_20880);
  not g50879 (n_20881, n30094);
  and g50880 (n30095, n29921, n_20881);
  and g50881 (n30096, n_20745, n30094);
  or g50882 (\result[14] , n30095, n30096);
  and g50883 (n30098, n_20761, n_20772);
  and g50884 (n30099, n_20752, n_20755);
  and g50903 (n30118, n_20751, n30117);
  not g50904 (n_20882, n30117);
  and g50905 (n30119, n29946, n_20882);
  not g50906 (n_20883, n30099);
  not g50907 (n_20884, n30119);
  and g50908 (n30120, n_20883, n_20884);
  not g50909 (n_20885, n30118);
  and g50910 (n30121, n_20885, n30120);
  not g50911 (n_20886, n30121);
  and g50912 (n30122, n_20883, n_20886);
  and g50913 (n30123, n_20884, n_20886);
  and g50914 (n30124, n_20885, n30123);
  not g50915 (n_20887, n30122);
  not g50916 (n_20888, n30124);
  and g50917 (n30125, n_20887, n_20888);
  and g50918 (n30126, n75, n_18142);
  and g50919 (n30127, n3020, n22344);
  and g50920 (n30128, n3023, n22350);
  and g50921 (n30129, n3028, n22347);
  not g50929 (n_20893, n30125);
  not g50930 (n_20894, n30132);
  and g50931 (n30133, n_20893, n_20894);
  not g50932 (n_20895, n30133);
  and g50933 (n30134, n_20893, n_20895);
  and g50934 (n30135, n_20894, n_20895);
  not g50935 (n_20896, n30134);
  not g50936 (n_20897, n30135);
  and g50937 (n30136, n_20896, n_20897);
  and g50938 (n30137, n3457, n22335);
  and g50939 (n30138, n3542, n22341);
  and g50940 (n30139, n3606, n22338);
  not g50941 (n_20898, n30138);
  not g50942 (n_20899, n30139);
  and g50943 (n30140, n_20898, n_20899);
  not g50944 (n_20900, n30137);
  and g50945 (n30141, n_20900, n30140);
  and g50946 (n30142, n_489, n30141);
  and g50947 (n30143, n24167, n30141);
  not g50948 (n_20901, n30142);
  not g50949 (n_20902, n30143);
  and g50950 (n30144, n_20901, n_20902);
  not g50951 (n_20903, n30144);
  and g50952 (n30145, \a[29] , n_20903);
  and g50953 (n30146, n_15, n30144);
  not g50954 (n_20904, n30145);
  not g50955 (n_20905, n30146);
  and g50956 (n30147, n_20904, n_20905);
  not g50957 (n_20906, n30136);
  not g50958 (n_20907, n30147);
  and g50959 (n30148, n_20906, n_20907);
  and g50960 (n30149, n30136, n30147);
  not g50961 (n_20908, n30148);
  not g50962 (n_20909, n30149);
  and g50963 (n30150, n_20908, n_20909);
  not g50964 (n_20910, n30098);
  and g50965 (n30151, n_20910, n30150);
  not g50966 (n_20911, n30150);
  and g50967 (n30152, n30098, n_20911);
  not g50968 (n_20912, n30151);
  not g50969 (n_20913, n30152);
  and g50970 (n30153, n_20912, n_20913);
  and g50971 (n30154, n3884, n22326);
  and g50972 (n30155, n3967, n22332);
  and g50973 (n30156, n4046, n22329);
  and g50979 (n30159, n4050, n_18133);
  not g50982 (n_20918, n30160);
  and g50983 (n30161, \a[26] , n_20918);
  not g50984 (n_20919, n30161);
  and g50985 (n30162, \a[26] , n_20919);
  and g50986 (n30163, n_20918, n_20919);
  not g50987 (n_20920, n30162);
  not g50988 (n_20921, n30163);
  and g50989 (n30164, n_20920, n_20921);
  not g50990 (n_20922, n30164);
  and g50991 (n30165, n30153, n_20922);
  not g50992 (n_20923, n30165);
  and g50993 (n30166, n30153, n_20923);
  and g50994 (n30167, n_20922, n_20923);
  not g50995 (n_20924, n30166);
  not g50996 (n_20925, n30167);
  and g50997 (n30168, n_20924, n_20925);
  and g50998 (n30169, n_20776, n_20787);
  and g50999 (n30170, n30168, n30169);
  not g51000 (n_20926, n30168);
  not g51001 (n_20927, n30169);
  and g51002 (n30171, n_20926, n_20927);
  not g51003 (n_20928, n30170);
  not g51004 (n_20929, n30171);
  and g51005 (n30172, n_20928, n_20929);
  and g51006 (n30173, n4694, n22312);
  and g51007 (n30174, n4533, n22323);
  and g51008 (n30175, n4604, n22320);
  and g51014 (n30178, n4536, n_17004);
  not g51017 (n_20934, n30179);
  and g51018 (n30180, \a[23] , n_20934);
  not g51019 (n_20935, n30180);
  and g51020 (n30181, \a[23] , n_20935);
  and g51021 (n30182, n_20934, n_20935);
  not g51022 (n_20936, n30181);
  not g51023 (n_20937, n30182);
  and g51024 (n30183, n_20936, n_20937);
  not g51025 (n_20938, n30183);
  and g51026 (n30184, n30172, n_20938);
  not g51027 (n_20939, n30184);
  and g51028 (n30185, n30172, n_20939);
  and g51029 (n30186, n_20938, n_20939);
  not g51030 (n_20940, n30185);
  not g51031 (n_20941, n30186);
  and g51032 (n30187, n_20940, n_20941);
  and g51033 (n30188, n_20793, n_20803);
  and g51034 (n30189, n30187, n30188);
  not g51035 (n_20942, n30187);
  not g51036 (n_20943, n30188);
  and g51037 (n30190, n_20942, n_20943);
  not g51038 (n_20944, n30189);
  not g51039 (n_20945, n30190);
  and g51040 (n30191, n_20944, n_20945);
  and g51041 (n30192, n5496, n26063);
  and g51042 (n30193, n4935, n22315);
  and g51043 (n30194, n5407, n22309);
  and g51049 (n30197, n4938, n_18124);
  not g51052 (n_20950, n30198);
  and g51053 (n30199, \a[20] , n_20950);
  not g51054 (n_20951, n30199);
  and g51055 (n30200, \a[20] , n_20951);
  and g51056 (n30201, n_20950, n_20951);
  not g51057 (n_20952, n30200);
  not g51058 (n_20953, n30201);
  and g51059 (n30202, n_20952, n_20953);
  not g51060 (n_20954, n30202);
  and g51061 (n30203, n30191, n_20954);
  not g51062 (n_20955, n30203);
  and g51063 (n30204, n30191, n_20955);
  and g51064 (n30205, n_20954, n_20955);
  not g51065 (n_20956, n30204);
  not g51066 (n_20957, n30205);
  and g51067 (n30206, n_20956, n_20957);
  and g51068 (n30207, n_20809, n_20819);
  and g51069 (n30208, n30206, n30207);
  not g51070 (n_20958, n30206);
  not g51071 (n_20959, n30207);
  and g51072 (n30209, n_20958, n_20959);
  not g51073 (n_20960, n30208);
  not g51074 (n_20961, n30209);
  and g51075 (n30210, n_20960, n_20961);
  and g51076 (n30211, n6233, n26890);
  and g51077 (n30212, n5663, n26066);
  and g51078 (n30213, n5939, n26060);
  and g51084 (n30216, n5666, n_18823);
  not g51087 (n_20966, n30217);
  and g51088 (n30218, \a[17] , n_20966);
  not g51089 (n_20967, n30218);
  and g51090 (n30219, \a[17] , n_20967);
  and g51091 (n30220, n_20966, n_20967);
  not g51092 (n_20968, n30219);
  not g51093 (n_20969, n30220);
  and g51094 (n30221, n_20968, n_20969);
  not g51095 (n_20970, n30221);
  and g51096 (n30222, n30210, n_20970);
  not g51097 (n_20971, n30222);
  and g51098 (n30223, n30210, n_20971);
  and g51099 (n30224, n_20970, n_20971);
  not g51100 (n_20972, n30223);
  not g51101 (n_20973, n30224);
  and g51102 (n30225, n_20972, n_20973);
  and g51103 (n30226, n_20825, n_20835);
  and g51104 (n30227, n30225, n30226);
  not g51105 (n_20974, n30225);
  not g51106 (n_20975, n30226);
  and g51107 (n30228, n_20974, n_20975);
  not g51108 (n_20976, n30227);
  not g51109 (n_20977, n30228);
  and g51110 (n30229, n_20976, n_20977);
  and g51111 (n30230, n7101, n27698);
  and g51112 (n30231, n6402, n27173);
  and g51113 (n30232, n6951, n27442);
  and g51119 (n30235, n6397, n_19446);
  not g51122 (n_20982, n30236);
  and g51123 (n30237, \a[14] , n_20982);
  not g51124 (n_20983, n30237);
  and g51125 (n30238, \a[14] , n_20983);
  and g51126 (n30239, n_20982, n_20983);
  not g51127 (n_20984, n30238);
  not g51128 (n_20985, n30239);
  and g51129 (n30240, n_20984, n_20985);
  not g51130 (n_20986, n30240);
  and g51131 (n30241, n30229, n_20986);
  not g51132 (n_20987, n30241);
  and g51133 (n30242, n30229, n_20987);
  and g51134 (n30243, n_20986, n_20987);
  not g51135 (n_20988, n30242);
  not g51136 (n_20989, n30243);
  and g51137 (n30244, n_20988, n_20989);
  and g51138 (n30245, n_20840, n_20853);
  and g51139 (n30246, n_9481, n_19417);
  and g51140 (n30247, n7291, n27964);
  not g51141 (n_20990, n30246);
  not g51142 (n_20991, n30247);
  and g51143 (n30248, n_20990, n_20991);
  and g51144 (n30249, n_2446, n30248);
  and g51145 (n30250, n28221, n30248);
  not g51146 (n_20992, n30249);
  not g51147 (n_20993, n30250);
  and g51148 (n30251, n_20992, n_20993);
  not g51149 (n_20994, n30251);
  and g51150 (n30252, \a[11] , n_20994);
  and g51151 (n30253, n_1071, n30251);
  not g51152 (n_20995, n30252);
  not g51153 (n_20996, n30253);
  and g51154 (n30254, n_20995, n_20996);
  not g51155 (n_20997, n30245);
  not g51156 (n_20998, n30254);
  and g51157 (n30255, n_20997, n_20998);
  and g51158 (n30256, n30245, n30254);
  not g51159 (n_20999, n30255);
  not g51160 (n_21000, n30256);
  and g51161 (n30257, n_20999, n_21000);
  not g51162 (n_21001, n30244);
  and g51163 (n30258, n_21001, n30257);
  not g51164 (n_21002, n30258);
  and g51165 (n30259, n_21001, n_21002);
  and g51166 (n30260, n30257, n_21002);
  not g51167 (n_21003, n30259);
  not g51168 (n_21004, n30260);
  and g51169 (n30261, n_21003, n_21004);
  and g51170 (n30262, n_20859, n_20869);
  and g51171 (n30263, n30261, n30262);
  not g51172 (n_21005, n30261);
  not g51173 (n_21006, n30262);
  and g51174 (n30264, n_21005, n_21006);
  not g51175 (n_21007, n30263);
  not g51176 (n_21008, n30264);
  and g51177 (n30265, n_21007, n_21008);
  and g51178 (n30266, n_20874, n_20880);
  not g51179 (n_21009, n30265);
  and g51180 (n30267, n_21009, n30266);
  not g51181 (n_21010, n30266);
  and g51182 (n30268, n30265, n_21010);
  not g51183 (n_21011, n30267);
  not g51184 (n_21012, n30268);
  and g51185 (n30269, n_21011, n_21012);
  and g51186 (n30270, n29921, n30094);
  and g51187 (n30271, n30269, n30270);
  not g51188 (n_21013, n30269);
  not g51189 (n_21014, n30270);
  and g51190 (n30272, n_21013, n_21014);
  not g51191 (n_21015, n30271);
  not g51192 (n_21016, n30272);
  and g51193 (\result[15] , n_21015, n_21016);
  and g51194 (n30274, n_21008, n_21012);
  and g51195 (n30275, n_20999, n_21002);
  and g51196 (n30276, n_20895, n_20908);
  and g51197 (n30277, n75, n24142);
  and g51198 (n30278, n3020, n22341);
  and g51199 (n30279, n3023, n22347);
  and g51200 (n30280, n3028, n22344);
  and g51208 (n30284, n_8049, n_19417);
  not g51209 (n_21021, n30284);
  and g51210 (n30285, \a[11] , n_21021);
  and g51211 (n30286, n_1071, n30284);
  not g51212 (n_21022, n30285);
  not g51213 (n_21023, n30286);
  and g51214 (n30287, n_21022, n_21023);
  and g51231 (n30304, n29946, n30303);
  not g51232 (n_21024, n30303);
  and g51233 (n30305, n_20751, n_21024);
  not g51234 (n_21025, n30304);
  not g51235 (n_21026, n30305);
  and g51236 (n30306, n_21025, n_21026);
  and g51237 (n30307, n30287, n30306);
  not g51238 (n_21027, n30287);
  not g51239 (n_21028, n30306);
  and g51240 (n30308, n_21027, n_21028);
  not g51241 (n_21029, n30307);
  not g51242 (n_21030, n30308);
  and g51243 (n30309, n_21029, n_21030);
  not g51244 (n_21031, n30283);
  and g51245 (n30310, n_21031, n30309);
  not g51246 (n_21032, n30310);
  and g51247 (n30311, n30309, n_21032);
  and g51248 (n30312, n_21031, n_21032);
  not g51249 (n_21033, n30311);
  not g51250 (n_21034, n30312);
  and g51251 (n30313, n_21033, n_21034);
  not g51252 (n_21035, n30123);
  not g51253 (n_21036, n30313);
  and g51254 (n30314, n_21035, n_21036);
  not g51255 (n_21037, n30314);
  and g51256 (n30315, n_21036, n_21037);
  and g51257 (n30316, n_21035, n_21037);
  not g51258 (n_21038, n30315);
  not g51259 (n_21039, n30316);
  and g51260 (n30317, n_21038, n_21039);
  not g51261 (n_21040, n30276);
  not g51262 (n_21041, n30317);
  and g51263 (n30318, n_21040, n_21041);
  not g51264 (n_21042, n30318);
  and g51265 (n30319, n_21040, n_21042);
  and g51266 (n30320, n_21041, n_21042);
  not g51267 (n_21043, n30319);
  not g51268 (n_21044, n30320);
  and g51269 (n30321, n_21043, n_21044);
  and g51270 (n30322, n3457, n22332);
  and g51271 (n30323, n3542, n22338);
  and g51272 (n30324, n3606, n22335);
  and g51278 (n30327, n3368, n22542);
  not g51281 (n_21049, n30328);
  and g51282 (n30329, \a[29] , n_21049);
  not g51283 (n_21050, n30329);
  and g51284 (n30330, \a[29] , n_21050);
  and g51285 (n30331, n_21049, n_21050);
  not g51286 (n_21051, n30330);
  not g51287 (n_21052, n30331);
  and g51288 (n30332, n_21051, n_21052);
  not g51289 (n_21053, n30321);
  not g51290 (n_21054, n30332);
  and g51291 (n30333, n_21053, n_21054);
  not g51292 (n_21055, n30333);
  and g51293 (n30334, n_21053, n_21055);
  and g51294 (n30335, n_21054, n_21055);
  not g51295 (n_21056, n30334);
  not g51296 (n_21057, n30335);
  and g51297 (n30336, n_21056, n_21057);
  and g51298 (n30337, n3884, n22323);
  and g51299 (n30338, n3967, n22329);
  and g51300 (n30339, n4046, n22326);
  and g51306 (n30342, n4050, n24599);
  not g51309 (n_21062, n30343);
  and g51310 (n30344, \a[26] , n_21062);
  not g51311 (n_21063, n30344);
  and g51312 (n30345, \a[26] , n_21063);
  and g51313 (n30346, n_21062, n_21063);
  not g51314 (n_21064, n30345);
  not g51315 (n_21065, n30346);
  and g51316 (n30347, n_21064, n_21065);
  not g51317 (n_21066, n30336);
  not g51318 (n_21067, n30347);
  and g51319 (n30348, n_21066, n_21067);
  not g51320 (n_21068, n30348);
  and g51321 (n30349, n_21066, n_21068);
  and g51322 (n30350, n_21067, n_21068);
  not g51323 (n_21069, n30349);
  not g51324 (n_21070, n30350);
  and g51325 (n30351, n_21069, n_21070);
  and g51326 (n30352, n_20912, n_20923);
  and g51327 (n30353, n30351, n30352);
  not g51328 (n_21071, n30351);
  not g51329 (n_21072, n30352);
  and g51330 (n30354, n_21071, n_21072);
  not g51331 (n_21073, n30353);
  not g51332 (n_21074, n30354);
  and g51333 (n30355, n_21073, n_21074);
  and g51334 (n30356, n4694, n22315);
  and g51335 (n30357, n4533, n22320);
  and g51336 (n30358, n4604, n22312);
  and g51342 (n30361, n4536, n25294);
  not g51345 (n_21079, n30362);
  and g51346 (n30363, \a[23] , n_21079);
  not g51347 (n_21080, n30363);
  and g51348 (n30364, \a[23] , n_21080);
  and g51349 (n30365, n_21079, n_21080);
  not g51350 (n_21081, n30364);
  not g51351 (n_21082, n30365);
  and g51352 (n30366, n_21081, n_21082);
  not g51353 (n_21083, n30366);
  and g51354 (n30367, n30355, n_21083);
  not g51355 (n_21084, n30367);
  and g51356 (n30368, n30355, n_21084);
  and g51357 (n30369, n_21083, n_21084);
  not g51358 (n_21085, n30368);
  not g51359 (n_21086, n30369);
  and g51360 (n30370, n_21085, n_21086);
  and g51361 (n30371, n_20929, n_20939);
  and g51362 (n30372, n30370, n30371);
  not g51363 (n_21087, n30370);
  not g51364 (n_21088, n30371);
  and g51365 (n30373, n_21087, n_21088);
  not g51366 (n_21089, n30372);
  not g51367 (n_21090, n30373);
  and g51368 (n30374, n_21089, n_21090);
  and g51369 (n30375, n_20945, n_20955);
  and g51370 (n30376, n5496, n26066);
  and g51371 (n30377, n4935, n22309);
  and g51372 (n30378, n5407, n26063);
  and g51378 (n30381, n4938, n_18359);
  not g51381 (n_21095, n30382);
  and g51382 (n30383, \a[20] , n_21095);
  not g51383 (n_21096, n30383);
  and g51384 (n30384, \a[20] , n_21096);
  and g51385 (n30385, n_21095, n_21096);
  not g51386 (n_21097, n30384);
  not g51387 (n_21098, n30385);
  and g51388 (n30386, n_21097, n_21098);
  not g51389 (n_21099, n30375);
  not g51390 (n_21100, n30386);
  and g51391 (n30387, n_21099, n_21100);
  not g51392 (n_21101, n30387);
  and g51393 (n30388, n_21099, n_21101);
  and g51394 (n30389, n_21100, n_21101);
  not g51395 (n_21102, n30388);
  not g51396 (n_21103, n30389);
  and g51397 (n30390, n_21102, n_21103);
  not g51398 (n_21104, n30374);
  and g51399 (n30391, n_21104, n30390);
  not g51400 (n_21105, n30390);
  and g51401 (n30392, n30374, n_21105);
  not g51402 (n_21106, n30391);
  not g51403 (n_21107, n30392);
  and g51404 (n30393, n_21106, n_21107);
  and g51405 (n30394, n6233, n27173);
  and g51406 (n30395, n5663, n26060);
  and g51407 (n30396, n5939, n26890);
  and g51413 (n30399, n5666, n27185);
  not g51416 (n_21112, n30400);
  and g51417 (n30401, \a[17] , n_21112);
  not g51418 (n_21113, n30401);
  and g51419 (n30402, \a[17] , n_21113);
  and g51420 (n30403, n_21112, n_21113);
  not g51421 (n_21114, n30402);
  not g51422 (n_21115, n30403);
  and g51423 (n30404, n_21114, n_21115);
  not g51424 (n_21116, n30404);
  and g51425 (n30405, n30393, n_21116);
  not g51426 (n_21117, n30405);
  and g51427 (n30406, n30393, n_21117);
  and g51428 (n30407, n_21116, n_21117);
  not g51429 (n_21118, n30406);
  not g51430 (n_21119, n30407);
  and g51431 (n30408, n_21118, n_21119);
  and g51432 (n30409, n_20961, n_20971);
  and g51433 (n30410, n30408, n30409);
  not g51434 (n_21120, n30408);
  not g51435 (n_21121, n30409);
  and g51436 (n30411, n_21120, n_21121);
  not g51437 (n_21122, n30410);
  not g51438 (n_21123, n30411);
  and g51439 (n30412, n_21122, n_21123);
  and g51440 (n30413, n_20977, n_20987);
  and g51441 (n30414, n7101, n27964);
  and g51442 (n30415, n6402, n27442);
  and g51443 (n30416, n6951, n27698);
  and g51449 (n30419, n6397, n27976);
  not g51452 (n_21128, n30420);
  and g51453 (n30421, \a[14] , n_21128);
  not g51454 (n_21129, n30421);
  and g51455 (n30422, \a[14] , n_21129);
  and g51456 (n30423, n_21128, n_21129);
  not g51457 (n_21130, n30422);
  not g51458 (n_21131, n30423);
  and g51459 (n30424, n_21130, n_21131);
  not g51460 (n_21132, n30413);
  not g51461 (n_21133, n30424);
  and g51462 (n30425, n_21132, n_21133);
  not g51463 (n_21134, n30425);
  and g51464 (n30426, n_21132, n_21134);
  and g51465 (n30427, n_21133, n_21134);
  not g51466 (n_21135, n30426);
  not g51467 (n_21136, n30427);
  and g51468 (n30428, n_21135, n_21136);
  not g51469 (n_21137, n30412);
  and g51470 (n30429, n_21137, n30428);
  not g51471 (n_21138, n30428);
  and g51472 (n30430, n30412, n_21138);
  not g51473 (n_21139, n30429);
  not g51474 (n_21140, n30430);
  and g51475 (n30431, n_21139, n_21140);
  not g51476 (n_21141, n30275);
  and g51477 (n30432, n_21141, n30431);
  not g51478 (n_21142, n30431);
  and g51479 (n30433, n30275, n_21142);
  not g51480 (n_21143, n30432);
  not g51481 (n_21144, n30433);
  and g51482 (n30434, n_21143, n_21144);
  not g51483 (n_21145, n30274);
  and g51484 (n30435, n_21145, n30434);
  not g51485 (n_21146, n30434);
  and g51486 (n30436, n30274, n_21146);
  not g51487 (n_21147, n30435);
  not g51488 (n_21148, n30436);
  and g51489 (n30437, n_21147, n_21148);
  not g51490 (n_21149, n30437);
  and g51491 (n30438, n_21015, n_21149);
  and g51492 (n30439, n30271, n30437);
  not g51493 (n_21150, n30438);
  not g51494 (n_21151, n30439);
  and g51495 (\result[16] , n_21150, n_21151);
  and g51496 (n30441, n_21042, n_21055);
  and g51497 (n30442, n75, n_16033);
  and g51498 (n30443, n3020, n22338);
  and g51499 (n30444, n3023, n22344);
  and g51500 (n30445, n3028, n22341);
  and g51508 (n30449, n_21026, n_21029);
  not g51524 (n_21156, n30449);
  and g51525 (n30465, n_21156, n30464);
  not g51526 (n_21157, n30464);
  and g51527 (n30466, n30449, n_21157);
  not g51528 (n_21158, n30465);
  not g51529 (n_21159, n30466);
  and g51530 (n30467, n_21158, n_21159);
  not g51531 (n_21160, n30448);
  and g51532 (n30468, n_21160, n30467);
  not g51533 (n_21161, n30468);
  and g51534 (n30469, n_21160, n_21161);
  and g51535 (n30470, n30467, n_21161);
  not g51536 (n_21162, n30469);
  not g51537 (n_21163, n30470);
  and g51538 (n30471, n_21162, n_21163);
  and g51539 (n30472, n_21032, n_21037);
  and g51540 (n30473, n30471, n30472);
  not g51541 (n_21164, n30471);
  not g51542 (n_21165, n30472);
  and g51543 (n30474, n_21164, n_21165);
  not g51544 (n_21166, n30473);
  not g51545 (n_21167, n30474);
  and g51546 (n30475, n_21166, n_21167);
  and g51547 (n30476, n3457, n22329);
  and g51548 (n30477, n3542, n22335);
  and g51549 (n30478, n3606, n22332);
  not g51550 (n_21168, n30477);
  not g51551 (n_21169, n30478);
  and g51552 (n30479, n_21168, n_21169);
  not g51553 (n_21170, n30476);
  and g51554 (n30480, n_21170, n30479);
  and g51555 (n30481, n_489, n30480);
  and g51556 (n30482, n24633, n30480);
  not g51557 (n_21171, n30481);
  not g51558 (n_21172, n30482);
  and g51559 (n30483, n_21171, n_21172);
  not g51560 (n_21173, n30483);
  and g51561 (n30484, \a[29] , n_21173);
  and g51562 (n30485, n_15, n30483);
  not g51563 (n_21174, n30484);
  not g51564 (n_21175, n30485);
  and g51565 (n30486, n_21174, n_21175);
  not g51566 (n_21176, n30486);
  and g51567 (n30487, n30475, n_21176);
  not g51568 (n_21177, n30475);
  and g51569 (n30488, n_21177, n30486);
  not g51570 (n_21178, n30487);
  not g51571 (n_21179, n30488);
  and g51572 (n30489, n_21178, n_21179);
  not g51573 (n_21180, n30441);
  and g51574 (n30490, n_21180, n30489);
  not g51575 (n_21181, n30489);
  and g51576 (n30491, n30441, n_21181);
  not g51577 (n_21182, n30490);
  not g51578 (n_21183, n30491);
  and g51579 (n30492, n_21182, n_21183);
  and g51580 (n30493, n3884, n22320);
  and g51581 (n30494, n3967, n22326);
  and g51582 (n30495, n4046, n22323);
  and g51588 (n30498, n4050, n_17020);
  not g51591 (n_21188, n30499);
  and g51592 (n30500, \a[26] , n_21188);
  not g51593 (n_21189, n30500);
  and g51594 (n30501, \a[26] , n_21189);
  and g51595 (n30502, n_21188, n_21189);
  not g51596 (n_21190, n30501);
  not g51597 (n_21191, n30502);
  and g51598 (n30503, n_21190, n_21191);
  not g51599 (n_21192, n30503);
  and g51600 (n30504, n30492, n_21192);
  not g51601 (n_21193, n30504);
  and g51602 (n30505, n30492, n_21193);
  and g51603 (n30506, n_21192, n_21193);
  not g51604 (n_21194, n30505);
  not g51605 (n_21195, n30506);
  and g51606 (n30507, n_21194, n_21195);
  and g51607 (n30508, n_21068, n_21074);
  and g51608 (n30509, n30507, n30508);
  not g51609 (n_21196, n30507);
  not g51610 (n_21197, n30508);
  and g51611 (n30510, n_21196, n_21197);
  not g51612 (n_21198, n30509);
  not g51613 (n_21199, n30510);
  and g51614 (n30511, n_21198, n_21199);
  and g51615 (n30512, n4694, n22309);
  and g51616 (n30513, n4533, n22312);
  and g51617 (n30514, n4604, n22315);
  and g51623 (n30517, n4536, n_14657);
  not g51626 (n_21204, n30518);
  and g51627 (n30519, \a[23] , n_21204);
  not g51628 (n_21205, n30519);
  and g51629 (n30520, \a[23] , n_21205);
  and g51630 (n30521, n_21204, n_21205);
  not g51631 (n_21206, n30520);
  not g51632 (n_21207, n30521);
  and g51633 (n30522, n_21206, n_21207);
  not g51634 (n_21208, n30522);
  and g51635 (n30523, n30511, n_21208);
  not g51636 (n_21209, n30523);
  and g51637 (n30524, n30511, n_21209);
  and g51638 (n30525, n_21208, n_21209);
  not g51639 (n_21210, n30524);
  not g51640 (n_21211, n30525);
  and g51641 (n30526, n_21210, n_21211);
  and g51642 (n30527, n_21084, n_21090);
  and g51643 (n30528, n30526, n30527);
  not g51644 (n_21212, n30526);
  not g51645 (n_21213, n30527);
  and g51646 (n30529, n_21212, n_21213);
  not g51647 (n_21214, n30528);
  not g51648 (n_21215, n30529);
  and g51649 (n30530, n_21214, n_21215);
  and g51650 (n30531, n5496, n26060);
  and g51651 (n30532, n4935, n26063);
  and g51652 (n30533, n5407, n26066);
  and g51658 (n30536, n4938, n_18596);
  not g51661 (n_21220, n30537);
  and g51662 (n30538, \a[20] , n_21220);
  not g51663 (n_21221, n30538);
  and g51664 (n30539, \a[20] , n_21221);
  and g51665 (n30540, n_21220, n_21221);
  not g51666 (n_21222, n30539);
  not g51667 (n_21223, n30540);
  and g51668 (n30541, n_21222, n_21223);
  not g51669 (n_21224, n30541);
  and g51670 (n30542, n30530, n_21224);
  not g51671 (n_21225, n30542);
  and g51672 (n30543, n30530, n_21225);
  and g51673 (n30544, n_21224, n_21225);
  not g51674 (n_21226, n30543);
  not g51675 (n_21227, n30544);
  and g51676 (n30545, n_21226, n_21227);
  and g51677 (n30546, n_21101, n_21107);
  not g51678 (n_21228, n30545);
  not g51679 (n_21229, n30546);
  and g51680 (n30547, n_21228, n_21229);
  not g51681 (n_21230, n30547);
  and g51682 (n30548, n_21228, n_21230);
  and g51683 (n30549, n_21229, n_21230);
  not g51684 (n_21231, n30548);
  not g51685 (n_21232, n30549);
  and g51686 (n30550, n_21231, n_21232);
  and g51687 (n30551, n6233, n27442);
  and g51688 (n30552, n5663, n26890);
  and g51689 (n30553, n5939, n27173);
  and g51695 (n30556, n5666, n27455);
  not g51698 (n_21237, n30557);
  and g51699 (n30558, \a[17] , n_21237);
  not g51700 (n_21238, n30558);
  and g51701 (n30559, \a[17] , n_21238);
  and g51702 (n30560, n_21237, n_21238);
  not g51703 (n_21239, n30559);
  not g51704 (n_21240, n30560);
  and g51705 (n30561, n_21239, n_21240);
  not g51706 (n_21241, n30550);
  not g51707 (n_21242, n30561);
  and g51708 (n30562, n_21241, n_21242);
  not g51709 (n_21243, n30562);
  and g51710 (n30563, n_21241, n_21243);
  and g51711 (n30564, n_21242, n_21243);
  not g51712 (n_21244, n30563);
  not g51713 (n_21245, n30564);
  and g51714 (n30565, n_21244, n_21245);
  and g51715 (n30566, n_21117, n_21123);
  and g51716 (n30567, n30565, n30566);
  not g51717 (n_21246, n30565);
  not g51718 (n_21247, n30566);
  and g51719 (n30568, n_21246, n_21247);
  not g51720 (n_21248, n30567);
  not g51721 (n_21249, n30568);
  and g51722 (n30569, n_21248, n_21249);
  and g51723 (n30570, n7101, n_19417);
  and g51724 (n30571, n6402, n27698);
  and g51725 (n30572, n6951, n27964);
  and g51731 (n30575, n6397, n_19940);
  not g51734 (n_21254, n30576);
  and g51735 (n30577, \a[14] , n_21254);
  not g51736 (n_21255, n30577);
  and g51737 (n30578, \a[14] , n_21255);
  and g51738 (n30579, n_21254, n_21255);
  not g51739 (n_21256, n30578);
  not g51740 (n_21257, n30579);
  and g51741 (n30580, n_21256, n_21257);
  not g51742 (n_21258, n30580);
  and g51743 (n30581, n30569, n_21258);
  not g51744 (n_21259, n30581);
  and g51745 (n30582, n30569, n_21259);
  and g51746 (n30583, n_21258, n_21259);
  not g51747 (n_21260, n30582);
  not g51748 (n_21261, n30583);
  and g51749 (n30584, n_21260, n_21261);
  and g51750 (n30585, n_21134, n_21140);
  not g51751 (n_21262, n30584);
  not g51752 (n_21263, n30585);
  and g51753 (n30586, n_21262, n_21263);
  not g51754 (n_21264, n30586);
  and g51755 (n30587, n_21262, n_21264);
  and g51756 (n30588, n_21263, n_21264);
  not g51757 (n_21265, n30587);
  not g51758 (n_21266, n30588);
  and g51759 (n30589, n_21265, n_21266);
  and g51760 (n30590, n_21143, n_21147);
  and g51761 (n30591, n30589, n30590);
  not g51762 (n_21267, n30589);
  not g51763 (n_21268, n30590);
  and g51764 (n30592, n_21267, n_21268);
  not g51765 (n_21269, n30591);
  not g51766 (n_21270, n30592);
  and g51767 (n30593, n_21269, n_21270);
  and g51768 (n30594, n_21151, n30593);
  not g51769 (n_21271, n30593);
  and g51770 (n30595, n30439, n_21271);
  or g51771 (\result[17] , n30594, n30595);
  and g51772 (n30597, n30439, n30593);
  and g51773 (n30598, n75, n_16015);
  and g51774 (n30599, n3020, n22335);
  and g51775 (n30600, n3023, n22341);
  and g51776 (n30601, n3028, n22338);
  and g51801 (n30622, n_21157, n30621);
  not g51802 (n_21276, n30621);
  and g51803 (n30623, n30464, n_21276);
  not g51804 (n_21277, n30604);
  not g51805 (n_21278, n30623);
  and g51806 (n30624, n_21277, n_21278);
  not g51807 (n_21279, n30622);
  and g51808 (n30625, n_21279, n30624);
  not g51809 (n_21280, n30625);
  and g51810 (n30626, n_21277, n_21280);
  and g51811 (n30627, n_21278, n_21280);
  and g51812 (n30628, n_21279, n30627);
  not g51813 (n_21281, n30626);
  not g51814 (n_21282, n30628);
  and g51815 (n30629, n_21281, n_21282);
  and g51816 (n30630, n_21158, n_21161);
  and g51817 (n30631, n30629, n30630);
  not g51818 (n_21283, n30629);
  not g51819 (n_21284, n30630);
  and g51820 (n30632, n_21283, n_21284);
  not g51821 (n_21285, n30631);
  not g51822 (n_21286, n30632);
  and g51823 (n30633, n_21285, n_21286);
  and g51824 (n30634, n_21167, n_21178);
  not g51825 (n_21287, n30633);
  and g51826 (n30635, n_21287, n30634);
  not g51827 (n_21288, n30634);
  and g51828 (n30636, n30633, n_21288);
  not g51829 (n_21289, n30635);
  not g51830 (n_21290, n30636);
  and g51831 (n30637, n_21289, n_21290);
  and g51832 (n30638, n3457, n22326);
  and g51833 (n30639, n3542, n22332);
  and g51834 (n30640, n3606, n22329);
  and g51840 (n30643, n3368, n_18133);
  not g51843 (n_21295, n30644);
  and g51844 (n30645, \a[29] , n_21295);
  not g51845 (n_21296, n30645);
  and g51846 (n30646, \a[29] , n_21296);
  and g51847 (n30647, n_21295, n_21296);
  not g51848 (n_21297, n30646);
  not g51849 (n_21298, n30647);
  and g51850 (n30648, n_21297, n_21298);
  not g51851 (n_21299, n30648);
  and g51852 (n30649, n30637, n_21299);
  not g51853 (n_21300, n30649);
  and g51854 (n30650, n30637, n_21300);
  and g51855 (n30651, n_21299, n_21300);
  not g51856 (n_21301, n30650);
  not g51857 (n_21302, n30651);
  and g51858 (n30652, n_21301, n_21302);
  and g51859 (n30653, n3884, n22312);
  and g51860 (n30654, n3967, n22323);
  and g51861 (n30655, n4046, n22320);
  and g51867 (n30658, n4050, n_17004);
  not g51870 (n_21307, n30659);
  and g51871 (n30660, \a[26] , n_21307);
  not g51872 (n_21308, n30660);
  and g51873 (n30661, \a[26] , n_21308);
  and g51874 (n30662, n_21307, n_21308);
  not g51875 (n_21309, n30661);
  not g51876 (n_21310, n30662);
  and g51877 (n30663, n_21309, n_21310);
  not g51878 (n_21311, n30652);
  not g51879 (n_21312, n30663);
  and g51880 (n30664, n_21311, n_21312);
  not g51881 (n_21313, n30664);
  and g51882 (n30665, n_21311, n_21313);
  and g51883 (n30666, n_21312, n_21313);
  not g51884 (n_21314, n30665);
  not g51885 (n_21315, n30666);
  and g51886 (n30667, n_21314, n_21315);
  and g51887 (n30668, n_21182, n_21193);
  and g51888 (n30669, n30667, n30668);
  not g51889 (n_21316, n30667);
  not g51890 (n_21317, n30668);
  and g51891 (n30670, n_21316, n_21317);
  not g51892 (n_21318, n30669);
  not g51893 (n_21319, n30670);
  and g51894 (n30671, n_21318, n_21319);
  and g51895 (n30672, n4694, n26063);
  and g51896 (n30673, n4533, n22315);
  and g51897 (n30674, n4604, n22309);
  and g51903 (n30677, n4536, n_18124);
  not g51906 (n_21324, n30678);
  and g51907 (n30679, \a[23] , n_21324);
  not g51908 (n_21325, n30679);
  and g51909 (n30680, \a[23] , n_21325);
  and g51910 (n30681, n_21324, n_21325);
  not g51911 (n_21326, n30680);
  not g51912 (n_21327, n30681);
  and g51913 (n30682, n_21326, n_21327);
  not g51914 (n_21328, n30682);
  and g51915 (n30683, n30671, n_21328);
  not g51916 (n_21329, n30683);
  and g51917 (n30684, n30671, n_21329);
  and g51918 (n30685, n_21328, n_21329);
  not g51919 (n_21330, n30684);
  not g51920 (n_21331, n30685);
  and g51921 (n30686, n_21330, n_21331);
  and g51922 (n30687, n_21199, n_21209);
  and g51923 (n30688, n30686, n30687);
  not g51924 (n_21332, n30686);
  not g51925 (n_21333, n30687);
  and g51926 (n30689, n_21332, n_21333);
  not g51927 (n_21334, n30688);
  not g51928 (n_21335, n30689);
  and g51929 (n30690, n_21334, n_21335);
  and g51930 (n30691, n5496, n26890);
  and g51931 (n30692, n4935, n26066);
  and g51932 (n30693, n5407, n26060);
  and g51938 (n30696, n4938, n_18823);
  not g51941 (n_21340, n30697);
  and g51942 (n30698, \a[20] , n_21340);
  not g51943 (n_21341, n30698);
  and g51944 (n30699, \a[20] , n_21341);
  and g51945 (n30700, n_21340, n_21341);
  not g51946 (n_21342, n30699);
  not g51947 (n_21343, n30700);
  and g51948 (n30701, n_21342, n_21343);
  not g51949 (n_21344, n30701);
  and g51950 (n30702, n30690, n_21344);
  not g51951 (n_21345, n30702);
  and g51952 (n30703, n30690, n_21345);
  and g51953 (n30704, n_21344, n_21345);
  not g51954 (n_21346, n30703);
  not g51955 (n_21347, n30704);
  and g51956 (n30705, n_21346, n_21347);
  and g51957 (n30706, n_21215, n_21225);
  and g51958 (n30707, n30705, n30706);
  not g51959 (n_21348, n30705);
  not g51960 (n_21349, n30706);
  and g51961 (n30708, n_21348, n_21349);
  not g51962 (n_21350, n30707);
  not g51963 (n_21351, n30708);
  and g51964 (n30709, n_21350, n_21351);
  and g51965 (n30710, n6233, n27698);
  and g51966 (n30711, n5663, n27173);
  and g51967 (n30712, n5939, n27442);
  and g51973 (n30715, n5666, n_19446);
  not g51976 (n_21356, n30716);
  and g51977 (n30717, \a[17] , n_21356);
  not g51978 (n_21357, n30717);
  and g51979 (n30718, \a[17] , n_21357);
  and g51980 (n30719, n_21356, n_21357);
  not g51981 (n_21358, n30718);
  not g51982 (n_21359, n30719);
  and g51983 (n30720, n_21358, n_21359);
  not g51984 (n_21360, n30720);
  and g51985 (n30721, n30709, n_21360);
  not g51986 (n_21361, n30721);
  and g51987 (n30722, n30709, n_21361);
  and g51988 (n30723, n_21360, n_21361);
  not g51989 (n_21362, n30722);
  not g51990 (n_21363, n30723);
  and g51991 (n30724, n_21362, n_21363);
  and g51992 (n30725, n_21230, n_21243);
  and g51993 (n30726, n_8877, n_19417);
  and g51994 (n30727, n6402, n27964);
  not g51995 (n_21364, n30726);
  not g51996 (n_21365, n30727);
  and g51997 (n30728, n_21364, n_21365);
  and g51998 (n30729, n_1885, n30728);
  and g51999 (n30730, n28221, n30728);
  not g52000 (n_21366, n30729);
  not g52001 (n_21367, n30730);
  and g52002 (n30731, n_21366, n_21367);
  not g52003 (n_21368, n30731);
  and g52004 (n30732, \a[14] , n_21368);
  and g52005 (n30733, n_652, n30731);
  not g52006 (n_21369, n30732);
  not g52007 (n_21370, n30733);
  and g52008 (n30734, n_21369, n_21370);
  not g52009 (n_21371, n30725);
  not g52010 (n_21372, n30734);
  and g52011 (n30735, n_21371, n_21372);
  and g52012 (n30736, n30725, n30734);
  not g52013 (n_21373, n30735);
  not g52014 (n_21374, n30736);
  and g52015 (n30737, n_21373, n_21374);
  not g52016 (n_21375, n30724);
  and g52017 (n30738, n_21375, n30737);
  not g52018 (n_21376, n30738);
  and g52019 (n30739, n_21375, n_21376);
  and g52020 (n30740, n30737, n_21376);
  not g52021 (n_21377, n30739);
  not g52022 (n_21378, n30740);
  and g52023 (n30741, n_21377, n_21378);
  and g52024 (n30742, n_21249, n_21259);
  and g52025 (n30743, n30741, n30742);
  not g52026 (n_21379, n30741);
  not g52027 (n_21380, n30742);
  and g52028 (n30744, n_21379, n_21380);
  not g52029 (n_21381, n30743);
  not g52030 (n_21382, n30744);
  and g52031 (n30745, n_21381, n_21382);
  and g52032 (n30746, n_21264, n_21270);
  not g52033 (n_21383, n30745);
  and g52034 (n30747, n_21383, n30746);
  not g52035 (n_21384, n30746);
  and g52036 (n30748, n30745, n_21384);
  not g52037 (n_21385, n30747);
  not g52038 (n_21386, n30748);
  and g52039 (n30749, n_21385, n_21386);
  and g52040 (n30750, n30597, n30749);
  not g52041 (n_21387, n30597);
  not g52042 (n_21388, n30749);
  and g52043 (n30751, n_21387, n_21388);
  not g52044 (n_21389, n30750);
  not g52045 (n_21390, n30751);
  and g52046 (\result[18] , n_21389, n_21390);
  and g52047 (n30753, n_21382, n_21386);
  and g52048 (n30754, n_21373, n_21376);
  and g52049 (n30755, n75, n22542);
  and g52050 (n30756, n3020, n22332);
  and g52051 (n30757, n3023, n22338);
  and g52052 (n30758, n3028, n22335);
  and g52060 (n30762, n_7622, n_19417);
  not g52061 (n_21395, n30762);
  and g52062 (n30763, \a[14] , n_21395);
  and g52063 (n30764, n_652, n30762);
  not g52064 (n_21396, n30763);
  not g52065 (n_21397, n30764);
  and g52066 (n30765, n_21396, n_21397);
  and g52079 (n30778, n30464, n30777);
  not g52080 (n_21398, n30777);
  and g52081 (n30779, n_21157, n_21398);
  not g52082 (n_21399, n30778);
  not g52083 (n_21400, n30779);
  and g52084 (n30780, n_21399, n_21400);
  and g52085 (n30781, n30765, n30780);
  not g52086 (n_21401, n30765);
  not g52087 (n_21402, n30780);
  and g52088 (n30782, n_21401, n_21402);
  not g52089 (n_21403, n30781);
  not g52090 (n_21404, n30782);
  and g52091 (n30783, n_21403, n_21404);
  not g52092 (n_21405, n30627);
  and g52093 (n30784, n_21405, n30783);
  not g52094 (n_21406, n30783);
  and g52095 (n30785, n30627, n_21406);
  not g52096 (n_21407, n30784);
  not g52097 (n_21408, n30785);
  and g52098 (n30786, n_21407, n_21408);
  not g52099 (n_21409, n30761);
  and g52100 (n30787, n_21409, n30786);
  not g52101 (n_21410, n30787);
  and g52102 (n30788, n30786, n_21410);
  and g52103 (n30789, n_21409, n_21410);
  not g52104 (n_21411, n30788);
  not g52105 (n_21412, n30789);
  and g52106 (n30790, n_21411, n_21412);
  and g52107 (n30791, n3457, n22323);
  and g52108 (n30792, n3542, n22329);
  and g52109 (n30793, n3606, n22326);
  and g52115 (n30796, n3368, n24599);
  not g52118 (n_21417, n30797);
  and g52119 (n30798, \a[29] , n_21417);
  not g52120 (n_21418, n30798);
  and g52121 (n30799, \a[29] , n_21418);
  and g52122 (n30800, n_21417, n_21418);
  not g52123 (n_21419, n30799);
  not g52124 (n_21420, n30800);
  and g52125 (n30801, n_21419, n_21420);
  not g52126 (n_21421, n30790);
  not g52127 (n_21422, n30801);
  and g52128 (n30802, n_21421, n_21422);
  not g52129 (n_21423, n30802);
  and g52130 (n30803, n_21421, n_21423);
  and g52131 (n30804, n_21422, n_21423);
  not g52132 (n_21424, n30803);
  not g52133 (n_21425, n30804);
  and g52134 (n30805, n_21424, n_21425);
  and g52135 (n30806, n_21286, n_21290);
  and g52136 (n30807, n30805, n30806);
  not g52137 (n_21426, n30805);
  not g52138 (n_21427, n30806);
  and g52139 (n30808, n_21426, n_21427);
  not g52140 (n_21428, n30807);
  not g52141 (n_21429, n30808);
  and g52142 (n30809, n_21428, n_21429);
  and g52143 (n30810, n3884, n22315);
  and g52144 (n30811, n3967, n22320);
  and g52145 (n30812, n4046, n22312);
  and g52151 (n30815, n4050, n25294);
  not g52154 (n_21434, n30816);
  and g52155 (n30817, \a[26] , n_21434);
  not g52156 (n_21435, n30817);
  and g52157 (n30818, \a[26] , n_21435);
  and g52158 (n30819, n_21434, n_21435);
  not g52159 (n_21436, n30818);
  not g52160 (n_21437, n30819);
  and g52161 (n30820, n_21436, n_21437);
  not g52162 (n_21438, n30820);
  and g52163 (n30821, n30809, n_21438);
  not g52164 (n_21439, n30821);
  and g52165 (n30822, n30809, n_21439);
  and g52166 (n30823, n_21438, n_21439);
  not g52167 (n_21440, n30822);
  not g52168 (n_21441, n30823);
  and g52169 (n30824, n_21440, n_21441);
  and g52170 (n30825, n_21300, n_21313);
  and g52171 (n30826, n30824, n30825);
  not g52172 (n_21442, n30824);
  not g52173 (n_21443, n30825);
  and g52174 (n30827, n_21442, n_21443);
  not g52175 (n_21444, n30826);
  not g52176 (n_21445, n30827);
  and g52177 (n30828, n_21444, n_21445);
  and g52178 (n30829, n_21319, n_21329);
  and g52179 (n30830, n4694, n26066);
  and g52180 (n30831, n4533, n22309);
  and g52181 (n30832, n4604, n26063);
  and g52187 (n30835, n4536, n_18359);
  not g52190 (n_21450, n30836);
  and g52191 (n30837, \a[23] , n_21450);
  not g52192 (n_21451, n30837);
  and g52193 (n30838, \a[23] , n_21451);
  and g52194 (n30839, n_21450, n_21451);
  not g52195 (n_21452, n30838);
  not g52196 (n_21453, n30839);
  and g52197 (n30840, n_21452, n_21453);
  not g52198 (n_21454, n30829);
  not g52199 (n_21455, n30840);
  and g52200 (n30841, n_21454, n_21455);
  not g52201 (n_21456, n30841);
  and g52202 (n30842, n_21454, n_21456);
  and g52203 (n30843, n_21455, n_21456);
  not g52204 (n_21457, n30842);
  not g52205 (n_21458, n30843);
  and g52206 (n30844, n_21457, n_21458);
  not g52207 (n_21459, n30828);
  and g52208 (n30845, n_21459, n30844);
  not g52209 (n_21460, n30844);
  and g52210 (n30846, n30828, n_21460);
  not g52211 (n_21461, n30845);
  not g52212 (n_21462, n30846);
  and g52213 (n30847, n_21461, n_21462);
  and g52214 (n30848, n5496, n27173);
  and g52215 (n30849, n4935, n26060);
  and g52216 (n30850, n5407, n26890);
  and g52222 (n30853, n4938, n27185);
  not g52225 (n_21467, n30854);
  and g52226 (n30855, \a[20] , n_21467);
  not g52227 (n_21468, n30855);
  and g52228 (n30856, \a[20] , n_21468);
  and g52229 (n30857, n_21467, n_21468);
  not g52230 (n_21469, n30856);
  not g52231 (n_21470, n30857);
  and g52232 (n30858, n_21469, n_21470);
  not g52233 (n_21471, n30858);
  and g52234 (n30859, n30847, n_21471);
  not g52235 (n_21472, n30859);
  and g52236 (n30860, n30847, n_21472);
  and g52237 (n30861, n_21471, n_21472);
  not g52238 (n_21473, n30860);
  not g52239 (n_21474, n30861);
  and g52240 (n30862, n_21473, n_21474);
  and g52241 (n30863, n_21335, n_21345);
  and g52242 (n30864, n30862, n30863);
  not g52243 (n_21475, n30862);
  not g52244 (n_21476, n30863);
  and g52245 (n30865, n_21475, n_21476);
  not g52246 (n_21477, n30864);
  not g52247 (n_21478, n30865);
  and g52248 (n30866, n_21477, n_21478);
  and g52249 (n30867, n_21351, n_21361);
  and g52250 (n30868, n6233, n27964);
  and g52251 (n30869, n5663, n27442);
  and g52252 (n30870, n5939, n27698);
  and g52258 (n30873, n5666, n27976);
  not g52261 (n_21483, n30874);
  and g52262 (n30875, \a[17] , n_21483);
  not g52263 (n_21484, n30875);
  and g52264 (n30876, \a[17] , n_21484);
  and g52265 (n30877, n_21483, n_21484);
  not g52266 (n_21485, n30876);
  not g52267 (n_21486, n30877);
  and g52268 (n30878, n_21485, n_21486);
  not g52269 (n_21487, n30867);
  not g52270 (n_21488, n30878);
  and g52271 (n30879, n_21487, n_21488);
  not g52272 (n_21489, n30879);
  and g52273 (n30880, n_21487, n_21489);
  and g52274 (n30881, n_21488, n_21489);
  not g52275 (n_21490, n30880);
  not g52276 (n_21491, n30881);
  and g52277 (n30882, n_21490, n_21491);
  not g52278 (n_21492, n30866);
  and g52279 (n30883, n_21492, n30882);
  not g52280 (n_21493, n30882);
  and g52281 (n30884, n30866, n_21493);
  not g52282 (n_21494, n30883);
  not g52283 (n_21495, n30884);
  and g52284 (n30885, n_21494, n_21495);
  not g52285 (n_21496, n30754);
  and g52286 (n30886, n_21496, n30885);
  not g52287 (n_21497, n30885);
  and g52288 (n30887, n30754, n_21497);
  not g52289 (n_21498, n30886);
  not g52290 (n_21499, n30887);
  and g52291 (n30888, n_21498, n_21499);
  not g52292 (n_21500, n30753);
  and g52293 (n30889, n_21500, n30888);
  not g52294 (n_21501, n30888);
  and g52295 (n30890, n30753, n_21501);
  not g52296 (n_21502, n30889);
  not g52297 (n_21503, n30890);
  and g52298 (n30891, n_21502, n_21503);
  not g52299 (n_21504, n30891);
  and g52300 (n30892, n_21389, n_21504);
  and g52301 (n30893, n30750, n30891);
  not g52302 (n_21505, n30892);
  not g52303 (n_21506, n30893);
  and g52304 (\result[19] , n_21505, n_21506);
  and g52305 (n30895, n_21423, n_21429);
  and g52306 (n30896, n75, n_16827);
  and g52307 (n30897, n3020, n22329);
  and g52308 (n30898, n3023, n22335);
  and g52309 (n30899, n3028, n22332);
  and g52317 (n30903, n_21400, n_21403);
  not g52334 (n_21511, n30903);
  and g52335 (n30920, n_21511, n30919);
  not g52336 (n_21512, n30919);
  and g52337 (n30921, n30903, n_21512);
  not g52338 (n_21513, n30920);
  not g52339 (n_21514, n30921);
  and g52340 (n30922, n_21513, n_21514);
  not g52341 (n_21515, n30902);
  and g52342 (n30923, n_21515, n30922);
  not g52343 (n_21516, n30923);
  and g52344 (n30924, n_21515, n_21516);
  and g52345 (n30925, n30922, n_21516);
  not g52346 (n_21517, n30924);
  not g52347 (n_21518, n30925);
  and g52348 (n30926, n_21517, n_21518);
  and g52349 (n30927, n_21407, n_21410);
  and g52350 (n30928, n30926, n30927);
  not g52351 (n_21519, n30926);
  not g52352 (n_21520, n30927);
  and g52353 (n30929, n_21519, n_21520);
  not g52354 (n_21521, n30928);
  not g52355 (n_21522, n30929);
  and g52356 (n30930, n_21521, n_21522);
  and g52357 (n30931, n3457, n22320);
  and g52358 (n30932, n3542, n22326);
  and g52359 (n30933, n3606, n22323);
  not g52360 (n_21523, n30932);
  not g52361 (n_21524, n30933);
  and g52362 (n30934, n_21523, n_21524);
  not g52363 (n_21525, n30931);
  and g52364 (n30935, n_21525, n30934);
  and g52365 (n30936, n_489, n30935);
  and g52366 (n30937, n25270, n30935);
  not g52367 (n_21526, n30936);
  not g52368 (n_21527, n30937);
  and g52369 (n30938, n_21526, n_21527);
  not g52370 (n_21528, n30938);
  and g52371 (n30939, \a[29] , n_21528);
  and g52372 (n30940, n_15, n30938);
  not g52373 (n_21529, n30939);
  not g52374 (n_21530, n30940);
  and g52375 (n30941, n_21529, n_21530);
  not g52376 (n_21531, n30941);
  and g52377 (n30942, n30930, n_21531);
  not g52378 (n_21532, n30930);
  and g52379 (n30943, n_21532, n30941);
  not g52380 (n_21533, n30942);
  not g52381 (n_21534, n30943);
  and g52382 (n30944, n_21533, n_21534);
  not g52383 (n_21535, n30895);
  and g52384 (n30945, n_21535, n30944);
  not g52385 (n_21536, n30944);
  and g52386 (n30946, n30895, n_21536);
  not g52387 (n_21537, n30945);
  not g52388 (n_21538, n30946);
  and g52389 (n30947, n_21537, n_21538);
  and g52390 (n30948, n3884, n22309);
  and g52391 (n30949, n3967, n22312);
  and g52392 (n30950, n4046, n22315);
  and g52398 (n30953, n4050, n_14657);
  not g52401 (n_21543, n30954);
  and g52402 (n30955, \a[26] , n_21543);
  not g52403 (n_21544, n30955);
  and g52404 (n30956, \a[26] , n_21544);
  and g52405 (n30957, n_21543, n_21544);
  not g52406 (n_21545, n30956);
  not g52407 (n_21546, n30957);
  and g52408 (n30958, n_21545, n_21546);
  not g52409 (n_21547, n30958);
  and g52410 (n30959, n30947, n_21547);
  not g52411 (n_21548, n30959);
  and g52412 (n30960, n30947, n_21548);
  and g52413 (n30961, n_21547, n_21548);
  not g52414 (n_21549, n30960);
  not g52415 (n_21550, n30961);
  and g52416 (n30962, n_21549, n_21550);
  and g52417 (n30963, n_21439, n_21445);
  and g52418 (n30964, n30962, n30963);
  not g52419 (n_21551, n30962);
  not g52420 (n_21552, n30963);
  and g52421 (n30965, n_21551, n_21552);
  not g52422 (n_21553, n30964);
  not g52423 (n_21554, n30965);
  and g52424 (n30966, n_21553, n_21554);
  and g52425 (n30967, n4694, n26060);
  and g52426 (n30968, n4533, n26063);
  and g52427 (n30969, n4604, n26066);
  and g52433 (n30972, n4536, n_18596);
  not g52436 (n_21559, n30973);
  and g52437 (n30974, \a[23] , n_21559);
  not g52438 (n_21560, n30974);
  and g52439 (n30975, \a[23] , n_21560);
  and g52440 (n30976, n_21559, n_21560);
  not g52441 (n_21561, n30975);
  not g52442 (n_21562, n30976);
  and g52443 (n30977, n_21561, n_21562);
  not g52444 (n_21563, n30977);
  and g52445 (n30978, n30966, n_21563);
  not g52446 (n_21564, n30978);
  and g52447 (n30979, n30966, n_21564);
  and g52448 (n30980, n_21563, n_21564);
  not g52449 (n_21565, n30979);
  not g52450 (n_21566, n30980);
  and g52451 (n30981, n_21565, n_21566);
  and g52452 (n30982, n_21456, n_21462);
  not g52453 (n_21567, n30981);
  not g52454 (n_21568, n30982);
  and g52455 (n30983, n_21567, n_21568);
  not g52456 (n_21569, n30983);
  and g52457 (n30984, n_21567, n_21569);
  and g52458 (n30985, n_21568, n_21569);
  not g52459 (n_21570, n30984);
  not g52460 (n_21571, n30985);
  and g52461 (n30986, n_21570, n_21571);
  and g52462 (n30987, n5496, n27442);
  and g52463 (n30988, n4935, n26890);
  and g52464 (n30989, n5407, n27173);
  and g52470 (n30992, n4938, n27455);
  not g52473 (n_21576, n30993);
  and g52474 (n30994, \a[20] , n_21576);
  not g52475 (n_21577, n30994);
  and g52476 (n30995, \a[20] , n_21577);
  and g52477 (n30996, n_21576, n_21577);
  not g52478 (n_21578, n30995);
  not g52479 (n_21579, n30996);
  and g52480 (n30997, n_21578, n_21579);
  not g52481 (n_21580, n30986);
  not g52482 (n_21581, n30997);
  and g52483 (n30998, n_21580, n_21581);
  not g52484 (n_21582, n30998);
  and g52485 (n30999, n_21580, n_21582);
  and g52486 (n31000, n_21581, n_21582);
  not g52487 (n_21583, n30999);
  not g52488 (n_21584, n31000);
  and g52489 (n31001, n_21583, n_21584);
  and g52490 (n31002, n_21472, n_21478);
  and g52491 (n31003, n31001, n31002);
  not g52492 (n_21585, n31001);
  not g52493 (n_21586, n31002);
  and g52494 (n31004, n_21585, n_21586);
  not g52495 (n_21587, n31003);
  not g52496 (n_21588, n31004);
  and g52497 (n31005, n_21587, n_21588);
  and g52498 (n31006, n6233, n_19417);
  and g52499 (n31007, n5663, n27698);
  and g52500 (n31008, n5939, n27964);
  and g52506 (n31011, n5666, n_19940);
  not g52509 (n_21593, n31012);
  and g52510 (n31013, \a[17] , n_21593);
  not g52511 (n_21594, n31013);
  and g52512 (n31014, \a[17] , n_21594);
  and g52513 (n31015, n_21593, n_21594);
  not g52514 (n_21595, n31014);
  not g52515 (n_21596, n31015);
  and g52516 (n31016, n_21595, n_21596);
  not g52517 (n_21597, n31016);
  and g52518 (n31017, n31005, n_21597);
  not g52519 (n_21598, n31017);
  and g52520 (n31018, n31005, n_21598);
  and g52521 (n31019, n_21597, n_21598);
  not g52522 (n_21599, n31018);
  not g52523 (n_21600, n31019);
  and g52524 (n31020, n_21599, n_21600);
  and g52525 (n31021, n_21489, n_21495);
  not g52526 (n_21601, n31020);
  not g52527 (n_21602, n31021);
  and g52528 (n31022, n_21601, n_21602);
  not g52529 (n_21603, n31022);
  and g52530 (n31023, n_21601, n_21603);
  and g52531 (n31024, n_21602, n_21603);
  not g52532 (n_21604, n31023);
  not g52533 (n_21605, n31024);
  and g52534 (n31025, n_21604, n_21605);
  and g52535 (n31026, n_21498, n_21502);
  and g52536 (n31027, n31025, n31026);
  not g52537 (n_21606, n31025);
  not g52538 (n_21607, n31026);
  and g52539 (n31028, n_21606, n_21607);
  not g52540 (n_21608, n31027);
  not g52541 (n_21609, n31028);
  and g52542 (n31029, n_21608, n_21609);
  not g52543 (n_21610, n31029);
  and g52544 (n31030, n30893, n_21610);
  and g52545 (n31031, n_21506, n31029);
  or g52546 (\result[20] , n31030, n31031);
  and g52547 (n31033, n_21522, n_21533);
  and g52548 (n31034, n_21513, n_21516);
  and g52549 (n31035, n_97, n1253);
  and g52550 (n31036, n_46, n31035);
  not g52567 (n_21611, n31052);
  and g52568 (n31053, n30919, n_21611);
  and g52569 (n31054, n_21512, n31052);
  not g52570 (n_21612, n31034);
  not g52571 (n_21613, n31054);
  and g52572 (n31055, n_21612, n_21613);
  not g52573 (n_21614, n31053);
  and g52574 (n31056, n_21614, n31055);
  not g52575 (n_21615, n31056);
  and g52576 (n31057, n_21612, n_21615);
  and g52577 (n31058, n_21613, n_21615);
  and g52578 (n31059, n_21614, n31058);
  not g52579 (n_21616, n31057);
  not g52580 (n_21617, n31059);
  and g52581 (n31060, n_21616, n_21617);
  and g52582 (n31061, n75, n_18133);
  and g52583 (n31062, n3020, n22326);
  and g52584 (n31063, n3023, n22332);
  and g52585 (n31064, n3028, n22329);
  not g52593 (n_21622, n31060);
  not g52594 (n_21623, n31067);
  and g52595 (n31068, n_21622, n_21623);
  not g52596 (n_21624, n31068);
  and g52597 (n31069, n_21622, n_21624);
  and g52598 (n31070, n_21623, n_21624);
  not g52599 (n_21625, n31069);
  not g52600 (n_21626, n31070);
  and g52601 (n31071, n_21625, n_21626);
  and g52602 (n31072, n3457, n22312);
  and g52603 (n31073, n3542, n22323);
  and g52604 (n31074, n3606, n22320);
  not g52605 (n_21627, n31073);
  not g52606 (n_21628, n31074);
  and g52607 (n31075, n_21627, n_21628);
  not g52608 (n_21629, n31072);
  and g52609 (n31076, n_21629, n31075);
  and g52610 (n31077, n_489, n31076);
  and g52611 (n31078, n25315, n31076);
  not g52612 (n_21630, n31077);
  not g52613 (n_21631, n31078);
  and g52614 (n31079, n_21630, n_21631);
  not g52615 (n_21632, n31079);
  and g52616 (n31080, \a[29] , n_21632);
  and g52617 (n31081, n_15, n31079);
  not g52618 (n_21633, n31080);
  not g52619 (n_21634, n31081);
  and g52620 (n31082, n_21633, n_21634);
  not g52621 (n_21635, n31071);
  not g52622 (n_21636, n31082);
  and g52623 (n31083, n_21635, n_21636);
  and g52624 (n31084, n31071, n31082);
  not g52625 (n_21637, n31083);
  not g52626 (n_21638, n31084);
  and g52627 (n31085, n_21637, n_21638);
  not g52628 (n_21639, n31033);
  and g52629 (n31086, n_21639, n31085);
  not g52630 (n_21640, n31085);
  and g52631 (n31087, n31033, n_21640);
  not g52632 (n_21641, n31086);
  not g52633 (n_21642, n31087);
  and g52634 (n31088, n_21641, n_21642);
  and g52635 (n31089, n3884, n26063);
  and g52636 (n31090, n3967, n22315);
  and g52637 (n31091, n4046, n22309);
  and g52643 (n31094, n4050, n_18124);
  not g52646 (n_21647, n31095);
  and g52647 (n31096, \a[26] , n_21647);
  not g52648 (n_21648, n31096);
  and g52649 (n31097, \a[26] , n_21648);
  and g52650 (n31098, n_21647, n_21648);
  not g52651 (n_21649, n31097);
  not g52652 (n_21650, n31098);
  and g52653 (n31099, n_21649, n_21650);
  not g52654 (n_21651, n31099);
  and g52655 (n31100, n31088, n_21651);
  not g52656 (n_21652, n31100);
  and g52657 (n31101, n31088, n_21652);
  and g52658 (n31102, n_21651, n_21652);
  not g52659 (n_21653, n31101);
  not g52660 (n_21654, n31102);
  and g52661 (n31103, n_21653, n_21654);
  and g52662 (n31104, n_21537, n_21548);
  and g52663 (n31105, n31103, n31104);
  not g52664 (n_21655, n31103);
  not g52665 (n_21656, n31104);
  and g52666 (n31106, n_21655, n_21656);
  not g52667 (n_21657, n31105);
  not g52668 (n_21658, n31106);
  and g52669 (n31107, n_21657, n_21658);
  and g52670 (n31108, n4694, n26890);
  and g52671 (n31109, n4533, n26066);
  and g52672 (n31110, n4604, n26060);
  and g52678 (n31113, n4536, n_18823);
  not g52681 (n_21663, n31114);
  and g52682 (n31115, \a[23] , n_21663);
  not g52683 (n_21664, n31115);
  and g52684 (n31116, \a[23] , n_21664);
  and g52685 (n31117, n_21663, n_21664);
  not g52686 (n_21665, n31116);
  not g52687 (n_21666, n31117);
  and g52688 (n31118, n_21665, n_21666);
  not g52689 (n_21667, n31118);
  and g52690 (n31119, n31107, n_21667);
  not g52691 (n_21668, n31119);
  and g52692 (n31120, n31107, n_21668);
  and g52693 (n31121, n_21667, n_21668);
  not g52694 (n_21669, n31120);
  not g52695 (n_21670, n31121);
  and g52696 (n31122, n_21669, n_21670);
  and g52697 (n31123, n_21554, n_21564);
  and g52698 (n31124, n31122, n31123);
  not g52699 (n_21671, n31122);
  not g52700 (n_21672, n31123);
  and g52701 (n31125, n_21671, n_21672);
  not g52702 (n_21673, n31124);
  not g52703 (n_21674, n31125);
  and g52704 (n31126, n_21673, n_21674);
  and g52705 (n31127, n5496, n27698);
  and g52706 (n31128, n4935, n27173);
  and g52707 (n31129, n5407, n27442);
  and g52713 (n31132, n4938, n_19446);
  not g52716 (n_21679, n31133);
  and g52717 (n31134, \a[20] , n_21679);
  not g52718 (n_21680, n31134);
  and g52719 (n31135, \a[20] , n_21680);
  and g52720 (n31136, n_21679, n_21680);
  not g52721 (n_21681, n31135);
  not g52722 (n_21682, n31136);
  and g52723 (n31137, n_21681, n_21682);
  not g52724 (n_21683, n31137);
  and g52725 (n31138, n31126, n_21683);
  not g52726 (n_21684, n31138);
  and g52727 (n31139, n31126, n_21684);
  and g52728 (n31140, n_21683, n_21684);
  not g52729 (n_21685, n31139);
  not g52730 (n_21686, n31140);
  and g52731 (n31141, n_21685, n_21686);
  and g52732 (n31142, n_21569, n_21582);
  and g52733 (n31143, n_8391, n_19417);
  and g52734 (n31144, n5663, n27964);
  not g52735 (n_21687, n31143);
  not g52736 (n_21688, n31144);
  and g52737 (n31145, n_21687, n_21688);
  and g52738 (n31146, n_1409, n31145);
  and g52739 (n31147, n28221, n31145);
  not g52740 (n_21689, n31146);
  not g52741 (n_21690, n31147);
  and g52742 (n31148, n_21689, n_21690);
  not g52743 (n_21691, n31148);
  and g52744 (n31149, \a[17] , n_21691);
  and g52745 (n31150, n_617, n31148);
  not g52746 (n_21692, n31149);
  not g52747 (n_21693, n31150);
  and g52748 (n31151, n_21692, n_21693);
  not g52749 (n_21694, n31142);
  not g52750 (n_21695, n31151);
  and g52751 (n31152, n_21694, n_21695);
  and g52752 (n31153, n31142, n31151);
  not g52753 (n_21696, n31152);
  not g52754 (n_21697, n31153);
  and g52755 (n31154, n_21696, n_21697);
  not g52756 (n_21698, n31141);
  and g52757 (n31155, n_21698, n31154);
  not g52758 (n_21699, n31155);
  and g52759 (n31156, n_21698, n_21699);
  and g52760 (n31157, n31154, n_21699);
  not g52761 (n_21700, n31156);
  not g52762 (n_21701, n31157);
  and g52763 (n31158, n_21700, n_21701);
  and g52764 (n31159, n_21588, n_21598);
  and g52765 (n31160, n31158, n31159);
  not g52766 (n_21702, n31158);
  not g52767 (n_21703, n31159);
  and g52768 (n31161, n_21702, n_21703);
  not g52769 (n_21704, n31160);
  not g52770 (n_21705, n31161);
  and g52771 (n31162, n_21704, n_21705);
  and g52772 (n31163, n_21603, n_21609);
  not g52773 (n_21706, n31162);
  and g52774 (n31164, n_21706, n31163);
  not g52775 (n_21707, n31163);
  and g52776 (n31165, n31162, n_21707);
  not g52777 (n_21708, n31164);
  not g52778 (n_21709, n31165);
  and g52779 (n31166, n_21708, n_21709);
  and g52780 (n31167, n30893, n31029);
  and g52781 (n31168, n31166, n31167);
  not g52782 (n_21710, n31166);
  not g52783 (n_21711, n31167);
  and g52784 (n31169, n_21710, n_21711);
  not g52785 (n_21712, n31168);
  not g52786 (n_21713, n31169);
  and g52787 (\result[21] , n_21712, n_21713);
  and g52788 (n31171, n_21705, n_21709);
  and g52789 (n31172, n_21696, n_21699);
  and g52790 (n31173, n_21658, n_21668);
  and g52791 (n31174, n_21641, n_21652);
  and g52792 (n31175, n3884, n26066);
  and g52793 (n31176, n3967, n22309);
  and g52794 (n31177, n4046, n26063);
  and g52800 (n31180, n4050, n_18359);
  not g52803 (n_21718, n31181);
  and g52804 (n31182, \a[26] , n_21718);
  not g52805 (n_21719, n31182);
  and g52806 (n31183, \a[26] , n_21719);
  and g52807 (n31184, n_21718, n_21719);
  not g52808 (n_21720, n31183);
  not g52809 (n_21721, n31184);
  and g52810 (n31185, n_21720, n_21721);
  not g52811 (n_21722, n31174);
  not g52812 (n_21723, n31185);
  and g52813 (n31186, n_21722, n_21723);
  not g52814 (n_21724, n31186);
  and g52815 (n31187, n_21722, n_21724);
  and g52816 (n31188, n_21723, n_21724);
  not g52817 (n_21725, n31187);
  not g52818 (n_21726, n31188);
  and g52819 (n31189, n_21725, n_21726);
  and g52820 (n31190, n_21624, n_21637);
  and g52821 (n31191, n75, n24599);
  and g52822 (n31192, n3020, n22323);
  and g52823 (n31193, n3023, n22329);
  and g52824 (n31194, n3028, n22326);
  and g52832 (n31198, n_7582, n_19417);
  not g52833 (n_21731, n31198);
  and g52834 (n31199, \a[17] , n_21731);
  and g52835 (n31200, n_617, n31198);
  not g52836 (n_21732, n31199);
  not g52837 (n_21733, n31200);
  and g52838 (n31201, n_21732, n_21733);
  and g52852 (n31215, n31052, n31214);
  not g52853 (n_21734, n31214);
  and g52854 (n31216, n_21611, n_21734);
  not g52855 (n_21735, n31215);
  not g52856 (n_21736, n31216);
  and g52857 (n31217, n_21735, n_21736);
  and g52858 (n31218, n31201, n31217);
  not g52859 (n_21737, n31201);
  not g52860 (n_21738, n31217);
  and g52861 (n31219, n_21737, n_21738);
  not g52862 (n_21739, n31218);
  not g52863 (n_21740, n31219);
  and g52864 (n31220, n_21739, n_21740);
  not g52865 (n_21741, n31197);
  and g52866 (n31221, n_21741, n31220);
  not g52867 (n_21742, n31221);
  and g52868 (n31222, n31220, n_21742);
  and g52869 (n31223, n_21741, n_21742);
  not g52870 (n_21743, n31222);
  not g52871 (n_21744, n31223);
  and g52872 (n31224, n_21743, n_21744);
  not g52873 (n_21745, n31058);
  not g52874 (n_21746, n31224);
  and g52875 (n31225, n_21745, n_21746);
  not g52876 (n_21747, n31225);
  and g52877 (n31226, n_21746, n_21747);
  and g52878 (n31227, n_21745, n_21747);
  not g52879 (n_21748, n31226);
  not g52880 (n_21749, n31227);
  and g52881 (n31228, n_21748, n_21749);
  not g52882 (n_21750, n31190);
  not g52883 (n_21751, n31228);
  and g52884 (n31229, n_21750, n_21751);
  not g52885 (n_21752, n31229);
  and g52886 (n31230, n_21750, n_21752);
  and g52887 (n31231, n_21751, n_21752);
  not g52888 (n_21753, n31230);
  not g52889 (n_21754, n31231);
  and g52890 (n31232, n_21753, n_21754);
  and g52891 (n31233, n3457, n22315);
  and g52892 (n31234, n3542, n22320);
  and g52893 (n31235, n3606, n22312);
  and g52899 (n31238, n3368, n25294);
  not g52902 (n_21759, n31239);
  and g52903 (n31240, \a[29] , n_21759);
  not g52904 (n_21760, n31240);
  and g52905 (n31241, \a[29] , n_21760);
  and g52906 (n31242, n_21759, n_21760);
  not g52907 (n_21761, n31241);
  not g52908 (n_21762, n31242);
  and g52909 (n31243, n_21761, n_21762);
  not g52910 (n_21763, n31232);
  not g52911 (n_21764, n31243);
  and g52912 (n31244, n_21763, n_21764);
  not g52913 (n_21765, n31244);
  and g52914 (n31245, n_21763, n_21765);
  and g52915 (n31246, n_21764, n_21765);
  not g52916 (n_21766, n31245);
  not g52917 (n_21767, n31246);
  and g52918 (n31247, n_21766, n_21767);
  not g52919 (n_21768, n31189);
  and g52920 (n31248, n_21768, n31247);
  not g52921 (n_21769, n31247);
  and g52922 (n31249, n31189, n_21769);
  not g52923 (n_21770, n31248);
  not g52924 (n_21771, n31249);
  and g52925 (n31250, n_21770, n_21771);
  and g52926 (n31251, n4694, n27173);
  and g52927 (n31252, n4533, n26060);
  and g52928 (n31253, n4604, n26890);
  and g52934 (n31256, n4536, n27185);
  not g52937 (n_21776, n31257);
  and g52938 (n31258, \a[23] , n_21776);
  not g52939 (n_21777, n31258);
  and g52940 (n31259, \a[23] , n_21777);
  and g52941 (n31260, n_21776, n_21777);
  not g52942 (n_21778, n31259);
  not g52943 (n_21779, n31260);
  and g52944 (n31261, n_21778, n_21779);
  not g52945 (n_21780, n31250);
  not g52946 (n_21781, n31261);
  and g52947 (n31262, n_21780, n_21781);
  and g52948 (n31263, n31250, n31261);
  not g52949 (n_21782, n31262);
  not g52950 (n_21783, n31263);
  and g52951 (n31264, n_21782, n_21783);
  not g52952 (n_21784, n31264);
  and g52953 (n31265, n31173, n_21784);
  not g52954 (n_21785, n31173);
  and g52955 (n31266, n_21785, n31264);
  not g52956 (n_21786, n31265);
  not g52957 (n_21787, n31266);
  and g52958 (n31267, n_21786, n_21787);
  and g52959 (n31268, n_21674, n_21684);
  and g52960 (n31269, n5496, n27964);
  and g52961 (n31270, n4935, n27442);
  and g52962 (n31271, n5407, n27698);
  and g52968 (n31274, n4938, n27976);
  not g52971 (n_21792, n31275);
  and g52972 (n31276, \a[20] , n_21792);
  not g52973 (n_21793, n31276);
  and g52974 (n31277, \a[20] , n_21793);
  and g52975 (n31278, n_21792, n_21793);
  not g52976 (n_21794, n31277);
  not g52977 (n_21795, n31278);
  and g52978 (n31279, n_21794, n_21795);
  not g52979 (n_21796, n31268);
  not g52980 (n_21797, n31279);
  and g52981 (n31280, n_21796, n_21797);
  not g52982 (n_21798, n31280);
  and g52983 (n31281, n_21796, n_21798);
  and g52984 (n31282, n_21797, n_21798);
  not g52985 (n_21799, n31281);
  not g52986 (n_21800, n31282);
  and g52987 (n31283, n_21799, n_21800);
  not g52988 (n_21801, n31267);
  and g52989 (n31284, n_21801, n31283);
  not g52990 (n_21802, n31283);
  and g52991 (n31285, n31267, n_21802);
  not g52992 (n_21803, n31284);
  not g52993 (n_21804, n31285);
  and g52994 (n31286, n_21803, n_21804);
  not g52995 (n_21805, n31172);
  and g52996 (n31287, n_21805, n31286);
  not g52997 (n_21806, n31286);
  and g52998 (n31288, n31172, n_21806);
  not g52999 (n_21807, n31287);
  not g53000 (n_21808, n31288);
  and g53001 (n31289, n_21807, n_21808);
  not g53002 (n_21809, n31171);
  and g53003 (n31290, n_21809, n31289);
  not g53004 (n_21810, n31289);
  and g53005 (n31291, n31171, n_21810);
  not g53006 (n_21811, n31290);
  not g53007 (n_21812, n31291);
  and g53008 (n31292, n_21811, n_21812);
  not g53009 (n_21813, n31292);
  and g53010 (n31293, n_21712, n_21813);
  and g53011 (n31294, n31168, n31292);
  not g53012 (n_21814, n31293);
  not g53013 (n_21815, n31294);
  and g53014 (\result[22] , n_21814, n_21815);
  and g53015 (n31296, n_21752, n_21765);
  and g53016 (n31297, n75, n_17020);
  and g53017 (n31298, n3020, n22320);
  and g53018 (n31299, n3023, n22326);
  and g53019 (n31300, n3028, n22323);
  and g53027 (n31304, n_21736, n_21739);
  not g53043 (n_21820, n31304);
  and g53044 (n31320, n_21820, n31319);
  not g53045 (n_21821, n31319);
  and g53046 (n31321, n31304, n_21821);
  not g53047 (n_21822, n31320);
  not g53048 (n_21823, n31321);
  and g53049 (n31322, n_21822, n_21823);
  not g53050 (n_21824, n31303);
  and g53051 (n31323, n_21824, n31322);
  not g53052 (n_21825, n31323);
  and g53053 (n31324, n_21824, n_21825);
  and g53054 (n31325, n31322, n_21825);
  not g53055 (n_21826, n31324);
  not g53056 (n_21827, n31325);
  and g53057 (n31326, n_21826, n_21827);
  and g53058 (n31327, n_21742, n_21747);
  and g53059 (n31328, n31326, n31327);
  not g53060 (n_21828, n31326);
  not g53061 (n_21829, n31327);
  and g53062 (n31329, n_21828, n_21829);
  not g53063 (n_21830, n31328);
  not g53064 (n_21831, n31329);
  and g53065 (n31330, n_21830, n_21831);
  and g53066 (n31331, n3457, n22309);
  and g53067 (n31332, n3542, n22312);
  and g53068 (n31333, n3606, n22315);
  not g53069 (n_21832, n31332);
  not g53070 (n_21833, n31333);
  and g53071 (n31334, n_21832, n_21833);
  not g53072 (n_21834, n31331);
  and g53073 (n31335, n_21834, n31334);
  and g53074 (n31336, n_489, n31335);
  and g53075 (n31337, n22529, n31335);
  not g53076 (n_21835, n31336);
  not g53077 (n_21836, n31337);
  and g53078 (n31338, n_21835, n_21836);
  not g53079 (n_21837, n31338);
  and g53080 (n31339, \a[29] , n_21837);
  and g53081 (n31340, n_15, n31338);
  not g53082 (n_21838, n31339);
  not g53083 (n_21839, n31340);
  and g53084 (n31341, n_21838, n_21839);
  not g53085 (n_21840, n31341);
  and g53086 (n31342, n31330, n_21840);
  not g53087 (n_21841, n31330);
  and g53088 (n31343, n_21841, n31341);
  not g53089 (n_21842, n31342);
  not g53090 (n_21843, n31343);
  and g53091 (n31344, n_21842, n_21843);
  not g53092 (n_21844, n31296);
  and g53093 (n31345, n_21844, n31344);
  not g53094 (n_21845, n31344);
  and g53095 (n31346, n31296, n_21845);
  not g53096 (n_21846, n31345);
  not g53097 (n_21847, n31346);
  and g53098 (n31347, n_21846, n_21847);
  and g53099 (n31348, n3884, n26060);
  and g53100 (n31349, n3967, n26063);
  and g53101 (n31350, n4046, n26066);
  and g53107 (n31353, n4050, n_18596);
  not g53110 (n_21852, n31354);
  and g53111 (n31355, \a[26] , n_21852);
  not g53112 (n_21853, n31355);
  and g53113 (n31356, \a[26] , n_21853);
  and g53114 (n31357, n_21852, n_21853);
  not g53115 (n_21854, n31356);
  not g53116 (n_21855, n31357);
  and g53117 (n31358, n_21854, n_21855);
  not g53118 (n_21856, n31358);
  and g53119 (n31359, n31347, n_21856);
  not g53120 (n_21857, n31359);
  and g53121 (n31360, n31347, n_21857);
  and g53122 (n31361, n_21856, n_21857);
  not g53123 (n_21858, n31360);
  not g53124 (n_21859, n31361);
  and g53125 (n31362, n_21858, n_21859);
  and g53126 (n31363, n_21768, n_21769);
  not g53127 (n_21860, n31363);
  and g53128 (n31364, n_21724, n_21860);
  not g53129 (n_21861, n31362);
  not g53130 (n_21862, n31364);
  and g53131 (n31365, n_21861, n_21862);
  not g53132 (n_21863, n31365);
  and g53133 (n31366, n_21861, n_21863);
  and g53134 (n31367, n_21862, n_21863);
  not g53135 (n_21864, n31366);
  not g53136 (n_21865, n31367);
  and g53137 (n31368, n_21864, n_21865);
  and g53138 (n31369, n4694, n27442);
  and g53139 (n31370, n4533, n26890);
  and g53140 (n31371, n4604, n27173);
  and g53146 (n31374, n4536, n27455);
  not g53149 (n_21870, n31375);
  and g53150 (n31376, \a[23] , n_21870);
  not g53151 (n_21871, n31376);
  and g53152 (n31377, \a[23] , n_21871);
  and g53153 (n31378, n_21870, n_21871);
  not g53154 (n_21872, n31377);
  not g53155 (n_21873, n31378);
  and g53156 (n31379, n_21872, n_21873);
  not g53157 (n_21874, n31368);
  not g53158 (n_21875, n31379);
  and g53159 (n31380, n_21874, n_21875);
  not g53160 (n_21876, n31380);
  and g53161 (n31381, n_21874, n_21876);
  and g53162 (n31382, n_21875, n_21876);
  not g53163 (n_21877, n31381);
  not g53164 (n_21878, n31382);
  and g53165 (n31383, n_21877, n_21878);
  and g53166 (n31384, n_21782, n_21787);
  and g53167 (n31385, n31383, n31384);
  not g53168 (n_21879, n31383);
  not g53169 (n_21880, n31384);
  and g53170 (n31386, n_21879, n_21880);
  not g53171 (n_21881, n31385);
  not g53172 (n_21882, n31386);
  and g53173 (n31387, n_21881, n_21882);
  and g53174 (n31388, n5496, n_19417);
  and g53175 (n31389, n4935, n27698);
  and g53176 (n31390, n5407, n27964);
  and g53182 (n31393, n4938, n_19940);
  not g53185 (n_21887, n31394);
  and g53186 (n31395, \a[20] , n_21887);
  not g53187 (n_21888, n31395);
  and g53188 (n31396, \a[20] , n_21888);
  and g53189 (n31397, n_21887, n_21888);
  not g53190 (n_21889, n31396);
  not g53191 (n_21890, n31397);
  and g53192 (n31398, n_21889, n_21890);
  not g53193 (n_21891, n31398);
  and g53194 (n31399, n31387, n_21891);
  not g53195 (n_21892, n31399);
  and g53196 (n31400, n31387, n_21892);
  and g53197 (n31401, n_21891, n_21892);
  not g53198 (n_21893, n31400);
  not g53199 (n_21894, n31401);
  and g53200 (n31402, n_21893, n_21894);
  and g53201 (n31403, n_21798, n_21804);
  not g53202 (n_21895, n31402);
  not g53203 (n_21896, n31403);
  and g53204 (n31404, n_21895, n_21896);
  not g53205 (n_21897, n31404);
  and g53206 (n31405, n_21895, n_21897);
  and g53207 (n31406, n_21896, n_21897);
  not g53208 (n_21898, n31405);
  not g53209 (n_21899, n31406);
  and g53210 (n31407, n_21898, n_21899);
  and g53211 (n31408, n_21807, n_21811);
  and g53212 (n31409, n31407, n31408);
  not g53213 (n_21900, n31407);
  not g53214 (n_21901, n31408);
  and g53215 (n31410, n_21900, n_21901);
  not g53216 (n_21902, n31409);
  not g53217 (n_21903, n31410);
  and g53218 (n31411, n_21902, n_21903);
  and g53219 (n31412, n_21815, n31411);
  not g53220 (n_21904, n31411);
  and g53221 (n31413, n31294, n_21904);
  or g53222 (\result[23] , n31412, n31413);
  and g53223 (n31415, n31294, n31411);
  and g53224 (n31416, n75, n_17004);
  and g53225 (n31417, n3020, n22312);
  and g53226 (n31418, n3023, n22323);
  and g53227 (n31419, n3028, n22320);
  and g53248 (n31436, n_21821, n31435);
  not g53249 (n_21909, n31435);
  and g53250 (n31437, n31319, n_21909);
  not g53251 (n_21910, n31422);
  not g53252 (n_21911, n31437);
  and g53253 (n31438, n_21910, n_21911);
  not g53254 (n_21912, n31436);
  and g53255 (n31439, n_21912, n31438);
  not g53256 (n_21913, n31439);
  and g53257 (n31440, n_21910, n_21913);
  and g53258 (n31441, n_21911, n_21913);
  and g53259 (n31442, n_21912, n31441);
  not g53260 (n_21914, n31440);
  not g53261 (n_21915, n31442);
  and g53262 (n31443, n_21914, n_21915);
  and g53263 (n31444, n_21822, n_21825);
  and g53264 (n31445, n31443, n31444);
  not g53265 (n_21916, n31443);
  not g53266 (n_21917, n31444);
  and g53267 (n31446, n_21916, n_21917);
  not g53268 (n_21918, n31445);
  not g53269 (n_21919, n31446);
  and g53270 (n31447, n_21918, n_21919);
  and g53271 (n31448, n_21831, n_21842);
  not g53272 (n_21920, n31447);
  and g53273 (n31449, n_21920, n31448);
  not g53274 (n_21921, n31448);
  and g53275 (n31450, n31447, n_21921);
  not g53276 (n_21922, n31449);
  not g53277 (n_21923, n31450);
  and g53278 (n31451, n_21922, n_21923);
  and g53279 (n31452, n3457, n26063);
  and g53280 (n31453, n3542, n22315);
  and g53281 (n31454, n3606, n22309);
  and g53287 (n31457, n3368, n_18124);
  not g53290 (n_21928, n31458);
  and g53291 (n31459, \a[29] , n_21928);
  not g53292 (n_21929, n31459);
  and g53293 (n31460, \a[29] , n_21929);
  and g53294 (n31461, n_21928, n_21929);
  not g53295 (n_21930, n31460);
  not g53296 (n_21931, n31461);
  and g53297 (n31462, n_21930, n_21931);
  not g53298 (n_21932, n31462);
  and g53299 (n31463, n31451, n_21932);
  not g53300 (n_21933, n31463);
  and g53301 (n31464, n31451, n_21933);
  and g53302 (n31465, n_21932, n_21933);
  not g53303 (n_21934, n31464);
  not g53304 (n_21935, n31465);
  and g53305 (n31466, n_21934, n_21935);
  and g53306 (n31467, n3884, n26890);
  and g53307 (n31468, n3967, n26066);
  and g53308 (n31469, n4046, n26060);
  and g53314 (n31472, n4050, n_18823);
  not g53317 (n_21940, n31473);
  and g53318 (n31474, \a[26] , n_21940);
  not g53319 (n_21941, n31474);
  and g53320 (n31475, \a[26] , n_21941);
  and g53321 (n31476, n_21940, n_21941);
  not g53322 (n_21942, n31475);
  not g53323 (n_21943, n31476);
  and g53324 (n31477, n_21942, n_21943);
  not g53325 (n_21944, n31466);
  not g53326 (n_21945, n31477);
  and g53327 (n31478, n_21944, n_21945);
  not g53328 (n_21946, n31478);
  and g53329 (n31479, n_21944, n_21946);
  and g53330 (n31480, n_21945, n_21946);
  not g53331 (n_21947, n31479);
  not g53332 (n_21948, n31480);
  and g53333 (n31481, n_21947, n_21948);
  and g53334 (n31482, n_21846, n_21857);
  and g53335 (n31483, n31481, n31482);
  not g53336 (n_21949, n31481);
  not g53337 (n_21950, n31482);
  and g53338 (n31484, n_21949, n_21950);
  not g53339 (n_21951, n31483);
  not g53340 (n_21952, n31484);
  and g53341 (n31485, n_21951, n_21952);
  and g53342 (n31486, n4694, n27698);
  and g53343 (n31487, n4533, n27173);
  and g53344 (n31488, n4604, n27442);
  and g53350 (n31491, n4536, n_19446);
  not g53353 (n_21957, n31492);
  and g53354 (n31493, \a[23] , n_21957);
  not g53355 (n_21958, n31493);
  and g53356 (n31494, \a[23] , n_21958);
  and g53357 (n31495, n_21957, n_21958);
  not g53358 (n_21959, n31494);
  not g53359 (n_21960, n31495);
  and g53360 (n31496, n_21959, n_21960);
  not g53361 (n_21961, n31496);
  and g53362 (n31497, n31485, n_21961);
  not g53363 (n_21962, n31497);
  and g53364 (n31498, n31485, n_21962);
  and g53365 (n31499, n_21961, n_21962);
  not g53366 (n_21963, n31498);
  not g53367 (n_21964, n31499);
  and g53368 (n31500, n_21963, n_21964);
  and g53369 (n31501, n_21863, n_21876);
  and g53370 (n31502, n_7989, n_19417);
  and g53371 (n31503, n4935, n27964);
  not g53372 (n_21965, n31502);
  not g53373 (n_21966, n31503);
  and g53374 (n31504, n_21965, n_21966);
  and g53375 (n31505, n_1011, n31504);
  and g53376 (n31506, n28221, n31504);
  not g53377 (n_21967, n31505);
  not g53378 (n_21968, n31506);
  and g53379 (n31507, n_21967, n_21968);
  not g53380 (n_21969, n31507);
  and g53381 (n31508, \a[20] , n_21969);
  and g53382 (n31509, n_435, n31507);
  not g53383 (n_21970, n31508);
  not g53384 (n_21971, n31509);
  and g53385 (n31510, n_21970, n_21971);
  not g53386 (n_21972, n31501);
  not g53387 (n_21973, n31510);
  and g53388 (n31511, n_21972, n_21973);
  and g53389 (n31512, n31501, n31510);
  not g53390 (n_21974, n31511);
  not g53391 (n_21975, n31512);
  and g53392 (n31513, n_21974, n_21975);
  not g53393 (n_21976, n31500);
  and g53394 (n31514, n_21976, n31513);
  not g53395 (n_21977, n31514);
  and g53396 (n31515, n_21976, n_21977);
  and g53397 (n31516, n31513, n_21977);
  not g53398 (n_21978, n31515);
  not g53399 (n_21979, n31516);
  and g53400 (n31517, n_21978, n_21979);
  and g53401 (n31518, n_21882, n_21892);
  and g53402 (n31519, n31517, n31518);
  not g53403 (n_21980, n31517);
  not g53404 (n_21981, n31518);
  and g53405 (n31520, n_21980, n_21981);
  not g53406 (n_21982, n31519);
  not g53407 (n_21983, n31520);
  and g53408 (n31521, n_21982, n_21983);
  and g53409 (n31522, n_21897, n_21903);
  not g53410 (n_21984, n31521);
  and g53411 (n31523, n_21984, n31522);
  not g53412 (n_21985, n31522);
  and g53413 (n31524, n31521, n_21985);
  not g53414 (n_21986, n31523);
  not g53415 (n_21987, n31524);
  and g53416 (n31525, n_21986, n_21987);
  and g53417 (n31526, n31415, n31525);
  not g53418 (n_21988, n31415);
  not g53419 (n_21989, n31525);
  and g53420 (n31527, n_21988, n_21989);
  not g53421 (n_21990, n31526);
  not g53422 (n_21991, n31527);
  and g53423 (\result[24] , n_21990, n_21991);
  and g53424 (n31529, n_21983, n_21987);
  and g53425 (n31530, n_21974, n_21977);
  and g53426 (n31531, n75, n25294);
  and g53427 (n31532, n3020, n22315);
  and g53428 (n31533, n3023, n22320);
  and g53429 (n31534, n3028, n22312);
  and g53437 (n31538, n_7418, n_19417);
  not g53438 (n_21996, n31538);
  and g53439 (n31539, \a[20] , n_21996);
  and g53440 (n31540, n_435, n31538);
  not g53441 (n_21997, n31539);
  not g53442 (n_21998, n31540);
  and g53443 (n31541, n_21997, n_21998);
  and g53461 (n31559, n31319, n31558);
  not g53462 (n_21999, n31558);
  and g53463 (n31560, n_21821, n_21999);
  not g53464 (n_22000, n31559);
  not g53465 (n_22001, n31560);
  and g53466 (n31561, n_22000, n_22001);
  and g53467 (n31562, n31541, n31561);
  not g53468 (n_22002, n31541);
  not g53469 (n_22003, n31561);
  and g53470 (n31563, n_22002, n_22003);
  not g53471 (n_22004, n31562);
  not g53472 (n_22005, n31563);
  and g53473 (n31564, n_22004, n_22005);
  not g53474 (n_22006, n31441);
  and g53475 (n31565, n_22006, n31564);
  not g53476 (n_22007, n31564);
  and g53477 (n31566, n31441, n_22007);
  not g53478 (n_22008, n31565);
  not g53479 (n_22009, n31566);
  and g53480 (n31567, n_22008, n_22009);
  not g53481 (n_22010, n31537);
  and g53482 (n31568, n_22010, n31567);
  not g53483 (n_22011, n31568);
  and g53484 (n31569, n31567, n_22011);
  and g53485 (n31570, n_22010, n_22011);
  not g53486 (n_22012, n31569);
  not g53487 (n_22013, n31570);
  and g53488 (n31571, n_22012, n_22013);
  and g53489 (n31572, n_21919, n_21923);
  and g53490 (n31573, n31571, n31572);
  not g53491 (n_22014, n31571);
  not g53492 (n_22015, n31572);
  and g53493 (n31574, n_22014, n_22015);
  not g53494 (n_22016, n31573);
  not g53495 (n_22017, n31574);
  and g53496 (n31575, n_22016, n_22017);
  and g53497 (n31576, n3457, n26066);
  and g53498 (n31577, n3542, n22309);
  and g53499 (n31578, n3606, n26063);
  and g53505 (n31581, n3368, n_18359);
  not g53508 (n_22022, n31582);
  and g53509 (n31583, \a[29] , n_22022);
  not g53510 (n_22023, n31583);
  and g53511 (n31584, \a[29] , n_22023);
  and g53512 (n31585, n_22022, n_22023);
  not g53513 (n_22024, n31584);
  not g53514 (n_22025, n31585);
  and g53515 (n31586, n_22024, n_22025);
  not g53516 (n_22026, n31586);
  and g53517 (n31587, n31575, n_22026);
  not g53518 (n_22027, n31587);
  and g53519 (n31588, n31575, n_22027);
  and g53520 (n31589, n_22026, n_22027);
  not g53521 (n_22028, n31588);
  not g53522 (n_22029, n31589);
  and g53523 (n31590, n_22028, n_22029);
  and g53524 (n31591, n3884, n27173);
  and g53525 (n31592, n3967, n26060);
  and g53526 (n31593, n4046, n26890);
  and g53532 (n31596, n4050, n27185);
  not g53535 (n_22034, n31597);
  and g53536 (n31598, \a[26] , n_22034);
  not g53537 (n_22035, n31598);
  and g53538 (n31599, \a[26] , n_22035);
  and g53539 (n31600, n_22034, n_22035);
  not g53540 (n_22036, n31599);
  not g53541 (n_22037, n31600);
  and g53542 (n31601, n_22036, n_22037);
  not g53543 (n_22038, n31590);
  not g53544 (n_22039, n31601);
  and g53545 (n31602, n_22038, n_22039);
  not g53546 (n_22040, n31602);
  and g53547 (n31603, n_22038, n_22040);
  and g53548 (n31604, n_22039, n_22040);
  not g53549 (n_22041, n31603);
  not g53550 (n_22042, n31604);
  and g53551 (n31605, n_22041, n_22042);
  and g53552 (n31606, n_21933, n_21946);
  and g53553 (n31607, n31605, n31606);
  not g53554 (n_22043, n31605);
  not g53555 (n_22044, n31606);
  and g53556 (n31608, n_22043, n_22044);
  not g53557 (n_22045, n31607);
  not g53558 (n_22046, n31608);
  and g53559 (n31609, n_22045, n_22046);
  and g53560 (n31610, n_21952, n_21962);
  and g53561 (n31611, n4694, n27964);
  and g53562 (n31612, n4533, n27442);
  and g53563 (n31613, n4604, n27698);
  and g53569 (n31616, n4536, n27976);
  not g53572 (n_22051, n31617);
  and g53573 (n31618, \a[23] , n_22051);
  not g53574 (n_22052, n31618);
  and g53575 (n31619, \a[23] , n_22052);
  and g53576 (n31620, n_22051, n_22052);
  not g53577 (n_22053, n31619);
  not g53578 (n_22054, n31620);
  and g53579 (n31621, n_22053, n_22054);
  not g53580 (n_22055, n31610);
  not g53581 (n_22056, n31621);
  and g53582 (n31622, n_22055, n_22056);
  not g53583 (n_22057, n31622);
  and g53584 (n31623, n_22055, n_22057);
  and g53585 (n31624, n_22056, n_22057);
  not g53586 (n_22058, n31623);
  not g53587 (n_22059, n31624);
  and g53588 (n31625, n_22058, n_22059);
  not g53589 (n_22060, n31609);
  and g53590 (n31626, n_22060, n31625);
  not g53591 (n_22061, n31625);
  and g53592 (n31627, n31609, n_22061);
  not g53593 (n_22062, n31626);
  not g53594 (n_22063, n31627);
  and g53595 (n31628, n_22062, n_22063);
  not g53596 (n_22064, n31530);
  and g53597 (n31629, n_22064, n31628);
  not g53598 (n_22065, n31628);
  and g53599 (n31630, n31530, n_22065);
  not g53600 (n_22066, n31629);
  not g53601 (n_22067, n31630);
  and g53602 (n31631, n_22066, n_22067);
  not g53603 (n_22068, n31529);
  and g53604 (n31632, n_22068, n31631);
  not g53605 (n_22069, n31631);
  and g53606 (n31633, n31529, n_22069);
  not g53607 (n_22070, n31632);
  not g53608 (n_22071, n31633);
  and g53609 (n31634, n_22070, n_22071);
  not g53610 (n_22072, n31634);
  and g53611 (n31635, n_21990, n_22072);
  and g53612 (n31636, n31526, n31634);
  not g53613 (n_22073, n31635);
  not g53614 (n_22074, n31636);
  and g53615 (\result[25] , n_22073, n_22074);
  and g53616 (n31638, n_22017, n_22027);
  and g53617 (n31639, n75, n_14657);
  and g53618 (n31640, n3020, n22309);
  and g53619 (n31641, n3023, n22312);
  and g53620 (n31642, n3028, n22315);
  and g53628 (n31646, n_22001, n_22004);
  not g53644 (n_22079, n31646);
  and g53645 (n31662, n_22079, n31661);
  not g53646 (n_22080, n31661);
  and g53647 (n31663, n31646, n_22080);
  not g53648 (n_22081, n31662);
  not g53649 (n_22082, n31663);
  and g53650 (n31664, n_22081, n_22082);
  not g53651 (n_22083, n31645);
  and g53652 (n31665, n_22083, n31664);
  not g53653 (n_22084, n31665);
  and g53654 (n31666, n_22083, n_22084);
  and g53655 (n31667, n31664, n_22084);
  not g53656 (n_22085, n31666);
  not g53657 (n_22086, n31667);
  and g53658 (n31668, n_22085, n_22086);
  and g53659 (n31669, n_22008, n_22011);
  and g53660 (n31670, n31668, n31669);
  not g53661 (n_22087, n31668);
  not g53662 (n_22088, n31669);
  and g53663 (n31671, n_22087, n_22088);
  not g53664 (n_22089, n31670);
  not g53665 (n_22090, n31671);
  and g53666 (n31672, n_22089, n_22090);
  and g53667 (n31673, n3457, n26060);
  and g53668 (n31674, n3542, n26063);
  and g53669 (n31675, n3606, n26066);
  not g53670 (n_22091, n31674);
  not g53671 (n_22092, n31675);
  and g53672 (n31676, n_22091, n_22092);
  not g53673 (n_22093, n31673);
  and g53674 (n31677, n_22093, n31676);
  and g53675 (n31678, n_489, n31677);
  and g53676 (n31679, n26088, n31677);
  not g53677 (n_22094, n31678);
  not g53678 (n_22095, n31679);
  and g53679 (n31680, n_22094, n_22095);
  not g53680 (n_22096, n31680);
  and g53681 (n31681, \a[29] , n_22096);
  and g53682 (n31682, n_15, n31680);
  not g53683 (n_22097, n31681);
  not g53684 (n_22098, n31682);
  and g53685 (n31683, n_22097, n_22098);
  not g53686 (n_22099, n31683);
  and g53687 (n31684, n31672, n_22099);
  not g53688 (n_22100, n31672);
  and g53689 (n31685, n_22100, n31683);
  not g53690 (n_22101, n31684);
  not g53691 (n_22102, n31685);
  and g53692 (n31686, n_22101, n_22102);
  not g53693 (n_22103, n31638);
  and g53694 (n31687, n_22103, n31686);
  not g53695 (n_22104, n31686);
  and g53696 (n31688, n31638, n_22104);
  not g53697 (n_22105, n31687);
  not g53698 (n_22106, n31688);
  and g53699 (n31689, n_22105, n_22106);
  and g53700 (n31690, n3884, n27442);
  and g53701 (n31691, n3967, n26890);
  and g53702 (n31692, n4046, n27173);
  and g53708 (n31695, n4050, n27455);
  not g53711 (n_22111, n31696);
  and g53712 (n31697, \a[26] , n_22111);
  not g53713 (n_22112, n31697);
  and g53714 (n31698, \a[26] , n_22112);
  and g53715 (n31699, n_22111, n_22112);
  not g53716 (n_22113, n31698);
  not g53717 (n_22114, n31699);
  and g53718 (n31700, n_22113, n_22114);
  not g53719 (n_22115, n31700);
  and g53720 (n31701, n31689, n_22115);
  not g53721 (n_22116, n31701);
  and g53722 (n31702, n31689, n_22116);
  and g53723 (n31703, n_22115, n_22116);
  not g53724 (n_22117, n31702);
  not g53725 (n_22118, n31703);
  and g53726 (n31704, n_22117, n_22118);
  and g53727 (n31705, n_22040, n_22046);
  and g53728 (n31706, n31704, n31705);
  not g53729 (n_22119, n31704);
  not g53730 (n_22120, n31705);
  and g53731 (n31707, n_22119, n_22120);
  not g53732 (n_22121, n31706);
  not g53733 (n_22122, n31707);
  and g53734 (n31708, n_22121, n_22122);
  and g53735 (n31709, n4694, n_19417);
  and g53736 (n31710, n4533, n27698);
  and g53737 (n31711, n4604, n27964);
  and g53743 (n31714, n4536, n_19940);
  not g53746 (n_22127, n31715);
  and g53747 (n31716, \a[23] , n_22127);
  not g53748 (n_22128, n31716);
  and g53749 (n31717, \a[23] , n_22128);
  and g53750 (n31718, n_22127, n_22128);
  not g53751 (n_22129, n31717);
  not g53752 (n_22130, n31718);
  and g53753 (n31719, n_22129, n_22130);
  not g53754 (n_22131, n31719);
  and g53755 (n31720, n31708, n_22131);
  not g53756 (n_22132, n31720);
  and g53757 (n31721, n31708, n_22132);
  and g53758 (n31722, n_22131, n_22132);
  not g53759 (n_22133, n31721);
  not g53760 (n_22134, n31722);
  and g53761 (n31723, n_22133, n_22134);
  and g53762 (n31724, n_22057, n_22063);
  not g53763 (n_22135, n31723);
  not g53764 (n_22136, n31724);
  and g53765 (n31725, n_22135, n_22136);
  not g53766 (n_22137, n31725);
  and g53767 (n31726, n_22135, n_22137);
  and g53768 (n31727, n_22136, n_22137);
  not g53769 (n_22138, n31726);
  not g53770 (n_22139, n31727);
  and g53771 (n31728, n_22138, n_22139);
  and g53772 (n31729, n_22066, n_22070);
  and g53773 (n31730, n31728, n31729);
  not g53774 (n_22140, n31728);
  not g53775 (n_22141, n31729);
  and g53776 (n31731, n_22140, n_22141);
  not g53777 (n_22142, n31730);
  not g53778 (n_22143, n31731);
  and g53779 (n31732, n_22142, n_22143);
  not g53780 (n_22144, n31732);
  and g53781 (n31733, n31636, n_22144);
  and g53782 (n31734, n_22074, n31732);
  or g53783 (\result[26] , n31733, n31734);
  and g53784 (n31736, n_22081, n_22084);
  not g53800 (n_22145, n31751);
  and g53801 (n31752, n31661, n_22145);
  and g53802 (n31753, n_22080, n31751);
  not g53803 (n_22146, n31736);
  not g53804 (n_22147, n31753);
  and g53805 (n31754, n_22146, n_22147);
  not g53806 (n_22148, n31752);
  and g53807 (n31755, n_22148, n31754);
  not g53808 (n_22149, n31755);
  and g53809 (n31756, n_22146, n_22149);
  and g53810 (n31757, n_22147, n_22149);
  and g53811 (n31758, n_22148, n31757);
  not g53812 (n_22150, n31756);
  not g53813 (n_22151, n31758);
  and g53814 (n31759, n_22150, n_22151);
  and g53815 (n31760, n75, n_18124);
  and g53816 (n31761, n3020, n26063);
  and g53817 (n31762, n3023, n22315);
  and g53818 (n31763, n3028, n22309);
  not g53826 (n_22156, n31759);
  not g53827 (n_22157, n31766);
  and g53828 (n31767, n_22156, n_22157);
  not g53829 (n_22158, n31767);
  and g53830 (n31768, n_22156, n_22158);
  and g53831 (n31769, n_22157, n_22158);
  not g53832 (n_22159, n31768);
  not g53833 (n_22160, n31769);
  and g53834 (n31770, n_22159, n_22160);
  and g53835 (n31771, n_22090, n_22101);
  and g53836 (n31772, n31770, n31771);
  not g53837 (n_22161, n31770);
  not g53838 (n_22162, n31771);
  and g53839 (n31773, n_22161, n_22162);
  not g53840 (n_22163, n31772);
  not g53841 (n_22164, n31773);
  and g53842 (n31774, n_22163, n_22164);
  and g53843 (n31775, n3457, n26890);
  and g53844 (n31776, n3542, n26066);
  and g53845 (n31777, n3606, n26060);
  and g53851 (n31780, n3368, n_18823);
  not g53854 (n_22169, n31781);
  and g53855 (n31782, \a[29] , n_22169);
  not g53856 (n_22170, n31782);
  and g53857 (n31783, \a[29] , n_22170);
  and g53858 (n31784, n_22169, n_22170);
  not g53859 (n_22171, n31783);
  not g53860 (n_22172, n31784);
  and g53861 (n31785, n_22171, n_22172);
  not g53862 (n_22173, n31785);
  and g53863 (n31786, n31774, n_22173);
  not g53864 (n_22174, n31786);
  and g53865 (n31787, n31774, n_22174);
  and g53866 (n31788, n_22173, n_22174);
  not g53867 (n_22175, n31787);
  not g53868 (n_22176, n31788);
  and g53869 (n31789, n_22175, n_22176);
  and g53870 (n31790, n3884, n27698);
  and g53871 (n31791, n3967, n27173);
  and g53872 (n31792, n4046, n27442);
  and g53878 (n31795, n4050, n_19446);
  not g53881 (n_22181, n31796);
  and g53882 (n31797, \a[26] , n_22181);
  not g53883 (n_22182, n31797);
  and g53884 (n31798, \a[26] , n_22182);
  and g53885 (n31799, n_22181, n_22182);
  not g53886 (n_22183, n31798);
  not g53887 (n_22184, n31799);
  and g53888 (n31800, n_22183, n_22184);
  not g53889 (n_22185, n31789);
  not g53890 (n_22186, n31800);
  and g53891 (n31801, n_22185, n_22186);
  not g53892 (n_22187, n31801);
  and g53893 (n31802, n_22185, n_22187);
  and g53894 (n31803, n_22186, n_22187);
  not g53895 (n_22188, n31802);
  not g53896 (n_22189, n31803);
  and g53897 (n31804, n_22188, n_22189);
  and g53898 (n31805, n_22105, n_22116);
  and g53899 (n31806, n_7705, n_19417);
  and g53900 (n31807, n4533, n27964);
  not g53901 (n_22190, n31806);
  not g53902 (n_22191, n31807);
  and g53903 (n31808, n_22190, n_22191);
  and g53904 (n31809, n_732, n31808);
  and g53905 (n31810, n28221, n31808);
  not g53906 (n_22192, n31809);
  not g53907 (n_22193, n31810);
  and g53908 (n31811, n_22192, n_22193);
  not g53909 (n_22194, n31811);
  and g53910 (n31812, \a[23] , n_22194);
  and g53911 (n31813, n_27, n31811);
  not g53912 (n_22195, n31812);
  not g53913 (n_22196, n31813);
  and g53914 (n31814, n_22195, n_22196);
  not g53915 (n_22197, n31805);
  not g53916 (n_22198, n31814);
  and g53917 (n31815, n_22197, n_22198);
  and g53918 (n31816, n31805, n31814);
  not g53919 (n_22199, n31815);
  not g53920 (n_22200, n31816);
  and g53921 (n31817, n_22199, n_22200);
  not g53922 (n_22201, n31804);
  and g53923 (n31818, n_22201, n31817);
  not g53924 (n_22202, n31818);
  and g53925 (n31819, n_22201, n_22202);
  and g53926 (n31820, n31817, n_22202);
  not g53927 (n_22203, n31819);
  not g53928 (n_22204, n31820);
  and g53929 (n31821, n_22203, n_22204);
  and g53930 (n31822, n_22122, n_22132);
  and g53931 (n31823, n31821, n31822);
  not g53932 (n_22205, n31821);
  not g53933 (n_22206, n31822);
  and g53934 (n31824, n_22205, n_22206);
  not g53935 (n_22207, n31823);
  not g53936 (n_22208, n31824);
  and g53937 (n31825, n_22207, n_22208);
  and g53938 (n31826, n_22137, n_22143);
  not g53939 (n_22209, n31825);
  and g53940 (n31827, n_22209, n31826);
  not g53941 (n_22210, n31826);
  and g53942 (n31828, n31825, n_22210);
  not g53943 (n_22211, n31827);
  not g53944 (n_22212, n31828);
  and g53945 (n31829, n_22211, n_22212);
  and g53946 (n31830, n31636, n31732);
  and g53947 (n31831, n31829, n31830);
  not g53948 (n_22213, n31829);
  not g53949 (n_22214, n31830);
  and g53950 (n31832, n_22213, n_22214);
  not g53951 (n_22215, n31831);
  not g53952 (n_22216, n31832);
  and g53953 (\result[27] , n_22215, n_22216);
  and g53954 (n31834, n_22208, n_22212);
  and g53955 (n31835, n_22199, n_22202);
  and g53956 (n31836, n_22174, n_22187);
  and g53957 (n31837, n3884, n27964);
  and g53958 (n31838, n3967, n27442);
  and g53959 (n31839, n4046, n27698);
  and g53965 (n31842, n4050, n27976);
  not g53968 (n_22221, n31843);
  and g53969 (n31844, \a[26] , n_22221);
  not g53970 (n_22222, n31844);
  and g53971 (n31845, \a[26] , n_22222);
  and g53972 (n31846, n_22221, n_22222);
  not g53973 (n_22223, n31845);
  not g53974 (n_22224, n31846);
  and g53975 (n31847, n_22223, n_22224);
  not g53976 (n_22225, n31836);
  not g53977 (n_22226, n31847);
  and g53978 (n31848, n_22225, n_22226);
  not g53979 (n_22227, n31848);
  and g53980 (n31849, n_22225, n_22227);
  and g53981 (n31850, n_22226, n_22227);
  not g53982 (n_22228, n31849);
  not g53983 (n_22229, n31850);
  and g53984 (n31851, n_22228, n_22229);
  and g53985 (n31852, n75, n_18359);
  and g53986 (n31853, n3020, n26066);
  and g53987 (n31854, n3023, n22309);
  and g53988 (n31855, n3028, n26063);
  and g53996 (n31859, n_14400, n_19417);
  not g53997 (n_22234, n31859);
  and g53998 (n31860, \a[23] , n_22234);
  and g53999 (n31861, n_27, n31859);
  not g54000 (n_22235, n31860);
  not g54001 (n_22236, n31861);
  and g54002 (n31862, n_22235, n_22236);
  and g54017 (n31877, n31751, n31876);
  not g54018 (n_22237, n31876);
  and g54019 (n31878, n_22145, n_22237);
  not g54020 (n_22238, n31877);
  not g54021 (n_22239, n31878);
  and g54022 (n31879, n_22238, n_22239);
  and g54023 (n31880, n31862, n31879);
  not g54024 (n_22240, n31862);
  not g54025 (n_22241, n31879);
  and g54026 (n31881, n_22240, n_22241);
  not g54027 (n_22242, n31880);
  not g54028 (n_22243, n31881);
  and g54029 (n31882, n_22242, n_22243);
  not g54030 (n_22244, n31757);
  and g54031 (n31883, n_22244, n31882);
  not g54032 (n_22245, n31882);
  and g54033 (n31884, n31757, n_22245);
  not g54034 (n_22246, n31883);
  not g54035 (n_22247, n31884);
  and g54036 (n31885, n_22246, n_22247);
  not g54037 (n_22248, n31858);
  and g54038 (n31886, n_22248, n31885);
  not g54039 (n_22249, n31886);
  and g54040 (n31887, n31885, n_22249);
  and g54041 (n31888, n_22248, n_22249);
  not g54042 (n_22250, n31887);
  not g54043 (n_22251, n31888);
  and g54044 (n31889, n_22250, n_22251);
  and g54045 (n31890, n_22158, n_22164);
  and g54046 (n31891, n31889, n31890);
  not g54047 (n_22252, n31889);
  not g54048 (n_22253, n31890);
  and g54049 (n31892, n_22252, n_22253);
  not g54050 (n_22254, n31891);
  not g54051 (n_22255, n31892);
  and g54052 (n31893, n_22254, n_22255);
  and g54053 (n31894, n3457, n27173);
  and g54054 (n31895, n3542, n26060);
  and g54055 (n31896, n3606, n26890);
  and g54061 (n31899, n3368, n27185);
  not g54064 (n_22260, n31900);
  and g54065 (n31901, \a[29] , n_22260);
  not g54066 (n_22261, n31901);
  and g54067 (n31902, \a[29] , n_22261);
  and g54068 (n31903, n_22260, n_22261);
  not g54069 (n_22262, n31902);
  not g54070 (n_22263, n31903);
  and g54071 (n31904, n_22262, n_22263);
  not g54072 (n_22264, n31904);
  and g54073 (n31905, n31893, n_22264);
  not g54074 (n_22265, n31905);
  and g54075 (n31906, n31893, n_22265);
  and g54076 (n31907, n_22264, n_22265);
  not g54077 (n_22266, n31906);
  not g54078 (n_22267, n31907);
  and g54079 (n31908, n_22266, n_22267);
  not g54080 (n_22268, n31851);
  and g54081 (n31909, n_22268, n31908);
  not g54082 (n_22269, n31908);
  and g54083 (n31910, n31851, n_22269);
  not g54084 (n_22270, n31909);
  not g54085 (n_22271, n31910);
  and g54086 (n31911, n_22270, n_22271);
  not g54087 (n_22272, n31835);
  not g54088 (n_22273, n31911);
  and g54089 (n31912, n_22272, n_22273);
  and g54090 (n31913, n31835, n31911);
  not g54091 (n_22274, n31912);
  not g54092 (n_22275, n31913);
  and g54093 (n31914, n_22274, n_22275);
  not g54094 (n_22276, n31834);
  and g54095 (n31915, n_22276, n31914);
  not g54096 (n_22277, n31914);
  and g54097 (n31916, n31834, n_22277);
  not g54098 (n_22278, n31915);
  not g54099 (n_22279, n31916);
  and g54100 (n31917, n_22278, n_22279);
  not g54101 (n_22280, n31917);
  and g54102 (n31918, n_22215, n_22280);
  and g54103 (n31919, n31831, n31917);
  not g54104 (n_22281, n31918);
  not g54105 (n_22282, n31919);
  and g54106 (\result[28] , n_22281, n_22282);
  and g54107 (n31921, n_22255, n_22265);
  and g54108 (n31922, n75, n_18596);
  and g54109 (n31923, n3020, n26060);
  and g54110 (n31924, n3023, n26063);
  and g54111 (n31925, n3028, n26066);
  and g54119 (n31929, n_22239, n_22242);
  not g54136 (n_22287, n31929);
  and g54137 (n31946, n_22287, n31945);
  not g54138 (n_22288, n31945);
  and g54139 (n31947, n31929, n_22288);
  not g54140 (n_22289, n31946);
  not g54141 (n_22290, n31947);
  and g54142 (n31948, n_22289, n_22290);
  not g54143 (n_22291, n31928);
  and g54144 (n31949, n_22291, n31948);
  not g54145 (n_22292, n31949);
  and g54146 (n31950, n_22291, n_22292);
  and g54147 (n31951, n31948, n_22292);
  not g54148 (n_22293, n31950);
  not g54149 (n_22294, n31951);
  and g54150 (n31952, n_22293, n_22294);
  and g54151 (n31953, n_22246, n_22249);
  and g54152 (n31954, n31952, n31953);
  not g54153 (n_22295, n31952);
  not g54154 (n_22296, n31953);
  and g54155 (n31955, n_22295, n_22296);
  not g54156 (n_22297, n31954);
  not g54157 (n_22298, n31955);
  and g54158 (n31956, n_22297, n_22298);
  and g54159 (n31957, n3457, n27442);
  and g54160 (n31958, n3542, n26890);
  and g54161 (n31959, n3606, n27173);
  not g54162 (n_22299, n31958);
  not g54163 (n_22300, n31959);
  and g54164 (n31960, n_22299, n_22300);
  not g54165 (n_22301, n31957);
  and g54166 (n31961, n_22301, n31960);
  and g54167 (n31962, n_489, n31961);
  and g54168 (n31963, n_18803, n31961);
  not g54169 (n_22302, n31962);
  not g54170 (n_22303, n31963);
  and g54171 (n31964, n_22302, n_22303);
  not g54172 (n_22304, n31964);
  and g54173 (n31965, \a[29] , n_22304);
  and g54174 (n31966, n_15, n31964);
  not g54175 (n_22305, n31965);
  not g54176 (n_22306, n31966);
  and g54177 (n31967, n_22305, n_22306);
  not g54178 (n_22307, n31967);
  and g54179 (n31968, n31956, n_22307);
  not g54180 (n_22308, n31956);
  and g54181 (n31969, n_22308, n31967);
  not g54182 (n_22309, n31968);
  not g54183 (n_22310, n31969);
  and g54184 (n31970, n_22309, n_22310);
  not g54185 (n_22311, n31921);
  and g54186 (n31971, n_22311, n31970);
  not g54187 (n_22312, n31970);
  and g54188 (n31972, n31921, n_22312);
  not g54189 (n_22313, n31971);
  not g54190 (n_22314, n31972);
  and g54191 (n31973, n_22313, n_22314);
  and g54192 (n31974, n3884, n_19417);
  and g54193 (n31975, n3967, n27698);
  and g54194 (n31976, n4046, n27964);
  and g54200 (n31979, n4050, n_19940);
  not g54203 (n_22319, n31980);
  and g54204 (n31981, \a[26] , n_22319);
  not g54205 (n_22320, n31981);
  and g54206 (n31982, \a[26] , n_22320);
  and g54207 (n31983, n_22319, n_22320);
  not g54208 (n_22321, n31982);
  not g54209 (n_22322, n31983);
  and g54210 (n31984, n_22321, n_22322);
  not g54211 (n_22323, n31984);
  and g54212 (n31985, n31973, n_22323);
  not g54213 (n_22324, n31985);
  and g54214 (n31986, n31973, n_22324);
  and g54215 (n31987, n_22323, n_22324);
  not g54216 (n_22325, n31986);
  not g54217 (n_22326, n31987);
  and g54218 (n31988, n_22325, n_22326);
  and g54219 (n31989, n_22268, n_22269);
  not g54220 (n_22327, n31989);
  and g54221 (n31990, n_22227, n_22327);
  not g54222 (n_22328, n31988);
  not g54223 (n_22329, n31990);
  and g54224 (n31991, n_22328, n_22329);
  not g54225 (n_22330, n31991);
  and g54226 (n31992, n_22328, n_22330);
  and g54227 (n31993, n_22329, n_22330);
  not g54228 (n_22331, n31992);
  not g54229 (n_22332, n31993);
  and g54230 (n31994, n_22331, n_22332);
  and g54231 (n31995, n_22274, n_22278);
  and g54232 (n31996, n31994, n31995);
  not g54233 (n_22333, n31994);
  not g54234 (n_22334, n31995);
  and g54235 (n31997, n_22333, n_22334);
  not g54236 (n_22335, n31996);
  not g54237 (n_22336, n31997);
  and g54238 (n31998, n_22335, n_22336);
  and g54239 (n31999, n_22282, n31998);
  not g54240 (n_22337, n31998);
  and g54241 (n32000, n31919, n_22337);
  or g54242 (\result[29] , n31999, n32000);
  and g54243 (n32002, n31919, n31998);
  and g54244 (n32003, n_22330, n_22336);
  and g54245 (n32004, n_22313, n_22324);
  and g54246 (n32005, n_22289, n_22292);
  and g54254 (n32013, n_22288, n32012);
  not g54255 (n_22338, n32012);
  and g54256 (n32014, n31945, n_22338);
  not g54257 (n_22339, n32005);
  not g54258 (n_22340, n32014);
  and g54259 (n32015, n_22339, n_22340);
  not g54260 (n_22341, n32013);
  and g54261 (n32016, n_22341, n32015);
  not g54262 (n_22342, n32016);
  and g54263 (n32017, n_22339, n_22342);
  and g54264 (n32018, n_22340, n_22342);
  and g54265 (n32019, n_22341, n32018);
  not g54266 (n_22343, n32017);
  not g54267 (n_22344, n32019);
  and g54268 (n32020, n_22343, n_22344);
  and g54269 (n32021, n75, n_18823);
  and g54270 (n32022, n3020, n26890);
  and g54271 (n32023, n3023, n26066);
  and g54272 (n32024, n3028, n26060);
  not g54280 (n_22349, n32020);
  not g54281 (n_22350, n32027);
  and g54282 (n32028, n_22349, n_22350);
  not g54283 (n_22351, n32028);
  and g54284 (n32029, n_22349, n_22351);
  and g54285 (n32030, n_22350, n_22351);
  not g54286 (n_22352, n32029);
  not g54287 (n_22353, n32030);
  and g54288 (n32031, n_22352, n_22353);
  and g54289 (n32032, n_22298, n_22309);
  and g54290 (n32033, n32031, n32032);
  not g54291 (n_22354, n32031);
  not g54292 (n_22355, n32032);
  and g54293 (n32034, n_22354, n_22355);
  not g54294 (n_22356, n32033);
  not g54295 (n_22357, n32034);
  and g54296 (n32035, n_22356, n_22357);
  and g54297 (n32036, n_17540, n_19417);
  and g54298 (n32037, n3967, n27964);
  not g54299 (n_22358, n32036);
  not g54300 (n_22359, n32037);
  and g54301 (n32038, n_22358, n_22359);
  and g54302 (n32039, n4050, n_19600);
  not g54303 (n_22360, n32039);
  and g54304 (n32040, n32038, n_22360);
  not g54305 (n_22361, n32040);
  and g54306 (n32041, \a[26] , n_22361);
  not g54307 (n_22362, n32041);
  and g54308 (n32042, n_22361, n_22362);
  and g54309 (n32043, \a[26] , n_22362);
  not g54310 (n_22363, n32042);
  not g54311 (n_22364, n32043);
  and g54312 (n32044, n_22363, n_22364);
  and g54313 (n32045, n3457, n27698);
  and g54314 (n32046, n3542, n27173);
  and g54315 (n32047, n3606, n27442);
  and g54321 (n32050, n3368, n_19446);
  not g54324 (n_22369, n32051);
  and g54325 (n32052, \a[29] , n_22369);
  not g54326 (n_22370, n32052);
  and g54327 (n32053, \a[29] , n_22370);
  and g54328 (n32054, n_22369, n_22370);
  not g54329 (n_22371, n32053);
  not g54330 (n_22372, n32054);
  and g54331 (n32055, n_22371, n_22372);
  not g54332 (n_22373, n32044);
  not g54333 (n_22374, n32055);
  and g54334 (n32056, n_22373, n_22374);
  not g54335 (n_22375, n32056);
  and g54336 (n32057, n_22373, n_22375);
  and g54337 (n32058, n_22374, n_22375);
  not g54338 (n_22376, n32057);
  not g54339 (n_22377, n32058);
  and g54340 (n32059, n_22376, n_22377);
  not g54341 (n_22378, n32035);
  and g54342 (n32060, n_22378, n32059);
  not g54343 (n_22379, n32059);
  and g54344 (n32061, n32035, n_22379);
  not g54345 (n_22380, n32060);
  not g54346 (n_22381, n32061);
  and g54347 (n32062, n_22380, n_22381);
  not g54348 (n_22382, n32004);
  and g54349 (n32063, n_22382, n32062);
  not g54350 (n_22383, n32062);
  and g54351 (n32064, n32004, n_22383);
  not g54352 (n_22384, n32063);
  not g54353 (n_22385, n32064);
  and g54354 (n32065, n_22384, n_22385);
  not g54355 (n_22386, n32003);
  and g54356 (n32066, n_22386, n32065);
  not g54357 (n_22387, n32065);
  and g54358 (n32067, n32003, n_22387);
  not g54359 (n_22388, n32066);
  not g54360 (n_22389, n32067);
  and g54361 (n32068, n_22388, n_22389);
  not g54362 (n_22390, n32002);
  not g54363 (n_22391, n32068);
  and g54364 (n32069, n_22390, n_22391);
  and g54365 (n32070, n32002, n32068);
  not g54366 (n_22392, n32069);
  not g54367 (n_22393, n32070);
  and g54368 (\result[30] , n_22392, n_22393);
  and g54369 (n32072, n_22384, n_22388);
  and g54370 (n32073, n3457, n27964);
  and g54371 (n32074, n3542, n27442);
  and g54372 (n32075, n3606, n27698);
  and g54378 (n32078, n3368, n27976);
  and g54381 (n32080, n_22351, n_22357);
  not g54382 (n_22398, n32080);
  and g54383 (n32081, \a[29] , n_22398);
  and g54384 (n32082, n_15, n32080);
  not g54385 (n_22399, n32081);
  not g54386 (n_22400, n32082);
  and g54387 (n32083, n_22399, n_22400);
  and g54388 (n32084, n32079, n32083);
  not g54389 (n_22401, n32079);
  not g54390 (n_22402, n32083);
  and g54391 (n32085, n_22401, n_22402);
  not g54392 (n_22403, n32084);
  not g54393 (n_22404, n32085);
  and g54394 (n32086, n_22403, n_22404);
  and g54395 (n32087, n75, n27185);
  and g54396 (n32088, n3020, n27173);
  and g54397 (n32089, n3023, n26060);
  and g54398 (n32090, n3028, n26890);
  not g54406 (n_22409, n32093);
  and g54407 (n32094, n32018, n_22409);
  not g54408 (n_22410, n32018);
  and g54409 (n32095, n_22410, n32093);
  not g54410 (n_22411, n32094);
  not g54411 (n_22412, n32095);
  and g54412 (n32096, n_22411, n_22412);
  not g54413 (n_22413, n32096);
  and g54414 (n32097, n32086, n_22413);
  not g54415 (n_22414, n32086);
  and g54416 (n32098, n_22414, n32096);
  not g54417 (n_22415, n32097);
  not g54418 (n_22416, n32098);
  and g54419 (n32099, n_22415, n_22416);
  and g54420 (n32100, n_22375, n_22381);
  and g54421 (n32101, n3874, n4511);
  and g54422 (n32102, n_242, n32101);
  not g54423 (n_22417, n32102);
  and g54424 (n32103, \a[26] , n_22417);
  and g54425 (n32104, n_33, n32102);
  not g54426 (n_22418, n32103);
  not g54427 (n_22419, n32104);
  and g54428 (n32105, n_22418, n_22419);
  and g54429 (n32106, n_17587, n_19417);
  not g54430 (n_22420, n32106);
  and g54431 (n32107, n31945, n_22420);
  and g54432 (n32108, n_22288, n32106);
  not g54433 (n_22421, n32107);
  not g54434 (n_22422, n32108);
  and g54435 (n32109, n_22421, n_22422);
  and g54436 (n32110, n32105, n32109);
  not g54437 (n_22423, n32105);
  not g54438 (n_22424, n32109);
  and g54439 (n32111, n_22423, n_22424);
  not g54440 (n_22425, n32110);
  not g54441 (n_22426, n32111);
  and g54442 (n32112, n_22425, n_22426);
  not g54443 (n_22427, n32112);
  and g54444 (n32113, n32100, n_22427);
  not g54445 (n_22428, n32100);
  and g54446 (n32114, n_22428, n32112);
  not g54447 (n_22429, n32113);
  not g54448 (n_22430, n32114);
  and g54449 (n32115, n_22429, n_22430);
  and g54450 (n32116, n32099, n32115);
  not g54451 (n_22431, n32099);
  not g54452 (n_22432, n32115);
  and g54453 (n32117, n_22431, n_22432);
  not g54454 (n_22433, n32116);
  not g54455 (n_22434, n32117);
  and g54456 (n32118, n_22433, n_22434);
  not g54457 (n_22435, n32072);
  not g54458 (n_22436, n32118);
  and g54459 (n32119, n_22435, n_22436);
  and g54460 (n32120, n32072, n32118);
  not g54461 (n_22437, n32119);
  not g54462 (n_22438, n32120);
  and g54463 (n32121, n_22437, n_22438);
  and g54464 (n32122, n32070, n32121);
  not g54465 (n_22439, n32121);
  and g54466 (n32123, n_22393, n_22439);
  or g54467 (\result[31] , n32122, n32123);
  nor g54468 (n26647, n26641, n26642, n26643, n26646);
  nor g54469 (n25296, n25288, n25289, n25290, n25295);
  nor g54470 (n22531, n22310, n22313, n22316, n22530);
  nor g54471 (n25317, n25308, n25309, n25310, n25316);
  nor g54472 (n26573, n26567, n26568, n26569, n26572);
  nor g54473 (n25335, n25329, n25330, n25331, n25334);
  nor g54474 (n26559, n26553, n26554, n26555, n26558);
  nor g54475 (n26008, n26002, n26003, n26004, n26005);
  nor g54476 (n26041, n26035, n26036, n26037, n26040);
  nor g54477 (n26855, n26849, n26850, n26851, n26852);
  nor g54478 (n25914, n25908, n25909, n25910, n25913);
  nor g54479 (n25973, n25967, n25968, n25969, n25972);
  nor g54480 (n24646, n24640, n24641, n24642, n24645);
  nor g54481 (n26659, n26653, n26654, n26655, n26658);
  nor g54482 (n25927, n25921, n25922, n25923, n25924);
  and g54483 (n_22472, n_123, n_207, n_159);
  and g54484 (n_22473, n1367, n2276, n25863);
  and g54485 (n_22474, n1601, n3405, n3764);
  and g54486 (n_22475, n3432, n792, n13063);
  and g54487 (n25874, n_22472, n_22473, n_22474, n_22475);
  nor g54488 (n25884, n25878, n25879, n25880, n25881);
  nor g54489 (n22544, n22536, n22537, n22538, n22543);
  nor g54490 (n24663, n24657, n24658, n24659, n24662);
  nor g54491 (n25381, n25375, n25376, n25377, n25380);
  nor g54492 (n25102, n25096, n25097, n25098, n25101);
  and g54493 (n26859, n_148, n26016, n4030, n4511);
  nor g54494 (n22231, n22225, n22226, n22227, n22230);
  nor g54495 (n22246, n22240, n22241, n22242, n22243);
  and g54496 (n_22476, n_85, n_99, n_242, n_58);
  and g54497 (n_22477, n_123, n_262, n3757, n2170);
  and g54498 (n_22478, n1731, n13063, n3782);
  and g54499 (n_22479, n3978, n473, n1047);
  and g54500 (n25940, n_22476, n_22477, n_22478, n_22479);
  and g54501 (n_22480, n_94, n_294);
  and g54502 (n_22481, n_192, n_244);
  and g54503 (n_22482, n3886, n1824);
  and g54504 (n_22483, n774, n6716);
  and g54505 (n25863, n_22480, n_22481, n_22482, n_22483);
  and g54506 (n_22484, n_276, n_145, n_194, n_197);
  and g54507 (n_22485, n_46, n_243, n291);
  and g54508 (n_22486, n3386, n3389, n3391);
  and g54509 (n_22487, n3393, n1392, n1739);
  and g54510 (n3405, n_22484, n_22485, n_22486, n_22487);
  and g54511 (n_22488, n_228, n_185);
  and g54512 (n_22489, n_143, n_202);
  and g54513 (n_22490, n_65, n_75);
  and g54514 (n_22491, n_245, n2293);
  and g54515 (n3764, n_22488, n_22489, n_22490, n_22491);
  and g54516 (n_22492, n_209, n_76);
  and g54517 (n_22493, n_173, n_87, n_128, n_49);
  and g54518 (n_22494, n720, n1182, n873, n1528);
  and g54519 (n_22495, n3408, n3415, n1132, n1388);
  and g54520 (n_22496, n3266, n1045, n3416, n_22492);
  and g54521 (n3432, n_22493, n_22494, n_22495, n_22496);
  and g54522 (n_22497, n_191, n_259);
  and g54523 (n13063, n3984, n1255, n1781, n_22497);
  nor g54524 (n24169, n24160, n24161, n24162, n24168);
  nor g54525 (n25398, n25392, n25393, n25394, n25397);
  nor g54526 (n26491, n26485, n26486, n26487, n26490);
  nor g54527 (n14030, n14022, n14023, n14024, n14029);
  nor g54528 (n22292, n22286, n22287, n22288, n22291);
  and g54529 (n_22498, n_78, n_213, n_69, n_284);
  and g54530 (n_22499, n_211, n_196, n_262, n_38);
  and g54531 (n_22500, n_68, n_48, n3947);
  and g54532 (n_22501, n3128, n3914, n3931);
  and g54533 (n4030, n_22498, n_22499, n_22500, n_22501);
  and g54534 (n_22502, n_201, n_259, n_133);
  and g54535 (n_22503, n1367, n1761, n1046);
  and g54536 (n_22504, n2346, n4493);
  and g54537 (n_22505, n133, n4502);
  and g54538 (n4511, n_22502, n_22503, n_22504, n_22505);
  nor g54539 (n13591, n13585, n13586, n13587, n13588);
  and g54540 (n_22506, n_189, n_81, n_57, n_212);
  and g54541 (n_22507, n_271, n1367, n515, n1141);
  and g54542 (n_22508, n720, n2582, n3733, n3739);
  and g54543 (n_22509, n3743, n401, n2556);
  and g54544 (n3757, n_22506, n_22507, n_22508, n_22509);
  and g54545 (n_22510, n_204, n_133);
  and g54546 (n1731, n_181, n_68, n1727, n_22510);
  and g54547 (n_22511, n_183, n_136, n_151);
  and g54548 (n_22512, n_234, n_278, n_241);
  and g54549 (n_22513, n_131, n872, n2512);
  and g54550 (n_22514, n3768, n1784, n3771);
  and g54551 (n3782, n_22511, n_22512, n_22513, n_22514);
  and g54552 (n_22515, n_238, n_194);
  and g54553 (n_22516, n_274, n_94);
  and g54554 (n_22517, n_244, n2470);
  and g54555 (n3978, n3832, n_22515, n_22516, n_22517);
  and g54556 (n_22518, n_72, n_258);
  and g54557 (n_22519, n_227, n_195);
  and g54558 (n_22520, n_212, n_126);
  and g54559 (n3386, n3380, n_22518, n_22519, n_22520);
  and g54560 (n3389, n_177, n_50, n_297, n2508);
  and g54561 (n3408, n_40, n_263, n_254, n2073);
  and g54562 (n_22521, n_274, n_66);
  and g54563 (n_22522, n_216, n_287);
  and g54564 (n_22523, n3409, n300);
  and g54565 (n3415, n962, n_22521, n_22522, n_22523);
  and g54566 (n_22524, n_117, n_36);
  and g54567 (n_22525, n_264, n_167);
  and g54568 (n_22526, n_149, n1478);
  and g54569 (n3984, n1726, n_22524, n_22525, n_22526);
  nor g54570 (n24190, n24181, n24182, n24183, n24189);
  and g54571 (n_22527, n_191, n968);
  and g54572 (n3873, n1480, n3570, n3869, n_22527);
  and g54573 (n_22528, n_189, n_223);
  and g54574 (n3972, n_181, n_209, n_208, n_22528);
  and g54575 (n_22529, n_212, n_289, n_188);
  and g54576 (n_22530, n_60, n_131);
  and g54577 (n_22531, n1292, n3409);
  and g54578 (n_22532, n1440, n3729);
  and g54579 (n3947, n_22529, n_22530, n_22531, n_22532);
  and g54580 (n_22533, n_75, n_198);
  and g54581 (n_22534, n_83, n_98);
  and g54582 (n4493, n_265, n2014, n_22533, n_22534);
  and g54583 (n_22535, n_166, n_52, n_129);
  and g54584 (n_22536, n_234, n_84, n_58);
  and g54585 (n_22537, n2170, n604);
  and g54586 (n_22538, n1388, n1785);
  and g54587 (n4502, n_22535, n_22536, n_22537, n_22538);
  and g54588 (n_22539, n_242, n_148);
  and g54589 (n_22540, n26016, n2740);
  and g54590 (n26021, n4017, n4040, n_22539, n_22540);
  and g54591 (n13059, n_192, n193, n3831, n13056);
  and g54592 (n_22541, n_233, n_205);
  and g54593 (n3733, n_80, n_59, n3729, n_22541);
  and g54594 (n_22542, n_246, n_108);
  and g54595 (n_22543, n_225, n_263);
  and g54596 (n_22544, n_254, n_226);
  and g54597 (n3739, n1839, n_22542, n_22543, n_22544);
  and g54598 (n_22545, n_92, n_79);
  and g54599 (n3743, n_48, n640, n895, n_22545);
  and g54600 (n872, n_130, n_267, n_51, n_105);
  and g54601 (n_22546, n_214, n_120);
  and g54602 (n2512, n_184, n642, n2508, n_22546);
  and g54603 (n_22547, n_218, n_40);
  and g54604 (n3768, n590, n1392, n3115, n_22547);
  and g54605 (n3771, n_231, n_285, n_180, n747);
  and g54606 (n_22548, n_137, n_53);
  and g54607 (n_22549, n_129, n_87, n_160, n_272);
  and g54608 (n_22550, n1269, n3733, n471, n774);
  and g54609 (n_22551, n14534, n13787, n16031, n4827);
  and g54610 (n_22552, n6567, n303, n3042, n_22548);
  and g54611 (n22268, n_22549, n_22550, n_22551, n_22552);
  nor g54612 (n25416, n25410, n25411, n25412, n25415);
  nor g54613 (n26477, n26471, n26472, n26473, n26476);
  nor g54614 (n13656, n13628, n13631, n13634, n13655);
  nor g54615 (n13931, n13923, n13924, n13925, n13930);
  and g54616 (n3869, n_137, n_247, n3858, n3866);
  and g54617 (n_22553, n_170, n_174);
  and g54618 (n_22554, n_297, n_200);
  and g54619 (n_22555, n_47, n_93);
  and g54620 (n3912, n_126, n_22553, n_22554, n_22555);
  and g54621 (n_22556, n_193, n421);
  and g54622 (n_22557, n1783, n4003);
  and g54623 (n_22558, n4009, n3408);
  and g54624 (n4017, n4011, n_22556, n_22557, n_22558);
  and g54625 (n_22559, n_44, n159);
  and g54626 (n_22560, n1046, n604);
  and g54627 (n_22561, n3790, n1204);
  and g54628 (n4040, n3852, n_22559, n_22560, n_22561);
  and g54629 (n_22562, n_180, n_268);
  and g54630 (n3831, n_99, n3437, n3827, n_22562);
  and g54631 (n_22563, n_292, n_289, n341, n1389);
  and g54632 (n_22564, n826, n1139, n291, n1029);
  and g54633 (n_22565, n13031, n1521, n13041, n12828);
  and g54634 (n_22566, n6607, n593, n2020, n6664);
  and g54635 (n13056, n_22563, n_22564, n_22565, n_22566);
  and g54636 (n_22567, n_182, n_277);
  and g54637 (n_22568, n_177, n_178);
  and g54638 (n_22569, n_239, n887);
  and g54639 (n895, n889, n_22567, n_22568, n_22569);
  and g54640 (n_22570, n_161, n_227, n_116, n_56);
  and g54641 (n_22571, n_272, n3886, n896, n2021);
  and g54642 (n_22572, n4293, n13560, n12939, n3389);
  and g54643 (n_22573, n12390, n3549, n5734);
  and g54644 (n13574, n_22570, n_22571, n_22572, n_22573);
  and g54645 (n_22574, n_202, n_257, n_258);
  and g54646 (n_22575, n_138, n_269, n_288);
  and g54647 (n_22576, n3409, n1070);
  and g54648 (n_22577, n343, n13700);
  and g54649 (n14534, n_22574, n_22575, n_22576, n_22577);
  and g54650 (n_22578, n_277, n_135, n_167, n_101);
  and g54651 (n_22579, n_184, n_207, n_90, n_254);
  and g54652 (n_22580, n1366, n6020, n4325);
  and g54653 (n_22581, n13773, n3160, n13774);
  and g54654 (n13787, n_22578, n_22579, n_22580, n_22581);
  and g54655 (n_22582, n_182, n_121, n_181);
  and g54656 (n_22583, n_149, n_38, n731);
  and g54657 (n_22584, n1480, n808, n877);
  and g54658 (n_22585, n1103, n1409, n16020);
  and g54659 (n16031, n_22582, n_22583, n_22584, n_22585);
  and g54660 (n_22586, n_235, n_100, n_119);
  and g54661 (n_22587, n_284, n570);
  and g54662 (n_22588, n1726, n4819);
  and g54663 (n_22589, n2584, n2721);
  and g54664 (n4827, n_22586, n_22587, n_22588, n_22589);
  nor g54665 (n14687, n14681, n14682, n14683, n14686);
  nor g54666 (n14138, n14130, n14131, n14132, n14137);
  nor g54667 (n13978, n13970, n13971, n13972, n13977);
  and g54668 (n_22590, n_225, n_115, n_118);
  and g54669 (n_22591, n356, n979);
  and g54670 (n_22592, n1254, n2963);
  and g54671 (n_22593, n624, n3206);
  and g54672 (n3866, n_22590, n_22591, n_22592, n_22593);
  and g54673 (n_22594, n_164, n_114);
  and g54674 (n_22595, n_120, n_184);
  and g54675 (n_22596, n538, n3990);
  and g54676 (n4003, n3997, n_22594, n_22595, n_22596);
  and g54677 (n_22597, n_37, n_210);
  and g54678 (n_22598, n1389, n1248);
  and g54679 (n_22599, n2739, n2133);
  and g54680 (n4009, n2703, n_22597, n_22598, n_22599);
  and g54681 (n_22600, n_168, n_290, n_251);
  and g54682 (n_22601, n_220, n_86);
  and g54683 (n_22602, n_45, n_227);
  and g54684 (n_22603, n1388, n1577);
  and g54685 (n3790, n_22600, n_22601, n_22602, n_22603);
  and g54686 (n_22604, n_41, n_204);
  and g54687 (n3852, n128, n2208, n2573, n_22604);
  and g54688 (n_22605, n_185, n_224, n_167, n_39);
  and g54689 (n_22606, n_111, n_126, n1248, n1827);
  and g54690 (n_22607, n2507, n2782, n1511, n12795);
  and g54691 (n_22608, n13012, n1693, n13014, n13016);
  and g54692 (n13031, n_22605, n_22606, n_22607, n_22608);
  and g54693 (n_22609, n_266, n_135, n_96);
  and g54694 (n_22610, n_270, n_132, n_57);
  and g54695 (n_22611, n_149, n_273, n_48);
  and g54696 (n_22612, n_159, n960);
  and g54697 (n1521, n_22609, n_22610, n_22611, n_22612);
  and g54698 (n_22613, n_121, n_256, n_62);
  and g54699 (n_22614, n_218, n_177, n_239);
  and g54700 (n_22615, n_252, n591, n897);
  and g54701 (n_22616, n1556, n4151);
  and g54702 (n13041, n_22613, n_22614, n_22615, n_22616);
  and g54703 (n_22617, n_182, n_136);
  and g54704 (n_22618, n_214, n_98, n_127, n_117);
  and g54705 (n_22619, n_172, n_49, n_95, n_106);
  and g54706 (n_22620, n_69, n202, n4794, n12805);
  and g54707 (n_22621, n12810, n1527, n12812, n_22617);
  and g54708 (n12828, n_22618, n_22619, n_22620, n_22621);
  and g54709 (n6607, n_201, n_175, n_148, n515);
  and g54710 (n2020, n_163, n_81, n_153, n_211);
  and g54711 (n_22622, n_163, n_72, n_280, n_36);
  and g54712 (n_22623, n_82, n_128, n_111, n1237);
  and g54713 (n_22624, n773, n1917, n4274, n4215);
  and g54714 (n_22625, n4279, n1944, n2684);
  and g54715 (n4293, n_22622, n_22623, n_22624, n_22625);
  and g54716 (n_22626, n_42, n_136, n_199);
  and g54717 (n_22627, n_244, n_288, n_170);
  and g54718 (n_22628, n285, n3544, n2371);
  and g54719 (n_22629, n989, n3792, n4788);
  and g54720 (n13560, n_22626, n_22627, n_22628, n_22629);
  and g54722 (n_22631, n_47, n2443);
  and g54723 (n_22632, n12924, n12932);
  and g54724 (n_22633, n640, n5040);
  and g54725 (n12939, n_22630, n_22631, n_22632, n_22633);
  and g54726 (n12390, n_75, n_160, n_207, n508);
  and g54727 (n_22634, n_240, n_234);
  and g54728 (n_22635, n_157, n_245);
  and g54729 (n6020, n_118, n2059, n_22634, n_22635);
  and g54730 (n_22636, n_268, n_124, n_189, n_150);
  and g54731 (n_22637, n_267, n_175, n_239);
  and g54732 (n_22638, n_49, n_244, n_50);
  and g54733 (n_22639, n1602, n941, n4313);
  and g54734 (n4325, n_22636, n_22637, n_22638, n_22639);
  and g54735 (n_22640, n_219, n_116);
  and g54736 (n_22641, n_241, n_263);
  and g54737 (n13773, n_243, n_297, n_22640, n_22641);
  and g54738 (n808, n_166, n_180, n_123, n_209);
  and g54739 (n_22642, n_256, n_72);
  and g54740 (n4819, n_221, n_63, n_226, n_22642);
  nor g54741 (n26460, n26454, n26455, n26456, n26459);
  nor g54742 (n12902, n12896, n12897, n12898, n12899);
  nor g54743 (n13507, n13492, n13493, n13494, n13504);
  and g54744 (n3990, n_175, n_51, n1347, n3987);
  and g54745 (n_22643, n_87, n_128);
  and g54746 (n_22644, n_172, n_108);
  and g54747 (n_22645, n_239, n_80);
  and g54748 (n_22646, n1916, n2297);
  and g54749 (n3997, n_22643, n_22644, n_22645, n_22646);
  and g54750 (n_22647, n_101, n_91);
  and g54751 (n_22648, n_142, n_215);
  and g54752 (n2703, n_232, n_269, n_22647, n_22648);
  and g54753 (n_22630, n_155, n_277);
  and g54754 (n_22650, n_34, n_136);
  and g54755 (n_22651, n_224, n720);
  and g54756 (n2208, n1531, n_22630, n_22650, n_22651);
  and g54757 (n_22652, n_83, n_160);
  and g54758 (n2782, n_188, n566, n1727, n_22652);
  and g54759 (n_22653, n_137, n_231, n_251, n_58);
  and g54760 (n_22654, n_140, n_241, n1478);
  and g54761 (n_22655, n1479, n1480, n1488);
  and g54762 (n_22656, n1496, n1497, n1499);
  and g54763 (n1511, n_22653, n_22654, n_22655, n_22656);
  and g54764 (n_22657, n_92, n_274, n_86);
  and g54765 (n_22658, n_134, n_280, n_197);
  and g54766 (n_22659, n_131, n2582, n2573);
  and g54767 (n_22660, n653, n12785);
  and g54768 (n12795, n_22657, n_22658, n_22659, n_22660);
  and g54769 (n13012, n_41, n_215, n_59, n238);
  and g54770 (n4151, n_71, n_277, n_60, n_294);
  and g54771 (n_22661, n_65, n_91);
  and g54772 (n_22662, n_70, n_174);
  and g54773 (n_22663, n_297, n2154);
  and g54774 (n4794, n4788, n_22661, n_22662, n_22663);
  and g54775 (n_22664, n_290, n_220, n_257);
  and g54776 (n_22665, n_76, n1247, n282);
  and g54777 (n_22666, n2170, n968, n1476);
  and g54778 (n_22667, n561, n5808);
  and g54779 (n12805, n_22664, n_22665, n_22666, n_22667);
  and g54780 (n_22668, n_42, n_194);
  and g54781 (n_22669, n_288, n_78);
  and g54782 (n12810, n_196, n_254, n_22668, n_22669);
  and g54783 (n1527, n_204, n_240, n_61, n1524);
  and g54784 (n_22670, n_213, n_97, n2583);
  and g54785 (n_22671, n2738, n3848, n4502);
  and g54786 (n_22672, n13063, n4017, n5233);
  and g54787 (n_22673, n3580, n2265, n3906);
  and g54788 (n13074, n_22670, n_22671, n_22672, n_22673);
  and g54789 (n_22674, n_233, n_222);
  and g54790 (n_22675, n_148, n3869);
  and g54791 (n_22676, n13075, n3832);
  and g54792 (n13081, n4034, n_22674, n_22675, n_22676);
  and g54793 (n_22677, n_183, n_181);
  and g54794 (n_22678, n_172, n_263);
  and g54795 (n4274, n250, n4269, n_22677, n_22678);
  and g54796 (n_22679, n_191, n_158);
  and g54797 (n_22680, n_34, n2090);
  and g54798 (n_22681, n977, n2348);
  and g54799 (n4215, n2515, n_22679, n_22680, n_22681);
  and g54800 (n_22682, n_279, n_54);
  and g54801 (n_22683, n_190, n_173);
  and g54802 (n4279, n_131, n_178, n_22682, n_22683);
  and g54803 (n_22684, n_121, n_233);
  and g54804 (n_22685, n_242, n_270);
  and g54805 (n12924, n_95, n2092, n_22684, n_22685);
  and g54806 (n_22686, n_168, n_176, n_81);
  and g54807 (n_22687, n_149, n_97);
  and g54808 (n_22688, n_38, n1782);
  and g54809 (n_22689, n1994, n6520);
  and g54810 (n12932, n_22686, n_22687, n_22688, n_22689);
  nor g54811 (n14123, n14117, n14118, n14119, n14122);
  nor g54812 (n14298, n14292, n14293, n14294, n14297);
  nor g54813 (n14793, n14787, n14788, n14789, n14792);
  nor g54814 (n13911, n13902, n13903, n13904, n13910);
  nor g54815 (n13311, n13305, n13306, n13307, n13308);
  and g54816 (n_22690, n_53, n_285, n_199);
  and g54817 (n_22691, n_45, n_234);
  and g54818 (n_22692, n_264, n_115);
  and g54819 (n_22693, n253, n1384);
  and g54820 (n1488, n_22690, n_22691, n_22692, n_22693);
  and g54821 (n_22694, n_43, n_122);
  and g54822 (n_22695, n_52, n_138);
  and g54823 (n_22696, n_278, n_184);
  and g54824 (n1496, n1490, n_22694, n_22695, n_22696);
  and g54825 (n_22697, n_108, n_80, n_170);
  and g54826 (n_22698, n618, n621, n622);
  and g54827 (n_22699, n631, n632, n636);
  and g54828 (n_22700, n638, n640, n642);
  and g54829 (n653, n_22697, n_22698, n_22699, n_22700);
  and g54830 (n561, n_110, n_87, n_225, n_226);
  and g54831 (n_22701, n_292, n_139, n_110);
  and g54832 (n_22702, n_238, n_104, n_251);
  and g54833 (n_22703, n827, n471);
  and g54834 (n_22704, n772, n1105);
  and g54835 (n3848, n_22701, n_22702, n_22703, n_22704);
  and g54836 (n_22705, n_169, n_219, n_274);
  and g54837 (n_22706, n_44, n_124, n_146);
  and g54838 (n_22707, n1367, n1155);
  and g54839 (n_22708, n1085, n2752);
  and g54840 (n5233, n_22705, n_22706, n_22707, n_22708);
  and g54841 (n_22709, n_145, n_144, n_45);
  and g54842 (n_22710, n_222, n_227, n_196);
  and g54843 (n_22711, n3569, n2348, n2013);
  and g54844 (n_22712, n2267, n3570);
  and g54845 (n3580, n_22709, n_22710, n_22711, n_22712);
  and g54846 (n_22713, n_35, n_270);
  and g54847 (n4034, n3984, n4017, n4030, n_22713);
  and g54848 (n2515, n_92, n_273, n_90, n282);
  and g54849 (n6520, n_137, n_52, n_48, n_213);
  nor g54850 (n14339, n14333, n14334, n14335, n14338);
  nor g54851 (n13995, n13989, n13990, n13991, n13994);
  nor g54852 (n14010, n14004, n14005, n14006, n14009);
  nor g54853 (n23674, n23666, n23667, n23668, n23673);
  nor g54854 (n24236, n24230, n24231, n24232, n24235);
  and g54855 (n_22714, n_259, n_123);
  and g54856 (n1384, n_152, n_89, n1380, n_22714);
  and g54857 (n_22715, n_168, n_219);
  and g54858 (n_22716, n_246, n_63);
  and g54859 (n_22717, n_101, n_79);
  and g54860 (n_22718, n_141, n624);
  and g54861 (n631, n_22715, n_22716, n_22717, n_22718);
  and g54862 (n_22719, n_205, n_267);
  and g54863 (n3569, n_154, n_207, n_244, n_22719);
  nor g54864 (n14107, n14101, n14102, n14103, n14106);
  nor g54865 (n23691, n23685, n23686, n23687, n23690);
  nor g54866 (n24253, n24247, n24248, n24249, n24252);
  nor g54867 (n13006, n13000, n13001, n13002, n13003);
  and g54868 (n_22720, n_167, n_120, n_105, n_146);
  and g54869 (n_22721, n4295, n1129, n12909, n12919);
  and g54870 (n_22722, n2623, n12939, n12944, n2468);
  and g54871 (n_22723, n1249, n638, n2230);
  and g54872 (n12958, n_22720, n_22721, n_22722, n_22723);
  nor g54873 (n13740, n13731, n13732, n13733, n13737);
  and g54874 (n_22724, n_35, n_257, n_242);
  and g54875 (n_22725, n1761, n665);
  and g54876 (n_22726, n4493, n3856);
  and g54877 (n_22727, n3949, n13087);
  and g54878 (n13095, n_22724, n_22725, n_22726, n_22727);
  nor g54879 (n13332, n13326, n13327, n13328, n13329);
  nor g54880 (n14167, n14161, n14162, n14163, n14166);
  nor g54881 (n15194, n15188, n15189, n15190, n15193);
  nor g54882 (n24723, n24717, n24718, n24719, n24722);
  and g54883 (n_22728, n_228, n_94);
  and g54884 (n_22729, n_166, n6706);
  and g54885 (n_22730, n_100, n_207);
  and g54886 (n_22731, n_153, n_97, n1252, n1825);
  and g54887 (n_22732, n2633, n1523, n12973, n1969);
  and g54888 (n_22733, n5224, n1216, n12977, n3985);
  and g54889 (n_22734, n4334, n_22728, n_22729, n_22730);
  and g54890 (n12995, n_22731, n_22732, n_22733, n_22734);
  and g54891 (n_22735, n_45, n_180);
  and g54892 (n_22736, n_193, n_175);
  and g54893 (n_22737, n_291, n_69);
  and g54894 (n_22738, n_131, n_254);
  and g54895 (n12909, n_22735, n_22736, n_22737, n_22738);
  and g54896 (n_22739, n_71, n_145, n_279);
  and g54897 (n_22740, n_290, n_172);
  and g54898 (n_22741, n_51, n12911);
  and g54899 (n_22742, n1611, n4327);
  and g54900 (n12919, n_22739, n_22740, n_22741, n_22742);
  and g54901 (n_22743, n_257, n_190, n_40, n_157);
  and g54902 (n_22744, n_60, n_159, n2582, n2583);
  and g54903 (n_22745, n1602, n2591, n2605, n790);
  and g54904 (n_22746, n595, n2607, n1800, n2608);
  and g54905 (n2623, n_22743, n_22744, n_22745, n_22746);
  and g54906 (n12944, n_228, n1237, n373, n12941);
  nor g54907 (n26671, n26665, n26666, n26667, n26670);
  and g54908 (n_22747, n_231, n_168);
  and g54909 (n3856, n3848, n2275, n3852, n_22747);
  and g54910 (n_22748, n_193, n968);
  and g54911 (n13087, n539, n3570, n3832, n_22748);
  and g54912 (n_22749, n_259, n471);
  and g54913 (n_22750, n3972, n3978);
  and g54914 (n4045, n4034, n4040, n_22749, n_22750);
  and g54915 (n3877, n_123, n_148, n3839, n3874);
  nor g54916 (n14669, n14663, n14664, n14665, n14668);
  nor g54917 (n24010, n24004, n24005, n24006, n24009);
  nor g54918 (n14780, n14774, n14775, n14776, n14779);
  nor g54919 (n14927, n14921, n14922, n14923, n14926);
  nor g54920 (n24271, n24265, n24266, n24267, n24270);
  nor g54921 (n24740, n24734, n24735, n24736, n24739);
  and g54922 (n_22751, n_139, n_86, n_234, n_283);
  and g54923 (n_22752, n_248, n_51, n_244, n_272);
  and g54924 (n_22753, n1161, n1827, n1254, n789);
  and g54925 (n_22754, n1925, n530, n2684, n3438);
  and g54926 (n12973, n_22751, n_22752, n_22753, n_22754);
  and g54927 (n_22755, n_155, n_217, n_176);
  and g54928 (n_22756, n_160, n_243, n896);
  and g54929 (n_22757, n1183, n512);
  and g54930 (n_22758, n772, n1960);
  and g54931 (n1969, n_22755, n_22756, n_22757, n_22758);
  and g54932 (n_22759, n_231, n_202, n_290, n_246);
  and g54933 (n_22760, n_58, n_61, n_177, n_245);
  and g54934 (n_22761, n_38, n5199, n5209, n1131);
  and g54935 (n_22762, n1024, n593, n2297, n4313);
  and g54936 (n5224, n_22759, n_22760, n_22761, n_22762);
  and g54937 (n_22763, n_259, n_138);
  and g54938 (n_22764, n_36, n_171);
  and g54939 (n1216, n_50, n_105, n_22763, n_22764);
  and g54940 (n_22765, n_92, n_195);
  and g54941 (n12977, n_70, n_113, n_188, n_22765);
  and g54942 (n_22766, n_276, n_266);
  and g54943 (n_22767, n_231, n_279, n_104, n_106);
  and g54944 (n_22768, n_225, n869, n450, n621);
  and g54945 (n_22769, n1708, n13458, n805, n988);
  and g54946 (n_22770, n2806, n694, n3192, n_22766);
  and g54947 (n13474, n_22767, n_22768, n_22769, n_22770);
  and g54948 (n_22771, n_292, n_143);
  and g54949 (n_22772, n_230, n_108);
  and g54950 (n_22773, n_56, n_272);
  and g54951 (n_22774, n2090, n2584);
  and g54952 (n2591, n_22771, n_22772, n_22773, n_22774);
  and g54953 (n_22775, n_169, n_219, n_86);
  and g54954 (n_22776, n_184, n_215, n_39);
  and g54955 (n_22777, n977, n1839, n2349);
  and g54956 (n_22778, n2593, n2595);
  and g54957 (n2605, n_22775, n_22776, n_22777, n_22778);
  nor g54958 (n25114, n25108, n25109, n25110, n25113);
  and g54959 (n_22779, n_121, n_217, n_233);
  and g54960 (n_22780, n1046, n4009, n13063);
  and g54961 (n_22781, n3947, n13087, n13161);
  and g54962 (n_22782, n1249, n1425, n1740);
  and g54963 (n13172, n_22779, n_22780, n_22781, n_22782);
  and g54964 (n_22783, n_164, n_35);
  and g54965 (n_22784, n193, n454);
  and g54966 (n_22785, n539, n665);
  and g54967 (n_22786, n3831, n3832);
  and g54968 (n3839, n_22783, n_22784, n_22785, n_22786);
  and g54969 (n4514, n_242, n_123, n3972, n4511);
  and g54970 (n_22787, n_256, n_217);
  and g54971 (n_22788, n_133, n_120);
  and g54972 (n_22789, n_160, n_115);
  and g54973 (n_22790, n_272, n_48);
  and g54974 (n_22791, n978, n2466);
  and g54975 (n_22792, n1252, n730, n1366, n2635);
  and g54976 (n_22793, n5085, n13123, n1202, n1735);
  and g54977 (n_22794, n13138, n1163, n2544, n_22787);
  and g54978 (n_22795, n_22788, n_22789, n_22790, n_22791);
  and g54979 (n13158, n_22792, n_22793, n_22794, n_22795);
  nor g54980 (n22558, n22549, n22550, n22551, n22557);
  and g54981 (n_22796, n_130, n_104, n_45);
  and g54982 (n_22797, n_261, n_127);
  and g54983 (n_22798, n_269, n_147);
  and g54984 (n_22799, n_273, n_287);
  and g54985 (n1925, n_22796, n_22797, n_22798, n_22799);
  and g54986 (n_22800, n_277, n_162);
  and g54987 (n_22801, n_240, n_282);
  and g54988 (n_22802, n_257, n_150);
  and g54989 (n5199, n2240, n_22800, n_22801, n_22802);
  and g54990 (n_22803, n_253, n_164, n_98);
  and g54991 (n_22804, n_186, n_79);
  and g54992 (n_22805, n_89, n_262);
  and g54993 (n_22806, n_93, n5201);
  and g54994 (n5209, n_22803, n_22804, n_22805, n_22806);
  and g54995 (n1024, n_102, n_205, n_91, n1021);
  and g54996 (n_22807, n_143, n_164, n_117);
  and g54997 (n_22808, n_60, n1667, n1679);
  and g54998 (n_22809, n1687, n1691, n1692);
  and g54999 (n_22810, n778, n1695, n1697);
  and g55000 (n1708, n_22807, n_22808, n_22809, n_22810);
  and g55001 (n_22811, n_229, n_274, n_115, n_90);
  and g55002 (n_22812, n_89, n1252, n294, n241);
  and g55003 (n_22813, n1245, n1894, n3435);
  and g55004 (n_22814, n2595, n336, n5002);
  and g55005 (n13458, n_22811, n_22812, n_22813, n_22814);
  and g55006 (n_22815, n_58, n_67);
  and g55007 (n_22816, n_283, n_40);
  and g55008 (n_22817, n_142, n515);
  and g55009 (n988, n982, n_22815, n_22816, n_22817);
  and g55010 (n_22818, n_253, n_43, n_217);
  and g55011 (n_22819, n_44, n_81, n_211);
  and g55012 (n_22820, n_287, n654, n1426);
  and g55013 (n_22821, n1025, n1602);
  and g55014 (n2806, n_22818, n_22819, n_22820, n_22821);
  and g55015 (n_22822, n_137, n_235, n_149, n_47);
  and g55016 (n_22823, n1380, n202, n2406, n1575);
  and g55017 (n_22824, n2605, n4815, n12919, n13698);
  and g55018 (n_22825, n13138, n6672, n2753, n13700);
  and g55019 (n13715, n_22822, n_22823, n_22824, n_22825);
  and g55020 (n_22826, n_185, n_274);
  and g55021 (n_22827, n_246, n1155);
  and g55022 (n_22828, n535, n2265);
  and g55023 (n2273, n2267, n_22826, n_22827, n_22828);
  and g55024 (n13161, n_84, n885, n3929, n5064);
  nor g55025 (n13296, n13290, n13291, n13292, n13293);
  and g55026 (n_22829, n_54, n_193);
  and g55027 (n_22830, n_224, n_209);
  and g55028 (n_22831, n_230, n_264, n_107, n1531);
  and g55029 (n_22832, n1254, n4232, n6707, n13210);
  and g55030 (n_22833, n13221, n2987, n494, n624);
  and g55031 (n_22834, n3115, n5787, n_22829, n_22830);
  and g55032 (n13238, n_22831, n_22832, n_22833, n_22834);
  and g55033 (n_22835, n_144, n_114, n_222, n_192);
  and g55034 (n_22836, n_283, n_284, n720, n2583);
  and g55035 (n_22837, n520, n1046, n3929, n3939);
  and g55036 (n_22838, n2740, n3947, n1155, n3949);
  and g55037 (n3964, n_22835, n_22836, n_22837, n_22838);
  and g55038 (n_22839, n_144, n_235);
  and g55039 (n_22840, n_233, n_116);
  and g55040 (n_22841, n_82, n_153);
  and g55041 (n_22842, n722, n723);
  and g55042 (n730, n_22839, n_22840, n_22841, n_22842);
  and g55043 (n5085, n_206, n_44, n_124, n_270);
  and g55044 (n_22843, n_121, n_42, n_214);
  and g55045 (n_22844, n_100, n_173, n_128);
  and g55046 (n_22845, n1916, n4216);
  and g55047 (n_22846, n12397, n13114);
  and g55048 (n13123, n_22843, n_22844, n_22845, n_22846);
  and g55049 (n_22847, n_253, n_240);
  and g55050 (n_22848, n_222, n_63);
  and g55051 (n_22849, n_58, n_278, n_107, n_152);
  and g55052 (n_22850, n_38, n_47, n_126, n1182);
  and g55053 (n_22851, n1183, n787, n1155, n751);
  and g55054 (n_22852, n675, n1185, n_22847, n_22848);
  and g55055 (n1202, n_22849, n_22850, n_22851, n_22852);
  and g55056 (n1735, n_191, n_64, n_174, n1732);
  and g55057 (n13138, n_53, n_62, n_61, n13135);
  nor g55058 (n14280, n14274, n14275, n14276, n14279);
  nor g55059 (n14089, n14083, n14084, n14085, n14088);
  nor g55060 (n13755, n13749, n13750, n13751, n13752);
  nor g55061 (n23347, n23338, n23339, n23340, n23346);
  nor g55062 (n14764, n14758, n14759, n14760, n14763);
  nor g55063 (n14968, n14962, n14963, n14964, n14967);
  nor g55064 (n25476, n25470, n25471, n25472, n25475);
  and g55065 (n2240, n_64, n_223, n_157, n_179);
  and g55066 (n_22853, n_92, n_220, n_259);
  and g55067 (n_22854, n_189, n_261, n_38);
  and g55068 (n_22855, n1668, n1475, n933);
  and g55069 (n_22856, n849, n1669);
  and g55070 (n1679, n_22853, n_22854, n_22855, n_22856);
  and g55071 (n_22857, n_119, n_184);
  and g55072 (n_22858, n_239, n_159);
  and g55073 (n_22859, n790, n303);
  and g55074 (n1687, n1681, n_22857, n_22858, n_22859);
  and g55075 (n_22860, n_235, n_242);
  and g55076 (n1691, n_176, n_59, n_70, n_22860);
  and g55077 (n_22861, n_110, n_190);
  and g55078 (n_22862, n_208, n_172);
  and g55079 (n1245, n590, n1240, n_22861, n_22862);
  and g55080 (n3435, n_240, n_221, n_157, n1141);
  and g55081 (n_22863, n_168, n_199);
  and g55082 (n_22864, n_73, n_209);
  and g55083 (n_22865, n_252, n13671);
  and g55084 (n_22866, n_70, n2466, n2583, n1824);
  and g55085 (n_22867, n4786, n5264, n3108, n772);
  and g55086 (n_22868, n13677, n2345, n2487, n1437);
  and g55087 (n_22869, n2220, n_22863, n_22864, n_22865);
  and g55088 (n13695, n_22866, n_22867, n_22868, n_22869);
  and g55089 (n_22870, n_268, n_66);
  and g55090 (n_22871, n_203, n_79, n_241, n_225);
  and g55091 (n_22872, n_131, n_200, n341, n2219);
  and g55092 (n_22873, n933, n4786, n4794, n439);
  and g55093 (n_22874, n297, n4797, n4799, n_22870);
  and g55094 (n4815, n_22871, n_22872, n_22873, n_22874);
  and g55095 (n13698, n_204, n_83, n_252, n_269);
  and g55096 (n_22875, n_231, n_277, n_219, n_122);
  and g55097 (n_22876, n_134, n_201, n_189, n_205);
  and g55098 (n_22877, n_243, n1731, n3901, n3905);
  and g55099 (n_22878, n732, n3906, n517, n3914);
  and g55100 (n3929, n_22875, n_22876, n_22877, n_22878);
  nor g55101 (n13358, n13352, n13353, n13354, n13355);
  and g55102 (n_22879, n_274, n_70, n_289, n_254);
  and g55103 (n_22880, n_47, n885, n227, n399);
  and g55104 (n_22881, n805, n2202, n2301, n2132);
  and g55105 (n_22882, n4216, n3085, n4218);
  and g55106 (n4232, n_22879, n_22880, n_22881, n_22882);
  and g55107 (n_22883, n_34, n_139, n_282, n_198);
  and g55108 (n_22884, n_223, n_172, n_152, n_263);
  and g55109 (n_22885, n1040, n1726, n471, n288);
  and g55110 (n_22886, n775, n1138, n3300);
  and g55111 (n13210, n_22883, n_22884, n_22885, n_22886);
  and g55112 (n_22887, n_253, n_72, n_45);
  and g55113 (n_22888, n_167, n_160, n_177);
  and g55114 (n_22889, n_148, n_78, n_273);
  and g55115 (n_22890, n826, n621, n3459);
  and g55116 (n13221, n_22887, n_22888, n_22889, n_22890);
  and g55117 (n_22891, n_214, n_285, n_164);
  and g55118 (n_22892, n_114, n_138);
  and g55119 (n_22893, n_36, n_128);
  and g55120 (n_22894, n_55, n2409);
  and g55121 (n2987, n_22891, n_22892, n_22893, n_22894);
  and g55122 (n_22895, n_266, n_136, n_233);
  and g55123 (n_22896, n_268, n_85);
  and g55124 (n_22897, n_99, n_224);
  and g55125 (n_22898, n2698, n3931);
  and g55126 (n3939, n_22895, n_22896, n_22897, n_22898);
  and g55127 (n_22899, n_136, n_164, n_203);
  and g55128 (n_22900, n_154, n_119, n773);
  and g55129 (n_22901, n774, n775);
  and g55130 (n_22902, n776, n778);
  and g55131 (n787, n_22899, n_22900, n_22901, n_22902);
  and g55132 (n_22903, n_238, n_35);
  and g55133 (n751, n_189, n_262, n747, n_22903);
  and g55134 (n_22904, n_266, n_168, n_246, n_52);
  and g55135 (n_22905, n_208, n_205, n_87);
  and g55136 (n_22906, n_80, n_118, n_90);
  and g55137 (n_22907, n2740, n530, n3570);
  and g55138 (n13135, n_22904, n_22905, n_22906, n_22907);
  nor g55139 (n13398, n13392, n13393, n13394, n13397);
  nor g55140 (n13867, n13859, n13860, n13861, n13864);
  nor g55141 (n14058, n14052, n14053, n14054, n14055);
  nor g55142 (n14653, n14647, n14648, n14649, n14652);
  nor g55143 (n15492, n15486, n15487, n15488, n15491);
  nor g55144 (n14821, n14815, n14816, n14817, n14820);
  nor g55145 (n16263, n16257, n16258, n16259, n16262);
  nor g55146 (n23395, n23389, n23390, n23391, n23394);
  nor g55147 (n24758, n24752, n24753, n24754, n24757);
  nor g55148 (n25493, n25487, n25488, n25489, n25492);
  nor g55149 (n26392, n26386, n26387, n26388, n26391);
  and g55150 (n1240, n_165, n_128, n_79, n_177);
  and g55151 (n_22908, n_191, n_290, n_66);
  and g55152 (n_22909, n_278, n_39, n_77);
  and g55153 (n_22910, n_153, n_159, n2021);
  and g55154 (n_22911, n2424, n3040);
  and g55155 (n5264, n_22908, n_22909, n_22910, n_22911);
  and g55156 (n_22912, n_255, n_54, n_223, n_117);
  and g55157 (n_22913, n_88, n_40, n_57, n_47);
  and g55158 (n_22914, n1884, n1827, n2573, n2698);
  and g55159 (n_22915, n3094, n497, n3059);
  and g55160 (n3108, n_22912, n_22913, n_22914, n_22915);
  and g55161 (n_22916, n_75, n_230);
  and g55162 (n_22917, n_177, n_225);
  and g55163 (n_22918, n_272, n_287);
  and g55164 (n13677, n2809, n_22916, n_22917, n_22918);
  and g55165 (n_22919, n_292, n_51, n_156);
  and g55166 (n_22920, n_179, n896, n2325);
  and g55167 (n_22921, n238, n2330, n632);
  and g55168 (n_22922, n2332, n887, n2334);
  and g55169 (n2345, n_22919, n_22920, n_22921, n_22922);
  and g55170 (n2487, n_240, n_165, n_205, n_215);
  and g55171 (n4797, n_102, n_282, n_75, n_132);
  and g55172 (n_22923, n_155, n_185, n_256, n_143);
  and g55173 (n_22924, n_54, n_64, n_209, n_267);
  and g55174 (n_22925, n_272, n_69, n3886, n1824);
  and g55175 (n_22926, n1479, n2633, n2390, n3041);
  and g55176 (n3901, n_22923, n_22924, n_22925, n_22926);
  and g55177 (n_22927, n_279, n_166);
  and g55178 (n3905, n_234, n_38, n_223, n_22927);
  and g55179 (n_22928, n_58, n_132, n_49);
  and g55180 (n_22929, n_111, n_69, n2073);
  and g55181 (n_22930, n1550, n1825, n2154);
  and g55182 (n_22931, n2191, n2192);
  and g55183 (n2202, n_22928, n_22929, n_22930, n_22931);
  and g55184 (n_22932, n_119, n_79);
  and g55185 (n2301, n_272, n827, n2297, n_22932);
  and g55186 (n_22933, n_144, n_246);
  and g55187 (n_22934, n_233, n_99);
  and g55188 (n2132, n_174, n_218, n_22933, n_22934);
  and g55189 (n1138, n_234, n_257, n_125, n_188);
  and g55190 (n2409, n_183, n_279, n_134, n_120);
  nor g55191 (n23412, n23406, n23407, n23408, n23411);
  and g55192 (n_22935, n_274, n_35);
  and g55193 (n_22936, n_170, n1247);
  and g55194 (n1884, n1438, n1879, n_22935, n_22936);
  and g55195 (n_22937, n_155, n_85, n_282);
  and g55196 (n_22938, n_119, n_148, n_46);
  and g55197 (n_22939, n_296, n615);
  and g55198 (n_22940, n723, n3085);
  and g55199 (n3094, n_22937, n_22938, n_22939, n_22940);
  and g55200 (n_22941, n_233, n_63, n_67);
  and g55201 (n_22942, n_203, n_120);
  and g55202 (n_22943, n_132, n_112);
  and g55203 (n_22944, n_55, n_152);
  and g55204 (n2325, n_22941, n_22942, n_22943, n_22944);
  and g55205 (n_22945, n_71, n_251);
  and g55206 (n_22946, n_154, n_142);
  and g55207 (n2330, n_126, n437, n_22945, n_22946);
  and g55208 (n_22947, n_121, n_110, n_172, n_196);
  and g55209 (n_22948, n538, n1761, n3757, n937);
  and g55210 (n_22949, n2740, n3764, n3782);
  and g55211 (n_22950, n3790, n3040, n3792);
  and g55212 (n3805, n_22947, n_22948, n_22949, n_22950);
  and g55213 (n_22951, n_137, n_110);
  and g55214 (n_22952, n_36, n_264);
  and g55215 (n_22953, n_50, n116);
  and g55216 (n_22954, n356, n4786, n120, n12710);
  and g55217 (n_22955, n2573, n1577, n2507, n1549);
  and g55218 (n_22956, n5806, n6054, n1879, n2361);
  and g55219 (n_22957, n12712, n_22951, n_22952, n_22953);
  and g55220 (n12730, n_22954, n_22955, n_22956, n_22957);
  and g55221 (n_22958, n_202, n_192, n_66, n_115);
  and g55222 (n_22959, n570, n1667, n159);
  and g55223 (n_22960, n1479, n12795, n12828);
  and g55224 (n_22961, n6084, n3827, n12830);
  and g55225 (n12842, n_22958, n_22959, n_22960, n_22961);
  nor g55226 (n12872, n12866, n12867, n12868, n12871);
  nor g55227 (n14184, n14178, n14179, n14180, n14181);
  nor g55228 (n23008, n23000, n23001, n23002, n23007);
  nor g55229 (n15479, n15473, n15474, n15475, n15478);
  nor g55230 (n15627, n15621, n15622, n15623, n15626);
  nor g55231 (n16427, n16421, n16422, n16423, n16426);
  nor g55232 (n15176, n15170, n15171, n15172, n15175);
  nor g55233 (n25511, n25505, n25506, n25507, n25510);
  nor g55234 (n26378, n26372, n26373, n26374, n26377);
  and g55235 (n_22962, n_62, n_83, n_149, n_90);
  and g55236 (n_22963, n279, n156, n2406, n1330);
  and g55237 (n_22964, n2090, n13247, n13265, n2772);
  and g55238 (n_22965, n13268, n1557, n3645, n6104);
  and g55239 (n13283, n_22962, n_22963, n_22964, n_22965);
  and g55240 (n_22966, n_65, n_251);
  and g55241 (n_22967, n_234, n_178);
  and g55242 (n_22968, n_291, n_271);
  and g55243 (n_22969, n_59, n_68);
  and g55244 (n12710, n_22966, n_22967, n_22968, n_22969);
  and g55245 (n_22970, n_217, n_130);
  and g55246 (n_22971, n_129, n_223, n_142, n1522);
  and g55247 (n_22972, n590, n1426, n1523, n1305);
  and g55248 (n_22973, n1105, n1527, n439, n723);
  and g55249 (n_22974, n1530, n1331, n1533, n_22970);
  and g55250 (n1549, n_22971, n_22972, n_22973, n_22974);
  and g55251 (n_22975, n_292, n_206, n_84, n_218);
  and g55252 (n_22976, n_49, n_210, n_245, n2758);
  and g55253 (n_22977, n100, n227, n1237);
  and g55254 (n_22978, n5785, n5791, n5793);
  and g55255 (n5806, n_22975, n_22976, n_22977, n_22978);
  and g55256 (n_22979, n_98, n_265, n_189);
  and g55257 (n_22980, n_227, n_67, n_203);
  and g55258 (n_22981, n_171, n_177, n_288);
  and g55259 (n_22982, n_179, n467, n1611);
  and g55260 (n6054, n_22979, n_22980, n_22981, n_22982);
  nor g55261 (n12783, n12777, n12778, n12779, n12780);
  and g55262 (n_22983, n_214, n_122);
  and g55263 (n_22984, n_130, n_86);
  and g55264 (n_22985, n_267, n_196);
  and g55265 (n_22986, n810, n978, n491, n1917);
  and g55266 (n_22987, n247, n3378, n2740, n3405);
  and g55267 (n_22988, n3432, n3225, n3435, n3437);
  and g55268 (n_22989, n3438, n_22983, n_22984, n_22985);
  and g55269 (n3456, n_22986, n_22987, n_22988, n_22989);
  and g55270 (n_22990, n_130, n_274);
  and g55271 (n_22991, n_233, n_249, n_156, n_147);
  and g55272 (n_22992, n_89, n1161, n159, n2484);
  and g55273 (n_22993, n1575, n13768, n2796, n5791);
  and g55274 (n_22994, n1942, n1308, n13789, n_22990);
  and g55275 (n13805, n_22991, n_22992, n_22993, n_22994);
  nor g55276 (n14360, n14354, n14355, n14356, n14359);
  nor g55277 (n14714, n14708, n14709, n14710, n14713);
  nor g55278 (n23027, n23019, n23020, n23021, n23026);
  nor g55279 (n14909, n14903, n14904, n14905, n14908);
  nor g55280 (n15668, n15662, n15663, n15664, n15667);
  and g55281 (n_22995, n_191, n_151);
  and g55282 (n_22996, n_84, n_157);
  and g55283 (n_22997, n418, n1826);
  and g55284 (n_22998, n4797, n12412);
  and g55285 (n13247, n_22995, n_22996, n_22997, n_22998);
  and g55286 (n_22999, n_255, n_100);
  and g55287 (n_23000, n_67, n_205, n_117, n_289);
  and g55288 (n_23001, n_297, n_93, n1366, n1825);
  and g55289 (n_23002, n285, n3544, n1292, n6083);
  and g55290 (n_23003, n6084, n691, n13249, n_22999);
  and g55291 (n13265, n_23000, n_23001, n_23002, n_23003);
  and g55292 (n_23004, n_220, n_98);
  and g55293 (n_23005, n_230, n_125, n_148, n_105);
  and g55294 (n_23006, n507, n2651, n1253, n2738);
  and g55295 (n_23007, n2751, n494, n2544, n2445);
  and g55296 (n_23008, n2752, n2753, n2760, n_23004);
  and g55297 (n2772, n_23005, n_23006, n_23007, n_23008);
  and g55298 (n13268, n_183, n_42, n_162, n590);
  and g55299 (n_23009, n_247, n_169, n_42);
  and g55300 (n_23010, n_185, n_66, n_242);
  and g55301 (n_23011, n_195, n_69, n_211);
  and g55302 (n_23012, n359, n735, n1294);
  and g55303 (n1305, n_23009, n_23010, n_23011, n_23012);
  and g55304 (n_23013, n_53, n_168, n_282);
  and g55305 (n_23014, n_117, n_278);
  and g55306 (n_23015, n_60, n_97);
  and g55307 (n_23016, n5775, n5777);
  and g55308 (n5785, n_23013, n_23014, n_23015, n_23016);
  and g55309 (n_23017, n_88, n_132);
  and g55310 (n5791, n_212, n_47, n5787, n_23017);
  and g55311 (n_23018, n_235, n_233, n_83);
  and g55312 (n_23019, n_142, n_262);
  and g55313 (n_23020, n_68, n2361);
  and g55314 (n_23021, n2426, n3370);
  and g55315 (n3378, n_23018, n_23019, n_23020, n_23021);
  and g55316 (n_23022, n_182, n_34);
  and g55317 (n_23023, n_292, n_201);
  and g55318 (n_23024, n_44, n674);
  and g55319 (n3225, n1531, n_23022, n_23023, n_23024);
  nor g55320 (n12703, n12697, n12698, n12699, n12700);
  and g55321 (n_23025, n_42, n_228, n_257, n888);
  and g55322 (n_23026, n_82, n_241, n_213, n1080);
  and g55323 (n_23027, n4367, n3489, n2716);
  and g55324 (n_23028, n3041, n5271, n13808);
  and g55325 (n13821, n_23025, n_23026, n_23027, n_23028);
  and g55326 (n_23029, n_53, n_251);
  and g55327 (n_23030, n_73, n_181);
  and g55328 (n_23031, n_67, n_127);
  and g55329 (n_23032, n_288, n_47, n1522, n4101);
  and g55330 (n_23033, n2088, n937, n450, n1046);
  and g55331 (n_23034, n14202, n2296, n3681, n529);
  and g55332 (n_23035, n14210, n_23029, n_23030, n_23031);
  and g55333 (n14228, n_23032, n_23033, n_23034, n_23035);
  and g55334 (n_23036, n_168, n_251, n_197);
  and g55335 (n_23037, n_95, n_112, n_141);
  and g55336 (n_23038, n_187, n238, n2090);
  and g55337 (n_23039, n1253, n2739);
  and g55338 (n13768, n_23036, n_23037, n_23038, n_23039);
  and g55339 (n_23040, n_204, n_235, n_265, n_203);
  and g55340 (n_23041, n634, n1237, n515);
  and g55341 (n_23042, n1994, n2778, n2782);
  and g55342 (n_23043, n204, n632, n2784);
  and g55343 (n2796, n_23040, n_23041, n_23042, n_23043);
  nor g55344 (n16992, n16986, n16987, n16988, n16991);
  nor g55345 (n15463, n15457, n15458, n15459, n15462);
  nor g55346 (n23430, n23424, n23425, n23426, n23429);
  nor g55347 (n23751, n23745, n23746, n23747, n23750);
  nor g55348 (n26361, n26355, n26356, n26357, n26360);
  and g55349 (n12412, n_129, n_192, n_119, n2346);
  and g55350 (n_23044, n_285, n_44);
  and g55351 (n_23045, n_128, n_248);
  and g55352 (n_23046, n_95, n_69);
  and g55353 (n_23047, n1426, n1644);
  and g55354 (n6083, n_23044, n_23045, n_23046, n_23047);
  and g55355 (n_23048, n_104, n_186, n_264);
  and g55356 (n_23049, n_108, n_269, n_46);
  and g55357 (n_23050, n1128, n2739);
  and g55358 (n_23051, n2740, n2742);
  and g55359 (n2751, n_23048, n_23049, n_23050, n_23051);
  nor g55360 (n12463, n12457, n12458, n12459, n12460);
  nor g55361 (n12379, n12373, n12374, n12375, n12378);
  and g55362 (n_23052, n_58, n_37);
  and g55363 (n_23053, n_80, n_250);
  and g55364 (n_23054, n_126, n1070);
  and g55365 (n_23055, n1071, n1073);
  and g55366 (n1080, n_23052, n_23053, n_23054, n_23055);
  and g55367 (n_23056, n_63, n_127, n_146, n570);
  and g55368 (n_23057, n1576, n3470, n1046, n615);
  and g55369 (n_23058, n3472, n1601, n437, n593);
  and g55370 (n_23059, n2556, n3474, n754, n3226);
  and g55371 (n3489, n_23056, n_23057, n_23058, n_23059);
  and g55372 (n_23060, n_137, n_277, n_234);
  and g55373 (n_23061, n_267, n_171, n_40);
  and g55374 (n_23062, n_207, n_284, n2507);
  and g55375 (n_23063, n2704, n1636, n2705);
  and g55376 (n2716, n_23060, n_23061, n_23062, n_23063);
  and g55377 (n_23064, n_242, n_175, n_178, n_225);
  and g55378 (n_23065, n515, n2068, n2072, n918);
  and g55379 (n_23066, n1085, n207, n1132);
  and g55380 (n_23067, n812, n1784, n2075);
  and g55381 (n2088, n_23064, n_23065, n_23066, n_23067);
  and g55382 (n_23068, n_253, n_65, n_173, n_297);
  and g55383 (n_23069, n356, n872, n774, n874);
  and g55384 (n_23070, n622, n2022, n14189);
  and g55385 (n_23071, n5777, n1109, n3523);
  and g55386 (n14202, n_23068, n_23069, n_23070, n_23071);
  and g55387 (n2296, n_199, n_221, n_88, n2293);
  and g55388 (n_23072, n_104, n_294);
  and g55389 (n_23073, n_203, n_195);
  and g55390 (n_23074, n_132, n_89);
  and g55391 (n3681, n_287, n_23072, n_23073, n_23074);
  and g55392 (n_23075, n_45, n_138, n_272);
  and g55393 (n_23076, n_284, n1782);
  and g55394 (n_23077, n989, n2390);
  and g55395 (n_23078, n642, n3165);
  and g55396 (n14210, n_23075, n_23076, n_23077, n_23078);
  nor g55397 (n14240, n14234, n14235, n14236, n14237);
  and g55399 (n_23080, n_124, n_127, n_88, n_248);
  and g55400 (n_23081, n_90, n1838, n774, n6514);
  and g55401 (n_23082, n1814, n13826, n434, n3068);
  and g55402 (n_23083, n4298, n1346, n13827, n_22694);
  and g55403 (n13843, n_23080, n_23081, n_23082, n_23083);
  and g55404 (n_23084, n_163, n_256);
  and g55405 (n_23085, n_270, n_128);
  and g55406 (n_23086, n_172, n_262);
  and g55407 (n2778, n_284, n_23084, n_23085, n_23086);
  nor g55408 (n14447, n14438, n14439, n14440, n14444);
  nor g55409 (n14731, n14725, n14726, n14727, n14730);
  nor g55410 (n14746, n14740, n14741, n14742, n14745);
  nor g55411 (n15520, n15514, n15515, n15516, n15519);
  nor g55412 (n15160, n15154, n15155, n15156, n15159);
  nor g55413 (n23768, n23762, n23763, n23764, n23767);
  and g55414 (n_23087, n_266, n_204);
  and g55415 (n_23088, n_168, n_130);
  and g55416 (n_23089, n_258, n_128);
  and g55417 (n_23090, n_215, n_291, n_112, n_46);
  and g55418 (n_23091, n_93, n3559, n1687, n221);
  and g55419 (n_23092, n3565, n1928, n3580, n3583);
  and g55420 (n_23093, n3587, n_23087, n_23088, n_23089);
  and g55421 (n3605, n_23090, n_23091, n_23092, n_23093);
  nor g55422 (n3719, n3711, n3712, n3713, n3716);
  and g55423 (n_23094, n_182, n_231);
  and g55424 (n_23095, n_41, n_163);
  and g55425 (n_23096, n_154, n_252, n_232, n_90);
  and g55426 (n_23097, n_297, n3163, n12396, n6769);
  and g55427 (n_23098, n12404, n12428, n12431, n1158);
  and g55428 (n_23099, n253, n722, n_23094, n_23095);
  and g55429 (n12448, n_23096, n_23097, n_23098, n_23099);
  and g55430 (n_23100, n_217, n_246);
  and g55431 (n_23101, n_283, n_123);
  and g55432 (n_23102, n_291, n792);
  and g55433 (n3470, n2091, n_23100, n_23101, n_23102);
  and g55434 (n_23103, n_53, n_166);
  and g55435 (n_23104, n_294, n_271, n_141, n_147);
  and g55436 (n_23105, n_59, n_243, n1040, n356);
  and g55437 (n_23106, n1667, n1668, n664, n5063);
  and g55438 (n_23107, n1249, n5064, n5066, n_23103);
  and g55439 (n5082, n_23104, n_23105, n_23106, n_23107);
  and g55440 (n_23108, n_247, n_145, n_124);
  and g55441 (n_23109, n_84, n_208, n_269);
  and g55442 (n_23110, n_90, n591);
  and g55443 (n_23111, n735, n2059);
  and g55444 (n2068, n_23108, n_23109, n_23110, n_23111);
  and g55445 (n_23112, n_204, n_106);
  and g55446 (n2072, n_118, n1248, n1252, n_23112);
  and g55447 (n_23113, n_139, n_44);
  and g55448 (n_23114, n_240, n_180);
  and g55449 (n14189, n_85, n_210, n_23113, n_23114);
  and g55450 (n_23115, n_145, n_231, n_163);
  and g55451 (n_23116, n_220, n_223, n_119);
  and g55452 (n_23117, n_288, n591, n1827);
  and g55453 (n_23118, n1667, n1828);
  and g55454 (n1838, n_23115, n_23116, n_23117, n_23118);
  and g55455 (n_23119, n_268, n_161, n_269, n_105);
  and g55456 (n_23120, n_243, n116, n2993, n1139);
  and g55457 (n_23121, n874, n1292, n1794, n4279);
  and g55458 (n_23122, n4828, n2608, n4357);
  and g55459 (n6514, n_23119, n_23120, n_23121, n_23122);
  and g55460 (n_23123, n_71, n_277, n_164, n_133);
  and g55461 (n_23124, n_123, n_177, n_55, n_47);
  and g55462 (n_23125, n193, n515, n1020, n1798);
  and g55463 (n_23126, n494, n1408, n1800);
  and g55464 (n1814, n_23123, n_23124, n_23125, n_23126);
  and g55465 (n_23127, n_109, n_166);
  and g55466 (n_23128, n_221, n_78);
  and g55467 (n13826, n423, n1366, n_23127, n_23128);
  and g55468 (n434, n_183, n_182, n_73, n431);
  and g55469 (n3068, n_229, n_46, n_296, n2633);
  and g55470 (n4298, n_199, n_52, n_35, n_146);
  nor g55471 (n16581, n16575, n16576, n16577, n16580);
  nor g55472 (n16414, n16408, n16409, n16410, n16413);
  nor g55473 (n14893, n14887, n14888, n14889, n14892);
  nor g55474 (n16245, n16239, n16240, n16241, n16244);
  nor g55475 (n23786, n23780, n23781, n23782, n23785);
  nor g55476 (n24331, n24325, n24326, n24327, n24330);
  nor g55477 (n26683, n26677, n26678, n26679, n26682);
  and g55478 (n_23129, n_246, n_140, n_152);
  and g55479 (n_23130, n421, n1574, n3544);
  and g55480 (n_23131, n1479, n2010, n3548);
  and g55481 (n_23132, n1960, n3549);
  and g55482 (n3559, n_23129, n_23130, n_23131, n_23132);
  and g55483 (n_23133, n_85, n_84, n_83, n_82);
  and g55484 (n_23134, n_81, n_80, n_79, n_78);
  and g55485 (n_23135, n_77, n156, n159, n187);
  and g55486 (n_23136, n198, n204, n207);
  and g55487 (n221, n_23133, n_23134, n_23135, n_23136);
  and g55488 (n_23137, n_180, n_181);
  and g55490 (n_23139, n_210, n116);
  and g55491 (n3565, n_297, n_23137, n_23138, n_23139);
  and g55492 (n1928, n_257, n_289, n_90, n_263);
  and g55493 (n_23140, n_155, n_34);
  and g55494 (n3587, n_170, n1330, n1826, n_23140);
  and g55495 (n_23141, n_192, n_76, n_40, n_78);
  and g55496 (n_23142, n_272, n_59, n1366, n1046);
  and g55497 (n_23143, n1915, n3675, n3681, n1323);
  and g55498 (n_23144, n3685, n723, n2427, n3687);
  and g55499 (n3702, n_23141, n_23142, n_23143, n_23144);
  nor g55500 (n4069, n3885, n3968, n4047, n4068);
  and g55501 (n_23145, n_64, n_49);
  and g55502 (n_23146, n_55, n2582);
  and g55503 (n_23147, n12387, n2584);
  and g55504 (n12396, n12390, n_23145, n_23146, n_23147);
  and g55505 (n_23148, n_279, n_240, n_234, n_180);
  and g55506 (n_23149, n_261, n2073, n1824, n2010);
  and g55507 (n_23150, n873, n2738, n6670, n467);
  and g55508 (n_23151, n776, n5201, n5793);
  and g55509 (n6769, n_23148, n_23149, n_23150, n_23151);
  and g55510 (n_23152, n_136, n_199);
  and g55511 (n_23153, n_280, n_188);
  and g55512 (n_23154, n_118, n_38);
  and g55513 (n_23155, n1550, n12397);
  and g55514 (n12404, n_23152, n_23153, n_23154, n_23155);
  and g55515 (n_23156, n_169, n_194);
  and g55516 (n_23157, n_190, n_167, n_153, n_272);
  and g55517 (n_23158, n_131, n885, n1994, n1253);
  and g55518 (n_23159, n774, n811, n2961, n1496);
  and g55519 (n_23160, n12409, n1644, n12412, n_23156);
  and g55520 (n12428, n_23157, n_23158, n_23159, n_23160);
  and g55521 (n12431, n_247, n_228, n_85, n_126);
  and g55522 (n1158, n_253, n_45, n773, n979);
  and g55523 (n_23161, n_163, n_67, n_140, n591);
  and g55524 (n_23162, n1254, n1528, n1029, n3464);
  and g55525 (n_23163, n3489, n3521, n465, n1586);
  and g55526 (n_23164, n530, n3523, n3298, n3524);
  and g55527 (n3539, n_23161, n_23162, n_23163, n_23164);
  and g55528 (n_23165, n_253, n_120);
  and g55529 (n_23166, n_252, n_188);
  and g55530 (n_23167, n_156, n_187);
  and g55531 (n664, n658, n_23165, n_23166, n_23167);
  and g55532 (n_23168, n_84, n_203);
  and g55533 (n_23169, n_173, n896);
  and g55534 (n_23170, n621, n5056);
  and g55535 (n_23171, n2608, n3043);
  and g55536 (n5063, n_23168, n_23169, n_23170, n_23171);
  and g55537 (n_23172, n_258, n_138, n_218);
  and g55538 (n_23173, n_197, n1755, n_210);
  and g55539 (n_23174, n1782, n896);
  and g55540 (n_23175, n1784, n1785);
  and g55541 (n1794, n_23172, n_23173, n_23174, n_23175);
  and g55542 (n_23176, n_228, n_285, n_246);
  and g55543 (n_23177, n_44, n_280);
  and g55544 (n_23178, n_184, n_284);
  and g55545 (n_23179, n_187, n1012);
  and g55546 (n1020, n_23176, n_23177, n_23178, n_23179);
  and g55547 (n1798, n_158, n_216, n_108, n1795);
  nor g55548 (n24022, n24016, n24017, n24018, n24021);
  nor g55549 (n16622, n16616, n16617, n16618, n16621);
  nor g55550 (n17412, n17406, n17407, n17408, n17411);
  nor g55551 (n24348, n24342, n24343, n24344, n24347);
  nor g55552 (n4479, n4471, n4472, n4473, n4478);
  nor g55553 (n25126, n25120, n25121, n25122, n25125);
  and g55554 (n2010, n_44, n_197, n_254, n2007);
  and g55555 (n_23180, n_231, n_139);
  and g55556 (n3548, n_166, n_273, n_268, n_23180);
  and g55557 (n_23181, n_65, n_64, n_63);
  and g55558 (n_23182, n_62, n_61);
  and g55559 (n_23183, n_60, n_59);
  and g55560 (n_23184, n172, n179);
  and g55561 (n187, n_23181, n_23182, n_23183, n_23184);
  and g55562 (n_23185, n_71, n_70);
  and g55563 (n198, n_69, n193, n_68, n_23185);
  and g55564 (n_23186, n_96, n_74, n_289, n_156);
  and g55565 (n_23187, n_187, n804, n3057, n3065);
  and g55566 (n_23188, n2651, n2317, n931, n494);
  and g55567 (n_23189, n3068, n1438, n373, n573);
  and g55568 (n3083, n_23186, n_23187, n_23188, n_23189);
  and g55569 (n_23190, n_253, n_144, n_180, n_198);
  and g55570 (n_23191, n_133, n_189, n3636);
  and g55571 (n_23192, n_47, n241, n3644);
  and g55572 (n_23193, n2581, n3651, n3663);
  and g55573 (n3675, n_23190, n_23191, n_23192, n_23193);
  and g55574 (n_23194, n_145, n_130, n_265);
  and g55575 (n_23195, n_209, n_82);
  and g55576 (n_23196, n_142, n_146);
  and g55577 (n_23197, n1139, n1315);
  and g55578 (n1323, n_23194, n_23195, n_23196, n_23197);
  and g55579 (n_23198, n_109, n_135);
  and g55580 (n3685, n_129, n_224, n_250, n_23198);
  and g55581 (n_23199, n_163, n_72);
  and g55582 (n_23200, n_294, n_150);
  and g55583 (n_23201, n_154, n_210, n_47, n1389);
  and g55584 (n_23202, n590, n2958, n244, n2979);
  and g55585 (n_23203, n2987, n1823, n2990, n2992);
  and g55586 (n_23204, n2113, n2995, n_23199, n_23200);
  and g55587 (n3012, n_23201, n_23202, n_23203, n_23204);
  and g55588 (n12387, n_92, n_48, n288, n2276);
  and g55589 (n6670, n_109, n_130, n_65, n_220);
  and g55590 (n2961, n_283, n_196, n2263, n2752);
  and g55591 (n_23205, n_173, n_81);
  and g55592 (n_23206, n_74, n_68);
  and g55593 (n12409, n533, n1071, n_23205, n_23206);
  and g55594 (n_23207, n_285, n_274);
  and g55595 (n_23208, n_222, n_208);
  and g55596 (n3464, n_105, n3459, n_23207, n_23208);
  and g55597 (n_23209, n_99, n_282);
  and g55598 (n_23210, n_272, n3510);
  and g55599 (n_23211, n2022, n3512);
  and g55600 (n_23212, n172, n3514);
  and g55601 (n3521, n_23209, n_23210, n_23211, n_23212);
  and g55602 (n465, n_114, n_197, n_195, n_196);
  and g55603 (n5056, n_229, n_114, n_212, n_262);
  and g55604 (n_23213, n_83, n_76, n_171, n_60);
  and g55605 (n_23214, n4295, n933, n14407, n3472);
  and g55606 (n_23215, n3405, n268, n1119, n5746);
  and g55607 (n_23216, n1085, n2544, n889, n2363);
  and g55608 (n14422, n_23213, n_23214, n_23215, n_23216);
  nor g55609 (n23226, n23220, n23221, n23222, n23225);
  nor g55610 (n16398, n16392, n16393, n16394, n16397);
  nor g55611 (n18387, n18381, n18382, n18383, n18386);
  nor g55612 (n22863, n22857, n22858, n22859, n22862);
  nor g55613 (n15609, n15603, n15604, n15605, n15608);
  nor g55614 (n14992, n14986, n14987, n14988, n14991);
  nor g55615 (n24818, n24812, n24813, n24814, n24817);
  and g55616 (n_23217, n_169, n_168);
  and g55617 (n_23218, n_167, n100, n108, n116);
  and g55618 (n_23219, n120, n141, n221, n268);
  and g55619 (n_23220, n324, n351, n362, n365);
  and g55620 (n_23221, n370, n373, n376, n_23217);
  and g55621 (n392, n_23218, n_23219, n_23220, n_23221);
  and g55622 (n_23222, n_227, n_254, n_211, n1141);
  and g55623 (n_23223, n533, n3039, n285);
  and g55624 (n_23224, n1781, n3040, n3041);
  and g55625 (n_23225, n3042, n3043, n3045);
  and g55626 (n3057, n_23222, n_23223, n_23224, n_23225);
  and g55627 (n_23226, n_285, n_65);
  and g55628 (n_23227, n_72, n_205);
  and g55629 (n_23228, n_174, n_131);
  and g55630 (n3065, n3059, n_23226, n_23227, n_23228);
  and g55631 (n_23229, n_290, n_240, n_117, n_267);
  and g55632 (n_23230, n_89, n1825, n2169, n2296);
  and g55633 (n_23231, n2301, n2091, n207, n816);
  and g55634 (n_23232, n1533, n1025, n2303);
  and g55635 (n2317, n_23229, n_23230, n_23231, n_23232);
  and g55636 (n_23233, n_103, n_83, n_176);
  and g55637 (n_23234, n_195, n_269, n_148);
  and g55638 (n_23235, n_70, n_106, n918);
  and g55639 (n_23236, n179, n921);
  and g55640 (n931, n_23233, n_23234, n_23235, n_23236);
  and g55641 (n_23237, n_169, n_99, n_160);
  and g55642 (n_23238, n_80, n_252);
  and g55643 (n_23239, n_288, n_212);
  and g55644 (n_23240, n_211, n3226);
  and g55645 (n3644, n_23237, n_23238, n_23239, n_23240);
  and g55646 (n_23241, n_204, n_162, n_114);
  and g55647 (n_23242, n_66, n_88);
  and g55648 (n_23243, n_271, n_105);
  and g55649 (n_23244, n_187, n_243);
  and g55650 (n2581, n_23241, n_23242, n_23243, n_23244);
  and g55651 (n_23245, n_231, n_98);
  and g55652 (n_23246, n_56, n_156);
  and g55653 (n_23247, n_225, n202);
  and g55654 (n3651, n3645, n_23245, n_23246, n_23247);
  and g55655 (n_23248, n_247, n_34, n_161, n_165);
  and g55656 (n_23249, n_154, n_125, n_55);
  and g55657 (n_23250, n_90, n_170, n3252);
  and g55658 (n_23251, n3472, n1408, n1458);
  and g55659 (n3663, n_23248, n_23249, n_23250, n_23251);
  and g55660 (n_23252, n_151, n_110, n_96, n_133);
  and g55661 (n_23253, n_265, n_249, n_141, n_153);
  and g55662 (n_23254, n_131, n_126, n1180, n2219);
  and g55663 (n_23255, n2940, n2943, n990, n1408);
  and g55664 (n2958, n_23252, n_23253, n_23254, n_23255);
  and g55665 (n_23256, n_102, n_204);
  and g55666 (n_23257, n_255, n_238, n_199, n_239);
  and g55667 (n_23258, n2466, n1825, n533, n288);
  and g55668 (n_23259, n2021, n1916, n2961, n2963);
  and g55669 (n_23260, n2230, n832, n1423, n_23256);
  and g55670 (n2979, n_23257, n_23258, n_23259, n_23260);
  and g55671 (n_23261, n_34, n_290);
  and g55672 (n1823, n_227, n454, n508, n_23261);
  and g55673 (n2990, n_220, n_118, n634, n1009);
  and g55674 (n_23262, n_162, n3490, n_178, n_107);
  and g55675 (n_23263, n_243, n1269, n291, n2021);
  and g55676 (n_23264, n614, n3497, n2007);
  and g55677 (n_23265, n2220, n941, n1255);
  and g55678 (n3510, n_23262, n_23263, n_23264, n_23265);
  and g55680 (n_23267, n_135, n_235);
  and g55681 (n_23268, n4294, n_113, n_179, n1389);
  and g55682 (n_23269, n1367, n2583, n14381, n6097);
  and g55683 (n_23270, n2772, n14386, n2022, n4130);
  and g55684 (n_23271, n1996, n13114, n_23084, n_23267);
  and g55685 (n14403, n_23268, n_23269, n_23270, n_23271);
  and g55686 (n_23272, n_42, n_52);
  and g55687 (n14407, n_244, n1140, n2210, n_23272);
  and g55688 (n_23273, n_109, n_108, n_107, n227);
  and g55689 (n_23274, n230, n235, n238);
  and g55690 (n_23275, n241, n244, n247);
  and g55691 (n_23276, n250, n253, n256);
  and g55692 (n268, n_23273, n_23274, n_23275, n_23276);
  and g55693 (n_23277, n_43, n_176, n_184);
  and g55694 (n_23278, n_291, n_272, n_196);
  and g55695 (n_23279, n_174, n_47, n1103);
  and g55696 (n_23280, n1107, n1109);
  and g55697 (n1119, n_23277, n_23278, n_23279, n_23280);
  and g55698 (n_23281, n_253, n_191, n_294, n_221);
  and g55699 (n_23282, n_278, n_200, n1575);
  and g55700 (n_23283, n977, n3160, n1424);
  and g55701 (n_23284, n3583, n3687, n5734);
  and g55702 (n5746, n_23281, n_23282, n_23283, n_23284);
  nor g55703 (n14461, n14455, n14456, n14457, n14458);
  nor g55704 (n22571, n22563, n22564, n22565, n22570);
  nor g55705 (n16455, n16449, n16450, n16451, n16454);
  nor g55706 (n14875, n14869, n14870, n14871, n14874);
  nor g55707 (n16229, n16223, n16224, n16225, n16228);
  nor g55708 (n15221, n15215, n15216, n15217, n15220);
  nor g55709 (n24366, n24360, n24361, n24362, n24365);
  nor g55710 (n24835, n24829, n24830, n24831, n24834);
  and g55711 (n_23285, n_49, n_48);
  and g55712 (n141, n128, n133, n137, n_23285);
  and g55713 (n_23286, n_137, n_136);
  and g55714 (n_23287, n_135, n_134, n_133, n_132);
  and g55715 (n_23288, n_131, n279, n282, n285);
  and g55716 (n_23289, n288, n291, n294, n297);
  and g55717 (n_23290, n300, n303, n308, n_23286);
  and g55718 (n324, n_23287, n_23288, n_23289, n_23290);
  and g55719 (n_23291, n_151, n_150, n_149);
  and g55720 (n_23292, n_148, n_147);
  and g55721 (n_23293, n_146, n333);
  and g55722 (n_23294, n336, n343);
  and g55723 (n351, n_23291, n_23292, n_23293, n_23294);
  and g55724 (n362, n_157, n_156, n356, n359);
  and g55725 (n_23295, n_204, n_246);
  and g55726 (n_23296, n_99, n_133);
  and g55727 (n_23297, n_154, n_120);
  and g55728 (n_23298, n_132, n2760);
  and g55729 (n3039, n_23295, n_23296, n_23297, n_23298);
  and g55730 (n921, n_247, n_44, n_68, n_259);
  and g55731 (n_23299, n_266, n_145, n_256);
  and g55732 (n_23300, n_129, n_248, n_188);
  and g55733 (n_23301, n_225, n_287);
  and g55734 (n_23302, n2090, n2931);
  and g55735 (n2940, n_23299, n_23300, n_23301, n_23302);
  and g55736 (n2943, n_35, n_230, n_80, n1556);
  and g55737 (n_23303, n_143, n_135, n_199);
  and g55738 (n_23304, n_235, n_242, n_98);
  and g55739 (n_23305, n_37, n_125, n_241);
  and g55740 (n_23306, n359, n604);
  and g55741 (n614, n_23303, n_23304, n_23305, n_23306);
  and g55742 (n_23307, n_94, n_76);
  and g55743 (n_23308, n_267, n_115);
  and g55744 (n_23309, n_153, n1531);
  and g55745 (n_23310, n401, n2113);
  and g55746 (n3497, n_23307, n_23308, n_23309, n_23310);
  and g55747 (n_23311, n_164, n_66, n_127);
  and g55748 (n_23312, n_205, n_216, n_232);
  and g55749 (n_23313, n_225, n_48, n2698);
  and g55750 (n_23314, n1271, n1602);
  and g55751 (n14381, n_23311, n_23312, n_23313, n_23314);
  and g55752 (n_23315, n_194, n_87, n_132, n_107);
  and g55753 (n_23316, n_263, n979, n454, n1029);
  and g55754 (n_23317, n1601, n5193, n6084);
  and g55755 (n_23318, n1438, n2593, n5150);
  and g55756 (n6097, n_23315, n_23316, n_23317, n_23318);
  and g55757 (n_23319, n_162, n_63);
  and g55758 (n_23320, n_173, n_101);
  and g55759 (n14386, n_111, n5064, n_23319, n_23320);
  and g55760 (n4130, n_229, n_97, n1139, n1781);
  nor g55761 (n17399, n17393, n17394, n17395, n17398);
  nor g55762 (n17869, n17863, n17864, n17865, n17868);
  nor g55763 (n22584, n22576, n22577, n22578, n22583);
  nor g55764 (n18930, n18924, n18925, n18926, n18929);
  nor g55765 (n16974, n16968, n16969, n16970, n16973);
  nor g55766 (n14844, n14838, n14839, n14840, n14841);
  nor g55767 (n15445, n15439, n15440, n15441, n15444);
  nor g55768 (n22895, n22889, n22890, n22891, n22894);
  and g55769 (n2931, n_253, n_201, n_76, n_149);
  and g55770 (n5193, n_149, n_284, n2423, n5190);
  nor g55771 (n17910, n17904, n17905, n17906, n17909);
  nor g55772 (n22712, n22706, n22707, n22708, n22711);
  nor g55773 (n22651, n22643, n22644, n22645, n22650);
  nor g55774 (n22597, n22589, n22590, n22591, n22596);
  nor g55775 (n15593, n15587, n15588, n15589, n15592);
  nor g55776 (n23087, n23081, n23082, n23083, n23086);
  nor g55777 (n15142, n15136, n15137, n15138, n15141);
  nor g55778 (n25571, n25565, n25566, n25567, n25570);
  nor g55779 (n3032, n3019, n3021, n3024, n3029);
  nor g55780 (n4701, n4695, n4696, n4697, n4700);
  and g55781 (n_23321, n_41, n_94);
  and g55782 (n_23322, n_203, n_101, n_245, n_89);
  and g55783 (n_23323, n356, n159, n2739, n622);
  and g55784 (n_23324, n14476, n4247, n14498, n207);
  and g55785 (n_23325, n3985, n674, n1646, n_23321);
  and g55786 (n14514, n_23322, n_23323, n_23324, n_23325);
  nor g55787 (n16563, n16557, n16558, n16559, n16562);
  nor g55788 (n17383, n17377, n17378, n17379, n17382);
  nor g55789 (n20136, n20130, n20131, n20132, n20135);
  nor g55790 (n15691, n15685, n15686, n15687, n15690);
  nor g55791 (n16290, n16284, n16285, n16286, n16289);
  nor g55792 (n14612, n14604, n14605, n14606, n14609);
  nor g55793 (n24853, n24847, n24848, n24849, n24852);
  nor g55794 (n25588, n25582, n25583, n25584, n25587);
  nor g55795 (n26293, n26287, n26288, n26289, n26292);
  nor g55796 (n4086, n4078, n4079, n4080, n4085);
  nor g55797 (n3354, n3348, n3349, n3350, n3351);
  nor g55798 (n4918, n4912, n4913, n4914, n4917);
  and g55799 (n_23326, n_45, n_165, n_205);
  and g55800 (n_23327, n_172, n_254, n_59);
  and g55801 (n_23328, n_243, n665);
  and g55802 (n_23329, n1204, n2154);
  and g55803 (n14476, n_23326, n_23327, n_23328, n_23329);
  and g55804 (n_23330, n_129, n_35, n_189, n_249);
  and g55805 (n_23331, n_91, n_39, n_156, n_48);
  and g55806 (n_23332, n156, n2740, n2017);
  and g55807 (n_23333, n778, n3827, n4234);
  and g55808 (n4247, n_23330, n_23331, n_23332, n_23333);
  and g55809 (n_23334, n_42, n_34);
  and g55810 (n_23335, n_111, n_296, n_174, n1269);
  and g55811 (n_23336, n1380, n827, n1330, n1292);
  and g55812 (n_23337, n14479, n1940, n198, n14482);
  and g55813 (n_23338, n2653, n1425, n3549, n_23334);
  and g55814 (n14498, n_23335, n_23336, n_23337, n_23338);
  nor g55815 (n17440, n17434, n17435, n17436, n17439);
  nor g55816 (n16958, n16952, n16953, n16954, n16957);
  nor g55817 (n15429, n15423, n15424, n15425, n15428);
  nor g55818 (n20791, n20785, n20786, n20787, n20790);
  nor g55819 (n19493, n19487, n19488, n19489, n19492);
  nor g55820 (n18917, n18911, n18912, n18913, n18916);
  nor g55821 (n23490, n23484, n23485, n23486, n23489);
  nor g55822 (n3338, n3332, n3333, n3334, n3335);
  and g55823 (n_23339, n_136, n_64);
  and g55824 (n_23340, n_209, n_173);
  and g55825 (n_23341, n_195, n_297);
  and g55826 (n_23342, n341, n1237, n1994, n3108);
  and g55827 (n_23343, n512, n3127, n1488, n1126);
  and g55828 (n_23344, n2091, n690, n439, n897);
  and g55829 (n_23345, n3128, n_23339, n_23340, n_23341);
  and g55830 (n3146, n_23342, n_23343, n_23344, n_23345);
  nor g55831 (n4571, n4565, n4566, n4567, n4570);
  and g55832 (n_23346, n_102, n_53, n_155, n_273);
  and g55833 (n_23347, n1574, n621, n120, n3155);
  and g55834 (n_23348, n3180, n3205, n3219);
  and g55835 (n_23349, n3225, n2332, n3226);
  and g55836 (n3239, n_23346, n_23347, n_23348, n_23349);
  and g55837 (n2017, n_193, n1105, n2013, n2014);
  and g55838 (n14479, n_137, n_103, n_242, n_291);
  and g55839 (n_23350, n_151, n_110, n_134);
  and g55840 (n_23351, n_142, n_215, n_250);
  and g55841 (n_23352, n1426, n874);
  and g55842 (n_23353, n1557, n1931);
  and g55843 (n1940, n_23350, n_23351, n_23352, n_23353);
  and g55844 (n14482, n_190, n_230, n510, n_269);
  nor g55845 (n16380, n16374, n16375, n16376, n16379);
  nor g55846 (n18369, n18363, n18364, n18365, n18368);
  nor g55847 (n15543, n15537, n15538, n15539, n15542);
  nor g55848 (n20810, n20804, n20805, n20806, n20809);
  nor g55849 (n22954, n22948, n22949, n22950, n22953);
  nor g55850 (n15010, n15004, n15005, n15006, n15007);
  nor g55851 (n23119, n23113, n23114, n23115, n23118);
  nor g55852 (n25606, n25600, n25601, n25602, n25605);
  nor g55853 (n26279, n26273, n26274, n26275, n26278);
  and g55854 (n_23354, n_53, n_239, n_91, n570);
  and g55855 (n_23355, n804, n3252, n872, n3282);
  and g55856 (n_23356, n3312, n2237, n524);
  and g55857 (n_23357, n1931, n1071, n3314);
  and g55858 (n3327, n_23354, n_23355, n_23356, n_23357);
  and g55859 (n_23358, n_43, n_66, n_97, n1248);
  and g55860 (n_23359, n1366, n1781, n2678);
  and g55861 (n_23360, n1917, n3113, n1132);
  and g55862 (n_23361, n3114, n1333, n3115);
  and g55863 (n3127, n_23358, n_23359, n_23360, n_23361);
  and g55864 (n_23362, n_139, n_73);
  and g55865 (n_23363, n_84, n_261);
  and g55866 (n1126, n_172, n1121, n_23362, n_23363);
  nor g55867 (n4186, n4180, n4181, n4182, n4183);
  and g55868 (n_23364, n_102, n_235, n_234, n_98);
  and g55869 (n_23365, n_127, n_77, n193, n415);
  and g55870 (n_23366, n488, n491, n503, n556);
  and g55871 (n_23367, n561, n566, n573);
  and g55872 (n587, n_23364, n_23365, n_23366, n_23367);
  nor g55873 (n4684, n4678, n4679, n4680, n4683);
  and g55874 (n_23368, n_158, n_103);
  and g55875 (n_23369, n_214, n_198);
  and g55876 (n_23370, n_223, n2467);
  and g55877 (n_23371, n128, n3148);
  and g55878 (n3155, n_23368, n_23369, n_23370, n_23371);
  and g55879 (n_23372, n_177, n_252, n_106, n_47);
  and g55880 (n_23373, n341, n810, n3159, n804);
  and g55881 (n_23374, n1139, n1063, n2633, n665);
  and g55882 (n_23375, n3160, n3162, n2349, n3165);
  and g55883 (n3180, n_23372, n_23373, n_23374, n_23375);
  and g55884 (n_23376, n_35, n_85, n_149);
  and g55885 (n_23377, n_215, n1252, n731);
  and g55886 (n_23378, n1825, n3191, n1555);
  and g55887 (n_23379, n1423, n3192, n3194);
  and g55888 (n3205, n_23376, n_23377, n_23378, n_23379);
  and g55889 (n_23380, n_71, n_238, n_144, n_268);
  and g55890 (n_23381, n_61, n_270, n_36, n_101);
  and g55891 (n_23382, n_291, n_263, n_179);
  and g55892 (n_23383, n_93, n_243, n3206);
  and g55893 (n3219, n_23380, n_23381, n_23382, n_23383);
  and g55894 (n1931, n_164, n_195, n244, n_188);
  nor g55895 (n16547, n16541, n16542, n16543, n16546);
  nor g55896 (n20120, n20114, n20115, n20116, n20119);
  nor g55897 (n16211, n16205, n16206, n16207, n16210);
  nor g55898 (n20845, n20839, n20840, n20841, n20844);
  nor g55899 (n18901, n18895, n18896, n18897, n18900);
  and g55900 (n_23384, n_71, n_247, n_227, n_157);
  and g55901 (n_23385, n_250, n_156, n291, n773);
  and g55902 (n_23386, n3259, n3261, n1012, n2931);
  and g55903 (n_23387, n3264, n3266, n3268);
  and g55904 (n3282, n_23384, n_23385, n_23386, n_23387);
  and g55905 (n_23388, n_92, n_194, n_235, n507);
  and g55906 (n_23389, n731, n423, n128);
  and g55907 (n_23390, n1479, n3290, n1523);
  and g55908 (n_23391, n3296, n3298, n3300);
  and g55909 (n3312, n_23388, n_23389, n_23390, n_23391);
  and g55910 (n_23392, n_234, n_193);
  and g55911 (n_23393, n_177, n_70);
  and g55912 (n_23394, n_263, n1942);
  and g55913 (n_23395, n133, n2230);
  and g55914 (n2237, n_23392, n_23393, n_23394, n_23395);
  and g55915 (n_23396, n_133, n_216);
  and g55916 (n524, n_215, n517, n520, n_23396);
  and g55917 (n2678, n_130, n_96, n_153, n_224);
  and g55918 (n_23397, n_294, n_58);
  and g55919 (n_23398, n_113, n_273);
  and g55920 (n3113, n_196, n2191, n_23397, n_23398);
  and g55921 (n_23399, n_259, n_150);
  and g55922 (n_23400, n_215, n590, n202, n591);
  and g55923 (n_23401, n600, n614, n615, n333);
  and g55924 (n_23402, n616, n653, n688, n690);
  and g55925 (n_23403, n691, n693, n694, n_23399);
  and g55926 (n710, n_23400, n_23401, n_23402, n_23403);
  and g55927 (n_23404, n_121, n_151, n_176);
  and g55928 (n_23405, n_175, n_125, n_57);
  and g55929 (n_23406, n_174, n_38, n399);
  and g55930 (n_23407, n401, n405);
  and g55931 (n415, n_23404, n_23405, n_23406, n_23407);
  and g55932 (n_23408, n_145, n_203, n_105, n418);
  and g55933 (n_23409, n421, n423, n159, n448);
  and g55934 (n_23410, n450, n459, n465);
  and g55935 (n_23411, n467, n473, n475);
  and g55936 (n488, n_23408, n_23409, n_23410, n_23411);
  and g55937 (n_23412, n_92, n_209);
  and g55938 (n_23413, n_119, n_70);
  and g55939 (n_23414, n_97, n494);
  and g55940 (n503, n497, n_23412, n_23413, n_23414);
  and g55941 (n_23415, n_99, n_224, n_223, n_81);
  and g55942 (n_23416, n_59, n108, n507, n508);
  and g55943 (n_23417, n510, n512, n524, n526);
  and g55944 (n_23418, n529, n530, n535, n541);
  and g55945 (n556, n_23415, n_23416, n_23417, n_23418);
  nor g55946 (n4967, n4961, n4962, n4963, n4966);
  and g55947 (n_23419, n_124, n_197);
  and g55948 (n3159, n_172, n876, n2808, n_23419);
  and g55949 (n_23420, n_137, n_122, n_86);
  and g55950 (n_23421, n_94, n_134, n_64);
  and g55951 (n_23422, n_161, n_74, n_38);
  and g55952 (n_23423, n193, n401, n510);
  and g55953 (n3191, n_23420, n_23421, n_23422, n_23423);
  and g55954 (n_23424, n_110, n_193);
  and g55955 (n_23425, n_283, n1550);
  and g55956 (n1555, n202, n282, n_23424, n_23425);
  nor g55957 (n5503, n5497, n5498, n5499, n5502);
  nor g55958 (n17851, n17845, n17846, n17847, n17850);
  nor g55959 (n16645, n16639, n16640, n16641, n16644);
  nor g55960 (n15262, n15256, n15257, n15258, n15259);
  nor g55961 (n15242, n15236, n15237, n15238, n15241);
  nor g55962 (n19477, n19471, n19472, n19473, n19476);
  and g55963 (n_23426, n_42, n_140, n_68, n1180);
  and g55964 (n_23427, n356, n720, n2443, n2633);
  and g55965 (n_23428, n14525, n14534, n14544, n3113);
  and g55966 (n_23429, n2317, n3512, n2026, n2995);
  and g55967 (n14559, n_23426, n_23427, n_23428, n_23429);
  and g55968 (n_23430, n_73, n_94);
  and g55969 (n_23431, n_225, n_113, n_118, n_187);
  and g55970 (n_23432, n1857, n471, n2170, n187);
  and g55971 (n_23433, n2738, n3565, n1958, n2093);
  and g55972 (n_23434, n15012, n256, n5173, n_23430);
  and g55973 (n15028, n_23431, n_23432, n_23433, n_23434);
  nor g55974 (n23178, n23172, n23173, n23174, n23177);
  nor g55975 (n23846, n23840, n23841, n23842, n23845);
  nor g55976 (n26262, n26256, n26257, n26258, n26261);
  nor g55977 (n23522, n23516, n23517, n23518, n23521);
  and g55978 (n_23435, n_71, n_204);
  and g55979 (n_23436, n_274, n_201, n_85, n_208);
  and g55980 (n_23437, n_249, n_125, n_78, n_273);
  and g55981 (n_23438, n770, n772, n787, n802);
  and g55982 (n_23439, n844, n846, n851, n_23435);
  and g55983 (n867, n_23436, n_23437, n_23438, n_23439);
  and g55984 (n_23440, n_268, n_67);
  and g55985 (n_23441, n_248, n_252);
  and g55986 (n_23442, n_113, n_50);
  and g55987 (n_23443, n_170, n2705);
  and g55988 (n3259, n_23440, n_23441, n_23442, n_23443);
  and g55989 (n3264, n_255, n_107, n_152, n539);
  and g55990 (n_23444, n_137, n_217, n_249);
  and g55991 (n_23445, n_218, n_125);
  and g55992 (n_23446, n_140, n_271);
  and g55993 (n_23447, n_225, n_296);
  and g55994 (n3290, n_23444, n_23445, n_23446, n_23447);
  and g55995 (n_23448, n_220, n_280);
  and g55996 (n_23449, n_85, n_282);
  and g55997 (n_23450, n_264, n_112);
  and g55998 (n3296, n720, n_23448, n_23449, n_23450);
  and g55999 (n_23451, n_73, n_186);
  and g56000 (n_23452, n_150, n1524);
  and g56001 (n_23453, n_173, n_149);
  and g56002 (n_23454, n_289, n_152, n_174, n1040);
  and g56003 (n_23455, n454, n235, n773, n3408);
  and g56004 (n_23456, n4148, n3521, n2371, n4151);
  and g56005 (n_23457, n4153, n_23451, n_23452, n_23453);
  and g56006 (n4171, n_23454, n_23455, n_23456, n_23457);
  nor g56007 (n4208, n4200, n4201, n4202, n4205);
  and g56008 (n_23458, n_41, n_234);
  and g56009 (n_23459, n_57, n_47);
  and g56010 (n600, n593, n595, n_23458, n_23459);
  and g56011 (n_23460, n_229, n_54, n_180, n_218);
  and g56012 (n_23461, n_195, n_178, n_146, n450);
  and g56013 (n_23462, n654, n664, n665);
  and g56014 (n_23463, n671, n674, n675);
  and g56015 (n688, n_23460, n_23461, n_23462, n_23463);
  and g56016 (n_23464, n_190, n_189, n_160);
  and g56017 (n_23465, n_112, n_188, n_68);
  and g56018 (n_23466, n_187, n434);
  and g56019 (n_23467, n437, n439);
  and g56020 (n448, n_23464, n_23465, n_23466, n_23467);
  and g56021 (n_23468, n_194, n_86);
  and g56022 (n_23469, n_116, n_120);
  and g56023 (n459, n_118, n454, n_23468, n_23469);
  nor g56024 (n26695, n26689, n26690, n26691, n26694);
  nor g56025 (n5646, n5640, n5641, n5642, n5645);
  nor g56026 (n16364, n16358, n16359, n16360, n16363);
  nor g56027 (n24034, n24028, n24029, n24030, n24033);
  nor g56028 (n18353, n18347, n18348, n18349, n18352);
  nor g56029 (n17019, n17013, n17014, n17015, n17018);
  nor g56030 (n15560, n15554, n15555, n15556, n15559);
  nor g56031 (n15575, n15569, n15570, n15571, n15574);
  and g56032 (n_23470, n_137, n_285);
  and g56033 (n_23471, n_45, n_239);
  and g56034 (n_23472, n_232, n1576);
  and g56035 (n_23473, n2348, n14518);
  and g56036 (n14525, n_23470, n_23471, n_23472, n_23473);
  and g56037 (n_23474, n_94, n_129, n_195);
  and g56038 (n_23475, n_184, n_271, n227);
  and g56039 (n_23476, n450, n2192, n4132);
  and g56040 (n_23477, n497, n1315);
  and g56041 (n14544, n_23474, n_23475, n_23476, n_23477);
  and g56042 (n_23478, n_72, n_207, n_232, n_271);
  and g56043 (n_23479, n_147, n_272, n1824, n1825);
  and g56044 (n_23480, n826, n1576, n520);
  and g56045 (n_23481, n1826, n1838, n1844);
  and g56046 (n1857, n_23478, n_23479, n_23480, n_23481);
  and g56047 (n_23482, n_109, n_169, n_285, n_294);
  and g56048 (n_23483, n_268, n_114, n_96, n_40);
  and g56049 (n_23484, n538, n977, n1928, n1940);
  and g56050 (n_23485, n1942, n989, n1944);
  and g56051 (n1958, n_23482, n_23483, n_23484, n_23485);
  and g56052 (n_23486, n_206, n_54);
  and g56053 (n_23487, n_223, n_76, n_174, n_187);
  and g56054 (n_23488, n359, n14565, n120, n1100);
  and g56055 (n_23489, n14572, n13265, n1692, n5036);
  and g56056 (n_23490, n693, n1896, n2293, n_23486);
  and g56057 (n14588, n_23487, n_23488, n_23489, n_23490);
  and g56058 (n_23491, n_182, n_62, n_265, n_264);
  and g56059 (n_23492, n_74, n227, n719, n720);
  and g56060 (n_23493, n730, n731, n745);
  and g56061 (n_23494, n751, n754, n757);
  and g56062 (n770, n_23491, n_23492, n_23493, n_23494);
  and g56063 (n_23495, n_191, n788, n_110);
  and g56064 (n_23496, n_175, n_57, n622);
  and g56065 (n_23497, n789, n790);
  and g56066 (n_23498, n792, n793);
  and g56067 (n802, n_23495, n_23496, n_23497, n_23498);
  and g56068 (n_23499, n_219, n_112, n_271, n_105);
  and g56069 (n_23500, n_225, n_211, n804);
  and g56070 (n_23501, n805, n808, n824);
  and g56071 (n_23502, n830, n467, n832);
  and g56072 (n844, n_23499, n_23500, n_23501, n_23502);
  and g56073 (n_23503, n_290, n_116);
  and g56074 (n_23504, n_120, n_149);
  and g56075 (n_23505, n4101, n507, n1183, n2500);
  and g56076 (n_23506, n3901, n3405, n2217, n877);
  and g56077 (n_23507, n2943, n4104, n2192, n792);
  and g56078 (n_23508, n250, n1760, n_23503, n_23504);
  and g56079 (n4121, n_23505, n_23506, n_23507, n_23508);
  and g56080 (n_23509, n_290, n_72);
  and g56081 (n_23510, n_258, n_218, n_239, n_291);
  and g56082 (n_23511, n_140, n_48, n1141, n1251);
  and g56083 (n_23512, n491, n4127, n4130, n1692);
  and g56084 (n_23513, n812, n1045, n4132, n_23509);
  and g56085 (n4148, n_23510, n_23511, n_23512, n_23513);
  and g56086 (n_23514, n_53, n_209);
  and g56087 (n_23515, n_165, n_171);
  and g56088 (n_23516, n_153, n_262, n869, n423);
  and g56089 (n_23517, n872, n873, n874, n882);
  and g56090 (n_23518, n916, n931, n936, n940);
  and g56091 (n_23519, n475, n941, n_23514, n_23515);
  and g56092 (n958, n_23516, n_23517, n_23518, n_23519);
  and g56093 (n_23520, n_255, n_214);
  and g56094 (n671, n_181, n_113, n_254, n_23520);
  nor g56095 (n4664, n4658, n4659, n4660, n4663);
  nor g56096 (n4637, n4629, n4630, n4631, n4634);
  nor g56097 (n25138, n25132, n25133, n25134, n25137);
  nor g56098 (n5394, n5388, n5389, n5390, n5393);
  nor g56099 (n23238, n23232, n23233, n23234, n23237);
  nor g56100 (n23249, n23243, n23244, n23245, n23246);
  nor g56101 (n16478, n16472, n16473, n16474, n16477);
  nor g56102 (n17365, n17359, n17360, n17361, n17364);
  nor g56103 (n22124, n22118, n22119, n22120, n22123);
  nor g56104 (n19535, n19529, n19530, n19531, n19534);
  nor g56105 (n16195, n16189, n16190, n16191, n16194);
  nor g56106 (n20863, n20857, n20858, n20859, n20862);
  nor g56107 (n18885, n18879, n18880, n18881, n18884);
  and g56108 (n_23521, n_240, n_178);
  and g56109 (n_23522, n_79, n_153);
  and g56110 (n1844, n962, n1839, n_23521, n_23522);
  and g56111 (n_23523, n_73, n_218);
  and g56112 (n14565, n_118, n_296, n14561, n_23523);
  and g56113 (n_23524, n_136, n_163, n_143, n_162);
  and g56114 (n_23525, n_259, n_124, n_288, n_39);
  and g56115 (n_23526, n570, n159, n1063, n1069);
  and g56116 (n_23527, n1080, n1084, n256, n1085);
  and g56117 (n1100, n_23524, n_23525, n_23526, n_23527);
  and g56118 (n_23528, n_135, n_208);
  and g56119 (n_23529, n_116, n_78);
  and g56120 (n_23530, n810, n1602);
  and g56121 (n_23531, n1695, n2012);
  and g56122 (n14572, n_23528, n_23529, n_23530, n_23531);
  nor g56123 (n23878, n23872, n23873, n23874, n23877);
  nor g56124 (n24426, n24420, n24421, n24422, n24425);
  and g56125 (n719, n_261, n_160, n137, n_196);
  and g56126 (n_23532, n_158, n_34, n_234);
  and g56127 (n_23533, n_193, n_101, n_128);
  and g56128 (n_23534, n_118, n_97, n732);
  and g56129 (n_23535, n734, n735);
  and g56130 (n745, n_23532, n_23533, n_23534, n_23535);
  and g56131 (n757, n_130, n_94, n193, n_205);
  and g56132 (n_23536, n_229, n_162, n_98);
  and g56133 (n_23537, n_88, n810);
  and g56134 (n_23538, n811, n812);
  and g56135 (n_23539, n814, n816);
  and g56136 (n824, n_23536, n_23537, n_23538, n_23539);
  and g56137 (n830, n_270, n_49, n826, n827);
  and g56138 (n_23540, n_266, n_285, n_49, n_269);
  and g56139 (n_23541, n_38, n_287, n885, n896);
  and g56140 (n_23542, n621, n1915, n2487);
  and g56141 (n_23543, n300, n365, n1204);
  and g56142 (n2500, n_23540, n_23541, n_23542, n_23543);
  and g56143 (n_23544, n_261, n_88);
  and g56144 (n_23545, n_232, n_225);
  and g56145 (n_23546, n_113, n887);
  and g56146 (n_23547, n2209, n2210);
  and g56147 (n2217, n_23544, n_23545, n_23546, n_23547);
  and g56148 (n4104, n_160, n_57, n_152, n_284);
  and g56149 (n_23548, n_168, n_166);
  and g56150 (n_23549, n_280, n_62);
  and g56151 (n_23550, n_283, n_176);
  and g56152 (n4127, n1073, n_23548, n_23549, n_23550);
  and g56153 (n_23551, n_276, n_151);
  and g56154 (n_23552, n_75, n_241);
  and g56155 (n882, n876, n877, n_23551, n_23552);
  and g56156 (n_23553, n_183, n_279);
  and g56157 (n_23554, n_138, n_270);
  and g56158 (n_23555, n_278, n_244, n572, n_89);
  and g56159 (n_23556, n885, n507, n895, n399);
  and g56160 (n_23557, n896, n128, n539, n851);
  and g56161 (n_23558, n897, n899, n_23553, n_23554);
  and g56162 (n916, n_23555, n_23556, n_23557, n_23558);
  and g56163 (n936, n_85, n454, n235, n933);
  and g56164 (n940, n_246, n_157, n_113, n937);
  nor g56165 (n4898, n4892, n4893, n4894, n4897);
  nor g56166 (n5486, n5480, n5481, n5482, n5485);
  and g56167 (n_23559, n_233, n_257);
  and g56168 (n_23560, n_283, n_88);
  and g56169 (n_23561, n_112, n_179);
  and g56170 (n_23562, n15867, n731, n1129, n294);
  and g56171 (n_23563, n967, n5209, n6625, n3261);
  and g56172 (n_23564, n732, n12387, n3041, n13774);
  and g56173 (n_23565, n23251, n_23559, n_23560, n_23561);
  and g56174 (n23269, n_23562, n_23563, n_23564, n_23565);
  nor g56175 (n22733, n22727, n22728, n22729, n22732);
  and g56176 (n_23566, n_162, n_84);
  and g56177 (n_23567, n_138, n_70);
  and g56178 (n_23568, n_174, n341, n1128, n810);
  and g56179 (n_23569, n1180, n1269, n1161, n15867);
  and g56180 (n_23570, n22748, n22762, n15956, n1044);
  and g56181 (n_23571, n735, n2075, n_23566, n_23567);
  and g56182 (n22779, n_23568, n_23569, n_23570, n_23571);
  nor g56183 (n17835, n17829, n17830, n17831, n17834);
  nor g56184 (n16940, n16934, n16935, n16936, n16939);
  nor g56185 (n15392, n15386, n15387, n15388, n15389);
  and g56186 (n_23572, n_276, n_61);
  and g56187 (n1069, n_171, n_170, n1065, n_23572);
  and g56188 (n_23573, n_194, n_180);
  and g56189 (n1084, n_221, n_70, n_123, n_23573);
  nor g56190 (n23581, n23575, n23576, n23577, n23580);
  and g56191 (n_23574, n_52, n_189, n_210, n_241);
  and g56192 (n_23575, n885, n967, n976, n622);
  and g56193 (n_23576, n977, n1008, n1039);
  and g56194 (n_23577, n1044, n1045, n1047);
  and g56195 (n1060, n_23574, n_23575, n_23576, n_23577);
  and g56196 (n_23578, n_266, n_277);
  and g56197 (n_23579, n_255, n_130);
  and g56198 (n_23580, n_265, n_176);
  and g56199 (n_23581, n_150, n_88);
  and g56200 (n_23582, n_195, n_187, n1781, n2682);
  and g56201 (n_23583, n2635, n4215, n4232, n4247);
  and g56202 (n_23584, n2507, n2330, n541, n2241);
  and g56203 (n_23585, n_23578, n_23579, n_23580, n_23581);
  and g56204 (n4266, n_23582, n_23583, n_23584, n_23585);
  and g56205 (n_23586, n_183, n_206, n_180, n_291);
  and g56206 (n_23587, n116, n1237, n933, n244);
  and g56207 (n_23588, n3155, n4311, n13677, n790);
  and g56208 (n_23589, n1887, n4771, n12397, n13789);
  and g56209 (n26715, n_23586, n_23587, n_23588, n_23589);
  nor g56210 (n26722, n26716, n26717, n26718, n26719);
  nor g56211 (n5540, n5534, n5535, n5536, n5539);
  and g56212 (n_23590, n_102, n_122, n_144, n_61);
  and g56213 (n_23591, n_264, n_95, n_241, n1522);
  and g56214 (n_23592, n6604, n3159, n4101);
  and g56215 (n_23593, n690, n1391, n15854);
  and g56216 (n15867, n_23590, n_23591, n_23592, n_23593);
  and g56217 (n_23594, n_96, n_36);
  and g56218 (n_23595, n_278, n_157);
  and g56219 (n967, n960, n962, n_23594, n_23595);
  and g56220 (n_23596, n_274, n_135, n_280, n_161);
  and g56221 (n_23597, n_203, n_267, n_152, n_77);
  and g56222 (n_23598, n_170, n634, n720, n5148);
  and g56223 (n_23599, n6607, n6610, n1424, n1588);
  and g56224 (n6625, n_23596, n_23597, n_23598, n_23599);
  and g56225 (n_23600, n_274, n_268, n_283);
  and g56226 (n_23601, n_203, n_88, n_80);
  and g56227 (n_23602, n_196, n1367, n108);
  and g56228 (n_23603, n885, n437, n2091);
  and g56229 (n22748, n_23600, n_23601, n_23602, n_23603);
  and g56230 (n_23604, n_194, n_64, n_259, n_205);
  and g56231 (n_23605, n538, n418, n634, n2276);
  and g56232 (n_23606, n3163, n804, n14189, n4104);
  and g56233 (n_23607, n2809, n3206, n3858);
  and g56234 (n22762, n_23604, n_23605, n_23606, n_23607);
  and g56235 (n15956, n_58, n_270, n_49, n13671);
  and g56236 (n_23608, n_55, n_77);
  and g56237 (n1044, n_272, n570, n1040, n_23608);
  nor g56238 (n16314, n16308, n16309, n16310, n16313);
  and g56239 (n_23609, n_86, n_268);
  and g56240 (n_23610, n_36, n_40, n520, n1531);
  and g56241 (n_23611, n471, n291, n2346, n3290);
  and g56242 (n_23612, n916, n5296, n1621, n4216);
  and g56243 (n_23613, n24041, n1971, n5002, n_23609);
  and g56244 (n24057, n_23610, n_23611, n_23612, n_23613);
  nor g56245 (n24064, n24058, n24059, n24060, n24061);
  nor g56246 (n18337, n18331, n18332, n18333, n18336);
  nor g56247 (n22110, n22104, n22105, n22106, n22109);
  nor g56248 (n20881, n20875, n20876, n20877, n20880);
  nor g56249 (n15100, n15091, n15092, n15093, n15097);
  nor g56250 (n24913, n24907, n24908, n24909, n24912);
  and g56251 (n_23614, n_279, n_204, n_220);
  and g56252 (n_23615, n_268, n_62);
  and g56253 (n_23616, n_216, n_125);
  and g56254 (n_23617, n_131, n968);
  and g56255 (n976, n_23614, n_23615, n_23616, n_23617);
  and g56256 (n_23618, n_42, n_144);
  and g56257 (n_23619, n_63, n_258, n_57, n_262);
  and g56258 (n_23620, n418, n227, n978, n979);
  and g56259 (n_23621, n238, n294, n510, n988);
  and g56260 (n_23622, n989, n990, n992, n_23618);
  and g56261 (n1008, n_23619, n_23620, n_23621, n_23622);
  and g56262 (n_23623, n_103, n_180, n_85, n_203);
  and g56263 (n_23624, n_188, n_48, n747, n1009);
  and g56264 (n_23625, n244, n1020, n1024);
  and g56265 (n_23626, n405, n1025, n1029);
  and g56266 (n1039, n_23623, n_23624, n_23625, n_23626);
  nor g56267 (n4645, n4639, n4640, n4641, n4644);
  nor g56268 (n4436, n4430, n4431, n4432, n4433);
  and g56269 (n_23627, n_229, n_197, n_207, n_243);
  and g56270 (n_23628, n937, n896, n1100, n665);
  and g56271 (n_23629, n1119, n1126, n1154, n1155);
  and g56272 (n_23630, n1158, n776, n1160, n1163);
  and g56273 (n1178, n_23627, n_23628, n_23629, n_23630);
  and g56274 (n_23631, n_220, n_294);
  and g56275 (n2682, n_240, n128, n1121, n_23631);
  and g56276 (n_23632, n_86, n_138, n_230, n_46);
  and g56277 (n_23633, n_111, n515, n15924, n12909);
  and g56278 (n_23634, n12932, n13560, n204, n691);
  and g56279 (n_23635, n4269, n1611, n5748);
  and g56280 (n25157, n_23632, n_23633, n_23634, n_23635);
  nor g56281 (n25164, n25158, n25159, n25160, n25161);
  and g56282 (n_23636, n_228, n_134, n_224, n_218);
  and g56283 (n_23637, n_80, n_226, n_48, n4295);
  and g56284 (n_23638, n2738, n3464, n4298);
  and g56285 (n_23639, n4218, n1047, n2637);
  and g56286 (n4311, n_23636, n_23637, n_23638, n_23639);
  and g56287 (n1887, n_99, n_278, n_111, n_269);
  nor g56288 (n5378, n5372, n5373, n5374, n5377);
  nor g56289 (n6240, n6234, n6235, n6236, n6239);
  and g56290 (n_23640, n_256, n_198, n_100);
  and g56291 (n_23641, n_271, n_118);
  and g56292 (n_23642, n100, n279);
  and g56293 (n_23643, n918, n2191);
  and g56294 (n6604, n_23640, n_23641, n_23642, n_23643);
  and g56295 (n_23644, n_228, n_75);
  and g56296 (n5148, n_37, n_39, n1183, n_23644);
  and g56297 (n6610, n_204, n_261, n_263, n1824);
  nor g56298 (n16529, n16523, n16524, n16525, n16528);
  and g56299 (n_23645, n_110, n_166, n_205);
  and g56300 (n_23646, n_117, n_128, n_37);
  and g56301 (n_23647, n_48, n665, n1103);
  and g56302 (n_23648, n1604, n2508);
  and g56303 (n5296, n_23645, n_23646, n_23647, n_23648);
  and g56304 (n_23649, n_191, n_145);
  and g56305 (n1621, n_283, n_147, n_245, n_23649);
  nor g56306 (n17349, n17343, n17344, n17345, n17348);
  nor g56307 (n19552, n19546, n19547, n19548, n19551);
  nor g56308 (n15715, n15709, n15710, n15711, n15712);
  nor g56309 (n16177, n16171, n16172, n16173, n16176);
  nor g56310 (n24458, n24452, n24453, n24454, n24457);
  nor g56311 (n23937, n23931, n23932, n23933, n23936);
  nor g56312 (n4868, n4862, n4863, n4864, n4865);
  and g56313 (n_23650, n_160, n_248, n1128);
  and g56314 (n_23651, n654, n1129, n1131);
  and g56315 (n_23652, n936, n1132, n1135);
  and g56316 (n_23653, n1138, n1140, n1143);
  and g56317 (n1154, n_23650, n_23651, n_23652, n_23653);
  and g56318 (n_23654, n_234, n_268, n_258, n_153);
  and g56319 (n_23655, n634, n2467, n1781, n1063);
  and g56320 (n_23656, n1183, n1264, n622, n247);
  and g56321 (n_23657, n14572, n12812, n13249);
  and g56322 (n15924, n_23654, n_23655, n_23656, n_23657);
  nor g56323 (n5924, n5918, n5919, n5920, n5923);
  nor g56324 (n6384, n6378, n6379, n6380, n6383);
  nor g56325 (n17819, n17813, n17814, n17815, n17818);
  nor g56326 (n20899, n20893, n20894, n20895, n20898);
  nor g56327 (n16924, n16918, n16919, n16920, n16923);
  and g56328 (n1135, n_255, n_205, n_49, n_131);
  and g56329 (n_23658, n_233, n_282, n_123);
  and g56330 (n_23659, n_207, n1252, n1253);
  and g56331 (n_23660, n1254, n734);
  and g56332 (n_23661, n814, n1255);
  and g56333 (n1264, n_23658, n_23659, n_23660, n_23661);
  nor g56334 (n5628, n5622, n5623, n5624, n5627);
  nor g56335 (n16331, n16325, n16326, n16327, n16330);
  nor g56336 (n16346, n16340, n16341, n16342, n16345);
  nor g56337 (n20917, n20911, n20912, n20913, n20916);
  nor g56338 (n18415, n18409, n18410, n18411, n18414);
  and g56339 (n_23662, n_219, n_40, n_157, n_245);
  and g56340 (n_23663, n3252, n247, n1523, n15061);
  and g56341 (n_23664, n12404, n14381, n6667);
  and g56342 (n_23665, n6102, n137, n3192);
  and g56343 (n15074, n_23662, n_23663, n_23664, n_23665);
  nor g56344 (n24517, n24511, n24512, n24513, n24516);
  nor g56345 (n25666, n25660, n25661, n25662, n25665);
  and g56346 (n_23666, n_122, n_72, n_242, n_165);
  and g56347 (n_23667, n_213, n1180, n1181, n1202);
  and g56348 (n_23668, n1211, n802, n1154, n1216);
  and g56349 (n_23669, n1219, n982, n1221);
  and g56350 (n1235, n_23666, n_23667, n_23668, n_23669);
  and g56351 (n_23670, n_71, n_168);
  and g56352 (n_23671, n_256, n_110, n_258, n_40);
  and g56353 (n_23672, n1182, n491, n4293, n4311);
  and g56354 (n_23673, n4325, n2169, n2740, n4332);
  and g56355 (n_23674, n4334, n3114, n4335, n_23670);
  and g56356 (n4351, n_23671, n_23672, n_23673, n_23674);
  and g56357 (n_23675, n_136, n_94);
  and g56358 (n_23676, n_114, n_222, n_98, n_167);
  and g56359 (n_23677, n_254, n2467, n423, n1576);
  and g56360 (n_23678, n4767, n4785, n1928, n4815);
  and g56361 (n_23679, n4827, n1973, n4828, n_23675);
  and g56362 (n4844, n_23676, n_23677, n_23678, n_23679);
  nor g56363 (n4987, n4981, n4982, n4983, n4986);
  nor g56364 (n6223, n6217, n6218, n6219, n6222);
  nor g56365 (n16498, n16492, n16493, n16494, n16497);
  nor g56366 (n16513, n16507, n16508, n16509, n16512);
  nor g56367 (n17333, n17327, n17328, n17329, n17332);
  nor g56368 (n20935, n20929, n20930, n20931, n20934);
  nor g56369 (n20989, n20983, n20984, n20985, n20988);
  nor g56370 (n19570, n19564, n19565, n19566, n19569);
  and g56371 (n_23680, n_217, n_122);
  and g56372 (n_23681, n_238, n_290);
  and g56373 (n_23682, n_52, n_164, n_124, n_216);
  and g56374 (n_23683, n_291, n_200, n1180, n2778);
  and g56375 (n_23684, n5785, n3675, n3743, n1894);
  and g56376 (n_23685, n1185, n2349, n_23680, n_23681);
  and g56377 (n15283, n_23682, n_23683, n_23684, n_23685);
  nor g56378 (n15731, n15725, n15726, n15727, n15728);
  nor g56379 (n18432, n18426, n18427, n18428, n18431);
  and g56380 (n_23686, n_177, n1389, n15047);
  and g56381 (n_23687, n1781, n294, n2591);
  and g56382 (n_23688, n12810, n15050, n2241);
  and g56383 (n_23689, n370, n3194, n13827);
  and g56384 (n15061, n_23686, n_23687, n_23688, n_23689);
  and g56385 (n6667, n_53, n_129, n827, n6664);
  and g56386 (n_23690, n_202, n_258);
  and g56387 (n_23691, n_265, n_76);
  and g56388 (n6102, n590, n_287, n_23690, n_23691);
  nor g56389 (n24945, n24939, n24940, n24941, n24944);
  nor g56390 (n26194, n26188, n26189, n26190, n26193);
  and g56391 (n_23692, n_151, n_294);
  and g56392 (n_23693, n_88, n_149);
  and g56393 (n1211, n1204, n1206, n_23692, n_23693);
  and g56394 (n1219, n_103, n_129, n_61, n_227);
  and g56395 (n_23694, n_204, n_227);
  and g56396 (n_23695, n_141, n_174, n_93, n285);
  and g56397 (n_23696, n2698, n774, n4356, n4366);
  and g56398 (n_23697, n4388, n4405, n1785, n992);
  and g56399 (n_23698, n1346, n2014, n3416, n_23694);
  and g56400 (n4421, n_23695, n_23696, n_23697, n_23698);
  and g56401 (n_23699, n_251, n_252);
  and g56402 (n_23700, n_212, n2073);
  and g56403 (n4332, n2371, n4327, n_23699, n_23700);
  and g56404 (n_23701, n_255, n_234);
  and g56405 (n_23702, n_148, n_250);
  and g56406 (n_23703, n_50, n_243);
  and g56407 (n4767, n3043, n_23701, n_23702, n_23703);
  and g56408 (n_23704, n_104, n_259, n_116, n_59);
  and g56409 (n_23705, n4101, n2583, n1827, n3252);
  and g56410 (n_23706, n968, n874, n1181, n141);
  and g56411 (n_23707, n4769, n2361, n4771);
  and g56412 (n4785, n_23704, n_23705, n_23706, n_23707);
  nor g56413 (n4855, n4849, n4850, n4851, n4852);
  and g56414 (n_23708, n_162, n_220);
  and g56415 (n_23709, n_201, n_180);
  and g56416 (n_23710, n_248, n_56, n_148, n_68);
  and g56417 (n_23711, n1237, n937, n1245, n1291);
  and g56418 (n_23712, n1292, n1305, n1345, n830);
  and g56419 (n_23713, n1346, n1347, n_23708, n_23709);
  and g56420 (n1364, n_23710, n_23711, n_23712, n_23713);
  nor g56421 (n5908, n5902, n5903, n5904, n5907);
  nor g56422 (n5450, n5444, n5445, n5446, n5449);
  nor g56423 (n6432, n6426, n6427, n6428, n6431);
  nor g56424 (n17464, n17458, n17459, n17460, n17463);
  nor g56425 (n20971, n20965, n20966, n20967, n20970);
  nor g56426 (n20953, n20947, n20948, n20949, n20952);
  nor g56427 (n16908, n16902, n16903, n16904, n16907);
  and g56428 (n_23714, n_266, n_204, n_285, n_54);
  and g56429 (n_23715, n_282, n_172, n_60);
  and g56430 (n_23716, n508, n439, n3548);
  and g56431 (n_23717, n1070, n1738, n3645);
  and g56432 (n15047, n_23714, n_23715, n_23716, n_23717);
  and g56433 (n15050, n_89, n_126, n2651, n14479);
  and g56434 (n_23718, n_229, n_158);
  and g56435 (n_23719, n_195, n_118);
  and g56436 (n4356, n_296, n1669, n_23718, n_23719);
  and g56437 (n_23720, n_164, n_95, n_269);
  and g56438 (n_23721, n_74, n_106, n_90);
  and g56439 (n_23722, n1040, n4357);
  and g56440 (n_23723, n1135, n2334);
  and g56441 (n4366, n_23720, n_23721, n_23722, n_23723);
  and g56442 (n_23724, n_102, n_136, n_73, n_283);
  and g56443 (n_23725, n_123, n_82, n_179, n_187);
  and g56444 (n_23726, n1550, n3378, n4375);
  and g56445 (n_23727, n439, n1272, n4234);
  and g56446 (n4388, n_23724, n_23725, n_23726, n_23727);
  and g56447 (n_23728, n_144, n_240);
  and g56448 (n_23729, n_242, n_37);
  and g56449 (n_23730, n_248, n_239, n_212, n_77);
  and g56450 (n_23731, n_153, n_254, n590, n978);
  and g56451 (n_23732, n827, n1330, n615, n2296);
  and g56452 (n_23733, n793, n3296, n_23728, n_23729);
  and g56453 (n4405, n_23730, n_23731, n_23732, n_23733);
  and g56454 (n_23734, n_231, n_280);
  and g56455 (n_23735, n_117, n_197);
  and g56456 (n_23736, n_70, n_188, n_296, n1247);
  and g56457 (n_23737, n1248, n285, n235, n1251);
  and g56458 (n_23738, n1264, n1268, n1103, n1271);
  and g56459 (n_23739, n1272, n1274, n_23734, n_23735);
  and g56460 (n1291, n_23736, n_23737, n_23738, n_23739);
  and g56461 (n_23740, n_87, n_95, n_39, n_141);
  and g56462 (n_23741, n_113, n_262, n1313);
  and g56463 (n_23742, n731, n1323, n1328);
  and g56464 (n_23743, n1329, n1331, n1333);
  and g56465 (n1345, n_23740, n_23741, n_23742, n_23743);
  nor g56466 (n5612, n5606, n5607, n5608, n5611);
  nor g56467 (n25004, n24998, n24999, n25000, n25003);
  nor g56468 (n25698, n25692, n25693, n25694, n25697);
  and g56469 (n_23744, n_184, n_69, n_59);
  and g56470 (n_23745, n4367, n2807);
  and g56471 (n_23746, n2013, n4153);
  and g56472 (n_23747, n876, n2210);
  and g56473 (n4375, n_23744, n_23745, n_23746, n_23747);
  and g56474 (n_23748, n_168, n_54);
  and g56475 (n1268, n_221, n244, n_283, n_23748);
  and g56476 (n_23749, n_137, n_138);
  and g56477 (n_23750, n_119, n_244);
  and g56478 (n1313, n_297, n1308, n_23749, n_23750);
  and g56479 (n_23751, n_183, n_251);
  and g56480 (n1328, n_199, n_52, n1324, n_23751);
  nor g56481 (n5121, n5115, n5116, n5117, n5118);
  nor g56482 (n5968, n5962, n5963, n5964, n5967);
  nor g56483 (n21035, n21029, n21030, n21031, n21034);
  nor g56484 (n19588, n19582, n19583, n19584, n19587);
  and g56485 (n_23752, n_145, n_277);
  and g56486 (n_23753, n_279, n_193);
  and g56487 (n_23754, n_67, n_95);
  and g56488 (n_23755, n_262, n4101);
  and g56489 (n_23756, n202, n1783, n730, n285);
  and g56490 (n_23757, n1183, n1915, n512, n503);
  and g56491 (n_23758, n15061, n1709, n13012, n15286);
  and g56492 (n_23759, n_23752, n_23753, n_23754, n_23755);
  and g56493 (n15305, n_23756, n_23757, n_23758, n_23759);
  nor g56494 (n18450, n18444, n18445, n18446, n18449);
  and g56495 (n_23760, n_45, n_267, n_172, n_80);
  and g56496 (n_23761, n_211, n_226, n1269, n1366);
  and g56497 (n_23762, n1378, n1407, n1419, n1422);
  and g56498 (n_23763, n1423, n1456, n1458);
  and g56499 (n1472, n_23760, n_23761, n_23762, n_23763);
  nor g56500 (n6364, n6358, n6359, n6360, n6363);
  nor g56501 (n6941, n6935, n6936, n6937, n6940);
  nor g56502 (n15363, n15357, n15358, n15359, n15360);
  nor g56503 (n17481, n17475, n17476, n17477, n17480);
  nor g56504 (n20298, n20292, n20293, n20294, n20297);
  nor g56505 (n21052, n21046, n21047, n21048, n21051);
  nor g56506 (n22042, n22036, n22037, n22038, n22041);
  nor g56507 (n7108, n7102, n7103, n7104, n7107);
  nor g56508 (n26163, n26157, n26158, n26159, n26162);
  nor g56509 (n25757, n25751, n25752, n25753, n25756);
  and g56510 (n_23764, n_127, n_278);
  and g56511 (n_23765, n_81, n_38);
  and g56512 (n_23766, n1367, n1369);
  and g56513 (n1378, n1372, n_23764, n_23765, n_23766);
  and g56514 (n_23767, n_246, n_108, n_90, n_196);
  and g56515 (n_23768, n1128, n1180, n1379, n1384);
  and g56516 (n_23769, n1387, n1388, n1391);
  and g56517 (n_23770, n846, n1392, n1394);
  and g56518 (n1407, n_23767, n_23768, n_23769, n_23770);
  and g56519 (n_23771, n_136, n_256, n_35);
  and g56520 (n_23772, n_83, n_205, n_150);
  and g56521 (n_23773, n_111, n_263, n789);
  and g56522 (n_23774, n1408, n1409);
  and g56523 (n1419, n_23771, n_23772, n_23773, n_23774);
  and g56524 (n1422, n_168, n_257, n_160, n_208);
  and g56525 (n_23775, n_182, n_145);
  and g56526 (n_23776, n_143, n_280);
  and g56527 (n_23777, n_190, n_116);
  and g56528 (n_23778, n_239, n_210);
  and g56529 (n_23779, n_111, n418);
  and g56530 (n_23780, n116, n508);
  and g56531 (n_23781, n5013, n5082, n2170, n5085);
  and g56532 (n_23782, n3094, n811, n789, n3663);
  and g56533 (n_23783, n1012, n1107, n_23775, n_23776);
  and g56534 (n_23784, n_23777, n_23778, n_23779, n_23780);
  and g56535 (n5106, n_23781, n_23782, n_23783, n_23784);
  nor g56536 (n5143, n5135, n5136, n5137, n5140);
  nor g56537 (n5565, n5557, n5558, n5559, n5562);
  nor g56538 (n5592, n5586, n5587, n5588, n5591);
  and g56539 (n_23785, n_238, n_116, n_37, n_40);
  and g56540 (n_23786, n_232, n_79, n_38, n1237);
  and g56541 (n_23787, n14479, n15330, n12973, n15337);
  and g56542 (n_23788, n1759, n2809, n475, n1530);
  and g56543 (n15352, n_23785, n_23786, n_23787, n_23788);
  and g56544 (n_23789, n_94, n_35);
  and g56545 (n_23790, n_61, n_175, n_80, n116);
  and g56546 (n_23791, n356, n288, n15743, n14386);
  and g56547 (n_23792, n4815, n688, n2091, n2262);
  and g56548 (n_23793, n2807, n2784, n3162, n_23789);
  and g56549 (n15759, n_23790, n_23791, n_23792, n_23793);
  nor g56550 (n15768, n15760, n15761, n15762, n15765);
  nor g56551 (n20315, n20309, n20310, n20311, n20314);
  nor g56552 (n7274, n7268, n7269, n7270, n7273);
  and g56553 (n1372, n_274, n_100, n_128, n_210);
  and g56554 (n1387, n_164, n_268, n_146, n_271);
  and g56555 (n_23794, n_34, n_58, n_88, n_177);
  and g56556 (n_23795, n_272, n1237, n827, n896);
  and g56557 (n_23796, n1139, n1435, n604, n1437);
  and g56558 (n_23797, n1438, n1065, n1440);
  and g56559 (n1454, n_23794, n_23795, n_23796, n_23797);
  and g56560 (n_23798, n_229, n_73, n_291, n_263);
  and g56561 (n_23799, n5013, n5034, n2979, n1610);
  and g56562 (n_23800, n4332, n4216, n5036);
  and g56563 (n_23801, n5038, n812, n5040);
  and g56564 (n5053, n_23798, n_23799, n_23800, n_23801);
  and g56565 (n_23802, n_279, n_201, n_259);
  and g56566 (n_23803, n_127, n_128, n1237);
  and g56567 (n_23804, n421, n3886, n3438);
  and g56568 (n_23805, n4357, n2546, n5002);
  and g56569 (n5013, n_23802, n_23803, n_23804, n_23805);
  and g56570 (n_23806, n_182, n_65, n_221, n_75);
  and g56571 (n_23807, n_190, n1379, n288, n1475);
  and g56572 (n_23808, n1476, n1511, n631, n1521);
  and g56573 (n_23809, n1549, n1555, n1556, n1557);
  and g56574 (n1572, n_23806, n_23807, n_23808, n_23809);
  and g56575 (n_23810, n_151, n_221);
  and g56576 (n_23811, n_257, n_270, n_119, n_215);
  and g56577 (n_23812, n_287, n770, n2484, n1915);
  and g56578 (n_23813, n1585, n3651, n1635, n5148);
  and g56579 (n_23814, n921, n5150, n5152, n_23810);
  and g56580 (n5168, n_23811, n_23812, n_23813, n_23814);
  nor g56581 (n6205, n6199, n6200, n6201, n6204);
  and g56582 (n_23815, n_219, n_290);
  and g56583 (n_23816, n_123, n_60);
  and g56584 (n_23817, n_152, n1692);
  and g56585 (n15330, n15324, n_23815, n_23816, n_23817);
  and g56586 (n_23818, n_280, n_99);
  and g56587 (n_23819, n_74, n_77);
  and g56588 (n_23820, n_90, n_262);
  and g56589 (n_23821, n_297, n3380);
  and g56590 (n15337, n_23818, n_23819, n_23820, n_23821);
  and g56591 (n_23822, n_253, n_256);
  and g56592 (n1759, n_268, n_84, n1755, n_23822);
  and g56593 (n_23823, n_137, n_129);
  and g56594 (n_23824, n_58, n_176);
  and g56595 (n15743, n_118, n12830, n_23823, n_23824);
  and g56596 (n_23825, n_182, n_216);
  and g56597 (n2262, n_95, n618, n1827, n_23825);
  nor g56598 (n21070, n21064, n21065, n21066, n21069);
  nor g56599 (n22028, n22022, n22023, n22024, n22027);
  nor g56600 (n19606, n19600, n19601, n19602, n19605);
  nor g56601 (n18468, n18462, n18463, n18464, n18467);
  nor g56602 (n_23826, n26107, n26108);
  nor g56603 (n_23827, n26114, n26115);
  nor g56604 (n_23828, n26116, n26117);
  and g56605 (n26123, \a[2] , n_23826, n_23827, n_23828);
  and g56606 (n_23829, n_92, n_36);
  and g56607 (n_23830, n_218, n1063);
  and g56608 (n_23831, n1424, n1219);
  and g56609 (n_23832, n1425, n1428);
  and g56610 (n1435, n_23829, n_23830, n_23831, n_23832);
  nor g56611 (n5888, n5882, n5883, n5884, n5887);
  and g56612 (n_23833, n_92, n_258, n_165, n_119);
  and g56613 (n_23834, n_172, n_289, n_46, n_50);
  and g56614 (n_23835, n3163, n5019, n811);
  and g56615 (n_23836, n5021, n1331, n1861);
  and g56616 (n5034, n_23833, n_23834, n_23835, n_23836);
  and g56617 (n_23837, n_100, n_208);
  and g56619 (n_23839, n294, n1603);
  and g56620 (n1610, n1604, n_23837, n_22764, n_23839);
  and g56621 (n_23840, n_168, n_132);
  and g56622 (n_23841, n_243, n235);
  and g56623 (n_23842, n873, n1181);
  and g56624 (n_23843, n1577, n1578);
  and g56625 (n1585, n_23840, n_23841, n_23842, n_23843);
  and g56626 (n_23844, n_204, n_110, n_246, n_201);
  and g56627 (n_23845, n_161, n_203, n_167, n_195);
  and g56628 (n_23846, n_226, n_126, n1602, n1610);
  and g56629 (n_23847, n1615, n1617, n1621);
  and g56630 (n1635, n_23844, n_23845, n_23846, n_23847);
  nor g56631 (n6348, n6342, n6343, n6344, n6347);
  nor g56632 (n6925, n6919, n6920, n6921, n6924);
  and g56633 (n_23848, n_246, n_294, n_186, n_132);
  and g56634 (n_23849, n_78, n2346, n15312);
  and g56635 (n_23850, n1725, n5085, n12431);
  and g56636 (n_23851, n2468, n365, n1329);
  and g56637 (n15324, n_23848, n_23849, n_23850, n_23851);
  nor g56638 (n17499, n17493, n17494, n17495, n17498);
  and g56639 (n_23852, n_182, n_168);
  and g56640 (n_23853, n_35, n_261, n_291, n_126);
  and g56641 (n_23854, n454, n230, n556, n1039);
  and g56642 (n_23855, n6026, n13221, n2422, n2808);
  and g56643 (n_23856, n2704, n1073, n3042, n_23852);
  and g56644 (n15785, n_23853, n_23854, n_23855, n_23856);
  nor g56645 (n15795, n15786, n15787, n15788, n15792);
  nor g56646 (n7091, n7085, n7086, n7087, n7090);
  and g56647 (n_23857, n_53, n_151);
  and g56648 (n_23858, n_44, n_180);
  and g56649 (n_23859, n_49, n_159);
  and g56650 (n5019, n1709, n_23857, n_23858, n_23859);
  and g56651 (n_23860, n_136, n_290);
  and g56653 (n_23138, n_230, n_150);
  and g56654 (n_23863, n_78, n359);
  and g56655 (n_23864, n1574, n1248, n745, n423);
  and g56656 (n_23865, n1575, n1600, n1601, n1635);
  and g56657 (n_23866, n1640, n1643, n1644, n1646);
  and g56658 (n_23867, n_23860, n_22840, n_23138, n_23863);
  and g56659 (n1665, n_23864, n_23865, n_23866, n_23867);
  and g56661 (n_23869, n_63, n_224, n_227, n_171);
  and g56662 (n_23870, n_46, n590, n1182, n1719);
  and g56663 (n_23871, n1725, n774, n1754, n1759);
  and g56664 (n_23872, n694, n1760, n1763, n_23551);
  and g56665 (n1779, n_23869, n_23870, n_23871, n_23872);
  nor g56666 (n5573, n5567, n5568, n5569, n5572);
  and g56667 (n_23873, n_186, n_248);
  and g56668 (n1615, n_149, n_296, n1611, n_23873);
  and g56669 (n_23874, n_231, n_259);
  and g56670 (n_23875, n_184, n_111);
  and g56671 (n_23876, n_179, n1557);
  and g56672 (n15312, n2209, n_23874, n_23875, n_23876);
  and g56673 (n_23877, n_153, n_296);
  and g56674 (n1725, n_48, n1294, n1721, n_23877);
  nor g56675 (n22011, n22005, n22006, n22007, n22010);
  nor g56676 (n19624, n19618, n19619, n19620, n19623);
  and g56677 (n_23878, n_137, n1680);
  and g56678 (n_23879, n_198, n_146);
  and g56679 (n_23880, n2556, n1727);
  and g56680 (n6026, n2705, n_23878, n_23879, n_23880);
  and g56681 (n_23881, n_238, n_199);
  and g56682 (n_23882, n_294, n_75);
  and g56683 (n2422, n_248, n_289, n_23881, n_23882);
  nor g56684 (n7146, n7140, n7141, n7142, n7145);
  nor g56685 (n26132, n26126, n26127, n26128, n26131);
  nor g56686 (n5335, n5329, n5330, n5331, n5332);
  and g56687 (n_23883, n_117, n_55, n_250, n_105);
  and g56688 (n_23884, n156, n731, n1576);
  and g56689 (n_23885, n120, n1480, n1585);
  and g56690 (n_23886, n1586, n1428, n1588);
  and g56691 (n1600, n_23883, n_23884, n_23885, n_23886);
  and g56692 (n_23887, n_103, n_165);
  and g56693 (n1640, n_244, n_111, n1636, n_23887);
  and g56694 (n1643, n_274, n_134, n_142, n_187);
  and g56695 (n_23888, n_53, n_99, n_76);
  and g56696 (n_23889, n_264, n_82, n_118);
  and g56697 (n_23890, n_77, n1161, n1708);
  and g56698 (n_23891, n1329, n1709);
  and g56699 (n1719, n_23888, n_23889, n_23890, n_23891);
  and g56700 (n_23892, n_233, n_57, n_291, n_55);
  and g56701 (n_23893, n_188, n_146, n227, n1726);
  and g56702 (n_23894, n1731, n1735, n1372, n1737);
  and g56703 (n_23895, n1738, n1739, n1740);
  and g56704 (n1754, n_23892, n_23893, n_23894, n_23895);
  nor g56705 (n6189, n6183, n6184, n6185, n6188);
  nor g56706 (n7990, n7984, n7985, n7986, n7989);
  nor g56707 (n18486, n18480, n18481, n18482, n18485);
  nor g56708 (n5858, n5852, n5853, n5854, n5855);
  nor g56709 (n6455, n6449, n6450, n6451, n6454);
  nor g56710 (n17517, n17511, n17512, n17513, n17516);
  nor g56711 (n19642, n19636, n19637, n19638, n19641);
  nor g56712 (n19742, n19736, n19737, n19738, n19741);
  nor g56713 (n19696, n19690, n19691, n19692, n19695);
  and g56714 (n_23896, n_266, n_251, n_54, n_250);
  and g56715 (n_23897, n_113, n1040, n4295, n1475);
  and g56716 (n_23898, n874, n15330, n2555, n1754);
  and g56717 (n_23899, n1604, n2607, n3987);
  and g56718 (n15810, n_23896, n_23897, n_23898, n_23899);
  nor g56719 (n15820, n15811, n15812, n15813, n15817);
  nor g56720 (n19660, n19654, n19655, n19656, n19659);
  nor g56721 (n19759, n19753, n19754, n19755, n19758);
  nor g56722 (n19678, n19672, n19673, n19674, n19677);
  and g56723 (n_23900, n_92, n_163, n_129);
  and g56724 (n_23901, n_117, n_244, n_106);
  and g56725 (n_23902, n2170, n2544);
  and g56726 (n_23903, n2427, n2546);
  and g56727 (n2555, n_23900, n_23901, n_23902, n_23903);
  nor g56728 (n7619, n7613, n7614, n7615, n7618);
  nor g56729 (n8401, n8395, n8396, n8397, n8400);
  nor g56730 (n7256, n7250, n7251, n7252, n7255);
  and g56731 (n_23904, n_103, n_117);
  and g56732 (n_23905, n_95, n_77, n1040, n399);
  and g56733 (n_23906, n282, n533, n1781, n1531);
  and g56734 (n_23907, n1794, n1814, n1819, n1823);
  and g56735 (n_23908, n776, n1859, n1861, n_23904);
  and g56736 (n1877, n_23905, n_23906, n_23907, n_23908);
  and g56737 (n_23909, n_182, n_145, n_255, n_73);
  and g56738 (n_23910, n_83, n_142, n5171, n_241);
  and g56739 (n_23911, n5188, n5193, n5224, n5233);
  and g56740 (n_23912, n5239, n1819, n636, n5066);
  and g56741 (n5254, n_23909, n_23910, n_23911, n_23912);
  and g56742 (n_23913, n_114, n_242);
  and g56743 (n_23914, n_58, n_227);
  and g56744 (n_23915, n_154, n_57, n_39, n_152);
  and g56745 (n_23916, n570, n108, n2633, n5746);
  and g56746 (n_23917, n3205, n5239, n824, n5269);
  and g56747 (n_23918, n658, n5748, n_23913, n_23914);
  and g56748 (n5765, n_23915, n_23916, n_23917, n_23918);
  nor g56749 (n5988, n5982, n5983, n5984, n5987);
  nor g56750 (n6011, n6003, n6004, n6005, n6008);
  nor g56751 (n19099, n19093, n19094, n19095, n19098);
  nor g56752 (n20375, n20369, n20370, n20371, n20374);
  nor g56753 (n7973, n7967, n7968, n7969, n7972);
  nor g56754 (n18504, n18498, n18499, n18500, n18503);
  and g56755 (n_23919, n_276, n_136);
  and g56756 (n_23920, n_128, n_74);
  and g56757 (n1819, n_200, n_250, n_23919, n_23920);
  and g56758 (n_23921, n_182, n_67);
  and g56759 (n_23922, n_123, n_270, n_172, n_141);
  and g56760 (n_23923, n100, n5286, n615, n1254);
  and g56761 (n_23924, n5296, n247, n1577, n5304);
  and g56762 (n_23925, n3312, n2627, n3264, n_23921);
  and g56763 (n5320, n_23922, n_23923, n_23924, n_23925);
  and g56764 (n_23926, n_122, n_135, n_72, n_283);
  and g56765 (n_23927, n_249, n_87, n_175, n_232);
  and g56766 (n_23928, n3163, n356, n654, n512);
  and g56767 (n_23929, n4356, n897, n2278, n5173);
  and g56768 (n5188, n_23926, n_23927, n_23928, n_23929);
  and g56769 (n_23930, n_53, n_218);
  and g56770 (n_23931, n_125, n_106);
  and g56771 (n_23932, n_90, n1732);
  and g56772 (n5239, n2133, n_23930, n_23931, n_23932);
  and g56773 (n_23933, n_102, n_71);
  and g56774 (n_23934, n_96, n_132);
  and g56775 (n5269, n634, n937, n_23933, n_23934);
  and g56776 (n_23935, n_238, n_264, n_178, n_239);
  and g56777 (n_23936, n_289, n1884, n1890, n1893);
  and g56778 (n_23937, n1476, n1601, n1039, n1211);
  and g56779 (n_23938, n1345, n1697, n1896, n1898);
  and g56780 (n1913, n_23935, n_23936, n_23937, n_23938);
  nor g56781 (n6328, n6322, n6323, n6324, n6327);
  nor g56782 (n6907, n6901, n6902, n6903, n6906);
  nor g56783 (n17535, n17529, n17530, n17531, n17534);
  nor g56784 (n19116, n19110, n19111, n19112, n19115);
  nor g56785 (n19777, n19771, n19772, n19773, n19776);
  nor g56786 (n20392, n20386, n20387, n20388, n20391);
  and g56787 (n_23939, n_110, n_35);
  and g56788 (n_23940, n_258, n_195, n_157, n_211);
  and g56789 (n_23941, n15826, n1531, n1475, n1916);
  and g56790 (n_23942, n6707, n6769, n3415, n3219);
  and g56791 (n_23943, n12428, n1272, n1586, n_23939);
  and g56792 (n15842, n_23940, n_23941, n_23942, n_23943);
  nor g56793 (n15851, n15843, n15844, n15845, n15848);
  nor g56794 (n7071, n7065, n7066, n7067, n7070);
  and g56795 (n_23944, n_214, n_52, n_129, n_189);
  and g56796 (n_23945, n_115, n_297, n621, n1575);
  and g56797 (n_23946, n2346, n872, n873, n5264);
  and g56798 (n_23947, n5269, n593, n3268, n5271);
  and g56799 (n5286, n_23944, n_23945, n_23946, n_23947);
  and g56800 (n_23948, n_155, n_228, n_144);
  and g56801 (n_23949, n_274, n_259);
  and g56802 (n_23950, n_111, n_254);
  and g56803 (n_23951, n_50, n1248);
  and g56804 (n5304, n_23948, n_23949, n_23950, n_23951);
  and g56805 (n1890, n_43, n_114, n_267, n1887);
  and g56806 (n1893, n_73, n_124, n_47, n_117);
  and g56807 (n_23952, n_86, n_206);
  and g56808 (n_23953, n_142, n_159);
  and g56809 (n15826, n202, n877, n_23952, n_23953);
  nor g56810 (n7603, n7597, n7598, n7599, n7602);
  nor g56811 (n7240, n7234, n7235, n7236, n7239);
  and g56812 (n_23954, n_137, n_121);
  and g56813 (n_23955, n_190, n_223);
  and g56814 (n_23956, n_123, n_203);
  and g56815 (n_23957, n_112, n_226);
  and g56816 (n_23958, n1574, n515, n1915, n1916);
  and g56817 (n_23959, n1917, n1925, n1958, n1969);
  and g56818 (n_23960, n877, n658, n1971, n1973);
  and g56819 (n_23961, n_23954, n_23955, n_23956, n_23957);
  and g56820 (n1992, n_23958, n_23959, n_23960, n_23961);
  nor g56821 (n21130, n21124, n21125, n21126, n21129);
  nor g56822 (n7664, n7658, n7659, n7660, n7663);
  nor g56823 (n9338, n9332, n9333, n9334, n9337);
  nor g56824 (n8834, n8828, n8829, n8830, n8833);
  nor g56825 (n18522, n18516, n18517, n18518, n18521);
  nor g56826 (n6891, n6885, n6886, n6887, n6890);
  nor g56827 (n17553, n17547, n17548, n17549, n17552);
  nor g56828 (n20410, n20404, n20405, n20406, n20409);
  nor g56829 (n21147, n21141, n21142, n21143, n21146);
  nor g56830 (n21943, n21937, n21938, n21939, n21942);
  and g56831 (n_23962, n_163, n_290);
  and g56832 (n_23963, n_166, n_207);
  and g56833 (n_23964, n_78, n_156, n15867, n202);
  and g56834 (n_23965, n2583, n1129, n1915, n15880);
  and g56835 (n_23966, n2703, n14210, n6517, n15882);
  and g56836 (n_23967, n1274, n2742, n_23962, n_23963);
  and g56837 (n15899, n_23964, n_23965, n_23966, n_23967);
  nor g56838 (n15909, n15900, n15901, n15902, n15906);
  nor g56839 (n7055, n7049, n7050, n7051, n7054);
  nor g56840 (n5841, n5835, n5836, n5837, n5838);
  and g56841 (n_23968, n_155, n_43, n_257, n_213);
  and g56842 (n_23969, n570, n193, n937, n2573);
  and g56843 (n_23970, n3990, n6707, n5190);
  and g56844 (n_23971, n4011, n2209, n14518);
  and g56845 (n15880, n_23968, n_23969, n_23970, n_23971);
  and g56846 (n6517, n_253, n_76, n_56, n5171);
  nor g56847 (n9856, n9850, n9851, n9852, n9855);
  nor g56848 (n8381, n8375, n8376, n8377, n8380);
  nor g56849 (n7169, n7163, n7164, n7165, n7168);
  nor g56850 (n6150, n6144, n6145, n6146, n6147);
  nor g56851 (n11038, n11032, n11033, n11034, n11037);
  nor g56852 (n18622, n18616, n18617, n18618, n18621);
  nor g56853 (n21165, n21159, n21160, n21161, n21164);
  nor g56854 (n21929, n21923, n21924, n21925, n21928);
  nor g56855 (n7955, n7949, n7950, n7951, n7954);
  nor g56856 (n9321, n9315, n9316, n9317, n9320);
  nor g56857 (n8818, n8812, n8813, n8814, n8817);
  nor g56858 (n18540, n18534, n18535, n18536, n18539);
  and g56859 (n_23972, n_92, n_169);
  and g56860 (n_23973, n_246, n_100);
  and g56861 (n_23974, n_138, n_197, n_55, n_273);
  and g56862 (n_23975, n_272, n520, n2940, n2651);
  and g56863 (n_23976, n5773, n616, n4388, n5806);
  and g56864 (n_23977, n2990, n5808, n_23972, n_23973);
  and g56865 (n5825, n_23974, n_23975, n_23976, n_23977);
  nor g56866 (n6483, n6475, n6476, n6477, n6480);
  nor g56867 (n6873, n6867, n6868, n6869, n6872);
  nor g56868 (n17571, n17565, n17566, n17567, n17570);
  nor g56869 (n18639, n18633, n18634, n18635, n18638);
  and g56870 (n_23978, n_54, n_221, n_67, n_171);
  and g56871 (n_23979, n_241, n_296, n_93, n978);
  and g56872 (n_23980, n731, n15924, n13041, n12805);
  and g56873 (n_23981, n2022, n1798, n2442);
  and g56874 (n15938, n_23978, n_23979, n_23980, n_23981);
  nor g56875 (n15948, n15939, n15940, n15941, n15945);
  nor g56876 (n16741, n16735, n16736, n16737, n16740);
  nor g56877 (n9838, n9832, n9833, n9834, n9837);
  nor g56878 (n10423, n10417, n10418, n10419, n10422);
  and g56879 (n_23982, n_255, n_221);
  and g56880 (n_23983, n_75, n_224);
  and g56881 (n_23984, n_93, n1497);
  and g56882 (n5773, n3524, n_23982, n_23983, n_23984);
  and g56883 (n_23985, n_229, n_199);
  and g56884 (n_23986, n_190, n_36);
  and g56885 (n_23987, n_119, n1795, n_74, n_115);
  and g56886 (n_23988, n_226, n720, n2006, n2010);
  and g56887 (n_23989, n1183, n2012, n1600, n2017);
  and g56888 (n_23990, n2020, n2040, n_23985, n_23986);
  and g56889 (n2057, n_23987, n_23988, n_23989, n_23990);
  nor g56890 (n18657, n18651, n18652, n18653, n18656);
  nor g56891 (n18074, n18068, n18069, n18070, n18073);
  nor g56892 (n19176, n19170, n19171, n19172, n19175);
  nor g56893 (n21912, n21906, n21907, n21908, n21911);
  nor g56894 (n18576, n18570, n18571, n18572, n18575);
  nor g56895 (n7583, n7577, n7578, n7579, n7582);
  nor g56896 (n9303, n9297, n9298, n9299, n9302);
  nor g56897 (n8365, n8359, n8360, n8361, n8364);
  nor g56898 (n8800, n8794, n8795, n8796, n8799);
  nor g56899 (n7222, n7216, n7217, n7218, n7221);
  and g56900 (n_23991, n_276, n_204, n_292);
  and g56901 (n_23992, n_66, n_75, n_291);
  and g56902 (n_23993, n1994, n297, n793);
  and g56903 (n_23994, n1898, n1996);
  and g56904 (n2006, n_23991, n_23992, n_23993, n_23994);
  and g56905 (n_23995, n_231, n_185, n_201, n_67);
  and g56906 (n_23996, n_244, n1009, n1668, n1330);
  and g56907 (n_23997, n2021, n2022, n1691, n2025);
  and g56908 (n_23998, n529, n1329, n2026);
  and g56909 (n2040, n_23995, n_23996, n_23997, n_23998);
  and g56910 (n_23999, n_169, n_43, n_214, n_98);
  and g56911 (n_24000, n618, n4786, n1029, n6020);
  and g56912 (n_24001, n2439, n6026, n3580, n2127);
  and g56913 (n_24002, n1084, n5056, n4335, n5152);
  and g56914 (n6041, n_23999, n_24000, n_24001, n_24002);
  and g56915 (n_24003, n_253, n_231);
  and g56916 (n_24004, n_44, n_161);
  and g56917 (n_24005, n_150, n_195);
  and g56918 (n_24006, n_184, n_51);
  and g56919 (n_24007, n_78, n_213, n356, n2088);
  and g56920 (n_24008, n120, n1251, n2104, n2127);
  and g56921 (n_24009, n2132, n2133, n475, n2013);
  and g56922 (n_24010, n_24003, n_24004, n_24005, n_24006);
  and g56923 (n2152, n_24007, n_24008, n_24009, n_24010);
  nor g56924 (n18091, n18085, n18086, n18087, n18090);
  nor g56925 (n19193, n19187, n19188, n19189, n19192);
  nor g56926 (n18558, n18552, n18553, n18554, n18557);
  nor g56927 (n11070, n11064, n11065, n11066, n11069);
  nor g56928 (n7939, n7933, n7934, n7935, n7938);
  and g56929 (n2025, n_162, n_180, n_76, n_159);
  and g56930 (n_24011, n_191, n_44, n_115, n_97);
  and g56931 (n_24012, n_93, n1247, n2417);
  and g56932 (n_24013, n1131, n2422, n2423);
  and g56933 (n_24014, n2424, n2426, n2427);
  and g56934 (n2439, n_24011, n_24012, n_24013, n_24014);
  and g56935 (n_24015, n_117, n_239, n2105, n_74);
  and g56936 (n_24016, n108, n1063, n2021);
  and g56937 (n_24017, n2112, n1012, n1879);
  and g56938 (n_24018, n1643, n2113, n2115);
  and g56939 (n2127, n_24015, n_24016, n_24017, n_24018);
  and g56940 (n_24019, n_217, n_235, n_164);
  and g56941 (n_24020, n_63, n_278, n_79);
  and g56942 (n_24021, n_147, n2089, n2090);
  and g56943 (n_24022, n2091, n2092, n2093);
  and g56944 (n2104, n_24019, n_24020, n_24021, n_24022);
  and g56945 (n_24023, n_98, n_273, n508, n1247);
  and g56946 (n_24024, n2167, n423, n1668, n2169);
  and g56947 (n_24025, n671, n757, n2172);
  and g56948 (n_24026, n2174, n1456, n2176);
  and g56949 (n2189, n_24023, n_24024, n_24025, n_24026);
  nor g56950 (n17589, n17583, n17584, n17585, n17588);
  nor g56951 (n19211, n19205, n19206, n19207, n19210);
  nor g56952 (n19837, n19831, n19832, n19833, n19836);
  nor g56953 (n16759, n16753, n16754, n16755, n16758);
  nor g56954 (n7035, n7029, n7030, n7031, n7034);
  nor g56955 (n8347, n8341, n8342, n8343, n8346);
  and g56956 (n_24027, n_259, n_164);
  and g56957 (n_24028, n_96, n_83);
  and g56958 (n_24029, n_270, n_249);
  and g56959 (n_24030, n1324, n2410);
  and g56960 (n2417, n_24027, n_24028, n_24029, n_24030);
  and g56961 (n_24031, n_54, n_100);
  and g56962 (n_24032, n_140, n_39);
  and g56963 (n_24033, n_241, n_188);
  and g56964 (n_24034, n_89, n_254);
  and g56965 (n2112, n_24031, n_24032, n_24033, n_24034);
  and g56966 (n_24035, n_136, n_85, n_154, n_184);
  and g56967 (n_24036, n_271, n_296, n_68, n341);
  and g56968 (n_24037, n2073, n1128, n1379);
  and g56969 (n_24038, n1890, n1328, n2154);
  and g56970 (n2167, n_24035, n_24036, n_24037, n_24038);
  nor g56971 (n6496, n6488, n6489, n6490, n6493);
  nor g56972 (n19854, n19848, n19849, n19850, n19853);
  and g56973 (n_24039, n_265, n_208, n_177, n_250);
  and g56974 (n_24040, n_46, n1253, n15970, n1131);
  and g56975 (n_24041, n2360, n1549, n459, n4819);
  and g56976 (n_24042, n1693, n1388, n2192);
  and g56977 (n15984, n_24039, n_24040, n_24041, n_24042);
  nor g56978 (n15993, n15985, n15986, n15987, n15990);
  nor g56979 (n7567, n7561, n7562, n7563, n7566);
  nor g56980 (n7921, n7915, n7916, n7917, n7920);
  nor g56981 (n7206, n7200, n7201, n7202, n7205);
  nor g56982 (n20470, n20464, n20465, n20466, n20469);
  nor g56983 (n11097, n11091, n11092, n11093, n11096);
  and g56984 (n_24043, n_158, n_246, n_198, n_133);
  and g56985 (n_24044, n_127, n_248, n_50, n_262);
  and g56986 (n_24045, n827, n2443, n1009, n471);
  and g56987 (n_24046, n15953, n14476, n15956);
  and g56988 (n15970, n_24043, n_24044, n_24045, n_24046);
  and g56989 (n_24047, n_202, n_294, n_181);
  and g56990 (n_24048, n_239, n_149, n2347);
  and g56991 (n_24049, n_289, n241, n2348);
  and g56992 (n_24050, n2349, n1636, n1739);
  and g56993 (n2360, n_24047, n_24048, n_24049, n_24050);
  nor g56994 (n8892, n8886, n8887, n8888, n8891);
  nor g56995 (n9897, n9891, n9892, n9893, n9896);
  and g56996 (n_24051, n_191, n_277);
  and g56997 (n_24052, n_238, n_268);
  and g56998 (n_24053, n_100, n_80);
  and g56999 (n_24054, n1379, n731, n423, n454);
  and g57000 (n_24055, n604, n4274, n2961, n2623);
  and g57001 (n_24056, n6054, n324, n204, n4828);
  and g57002 (n_24057, n6056, n_24051, n_24052, n_24053);
  and g57003 (n6074, n_24054, n_24055, n_24056, n_24057);
  nor g57004 (n17607, n17601, n17602, n17603, n17606);
  nor g57005 (n19872, n19866, n19867, n19868, n19871);
  nor g57006 (n20487, n20481, n20482, n20483, n20486);
  and g57007 (n_24058, n_209, n_60);
  and g57008 (n15953, n_284, n3160, n3391, n_24058);
  nor g57009 (n16777, n16771, n16772, n16773, n16776);
  nor g57010 (n7549, n7543, n7544, n7545, n7548);
  and g57011 (n_24059, n_245, n_106, n_153, n510);
  and g57012 (n_24060, n2202, n2208, n2217, n2258);
  and g57013 (n_24061, n1268, n2262, n2263);
  and g57014 (n_24062, n365, n2275, n2278);
  and g57015 (n2291, n_24059, n_24060, n_24061, n_24062);
  nor g57016 (n17671, n17665, n17666, n17667, n17670);
  and g57017 (n_24063, n_201, n_261, n_227, n_79);
  and g57018 (n_24064, n2073, n1916, n3912, n13135);
  and g57019 (n_24065, n13210, n3205, n5304, n6565);
  and g57020 (n_24066, n595, n2625, n3148);
  and g57021 (n16008, n_24063, n_24064, n_24065, n_24066);
  nor g57022 (n16017, n16009, n16010, n16011, n16014);
  nor g57023 (n8051, n8045, n8046, n8047, n8050);
  and g57024 (n_24067, n_233, n_119);
  and g57025 (n_24068, n_101, n_175);
  and g57026 (n_24069, n_120, n_250, n_273, n_47);
  and g57027 (n_24070, n1389, n116, n2219, n1994);
  and g57028 (n_24071, n2229, n808, n2237, n2240);
  and g57029 (n_24072, n1763, n2241, n_24067, n_24068);
  and g57030 (n2258, n_24069, n_24070, n_24071, n_24072);
  nor g57031 (n18151, n18145, n18146, n18147, n18150);
  nor g57032 (n21225, n21219, n21220, n21221, n21224);
  nor g57033 (n11115, n11109, n11110, n11111, n11114);
  and g57034 (n_24073, n_217, n_124);
  and g57035 (n6565, n_278, n423, n_288, n_24073);
  nor g57036 (n8910, n8904, n8905, n8906, n8909);
  nor g57037 (n9915, n9909, n9910, n9911, n9914);
  and g57038 (n_24074, n_99, n_116, n_82);
  and g57039 (n_24075, n_160, n_271, n_152);
  and g57040 (n_24076, n1069, n2093);
  and g57041 (n_24077, n595, n2220);
  and g57042 (n2229, n_24074, n_24075, n_24076, n_24077);
  nor g57043 (n17625, n17619, n17620, n17621, n17624);
  nor g57044 (n17703, n17697, n17698, n17699, n17702);
  nor g57045 (n17184, n17178, n17179, n17180, n17183);
  nor g57046 (n20505, n20499, n20500, n20501, n20504);
  nor g57047 (n21242, n21236, n21237, n21238, n21241);
  nor g57048 (n21844, n21838, n21839, n21840, n21843);
  and g57049 (n_24078, n_109, n_185);
  and g57050 (n_24079, n_261, n_176);
  and g57051 (n_24080, n_216, n_120);
  and g57052 (n_24081, n_81, n_212, n_148, n418);
  and g57053 (n_24082, n1247, n5085, n15337, n14498);
  and g57054 (n_24083, n16031, n3409, n658, n2992);
  and g57055 (n_24084, n12785, n_24078, n_24079, n_24080);
  and g57056 (n16049, n_24081, n_24082, n_24083, n_24084);
  nor g57057 (n16795, n16789, n16790, n16791, n16794);
  nor g57058 (n16101, n16095, n16096, n16097, n16098);
  nor g57059 (n6129, n6123, n6124, n6125, n6126);
  and g57060 (n_24085, n_277, n_204, n_228, n_73);
  and g57061 (n_24086, n4786, n1291, n333, n6083);
  and g57062 (n_24087, n6097, n2751, n6102, n2807);
  and g57063 (n_24088, n2241, n4269, n6104);
  and g57064 (n6118, n_24085, n_24086, n_24087, n_24088);
  nor g57065 (n17260, n17254, n17255, n17256, n17259);
  nor g57066 (n17201, n17195, n17196, n17197, n17200);
  nor g57067 (n16857, n16851, n16852, n16853, n16856);
  nor g57068 (n18717, n18711, n18712, n18713, n18716);
  nor g57069 (n8069, n8063, n8064, n8065, n8068);
  and g57070 (n_24089, n_185, n_134);
  and g57071 (n_24090, n_124, n_101, n_47, n1478);
  and g57072 (n_24091, n731, n454, n6514, n4375);
  and g57073 (n_24092, n4405, n1709, n6517, n6520);
  and g57074 (n_24093, n691, n3524, n5775, n_24089);
  and g57075 (n6536, n_24090, n_24091, n_24092, n_24093);
  nor g57076 (n6545, n6537, n6538, n6539, n6542);
  nor g57077 (n17762, n17756, n17757, n17758, n17761);
  nor g57078 (n18183, n18177, n18178, n18179, n18182);
  nor g57079 (n21260, n21254, n21255, n21256, n21259);
  nor g57080 (n21830, n21824, n21825, n21826, n21829);
  nor g57081 (n11133, n11127, n11128, n11129, n11132);
  and g57082 (n_24094, n_185, n_58, n_67, n_120);
  and g57083 (n_24095, n_262, n16067, n2346, n2112);
  and g57084 (n_24096, n6662, n2072, n3771, n2172);
  and g57085 (n_24097, n2441, n1409, n1644);
  and g57086 (n16081, n_24094, n_24095, n_24096, n_24097);
  nor g57087 (n8928, n8922, n8923, n8924, n8927);
  nor g57088 (n9933, n9927, n9928, n9929, n9932);
  and g57089 (n_24098, n_92, n_169, n_150, n_37);
  and g57090 (n_24099, n827, n282, n16055);
  and g57091 (n_24100, n15826, n790, n3905);
  and g57092 (n_24101, n13268, n2007, n3128);
  and g57093 (n16067, n_24098, n_24099, n_24100, n_24101);
  and g57094 (n_24102, n_143, n_181, n_172);
  and g57095 (n_24103, n_148, n_147, n_187);
  and g57096 (n_24104, n_48, n1523, n1105);
  and g57097 (n_24105, n3409, n3314, n3549);
  and g57098 (n6662, n_24102, n_24103, n_24104, n_24105);
  nor g57099 (n16813, n16807, n16808, n16809, n16812);
  and g57100 (n_24106, n_92, n_277);
  and g57101 (n_24107, n_151, n_52);
  and g57102 (n_24108, n_264, n1021, n_196, n1252);
  and g57103 (n_24109, n937, n1667, n2317, n2345);
  and g57104 (n_24110, n2360, n2370, n2371, n308);
  and g57105 (n_24111, n793, n1839, n_24106, n_24107);
  and g57106 (n2388, n_24108, n_24109, n_24110, n_24111);
  nor g57107 (n18242, n18236, n18237, n18238, n18241);
  nor g57108 (n19271, n19265, n19266, n19267, n19270);
  nor g57109 (n21813, n21807, n21808, n21809, n21812);
  nor g57110 (n18749, n18743, n18744, n18745, n18748);
  and g57111 (n_24112, n_65, n_192);
  and g57112 (n_24113, n_82, n_95);
  and g57113 (n_24114, n_263, n1160);
  and g57114 (n16055, n2191, n_24112, n_24113, n_24114);
  and g57115 (n_24115, n_72, n_206);
  and g57116 (n_24116, n_58, n_132);
  and g57117 (n_24117, n_78, n_68);
  and g57118 (n_24118, n1761, n450);
  and g57119 (n_24119, n5063, n6561, n4367, n268);
  and g57120 (n_24120, n1709, n877, n6565, n1692);
  and g57121 (n_24121, n6567, n2220, n1740, n3416);
  and g57122 (n_24122, n_24115, n_24116, n_24117, n_24118);
  and g57123 (n6586, n_24119, n_24120, n_24121, n_24122);
  nor g57124 (n6595, n6587, n6588, n6589, n6592);
  nor g57125 (n8087, n8081, n8082, n8083, n8086);
  and g57126 (n_24123, n_276, n_155);
  and g57127 (n_24124, n_206, n_268);
  and g57128 (n_24125, n_81, n_113);
  and g57129 (n_24126, n2361, n2363);
  and g57130 (n2370, n_24123, n_24124, n_24125, n_24126);
  and g57131 (n_24127, n_255, n_219);
  and g57133 (n_24129, n_52, n_195);
  and g57134 (n_24130, n_91, n_273);
  and g57135 (n_24131, n2405, n2068, n399, n1667);
  and g57136 (n_24132, n2406, n604, n665, n2040);
  and g57137 (n_24133, n790, n2409, n2441, n2445);
  and g57138 (n_24134, n_24127, n_22933, n_24129, n_24130);
  and g57139 (n2464, n_24131, n_24132, n_24133, n_24134);
  nor g57140 (n11151, n11145, n11146, n11147, n11150);
  and g57141 (n_24135, n_169, n_228, n_267, n_37);
  and g57142 (n_24136, n_70, n_250, n_254, n100);
  and g57143 (n_24137, n2583, n4127, n1586);
  and g57144 (n_24138, n1785, n5021, n6548);
  and g57145 (n6561, n_24135, n_24136, n_24137, n_24138);
  nor g57146 (n8946, n8940, n8941, n8942, n8945);
  nor g57147 (n9951, n9945, n9946, n9947, n9950);
  and g57148 (n_24139, n_292, n_135, n_72, n_221);
  and g57149 (n_24140, n_267, n_119, n_177, n_40);
  and g57150 (n_24141, n_212, n1108, n_48, n1761);
  and g57151 (n_24142, n1380, n1879, n362, n2390);
  and g57152 (n2405, n_24139, n_24140, n_24141, n_24142);
  nor g57153 (n19303, n19297, n19298, n19299, n19302);
  nor g57154 (n19932, n19926, n19927, n19928, n19931);
  nor g57155 (n18808, n18802, n18803, n18804, n18807);
  and g57156 (n_24143, n_121, n_122);
  and g57157 (n_24144, n_268, n_227);
  and g57158 (n_24145, n_186, n_87);
  and g57159 (n_24146, n_177, n_95, n_70, n2483);
  and g57160 (n_24147, n720, n2484, n2500, n2506);
  and g57161 (n_24148, n2439, n2507, n2512, n351);
  and g57162 (n_24149, n2515, n_24143, n_24144, n_24145);
  and g57163 (n2533, n_24146, n_24147, n_24148, n_24149);
  and g57164 (n_24150, n_185, n_86, n_66, n_270);
  and g57165 (n_24151, n_160, n_156, n6604, n6625);
  and g57166 (n_24152, n5224, n3768, n2370);
  and g57167 (n_24153, n6628, n172, n1497);
  and g57168 (n6641, n_24150, n_24151, n_24152, n_24153);
  nor g57169 (n6650, n6642, n6643, n6644, n6647);
  nor g57170 (n7391, n7385, n7386, n7387, n7390);
  nor g57171 (n8105, n8099, n8100, n8101, n8104);
  nor g57172 (n20565, n20559, n20560, n20561, n20564);
  nor g57173 (n11169, n11163, n11164, n11165, n11168);
  and g57174 (n_24154, n_253, n_53, n_217, n_114);
  and g57175 (n_24155, n_119, n_175, n2466, n193);
  and g57176 (n_24156, n2467, n2348, n2468);
  and g57177 (n_24157, n899, n990, n2470);
  and g57178 (n2483, n_24154, n_24155, n_24156, n_24157);
  and g57179 (n_24158, n_256, n_65);
  and g57180 (n_24159, n_251, n_98);
  and g57181 (n_24160, n_76, n_197);
  and g57182 (n2506, n_239, n_24158, n_24159, n_24160);
  and g57183 (n6628, n_149, n_142, n_226, n2169);
  nor g57184 (n8964, n8958, n8959, n8960, n8963);
  nor g57185 (n9969, n9963, n9964, n9965, n9968);
  nor g57186 (n19964, n19958, n19959, n19960, n19963);
  nor g57187 (n19362, n19356, n19357, n19358, n19361);
  nor g57188 (n12264, n12258, n12259, n12260, n12263);
  and g57189 (n_24161, n_231, n_261, n_37, n_140);
  and g57190 (n_24162, n_263, n_174, n1389, n1379);
  and g57191 (n_24163, n2543, n2555, n1202, n844);
  and g57192 (n_24164, n1879, n989, n638, n2556);
  and g57193 (n2571, n_24161, n_24162, n_24163, n_24164);
  nor g57194 (n7409, n7403, n7404, n7405, n7408);
  nor g57195 (n8123, n8117, n8118, n8119, n8122);
  nor g57196 (n20023, n20017, n20018, n20019, n20022);
  nor g57197 (n21320, n21314, n21315, n21316, n21319);
  nor g57198 (n11187, n11181, n11182, n11183, n11186);
  and g57199 (n_24165, n_34, n_104);
  and g57200 (n_24166, n_86, n_44);
  and g57201 (n_24167, n_282, n624);
  and g57202 (n2543, n2537, n_24165, n_24166, n_24167);
  and g57204 (n_24169, n_230, n_205);
  and g57205 (n_24170, n_125, n_156);
  and g57206 (n_24171, n1161, n978, n1141, n1531);
  and g57207 (n_24172, n2573, n805, n6662, n2258);
  and g57208 (n_24173, n6667, n6670, n4269, n1578);
  and g57209 (n_24174, n6672, n_22716, n_24169, n_24170);
  and g57210 (n6690, n_24171, n_24172, n_24173, n_24174);
  nor g57211 (n6699, n6691, n6692, n6693, n6696);
  nor g57212 (n8982, n8976, n8977, n8978, n8981);
  nor g57213 (n9987, n9981, n9982, n9983, n9986);
  nor g57214 (n12250, n12244, n12245, n12246, n12249);
  nor g57215 (n20597, n20591, n20592, n20593, n20596);
  nor g57216 (n21745, n21739, n21740, n21741, n21744);
  and g57217 (n2537, n_134, n_167, n_101, n_149);
  and g57218 (n_24175, n_253, n_229, n_290, n_194);
  and g57219 (n_24176, n_135, n_138, n6705, n2021);
  and g57220 (n_24177, n6707, n6732, n1454, n2632);
  and g57221 (n_24178, n1615, n1221, n6734);
  and g57222 (n6748, n_24175, n_24176, n_24177, n_24178);
  nor g57223 (n7427, n7421, n7422, n7423, n7426);
  nor g57224 (n6813, n6807, n6808, n6809, n6810);
  nor g57225 (n8141, n8135, n8136, n8137, n8140);
  nor g57226 (n20656, n20650, n20651, n20652, n20655);
  nor g57227 (n21352, n21346, n21347, n21348, n21351);
  and g57228 (n_24179, n_92, n_71);
  and g57229 (n_24180, n_163, n_228);
  and g57230 (n_24181, n_110, n_283);
  and g57231 (n_24182, n_213, n_200, n_287, n720);
  and g57232 (n_24183, n979, n159, n2573, n2581);
  and g57233 (n_24184, n2623, n2632, n2650, n2653);
  and g57234 (n_24185, n2656, n_24179, n_24180, n_24181);
  and g57235 (n2674, n_24182, n_24183, n_24184, n_24185);
  and g57236 (n_24186, n_117, n_150);
  and g57237 (n_24187, n_74, n_289);
  and g57238 (n6705, n300, n_126, n_24186, n_24187);
  and g57239 (n_24188, n_219, n_202, n_280, n_67);
  and g57240 (n_24189, n_291, n_213, n227, n826);
  and g57241 (n_24190, n1531, n6714, n665, n1476);
  and g57242 (n_24191, n897, n6716, n2423, n6717);
  and g57243 (n6732, n_24188, n_24189, n_24190, n_24191);
  and g57244 (n_24192, n_274, n_154);
  and g57245 (n_24193, n_97, n2371);
  and g57246 (n2632, n2625, n2627, n_24192, n_24193);
  nor g57247 (n9000, n8994, n8995, n8996, n8999);
  nor g57248 (n10005, n9999, n10000, n10001, n10004);
  and g57249 (n_24194, n_253, n_229, n_94, n_36);
  and g57250 (n_24195, n_174, n2484, n933, n2633);
  and g57251 (n_24196, n811, n1419, n1738);
  and g57252 (n_24197, n2637, n1578, n1828);
  and g57253 (n2650, n_24194, n_24195, n_24196, n_24197);
  and g57254 (n2656, n_206, n_58, n_179, n_241);
  and g57255 (n_24198, n_247, n_162);
  and g57256 (n_24199, n_164, n_264);
  and g57257 (n_24200, n3886, n2633);
  and g57258 (n_24201, n1528, n1617);
  and g57259 (n6714, n_24198, n_24199, n_24200, n_24201);
  and g57260 (n_24202, n_100, n_267);
  and g57261 (n_24203, n_160, n_74);
  and g57262 (n_24204, n_212, n_105);
  and g57263 (n_24205, n_118, n_93);
  and g57264 (n_24206, n810, n2466);
  and g57265 (n_24207, n869, n288, n1668, n510);
  and g57266 (n_24208, n6755, n6769, n2104, n4148);
  and g57267 (n_24209, n6771, n735, n1586, n_24202);
  and g57268 (n_24210, n_24203, n_24204, n_24205, n_24206);
  and g57269 (n6791, n_24207, n_24208, n_24209, n_24210);
  nor g57270 (n6802, n6792, n6793, n6794, n6799);
  nor g57271 (n21714, n21708, n21709, n21710, n21713);
  nor g57272 (n21411, n21405, n21406, n21407, n21410);
  and g57273 (n_24211, n_163, n_138);
  and g57274 (n_24212, n_227, n_165);
  and g57275 (n_24213, n_297, n_38);
  and g57276 (n_24214, n300, n2704);
  and g57277 (n6755, n_24211, n_24212, n_24213, n_24214);
  and g57278 (n_24215, n_285, n_72, n_249, n_244);
  and g57279 (n_24216, n937, n2678, n2697, n1183);
  and g57280 (n_24217, n2698, n2703, n2716, n2650);
  and g57281 (n_24218, n2719, n2230, n2303, n2721);
  and g57282 (n2736, n_24215, n_24216, n_24217, n_24218);
  nor g57283 (n7445, n7439, n7440, n7441, n7444);
  nor g57284 (n8159, n8153, n8154, n8155, n8158);
  and g57285 (n_24219, n_34, n_279, n_290, n_175);
  and g57286 (n_24220, n_59, n2583, n979, n1182);
  and g57287 (n_24221, n2325, n2682, n1387);
  and g57288 (n_24222, n2133, n2390, n2684);
  and g57289 (n2697, n_24219, n_24220, n_24221, n_24222);
  and g57290 (n2719, n_102, n_129, n_193, n1782);
  nor g57291 (n10558, n10552, n10553, n10554, n10557);
  nor g57292 (n_24223, n21658, n21659);
  nor g57293 (n_24224, n21665, n21666);
  nor g57294 (n_24225, n21667, n21668);
  and g57295 (n21674, \a[2] , n_24223, n_24224, n_24225);
  and g57296 (n_24226, n_133, n_138);
  and g57297 (n_24227, n_82, n_115);
  and g57298 (n_24228, n2276, n421);
  and g57299 (n_24229, n533, n1917, n1577, n789);
  and g57300 (n_24230, n2772, n2796, n2806, n1709);
  and g57301 (n_24231, n2807, n2808, n2809, n1828);
  and g57302 (n_24232, n2811, n_24226, n_24227, n_24228);
  and g57303 (n2829, n_24229, n_24230, n_24231, n_24232);
  nor g57304 (n10575, n10569, n10570, n10571, n10574);
  nor g57305 (n11233, n11227, n11228, n11229, n11232);
  nor g57306 (n7463, n7457, n7458, n7459, n7462);
  nor g57307 (n11250, n11244, n11245, n11246, n11249);
  nor g57308 (n12182, n12176, n12177, n12178, n12181);
  nor g57309 (n21683, n21677, n21678, n21679, n21682);
  nor g57310 (n8551, n8545, n8546, n8547, n8550);
  nor g57311 (n9474, n9468, n9469, n9470, n9473);
  nor g57312 (n11268, n11262, n11263, n11264, n11267);
  nor g57313 (n12168, n12162, n12163, n12164, n12167);
  nor g57314 (n7512, n7506, n7507, n7508, n7511);
  nor g57315 (n8568, n8562, n8563, n8564, n8567);
  nor g57316 (n9491, n9485, n9486, n9487, n9490);
  nor g57317 (n7786, n7780, n7781, n7782, n7785);
  nor g57318 (n12151, n12145, n12146, n12147, n12150);
  nor g57319 (n9046, n9040, n9041, n9042, n9045);
  nor g57320 (n10051, n10045, n10046, n10047, n10050);
  nor g57321 (n7803, n7797, n7798, n7799, n7802);
  nor g57322 (n8205, n8199, n8200, n8201, n8204);
  nor g57323 (n10068, n10062, n10063, n10064, n10067);
  nor g57324 (n9063, n9057, n9058, n9059, n9062);
  nor g57325 (n10635, n10629, n10630, n10631, n10634);
  nor g57326 (n10086, n10080, n10081, n10082, n10085);
  nor g57327 (n10652, n10646, n10647, n10648, n10651);
  nor g57328 (n9081, n9075, n9076, n9077, n9080);
  nor g57329 (n7862, n7856, n7857, n7858, n7861);
  nor g57330 (n11328, n11322, n11323, n11324, n11327);
  nor g57331 (n10670, n10664, n10665, n10666, n10669);
  nor g57332 (n11345, n11339, n11340, n11341, n11344);
  nor g57333 (n12083, n12077, n12078, n12079, n12082);
  nor g57334 (n8237, n8231, n8232, n8233, n8236);
  nor g57335 (n11363, n11357, n11358, n11359, n11362);
  nor g57336 (n12069, n12063, n12064, n12065, n12068);
  nor g57337 (n9551, n9545, n9546, n9547, n9550);
  nor g57338 (n12052, n12046, n12047, n12048, n12051);
  nor g57339 (n8628, n8622, n8623, n8624, n8627);
  nor g57340 (n9568, n9562, n9563, n9564, n9567);
  nor g57341 (n9586, n9580, n9581, n9582, n9585);
  nor g57342 (n10146, n10140, n10141, n10142, n10145);
  nor g57343 (n8296, n8290, n8291, n8292, n8295);
  nor g57344 (n10163, n10157, n10158, n10159, n10162);
  nor g57345 (n10730, n10724, n10725, n10726, n10729);
  nor g57346 (n10181, n10175, n10176, n10177, n10180);
  nor g57347 (n10747, n10741, n10742, n10743, n10746);
  nor g57348 (n8660, n8654, n8655, n8656, n8659);
  nor g57349 (n11423, n11417, n11418, n11419, n11422);
  nor g57350 (n10765, n10759, n10760, n10761, n10764);
  nor g57351 (n11440, n11434, n11435, n11436, n11439);
  nor g57352 (n11984, n11978, n11979, n11980, n11983);
  nor g57353 (n9141, n9135, n9136, n9137, n9140);
  nor g57354 (n11458, n11452, n11453, n11454, n11457);
  nor g57355 (n11970, n11964, n11965, n11966, n11969);
  nor g57356 (n8719, n8713, n8714, n8715, n8718);
  nor g57357 (n9646, n9640, n9641, n9642, n9645);
  nor g57358 (n11953, n11947, n11948, n11949, n11952);
  nor g57359 (n9173, n9167, n9168, n9169, n9172);
  nor g57360 (n9678, n9672, n9673, n9674, n9677);
  nor g57361 (n10241, n10235, n10236, n10237, n10240);
  nor g57362 (n9232, n9226, n9227, n9228, n9231);
  nor g57363 (n10825, n10819, n10820, n10821, n10824);
  nor g57364 (n10273, n10267, n10268, n10269, n10272);
  nor g57365 (n9737, n9731, n9732, n9733, n9736);
  nor g57366 (n10332, n10326, n10327, n10328, n10331);
  nor g57367 (n11518, n11512, n11513, n11514, n11517);
  nor g57368 (n10857, n10851, n10852, n10853, n10856);
  nor g57369 (n11885, n11879, n11880, n11881, n11884);
  nor g57370 (n10916, n10910, n10911, n10912, n10915);
  nor g57371 (n11550, n11544, n11545, n11546, n11549);
  nor g57372 (n11854, n11848, n11849, n11850, n11853);
  nor g57373 (n11609, n11603, n11604, n11605, n11608);
  nor g57374 (n_24233, n11795, n11797);
  nor g57375 (n_24234, n11803, n11804);
  nor g57376 (n_24235, n11806, n11808);
  and g57377 (n11814, \a[2] , n_24233, n_24234, n_24235);
  nor g57378 (n11823, n11817, n11818, n11819, n11822);
  nor g57379 (n26930, n26924, n26925, n26926, n26929);
  nor g57380 (n27160, n27154, n27155, n27156, n27157);
  nor g57381 (n26942, n26936, n26937, n26938, n26941);
  nor g57382 (n26954, n26948, n26949, n26950, n26953);
  nor g57383 (n26966, n26960, n26961, n26962, n26965);
  and g57384 (n_24236, n_266, n_280);
  and g57385 (n_24237, n_164, n_123);
  and g57386 (n_24238, n_146, n_296);
  and g57387 (n_24239, n1522, n2405, n1237, n2583);
  and g57388 (n_24240, n1575, n3544, n2979, n6755);
  and g57389 (n_24241, n14544, n6628, n2025, n1603);
  and g57390 (n_24242, n3514, n_24236, n_24237, n_24238);
  and g57391 (n26991, n_24239, n_24240, n_24241, n_24242);
  nor g57392 (n26998, n26992, n26993, n26994, n26995);
  nor g57393 (n27207, n27201, n27202, n27203, n27206);
  nor g57394 (n27417, n27411, n27412, n27413, n27414);
  nor g57395 (n27219, n27213, n27214, n27215, n27218);
  nor g57396 (n27231, n27225, n27226, n27227, n27230);
  nor g57397 (n27243, n27237, n27238, n27239, n27242);
  and g57398 (n_24243, n_199, n_99);
  and g57399 (n_24244, n_116, n_205);
  and g57400 (n_24245, n_37, n1269, n1726, n515);
  and g57401 (n_24246, n1844, n1479, n1600, n3191);
  and g57402 (n_24247, n3180, n616, n2410, n6717);
  and g57403 (n_24248, n13827, n14561, n_24243, n_24244);
  and g57404 (n27267, n_24245, n_24246, n_24247, n_24248);
  nor g57405 (n27274, n27268, n27269, n27270, n27271);
  nor g57406 (n27477, n27471, n27472, n27473, n27476);
  nor g57407 (n27682, n27676, n27677, n27678, n27679);
  nor g57408 (n27489, n27483, n27484, n27485, n27488);
  nor g57409 (n27501, n27495, n27496, n27497, n27500);
  nor g57410 (n27513, n27507, n27508, n27509, n27512);
  and g57411 (n_24249, n_143, n_66, n1182, n1826);
  and g57412 (n_24250, n510, n2229, n6769, n6732);
  and g57413 (n_24251, n15743, n4769, n2410);
  and g57414 (n_24252, n27522, n1721, n1737);
  and g57415 (n27535, n_24249, n_24250, n_24251, n_24252);
  nor g57416 (n27542, n27536, n27537, n27538, n27539);
  nor g57417 (n27735, n27729, n27730, n27731, n27734);
  nor g57418 (n27747, n27741, n27742, n27743, n27746);
  nor g57419 (n27759, n27753, n27754, n27755, n27758);
  nor g57420 (n27771, n27765, n27766, n27767, n27770);
  and g57421 (n_24253, n_182, n_99);
  and g57422 (n_24254, n_37, n_241);
  and g57423 (n_24255, n_146, n570);
  and g57424 (n_24256, n978, n120, n27789, n2012);
  and g57425 (n_24257, n4388, n3127, n1709, n3040);
  and g57426 (n_24258, n526, n1240, n1681, n1140);
  and g57427 (n_24259, n2092, n_24253, n_24254, n_24255);
  and g57428 (n27807, n_24256, n_24257, n_24258, n_24259);
  nor g57429 (n27814, n27808, n27809, n27810, n27811);
  and g57430 (n_24260, n_277, n_268, n_62);
  and g57431 (n_24261, n_205, n_76, n_87);
  and g57432 (n_24262, n_171, n_38, n1575);
  and g57433 (n_24263, n3544, n1423, n2093);
  and g57434 (n27789, n_24260, n_24261, n_24262, n_24263);
  nor g57435 (n27998, n27992, n27993, n27994, n27997);
  nor g57436 (n28010, n28004, n28005, n28006, n28009);
  nor g57437 (n28022, n28016, n28017, n28018, n28021);
  nor g57438 (n28034, n28028, n28029, n28030, n28033);
  and g57439 (n_24264, n_109, n_53);
  and g57440 (n_24265, n_103, n_65);
  and g57441 (n_24266, n_206, n_166);
  and g57442 (n_24267, n_242, n_55, n_97, n_38);
  and g57443 (n_24268, n_200, n1046, n5286, n3644);
  and g57444 (n_24269, n15970, n12409, n690, n207);
  and g57445 (n_24270, n3587, n_24264, n_24265, n_24266);
  and g57446 (n28059, n_24267, n_24268, n_24269, n_24270);
  nor g57447 (n28066, n28060, n28061, n28062, n28063);
  nor g57448 (n28244, n28238, n28239, n28240, n28243);
  nor g57449 (n28256, n28250, n28251, n28252, n28255);
  nor g57450 (n28268, n28262, n28263, n28264, n28267);
  nor g57451 (n28280, n28274, n28275, n28276, n28279);
  and g57452 (n_24271, n_183, n_277);
  and g57453 (n_24272, n_34, n_274);
  and g57454 (n_24273, n_251, n_164);
  and g57455 (n_24274, n_100, n_252);
  and g57456 (n_24275, n116, n2405);
  and g57457 (n_24276, n227, n978, n507, n15047);
  and g57458 (n_24277, n5013, n14565, n28294, n3040);
  and g57459 (n_24278, n437, n297, n27522, n_24271);
  and g57460 (n_24279, n_24272, n_24273, n_24274, n_24275);
  and g57461 (n28314, n_24276, n_24277, n_24278, n_24279);
  nor g57462 (n28321, n28315, n28316, n28317, n28318);
  and g57464 (n_24281, n_233, n_66);
  and g57465 (n_24282, n_88, n_59);
  and g57466 (n_24283, n1550, n1693);
  and g57467 (n28294, n_23857, n_24281, n_24282, n_24283);
  nor g57468 (n28665, n28659, n28660, n28661, n28664);
  nor g57469 (n28646, n28640, n28641, n28642, n28645);
  nor g57470 (n28627, n28621, n28622, n28623, n28626);
  nor g57471 (n28608, n28602, n28603, n28604, n28607);
  nor g57472 (n28589, n28583, n28584, n28585, n28588);
  nor g57473 (n28570, n28564, n28565, n28566, n28569);
  nor g57474 (n28551, n28545, n28546, n28547, n28550);
  nor g57475 (n28532, n28526, n28527, n28528, n28531);
  nor g57476 (n28474, n28468, n28469, n28470, n28471);
  and g57477 (n_24284, n_220, n_52);
  and g57478 (n_24285, n_221, n_242);
  and g57479 (n_24286, n_244, n_272);
  and g57480 (n_24287, n1389, n2483, n3984, n1574);
  and g57481 (n_24288, n1884, n3757, n1577, n12944);
  and g57482 (n_24289, n2022, n13698, n6734, n2115);
  and g57483 (n_24290, n2423, n_24284, n_24285, n_24286);
  and g57484 (n28492, n_24287, n_24288, n_24289, n_24290);
  nor g57485 (n28884, n28878, n28879, n28880, n28883);
  nor g57486 (n28865, n28859, n28860, n28861, n28864);
  nor g57487 (n28846, n28840, n28841, n28842, n28845);
  nor g57488 (n28827, n28821, n28822, n28823, n28826);
  nor g57489 (n28808, n28802, n28803, n28804, n28807);
  nor g57490 (n28789, n28783, n28784, n28785, n28788);
  nor g57491 (n28770, n28764, n28765, n28766, n28769);
  nor g57492 (n28751, n28745, n28746, n28747, n28750);
  nor g57493 (n28736, n28730, n28731, n28732, n28735);
  nor g57494 (n28721, n28715, n28716, n28717, n28718);
  and g57495 (n_24291, n_158, n_255);
  and g57496 (n_24292, n_114, n_49);
  and g57497 (n_24293, n279, n3163);
  and g57498 (n_24294, n2088, n2583, n399, n979);
  and g57499 (n_24295, n869, n1782, n1313, n16067);
  and g57500 (n_24296, n28688, n2410, n1424, n1347);
  and g57501 (n_24297, n23251, n_24291, n_24292, n_24293);
  and g57502 (n28706, n_24294, n_24295, n_24296, n_24297);
  and g57503 (n_24298, n_277, n_232);
  and g57504 (n28688, n_126, n720, n16020, n_24298);
  nor g57505 (n29078, n29072, n29073, n29074, n29077);
  nor g57506 (n29059, n29053, n29054, n29055, n29058);
  nor g57507 (n29040, n29034, n29035, n29036, n29039);
  nor g57508 (n29021, n29015, n29016, n29017, n29020);
  nor g57509 (n29002, n28996, n28997, n28998, n29001);
  nor g57510 (n28983, n28977, n28978, n28979, n28982);
  nor g57511 (n28964, n28958, n28959, n28960, n28963);
  nor g57512 (n28949, n28943, n28944, n28945, n28948);
  nor g57513 (n28934, n28928, n28929, n28930, n28931);
  and g57514 (n_24299, n_122, n_79);
  and g57515 (n_24300, n_106, n_284, n_131, n2167);
  and g57516 (n_24301, n937, n2443, n1182, n415);
  and g57517 (n_24302, n770, n5199, n3685, n1103);
  and g57518 (n_24303, n2704, n2424, n15286, n_24299);
  and g57519 (n28919, n_24300, n_24301, n_24302, n_24303);
  nor g57520 (n29297, n29291, n29292, n29293, n29296);
  nor g57521 (n29277, n29271, n29272, n29273, n29276);
  nor g57522 (n29259, n29253, n29254, n29255, n29258);
  nor g57523 (n29239, n29233, n29234, n29235, n29238);
  nor g57524 (n29220, n29214, n29215, n29216, n29219);
  nor g57525 (n29201, n29195, n29196, n29197, n29200);
  nor g57526 (n29182, n29176, n29177, n29178, n29181);
  nor g57527 (n29154, n29148, n29149, n29150, n29151);
  nor g57528 (n29167, n29161, n29162, n29163, n29166);
  and g57529 (n_24304, n_155, n_41, n_112, n_262);
  and g57530 (n_24305, n22748, n1761, n3886, n2467);
  and g57531 (n_24306, n3057, n13826, n526, n960);
  and g57532 (n_24307, n4357, n1073, n1859, n4335);
  and g57533 (n29132, n_24304, n_24305, n_24306, n_24307);
  nor g57534 (n29508, n29502, n29503, n29504, n29507);
  nor g57535 (n29489, n29483, n29484, n29485, n29488);
  nor g57536 (n29469, n29463, n29464, n29465, n29468);
  nor g57537 (n29450, n29444, n29445, n29446, n29449);
  nor g57538 (n29431, n29425, n29426, n29427, n29430);
  nor g57539 (n29412, n29406, n29407, n29408, n29411);
  nor g57540 (n29393, n29387, n29388, n29389, n29392);
  nor g57541 (n29325, n29319, n29320, n29321, n29322);
  and g57542 (n_24308, n_253, n_206);
  and g57543 (n_24309, n_62, n_154);
  and g57544 (n_24310, n_132, n_296);
  and g57545 (n_24311, n_284, n1522, n1825, n1009);
  and g57546 (n_24312, n488, n600, n2678, n1378);
  and g57547 (n_24313, n29337, n6771, n3160, n1732);
  and g57548 (n_24314, n2263, n_24308, n_24309, n_24310);
  and g57549 (n29355, n_24311, n_24312, n_24313, n_24314);
  and g57550 (n_24315, n_76, n_101, n_49, n_89);
  and g57551 (n_24316, n1141, n869, n3470);
  and g57552 (n_24317, n654, n6705, n1346);
  and g57553 (n_24318, n1206, n1324, n6056);
  and g57554 (n29337, n_24315, n_24316, n_24317, n_24318);
  nor g57555 (n29704, n29698, n29699, n29700, n29703);
  nor g57556 (n29685, n29679, n29680, n29681, n29684);
  nor g57557 (n29666, n29660, n29661, n29662, n29665);
  nor g57558 (n29647, n29641, n29642, n29643, n29646);
  nor g57559 (n29628, n29622, n29623, n29624, n29627);
  nor g57560 (n29609, n29603, n29604, n29605, n29608);
  nor g57561 (n29594, n29588, n29589, n29590, n29593);
  nor g57562 (n29579, n29573, n29574, n29575, n29576);
  and g57563 (n_24319, n_151, n_139, n_221, n_198);
  and g57564 (n_24320, n_98, n_184, n_105, n_68);
  and g57565 (n_24321, n12396, n3065, n29538, n29550);
  and g57566 (n_24322, n6548, n12911, n13808);
  and g57567 (n29564, n_24319, n_24320, n_24321, n_24322);
  and g57568 (n_24323, n_137, n_256, n_238);
  and g57569 (n_24324, n_62, n_209);
  and g57570 (n_24325, n_128, n_125);
  and g57571 (n_24326, n_56, n_106);
  and g57572 (n29538, n_24323, n_24324, n_24325, n_24326);
  and g57573 (n_24327, n_99, n_66, n_63, n_51);
  and g57574 (n_24328, n_118, n885, n2417);
  and g57575 (n_24329, n1046, n2406, n4295);
  and g57576 (n_24330, n940, n2442, n12712);
  and g57577 (n29550, n_24327, n_24328, n_24329, n_24330);
  nor g57578 (n29902, n29896, n29897, n29898, n29901);
  nor g57579 (n29882, n29876, n29877, n29878, n29881);
  nor g57580 (n29864, n29858, n29859, n29860, n29863);
  nor g57581 (n29844, n29838, n29839, n29840, n29843);
  nor g57582 (n29825, n29819, n29820, n29821, n29824);
  nor g57583 (n29806, n29800, n29801, n29802, n29805);
  nor g57584 (n29749, n29743, n29744, n29745, n29746);
  nor g57585 (n29787, n29781, n29782, n29783, n29786);
  and g57586 (n_24331, n_161, n_273, n156, n2170);
  and g57587 (n_24332, n2484, n2958, n235, n2697);
  and g57588 (n_24333, n1575, n2006, n13773, n300);
  and g57589 (n_24334, n1422, n960, n3474);
  and g57590 (n29767, n_24331, n_24332, n_24333, n_24334);
  nor g57591 (n30077, n30071, n30072, n30073, n30076);
  nor g57592 (n30058, n30052, n30053, n30054, n30057);
  nor g57593 (n30038, n30032, n30033, n30034, n30037);
  nor g57594 (n30019, n30013, n30014, n30015, n30018);
  nor g57595 (n30000, n29994, n29995, n29996, n29999);
  nor g57596 (n29981, n29975, n29976, n29977, n29980);
  nor g57597 (n29930, n29924, n29925, n29926, n29927);
  and g57598 (n_24335, n_137, n_285, n_283, n_116);
  and g57599 (n_24336, n_154, n_79, n_97, n2635);
  and g57600 (n_24337, n3559, n1719, n4786, n4767);
  and g57601 (n_24338, n14407, n15854, n962, n1490);
  and g57602 (n29946, n_24335, n_24336, n_24337, n_24338);
  nor g57603 (n30236, n30230, n30231, n30232, n30235);
  nor g57604 (n30217, n30211, n30212, n30213, n30216);
  nor g57605 (n30198, n30192, n30193, n30194, n30197);
  nor g57606 (n30179, n30173, n30174, n30175, n30178);
  nor g57607 (n30160, n30154, n30155, n30156, n30159);
  nor g57608 (n30132, n30126, n30127, n30128, n30129);
  and g57609 (n_24339, n_220, n_180);
  and g57610 (n_24340, n_36, n_120);
  and g57611 (n_24341, n_188, n1247);
  and g57612 (n_24342, n731, n29337, n1330, n291);
  and g57613 (n_24343, n2651, n5286, n15312, n13768);
  and g57614 (n_24344, n877, n1012, n2007, n2705);
  and g57615 (n_24345, n2811, n_24339, n_24340, n_24341);
  and g57616 (n30117, n_24342, n_24343, n_24344, n_24345);
  nor g57617 (n30420, n30414, n30415, n30416, n30419);
  nor g57618 (n30400, n30394, n30395, n30396, n30399);
  nor g57619 (n30382, n30376, n30377, n30378, n30381);
  nor g57620 (n30362, n30356, n30357, n30358, n30361);
  nor g57621 (n30343, n30337, n30338, n30339, n30342);
  nor g57622 (n30328, n30322, n30323, n30324, n30327);
  nor g57623 (n30283, n30277, n30278, n30279, n30280);
  and g57624 (n_24346, n_158, n_219);
  and g57625 (n_24347, n_184, n_97, n590, n3886);
  and g57626 (n_24348, n1252, n1576, n1435, n241);
  and g57627 (n_24349, n3510, n1407, n5019, n2808);
  and g57628 (n_24350, n5038, n675, n2174, n_24346);
  and g57629 (n30303, n_24347, n_24348, n_24349, n_24350);
  nor g57630 (n30576, n30570, n30571, n30572, n30575);
  nor g57631 (n30557, n30551, n30552, n30553, n30556);
  nor g57632 (n30537, n30531, n30532, n30533, n30536);
  nor g57633 (n30518, n30512, n30513, n30514, n30517);
  nor g57634 (n30499, n30493, n30494, n30495, n30498);
  nor g57635 (n30448, n30442, n30443, n30444, n30445);
  and g57636 (n_24351, n_199, n_175, n_289, n_262);
  and g57637 (n_24352, n_200, n810, n1380, n28294);
  and g57638 (n_24353, n15324, n13458, n27789, n12977);
  and g57639 (n_24354, n3128, n778, n1499, n2059);
  and g57640 (n30464, n_24351, n_24352, n_24353, n_24354);
  nor g57641 (n30716, n30710, n30711, n30712, n30715);
  nor g57642 (n30697, n30691, n30692, n30693, n30696);
  nor g57643 (n30678, n30672, n30673, n30674, n30677);
  nor g57644 (n30659, n30653, n30654, n30655, n30658);
  nor g57645 (n30644, n30638, n30639, n30640, n30643);
  nor g57646 (n30604, n30598, n30599, n30600, n30601);
  and g57647 (n_24355, n_169, n_185);
  and g57648 (n_24356, n_75, n_154);
  and g57649 (n_24357, n_101, n_51, n_289, n_226);
  and g57650 (n_24358, n2739, n5209, n2500, n3386);
  and g57651 (n_24359, n13123, n12710, n3108, n6084);
  and g57652 (n_24360, n694, n2176, n_24355, n_24356);
  and g57653 (n30621, n_24357, n_24358, n_24359, n_24360);
  nor g57654 (n30874, n30868, n30869, n30870, n30873);
  nor g57655 (n30854, n30848, n30849, n30850, n30853);
  nor g57656 (n30836, n30830, n30831, n30832, n30835);
  nor g57657 (n30816, n30810, n30811, n30812, n30815);
  nor g57658 (n30761, n30755, n30756, n30757, n30758);
  nor g57659 (n30797, n30791, n30792, n30793, n30796);
  and g57660 (n_24361, n_192, n_150, n_154, n2219);
  and g57661 (n_24362, n1139, n976, n1291);
  and g57662 (n_24363, n6714, n14202, n1894);
  and g57663 (n_24364, n14482, n2537, n3045);
  and g57664 (n30777, n_24361, n_24362, n_24363, n_24364);
  nor g57665 (n31012, n31006, n31007, n31008, n31011);
  nor g57666 (n30993, n30987, n30988, n30989, n30992);
  nor g57667 (n30973, n30967, n30968, n30969, n30972);
  nor g57668 (n30954, n30948, n30949, n30950, n30953);
  nor g57669 (n30902, n30896, n30897, n30898, n30899);
  and g57670 (n_24365, n_155, n_65);
  and g57671 (n_24366, n_82, n_107, n1782, n471);
  and g57672 (n_24367, n2697, n2346, n1183, n491);
  and g57673 (n_24368, n977, n5773, n5034, n14525);
  and g57674 (n_24369, n2361, n1369, n3393, n_24365);
  and g57675 (n30919, n_24366, n_24367, n_24368, n_24369);
  nor g57676 (n31133, n31127, n31128, n31129, n31132);
  nor g57677 (n31114, n31108, n31109, n31110, n31113);
  nor g57678 (n31095, n31089, n31090, n31091, n31094);
  nor g57679 (n31067, n31061, n31062, n31063, n31064);
  and g57680 (n_24370, n_204, n_217);
  and g57681 (n_24371, n_86, n_96, n_120, n_297);
  and g57682 (n_24372, n1380, n3739, n1781, n2506);
  and g57683 (n_24373, n1100, n13247, n5188, n2263);
  and g57684 (n_24374, n31036, n376, n2026, n_24370);
  and g57685 (n31052, n_24371, n_24372, n_24373, n_24374);
  nor g57686 (n31275, n31269, n31270, n31271, n31274);
  nor g57687 (n31257, n31251, n31252, n31253, n31256);
  nor g57688 (n31239, n31233, n31234, n31235, n31238);
  nor g57689 (n31181, n31175, n31176, n31177, n31180);
  nor g57690 (n31197, n31191, n31192, n31193, n31194);
  and g57691 (n_24375, n_266, n_217, n_125, n_141);
  and g57692 (n_24376, n_89, n279, n448, n882);
  and g57693 (n_24377, n12924, n3282, n4785);
  and g57694 (n_24378, n2719, n1143, n24041);
  and g57695 (n31214, n_24375, n_24376, n_24377, n_24378);
  nor g57696 (n31394, n31388, n31389, n31390, n31393);
  nor g57697 (n31375, n31369, n31370, n31371, n31374);
  nor g57698 (n31354, n31348, n31349, n31350, n31353);
  nor g57699 (n31303, n31297, n31298, n31299, n31300);
  and g57700 (n_24379, n_222, n_244, n_74, n_112);
  and g57701 (n_24380, n_147, n_146, n4101, n418);
  and g57702 (n_24381, n423, n29550, n3497, n2543);
  and g57703 (n_24382, n6514, n2656, n632, n13014);
  and g57704 (n31319, n_24379, n_24380, n_24381, n_24382);
  nor g57705 (n31492, n31486, n31487, n31488, n31491);
  nor g57706 (n31473, n31467, n31468, n31469, n31472);
  nor g57707 (n31458, n31452, n31453, n31454, n31457);
  nor g57708 (n31422, n31416, n31417, n31418, n31419);
  and g57709 (n_24383, n_42, n_85, n_291, n_241);
  and g57710 (n_24384, n28688, n488, n230, n2683);
  and g57711 (n_24385, n2651, n3259, n6561);
  and g57712 (n_24386, n4366, n12941, n31036);
  and g57713 (n31435, n_24383, n_24384, n_24385, n_24386);
  nor g57714 (n31617, n31611, n31612, n31613, n31616);
  nor g57715 (n31597, n31591, n31592, n31593, n31596);
  nor g57716 (n31582, n31576, n31577, n31578, n31581);
  nor g57717 (n31537, n31531, n31532, n31533, n31534);
  and g57718 (n_24387, n_73, n_192);
  and g57719 (n_24388, n_261, n_70);
  and g57720 (n_24389, n_179, n_226, n1574, n615);
  and g57721 (n_24390, n2506, n539, n805, n1008);
  and g57722 (n_24391, n4293, n15953, n15050, n530);
  and g57723 (n_24392, n2753, n3370, n_24387, n_24388);
  and g57724 (n31558, n_24389, n_24390, n_24391, n_24392);
  nor g57725 (n31715, n31709, n31710, n31711, n31714);
  nor g57726 (n31696, n31690, n31691, n31692, n31695);
  nor g57727 (n31645, n31639, n31640, n31641, n31642);
  and g57728 (n_24393, n_109, n_124, n_83, n_241);
  and g57729 (n_24394, n_296, n1252, n16055, n3039);
  and g57730 (n_24395, n1679, n3282, n1029, n14534);
  and g57731 (n_24396, n1640, n1604, n1740, n4828);
  and g57732 (n31661, n_24393, n_24394, n_24395, n_24396);
  nor g57733 (n31796, n31790, n31791, n31792, n31795);
  nor g57734 (n31781, n31775, n31776, n31777, n31780);
  nor g57735 (n31766, n31760, n31761, n31762, n31763);
  and g57736 (n_24397, n_265, n_127, n_91, n_140);
  and g57737 (n_24398, n22762, n720, n1252, n285);
  and g57738 (n_24399, n29538, n2651, n4232, n25863);
  and g57739 (n_24400, n15882, n1070, n3459, n13016);
  and g57740 (n31751, n_24397, n_24398, n_24399, n_24400);
  nor g57741 (n31900, n31894, n31895, n31896, n31899);
  nor g57742 (n31843, n31837, n31838, n31839, n31842);
  nor g57743 (n31858, n31852, n31853, n31854, n31855);
  and g57744 (n_24401, n_214, n_230, n_270, n_88);
  and g57745 (n_24402, n_284, n_211, n193, n1478);
  and g57746 (n_24403, n937, n288, n3866, n4003);
  and g57747 (n_24404, n1155, n4799, n13161);
  and g57748 (n31876, n_24401, n_24402, n_24403, n_24404);
  nor g57749 (n31980, n31974, n31975, n31976, n31979);
  nor g57750 (n31928, n31922, n31923, n31924, n31925);
  and g57751 (n_24405, n_103, n_124);
  and g57752 (n_24406, n_198, n_179, n100, n1783);
  and g57753 (n_24407, n1366, n1531, n1183, n3997);
  and g57754 (n_24408, n3939, n15880, n26016, n6610);
  and g57755 (n_24409, n3438, n1738, n15012, n_24405);
  and g57756 (n31945, n_24406, n_24407, n_24408, n_24409);
  nor g57757 (n32027, n32021, n32022, n32023, n32024);
  nor g57758 (n32051, n32045, n32046, n32047, n32050);
  and g57759 (n_24410, n_270, n3984);
  and g57760 (n_24411, n26016, n2273);
  and g57761 (n_24412, n3839, n3848);
  and g57762 (n_24413, n4009, n13075);
  and g57763 (n32012, n_24410, n_24411, n_24412, n_24413);
  nor g57764 (n32079, n32073, n32074, n32075, n32078);
  nor g57765 (n32093, n32087, n32088, n32089, n32090);
endmodule

