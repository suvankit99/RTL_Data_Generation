
module router(\dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] ,
     \dest_x[4] , \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] ,
     \dest_x[9] , \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13]
     , \dest_x[14] , \dest_x[15] , \dest_x[16] , \dest_x[17] ,
     \dest_x[18] , \dest_x[19] , \dest_x[20] , \dest_x[21] ,
     \dest_x[22] , \dest_x[23] , \dest_x[24] , \dest_x[25] ,
     \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] , \dest_y[0]
     , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] , \dest_y[5] ,
     \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] , \dest_y[10] ,
     \dest_y[11] , \dest_y[12] , \dest_y[13] , \dest_y[14] ,
     \dest_y[15] , \dest_y[16] , \dest_y[17] , \dest_y[18] ,
     \dest_y[19] , \dest_y[20] , \dest_y[21] , \dest_y[22] ,
     \dest_y[23] , \dest_y[24] , \dest_y[25] , \dest_y[26] ,
     \dest_y[27] , \dest_y[28] , \dest_y[29] , \outport[0] ,
     \outport[1] , \outport[2] , \outport[3] , \outport[4] ,
     \outport[5] , \outport[6] , \outport[7] , \outport[8] ,
     \outport[9] , \outport[10] , \outport[11] , \outport[12] ,
     \outport[13] , \outport[14] , \outport[15] , \outport[16] ,
     \outport[17] , \outport[18] , \outport[19] , \outport[20] ,
     \outport[21] , \outport[22] , \outport[23] , \outport[24] ,
     \outport[25] , \outport[26] , \outport[27] , \outport[28] ,
     \outport[29] );
  input \dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] , \dest_x[4]
       , \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] , \dest_x[9]
       , \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13] ,
       \dest_x[14] , \dest_x[15] , \dest_x[16] , \dest_x[17] ,
       \dest_x[18] , \dest_x[19] , \dest_x[20] , \dest_x[21] ,
       \dest_x[22] , \dest_x[23] , \dest_x[24] , \dest_x[25] ,
       \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] ,
       \dest_y[0] , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] ,
       \dest_y[5] , \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] ,
       \dest_y[10] , \dest_y[11] , \dest_y[12] , \dest_y[13] ,
       \dest_y[14] , \dest_y[15] , \dest_y[16] , \dest_y[17] ,
       \dest_y[18] , \dest_y[19] , \dest_y[20] , \dest_y[21] ,
       \dest_y[22] , \dest_y[23] , \dest_y[24] , \dest_y[25] ,
       \dest_y[26] , \dest_y[27] , \dest_y[28] , \dest_y[29] ;
  output \outport[0] , \outport[1] , \outport[2] , \outport[3] ,
       \outport[4] , \outport[5] , \outport[6] , \outport[7] ,
       \outport[8] , \outport[9] , \outport[10] , \outport[11] ,
       \outport[12] , \outport[13] , \outport[14] , \outport[15] ,
       \outport[16] , \outport[17] , \outport[18] , \outport[19] ,
       \outport[20] , \outport[21] , \outport[22] , \outport[23] ,
       \outport[24] , \outport[25] , \outport[26] , \outport[27] ,
       \outport[28] , \outport[29] ;
  wire \dest_x[0] , \dest_x[1] , \dest_x[2] , \dest_x[3] , \dest_x[4] ,
       \dest_x[5] , \dest_x[6] , \dest_x[7] , \dest_x[8] , \dest_x[9] ,
       \dest_x[10] , \dest_x[11] , \dest_x[12] , \dest_x[13] ,
       \dest_x[14] , \dest_x[15] , \dest_x[16] , \dest_x[17] ,
       \dest_x[18] , \dest_x[19] , \dest_x[20] , \dest_x[21] ,
       \dest_x[22] , \dest_x[23] , \dest_x[24] , \dest_x[25] ,
       \dest_x[26] , \dest_x[27] , \dest_x[28] , \dest_x[29] ,
       \dest_y[0] , \dest_y[1] , \dest_y[2] , \dest_y[3] , \dest_y[4] ,
       \dest_y[5] , \dest_y[6] , \dest_y[7] , \dest_y[8] , \dest_y[9] ,
       \dest_y[10] , \dest_y[11] , \dest_y[12] , \dest_y[13] ,
       \dest_y[14] , \dest_y[15] , \dest_y[16] , \dest_y[17] ,
       \dest_y[18] , \dest_y[19] , \dest_y[20] , \dest_y[21] ,
       \dest_y[22] , \dest_y[23] , \dest_y[24] , \dest_y[25] ,
       \dest_y[26] , \dest_y[27] , \dest_y[28] , \dest_y[29] ;
  wire \outport[0] , \outport[1] , \outport[2] , \outport[3] ,
       \outport[4] , \outport[5] , \outport[6] , \outport[7] ,
       \outport[8] , \outport[9] , \outport[10] , \outport[11] ,
       \outport[12] , \outport[13] , \outport[14] , \outport[15] ,
       \outport[16] , \outport[17] , \outport[18] , \outport[19] ,
       \outport[20] , \outport[21] , \outport[22] , \outport[23] ,
       \outport[24] , \outport[25] , \outport[26] , \outport[27] ,
       \outport[28] , \outport[29] ;
  wire n92, n93, n94, n95, n96, n97, n98, n99;
  wire n100, n101, n102, n103, n104, n105, n106, n107;
  wire n108, n109, n110, n111, n112, n113, n114, n115;
  wire n116, n117, n118, n119, n120, n121, n122, n123;
  wire n124, n125, n126, n127, n128, n129, n130, n131;
  wire n132, n133, n134, n135, n136, n137, n138, n139;
  wire n140, n141, n142, n143, n144, n145, n146, n147;
  wire n148, n149, n150, n151, n152, n153, n154, n155;
  wire n156, n185, n186, n187, n214, n215, n217, n218;
  wire n219, n220, n221, n222, n223, n224, n225, n226;
  wire n227, n228, n229, n230, n231, n232, n233, n234;
  wire n235, n236, n237, n238, n239, n240, n241, n242;
  wire n243, n244, n245, n246, n247, n248, n249, n250;
  wire n251, n252, n253, n254, n255, n256, n257, n258;
  wire n259, n260, n261, n262, n263, n264, n265, n266;
  wire n267, n268, n269, n270, n271, n272, n273, n274;
  wire n275, n276, n277, n278, n279, n280, n281, n282;
  wire n311, n338, n339, n340, n341, n342, n343, n345;
  wire n346, n347, n_30, n_31, n_32, n_33, n_35, n_36;
  wire n_37, n_39, n_40, n_41, n_43, n_44, n_45, n_47;
  wire n_48, n_49, n_51, n_52, n_53, n_55, n_56, n_57;
  wire n_58, n_60, n_61, n_62, n_64, n_65, n_66, n_68;
  wire n_69, n_70, n_72, n_73, n_74, n_76, n_77, n_78;
  wire n_79, n_81, n_82, n_83, n_85, n_86, n_87, n_89;
  wire n_90, n_91, n_93, n_94, n_95, n_96, n_98, n_99;
  wire n_100, n_101, n_103, n_104, n_105, n_107, n_108, n_109;
  wire n_111, n_112, n_113, n_114, n_138, n_139, n_154, n_157;
  wire n_158, n_160, n_162, n_163, n_165, n_167, n_170, n_171;
  wire n_173, n_175, n_176, n_178, n_181, n_182, n_184, n_186;
  wire n_190, n_191, n_193, n_196, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_289, n_290, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361;
  assign \outport[29]  = 1'b0;
//   assign \outport[28]  = 1'b0;
  assign \outport[27]  = 1'b0;
  assign \outport[26]  = 1'b0;
  assign \outport[25]  = 1'b0;
//   assign \outport[24]  = 1'b0;
  assign \outport[23]  = 1'b0;
  assign \outport[22]  = 1'b0;
  assign \outport[21]  = 1'b0;
  assign \outport[20]  = 1'b0;
//   assign \outport[19]  = 1'b0;
  assign \outport[18]  = 1'b0;
  assign \outport[17]  = 1'b0;
//   assign \outport[16]  = 1'b0;
//   assign \outport[15]  = 1'b0;
  assign \outport[14]  = 1'b0;
  assign \outport[13]  = 1'b0;
  assign \outport[12]  = 1'b0;
//   assign \outport[11]  = 1'b0;
  assign \outport[10]  = 1'b0;
  assign \outport[9]  = 1'b0;
  assign \outport[8]  = 1'b0;
  assign \outport[7]  = 1'b0;
  assign \outport[6]  = 1'b0;
  assign \outport[5]  = 1'b0;
  assign \outport[4]  = 1'b0;
  assign \outport[3]  = 1'b0;
  not g1 (n_30, \dest_x[9] );
  not g2 (n_31, \dest_x[10] );
  and g3 (n92, n_30, n_31);
  and g4 (n93, \dest_x[9] , \dest_x[10] );
  not g5 (n_32, n92);
  not g6 (n_33, n93);
  and g7 (n94, n_32, n_33);
  and g8 (n95, \dest_x[11] , n_32);
  not g9 (n_35, \dest_x[11] );
  and g10 (n96, n_35, n92);
  not g11 (n_36, n95);
  not g12 (n_37, n96);
  and g13 (n97, n_36, n_37);
  not g14 (n_39, \dest_x[12] );
  and g15 (n98, n_39, n_36);
  and g16 (n99, \dest_x[12] , n95);
  not g17 (n_40, n98);
  not g18 (n_41, n99);
  and g19 (n100, n_40, n_41);
  not g20 (n_43, \dest_x[13] );
  and g21 (n101, n_43, n98);
  and g22 (n102, \dest_x[13] , n_40);
  not g23 (n_44, n101);
  not g24 (n_45, n102);
  and g25 (n103, n_44, n_45);
  and g26 (n104, \dest_x[14] , n_44);
  not g27 (n_47, \dest_x[14] );
  and g28 (n105, n_47, n101);
  not g29 (n_48, n104);
  not g30 (n_49, n105);
  and g31 (n106, n_48, n_49);
  and g32 (n107, \dest_x[15] , n_48);
  not g33 (n_51, \dest_x[15] );
  and g34 (n108, n_51, n104);
  not g35 (n_52, n107);
  not g36 (n_53, n108);
  and g37 (n109, n_52, n_53);
  and g38 (n110, \dest_x[15] , n104);
  not g39 (n_55, \dest_x[16] );
  not g40 (n_56, n110);
  and g41 (n111, n_55, n_56);
  and g42 (n112, \dest_x[16] , n110);
  not g43 (n_57, n111);
  not g44 (n_58, n112);
  and g45 (n113, n_57, n_58);
  and g46 (n114, \dest_x[17] , n_57);
  not g47 (n_60, \dest_x[17] );
  and g48 (n115, n_60, n111);
  not g49 (n_61, n114);
  not g50 (n_62, n115);
  and g51 (n116, n_61, n_62);
  not g52 (n_64, \dest_x[18] );
  and g53 (n117, n_64, n_61);
  and g54 (n118, \dest_x[18] , n114);
  not g55 (n_65, n117);
  not g56 (n_66, n118);
  and g57 (n119, n_65, n_66);
  and g58 (n120, \dest_x[19] , n_65);
  not g59 (n_68, \dest_x[19] );
  and g60 (n121, n_68, n117);
  not g61 (n_69, n120);
  not g62 (n_70, n121);
  and g63 (n122, n_69, n_70);
  and g64 (n123, \dest_x[20] , n_69);
  not g65 (n_72, \dest_x[20] );
  and g66 (n124, n_72, n120);
  not g67 (n_73, n123);
  not g68 (n_74, n124);
  and g69 (n125, n_73, n_74);
  and g70 (n126, \dest_x[20] , n120);
  not g71 (n_76, \dest_x[21] );
  not g72 (n_77, n126);
  and g73 (n127, n_76, n_77);
  and g74 (n128, \dest_x[21] , n126);
  not g75 (n_78, n127);
  not g76 (n_79, n128);
  and g77 (n129, n_78, n_79);
  not g78 (n_81, \dest_x[22] );
  and g79 (n130, n_81, n127);
  and g80 (n131, \dest_x[22] , n_78);
  not g81 (n_82, n130);
  not g82 (n_83, n131);
  and g83 (n132, n_82, n_83);
  and g84 (n133, \dest_x[23] , n_82);
  not g85 (n_85, \dest_x[23] );
  and g86 (n134, n_85, n130);
  not g87 (n_86, n133);
  not g88 (n_87, n134);
  and g89 (n135, n_86, n_87);
  and g90 (n136, \dest_x[24] , n_86);
  not g91 (n_89, \dest_x[24] );
  and g92 (n137, n_89, n133);
  not g93 (n_90, n136);
  not g94 (n_91, n137);
  and g95 (n138, n_90, n_91);
  and g96 (n139, \dest_x[24] , n133);
  not g97 (n_93, n139);
  and g98 (n140, \dest_x[25] , n_93);
  not g99 (n_94, \dest_x[25] );
  and g100 (n141, n_94, n139);
  not g101 (n_95, n140);
  not g102 (n_96, n141);
  and g103 (n142, n_95, n_96);
  and g104 (n143, \dest_x[25] , n139);
  not g105 (n_98, \dest_x[26] );
  not g106 (n_99, n143);
  and g107 (n144, n_98, n_99);
  and g108 (n145, \dest_x[26] , n143);
  not g109 (n_100, n144);
  not g110 (n_101, n145);
  and g111 (n146, n_100, n_101);
  and g112 (n147, \dest_x[27] , n_100);
  not g113 (n_103, \dest_x[27] );
  and g114 (n148, n_103, n144);
  not g115 (n_104, n147);
  not g116 (n_105, n148);
  and g117 (n149, n_104, n_105);
  and g118 (n150, \dest_x[28] , n_104);
  not g119 (n_107, \dest_x[28] );
  and g120 (n151, n_107, n147);
  not g121 (n_108, n150);
  not g122 (n_109, n151);
  and g123 (n152, n_108, n_109);
  and g124 (n153, \dest_x[28] , n147);
  not g125 (n_111, \dest_x[29] );
  and g126 (n154, n_111, n153);
  not g127 (n_112, n153);
  and g128 (n155, \dest_x[29] , n_112);
  not g129 (n_113, n154);
  not g130 (n_114, n155);
  and g131 (n156, n_113, n_114);
  and g175 (n186, \dest_x[29] , n153);
  not g176 (n_138, n185);
  not g177 (n_139, n186);
  and g178 (n187, n_138, n_139);
  not g220 (n_154, n214);
  and g221 (n215, n186, n_154);
  or g222 (\outport[0] , n187, n215);
  not g223 (n_157, \dest_y[9] );
  not g224 (n_158, \dest_y[10] );
  and g225 (n217, n_157, n_158);
  not g226 (n_160, n217);
  and g227 (n218, \dest_y[11] , n_160);
  not g228 (n_162, \dest_y[12] );
  not g229 (n_163, n218);
  and g230 (n219, n_162, n_163);
  not g231 (n_165, \dest_y[13] );
  and g232 (n220, n_165, n219);
  not g233 (n_167, n220);
  and g234 (n221, \dest_y[14] , n_167);
  and g235 (n222, \dest_y[15] , n221);
  not g236 (n_170, \dest_y[16] );
  not g237 (n_171, n222);
  and g238 (n223, n_170, n_171);
  not g239 (n_173, n223);
  and g240 (n224, \dest_y[17] , n_173);
  not g241 (n_175, \dest_y[18] );
  not g242 (n_176, n224);
  and g243 (n225, n_175, n_176);
  not g244 (n_178, n225);
  and g245 (n226, \dest_y[19] , n_178);
  and g246 (n227, \dest_y[20] , n226);
  not g247 (n_181, \dest_y[21] );
  not g248 (n_182, n227);
  and g249 (n228, n_181, n_182);
  not g250 (n_184, \dest_y[22] );
  and g251 (n229, n_184, n228);
  not g252 (n_186, n229);
  and g253 (n230, \dest_y[23] , n_186);
  and g254 (n231, \dest_y[24] , n230);
  and g255 (n232, \dest_y[25] , n231);
  not g256 (n_190, \dest_y[26] );
  not g257 (n_191, n232);
  and g258 (n233, n_190, n_191);
  not g259 (n_193, n233);
  and g260 (n234, \dest_y[27] , n_193);
  and g261 (n235, \dest_y[28] , n234);
  and g262 (n236, \dest_y[29] , n235);
  not g263 (n_196, n236);
  and g264 (n237, \dest_x[0] , n_196);
  not g265 (n_198, \dest_x[0] );
  not g266 (n_199, \dest_y[0] );
  and g267 (n238, n_198, n_199);
  not g268 (n_200, n238);
  and g269 (n239, n236, n_200);
  and g270 (n240, \dest_y[9] , \dest_y[10] );
  not g271 (n_201, n240);
  and g272 (n241, n_160, n_201);
  not g273 (n_202, \dest_y[11] );
  and g274 (n242, n_202, n217);
  not g275 (n_203, n242);
  and g276 (n243, n_163, n_203);
  and g277 (n244, \dest_y[12] , n218);
  not g278 (n_204, n219);
  not g279 (n_205, n244);
  and g280 (n245, n_204, n_205);
  and g281 (n246, \dest_y[13] , n_204);
  not g282 (n_206, n246);
  and g283 (n247, n_167, n_206);
  not g284 (n_207, \dest_y[14] );
  and g285 (n248, n_207, n220);
  not g286 (n_208, n221);
  not g287 (n_209, n248);
  and g288 (n249, n_208, n_209);
  and g289 (n250, \dest_y[15] , n_208);
  not g290 (n_210, \dest_y[15] );
  and g291 (n251, n_210, n221);
  not g292 (n_211, n250);
  not g293 (n_212, n251);
  and g294 (n252, n_211, n_212);
  and g295 (n253, \dest_y[16] , n222);
  not g296 (n_213, n253);
  and g297 (n254, n_173, n_213);
  not g298 (n_214, \dest_y[17] );
  and g299 (n255, n_214, n223);
  not g300 (n_215, n255);
  and g301 (n256, n_176, n_215);
  and g302 (n257, \dest_y[18] , n224);
  not g303 (n_216, n257);
  and g304 (n258, n_178, n_216);
  not g305 (n_217, \dest_y[19] );
  and g306 (n259, n_217, n225);
  not g307 (n_218, n226);
  not g308 (n_219, n259);
  and g309 (n260, n_218, n_219);
  and g310 (n261, \dest_y[20] , n_218);
  not g311 (n_220, \dest_y[20] );
  and g312 (n262, n_220, n226);
  not g313 (n_221, n261);
  not g314 (n_222, n262);
  and g315 (n263, n_221, n_222);
  and g316 (n264, \dest_y[21] , n227);
  not g317 (n_223, n228);
  not g318 (n_224, n264);
  and g319 (n265, n_223, n_224);
  and g320 (n266, \dest_y[22] , n_223);
  not g321 (n_225, n266);
  and g322 (n267, n_186, n_225);
  not g323 (n_226, \dest_y[23] );
  and g324 (n268, n_226, n229);
  not g325 (n_227, n230);
  not g326 (n_228, n268);
  and g327 (n269, n_227, n_228);
  and g328 (n270, \dest_y[24] , n_227);
  not g329 (n_229, \dest_y[24] );
  and g330 (n271, n_229, n230);
  not g331 (n_230, n270);
  not g332 (n_231, n271);
  and g333 (n272, n_230, n_231);
  not g334 (n_232, n231);
  and g335 (n273, \dest_y[25] , n_232);
  not g336 (n_233, \dest_y[25] );
  and g337 (n274, n_233, n231);
  not g338 (n_234, n273);
  not g339 (n_235, n274);
  and g340 (n275, n_234, n_235);
  and g341 (n276, \dest_y[26] , n232);
  not g342 (n_236, n276);
  and g343 (n277, n_193, n_236);
  not g344 (n_237, \dest_y[27] );
  and g345 (n278, n_237, n233);
  not g346 (n_238, n234);
  not g347 (n_239, n278);
  and g348 (n279, n_238, n_239);
  and g349 (n280, \dest_y[28] , n_238);
  not g350 (n_240, \dest_y[28] );
  and g351 (n281, n_240, n234);
  not g352 (n_241, n280);
  not g353 (n_242, n281);
  and g354 (n282, n_241, n_242);
  not g438 (n_278, n338);
  and g439 (n339, n236, n_278);
  not g440 (n_279, n311);
  not g441 (n_280, n339);
  and g442 (n340, n_279, n_280);
  not g443 (n_281, n239);
  and g444 (n341, n_281, n340);
  not g445 (n_282, n187);
  not g446 (n_283, n341);
  and g447 (n342, n_282, n_283);
  not g448 (n_284, n237);
  and g449 (n343, n_284, n342);
  not g450 (n_285, n215);
  not g451 (n_286, n343);
  and g452 (\outport[1] , n_285, n_286);
  and g453 (n345, \dest_x[0] , n236);
  and g454 (n346, \dest_y[0] , n345);
  not g455 (n_287, n346);
  and g456 (n347, n_280, n_287);
  not g457 (n_289, \outport[0] );
  not g458 (n_290, n347);
  and g459 (\outport[2] , n_289, n_290);
  nor g460 (n_293, n94, n100);
  nor g461 (n_294, n103, n109);
  nor g462 (n_295, n113, n119);
  nor g463 (n_296, n125, n129);
  nor g464 (n_297, n132, n138);
  nor g465 (n_298, n142, n146);
  nor g466 (n_299, n152, n156);
  and g467 (n_300, \dest_x[0] , \dest_x[1] );
  and g468 (n_301, \dest_x[2] , \dest_x[3] );
  and g469 (n_302, \dest_x[4] , \dest_x[5] );
  and g470 (n_303, \dest_x[6] , \dest_x[7] );
  and g471 (n_304, \dest_x[8] , n97);
  and g472 (n_305, n106, n116);
  and g473 (n_306, n122, n135);
  and g474 (n_307, n149, n_30, n_293, n_294);
  and g475 (n_308, n_295, n_296, n_297, n_298);
  and g476 (n_309, n_299, n_300, n_301, n_302);
  and g477 (n_310, n_303, n_304, n_305, n_306);
  and g478 (n185, n_307, n_308, n_309, n_310);
  nor g479 (n_311, n149, n135);
  nor g480 (n_312, n122, n116);
  nor g481 (n_313, n106, n97);
  nor g482 (n_314, \dest_x[8] , \dest_x[7] );
  nor g483 (n_315, \dest_x[6] , \dest_x[5] );
  nor g484 (n_316, \dest_x[4] , \dest_x[3] );
  nor g485 (n_317, \dest_x[1] , \dest_x[2] );
  and g486 (n_318, \dest_x[9] , n152);
  and g487 (n_319, n146, n142);
  and g488 (n_320, n138, n132);
  and g489 (n_321, n129, n125);
  and g490 (n_322, n119, n113);
  and g491 (n_323, n109, n103, n100, n94);
  and g492 (n_324, n_311, n_312, n_313, n_314);
  and g493 (n_325, n_315, n_316, n_317, n_318);
  and g494 (n_326, n_319, n_320, n_321, n_322);
  and g495 (n214, n_323, n_324, n_325, n_326);
  nor g496 (n_328, n241, n245);
  nor g497 (n_329, n247, n252);
  nor g498 (n_330, n254, n258);
  nor g499 (n_331, n263, n265);
  nor g500 (n_332, n267, n272);
  nor g501 (n_333, n275, n277);
  and g502 (n_334, n_327, \dest_y[1] );
  not g503 (n_327, n282);
  and g504 (n_335, \dest_y[2] , \dest_y[3] );
  and g505 (n_336, \dest_y[4] , \dest_y[5] );
  and g506 (n_337, \dest_y[6] , \dest_y[7] );
  and g507 (n_338, \dest_y[8] , n243);
  and g508 (n_339, n249, n256);
  and g509 (n_340, n260, n269);
  and g510 (n_341, n279, \dest_y[29] );
  and g511 (n_342, \dest_y[0] , n_157, n_328, n_329);
  and g512 (n_343, n_330, n_331, n_332, n_333);
  and g513 (n_344, n_334, n_335, n_336, n_337);
  and g514 (n_345, n_338, n_339, n_340, n_341);
  and g515 (n311, n_342, n_343, n_344, n_345);
  nor g516 (n_346, n279, n269);
  nor g517 (n_347, n260, n256);
  nor g518 (n_348, n249, n243);
  nor g519 (n_349, \dest_y[8] , \dest_y[7] );
  nor g520 (n_350, \dest_y[6] , \dest_y[5] );
  nor g521 (n_351, \dest_y[4] , \dest_y[3] );
  nor g522 (n_352, \dest_y[1] , \dest_y[2] );
  and g523 (n_353, \dest_y[9] , n282);
  and g524 (n_354, n277, n275);
  and g525 (n_355, n272, n267);
  and g526 (n_356, n265, n263);
  and g527 (n_357, n258, n254);
  and g528 (n_358, n252, n247, n245, n241);
  and g529 (n_359, n_346, n_347, n_348, n_349);
  and g530 (n_360, n_350, n_351, n_352, n_353);
  and g531 (n_361, n_354, n_355, n_356, n_357);
  and g532 (n338, n_358, n_359, n_360, n_361);
endmodule

