
module sqrt(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] ,
     \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14]
     , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
     \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
     \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
     \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
     \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
     \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
     \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
     \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
     \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
     \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
     \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
     \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
     \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105]
     , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] ,
     \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
     \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
     \a[124] , \a[125] , \a[126] , \a[127] , \asqrt[0] , \asqrt[1] ,
     \asqrt[2] , \asqrt[3] , \asqrt[4] , \asqrt[5] , \asqrt[6] ,
     \asqrt[7] , \asqrt[8] , \asqrt[9] , \asqrt[10] , \asqrt[11] ,
     \asqrt[12] , \asqrt[13] , \asqrt[14] , \asqrt[15] , \asqrt[16] ,
     \asqrt[17] , \asqrt[18] , \asqrt[19] , \asqrt[20] , \asqrt[21] ,
     \asqrt[22] , \asqrt[23] , \asqrt[24] , \asqrt[25] , \asqrt[26] ,
     \asqrt[27] , \asqrt[28] , \asqrt[29] , \asqrt[30] , \asqrt[31] ,
     \asqrt[32] , \asqrt[33] , \asqrt[34] , \asqrt[35] , \asqrt[36] ,
     \asqrt[37] , \asqrt[38] , \asqrt[39] , \asqrt[40] , \asqrt[41] ,
     \asqrt[42] , \asqrt[43] , \asqrt[44] , \asqrt[45] , \asqrt[46] ,
     \asqrt[47] , \asqrt[48] , \asqrt[49] , \asqrt[50] , \asqrt[51] ,
     \asqrt[52] , \asqrt[53] , \asqrt[54] , \asqrt[55] , \asqrt[56] ,
     \asqrt[57] , \asqrt[58] , \asqrt[59] , \asqrt[60] , \asqrt[61] ,
     \asqrt[62] , \asqrt[63] );
//   input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
       \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
       \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
       \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
       \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
       \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] ,
       \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
       \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
       \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] ,
       \a[123] , \a[124] , \a[125] , \a[126] , \a[127] ;
//   output \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
       \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
       \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
       \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
       \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
       \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
       \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
       \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
       \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
       \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
       \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
       \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
       \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
       \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
       \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
       \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
       \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
       \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] ,
       \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
       \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
       \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] ,
       \a[123] , \a[124] , \a[125] , \a[126] , \a[127] ;
  wire \asqrt[0] , \asqrt[1] , \asqrt[2] , \asqrt[3] , \asqrt[4] ,
       \asqrt[5] , \asqrt[6] , \asqrt[7] , \asqrt[8] , \asqrt[9] ,
       \asqrt[10] , \asqrt[11] , \asqrt[12] , \asqrt[13] , \asqrt[14] ,
       \asqrt[15] , \asqrt[16] , \asqrt[17] , \asqrt[18] , \asqrt[19] ,
       \asqrt[20] , \asqrt[21] , \asqrt[22] , \asqrt[23] , \asqrt[24] ,
       \asqrt[25] , \asqrt[26] , \asqrt[27] , \asqrt[28] , \asqrt[29] ,
       \asqrt[30] , \asqrt[31] , \asqrt[32] , \asqrt[33] , \asqrt[34] ,
       \asqrt[35] , \asqrt[36] , \asqrt[37] , \asqrt[38] , \asqrt[39] ,
       \asqrt[40] , \asqrt[41] , \asqrt[42] , \asqrt[43] , \asqrt[44] ,
       \asqrt[45] , \asqrt[46] , \asqrt[47] , \asqrt[48] , \asqrt[49] ,
       \asqrt[50] , \asqrt[51] , \asqrt[52] , \asqrt[53] , \asqrt[54] ,
       \asqrt[55] , \asqrt[56] , \asqrt[57] , \asqrt[58] , \asqrt[59] ,
       \asqrt[60] , \asqrt[61] , \asqrt[62] , \asqrt[63] ;
  wire n194, n195, n196, n197, n199, n200, n201, n202;
  wire n203, n204, n205, n206, n207, n208, n209, n210;
  wire n211, n212, n213, n214, n216, n217, n218, n219;
  wire n220, n223, n224, n225, n226, n227, n228, n229;
  wire n232, n233, n234, n235, n236, n237, n238, n241;
  wire n242, n243, n244, n245, n246, n247, n250, n254;
  wire n255, n256, n257, n258, n259, n260, n261, n262;
  wire n266, n267, n268, n269, n270, n271, n275, n276;
  wire n277, n278, n279, n280, n281, n282, n283, n284;
  wire n285, n286, n287, n288, n289, n290, n293, n294;
  wire n295, n296, n297, n298, n299, n300, n305, n309;
  wire n310, n311, n312, n313, n318, n319, n320, n321;
  wire n322, n323, n324, n325, n326, n327, n331, n332;
  wire n333, n334, n335, n336, n337, n338, n339, n340;
  wire n341, n344, n345, n346, n347, n348, n349, n350;
  wire n353, n354, n355, n356, n357, n358, n359, n362;
  wire n363, n364, n365, n366, n367, n368, n369, n374;
  wire n378, n379, n380, n381, n382, n387, n388, n389;
  wire n390, n391, n392, n393, n394, n395, n396, n400;
  wire n401, n402, n403, n404, n405, n406, n407, n408;
  wire n409, n410, n411, n412, n413, n414, n415, n416;
  wire n417, n418, n419, n422, n423, n424, n425, n426;
  wire n427, n428, n429, n430, n433, n434, n435, n436;
  wire n437, n438, n439, n442, n443, n444, n445, n446;
  wire n447, n448, n449, n454, n458, n459, n460, n461;
  wire n462, n467, n468, n469, n470, n471, n472, n473;
  wire n474, n475, n476, n480, n481, n482, n483, n484;
  wire n485, n486, n487, n488, n489, n490, n491, n492;
  wire n493, n494, n495, n496, n497, n498, n499, n502;
  wire n503, n504, n505, n506, n507, n508, n509, n510;
  wire n511, n514, n515, n516, n517, n518, n519, n520;
  wire n521, n522, n525, n526, n527, n528, n529, n530;
  wire n531, n534, n535, n536, n537, n538, n539, n540;
  wire n541, n546, n550, n551, n552, n553, n554, n555;
  wire n556, n557, n558, n563, n564, n565, n566, n567;
  wire n568, n572, n573, n574, n575, n576, n577, n578;
  wire n579, n580, n581, n582, n583, n584, n585, n586;
  wire n587, n588, n589, n590, n591, n594, n595, n596;
  wire n597, n598, n599, n600, n601, n602, n603, n606;
  wire n607, n608, n609, n610, n611, n612, n613, n614;
  wire n615, n618, n619, n620, n621, n622, n623, n624;
  wire n625, n626, n629, n630, n631, n632, n633, n634;
  wire n635, n638, n639, n640, n641, n642, n643, n644;
  wire n645, n650, n654, n655, n656, n657, n658, n663;
  wire n664, n665, n666, n667, n668, n669, n670, n671;
  wire n672, n676, n677, n678, n679, n680, n681, n682;
  wire n683, n684, n685, n686, n689, n690, n691, n692;
  wire n693, n694, n695, n696, n699, n700, n701, n702;
  wire n703, n704, n705, n706, n707, n708, n711, n712;
  wire n713, n714, n715, n716, n717, n718, n719, n720;
  wire n723, n724, n725, n726, n727, n728, n729, n730;
  wire n731, n732, n735, n736, n737, n738, n739, n740;
  wire n741, n742, n743, n746, n747, n748, n749, n750;
  wire n751, n752, n755, n756, n757, n758, n759, n760;
  wire n761, n762, n767, n771, n772, n773, n774, n775;
  wire n780, n781, n782, n783, n784, n785, n786, n787;
  wire n788, n789, n793, n794, n795, n796, n797, n798;
  wire n799, n800, n801, n802, n803, n804, n805, n806;
  wire n807, n808, n809, n810, n811, n812, n815, n816;
  wire n817, n818, n819, n820, n821, n822, n823, n824;
  wire n825, n826, n829, n830, n831, n832, n833, n834;
  wire n835, n836, n839, n840, n841, n842, n843, n844;
  wire n845, n846, n847, n848, n851, n852, n853, n854;
  wire n855, n856, n857, n858, n859, n860, n863, n864;
  wire n865, n866, n867, n868, n869, n870, n871, n874;
  wire n875, n876, n877, n878, n879, n880, n883, n884;
  wire n885, n886, n887, n888, n889, n890, n895, n899;
  wire n900, n901, n902, n903, n908, n909, n910, n911;
  wire n912, n913, n914, n915, n916, n917, n921, n922;
  wire n923, n924, n925, n926, n927, n928, n929, n930;
  wire n931, n932, n933, n934, n935, n936, n937, n938;
  wire n939, n940, n943, n944, n945, n946, n947, n948;
  wire n949, n950, n951, n952, n955, n956, n957, n958;
  wire n959, n960, n961, n962, n963, n964, n967, n968;
  wire n969, n970, n971, n972, n973, n974, n975, n976;
  wire n977, n978, n981, n982, n983, n984, n985, n986;
  wire n987, n988, n991, n992, n993, n994, n995, n996;
  wire n997, n998, n999, n1000, n1003, n1004, n1005, n1006;
  wire n1007, n1008, n1009, n1010, n1011, n1014, n1015, n1016;
  wire n1017, n1018, n1019, n1020, n1023, n1024, n1025, n1026;
  wire n1027, n1028, n1029, n1030, n1035, n1039, n1040, n1041;
  wire n1042, n1043, n1048, n1049, n1050, n1051, n1052, n1053;
  wire n1054, n1055, n1056, n1057, n1061, n1062, n1063, n1064;
  wire n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072;
  wire n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;
  wire n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090;
  wire n1091, n1092, n1095, n1096, n1097, n1098, n1099, n1100;
  wire n1101, n1102, n1103, n1104, n1107, n1108, n1109, n1110;
  wire n1111, n1112, n1113, n1114, n1115, n1116, n1119, n1120;
  wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
  wire n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138;
  wire n1139, n1140, n1141, n1142, n1145, n1146, n1147, n1148;
  wire n1149, n1150, n1151, n1152, n1155, n1156, n1157, n1158;
  wire n1159, n1160, n1161, n1162, n1163, n1166, n1167, n1168;
  wire n1169, n1170, n1171, n1172, n1175, n1176, n1177, n1178;
  wire n1179, n1180, n1181, n1182, n1187, n1191, n1192, n1193;
  wire n1194, n1195, n1200, n1201, n1202, n1203, n1204, n1205;
  wire n1206, n1207, n1208, n1209, n1213, n1214, n1215, n1216;
  wire n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224;
  wire n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232;
  wire n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242;
  wire n1243, n1244, n1247, n1248, n1249, n1250, n1251, n1252;
  wire n1253, n1254, n1255, n1256, n1259, n1260, n1261, n1262;
  wire n1263, n1264, n1265, n1266, n1267, n1268, n1271, n1272;
  wire n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;
  wire n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290;
  wire n1291, n1292, n1295, n1296, n1297, n1298, n1299, n1300;
  wire n1301, n1302, n1303, n1304, n1307, n1308, n1309, n1310;
  wire n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318;
  wire n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1330;
  wire n1331, n1332, n1333, n1334, n1335, n1336, n1339, n1340;
  wire n1341, n1342, n1343, n1344, n1345, n1346, n1351, n1355;
  wire n1356, n1357, n1358, n1359, n1364, n1365, n1366, n1367;
  wire n1368, n1369, n1370, n1371, n1372, n1373, n1377, n1378;
  wire n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386;
  wire n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394;
  wire n1395, n1396, n1399, n1400, n1401, n1402, n1403, n1404;
  wire n1405, n1406, n1407, n1408, n1411, n1412, n1413, n1414;
  wire n1415, n1416, n1417, n1418, n1419, n1420, n1423, n1424;
  wire n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432;
  wire n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442;
  wire n1443, n1444, n1447, n1448, n1449, n1450, n1451, n1452;
  wire n1453, n1454, n1455, n1456, n1459, n1460, n1461, n1462;
  wire n1463, n1464, n1465, n1466, n1467, n1468, n1471, n1472;
  wire n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480;
  wire n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490;
  wire n1491, n1492, n1495, n1496, n1497, n1498, n1499, n1500;
  wire n1501, n1502, n1503, n1506, n1507, n1508, n1509, n1510;
  wire n1511, n1512, n1515, n1516, n1517, n1518, n1519, n1520;
  wire n1521, n1522, n1527, n1531, n1532, n1533, n1534, n1535;
  wire n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547;
  wire n1548, n1549, n1553, n1554, n1555, n1556, n1557, n1558;
  wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
  wire n1567, n1568, n1569, n1570, n1571, n1572, n1575, n1576;
  wire n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584;
  wire n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594;
  wire n1595, n1596, n1599, n1600, n1601, n1602, n1603, n1604;
  wire n1605, n1606, n1607, n1608, n1611, n1612, n1613, n1614;
  wire n1615, n1616, n1617, n1618, n1619, n1620, n1623, n1624;
  wire n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632;
  wire n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642;
  wire n1643, n1644, n1647, n1648, n1649, n1650, n1651, n1652;
  wire n1653, n1654, n1655, n1656, n1659, n1660, n1661, n1662;
  wire n1663, n1664, n1665, n1666, n1667, n1668, n1671, n1672;
  wire n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680;
  wire n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690;
  wire n1691, n1694, n1695, n1696, n1697, n1698, n1699, n1700;
  wire n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710;
  wire n1715, n1719, n1720, n1721, n1722, n1723, n1724, n1725;
  wire n1726, n1727, n1732, n1733, n1734, n1735, n1736, n1737;
  wire n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748;
  wire n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756;
  wire n1757, n1758, n1759, n1760, n1763, n1764, n1765, n1766;
  wire n1767, n1768, n1769, n1770, n1771, n1772, n1775, n1776;
  wire n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784;
  wire n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794;
  wire n1795, n1796, n1799, n1800, n1801, n1802, n1803, n1804;
  wire n1805, n1806, n1807, n1808, n1811, n1812, n1813, n1814;
  wire n1815, n1816, n1817, n1818, n1819, n1820, n1823, n1824;
  wire n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832;
  wire n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842;
  wire n1843, n1844, n1847, n1848, n1849, n1850, n1851, n1852;
  wire n1853, n1854, n1855, n1856, n1859, n1860, n1861, n1862;
  wire n1863, n1864, n1865, n1866, n1867, n1868, n1871, n1872;
  wire n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880;
  wire n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890;
  wire n1891, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
  wire n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910;
  wire n1915, n1919, n1920, n1921, n1922, n1923, n1928, n1929;
  wire n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937;
  wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
  wire n1949, n1950, n1951, n1954, n1955, n1956, n1957, n1958;
  wire n1959, n1960, n1961, n1964, n1965, n1966, n1967, n1968;
  wire n1969, n1970, n1971, n1972, n1973, n1976, n1977, n1978;
  wire n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1988;
  wire n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996;
  wire n1997, n2000, n2001, n2002, n2003, n2004, n2005, n2006;
  wire n2007, n2008, n2009, n2012, n2013, n2014, n2015, n2016;
  wire n2017, n2018, n2019, n2020, n2021, n2024, n2025, n2026;
  wire n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2036;
  wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
  wire n2045, n2048, n2049, n2050, n2051, n2052, n2053, n2054;
  wire n2055, n2056, n2057, n2060, n2061, n2062, n2063, n2064;
  wire n2065, n2066, n2067, n2068, n2069, n2072, n2073, n2074;
  wire n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2084;
  wire n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092;
  wire n2093, n2096, n2097, n2098, n2099, n2100, n2101, n2102;
  wire n2103, n2104, n2107, n2108, n2109, n2110, n2111, n2112;
  wire n2113, n2116, n2117, n2118, n2119, n2120, n2121, n2122;
  wire n2123, n2128, n2132, n2133, n2134, n2135, n2136, n2141;
  wire n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149;
  wire n2150, n2154, n2155, n2156, n2157, n2158, n2159, n2160;
  wire n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168;
  wire n2169, n2170, n2171, n2172, n2173, n2176, n2177, n2178;
  wire n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186;
  wire n2187, n2190, n2191, n2192, n2193, n2194, n2195, n2196;
  wire n2197, n2200, n2201, n2202, n2203, n2204, n2205, n2206;
  wire n2207, n2208, n2209, n2212, n2213, n2214, n2215, n2216;
  wire n2217, n2218, n2219, n2220, n2221, n2224, n2225, n2226;
  wire n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2236;
  wire n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244;
  wire n2245, n2248, n2249, n2250, n2251, n2252, n2253, n2254;
  wire n2255, n2256, n2257, n2260, n2261, n2262, n2263, n2264;
  wire n2265, n2266, n2267, n2268, n2269, n2272, n2273, n2274;
  wire n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2284;
  wire n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292;
  wire n2293, n2296, n2297, n2298, n2299, n2300, n2301, n2302;
  wire n2303, n2304, n2305, n2308, n2309, n2310, n2311, n2312;
  wire n2313, n2314, n2315, n2316, n2317, n2320, n2321, n2322;
  wire n2323, n2324, n2325, n2326, n2327, n2328, n2331, n2332;
  wire n2333, n2334, n2335, n2336, n2337, n2340, n2341, n2342;
  wire n2343, n2344, n2345, n2346, n2347, n2352, n2356, n2357;
  wire n2358, n2359, n2360, n2365, n2366, n2367, n2368, n2369;
  wire n2370, n2371, n2372, n2373, n2374, n2378, n2379, n2380;
  wire n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388;
  wire n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396;
  wire n2397, n2400, n2401, n2402, n2403, n2404, n2405, n2406;
  wire n2407, n2408, n2409, n2412, n2413, n2414, n2415, n2416;
  wire n2417, n2418, n2419, n2420, n2421, n2424, n2425, n2426;
  wire n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434;
  wire n2435, n2438, n2439, n2440, n2441, n2442, n2443, n2444;
  wire n2445, n2448, n2449, n2450, n2451, n2452, n2453, n2454;
  wire n2455, n2456, n2457, n2460, n2461, n2462, n2463, n2464;
  wire n2465, n2466, n2467, n2468, n2469, n2472, n2473, n2474;
  wire n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2484;
  wire n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492;
  wire n2493, n2496, n2497, n2498, n2499, n2500, n2501, n2502;
  wire n2503, n2504, n2505, n2508, n2509, n2510, n2511, n2512;
  wire n2513, n2514, n2515, n2516, n2517, n2520, n2521, n2522;
  wire n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2532;
  wire n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540;
  wire n2541, n2544, n2545, n2546, n2547, n2548, n2549, n2550;
  wire n2551, n2552, n2553, n2556, n2557, n2558, n2559, n2560;
  wire n2561, n2562, n2563, n2564, n2567, n2568, n2569, n2570;
  wire n2571, n2572, n2573, n2576, n2577, n2578, n2579, n2580;
  wire n2581, n2582, n2583, n2588, n2592, n2593, n2594, n2595;
  wire n2596, n2601, n2602, n2603, n2604, n2605, n2606, n2607;
  wire n2608, n2609, n2610, n2614, n2615, n2616, n2617, n2618;
  wire n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626;
  wire n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2636;
  wire n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644;
  wire n2645, n2648, n2649, n2650, n2651, n2652, n2653, n2654;
  wire n2655, n2656, n2657, n2660, n2661, n2662, n2663, n2664;
  wire n2665, n2666, n2667, n2668, n2669, n2672, n2673, n2674;
  wire n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2684;
  wire n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692;
  wire n2693, n2694, n2695, n2698, n2699, n2700, n2701, n2702;
  wire n2703, n2704, n2705, n2708, n2709, n2710, n2711, n2712;
  wire n2713, n2714, n2715, n2716, n2717, n2720, n2721, n2722;
  wire n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2732;
  wire n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740;
  wire n2741, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
  wire n2751, n2752, n2753, n2756, n2757, n2758, n2759, n2760;
  wire n2761, n2762, n2763, n2764, n2765, n2768, n2769, n2770;
  wire n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2780;
  wire n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788;
  wire n2789, n2792, n2793, n2794, n2795, n2796, n2797, n2798;
  wire n2799, n2800, n2801, n2804, n2805, n2806, n2807, n2808;
  wire n2809, n2810, n2811, n2812, n2815, n2816, n2817, n2818;
  wire n2819, n2820, n2821, n2824, n2825, n2826, n2827, n2828;
  wire n2829, n2830, n2831, n2836, n2840, n2841, n2842, n2843;
  wire n2844, n2849, n2850, n2851, n2852, n2853, n2854, n2855;
  wire n2856, n2857, n2858, n2862, n2863, n2864, n2865, n2866;
  wire n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874;
  wire n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2884;
  wire n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892;
  wire n2893, n2896, n2897, n2898, n2899, n2900, n2901, n2902;
  wire n2903, n2904, n2905, n2908, n2909, n2910, n2911, n2912;
  wire n2913, n2914, n2915, n2916, n2917, n2920, n2921, n2922;
  wire n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2932;
  wire n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940;
  wire n2941, n2944, n2945, n2946, n2947, n2948, n2949, n2950;
  wire n2951, n2952, n2953, n2956, n2957, n2958, n2959, n2960;
  wire n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2970;
  wire n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2980;
  wire n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988;
  wire n2989, n2992, n2993, n2994, n2995, n2996, n2997, n2998;
  wire n2999, n3000, n3001, n3004, n3005, n3006, n3007, n3008;
  wire n3009, n3010, n3011, n3012, n3013, n3016, n3017, n3018;
  wire n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3028;
  wire n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036;
  wire n3037, n3040, n3041, n3042, n3043, n3044, n3045, n3046;
  wire n3047, n3048, n3049, n3052, n3053, n3054, n3055, n3056;
  wire n3057, n3058, n3059, n3060, n3061, n3064, n3065, n3066;
  wire n3067, n3068, n3069, n3070, n3071, n3072, n3075, n3076;
  wire n3077, n3078, n3079, n3080, n3081, n3084, n3085, n3086;
  wire n3087, n3088, n3089, n3090, n3091, n3096, n3100, n3101;
  wire n3102, n3103, n3104, n3109, n3110, n3111, n3112, n3113;
  wire n3114, n3115, n3116, n3117, n3118, n3122, n3123, n3124;
  wire n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132;
  wire n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140;
  wire n3141, n3144, n3145, n3146, n3147, n3148, n3149, n3150;
  wire n3151, n3152, n3153, n3156, n3157, n3158, n3159, n3160;
  wire n3161, n3162, n3163, n3164, n3165, n3168, n3169, n3170;
  wire n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3180;
  wire n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188;
  wire n3189, n3192, n3193, n3194, n3195, n3196, n3197, n3198;
  wire n3199, n3200, n3201, n3204, n3205, n3206, n3207, n3208;
  wire n3209, n3210, n3211, n3212, n3213, n3216, n3217, n3218;
  wire n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3228;
  wire n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236;
  wire n3237, n3240, n3241, n3242, n3243, n3244, n3245, n3246;
  wire n3247, n3248, n3249, n3250, n3251, n3254, n3255, n3256;
  wire n3257, n3258, n3259, n3260, n3261, n3264, n3265, n3266;
  wire n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3276;
  wire n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284;
  wire n3285, n3288, n3289, n3290, n3291, n3292, n3293, n3294;
  wire n3295, n3296, n3297, n3300, n3301, n3302, n3303, n3304;
  wire n3305, n3306, n3307, n3308, n3309, n3312, n3313, n3314;
  wire n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3324;
  wire n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332;
  wire n3333, n3336, n3337, n3338, n3339, n3340, n3341, n3342;
  wire n3343, n3344, n3347, n3348, n3349, n3350, n3351, n3352;
  wire n3353, n3356, n3357, n3358, n3359, n3360, n3361, n3362;
  wire n3363, n3368, n3372, n3373, n3374, n3375, n3376, n3381;
  wire n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389;
  wire n3390, n3394, n3395, n3396, n3397, n3398, n3399, n3400;
  wire n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408;
  wire n3409, n3410, n3411, n3412, n3413, n3416, n3417, n3418;
  wire n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3428;
  wire n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436;
  wire n3437, n3440, n3441, n3442, n3443, n3444, n3445, n3446;
  wire n3447, n3448, n3449, n3452, n3453, n3454, n3455, n3456;
  wire n3457, n3458, n3459, n3460, n3461, n3464, n3465, n3466;
  wire n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3476;
  wire n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484;
  wire n3485, n3488, n3489, n3490, n3491, n3492, n3493, n3494;
  wire n3495, n3496, n3497, n3500, n3501, n3502, n3503, n3504;
  wire n3505, n3506, n3507, n3508, n3509, n3512, n3513, n3514;
  wire n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3524;
  wire n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532;
  wire n3533, n3536, n3537, n3538, n3539, n3540, n3541, n3542;
  wire n3543, n3544, n3545, n3546, n3547, n3550, n3551, n3552;
  wire n3553, n3554, n3555, n3556, n3557, n3560, n3561, n3562;
  wire n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3572;
  wire n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580;
  wire n3581, n3584, n3585, n3586, n3587, n3588, n3589, n3590;
  wire n3591, n3592, n3593, n3596, n3597, n3598, n3599, n3600;
  wire n3601, n3602, n3603, n3604, n3605, n3608, n3609, n3610;
  wire n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3620;
  wire n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628;
  wire n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3640;
  wire n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3652;
  wire n3656, n3657, n3658, n3659, n3660, n3665, n3666, n3667;
  wire n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3678;
  wire n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686;
  wire n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694;
  wire n3695, n3696, n3697, n3700, n3701, n3702, n3703, n3704;
  wire n3705, n3706, n3707, n3708, n3709, n3712, n3713, n3714;
  wire n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3724;
  wire n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732;
  wire n3733, n3736, n3737, n3738, n3739, n3740, n3741, n3742;
  wire n3743, n3744, n3745, n3748, n3749, n3750, n3751, n3752;
  wire n3753, n3754, n3755, n3756, n3757, n3760, n3761, n3762;
  wire n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3772;
  wire n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780;
  wire n3781, n3784, n3785, n3786, n3787, n3788, n3789, n3790;
  wire n3791, n3792, n3793, n3796, n3797, n3798, n3799, n3800;
  wire n3801, n3802, n3803, n3804, n3805, n3808, n3809, n3810;
  wire n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3820;
  wire n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828;
  wire n3829, n3832, n3833, n3834, n3835, n3836, n3837, n3838;
  wire n3839, n3840, n3841, n3844, n3845, n3846, n3847, n3848;
  wire n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3858;
  wire n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3868;
  wire n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876;
  wire n3877, n3880, n3881, n3882, n3883, n3884, n3885, n3886;
  wire n3887, n3888, n3889, n3892, n3893, n3894, n3895, n3896;
  wire n3897, n3898, n3899, n3900, n3901, n3904, n3905, n3906;
  wire n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3916;
  wire n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924;
  wire n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3936;
  wire n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3948;
  wire n3952, n3953, n3954, n3955, n3956, n3961, n3962, n3963;
  wire n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3974;
  wire n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982;
  wire n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990;
  wire n3991, n3992, n3993, n3996, n3997, n3998, n3999, n4000;
  wire n4001, n4002, n4003, n4004, n4005, n4008, n4009, n4010;
  wire n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4020;
  wire n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028;
  wire n4029, n4032, n4033, n4034, n4035, n4036, n4037, n4038;
  wire n4039, n4040, n4041, n4044, n4045, n4046, n4047, n4048;
  wire n4049, n4050, n4051, n4052, n4053, n4056, n4057, n4058;
  wire n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4068;
  wire n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076;
  wire n4077, n4080, n4081, n4082, n4083, n4084, n4085, n4086;
  wire n4087, n4088, n4089, n4092, n4093, n4094, n4095, n4096;
  wire n4097, n4098, n4099, n4100, n4101, n4104, n4105, n4106;
  wire n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4116;
  wire n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124;
  wire n4125, n4128, n4129, n4130, n4131, n4132, n4133, n4134;
  wire n4135, n4136, n4137, n4140, n4141, n4142, n4143, n4144;
  wire n4145, n4146, n4147, n4148, n4149, n4152, n4153, n4154;
  wire n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4164;
  wire n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172;
  wire n4173, n4174, n4175, n4178, n4179, n4180, n4181, n4182;
  wire n4183, n4184, n4185, n4188, n4189, n4190, n4191, n4192;
  wire n4193, n4194, n4195, n4196, n4197, n4200, n4201, n4202;
  wire n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4212;
  wire n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220;
  wire n4221, n4224, n4225, n4226, n4227, n4228, n4229, n4230;
  wire n4231, n4232, n4235, n4236, n4237, n4238, n4239, n4240;
  wire n4241, n4244, n4245, n4246, n4247, n4248, n4249, n4250;
  wire n4251, n4256, n4260, n4261, n4262, n4263, n4264, n4269;
  wire n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277;
  wire n4278, n4282, n4283, n4284, n4285, n4286, n4287, n4288;
  wire n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296;
  wire n4297, n4298, n4299, n4300, n4301, n4304, n4305, n4306;
  wire n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4316;
  wire n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324;
  wire n4325, n4328, n4329, n4330, n4331, n4332, n4333, n4334;
  wire n4335, n4336, n4337, n4340, n4341, n4342, n4343, n4344;
  wire n4345, n4346, n4347, n4348, n4349, n4352, n4353, n4354;
  wire n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4364;
  wire n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372;
  wire n4373, n4376, n4377, n4378, n4379, n4380, n4381, n4382;
  wire n4383, n4384, n4385, n4388, n4389, n4390, n4391, n4392;
  wire n4393, n4394, n4395, n4396, n4397, n4400, n4401, n4402;
  wire n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4412;
  wire n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420;
  wire n4421, n4424, n4425, n4426, n4427, n4428, n4429, n4430;
  wire n4431, n4432, n4433, n4436, n4437, n4438, n4439, n4440;
  wire n4441, n4442, n4443, n4444, n4445, n4448, n4449, n4450;
  wire n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4460;
  wire n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468;
  wire n4469, n4472, n4473, n4474, n4475, n4476, n4477, n4478;
  wire n4479, n4480, n4481, n4484, n4485, n4486, n4487, n4488;
  wire n4489, n4490, n4491, n4492, n4493, n4496, n4497, n4498;
  wire n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506;
  wire n4507, n4510, n4511, n4512, n4513, n4514, n4515, n4516;
  wire n4517, n4520, n4521, n4522, n4523, n4524, n4525, n4526;
  wire n4527, n4528, n4529, n4532, n4533, n4534, n4535, n4536;
  wire n4537, n4538, n4539, n4540, n4541, n4544, n4545, n4546;
  wire n4547, n4548, n4549, n4550, n4551, n4552, n4555, n4556;
  wire n4557, n4558, n4559, n4560, n4561, n4564, n4565, n4566;
  wire n4567, n4568, n4569, n4570, n4571, n4576, n4580, n4581;
  wire n4582, n4583, n4584, n4589, n4590, n4591, n4592, n4593;
  wire n4594, n4595, n4596, n4597, n4598, n4602, n4603, n4604;
  wire n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612;
  wire n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620;
  wire n4621, n4624, n4625, n4626, n4627, n4628, n4629, n4630;
  wire n4631, n4632, n4633, n4636, n4637, n4638, n4639, n4640;
  wire n4641, n4642, n4643, n4644, n4645, n4648, n4649, n4650;
  wire n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4660;
  wire n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668;
  wire n4669, n4672, n4673, n4674, n4675, n4676, n4677, n4678;
  wire n4679, n4680, n4681, n4684, n4685, n4686, n4687, n4688;
  wire n4689, n4690, n4691, n4692, n4693, n4696, n4697, n4698;
  wire n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4708;
  wire n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716;
  wire n4717, n4720, n4721, n4722, n4723, n4724, n4725, n4726;
  wire n4727, n4728, n4729, n4732, n4733, n4734, n4735, n4736;
  wire n4737, n4738, n4739, n4740, n4741, n4744, n4745, n4746;
  wire n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4756;
  wire n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764;
  wire n4765, n4768, n4769, n4770, n4771, n4772, n4773, n4774;
  wire n4775, n4776, n4777, n4780, n4781, n4782, n4783, n4784;
  wire n4785, n4786, n4787, n4788, n4789, n4792, n4793, n4794;
  wire n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4804;
  wire n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812;
  wire n4813, n4816, n4817, n4818, n4819, n4820, n4821, n4822;
  wire n4823, n4824, n4825, n4828, n4829, n4830, n4831, n4832;
  wire n4833, n4834, n4835, n4836, n4837, n4840, n4841, n4842;
  wire n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850;
  wire n4851, n4854, n4855, n4856, n4857, n4858, n4859, n4860;
  wire n4861, n4864, n4865, n4866, n4867, n4868, n4869, n4870;
  wire n4871, n4872, n4873, n4876, n4877, n4878, n4879, n4880;
  wire n4881, n4882, n4883, n4884, n4887, n4888, n4889, n4890;
  wire n4891, n4892, n4893, n4896, n4897, n4898, n4899, n4900;
  wire n4901, n4902, n4903, n4908, n4912, n4913, n4914, n4915;
  wire n4916, n4921, n4922, n4923, n4924, n4925, n4926, n4927;
  wire n4928, n4929, n4930, n4934, n4935, n4936, n4937, n4938;
  wire n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946;
  wire n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4956;
  wire n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964;
  wire n4965, n4968, n4969, n4970, n4971, n4972, n4973, n4974;
  wire n4975, n4976, n4977, n4980, n4981, n4982, n4983, n4984;
  wire n4985, n4986, n4987, n4988, n4989, n4992, n4993, n4994;
  wire n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5004;
  wire n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012;
  wire n5013, n5016, n5017, n5018, n5019, n5020, n5021, n5022;
  wire n5023, n5024, n5025, n5028, n5029, n5030, n5031, n5032;
  wire n5033, n5034, n5035, n5036, n5037, n5040, n5041, n5042;
  wire n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5052;
  wire n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060;
  wire n5061, n5064, n5065, n5066, n5067, n5068, n5069, n5070;
  wire n5071, n5072, n5073, n5076, n5077, n5078, n5079, n5080;
  wire n5081, n5082, n5083, n5084, n5085, n5088, n5089, n5090;
  wire n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5100;
  wire n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108;
  wire n5109, n5112, n5113, n5114, n5115, n5116, n5117, n5118;
  wire n5119, n5120, n5121, n5124, n5125, n5126, n5127, n5128;
  wire n5129, n5130, n5131, n5132, n5133, n5136, n5137, n5138;
  wire n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5148;
  wire n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156;
  wire n5157, n5160, n5161, n5162, n5163, n5164, n5165, n5166;
  wire n5167, n5168, n5169, n5172, n5173, n5174, n5175, n5176;
  wire n5177, n5178, n5179, n5180, n5181, n5184, n5185, n5186;
  wire n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5196;
  wire n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204;
  wire n5205, n5206, n5207, n5210, n5211, n5212, n5213, n5214;
  wire n5215, n5216, n5217, n5220, n5221, n5222, n5223, n5224;
  wire n5225, n5226, n5227, n5228, n5231, n5232, n5233, n5234;
  wire n5235, n5236, n5237, n5240, n5241, n5242, n5243, n5244;
  wire n5245, n5246, n5247, n5252, n5256, n5257, n5258, n5259;
  wire n5260, n5265, n5266, n5267, n5268, n5269, n5270, n5271;
  wire n5272, n5273, n5274, n5278, n5279, n5280, n5281, n5282;
  wire n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290;
  wire n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5300;
  wire n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308;
  wire n5309, n5312, n5313, n5314, n5315, n5316, n5317, n5318;
  wire n5319, n5320, n5321, n5324, n5325, n5326, n5327, n5328;
  wire n5329, n5330, n5331, n5332, n5333, n5336, n5337, n5338;
  wire n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5348;
  wire n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356;
  wire n5357, n5360, n5361, n5362, n5363, n5364, n5365, n5366;
  wire n5367, n5368, n5369, n5372, n5373, n5374, n5375, n5376;
  wire n5377, n5378, n5379, n5380, n5381, n5384, n5385, n5386;
  wire n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5396;
  wire n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404;
  wire n5405, n5408, n5409, n5410, n5411, n5412, n5413, n5414;
  wire n5415, n5416, n5417, n5420, n5421, n5422, n5423, n5424;
  wire n5425, n5426, n5427, n5428, n5429, n5432, n5433, n5434;
  wire n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5444;
  wire n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452;
  wire n5453, n5456, n5457, n5458, n5459, n5460, n5461, n5462;
  wire n5463, n5464, n5465, n5468, n5469, n5470, n5471, n5472;
  wire n5473, n5474, n5475, n5476, n5477, n5480, n5481, n5482;
  wire n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5492;
  wire n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500;
  wire n5501, n5504, n5505, n5506, n5507, n5508, n5509, n5510;
  wire n5511, n5512, n5513, n5516, n5517, n5518, n5519, n5520;
  wire n5521, n5522, n5523, n5524, n5525, n5528, n5529, n5530;
  wire n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5540;
  wire n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548;
  wire n5549, n5552, n5553, n5554, n5555, n5556, n5557, n5558;
  wire n5559, n5560, n5561, n5564, n5565, n5566, n5567, n5568;
  wire n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5578;
  wire n5579, n5580, n5581, n5582, n5583, n5584, n5587, n5588;
  wire n5589, n5590, n5591, n5592, n5593, n5596, n5597, n5598;
  wire n5599, n5600, n5601, n5602, n5603, n5608, n5612, n5613;
  wire n5614, n5615, n5616, n5621, n5622, n5623, n5624, n5625;
  wire n5626, n5627, n5628, n5629, n5630, n5634, n5635, n5636;
  wire n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644;
  wire n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652;
  wire n5653, n5656, n5657, n5658, n5659, n5660, n5661, n5662;
  wire n5663, n5664, n5665, n5668, n5669, n5670, n5671, n5672;
  wire n5673, n5674, n5675, n5676, n5677, n5680, n5681, n5682;
  wire n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5692;
  wire n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700;
  wire n5701, n5704, n5705, n5706, n5707, n5708, n5709, n5710;
  wire n5711, n5712, n5713, n5716, n5717, n5718, n5719, n5720;
  wire n5721, n5722, n5723, n5724, n5725, n5728, n5729, n5730;
  wire n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5740;
  wire n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748;
  wire n5749, n5752, n5753, n5754, n5755, n5756, n5757, n5758;
  wire n5759, n5760, n5761, n5764, n5765, n5766, n5767, n5768;
  wire n5769, n5770, n5771, n5772, n5773, n5776, n5777, n5778;
  wire n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5788;
  wire n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796;
  wire n5797, n5800, n5801, n5802, n5803, n5804, n5805, n5806;
  wire n5807, n5808, n5809, n5812, n5813, n5814, n5815, n5816;
  wire n5817, n5818, n5819, n5820, n5821, n5824, n5825, n5826;
  wire n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5836;
  wire n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844;
  wire n5845, n5848, n5849, n5850, n5851, n5852, n5853, n5854;
  wire n5855, n5856, n5857, n5860, n5861, n5862, n5863, n5864;
  wire n5865, n5866, n5867, n5868, n5869, n5872, n5873, n5874;
  wire n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5884;
  wire n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892;
  wire n5893, n5896, n5897, n5898, n5899, n5900, n5901, n5902;
  wire n5903, n5904, n5905, n5908, n5909, n5910, n5911, n5912;
  wire n5913, n5914, n5915, n5916, n5917, n5920, n5921, n5922;
  wire n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5932;
  wire n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940;
  wire n5941, n5944, n5945, n5946, n5947, n5948, n5949, n5950;
  wire n5951, n5952, n5955, n5956, n5957, n5958, n5959, n5960;
  wire n5961, n5964, n5965, n5966, n5967, n5968, n5969, n5970;
  wire n5971, n5976, n5980, n5981, n5982, n5983, n5984, n5989;
  wire n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997;
  wire n5998, n6002, n6003, n6004, n6005, n6006, n6007, n6008;
  wire n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016;
  wire n6017, n6018, n6019, n6020, n6021, n6024, n6025, n6026;
  wire n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6036;
  wire n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044;
  wire n6045, n6048, n6049, n6050, n6051, n6052, n6053, n6054;
  wire n6055, n6056, n6057, n6060, n6061, n6062, n6063, n6064;
  wire n6065, n6066, n6067, n6068, n6069, n6072, n6073, n6074;
  wire n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6084;
  wire n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092;
  wire n6093, n6096, n6097, n6098, n6099, n6100, n6101, n6102;
  wire n6103, n6104, n6105, n6108, n6109, n6110, n6111, n6112;
  wire n6113, n6114, n6115, n6116, n6117, n6120, n6121, n6122;
  wire n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6132;
  wire n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140;
  wire n6141, n6144, n6145, n6146, n6147, n6148, n6149, n6150;
  wire n6151, n6152, n6153, n6156, n6157, n6158, n6159, n6160;
  wire n6161, n6162, n6163, n6164, n6165, n6168, n6169, n6170;
  wire n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6180;
  wire n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188;
  wire n6189, n6192, n6193, n6194, n6195, n6196, n6197, n6198;
  wire n6199, n6200, n6201, n6204, n6205, n6206, n6207, n6208;
  wire n6209, n6210, n6211, n6212, n6213, n6216, n6217, n6218;
  wire n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6228;
  wire n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236;
  wire n6237, n6240, n6241, n6242, n6243, n6244, n6245, n6246;
  wire n6247, n6248, n6249, n6252, n6253, n6254, n6255, n6256;
  wire n6257, n6258, n6259, n6260, n6261, n6264, n6265, n6266;
  wire n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6276;
  wire n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284;
  wire n6285, n6288, n6289, n6290, n6291, n6292, n6293, n6294;
  wire n6295, n6296, n6297, n6300, n6301, n6302, n6303, n6304;
  wire n6305, n6306, n6307, n6308, n6309, n6312, n6313, n6314;
  wire n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6324;
  wire n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332;
  wire n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6344;
  wire n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6356;
  wire n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367;
  wire n6368, n6373, n6374, n6375, n6376, n6377, n6378, n6382;
  wire n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390;
  wire n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398;
  wire n6399, n6400, n6401, n6404, n6405, n6406, n6407, n6408;
  wire n6409, n6410, n6411, n6412, n6413, n6416, n6417, n6418;
  wire n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6428;
  wire n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436;
  wire n6437, n6440, n6441, n6442, n6443, n6444, n6445, n6446;
  wire n6447, n6448, n6449, n6452, n6453, n6454, n6455, n6456;
  wire n6457, n6458, n6459, n6460, n6461, n6464, n6465, n6466;
  wire n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6476;
  wire n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484;
  wire n6485, n6488, n6489, n6490, n6491, n6492, n6493, n6494;
  wire n6495, n6496, n6497, n6500, n6501, n6502, n6503, n6504;
  wire n6505, n6506, n6507, n6508, n6509, n6512, n6513, n6514;
  wire n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6524;
  wire n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532;
  wire n6533, n6536, n6537, n6538, n6539, n6540, n6541, n6542;
  wire n6543, n6544, n6545, n6548, n6549, n6550, n6551, n6552;
  wire n6553, n6554, n6555, n6556, n6557, n6560, n6561, n6562;
  wire n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6572;
  wire n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580;
  wire n6581, n6584, n6585, n6586, n6587, n6588, n6589, n6590;
  wire n6591, n6592, n6593, n6596, n6597, n6598, n6599, n6600;
  wire n6601, n6602, n6603, n6604, n6605, n6608, n6609, n6610;
  wire n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6620;
  wire n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628;
  wire n6629, n6632, n6633, n6634, n6635, n6636, n6637, n6638;
  wire n6639, n6640, n6641, n6644, n6645, n6646, n6647, n6648;
  wire n6649, n6650, n6651, n6652, n6653, n6656, n6657, n6658;
  wire n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6668;
  wire n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676;
  wire n6677, n6680, n6681, n6682, n6683, n6684, n6685, n6686;
  wire n6687, n6688, n6689, n6692, n6693, n6694, n6695, n6696;
  wire n6697, n6698, n6699, n6700, n6701, n6704, n6705, n6706;
  wire n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6716;
  wire n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724;
  wire n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6736;
  wire n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6748;
  wire n6752, n6753, n6754, n6755, n6756, n6761, n6762, n6763;
  wire n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6774;
  wire n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782;
  wire n6783, n6784, n6787, n6788, n6789, n6790, n6791, n6792;
  wire n6793, n6794, n6797, n6798, n6799, n6800, n6801, n6802;
  wire n6803, n6804, n6805, n6806, n6809, n6810, n6811, n6812;
  wire n6813, n6814, n6815, n6816, n6817, n6818, n6821, n6822;
  wire n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830;
  wire n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840;
  wire n6841, n6842, n6845, n6846, n6847, n6848, n6849, n6850;
  wire n6851, n6852, n6853, n6854, n6857, n6858, n6859, n6860;
  wire n6861, n6862, n6863, n6864, n6865, n6866, n6869, n6870;
  wire n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878;
  wire n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888;
  wire n6889, n6890, n6893, n6894, n6895, n6896, n6897, n6898;
  wire n6899, n6900, n6901, n6902, n6905, n6906, n6907, n6908;
  wire n6909, n6910, n6911, n6912, n6913, n6914, n6917, n6918;
  wire n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926;
  wire n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936;
  wire n6937, n6938, n6941, n6942, n6943, n6944, n6945, n6946;
  wire n6947, n6948, n6949, n6950, n6953, n6954, n6955, n6956;
  wire n6957, n6958, n6959, n6960, n6961, n6962, n6965, n6966;
  wire n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974;
  wire n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984;
  wire n6985, n6986, n6989, n6990, n6991, n6992, n6993, n6994;
  wire n6995, n6996, n6997, n6998, n7001, n7002, n7003, n7004;
  wire n7005, n7006, n7007, n7008, n7009, n7010, n7013, n7014;
  wire n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022;
  wire n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032;
  wire n7033, n7034, n7037, n7038, n7039, n7040, n7041, n7042;
  wire n7043, n7044, n7045, n7046, n7049, n7050, n7051, n7052;
  wire n7053, n7054, n7055, n7056, n7057, n7058, n7061, n7062;
  wire n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070;
  wire n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080;
  wire n7081, n7082, n7085, n7086, n7087, n7088, n7089, n7090;
  wire n7091, n7092, n7093, n7094, n7097, n7098, n7099, n7100;
  wire n7101, n7102, n7103, n7104, n7105, n7106, n7109, n7110;
  wire n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118;
  wire n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128;
  wire n7129, n7132, n7133, n7134, n7135, n7136, n7137, n7138;
  wire n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148;
  wire n7153, n7157, n7158, n7159, n7160, n7161, n7166, n7167;
  wire n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175;
  wire n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186;
  wire n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194;
  wire n7195, n7196, n7197, n7198, n7201, n7202, n7203, n7204;
  wire n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212;
  wire n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222;
  wire n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232;
  wire n7233, n7234, n7237, n7238, n7239, n7240, n7241, n7242;
  wire n7243, n7244, n7245, n7246, n7249, n7250, n7251, n7252;
  wire n7253, n7254, n7255, n7256, n7257, n7258, n7261, n7262;
  wire n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270;
  wire n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280;
  wire n7281, n7282, n7285, n7286, n7287, n7288, n7289, n7290;
  wire n7291, n7292, n7293, n7294, n7297, n7298, n7299, n7300;
  wire n7301, n7302, n7303, n7304, n7305, n7306, n7309, n7310;
  wire n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318;
  wire n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328;
  wire n7329, n7330, n7333, n7334, n7335, n7336, n7337, n7338;
  wire n7339, n7340, n7341, n7342, n7345, n7346, n7347, n7348;
  wire n7349, n7350, n7351, n7352, n7353, n7354, n7357, n7358;
  wire n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366;
  wire n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376;
  wire n7377, n7378, n7381, n7382, n7383, n7384, n7385, n7386;
  wire n7387, n7388, n7389, n7390, n7393, n7394, n7395, n7396;
  wire n7397, n7398, n7399, n7400, n7401, n7402, n7405, n7406;
  wire n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414;
  wire n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424;
  wire n7425, n7426, n7429, n7430, n7431, n7432, n7433, n7434;
  wire n7435, n7436, n7437, n7438, n7441, n7442, n7443, n7444;
  wire n7445, n7446, n7447, n7448, n7449, n7450, n7453, n7454;
  wire n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462;
  wire n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472;
  wire n7473, n7474, n7477, n7478, n7479, n7480, n7481, n7482;
  wire n7483, n7484, n7485, n7486, n7489, n7490, n7491, n7492;
  wire n7493, n7494, n7495, n7496, n7497, n7498, n7501, n7502;
  wire n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510;
  wire n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520;
  wire n7521, n7522, n7525, n7526, n7527, n7528, n7529, n7530;
  wire n7531, n7532, n7533, n7534, n7537, n7538, n7539, n7540;
  wire n7541, n7542, n7543, n7544, n7545, n7548, n7549, n7550;
  wire n7551, n7552, n7553, n7554, n7557, n7558, n7559, n7560;
  wire n7561, n7562, n7563, n7564, n7569, n7573, n7574, n7575;
  wire n7576, n7577, n7582, n7583, n7584, n7585, n7586, n7587;
  wire n7588, n7589, n7590, n7591, n7595, n7596, n7597, n7598;
  wire n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606;
  wire n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614;
  wire n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624;
  wire n7625, n7626, n7629, n7630, n7631, n7632, n7633, n7634;
  wire n7635, n7636, n7637, n7638, n7641, n7642, n7643, n7644;
  wire n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652;
  wire n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662;
  wire n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672;
  wire n7673, n7674, n7677, n7678, n7679, n7680, n7681, n7682;
  wire n7683, n7684, n7685, n7686, n7689, n7690, n7691, n7692;
  wire n7693, n7694, n7695, n7696, n7697, n7698, n7701, n7702;
  wire n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710;
  wire n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720;
  wire n7721, n7722, n7725, n7726, n7727, n7728, n7729, n7730;
  wire n7731, n7732, n7733, n7734, n7737, n7738, n7739, n7740;
  wire n7741, n7742, n7743, n7744, n7745, n7746, n7749, n7750;
  wire n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758;
  wire n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768;
  wire n7769, n7770, n7773, n7774, n7775, n7776, n7777, n7778;
  wire n7779, n7780, n7781, n7782, n7785, n7786, n7787, n7788;
  wire n7789, n7790, n7791, n7792, n7793, n7794, n7797, n7798;
  wire n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806;
  wire n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816;
  wire n7817, n7818, n7821, n7822, n7823, n7824, n7825, n7826;
  wire n7827, n7828, n7829, n7830, n7833, n7834, n7835, n7836;
  wire n7837, n7838, n7839, n7840, n7841, n7842, n7845, n7846;
  wire n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854;
  wire n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864;
  wire n7865, n7866, n7869, n7870, n7871, n7872, n7873, n7874;
  wire n7875, n7876, n7877, n7878, n7881, n7882, n7883, n7884;
  wire n7885, n7886, n7887, n7888, n7889, n7890, n7893, n7894;
  wire n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902;
  wire n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912;
  wire n7913, n7914, n7917, n7918, n7919, n7920, n7921, n7922;
  wire n7923, n7924, n7925, n7926, n7929, n7930, n7931, n7932;
  wire n7933, n7934, n7935, n7936, n7937, n7938, n7941, n7942;
  wire n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950;
  wire n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960;
  wire n7961, n7962, n7965, n7966, n7967, n7968, n7969, n7970;
  wire n7971, n7972, n7973, n7976, n7977, n7978, n7979, n7980;
  wire n7981, n7982, n7985, n7986, n7987, n7988, n7989, n7990;
  wire n7991, n7992, n7997, n8001, n8002, n8003, n8004, n8005;
  wire n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017;
  wire n8018, n8019, n8023, n8024, n8025, n8026, n8027, n8028;
  wire n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036;
  wire n8037, n8038, n8039, n8040, n8041, n8042, n8045, n8046;
  wire n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054;
  wire n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064;
  wire n8065, n8066, n8069, n8070, n8071, n8072, n8073, n8074;
  wire n8075, n8076, n8077, n8078, n8081, n8082, n8083, n8084;
  wire n8085, n8086, n8087, n8088, n8089, n8090, n8093, n8094;
  wire n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102;
  wire n8103, n8104, n8107, n8108, n8109, n8110, n8111, n8112;
  wire n8113, n8114, n8117, n8118, n8119, n8120, n8121, n8122;
  wire n8123, n8124, n8125, n8126, n8129, n8130, n8131, n8132;
  wire n8133, n8134, n8135, n8136, n8137, n8138, n8141, n8142;
  wire n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150;
  wire n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160;
  wire n8161, n8162, n8165, n8166, n8167, n8168, n8169, n8170;
  wire n8171, n8172, n8173, n8174, n8177, n8178, n8179, n8180;
  wire n8181, n8182, n8183, n8184, n8185, n8186, n8189, n8190;
  wire n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198;
  wire n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208;
  wire n8209, n8210, n8213, n8214, n8215, n8216, n8217, n8218;
  wire n8219, n8220, n8221, n8222, n8225, n8226, n8227, n8228;
  wire n8229, n8230, n8231, n8232, n8233, n8234, n8237, n8238;
  wire n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246;
  wire n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256;
  wire n8257, n8258, n8261, n8262, n8263, n8264, n8265, n8266;
  wire n8267, n8268, n8269, n8270, n8273, n8274, n8275, n8276;
  wire n8277, n8278, n8279, n8280, n8281, n8282, n8285, n8286;
  wire n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294;
  wire n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304;
  wire n8305, n8306, n8309, n8310, n8311, n8312, n8313, n8314;
  wire n8315, n8316, n8317, n8318, n8321, n8322, n8323, n8324;
  wire n8325, n8326, n8327, n8328, n8329, n8330, n8333, n8334;
  wire n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342;
  wire n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352;
  wire n8353, n8354, n8357, n8358, n8359, n8360, n8361, n8362;
  wire n8363, n8364, n8365, n8366, n8369, n8370, n8371, n8372;
  wire n8373, n8374, n8375, n8376, n8377, n8378, n8381, n8382;
  wire n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390;
  wire n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400;
  wire n8401, n8402, n8405, n8406, n8407, n8408, n8409, n8410;
  wire n8411, n8412, n8413, n8416, n8417, n8418, n8419, n8420;
  wire n8421, n8422, n8425, n8426, n8427, n8428, n8429, n8430;
  wire n8431, n8432, n8437, n8441, n8442, n8443, n8444, n8445;
  wire n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457;
  wire n8458, n8459, n8463, n8464, n8465, n8466, n8467, n8468;
  wire n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476;
  wire n8477, n8478, n8479, n8480, n8481, n8482, n8485, n8486;
  wire n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494;
  wire n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504;
  wire n8505, n8506, n8509, n8510, n8511, n8512, n8513, n8514;
  wire n8515, n8516, n8517, n8518, n8521, n8522, n8523, n8524;
  wire n8525, n8526, n8527, n8528, n8529, n8530, n8533, n8534;
  wire n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542;
  wire n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552;
  wire n8553, n8554, n8557, n8558, n8559, n8560, n8561, n8562;
  wire n8563, n8564, n8565, n8566, n8567, n8568, n8571, n8572;
  wire n8573, n8574, n8575, n8576, n8577, n8578, n8581, n8582;
  wire n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590;
  wire n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600;
  wire n8601, n8602, n8605, n8606, n8607, n8608, n8609, n8610;
  wire n8611, n8612, n8613, n8614, n8617, n8618, n8619, n8620;
  wire n8621, n8622, n8623, n8624, n8625, n8626, n8629, n8630;
  wire n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638;
  wire n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648;
  wire n8649, n8650, n8653, n8654, n8655, n8656, n8657, n8658;
  wire n8659, n8660, n8661, n8662, n8665, n8666, n8667, n8668;
  wire n8669, n8670, n8671, n8672, n8673, n8674, n8677, n8678;
  wire n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686;
  wire n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696;
  wire n8697, n8698, n8701, n8702, n8703, n8704, n8705, n8706;
  wire n8707, n8708, n8709, n8710, n8713, n8714, n8715, n8716;
  wire n8717, n8718, n8719, n8720, n8721, n8722, n8725, n8726;
  wire n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734;
  wire n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744;
  wire n8745, n8746, n8749, n8750, n8751, n8752, n8753, n8754;
  wire n8755, n8756, n8757, n8758, n8761, n8762, n8763, n8764;
  wire n8765, n8766, n8767, n8768, n8769, n8770, n8773, n8774;
  wire n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782;
  wire n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792;
  wire n8793, n8794, n8797, n8798, n8799, n8800, n8801, n8802;
  wire n8803, n8804, n8805, n8806, n8809, n8810, n8811, n8812;
  wire n8813, n8814, n8815, n8816, n8817, n8818, n8821, n8822;
  wire n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830;
  wire n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840;
  wire n8841, n8842, n8845, n8846, n8847, n8848, n8849, n8850;
  wire n8851, n8852, n8853, n8854, n8857, n8858, n8859, n8860;
  wire n8861, n8862, n8863, n8864, n8865, n8868, n8869, n8870;
  wire n8871, n8872, n8873, n8874, n8877, n8878, n8879, n8880;
  wire n8881, n8882, n8883, n8884, n8889, n8893, n8894, n8895;
  wire n8896, n8897, n8902, n8903, n8904, n8905, n8906, n8907;
  wire n8908, n8909, n8910, n8911, n8915, n8916, n8917, n8918;
  wire n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926;
  wire n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934;
  wire n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944;
  wire n8945, n8946, n8949, n8950, n8951, n8952, n8953, n8954;
  wire n8955, n8956, n8957, n8958, n8961, n8962, n8963, n8964;
  wire n8965, n8966, n8967, n8968, n8969, n8970, n8973, n8974;
  wire n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982;
  wire n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992;
  wire n8993, n8994, n8997, n8998, n8999, n9000, n9001, n9002;
  wire n9003, n9004, n9005, n9006, n9009, n9010, n9011, n9012;
  wire n9013, n9014, n9015, n9016, n9017, n9018, n9021, n9022;
  wire n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030;
  wire n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040;
  wire n9041, n9042, n9043, n9044, n9047, n9048, n9049, n9050;
  wire n9051, n9052, n9053, n9054, n9057, n9058, n9059, n9060;
  wire n9061, n9062, n9063, n9064, n9065, n9066, n9069, n9070;
  wire n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078;
  wire n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088;
  wire n9089, n9090, n9093, n9094, n9095, n9096, n9097, n9098;
  wire n9099, n9100, n9101, n9102, n9105, n9106, n9107, n9108;
  wire n9109, n9110, n9111, n9112, n9113, n9114, n9117, n9118;
  wire n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126;
  wire n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136;
  wire n9137, n9138, n9141, n9142, n9143, n9144, n9145, n9146;
  wire n9147, n9148, n9149, n9150, n9153, n9154, n9155, n9156;
  wire n9157, n9158, n9159, n9160, n9161, n9162, n9165, n9166;
  wire n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174;
  wire n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184;
  wire n9185, n9186, n9189, n9190, n9191, n9192, n9193, n9194;
  wire n9195, n9196, n9197, n9198, n9201, n9202, n9203, n9204;
  wire n9205, n9206, n9207, n9208, n9209, n9210, n9213, n9214;
  wire n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222;
  wire n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232;
  wire n9233, n9234, n9237, n9238, n9239, n9240, n9241, n9242;
  wire n9243, n9244, n9245, n9246, n9249, n9250, n9251, n9252;
  wire n9253, n9254, n9255, n9256, n9257, n9258, n9261, n9262;
  wire n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270;
  wire n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280;
  wire n9281, n9282, n9285, n9286, n9287, n9288, n9289, n9290;
  wire n9291, n9292, n9293, n9294, n9297, n9298, n9299, n9300;
  wire n9301, n9302, n9303, n9304, n9305, n9306, n9309, n9310;
  wire n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318;
  wire n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328;
  wire n9329, n9332, n9333, n9334, n9335, n9336, n9337, n9338;
  wire n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348;
  wire n9353, n9357, n9358, n9359, n9360, n9361, n9366, n9367;
  wire n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375;
  wire n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386;
  wire n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394;
  wire n9395, n9396, n9397, n9398, n9401, n9402, n9403, n9404;
  wire n9405, n9406, n9407, n9408, n9409, n9410, n9413, n9414;
  wire n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422;
  wire n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432;
  wire n9433, n9434, n9437, n9438, n9439, n9440, n9441, n9442;
  wire n9443, n9444, n9445, n9446, n9449, n9450, n9451, n9452;
  wire n9453, n9454, n9455, n9456, n9457, n9458, n9461, n9462;
  wire n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470;
  wire n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480;
  wire n9481, n9482, n9485, n9486, n9487, n9488, n9489, n9490;
  wire n9491, n9492, n9493, n9494, n9497, n9498, n9499, n9500;
  wire n9501, n9502, n9503, n9504, n9505, n9506, n9509, n9510;
  wire n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518;
  wire n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528;
  wire n9529, n9530, n9531, n9532, n9535, n9536, n9537, n9538;
  wire n9539, n9540, n9541, n9542, n9545, n9546, n9547, n9548;
  wire n9549, n9550, n9551, n9552, n9553, n9554, n9557, n9558;
  wire n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566;
  wire n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576;
  wire n9577, n9578, n9581, n9582, n9583, n9584, n9585, n9586;
  wire n9587, n9588, n9589, n9590, n9593, n9594, n9595, n9596;
  wire n9597, n9598, n9599, n9600, n9601, n9602, n9605, n9606;
  wire n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614;
  wire n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624;
  wire n9625, n9626, n9629, n9630, n9631, n9632, n9633, n9634;
  wire n9635, n9636, n9637, n9638, n9641, n9642, n9643, n9644;
  wire n9645, n9646, n9647, n9648, n9649, n9650, n9653, n9654;
  wire n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662;
  wire n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672;
  wire n9673, n9674, n9677, n9678, n9679, n9680, n9681, n9682;
  wire n9683, n9684, n9685, n9686, n9689, n9690, n9691, n9692;
  wire n9693, n9694, n9695, n9696, n9697, n9698, n9701, n9702;
  wire n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710;
  wire n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720;
  wire n9721, n9722, n9725, n9726, n9727, n9728, n9729, n9730;
  wire n9731, n9732, n9733, n9734, n9737, n9738, n9739, n9740;
  wire n9741, n9742, n9743, n9744, n9745, n9746, n9749, n9750;
  wire n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758;
  wire n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768;
  wire n9769, n9770, n9773, n9774, n9775, n9776, n9777, n9778;
  wire n9779, n9780, n9781, n9782, n9785, n9786, n9787, n9788;
  wire n9789, n9790, n9791, n9792, n9793, n9794, n9797, n9798;
  wire n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9808;
  wire n9809, n9810, n9811, n9812, n9813, n9814, n9817, n9818;
  wire n9819, n9820, n9821, n9822, n9823, n9824, n9829, n9833;
  wire n9834, n9835, n9836, n9837, n9842, n9843, n9844, n9845;
  wire n9846, n9847, n9848, n9849, n9850, n9851, n9855, n9856;
  wire n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864;
  wire n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872;
  wire n9873, n9874, n9877, n9878, n9879, n9880, n9881, n9882;
  wire n9883, n9884, n9885, n9886, n9889, n9890, n9891, n9892;
  wire n9893, n9894, n9895, n9896, n9897, n9898, n9901, n9902;
  wire n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910;
  wire n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920;
  wire n9921, n9922, n9925, n9926, n9927, n9928, n9929, n9930;
  wire n9931, n9932, n9933, n9934, n9937, n9938, n9939, n9940;
  wire n9941, n9942, n9943, n9944, n9945, n9946, n9949, n9950;
  wire n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958;
  wire n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968;
  wire n9969, n9970, n9973, n9974, n9975, n9976, n9977, n9978;
  wire n9979, n9980, n9981, n9982, n9985, n9986, n9987, n9988;
  wire n9989, n9990, n9991, n9992, n9993, n9994, n9997, n9998;
  wire n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006;
  wire n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016;
  wire n10017, n10018, n10021, n10022, n10023, n10024, n10025, n10026;
  wire n10027, n10028, n10029, n10030, n10031, n10032, n10035, n10036;
  wire n10037, n10038, n10039, n10040, n10041, n10042, n10045, n10046;
  wire n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054;
  wire n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064;
  wire n10065, n10066, n10069, n10070, n10071, n10072, n10073, n10074;
  wire n10075, n10076, n10077, n10078, n10081, n10082, n10083, n10084;
  wire n10085, n10086, n10087, n10088, n10089, n10090, n10093, n10094;
  wire n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102;
  wire n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112;
  wire n10113, n10114, n10117, n10118, n10119, n10120, n10121, n10122;
  wire n10123, n10124, n10125, n10126, n10129, n10130, n10131, n10132;
  wire n10133, n10134, n10135, n10136, n10137, n10138, n10141, n10142;
  wire n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150;
  wire n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160;
  wire n10161, n10162, n10165, n10166, n10167, n10168, n10169, n10170;
  wire n10171, n10172, n10173, n10174, n10177, n10178, n10179, n10180;
  wire n10181, n10182, n10183, n10184, n10185, n10186, n10189, n10190;
  wire n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198;
  wire n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208;
  wire n10209, n10210, n10213, n10214, n10215, n10216, n10217, n10218;
  wire n10219, n10220, n10221, n10222, n10225, n10226, n10227, n10228;
  wire n10229, n10230, n10231, n10232, n10233, n10234, n10237, n10238;
  wire n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246;
  wire n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256;
  wire n10257, n10258, n10261, n10262, n10263, n10264, n10265, n10266;
  wire n10267, n10268, n10269, n10270, n10273, n10274, n10275, n10276;
  wire n10277, n10278, n10279, n10280, n10281, n10282, n10285, n10286;
  wire n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10296;
  wire n10297, n10298, n10299, n10300, n10301, n10302, n10305, n10306;
  wire n10307, n10308, n10309, n10310, n10311, n10312, n10317, n10321;
  wire n10322, n10323, n10324, n10325, n10330, n10331, n10332, n10333;
  wire n10334, n10335, n10336, n10337, n10338, n10339, n10343, n10344;
  wire n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352;
  wire n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360;
  wire n10361, n10362, n10365, n10366, n10367, n10368, n10369, n10370;
  wire n10371, n10372, n10373, n10374, n10377, n10378, n10379, n10380;
  wire n10381, n10382, n10383, n10384, n10385, n10386, n10389, n10390;
  wire n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398;
  wire n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408;
  wire n10409, n10410, n10413, n10414, n10415, n10416, n10417, n10418;
  wire n10419, n10420, n10421, n10422, n10425, n10426, n10427, n10428;
  wire n10429, n10430, n10431, n10432, n10433, n10434, n10437, n10438;
  wire n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446;
  wire n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456;
  wire n10457, n10458, n10461, n10462, n10463, n10464, n10465, n10466;
  wire n10467, n10468, n10469, n10470, n10473, n10474, n10475, n10476;
  wire n10477, n10478, n10479, n10480, n10481, n10482, n10485, n10486;
  wire n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494;
  wire n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504;
  wire n10505, n10506, n10509, n10510, n10511, n10512, n10513, n10514;
  wire n10515, n10516, n10517, n10518, n10521, n10522, n10523, n10524;
  wire n10525, n10526, n10527, n10528, n10529, n10530, n10533, n10534;
  wire n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542;
  wire n10543, n10544, n10547, n10548, n10549, n10550, n10551, n10552;
  wire n10553, n10554, n10557, n10558, n10559, n10560, n10561, n10562;
  wire n10563, n10564, n10565, n10566, n10569, n10570, n10571, n10572;
  wire n10573, n10574, n10575, n10576, n10577, n10578, n10581, n10582;
  wire n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590;
  wire n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600;
  wire n10601, n10602, n10605, n10606, n10607, n10608, n10609, n10610;
  wire n10611, n10612, n10613, n10614, n10617, n10618, n10619, n10620;
  wire n10621, n10622, n10623, n10624, n10625, n10626, n10629, n10630;
  wire n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638;
  wire n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648;
  wire n10649, n10650, n10653, n10654, n10655, n10656, n10657, n10658;
  wire n10659, n10660, n10661, n10662, n10665, n10666, n10667, n10668;
  wire n10669, n10670, n10671, n10672, n10673, n10674, n10677, n10678;
  wire n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686;
  wire n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696;
  wire n10697, n10698, n10701, n10702, n10703, n10704, n10705, n10706;
  wire n10707, n10708, n10709, n10710, n10713, n10714, n10715, n10716;
  wire n10717, n10718, n10719, n10720, n10721, n10722, n10725, n10726;
  wire n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734;
  wire n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744;
  wire n10745, n10746, n10749, n10750, n10751, n10752, n10753, n10754;
  wire n10755, n10756, n10757, n10758, n10761, n10762, n10763, n10764;
  wire n10765, n10766, n10767, n10768, n10769, n10770, n10773, n10774;
  wire n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782;
  wire n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792;
  wire n10793, n10796, n10797, n10798, n10799, n10800, n10801, n10802;
  wire n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812;
  wire n10817, n10821, n10822, n10823, n10824, n10825, n10830, n10831;
  wire n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839;
  wire n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850;
  wire n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858;
  wire n10859, n10860, n10861, n10862, n10865, n10866, n10867, n10868;
  wire n10869, n10870, n10871, n10872, n10873, n10874, n10877, n10878;
  wire n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886;
  wire n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896;
  wire n10897, n10898, n10901, n10902, n10903, n10904, n10905, n10906;
  wire n10907, n10908, n10909, n10910, n10913, n10914, n10915, n10916;
  wire n10917, n10918, n10919, n10920, n10921, n10922, n10925, n10926;
  wire n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934;
  wire n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944;
  wire n10945, n10946, n10949, n10950, n10951, n10952, n10953, n10954;
  wire n10955, n10956, n10957, n10958, n10961, n10962, n10963, n10964;
  wire n10965, n10966, n10967, n10968, n10969, n10970, n10973, n10974;
  wire n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982;
  wire n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992;
  wire n10993, n10994, n10997, n10998, n10999, n11000, n11001, n11002;
  wire n11003, n11004, n11005, n11006, n11009, n11010, n11011, n11012;
  wire n11013, n11014, n11015, n11016, n11017, n11018, n11021, n11022;
  wire n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030;
  wire n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040;
  wire n11041, n11042, n11045, n11046, n11047, n11048, n11049, n11050;
  wire n11051, n11052, n11053, n11054, n11057, n11058, n11059, n11060;
  wire n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068;
  wire n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078;
  wire n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088;
  wire n11089, n11090, n11093, n11094, n11095, n11096, n11097, n11098;
  wire n11099, n11100, n11101, n11102, n11105, n11106, n11107, n11108;
  wire n11109, n11110, n11111, n11112, n11113, n11114, n11117, n11118;
  wire n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126;
  wire n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136;
  wire n11137, n11138, n11141, n11142, n11143, n11144, n11145, n11146;
  wire n11147, n11148, n11149, n11150, n11153, n11154, n11155, n11156;
  wire n11157, n11158, n11159, n11160, n11161, n11162, n11165, n11166;
  wire n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174;
  wire n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184;
  wire n11185, n11186, n11189, n11190, n11191, n11192, n11193, n11194;
  wire n11195, n11196, n11197, n11198, n11201, n11202, n11203, n11204;
  wire n11205, n11206, n11207, n11208, n11209, n11210, n11213, n11214;
  wire n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222;
  wire n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232;
  wire n11233, n11234, n11237, n11238, n11239, n11240, n11241, n11242;
  wire n11243, n11244, n11245, n11246, n11249, n11250, n11251, n11252;
  wire n11253, n11254, n11255, n11256, n11257, n11258, n11261, n11262;
  wire n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270;
  wire n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280;
  wire n11281, n11282, n11285, n11286, n11287, n11288, n11289, n11290;
  wire n11291, n11292, n11293, n11294, n11297, n11298, n11299, n11300;
  wire n11301, n11302, n11303, n11304, n11305, n11308, n11309, n11310;
  wire n11311, n11312, n11313, n11314, n11317, n11318, n11319, n11320;
  wire n11321, n11322, n11323, n11324, n11329, n11333, n11334, n11335;
  wire n11336, n11337, n11342, n11343, n11344, n11345, n11346, n11347;
  wire n11348, n11349, n11350, n11351, n11355, n11356, n11357, n11358;
  wire n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366;
  wire n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374;
  wire n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384;
  wire n11385, n11386, n11389, n11390, n11391, n11392, n11393, n11394;
  wire n11395, n11396, n11397, n11398, n11401, n11402, n11403, n11404;
  wire n11405, n11406, n11407, n11408, n11409, n11410, n11413, n11414;
  wire n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422;
  wire n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432;
  wire n11433, n11434, n11437, n11438, n11439, n11440, n11441, n11442;
  wire n11443, n11444, n11445, n11446, n11449, n11450, n11451, n11452;
  wire n11453, n11454, n11455, n11456, n11457, n11458, n11461, n11462;
  wire n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470;
  wire n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480;
  wire n11481, n11482, n11485, n11486, n11487, n11488, n11489, n11490;
  wire n11491, n11492, n11493, n11494, n11497, n11498, n11499, n11500;
  wire n11501, n11502, n11503, n11504, n11505, n11506, n11509, n11510;
  wire n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518;
  wire n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528;
  wire n11529, n11530, n11533, n11534, n11535, n11536, n11537, n11538;
  wire n11539, n11540, n11541, n11542, n11545, n11546, n11547, n11548;
  wire n11549, n11550, n11551, n11552, n11553, n11554, n11557, n11558;
  wire n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566;
  wire n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576;
  wire n11577, n11578, n11581, n11582, n11583, n11584, n11585, n11586;
  wire n11587, n11588, n11589, n11590, n11593, n11594, n11595, n11596;
  wire n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604;
  wire n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614;
  wire n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624;
  wire n11625, n11626, n11629, n11630, n11631, n11632, n11633, n11634;
  wire n11635, n11636, n11637, n11638, n11641, n11642, n11643, n11644;
  wire n11645, n11646, n11647, n11648, n11649, n11650, n11653, n11654;
  wire n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662;
  wire n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672;
  wire n11673, n11674, n11677, n11678, n11679, n11680, n11681, n11682;
  wire n11683, n11684, n11685, n11686, n11689, n11690, n11691, n11692;
  wire n11693, n11694, n11695, n11696, n11697, n11698, n11701, n11702;
  wire n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710;
  wire n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720;
  wire n11721, n11722, n11725, n11726, n11727, n11728, n11729, n11730;
  wire n11731, n11732, n11733, n11734, n11737, n11738, n11739, n11740;
  wire n11741, n11742, n11743, n11744, n11745, n11746, n11749, n11750;
  wire n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758;
  wire n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768;
  wire n11769, n11770, n11773, n11774, n11775, n11776, n11777, n11778;
  wire n11779, n11780, n11781, n11782, n11785, n11786, n11787, n11788;
  wire n11789, n11790, n11791, n11792, n11793, n11794, n11797, n11798;
  wire n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806;
  wire n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816;
  wire n11817, n11818, n11821, n11822, n11823, n11824, n11825, n11826;
  wire n11827, n11828, n11829, n11832, n11833, n11834, n11835, n11836;
  wire n11837, n11838, n11841, n11842, n11843, n11844, n11845, n11846;
  wire n11847, n11848, n11853, n11857, n11858, n11859, n11860, n11861;
  wire n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873;
  wire n11874, n11875, n11879, n11880, n11881, n11882, n11883, n11884;
  wire n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892;
  wire n11893, n11894, n11895, n11896, n11897, n11898, n11901, n11902;
  wire n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910;
  wire n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920;
  wire n11921, n11922, n11925, n11926, n11927, n11928, n11929, n11930;
  wire n11931, n11932, n11933, n11934, n11937, n11938, n11939, n11940;
  wire n11941, n11942, n11943, n11944, n11945, n11946, n11949, n11950;
  wire n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958;
  wire n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968;
  wire n11969, n11970, n11973, n11974, n11975, n11976, n11977, n11978;
  wire n11979, n11980, n11981, n11982, n11985, n11986, n11987, n11988;
  wire n11989, n11990, n11991, n11992, n11993, n11994, n11997, n11998;
  wire n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006;
  wire n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016;
  wire n12017, n12018, n12021, n12022, n12023, n12024, n12025, n12026;
  wire n12027, n12028, n12029, n12030, n12033, n12034, n12035, n12036;
  wire n12037, n12038, n12039, n12040, n12041, n12042, n12045, n12046;
  wire n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054;
  wire n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064;
  wire n12065, n12066, n12069, n12070, n12071, n12072, n12073, n12074;
  wire n12075, n12076, n12077, n12078, n12081, n12082, n12083, n12084;
  wire n12085, n12086, n12087, n12088, n12089, n12090, n12093, n12094;
  wire n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102;
  wire n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112;
  wire n12113, n12114, n12117, n12118, n12119, n12120, n12121, n12122;
  wire n12123, n12124, n12125, n12126, n12129, n12130, n12131, n12132;
  wire n12133, n12134, n12135, n12136, n12137, n12138, n12141, n12142;
  wire n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150;
  wire n12151, n12152, n12155, n12156, n12157, n12158, n12159, n12160;
  wire n12161, n12162, n12165, n12166, n12167, n12168, n12169, n12170;
  wire n12171, n12172, n12173, n12174, n12177, n12178, n12179, n12180;
  wire n12181, n12182, n12183, n12184, n12185, n12186, n12189, n12190;
  wire n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198;
  wire n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208;
  wire n12209, n12210, n12213, n12214, n12215, n12216, n12217, n12218;
  wire n12219, n12220, n12221, n12222, n12225, n12226, n12227, n12228;
  wire n12229, n12230, n12231, n12232, n12233, n12234, n12237, n12238;
  wire n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246;
  wire n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256;
  wire n12257, n12258, n12261, n12262, n12263, n12264, n12265, n12266;
  wire n12267, n12268, n12269, n12270, n12273, n12274, n12275, n12276;
  wire n12277, n12278, n12279, n12280, n12281, n12282, n12285, n12286;
  wire n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294;
  wire n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304;
  wire n12305, n12306, n12309, n12310, n12311, n12312, n12313, n12314;
  wire n12315, n12316, n12317, n12318, n12321, n12322, n12323, n12324;
  wire n12325, n12326, n12327, n12328, n12329, n12330, n12333, n12334;
  wire n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342;
  wire n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352;
  wire n12353, n12354, n12357, n12358, n12359, n12360, n12361, n12362;
  wire n12363, n12364, n12365, n12368, n12369, n12370, n12371, n12372;
  wire n12373, n12374, n12377, n12378, n12379, n12380, n12381, n12382;
  wire n12383, n12384, n12389, n12393, n12394, n12395, n12396, n12397;
  wire n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409;
  wire n12410, n12411, n12415, n12416, n12417, n12418, n12419, n12420;
  wire n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428;
  wire n12429, n12430, n12431, n12432, n12433, n12434, n12437, n12438;
  wire n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446;
  wire n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456;
  wire n12457, n12458, n12461, n12462, n12463, n12464, n12465, n12466;
  wire n12467, n12468, n12469, n12470, n12473, n12474, n12475, n12476;
  wire n12477, n12478, n12479, n12480, n12481, n12482, n12485, n12486;
  wire n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494;
  wire n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504;
  wire n12505, n12506, n12509, n12510, n12511, n12512, n12513, n12514;
  wire n12515, n12516, n12517, n12518, n12521, n12522, n12523, n12524;
  wire n12525, n12526, n12527, n12528, n12529, n12530, n12533, n12534;
  wire n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542;
  wire n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552;
  wire n12553, n12554, n12557, n12558, n12559, n12560, n12561, n12562;
  wire n12563, n12564, n12565, n12566, n12569, n12570, n12571, n12572;
  wire n12573, n12574, n12575, n12576, n12577, n12578, n12581, n12582;
  wire n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590;
  wire n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600;
  wire n12601, n12602, n12605, n12606, n12607, n12608, n12609, n12610;
  wire n12611, n12612, n12613, n12614, n12617, n12618, n12619, n12620;
  wire n12621, n12622, n12623, n12624, n12625, n12626, n12629, n12630;
  wire n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638;
  wire n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648;
  wire n12649, n12650, n12653, n12654, n12655, n12656, n12657, n12658;
  wire n12659, n12660, n12661, n12662, n12665, n12666, n12667, n12668;
  wire n12669, n12670, n12671, n12672, n12673, n12674, n12677, n12678;
  wire n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686;
  wire n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696;
  wire n12697, n12698, n12701, n12702, n12703, n12704, n12705, n12706;
  wire n12707, n12708, n12709, n12710, n12711, n12712, n12715, n12716;
  wire n12717, n12718, n12719, n12720, n12721, n12722, n12725, n12726;
  wire n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734;
  wire n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744;
  wire n12745, n12746, n12749, n12750, n12751, n12752, n12753, n12754;
  wire n12755, n12756, n12757, n12758, n12761, n12762, n12763, n12764;
  wire n12765, n12766, n12767, n12768, n12769, n12770, n12773, n12774;
  wire n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782;
  wire n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792;
  wire n12793, n12794, n12797, n12798, n12799, n12800, n12801, n12802;
  wire n12803, n12804, n12805, n12806, n12809, n12810, n12811, n12812;
  wire n12813, n12814, n12815, n12816, n12817, n12818, n12821, n12822;
  wire n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830;
  wire n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840;
  wire n12841, n12842, n12845, n12846, n12847, n12848, n12849, n12850;
  wire n12851, n12852, n12853, n12854, n12857, n12858, n12859, n12860;
  wire n12861, n12862, n12863, n12864, n12865, n12866, n12869, n12870;
  wire n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878;
  wire n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888;
  wire n12889, n12890, n12893, n12894, n12895, n12896, n12897, n12898;
  wire n12899, n12900, n12901, n12902, n12905, n12906, n12907, n12908;
  wire n12909, n12910, n12911, n12912, n12913, n12916, n12917, n12918;
  wire n12919, n12920, n12921, n12922, n12925, n12926, n12927, n12928;
  wire n12929, n12930, n12931, n12932, n12937, n12941, n12942, n12943;
  wire n12944, n12945, n12950, n12951, n12952, n12953, n12954, n12955;
  wire n12956, n12957, n12958, n12959, n12963, n12964, n12965, n12966;
  wire n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974;
  wire n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982;
  wire n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992;
  wire n12993, n12994, n12997, n12998, n12999, n13000, n13001, n13002;
  wire n13003, n13004, n13005, n13006, n13009, n13010, n13011, n13012;
  wire n13013, n13014, n13015, n13016, n13017, n13018, n13021, n13022;
  wire n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030;
  wire n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040;
  wire n13041, n13042, n13045, n13046, n13047, n13048, n13049, n13050;
  wire n13051, n13052, n13053, n13054, n13057, n13058, n13059, n13060;
  wire n13061, n13062, n13063, n13064, n13065, n13066, n13069, n13070;
  wire n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078;
  wire n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088;
  wire n13089, n13090, n13093, n13094, n13095, n13096, n13097, n13098;
  wire n13099, n13100, n13101, n13102, n13105, n13106, n13107, n13108;
  wire n13109, n13110, n13111, n13112, n13113, n13114, n13117, n13118;
  wire n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126;
  wire n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136;
  wire n13137, n13138, n13141, n13142, n13143, n13144, n13145, n13146;
  wire n13147, n13148, n13149, n13150, n13153, n13154, n13155, n13156;
  wire n13157, n13158, n13159, n13160, n13161, n13162, n13165, n13166;
  wire n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174;
  wire n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184;
  wire n13185, n13186, n13189, n13190, n13191, n13192, n13193, n13194;
  wire n13195, n13196, n13197, n13198, n13201, n13202, n13203, n13204;
  wire n13205, n13206, n13207, n13208, n13209, n13210, n13213, n13214;
  wire n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222;
  wire n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232;
  wire n13233, n13234, n13237, n13238, n13239, n13240, n13241, n13242;
  wire n13243, n13244, n13245, n13246, n13249, n13250, n13251, n13252;
  wire n13253, n13254, n13255, n13256, n13257, n13258, n13261, n13262;
  wire n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270;
  wire n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280;
  wire n13281, n13282, n13283, n13284, n13287, n13288, n13289, n13290;
  wire n13291, n13292, n13293, n13294, n13297, n13298, n13299, n13300;
  wire n13301, n13302, n13303, n13304, n13305, n13306, n13309, n13310;
  wire n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318;
  wire n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328;
  wire n13329, n13330, n13333, n13334, n13335, n13336, n13337, n13338;
  wire n13339, n13340, n13341, n13342, n13345, n13346, n13347, n13348;
  wire n13349, n13350, n13351, n13352, n13353, n13354, n13357, n13358;
  wire n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366;
  wire n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376;
  wire n13377, n13378, n13381, n13382, n13383, n13384, n13385, n13386;
  wire n13387, n13388, n13389, n13390, n13393, n13394, n13395, n13396;
  wire n13397, n13398, n13399, n13400, n13401, n13402, n13405, n13406;
  wire n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414;
  wire n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424;
  wire n13425, n13426, n13429, n13430, n13431, n13432, n13433, n13434;
  wire n13435, n13436, n13437, n13438, n13441, n13442, n13443, n13444;
  wire n13445, n13446, n13447, n13448, n13449, n13450, n13453, n13454;
  wire n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462;
  wire n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472;
  wire n13473, n13476, n13477, n13478, n13479, n13480, n13481, n13482;
  wire n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492;
  wire n13497, n13501, n13502, n13503, n13504, n13505, n13510, n13511;
  wire n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519;
  wire n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530;
  wire n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538;
  wire n13539, n13540, n13541, n13542, n13545, n13546, n13547, n13548;
  wire n13549, n13550, n13551, n13552, n13553, n13554, n13557, n13558;
  wire n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566;
  wire n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576;
  wire n13577, n13578, n13581, n13582, n13583, n13584, n13585, n13586;
  wire n13587, n13588, n13589, n13590, n13593, n13594, n13595, n13596;
  wire n13597, n13598, n13599, n13600, n13601, n13602, n13605, n13606;
  wire n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614;
  wire n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624;
  wire n13625, n13626, n13629, n13630, n13631, n13632, n13633, n13634;
  wire n13635, n13636, n13637, n13638, n13641, n13642, n13643, n13644;
  wire n13645, n13646, n13647, n13648, n13649, n13650, n13653, n13654;
  wire n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662;
  wire n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672;
  wire n13673, n13674, n13677, n13678, n13679, n13680, n13681, n13682;
  wire n13683, n13684, n13685, n13686, n13689, n13690, n13691, n13692;
  wire n13693, n13694, n13695, n13696, n13697, n13698, n13701, n13702;
  wire n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710;
  wire n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720;
  wire n13721, n13722, n13725, n13726, n13727, n13728, n13729, n13730;
  wire n13731, n13732, n13733, n13734, n13737, n13738, n13739, n13740;
  wire n13741, n13742, n13743, n13744, n13745, n13746, n13749, n13750;
  wire n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758;
  wire n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768;
  wire n13769, n13770, n13773, n13774, n13775, n13776, n13777, n13778;
  wire n13779, n13780, n13781, n13782, n13785, n13786, n13787, n13788;
  wire n13789, n13790, n13791, n13792, n13793, n13794, n13797, n13798;
  wire n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806;
  wire n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816;
  wire n13817, n13818, n13821, n13822, n13823, n13824, n13825, n13826;
  wire n13827, n13828, n13829, n13830, n13833, n13834, n13835, n13836;
  wire n13837, n13838, n13839, n13840, n13841, n13842, n13845, n13846;
  wire n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854;
  wire n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864;
  wire n13865, n13866, n13867, n13868, n13871, n13872, n13873, n13874;
  wire n13875, n13876, n13877, n13878, n13881, n13882, n13883, n13884;
  wire n13885, n13886, n13887, n13888, n13889, n13890, n13893, n13894;
  wire n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902;
  wire n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912;
  wire n13913, n13914, n13917, n13918, n13919, n13920, n13921, n13922;
  wire n13923, n13924, n13925, n13926, n13929, n13930, n13931, n13932;
  wire n13933, n13934, n13935, n13936, n13937, n13938, n13941, n13942;
  wire n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950;
  wire n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960;
  wire n13961, n13962, n13965, n13966, n13967, n13968, n13969, n13970;
  wire n13971, n13972, n13973, n13974, n13977, n13978, n13979, n13980;
  wire n13981, n13982, n13983, n13984, n13985, n13986, n13989, n13990;
  wire n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998;
  wire n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008;
  wire n14009, n14010, n14013, n14014, n14015, n14016, n14017, n14018;
  wire n14019, n14020, n14021, n14022, n14025, n14026, n14027, n14028;
  wire n14029, n14030, n14031, n14032, n14033, n14034, n14037, n14038;
  wire n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14048;
  wire n14049, n14050, n14051, n14052, n14053, n14054, n14057, n14058;
  wire n14059, n14060, n14061, n14062, n14063, n14064, n14069, n14073;
  wire n14074, n14075, n14076, n14077, n14082, n14083, n14084, n14085;
  wire n14086, n14087, n14088, n14089, n14090, n14091, n14095, n14096;
  wire n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104;
  wire n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112;
  wire n14113, n14114, n14117, n14118, n14119, n14120, n14121, n14122;
  wire n14123, n14124, n14125, n14126, n14129, n14130, n14131, n14132;
  wire n14133, n14134, n14135, n14136, n14137, n14138, n14141, n14142;
  wire n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150;
  wire n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160;
  wire n14161, n14162, n14165, n14166, n14167, n14168, n14169, n14170;
  wire n14171, n14172, n14173, n14174, n14177, n14178, n14179, n14180;
  wire n14181, n14182, n14183, n14184, n14185, n14186, n14189, n14190;
  wire n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198;
  wire n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208;
  wire n14209, n14210, n14213, n14214, n14215, n14216, n14217, n14218;
  wire n14219, n14220, n14221, n14222, n14225, n14226, n14227, n14228;
  wire n14229, n14230, n14231, n14232, n14233, n14234, n14237, n14238;
  wire n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246;
  wire n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256;
  wire n14257, n14258, n14261, n14262, n14263, n14264, n14265, n14266;
  wire n14267, n14268, n14269, n14270, n14273, n14274, n14275, n14276;
  wire n14277, n14278, n14279, n14280, n14281, n14282, n14285, n14286;
  wire n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294;
  wire n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304;
  wire n14305, n14306, n14309, n14310, n14311, n14312, n14313, n14314;
  wire n14315, n14316, n14317, n14318, n14321, n14322, n14323, n14324;
  wire n14325, n14326, n14327, n14328, n14329, n14330, n14333, n14334;
  wire n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342;
  wire n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352;
  wire n14353, n14354, n14357, n14358, n14359, n14360, n14361, n14362;
  wire n14363, n14364, n14365, n14366, n14369, n14370, n14371, n14372;
  wire n14373, n14374, n14375, n14376, n14377, n14378, n14381, n14382;
  wire n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390;
  wire n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400;
  wire n14401, n14402, n14405, n14406, n14407, n14408, n14409, n14410;
  wire n14411, n14412, n14413, n14414, n14417, n14418, n14419, n14420;
  wire n14421, n14422, n14423, n14424, n14425, n14426, n14429, n14430;
  wire n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438;
  wire n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448;
  wire n14449, n14450, n14453, n14454, n14455, n14456, n14457, n14458;
  wire n14459, n14460, n14461, n14462, n14463, n14464, n14467, n14468;
  wire n14469, n14470, n14471, n14472, n14473, n14474, n14477, n14478;
  wire n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486;
  wire n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496;
  wire n14497, n14498, n14501, n14502, n14503, n14504, n14505, n14506;
  wire n14507, n14508, n14509, n14510, n14513, n14514, n14515, n14516;
  wire n14517, n14518, n14519, n14520, n14521, n14522, n14525, n14526;
  wire n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534;
  wire n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544;
  wire n14545, n14546, n14549, n14550, n14551, n14552, n14553, n14554;
  wire n14555, n14556, n14557, n14558, n14561, n14562, n14563, n14564;
  wire n14565, n14566, n14567, n14568, n14569, n14570, n14573, n14574;
  wire n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582;
  wire n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592;
  wire n14593, n14594, n14597, n14598, n14599, n14600, n14601, n14602;
  wire n14603, n14604, n14605, n14606, n14609, n14610, n14611, n14612;
  wire n14613, n14614, n14615, n14616, n14617, n14618, n14621, n14622;
  wire n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14632;
  wire n14633, n14634, n14635, n14636, n14637, n14638, n14641, n14642;
  wire n14643, n14644, n14645, n14646, n14647, n14648, n14653, n14657;
  wire n14658, n14659, n14660, n14661, n14666, n14667, n14668, n14669;
  wire n14670, n14671, n14672, n14673, n14674, n14675, n14679, n14680;
  wire n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688;
  wire n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696;
  wire n14697, n14698, n14701, n14702, n14703, n14704, n14705, n14706;
  wire n14707, n14708, n14709, n14710, n14713, n14714, n14715, n14716;
  wire n14717, n14718, n14719, n14720, n14721, n14722, n14725, n14726;
  wire n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734;
  wire n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744;
  wire n14745, n14746, n14749, n14750, n14751, n14752, n14753, n14754;
  wire n14755, n14756, n14757, n14758, n14761, n14762, n14763, n14764;
  wire n14765, n14766, n14767, n14768, n14769, n14770, n14773, n14774;
  wire n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782;
  wire n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792;
  wire n14793, n14794, n14797, n14798, n14799, n14800, n14801, n14802;
  wire n14803, n14804, n14805, n14806, n14809, n14810, n14811, n14812;
  wire n14813, n14814, n14815, n14816, n14817, n14818, n14821, n14822;
  wire n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830;
  wire n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840;
  wire n14841, n14842, n14845, n14846, n14847, n14848, n14849, n14850;
  wire n14851, n14852, n14853, n14854, n14857, n14858, n14859, n14860;
  wire n14861, n14862, n14863, n14864, n14865, n14866, n14869, n14870;
  wire n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878;
  wire n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888;
  wire n14889, n14890, n14893, n14894, n14895, n14896, n14897, n14898;
  wire n14899, n14900, n14901, n14902, n14905, n14906, n14907, n14908;
  wire n14909, n14910, n14911, n14912, n14913, n14914, n14917, n14918;
  wire n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926;
  wire n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936;
  wire n14937, n14938, n14941, n14942, n14943, n14944, n14945, n14946;
  wire n14947, n14948, n14949, n14950, n14953, n14954, n14955, n14956;
  wire n14957, n14958, n14959, n14960, n14961, n14962, n14965, n14966;
  wire n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974;
  wire n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984;
  wire n14985, n14986, n14989, n14990, n14991, n14992, n14993, n14994;
  wire n14995, n14996, n14997, n14998, n15001, n15002, n15003, n15004;
  wire n15005, n15006, n15007, n15008, n15009, n15010, n15013, n15014;
  wire n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022;
  wire n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032;
  wire n15033, n15034, n15037, n15038, n15039, n15040, n15041, n15042;
  wire n15043, n15044, n15045, n15046, n15049, n15050, n15051, n15052;
  wire n15053, n15054, n15055, n15056, n15057, n15058, n15061, n15062;
  wire n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070;
  wire n15071, n15072, n15075, n15076, n15077, n15078, n15079, n15080;
  wire n15081, n15082, n15085, n15086, n15087, n15088, n15089, n15090;
  wire n15091, n15092, n15093, n15094, n15097, n15098, n15099, n15100;
  wire n15101, n15102, n15103, n15104, n15105, n15106, n15109, n15110;
  wire n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118;
  wire n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128;
  wire n15129, n15130, n15133, n15134, n15135, n15136, n15137, n15138;
  wire n15139, n15140, n15141, n15142, n15145, n15146, n15147, n15148;
  wire n15149, n15150, n15151, n15152, n15153, n15154, n15157, n15158;
  wire n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166;
  wire n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176;
  wire n15177, n15178, n15181, n15182, n15183, n15184, n15185, n15186;
  wire n15187, n15188, n15189, n15190, n15193, n15194, n15195, n15196;
  wire n15197, n15198, n15199, n15200, n15201, n15202, n15205, n15206;
  wire n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214;
  wire n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224;
  wire n15225, n15228, n15229, n15230, n15231, n15232, n15233, n15234;
  wire n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244;
  wire n15249, n15253, n15254, n15255, n15256, n15257, n15262, n15263;
  wire n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271;
  wire n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282;
  wire n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290;
  wire n15291, n15292, n15293, n15294, n15297, n15298, n15299, n15300;
  wire n15301, n15302, n15303, n15304, n15305, n15306, n15309, n15310;
  wire n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318;
  wire n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328;
  wire n15329, n15330, n15333, n15334, n15335, n15336, n15337, n15338;
  wire n15339, n15340, n15341, n15342, n15345, n15346, n15347, n15348;
  wire n15349, n15350, n15351, n15352, n15353, n15354, n15357, n15358;
  wire n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366;
  wire n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376;
  wire n15377, n15378, n15381, n15382, n15383, n15384, n15385, n15386;
  wire n15387, n15388, n15389, n15390, n15393, n15394, n15395, n15396;
  wire n15397, n15398, n15399, n15400, n15401, n15402, n15405, n15406;
  wire n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414;
  wire n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424;
  wire n15425, n15426, n15429, n15430, n15431, n15432, n15433, n15434;
  wire n15435, n15436, n15437, n15438, n15441, n15442, n15443, n15444;
  wire n15445, n15446, n15447, n15448, n15449, n15450, n15453, n15454;
  wire n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462;
  wire n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472;
  wire n15473, n15474, n15477, n15478, n15479, n15480, n15481, n15482;
  wire n15483, n15484, n15485, n15486, n15489, n15490, n15491, n15492;
  wire n15493, n15494, n15495, n15496, n15497, n15498, n15501, n15502;
  wire n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510;
  wire n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520;
  wire n15521, n15522, n15525, n15526, n15527, n15528, n15529, n15530;
  wire n15531, n15532, n15533, n15534, n15537, n15538, n15539, n15540;
  wire n15541, n15542, n15543, n15544, n15545, n15546, n15549, n15550;
  wire n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558;
  wire n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568;
  wire n15569, n15570, n15573, n15574, n15575, n15576, n15577, n15578;
  wire n15579, n15580, n15581, n15582, n15585, n15586, n15587, n15588;
  wire n15589, n15590, n15591, n15592, n15593, n15594, n15597, n15598;
  wire n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606;
  wire n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616;
  wire n15617, n15618, n15621, n15622, n15623, n15624, n15625, n15626;
  wire n15627, n15628, n15629, n15630, n15633, n15634, n15635, n15636;
  wire n15637, n15638, n15639, n15640, n15641, n15642, n15645, n15646;
  wire n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654;
  wire n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664;
  wire n15665, n15666, n15669, n15670, n15671, n15672, n15673, n15674;
  wire n15675, n15676, n15677, n15678, n15681, n15682, n15683, n15684;
  wire n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692;
  wire n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702;
  wire n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712;
  wire n15713, n15714, n15717, n15718, n15719, n15720, n15721, n15722;
  wire n15723, n15724, n15725, n15726, n15729, n15730, n15731, n15732;
  wire n15733, n15734, n15735, n15736, n15737, n15738, n15741, n15742;
  wire n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750;
  wire n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760;
  wire n15761, n15762, n15765, n15766, n15767, n15768, n15769, n15770;
  wire n15771, n15772, n15773, n15774, n15777, n15778, n15779, n15780;
  wire n15781, n15782, n15783, n15784, n15785, n15786, n15789, n15790;
  wire n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798;
  wire n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808;
  wire n15809, n15810, n15813, n15814, n15815, n15816, n15817, n15818;
  wire n15819, n15820, n15821, n15822, n15825, n15826, n15827, n15828;
  wire n15829, n15830, n15831, n15832, n15833, n15836, n15837, n15838;
  wire n15839, n15840, n15841, n15842, n15845, n15846, n15847, n15848;
  wire n15849, n15850, n15851, n15852, n15857, n15861, n15862, n15863;
  wire n15864, n15865, n15870, n15871, n15872, n15873, n15874, n15875;
  wire n15876, n15877, n15878, n15879, n15883, n15884, n15885, n15886;
  wire n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894;
  wire n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902;
  wire n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912;
  wire n15913, n15914, n15917, n15918, n15919, n15920, n15921, n15922;
  wire n15923, n15924, n15925, n15926, n15929, n15930, n15931, n15932;
  wire n15933, n15934, n15935, n15936, n15937, n15938, n15941, n15942;
  wire n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950;
  wire n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960;
  wire n15961, n15962, n15965, n15966, n15967, n15968, n15969, n15970;
  wire n15971, n15972, n15973, n15974, n15977, n15978, n15979, n15980;
  wire n15981, n15982, n15983, n15984, n15985, n15986, n15989, n15990;
  wire n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998;
  wire n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008;
  wire n16009, n16010, n16013, n16014, n16015, n16016, n16017, n16018;
  wire n16019, n16020, n16021, n16022, n16025, n16026, n16027, n16028;
  wire n16029, n16030, n16031, n16032, n16033, n16034, n16037, n16038;
  wire n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046;
  wire n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056;
  wire n16057, n16058, n16061, n16062, n16063, n16064, n16065, n16066;
  wire n16067, n16068, n16069, n16070, n16073, n16074, n16075, n16076;
  wire n16077, n16078, n16079, n16080, n16081, n16082, n16085, n16086;
  wire n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094;
  wire n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104;
  wire n16105, n16106, n16109, n16110, n16111, n16112, n16113, n16114;
  wire n16115, n16116, n16117, n16118, n16121, n16122, n16123, n16124;
  wire n16125, n16126, n16127, n16128, n16129, n16130, n16133, n16134;
  wire n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142;
  wire n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152;
  wire n16153, n16154, n16157, n16158, n16159, n16160, n16161, n16162;
  wire n16163, n16164, n16165, n16166, n16169, n16170, n16171, n16172;
  wire n16173, n16174, n16175, n16176, n16177, n16178, n16181, n16182;
  wire n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190;
  wire n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200;
  wire n16201, n16202, n16205, n16206, n16207, n16208, n16209, n16210;
  wire n16211, n16212, n16213, n16214, n16217, n16218, n16219, n16220;
  wire n16221, n16222, n16223, n16224, n16225, n16226, n16229, n16230;
  wire n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238;
  wire n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248;
  wire n16249, n16250, n16253, n16254, n16255, n16256, n16257, n16258;
  wire n16259, n16260, n16261, n16262, n16265, n16266, n16267, n16268;
  wire n16269, n16270, n16271, n16272, n16273, n16274, n16277, n16278;
  wire n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286;
  wire n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296;
  wire n16297, n16298, n16301, n16302, n16303, n16304, n16305, n16306;
  wire n16307, n16308, n16309, n16310, n16313, n16314, n16315, n16316;
  wire n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324;
  wire n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334;
  wire n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344;
  wire n16345, n16346, n16349, n16350, n16351, n16352, n16353, n16354;
  wire n16355, n16356, n16357, n16358, n16361, n16362, n16363, n16364;
  wire n16365, n16366, n16367, n16368, n16369, n16370, n16373, n16374;
  wire n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382;
  wire n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392;
  wire n16393, n16394, n16397, n16398, n16399, n16400, n16401, n16402;
  wire n16403, n16404, n16405, n16406, n16409, n16410, n16411, n16412;
  wire n16413, n16414, n16415, n16416, n16417, n16418, n16421, n16422;
  wire n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430;
  wire n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440;
  wire n16441, n16442, n16445, n16446, n16447, n16448, n16449, n16450;
  wire n16451, n16452, n16453, n16456, n16457, n16458, n16459, n16460;
  wire n16461, n16462, n16465, n16466, n16467, n16468, n16469, n16470;
  wire n16471, n16472, n16477, n16481, n16482, n16483, n16484, n16485;
  wire n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497;
  wire n16498, n16499, n16503, n16504, n16505, n16506, n16507, n16508;
  wire n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516;
  wire n16517, n16518, n16519, n16520, n16521, n16522, n16525, n16526;
  wire n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534;
  wire n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544;
  wire n16545, n16546, n16549, n16550, n16551, n16552, n16553, n16554;
  wire n16555, n16556, n16557, n16558, n16561, n16562, n16563, n16564;
  wire n16565, n16566, n16567, n16568, n16569, n16570, n16573, n16574;
  wire n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582;
  wire n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592;
  wire n16593, n16594, n16597, n16598, n16599, n16600, n16601, n16602;
  wire n16603, n16604, n16605, n16606, n16609, n16610, n16611, n16612;
  wire n16613, n16614, n16615, n16616, n16617, n16618, n16621, n16622;
  wire n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630;
  wire n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640;
  wire n16641, n16642, n16645, n16646, n16647, n16648, n16649, n16650;
  wire n16651, n16652, n16653, n16654, n16657, n16658, n16659, n16660;
  wire n16661, n16662, n16663, n16664, n16665, n16666, n16669, n16670;
  wire n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678;
  wire n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688;
  wire n16689, n16690, n16693, n16694, n16695, n16696, n16697, n16698;
  wire n16699, n16700, n16701, n16702, n16705, n16706, n16707, n16708;
  wire n16709, n16710, n16711, n16712, n16713, n16714, n16717, n16718;
  wire n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726;
  wire n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736;
  wire n16737, n16738, n16741, n16742, n16743, n16744, n16745, n16746;
  wire n16747, n16748, n16749, n16750, n16753, n16754, n16755, n16756;
  wire n16757, n16758, n16759, n16760, n16761, n16762, n16765, n16766;
  wire n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774;
  wire n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784;
  wire n16785, n16786, n16789, n16790, n16791, n16792, n16793, n16794;
  wire n16795, n16796, n16797, n16798, n16801, n16802, n16803, n16804;
  wire n16805, n16806, n16807, n16808, n16809, n16810, n16813, n16814;
  wire n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822;
  wire n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832;
  wire n16833, n16834, n16837, n16838, n16839, n16840, n16841, n16842;
  wire n16843, n16844, n16845, n16846, n16849, n16850, n16851, n16852;
  wire n16853, n16854, n16855, n16856, n16857, n16858, n16861, n16862;
  wire n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870;
  wire n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880;
  wire n16881, n16882, n16885, n16886, n16887, n16888, n16889, n16890;
  wire n16891, n16892, n16893, n16894, n16897, n16898, n16899, n16900;
  wire n16901, n16902, n16903, n16904, n16905, n16906, n16909, n16910;
  wire n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918;
  wire n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928;
  wire n16929, n16930, n16933, n16934, n16935, n16936, n16937, n16938;
  wire n16939, n16940, n16941, n16942, n16945, n16946, n16947, n16948;
  wire n16949, n16950, n16951, n16952, n16953, n16954, n16957, n16958;
  wire n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966;
  wire n16967, n16968, n16971, n16972, n16973, n16974, n16975, n16976;
  wire n16977, n16978, n16981, n16982, n16983, n16984, n16985, n16986;
  wire n16987, n16988, n16989, n16990, n16993, n16994, n16995, n16996;
  wire n16997, n16998, n16999, n17000, n17001, n17002, n17005, n17006;
  wire n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014;
  wire n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024;
  wire n17025, n17026, n17029, n17030, n17031, n17032, n17033, n17034;
  wire n17035, n17036, n17037, n17038, n17041, n17042, n17043, n17044;
  wire n17045, n17046, n17047, n17048, n17049, n17050, n17053, n17054;
  wire n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062;
  wire n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072;
  wire n17073, n17074, n17077, n17078, n17079, n17080, n17081, n17082;
  wire n17083, n17084, n17085, n17088, n17089, n17090, n17091, n17092;
  wire n17093, n17094, n17097, n17098, n17099, n17100, n17101, n17102;
  wire n17103, n17104, n17109, n17113, n17114, n17115, n17116, n17117;
  wire n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129;
  wire n17130, n17131, n17135, n17136, n17137, n17138, n17139, n17140;
  wire n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148;
  wire n17149, n17150, n17151, n17152, n17153, n17154, n17157, n17158;
  wire n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166;
  wire n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176;
  wire n17177, n17178, n17181, n17182, n17183, n17184, n17185, n17186;
  wire n17187, n17188, n17189, n17190, n17193, n17194, n17195, n17196;
  wire n17197, n17198, n17199, n17200, n17201, n17202, n17205, n17206;
  wire n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214;
  wire n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224;
  wire n17225, n17226, n17229, n17230, n17231, n17232, n17233, n17234;
  wire n17235, n17236, n17237, n17238, n17241, n17242, n17243, n17244;
  wire n17245, n17246, n17247, n17248, n17249, n17250, n17253, n17254;
  wire n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262;
  wire n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272;
  wire n17273, n17274, n17277, n17278, n17279, n17280, n17281, n17282;
  wire n17283, n17284, n17285, n17286, n17289, n17290, n17291, n17292;
  wire n17293, n17294, n17295, n17296, n17297, n17298, n17301, n17302;
  wire n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310;
  wire n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320;
  wire n17321, n17322, n17325, n17326, n17327, n17328, n17329, n17330;
  wire n17331, n17332, n17333, n17334, n17337, n17338, n17339, n17340;
  wire n17341, n17342, n17343, n17344, n17345, n17346, n17349, n17350;
  wire n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358;
  wire n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368;
  wire n17369, n17370, n17373, n17374, n17375, n17376, n17377, n17378;
  wire n17379, n17380, n17381, n17382, n17385, n17386, n17387, n17388;
  wire n17389, n17390, n17391, n17392, n17393, n17394, n17397, n17398;
  wire n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406;
  wire n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416;
  wire n17417, n17418, n17421, n17422, n17423, n17424, n17425, n17426;
  wire n17427, n17428, n17429, n17430, n17433, n17434, n17435, n17436;
  wire n17437, n17438, n17439, n17440, n17441, n17442, n17445, n17446;
  wire n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454;
  wire n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464;
  wire n17465, n17466, n17469, n17470, n17471, n17472, n17473, n17474;
  wire n17475, n17476, n17477, n17478, n17481, n17482, n17483, n17484;
  wire n17485, n17486, n17487, n17488, n17489, n17490, n17493, n17494;
  wire n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502;
  wire n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512;
  wire n17513, n17514, n17517, n17518, n17519, n17520, n17521, n17522;
  wire n17523, n17524, n17525, n17526, n17529, n17530, n17531, n17532;
  wire n17533, n17534, n17535, n17536, n17537, n17538, n17541, n17542;
  wire n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550;
  wire n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560;
  wire n17561, n17562, n17565, n17566, n17567, n17568, n17569, n17570;
  wire n17571, n17572, n17573, n17574, n17577, n17578, n17579, n17580;
  wire n17581, n17582, n17583, n17584, n17585, n17586, n17589, n17590;
  wire n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598;
  wire n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608;
  wire n17609, n17610, n17613, n17614, n17615, n17616, n17617, n17618;
  wire n17619, n17620, n17621, n17622, n17623, n17624, n17627, n17628;
  wire n17629, n17630, n17631, n17632, n17633, n17634, n17637, n17638;
  wire n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646;
  wire n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656;
  wire n17657, n17658, n17661, n17662, n17663, n17664, n17665, n17666;
  wire n17667, n17668, n17669, n17670, n17673, n17674, n17675, n17676;
  wire n17677, n17678, n17679, n17680, n17681, n17682, n17685, n17686;
  wire n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694;
  wire n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704;
  wire n17705, n17706, n17709, n17710, n17711, n17712, n17713, n17714;
  wire n17715, n17716, n17717, n17718, n17721, n17722, n17723, n17724;
  wire n17725, n17726, n17727, n17728, n17729, n17732, n17733, n17734;
  wire n17735, n17736, n17737, n17738, n17741, n17742, n17743, n17744;
  wire n17745, n17746, n17747, n17748, n17753, n17757, n17758, n17759;
  wire n17760, n17761, n17766, n17767, n17768, n17769, n17770, n17771;
  wire n17772, n17773, n17774, n17775, n17779, n17780, n17781, n17782;
  wire n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790;
  wire n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798;
  wire n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808;
  wire n17809, n17810, n17813, n17814, n17815, n17816, n17817, n17818;
  wire n17819, n17820, n17821, n17822, n17825, n17826, n17827, n17828;
  wire n17829, n17830, n17831, n17832, n17833, n17834, n17837, n17838;
  wire n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846;
  wire n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856;
  wire n17857, n17858, n17861, n17862, n17863, n17864, n17865, n17866;
  wire n17867, n17868, n17869, n17870, n17873, n17874, n17875, n17876;
  wire n17877, n17878, n17879, n17880, n17881, n17882, n17885, n17886;
  wire n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894;
  wire n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904;
  wire n17905, n17906, n17909, n17910, n17911, n17912, n17913, n17914;
  wire n17915, n17916, n17917, n17918, n17921, n17922, n17923, n17924;
  wire n17925, n17926, n17927, n17928, n17929, n17930, n17933, n17934;
  wire n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942;
  wire n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952;
  wire n17953, n17954, n17957, n17958, n17959, n17960, n17961, n17962;
  wire n17963, n17964, n17965, n17966, n17969, n17970, n17971, n17972;
  wire n17973, n17974, n17975, n17976, n17977, n17978, n17981, n17982;
  wire n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990;
  wire n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000;
  wire n18001, n18002, n18005, n18006, n18007, n18008, n18009, n18010;
  wire n18011, n18012, n18013, n18014, n18017, n18018, n18019, n18020;
  wire n18021, n18022, n18023, n18024, n18025, n18026, n18029, n18030;
  wire n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038;
  wire n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048;
  wire n18049, n18050, n18053, n18054, n18055, n18056, n18057, n18058;
  wire n18059, n18060, n18061, n18062, n18065, n18066, n18067, n18068;
  wire n18069, n18070, n18071, n18072, n18073, n18074, n18077, n18078;
  wire n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086;
  wire n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096;
  wire n18097, n18098, n18101, n18102, n18103, n18104, n18105, n18106;
  wire n18107, n18108, n18109, n18110, n18113, n18114, n18115, n18116;
  wire n18117, n18118, n18119, n18120, n18121, n18122, n18125, n18126;
  wire n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134;
  wire n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144;
  wire n18145, n18146, n18149, n18150, n18151, n18152, n18153, n18154;
  wire n18155, n18156, n18157, n18158, n18161, n18162, n18163, n18164;
  wire n18165, n18166, n18167, n18168, n18169, n18170, n18173, n18174;
  wire n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182;
  wire n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192;
  wire n18193, n18194, n18197, n18198, n18199, n18200, n18201, n18202;
  wire n18203, n18204, n18205, n18206, n18209, n18210, n18211, n18212;
  wire n18213, n18214, n18215, n18216, n18217, n18218, n18221, n18222;
  wire n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230;
  wire n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240;
  wire n18241, n18242, n18245, n18246, n18247, n18248, n18249, n18250;
  wire n18251, n18252, n18253, n18254, n18257, n18258, n18259, n18260;
  wire n18261, n18262, n18263, n18264, n18265, n18266, n18269, n18270;
  wire n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278;
  wire n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288;
  wire n18289, n18290, n18291, n18292, n18295, n18296, n18297, n18298;
  wire n18299, n18300, n18301, n18302, n18305, n18306, n18307, n18308;
  wire n18309, n18310, n18311, n18312, n18313, n18314, n18317, n18318;
  wire n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326;
  wire n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336;
  wire n18337, n18338, n18341, n18342, n18343, n18344, n18345, n18346;
  wire n18347, n18348, n18349, n18350, n18353, n18354, n18355, n18356;
  wire n18357, n18358, n18359, n18360, n18361, n18362, n18365, n18366;
  wire n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374;
  wire n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384;
  wire n18385, n18388, n18389, n18390, n18391, n18392, n18393, n18394;
  wire n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404;
  wire n18409, n18413, n18414, n18415, n18416, n18417, n18422, n18423;
  wire n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431;
  wire n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442;
  wire n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450;
  wire n18451, n18452, n18453, n18454, n18457, n18458, n18459, n18460;
  wire n18461, n18462, n18463, n18464, n18465, n18466, n18469, n18470;
  wire n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478;
  wire n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488;
  wire n18489, n18490, n18493, n18494, n18495, n18496, n18497, n18498;
  wire n18499, n18500, n18501, n18502, n18505, n18506, n18507, n18508;
  wire n18509, n18510, n18511, n18512, n18513, n18514, n18517, n18518;
  wire n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526;
  wire n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536;
  wire n18537, n18538, n18541, n18542, n18543, n18544, n18545, n18546;
  wire n18547, n18548, n18549, n18550, n18553, n18554, n18555, n18556;
  wire n18557, n18558, n18559, n18560, n18561, n18562, n18565, n18566;
  wire n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574;
  wire n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584;
  wire n18585, n18586, n18589, n18590, n18591, n18592, n18593, n18594;
  wire n18595, n18596, n18597, n18598, n18601, n18602, n18603, n18604;
  wire n18605, n18606, n18607, n18608, n18609, n18610, n18613, n18614;
  wire n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622;
  wire n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632;
  wire n18633, n18634, n18637, n18638, n18639, n18640, n18641, n18642;
  wire n18643, n18644, n18645, n18646, n18649, n18650, n18651, n18652;
  wire n18653, n18654, n18655, n18656, n18657, n18658, n18661, n18662;
  wire n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670;
  wire n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680;
  wire n18681, n18682, n18685, n18686, n18687, n18688, n18689, n18690;
  wire n18691, n18692, n18693, n18694, n18697, n18698, n18699, n18700;
  wire n18701, n18702, n18703, n18704, n18705, n18706, n18709, n18710;
  wire n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718;
  wire n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728;
  wire n18729, n18730, n18733, n18734, n18735, n18736, n18737, n18738;
  wire n18739, n18740, n18741, n18742, n18745, n18746, n18747, n18748;
  wire n18749, n18750, n18751, n18752, n18753, n18754, n18757, n18758;
  wire n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766;
  wire n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776;
  wire n18777, n18778, n18781, n18782, n18783, n18784, n18785, n18786;
  wire n18787, n18788, n18789, n18790, n18793, n18794, n18795, n18796;
  wire n18797, n18798, n18799, n18800, n18801, n18802, n18805, n18806;
  wire n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814;
  wire n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824;
  wire n18825, n18826, n18829, n18830, n18831, n18832, n18833, n18834;
  wire n18835, n18836, n18837, n18838, n18841, n18842, n18843, n18844;
  wire n18845, n18846, n18847, n18848, n18849, n18850, n18853, n18854;
  wire n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862;
  wire n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872;
  wire n18873, n18874, n18877, n18878, n18879, n18880, n18881, n18882;
  wire n18883, n18884, n18885, n18886, n18889, n18890, n18891, n18892;
  wire n18893, n18894, n18895, n18896, n18897, n18898, n18901, n18902;
  wire n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910;
  wire n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920;
  wire n18921, n18922, n18925, n18926, n18927, n18928, n18929, n18930;
  wire n18931, n18932, n18933, n18934, n18937, n18938, n18939, n18940;
  wire n18941, n18942, n18943, n18944, n18945, n18946, n18949, n18950;
  wire n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958;
  wire n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968;
  wire n18969, n18970, n18971, n18972, n18975, n18976, n18977, n18978;
  wire n18979, n18980, n18981, n18982, n18985, n18986, n18987, n18988;
  wire n18989, n18990, n18991, n18992, n18993, n18994, n18997, n18998;
  wire n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006;
  wire n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016;
  wire n19017, n19018, n19021, n19022, n19023, n19024, n19025, n19026;
  wire n19027, n19028, n19029, n19030, n19033, n19034, n19035, n19036;
  wire n19037, n19038, n19039, n19040, n19041, n19042, n19045, n19046;
  wire n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19056;
  wire n19057, n19058, n19059, n19060, n19061, n19062, n19065, n19066;
  wire n19067, n19068, n19069, n19070, n19071, n19072, n19077, n19081;
  wire n19082, n19083, n19084, n19085, n19090, n19091, n19092, n19093;
  wire n19094, n19095, n19096, n19097, n19098, n19099, n19103, n19104;
  wire n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112;
  wire n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120;
  wire n19121, n19122, n19125, n19126, n19127, n19128, n19129, n19130;
  wire n19131, n19132, n19133, n19134, n19137, n19138, n19139, n19140;
  wire n19141, n19142, n19143, n19144, n19145, n19146, n19149, n19150;
  wire n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158;
  wire n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168;
  wire n19169, n19170, n19173, n19174, n19175, n19176, n19177, n19178;
  wire n19179, n19180, n19181, n19182, n19185, n19186, n19187, n19188;
  wire n19189, n19190, n19191, n19192, n19193, n19194, n19197, n19198;
  wire n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206;
  wire n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216;
  wire n19217, n19218, n19221, n19222, n19223, n19224, n19225, n19226;
  wire n19227, n19228, n19229, n19230, n19233, n19234, n19235, n19236;
  wire n19237, n19238, n19239, n19240, n19241, n19242, n19245, n19246;
  wire n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254;
  wire n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264;
  wire n19265, n19266, n19269, n19270, n19271, n19272, n19273, n19274;
  wire n19275, n19276, n19277, n19278, n19281, n19282, n19283, n19284;
  wire n19285, n19286, n19287, n19288, n19289, n19290, n19293, n19294;
  wire n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302;
  wire n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312;
  wire n19313, n19314, n19317, n19318, n19319, n19320, n19321, n19322;
  wire n19323, n19324, n19325, n19326, n19329, n19330, n19331, n19332;
  wire n19333, n19334, n19335, n19336, n19337, n19338, n19341, n19342;
  wire n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350;
  wire n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360;
  wire n19361, n19362, n19365, n19366, n19367, n19368, n19369, n19370;
  wire n19371, n19372, n19373, n19374, n19377, n19378, n19379, n19380;
  wire n19381, n19382, n19383, n19384, n19385, n19386, n19389, n19390;
  wire n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398;
  wire n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408;
  wire n19409, n19410, n19413, n19414, n19415, n19416, n19417, n19418;
  wire n19419, n19420, n19421, n19422, n19425, n19426, n19427, n19428;
  wire n19429, n19430, n19431, n19432, n19433, n19434, n19437, n19438;
  wire n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446;
  wire n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456;
  wire n19457, n19458, n19461, n19462, n19463, n19464, n19465, n19466;
  wire n19467, n19468, n19469, n19470, n19473, n19474, n19475, n19476;
  wire n19477, n19478, n19479, n19480, n19481, n19482, n19485, n19486;
  wire n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494;
  wire n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504;
  wire n19505, n19506, n19509, n19510, n19511, n19512, n19513, n19514;
  wire n19515, n19516, n19517, n19518, n19521, n19522, n19523, n19524;
  wire n19525, n19526, n19527, n19528, n19529, n19530, n19533, n19534;
  wire n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542;
  wire n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552;
  wire n19553, n19554, n19557, n19558, n19559, n19560, n19561, n19562;
  wire n19563, n19564, n19565, n19566, n19569, n19570, n19571, n19572;
  wire n19573, n19574, n19575, n19576, n19577, n19578, n19581, n19582;
  wire n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590;
  wire n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600;
  wire n19601, n19602, n19605, n19606, n19607, n19608, n19609, n19610;
  wire n19611, n19612, n19613, n19614, n19617, n19618, n19619, n19620;
  wire n19621, n19622, n19623, n19624, n19625, n19626, n19629, n19630;
  wire n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638;
  wire n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648;
  wire n19649, n19650, n19653, n19654, n19655, n19656, n19657, n19658;
  wire n19659, n19660, n19661, n19662, n19663, n19664, n19667, n19668;
  wire n19669, n19670, n19671, n19672, n19673, n19674, n19677, n19678;
  wire n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686;
  wire n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696;
  wire n19697, n19698, n19701, n19702, n19703, n19704, n19705, n19706;
  wire n19707, n19708, n19709, n19710, n19713, n19714, n19715, n19716;
  wire n19717, n19718, n19719, n19720, n19721, n19722, n19725, n19726;
  wire n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19736;
  wire n19737, n19738, n19739, n19740, n19741, n19742, n19745, n19746;
  wire n19747, n19748, n19749, n19750, n19751, n19752, n19757, n19761;
  wire n19762, n19763, n19764, n19765, n19770, n19771, n19772, n19773;
  wire n19774, n19775, n19776, n19777, n19778, n19779, n19783, n19784;
  wire n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792;
  wire n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800;
  wire n19801, n19802, n19805, n19806, n19807, n19808, n19809, n19810;
  wire n19811, n19812, n19813, n19814, n19817, n19818, n19819, n19820;
  wire n19821, n19822, n19823, n19824, n19825, n19826, n19829, n19830;
  wire n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838;
  wire n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848;
  wire n19849, n19850, n19853, n19854, n19855, n19856, n19857, n19858;
  wire n19859, n19860, n19861, n19862, n19865, n19866, n19867, n19868;
  wire n19869, n19870, n19871, n19872, n19873, n19874, n19877, n19878;
  wire n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886;
  wire n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896;
  wire n19897, n19898, n19901, n19902, n19903, n19904, n19905, n19906;
  wire n19907, n19908, n19909, n19910, n19913, n19914, n19915, n19916;
  wire n19917, n19918, n19919, n19920, n19921, n19922, n19925, n19926;
  wire n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934;
  wire n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944;
  wire n19945, n19946, n19949, n19950, n19951, n19952, n19953, n19954;
  wire n19955, n19956, n19957, n19958, n19961, n19962, n19963, n19964;
  wire n19965, n19966, n19967, n19968, n19969, n19970, n19973, n19974;
  wire n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982;
  wire n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992;
  wire n19993, n19994, n19997, n19998, n19999, n20000, n20001, n20002;
  wire n20003, n20004, n20005, n20006, n20009, n20010, n20011, n20012;
  wire n20013, n20014, n20015, n20016, n20017, n20018, n20021, n20022;
  wire n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030;
  wire n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040;
  wire n20041, n20042, n20045, n20046, n20047, n20048, n20049, n20050;
  wire n20051, n20052, n20053, n20054, n20057, n20058, n20059, n20060;
  wire n20061, n20062, n20063, n20064, n20065, n20066, n20069, n20070;
  wire n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078;
  wire n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088;
  wire n20089, n20090, n20093, n20094, n20095, n20096, n20097, n20098;
  wire n20099, n20100, n20101, n20102, n20105, n20106, n20107, n20108;
  wire n20109, n20110, n20111, n20112, n20113, n20114, n20117, n20118;
  wire n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126;
  wire n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136;
  wire n20137, n20138, n20141, n20142, n20143, n20144, n20145, n20146;
  wire n20147, n20148, n20149, n20150, n20153, n20154, n20155, n20156;
  wire n20157, n20158, n20159, n20160, n20161, n20162, n20165, n20166;
  wire n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174;
  wire n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184;
  wire n20185, n20186, n20189, n20190, n20191, n20192, n20193, n20194;
  wire n20195, n20196, n20197, n20198, n20201, n20202, n20203, n20204;
  wire n20205, n20206, n20207, n20208, n20209, n20210, n20213, n20214;
  wire n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222;
  wire n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232;
  wire n20233, n20234, n20237, n20238, n20239, n20240, n20241, n20242;
  wire n20243, n20244, n20245, n20246, n20249, n20250, n20251, n20252;
  wire n20253, n20254, n20255, n20256, n20257, n20258, n20261, n20262;
  wire n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270;
  wire n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280;
  wire n20281, n20282, n20285, n20286, n20287, n20288, n20289, n20290;
  wire n20291, n20292, n20293, n20294, n20297, n20298, n20299, n20300;
  wire n20301, n20302, n20303, n20304, n20305, n20306, n20309, n20310;
  wire n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318;
  wire n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328;
  wire n20329, n20330, n20333, n20334, n20335, n20336, n20337, n20338;
  wire n20339, n20340, n20341, n20342, n20345, n20346, n20347, n20348;
  wire n20349, n20350, n20351, n20352, n20353, n20354, n20357, n20358;
  wire n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366;
  wire n20367, n20368, n20371, n20372, n20373, n20374, n20375, n20376;
  wire n20377, n20378, n20381, n20382, n20383, n20384, n20385, n20386;
  wire n20387, n20388, n20389, n20390, n20393, n20394, n20395, n20396;
  wire n20397, n20398, n20399, n20400, n20401, n20402, n20405, n20406;
  wire n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414;
  wire n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424;
  wire n20425, n20428, n20429, n20430, n20431, n20432, n20433, n20434;
  wire n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444;
  wire n20449, n20453, n20454, n20455, n20456, n20457, n20462, n20463;
  wire n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471;
  wire n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482;
  wire n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490;
  wire n20491, n20492, n20493, n20494, n20497, n20498, n20499, n20500;
  wire n20501, n20502, n20503, n20504, n20505, n20506, n20509, n20510;
  wire n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518;
  wire n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528;
  wire n20529, n20530, n20533, n20534, n20535, n20536, n20537, n20538;
  wire n20539, n20540, n20541, n20542, n20545, n20546, n20547, n20548;
  wire n20549, n20550, n20551, n20552, n20553, n20554, n20557, n20558;
  wire n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566;
  wire n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576;
  wire n20577, n20578, n20581, n20582, n20583, n20584, n20585, n20586;
  wire n20587, n20588, n20589, n20590, n20593, n20594, n20595, n20596;
  wire n20597, n20598, n20599, n20600, n20601, n20602, n20605, n20606;
  wire n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614;
  wire n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624;
  wire n20625, n20626, n20629, n20630, n20631, n20632, n20633, n20634;
  wire n20635, n20636, n20637, n20638, n20641, n20642, n20643, n20644;
  wire n20645, n20646, n20647, n20648, n20649, n20650, n20653, n20654;
  wire n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662;
  wire n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672;
  wire n20673, n20674, n20677, n20678, n20679, n20680, n20681, n20682;
  wire n20683, n20684, n20685, n20686, n20689, n20690, n20691, n20692;
  wire n20693, n20694, n20695, n20696, n20697, n20698, n20701, n20702;
  wire n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710;
  wire n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720;
  wire n20721, n20722, n20725, n20726, n20727, n20728, n20729, n20730;
  wire n20731, n20732, n20733, n20734, n20737, n20738, n20739, n20740;
  wire n20741, n20742, n20743, n20744, n20745, n20746, n20749, n20750;
  wire n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758;
  wire n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768;
  wire n20769, n20770, n20773, n20774, n20775, n20776, n20777, n20778;
  wire n20779, n20780, n20781, n20782, n20785, n20786, n20787, n20788;
  wire n20789, n20790, n20791, n20792, n20793, n20794, n20797, n20798;
  wire n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806;
  wire n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816;
  wire n20817, n20818, n20821, n20822, n20823, n20824, n20825, n20826;
  wire n20827, n20828, n20829, n20830, n20833, n20834, n20835, n20836;
  wire n20837, n20838, n20839, n20840, n20841, n20842, n20845, n20846;
  wire n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854;
  wire n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864;
  wire n20865, n20866, n20869, n20870, n20871, n20872, n20873, n20874;
  wire n20875, n20876, n20877, n20878, n20881, n20882, n20883, n20884;
  wire n20885, n20886, n20887, n20888, n20889, n20890, n20893, n20894;
  wire n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902;
  wire n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912;
  wire n20913, n20914, n20917, n20918, n20919, n20920, n20921, n20922;
  wire n20923, n20924, n20925, n20926, n20929, n20930, n20931, n20932;
  wire n20933, n20934, n20935, n20936, n20937, n20938, n20941, n20942;
  wire n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950;
  wire n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960;
  wire n20961, n20962, n20965, n20966, n20967, n20968, n20969, n20970;
  wire n20971, n20972, n20973, n20974, n20977, n20978, n20979, n20980;
  wire n20981, n20982, n20983, n20984, n20985, n20986, n20989, n20990;
  wire n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998;
  wire n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008;
  wire n21009, n21010, n21013, n21014, n21015, n21016, n21017, n21018;
  wire n21019, n21020, n21021, n21022, n21025, n21026, n21027, n21028;
  wire n21029, n21030, n21031, n21032, n21033, n21034, n21037, n21038;
  wire n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046;
  wire n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056;
  wire n21057, n21058, n21061, n21062, n21063, n21064, n21065, n21066;
  wire n21067, n21068, n21069, n21070, n21073, n21074, n21075, n21076;
  wire n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084;
  wire n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094;
  wire n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104;
  wire n21105, n21106, n21109, n21110, n21111, n21112, n21113, n21114;
  wire n21115, n21116, n21117, n21118, n21121, n21122, n21123, n21124;
  wire n21125, n21126, n21127, n21128, n21129, n21132, n21133, n21134;
  wire n21135, n21136, n21137, n21138, n21141, n21142, n21143, n21144;
  wire n21145, n21146, n21147, n21148, n21149, n21151, n21152, n21153;
  wire n21154, n21155, n21160, n21161, n21162, n21163, n21164, n21165;
  wire n21166, n21167, n21168, n21169, n21172, n21173, n21174, n21175;
  wire n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183;
  wire n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191;
  wire n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201;
  wire n21202, n21203, n21206, n21207, n21208, n21209, n21210, n21211;
  wire n21212, n21213, n21214, n21215, n21218, n21219, n21220, n21221;
  wire n21222, n21223, n21224, n21225, n21226, n21227, n21230, n21231;
  wire n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239;
  wire n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249;
  wire n21250, n21251, n21254, n21255, n21256, n21257, n21258, n21259;
  wire n21260, n21261, n21262, n21263, n21266, n21267, n21268, n21269;
  wire n21270, n21271, n21272, n21273, n21274, n21275, n21278, n21279;
  wire n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287;
  wire n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297;
  wire n21298, n21299, n21302, n21303, n21304, n21305, n21306, n21307;
  wire n21308, n21309, n21310, n21311, n21314, n21315, n21316, n21317;
  wire n21318, n21319, n21320, n21321, n21322, n21323, n21326, n21327;
  wire n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335;
  wire n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345;
  wire n21346, n21347, n21350, n21351, n21352, n21353, n21354, n21355;
  wire n21356, n21357, n21358, n21359, n21362, n21363, n21364, n21365;
  wire n21366, n21367, n21368, n21369, n21370, n21371, n21374, n21375;
  wire n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383;
  wire n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393;
  wire n21394, n21395, n21398, n21399, n21400, n21401, n21402, n21403;
  wire n21404, n21405, n21406, n21407, n21410, n21411, n21412, n21413;
  wire n21414, n21415, n21416, n21417, n21418, n21419, n21422, n21423;
  wire n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431;
  wire n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441;
  wire n21442, n21443, n21446, n21447, n21448, n21449, n21450, n21451;
  wire n21452, n21453, n21454, n21455, n21458, n21459, n21460, n21461;
  wire n21462, n21463, n21464, n21465, n21466, n21467, n21470, n21471;
  wire n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479;
  wire n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489;
  wire n21490, n21491, n21494, n21495, n21496, n21497, n21498, n21499;
  wire n21500, n21501, n21502, n21503, n21506, n21507, n21508, n21509;
  wire n21510, n21511, n21512, n21513, n21514, n21515, n21518, n21519;
  wire n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527;
  wire n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537;
  wire n21538, n21539, n21542, n21543, n21544, n21545, n21546, n21547;
  wire n21548, n21549, n21550, n21551, n21554, n21555, n21556, n21557;
  wire n21558, n21559, n21560, n21561, n21562, n21563, n21566, n21567;
  wire n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575;
  wire n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585;
  wire n21586, n21587, n21590, n21591, n21592, n21593, n21594, n21595;
  wire n21596, n21597, n21598, n21599, n21602, n21603, n21604, n21605;
  wire n21606, n21607, n21608, n21609, n21610, n21611, n21614, n21615;
  wire n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623;
  wire n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633;
  wire n21634, n21635, n21638, n21639, n21640, n21641, n21642, n21643;
  wire n21644, n21645, n21646, n21647, n21650, n21651, n21652, n21653;
  wire n21654, n21655, n21656, n21657, n21658, n21659, n21662, n21663;
  wire n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671;
  wire n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681;
  wire n21682, n21683, n21686, n21687, n21688, n21689, n21690, n21691;
  wire n21692, n21693, n21694, n21695, n21698, n21699, n21700, n21701;
  wire n21702, n21703, n21704, n21705, n21706, n21707, n21710, n21711;
  wire n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719;
  wire n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729;
  wire n21730, n21731, n21734, n21735, n21736, n21737, n21738, n21739;
  wire n21740, n21741, n21742, n21743, n21746, n21747, n21748, n21749;
  wire n21750, n21751, n21752, n21753, n21754, n21755, n21758, n21759;
  wire n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767;
  wire n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777;
  wire n21778, n21779, n21782, n21783, n21784, n21785, n21786, n21787;
  wire n21788, n21789, n21790, n21791, n21794, n21795, n21796, n21797;
  wire n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805;
  wire n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815;
  wire n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825;
  wire n21826, n21827, n21830, n21831, n21832, n21833, n21834, n21835;
  wire n21836, n21837, n21838, n21841, n21842, n21843, n21844, n21845;
  wire n21846, n21847, n21850, n21851, n21852, n21853, n21854, n21855;
  wire n21856, n21857, n21858, n21860, n21861, n21862, n21863, n21864;
  wire n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875;
  wire n21876, n21877, n21880, n21881, n21882, n21883, n21884, n21885;
  wire n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893;
  wire n21894, n21895, n21896, n21897, n21898, n21899, n21902, n21903;
  wire n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911;
  wire n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921;
  wire n21922, n21923, n21926, n21927, n21928, n21929, n21930, n21931;
  wire n21932, n21933, n21934, n21935, n21938, n21939, n21940, n21941;
  wire n21942, n21943, n21944, n21945, n21946, n21947, n21950, n21951;
  wire n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959;
  wire n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969;
  wire n21970, n21971, n21974, n21975, n21976, n21977, n21978, n21979;
  wire n21980, n21981, n21982, n21983, n21986, n21987, n21988, n21989;
  wire n21990, n21991, n21992, n21993, n21994, n21995, n21998, n21999;
  wire n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007;
  wire n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017;
  wire n22018, n22019, n22022, n22023, n22024, n22025, n22026, n22027;
  wire n22028, n22029, n22030, n22031, n22034, n22035, n22036, n22037;
  wire n22038, n22039, n22040, n22041, n22042, n22043, n22046, n22047;
  wire n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055;
  wire n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065;
  wire n22066, n22067, n22070, n22071, n22072, n22073, n22074, n22075;
  wire n22076, n22077, n22078, n22079, n22082, n22083, n22084, n22085;
  wire n22086, n22087, n22088, n22089, n22090, n22091, n22094, n22095;
  wire n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103;
  wire n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113;
  wire n22114, n22115, n22118, n22119, n22120, n22121, n22122, n22123;
  wire n22124, n22125, n22126, n22127, n22130, n22131, n22132, n22133;
  wire n22134, n22135, n22136, n22137, n22138, n22139, n22142, n22143;
  wire n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151;
  wire n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161;
  wire n22162, n22163, n22166, n22167, n22168, n22169, n22170, n22171;
  wire n22172, n22173, n22174, n22175, n22178, n22179, n22180, n22181;
  wire n22182, n22183, n22184, n22185, n22186, n22187, n22190, n22191;
  wire n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199;
  wire n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209;
  wire n22210, n22211, n22214, n22215, n22216, n22217, n22218, n22219;
  wire n22220, n22221, n22222, n22223, n22226, n22227, n22228, n22229;
  wire n22230, n22231, n22232, n22233, n22234, n22235, n22238, n22239;
  wire n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247;
  wire n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257;
  wire n22258, n22259, n22262, n22263, n22264, n22265, n22266, n22267;
  wire n22268, n22269, n22270, n22271, n22274, n22275, n22276, n22277;
  wire n22278, n22279, n22280, n22281, n22282, n22283, n22286, n22287;
  wire n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295;
  wire n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305;
  wire n22306, n22307, n22310, n22311, n22312, n22313, n22314, n22315;
  wire n22316, n22317, n22318, n22319, n22322, n22323, n22324, n22325;
  wire n22326, n22327, n22328, n22329, n22330, n22331, n22334, n22335;
  wire n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343;
  wire n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353;
  wire n22354, n22355, n22358, n22359, n22360, n22361, n22362, n22363;
  wire n22364, n22365, n22366, n22367, n22370, n22371, n22372, n22373;
  wire n22374, n22375, n22376, n22377, n22378, n22379, n22382, n22383;
  wire n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391;
  wire n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401;
  wire n22402, n22403, n22406, n22407, n22408, n22409, n22410, n22411;
  wire n22412, n22413, n22414, n22415, n22418, n22419, n22420, n22421;
  wire n22422, n22423, n22424, n22425, n22426, n22427, n22430, n22431;
  wire n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439;
  wire n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449;
  wire n22450, n22451, n22454, n22455, n22456, n22457, n22458, n22459;
  wire n22460, n22461, n22462, n22463, n22466, n22467, n22468, n22469;
  wire n22470, n22471, n22472, n22473, n22474, n22475, n22478, n22479;
  wire n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487;
  wire n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497;
  wire n22498, n22499, n22502, n22503, n22504, n22505, n22506, n22507;
  wire n22508, n22509, n22510, n22511, n22514, n22515, n22516, n22517;
  wire n22518, n22519, n22520, n22521, n22522, n22523, n22526, n22527;
  wire n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535;
  wire n22536, n22537, n22540, n22541, n22542, n22543, n22544, n22545;
  wire n22546, n22547, n22550, n22551, n22552, n22553, n22554, n22555;
  wire n22556, n22557, n22558, n22561, n22562, n22563, n22564, n22565;
  wire n22566, n22567, n22570, n22571, n22572, n22573, n22574, n22575;
  wire n22576, n22577, n22578, n22580, n22581, n22582, n22583, n22584;
  wire n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595;
  wire n22596, n22597, n22600, n22601, n22602, n22603, n22604, n22605;
  wire n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613;
  wire n22614, n22615, n22616, n22617, n22618, n22619, n22622, n22623;
  wire n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631;
  wire n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641;
  wire n22642, n22643, n22646, n22647, n22648, n22649, n22650, n22651;
  wire n22652, n22653, n22654, n22655, n22658, n22659, n22660, n22661;
  wire n22662, n22663, n22664, n22665, n22666, n22667, n22670, n22671;
  wire n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679;
  wire n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689;
  wire n22690, n22691, n22694, n22695, n22696, n22697, n22698, n22699;
  wire n22700, n22701, n22702, n22703, n22706, n22707, n22708, n22709;
  wire n22710, n22711, n22712, n22713, n22714, n22715, n22718, n22719;
  wire n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727;
  wire n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737;
  wire n22738, n22739, n22742, n22743, n22744, n22745, n22746, n22747;
  wire n22748, n22749, n22750, n22751, n22754, n22755, n22756, n22757;
  wire n22758, n22759, n22760, n22761, n22762, n22763, n22766, n22767;
  wire n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775;
  wire n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785;
  wire n22786, n22787, n22790, n22791, n22792, n22793, n22794, n22795;
  wire n22796, n22797, n22798, n22799, n22802, n22803, n22804, n22805;
  wire n22806, n22807, n22808, n22809, n22810, n22811, n22814, n22815;
  wire n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823;
  wire n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833;
  wire n22834, n22835, n22838, n22839, n22840, n22841, n22842, n22843;
  wire n22844, n22845, n22846, n22847, n22850, n22851, n22852, n22853;
  wire n22854, n22855, n22856, n22857, n22858, n22859, n22862, n22863;
  wire n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871;
  wire n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881;
  wire n22882, n22883, n22886, n22887, n22888, n22889, n22890, n22891;
  wire n22892, n22893, n22894, n22895, n22898, n22899, n22900, n22901;
  wire n22902, n22903, n22904, n22905, n22906, n22907, n22910, n22911;
  wire n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919;
  wire n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929;
  wire n22930, n22931, n22934, n22935, n22936, n22937, n22938, n22939;
  wire n22940, n22941, n22942, n22943, n22946, n22947, n22948, n22949;
  wire n22950, n22951, n22952, n22953, n22954, n22955, n22958, n22959;
  wire n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967;
  wire n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977;
  wire n22978, n22979, n22982, n22983, n22984, n22985, n22986, n22987;
  wire n22988, n22989, n22990, n22991, n22994, n22995, n22996, n22997;
  wire n22998, n22999, n23000, n23001, n23002, n23003, n23006, n23007;
  wire n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015;
  wire n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025;
  wire n23026, n23027, n23030, n23031, n23032, n23033, n23034, n23035;
  wire n23036, n23037, n23038, n23039, n23042, n23043, n23044, n23045;
  wire n23046, n23047, n23048, n23049, n23050, n23051, n23054, n23055;
  wire n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063;
  wire n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073;
  wire n23074, n23075, n23078, n23079, n23080, n23081, n23082, n23083;
  wire n23084, n23085, n23086, n23087, n23090, n23091, n23092, n23093;
  wire n23094, n23095, n23096, n23097, n23098, n23099, n23102, n23103;
  wire n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111;
  wire n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121;
  wire n23122, n23123, n23126, n23127, n23128, n23129, n23130, n23131;
  wire n23132, n23133, n23134, n23135, n23138, n23139, n23140, n23141;
  wire n23142, n23143, n23144, n23145, n23146, n23147, n23150, n23151;
  wire n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159;
  wire n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169;
  wire n23170, n23171, n23174, n23175, n23176, n23177, n23178, n23179;
  wire n23180, n23181, n23182, n23183, n23186, n23187, n23188, n23189;
  wire n23190, n23191, n23192, n23193, n23194, n23195, n23198, n23199;
  wire n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207;
  wire n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217;
  wire n23218, n23219, n23222, n23223, n23224, n23225, n23226, n23227;
  wire n23228, n23229, n23230, n23231, n23234, n23235, n23236, n23237;
  wire n23238, n23239, n23240, n23241, n23242, n23243, n23246, n23247;
  wire n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255;
  wire n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265;
  wire n23266, n23267, n23270, n23271, n23272, n23273, n23274, n23275;
  wire n23276, n23277, n23278, n23279, n23280, n23281, n23284, n23285;
  wire n23286, n23287, n23288, n23289, n23290, n23293, n23294, n23295;
  wire n23296, n23297, n23298, n23299, n23302, n23303, n23304, n23305;
  wire n23306, n23307, n23308, n23309, n23310, n23314, n23315, n23316;
  wire n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23327;
  wire n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335;
  wire n23336, n23339, n23340, n23341, n23342, n23343, n23344, n23345;
  wire n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353;
  wire n23354, n23355, n23356, n23357, n23358, n23361, n23362, n23363;
  wire n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23373;
  wire n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381;
  wire n23382, n23385, n23386, n23387, n23388, n23389, n23390, n23391;
  wire n23392, n23393, n23394, n23397, n23398, n23399, n23400, n23401;
  wire n23402, n23403, n23404, n23405, n23406, n23409, n23410, n23411;
  wire n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23421;
  wire n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429;
  wire n23430, n23433, n23434, n23435, n23436, n23437, n23438, n23439;
  wire n23440, n23441, n23442, n23445, n23446, n23447, n23448, n23449;
  wire n23450, n23451, n23452, n23453, n23454, n23457, n23458, n23459;
  wire n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23469;
  wire n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477;
  wire n23478, n23481, n23482, n23483, n23484, n23485, n23486, n23487;
  wire n23488, n23489, n23490, n23493, n23494, n23495, n23496, n23497;
  wire n23498, n23499, n23500, n23501, n23502, n23505, n23506, n23507;
  wire n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23517;
  wire n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525;
  wire n23526, n23529, n23530, n23531, n23532, n23533, n23534, n23535;
  wire n23536, n23537, n23538, n23541, n23542, n23543, n23544, n23545;
  wire n23546, n23547, n23548, n23549, n23550, n23553, n23554, n23555;
  wire n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23565;
  wire n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573;
  wire n23574, n23577, n23578, n23579, n23580, n23581, n23582, n23583;
  wire n23584, n23585, n23586, n23589, n23590, n23591, n23592, n23593;
  wire n23594, n23595, n23596, n23597, n23598, n23601, n23602, n23603;
  wire n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23613;
  wire n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621;
  wire n23622, n23625, n23626, n23627, n23628, n23629, n23630, n23631;
  wire n23632, n23633, n23634, n23637, n23638, n23639, n23640, n23641;
  wire n23642, n23643, n23644, n23645, n23646, n23649, n23650, n23651;
  wire n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23661;
  wire n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669;
  wire n23670, n23673, n23674, n23675, n23676, n23677, n23678, n23679;
  wire n23680, n23681, n23682, n23685, n23686, n23687, n23688, n23689;
  wire n23690, n23691, n23692, n23693, n23694, n23697, n23698, n23699;
  wire n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23709;
  wire n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717;
  wire n23718, n23721, n23722, n23723, n23724, n23725, n23726, n23727;
  wire n23728, n23729, n23730, n23733, n23734, n23735, n23736, n23737;
  wire n23738, n23739, n23740, n23741, n23742, n23745, n23746, n23747;
  wire n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23757;
  wire n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765;
  wire n23766, n23769, n23770, n23771, n23772, n23773, n23774, n23775;
  wire n23776, n23777, n23778, n23781, n23782, n23783, n23784, n23785;
  wire n23786, n23787, n23788, n23789, n23790, n23793, n23794, n23795;
  wire n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23805;
  wire n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813;
  wire n23814, n23817, n23818, n23819, n23820, n23821, n23822, n23823;
  wire n23824, n23825, n23826, n23829, n23830, n23831, n23832, n23833;
  wire n23834, n23835, n23836, n23837, n23838, n23841, n23842, n23843;
  wire n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23853;
  wire n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861;
  wire n23862, n23865, n23866, n23867, n23868, n23869, n23870, n23871;
  wire n23872, n23873, n23874, n23877, n23878, n23879, n23880, n23881;
  wire n23882, n23883, n23884, n23885, n23886, n23889, n23890, n23891;
  wire n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23901;
  wire n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909;
  wire n23910, n23913, n23914, n23915, n23916, n23917, n23918, n23919;
  wire n23920, n23921, n23922, n23925, n23926, n23927, n23928, n23929;
  wire n23930, n23931, n23932, n23933, n23934, n23937, n23938, n23939;
  wire n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23949;
  wire n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957;
  wire n23958, n23961, n23962, n23963, n23964, n23965, n23966, n23967;
  wire n23968, n23969, n23970, n23973, n23974, n23975, n23976, n23977;
  wire n23978, n23979, n23980, n23981, n23982, n23985, n23986, n23987;
  wire n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23997;
  wire n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005;
  wire n24006, n24009, n24010, n24011, n24012, n24013, n24014, n24015;
  wire n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023;
  wire n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033;
  wire n24034, n24037, n24038, n24039, n24040, n24041, n24042, n24043;
  wire n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053;
  wire n24054, n24056, n24057, n24058, n24061, n24062, n24063, n24064;
  wire n24065, n24068, n24069, n24070, n24071, n24072, n24075, n24076;
  wire n24077, n24078, n24079, n24082, n24083, n24084, n24085, n24086;
  wire n24089, n24090, n24091, n24092, n24093, n24096, n24097, n24098;
  wire n24099, n24100, n24103, n24104, n24105, n24106, n24107, n24110;
  wire n24111, n24112, n24113, n24114, n24117, n24118, n24119, n24120;
  wire n24121, n24124, n24125, n24126, n24127, n24128, n24131, n24132;
  wire n24133, n24134, n24135, n24138, n24139, n24140, n24141, n24142;
  wire n24145, n24146, n24147, n24148, n24149, n24152, n24153, n24154;
  wire n24155, n24156, n24159, n24160, n24161, n24162, n24163, n24166;
  wire n24167, n24168, n24169, n24170, n24173, n24174, n24175, n24176;
  wire n24177, n24180, n24181, n24182, n24183, n24184, n24187, n24188;
  wire n24189, n24190, n24191, n24194, n24195, n24196, n24197, n24198;
  wire n24201, n24202, n24203, n24204, n24205, n24208, n24209, n24210;
  wire n24211, n24212, n24215, n24216, n24217, n24218, n24219, n24222;
  wire n24223, n24224, n24225, n24226, n24229, n24230, n24231, n24232;
  wire n24233, n24236, n24237, n24238, n24239, n24240, n24243, n24244;
  wire n24245, n24246, n24247, n24250, n24251, n24254, n24255, n24256;
  wire n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264;
  wire n24265, n24268, n24269, n24270, n24271, n24272, n24273, n24274;
  wire n24275, n24276, n24277, n24280, n24281, n24282, n24283, n24284;
  wire n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292;
  wire n24293, n24294, n24295, n24296, n24297, n24298, n24301, n24302;
  wire n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310;
  wire n24311, n24312, n24313, n24314, n24315, n24318, n24319, n24320;
  wire n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328;
  wire n24329, n24330, n24331, n24332, n24335, n24336, n24337, n24338;
  wire n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346;
  wire n24347, n24348, n24349, n24352, n24353, n24354, n24355, n24356;
  wire n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364;
  wire n24365, n24366, n24369, n24370, n24371, n24372, n24373, n24374;
  wire n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382;
  wire n24383, n24386, n24387, n24388, n24389, n24390, n24391, n24392;
  wire n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400;
  wire n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410;
  wire n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24420;
  wire n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428;
  wire n24429, n24430, n24431, n24432, n24433, n24434, n24437, n24438;
  wire n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446;
  wire n24447, n24448, n24449, n24450, n24451, n24454, n24455, n24456;
  wire n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464;
  wire n24465, n24466, n24467, n24468, n24471, n24472, n24473, n24474;
  wire n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482;
  wire n24483, n24484, n24485, n24488, n24489, n24490, n24491, n24492;
  wire n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500;
  wire n24501, n24502, n24505, n24506, n24507, n24508, n24509, n24510;
  wire n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518;
  wire n24519, n24522, n24523, n24524, n24525, n24526, n24527, n24528;
  wire n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536;
  wire n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546;
  wire n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24556;
  wire n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564;
  wire n24565, n24566, n24567, n24568, n24569, n24570, n24573, n24574;
  wire n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582;
  wire n24583, n24584, n24585, n24586, n24587, n24590, n24591, n24592;
  wire n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600;
  wire n24601, n24602, n24603, n24604, n24607, n24608, n24609, n24610;
  wire n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618;
  wire n24619, n24620, n24621, n24624, n24625, n24626, n24627, n24628;
  wire n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636;
  wire n24637, n24638, n24641, n24642, n24643, n24644, n24645, n24646;
  wire n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654;
  wire n24655, n24658, n24659, n24660, n24661, n24662, n24663, n24664;
  wire n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672;
  wire n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682;
  wire n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24692;
  wire n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700;
  wire n24701, n24702, n24703, n24704, n24705, n24706, n24709, n24710;
  wire n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718;
  wire n24719, n24720, n24721, n24722, n24723, n24726, n24727, n24728;
  wire n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736;
  wire n24737, n24738, n24739, n24740, n24743, n24744, n24745, n24746;
  wire n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754;
  wire n24755, n24756, n24757, n24760, n24761, n24762, n24763, n24764;
  wire n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772;
  wire n24773, n24774, n24777, n24778, n24779, n24780, n24781, n24782;
  wire n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790;
  wire n24791, n24794, n24795, n24796, n24797, n24801, n24802, n24803;
  wire n24804, n24805, n24806, n24807, n24808, n24809, n_6, n_7;
  wire n_8, n_9, n_13, n_14, n_15, n_16, n_17, n_18;
  wire n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26;
  wire n_27, n_28, n_29, n_33, n_34, n_35, n_36, n_37;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_91, n_92, n_93;
  wire n_94, n_95, n_96, n_97, n_98, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492;
  wire n_493, n_494, n_495, n_497, n_498, n_499, n_500, n_501;
  wire n_502, n_503, n_504, n_505, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
  wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662;
  wire n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686;
  wire n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694;
  wire n_695, n_697, n_698, n_699, n_700, n_701, n_702, n_703;
  wire n_704, n_705, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  wire n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787;
  wire n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_833, n_834, n_835, n_836, n_837, n_838, n_839, n_840;
  wire n_841, n_842, n_843, n_844, n_845, n_846, n_847, n_848;
  wire n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864;
  wire n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872;
  wire n_873, n_874, n_875, n_876, n_877, n_878, n_879, n_880;
  wire n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_893, n_894, n_895, n_896;
  wire n_897, n_898, n_899, n_900, n_901, n_902, n_903, n_904;
  wire n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937;
  wire n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949;
  wire n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957;
  wire n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965;
  wire n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973;
  wire n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981;
  wire n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989;
  wire n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997;
  wire n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005;
  wire n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013;
  wire n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021;
  wire n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029;
  wire n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037;
  wire n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045;
  wire n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053;
  wire n_1054, n_1055, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062;
  wire n_1063, n_1064, n_1065, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082;
  wire n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
  wire n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154;
  wire n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186;
  wire n_1187, n_1188, n_1189, n_1190, n_1191, n_1193, n_1194, n_1195;
  wire n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1225, n_1226, n_1227, n_1228, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272;
  wire n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280;
  wire n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288;
  wire n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320;
  wire n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1337;
  wire n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
  wire n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437;
  wire n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469;
  wire n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477;
  wire n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485;
  wire n_1486, n_1487, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494;
  wire n_1495, n_1496, n_1497, n_1502, n_1503, n_1504, n_1505, n_1506;
  wire n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522;
  wire n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530;
  wire n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538;
  wire n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546;
  wire n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554;
  wire n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562;
  wire n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570;
  wire n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586;
  wire n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594;
  wire n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602;
  wire n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610;
  wire n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618;
  wire n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626;
  wire n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634;
  wire n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642;
  wire n_1643, n_1644, n_1645, n_1646, n_1647, n_1649, n_1650, n_1651;
  wire n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1662, n_1663;
  wire n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671;
  wire n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679;
  wire n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711;
  wire n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719;
  wire n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727;
  wire n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844;
  wire n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852;
  wire n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860;
  wire n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868;
  wire n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884;
  wire n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892;
  wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
  wire n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916;
  wire n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924;
  wire n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932;
  wire n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940;
  wire n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948;
  wire n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956;
  wire n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964;
  wire n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972;
  wire n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980;
  wire n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988;
  wire n_1989, n_1990, n_1991, n_1993, n_1994, n_1995, n_1996, n_1997;
  wire n_1998, n_1999, n_2000, n_2001, n_2006, n_2007, n_2008, n_2009;
  wire n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017;
  wire n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025;
  wire n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057;
  wire n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073;
  wire n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081;
  wire n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089;
  wire n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097;
  wire n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105;
  wire n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113;
  wire n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121;
  wire n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129;
  wire n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137;
  wire n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145;
  wire n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153;
  wire n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161;
  wire n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2190;
  wire n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198;
  wire n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206;
  wire n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214;
  wire n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222;
  wire n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230;
  wire n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238;
  wire n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246;
  wire n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254;
  wire n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262;
  wire n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270;
  wire n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278;
  wire n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286;
  wire n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294;
  wire n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302;
  wire n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310;
  wire n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318;
  wire n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326;
  wire n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334;
  wire n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342;
  wire n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350;
  wire n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358;
  wire n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366;
  wire n_2367, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375;
  wire n_2376, n_2377, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387;
  wire n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395;
  wire n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403;
  wire n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411;
  wire n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419;
  wire n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435;
  wire n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443;
  wire n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451;
  wire n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459;
  wire n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467;
  wire n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475;
  wire n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483;
  wire n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491;
  wire n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499;
  wire n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507;
  wire n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515;
  wire n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523;
  wire n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531;
  wire n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539;
  wire n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547;
  wire n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555;
  wire n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563;
  wire n_2564, n_2565, n_2566, n_2567, n_2569, n_2570, n_2571, n_2572;
  wire n_2573, n_2574, n_2575, n_2576, n_2577, n_2582, n_2583, n_2584;
  wire n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592;
  wire n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600;
  wire n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608;
  wire n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616;
  wire n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624;
  wire n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632;
  wire n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640;
  wire n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648;
  wire n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656;
  wire n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664;
  wire n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
  wire n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680;
  wire n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688;
  wire n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696;
  wire n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704;
  wire n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712;
  wire n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744;
  wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
  wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
  wire n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768;
  wire n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2777;
  wire n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785;
  wire n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797;
  wire n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805;
  wire n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813;
  wire n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821;
  wire n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829;
  wire n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837;
  wire n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845;
  wire n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853;
  wire n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861;
  wire n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869;
  wire n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877;
  wire n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885;
  wire n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893;
  wire n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901;
  wire n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909;
  wire n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917;
  wire n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925;
  wire n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933;
  wire n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941;
  wire n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949;
  wire n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957;
  wire n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965;
  wire n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973;
  wire n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981;
  wire n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989;
  wire n_2990, n_2991, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998;
  wire n_2999, n_3000, n_3001, n_3006, n_3007, n_3008, n_3009, n_3010;
  wire n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018;
  wire n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026;
  wire n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034;
  wire n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042;
  wire n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050;
  wire n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058;
  wire n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066;
  wire n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074;
  wire n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082;
  wire n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090;
  wire n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098;
  wire n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106;
  wire n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114;
  wire n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122;
  wire n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130;
  wire n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138;
  wire n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146;
  wire n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154;
  wire n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162;
  wire n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170;
  wire n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178;
  wire n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186;
  wire n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194;
  wire n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202;
  wire n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210;
  wire n_3211, n_3212, n_3213, n_3214, n_3215, n_3217, n_3218, n_3219;
  wire n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3230, n_3231;
  wire n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239;
  wire n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247;
  wire n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255;
  wire n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263;
  wire n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271;
  wire n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279;
  wire n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287;
  wire n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295;
  wire n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303;
  wire n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311;
  wire n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319;
  wire n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327;
  wire n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335;
  wire n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343;
  wire n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351;
  wire n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359;
  wire n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367;
  wire n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375;
  wire n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383;
  wire n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391;
  wire n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399;
  wire n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407;
  wire n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415;
  wire n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423;
  wire n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431;
  wire n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439;
  wire n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447;
  wire n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456;
  wire n_3457, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468;
  wire n_3469, n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476;
  wire n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484;
  wire n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492;
  wire n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500;
  wire n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508;
  wire n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516;
  wire n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524;
  wire n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532;
  wire n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540;
  wire n_3541, n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548;
  wire n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556;
  wire n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564;
  wire n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572;
  wire n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580;
  wire n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588;
  wire n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596;
  wire n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604;
  wire n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612;
  wire n_3613, n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620;
  wire n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628;
  wire n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636;
  wire n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644;
  wire n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652;
  wire n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660;
  wire n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668;
  wire n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676;
  wire n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684;
  wire n_3685, n_3686, n_3687, n_3689, n_3690, n_3691, n_3692, n_3693;
  wire n_3694, n_3695, n_3696, n_3697, n_3702, n_3703, n_3704, n_3705;
  wire n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713;
  wire n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721;
  wire n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729;
  wire n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737;
  wire n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745;
  wire n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753;
  wire n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761;
  wire n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769;
  wire n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777;
  wire n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785;
  wire n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793;
  wire n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801;
  wire n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809;
  wire n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817;
  wire n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825;
  wire n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833;
  wire n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841;
  wire n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849;
  wire n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857;
  wire n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865;
  wire n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873;
  wire n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881;
  wire n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889;
  wire n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897;
  wire n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905;
  wire n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913;
  wire n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921;
  wire n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929;
  wire n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3937, n_3938;
  wire n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3950;
  wire n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958;
  wire n_3959, n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966;
  wire n_3967, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974;
  wire n_3975, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981, n_3982;
  wire n_3983, n_3984, n_3985, n_3986, n_3987, n_3988, n_3989, n_3990;
  wire n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3998;
  wire n_3999, n_4000, n_4001, n_4002, n_4003, n_4004, n_4005, n_4006;
  wire n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014;
  wire n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022;
  wire n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4029, n_4030;
  wire n_4031, n_4032, n_4033, n_4034, n_4035, n_4036, n_4037, n_4038;
  wire n_4039, n_4040, n_4041, n_4042, n_4043, n_4044, n_4045, n_4046;
  wire n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054;
  wire n_4055, n_4056, n_4057, n_4058, n_4059, n_4060, n_4061, n_4062;
  wire n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4070;
  wire n_4071, n_4072, n_4073, n_4074, n_4075, n_4076, n_4077, n_4078;
  wire n_4079, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086;
  wire n_4087, n_4088, n_4089, n_4090, n_4091, n_4092, n_4093, n_4094;
  wire n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102;
  wire n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110;
  wire n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118;
  wire n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126;
  wire n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134;
  wire n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142;
  wire n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150;
  wire n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158;
  wire n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166;
  wire n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174;
  wire n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182;
  wire n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190;
  wire n_4191, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4199;
  wire n_4200, n_4201, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211;
  wire n_4212, n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219;
  wire n_4220, n_4221, n_4222, n_4223, n_4224, n_4225, n_4226, n_4227;
  wire n_4228, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235;
  wire n_4236, n_4237, n_4238, n_4239, n_4240, n_4241, n_4242, n_4243;
  wire n_4244, n_4245, n_4246, n_4247, n_4248, n_4249, n_4250, n_4251;
  wire n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258, n_4259;
  wire n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267;
  wire n_4268, n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275;
  wire n_4276, n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283;
  wire n_4284, n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291;
  wire n_4292, n_4293, n_4294, n_4295, n_4296, n_4297, n_4298, n_4299;
  wire n_4300, n_4301, n_4302, n_4303, n_4304, n_4305, n_4306, n_4307;
  wire n_4308, n_4309, n_4310, n_4311, n_4312, n_4313, n_4314, n_4315;
  wire n_4316, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323;
  wire n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4331;
  wire n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339;
  wire n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4347;
  wire n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355;
  wire n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363;
  wire n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371;
  wire n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379;
  wire n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387;
  wire n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395;
  wire n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403;
  wire n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411;
  wire n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419;
  wire n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427;
  wire n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4435;
  wire n_4436, n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4443;
  wire n_4444, n_4445, n_4446, n_4447, n_4448, n_4449, n_4450, n_4451;
  wire n_4452, n_4453, n_4454, n_4455, n_4457, n_4458, n_4459, n_4460;
  wire n_4461, n_4462, n_4463, n_4464, n_4465, n_4470, n_4471, n_4472;
  wire n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4479, n_4480;
  wire n_4481, n_4482, n_4483, n_4484, n_4485, n_4486, n_4487, n_4488;
  wire n_4489, n_4490, n_4491, n_4492, n_4494, n_4495, n_4496, n_4497;
  wire n_4498, n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4505;
  wire n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513;
  wire n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521;
  wire n_4522, n_4523, n_4524, n_4525, n_4526, n_4527, n_4528, n_4529;
  wire n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537;
  wire n_4538, n_4539, n_4540, n_4541, n_4542, n_4543, n_4544, n_4545;
  wire n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552, n_4553;
  wire n_4554, n_4555, n_4556, n_4557, n_4558, n_4559, n_4560, n_4561;
  wire n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569;
  wire n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4576, n_4577;
  wire n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4585;
  wire n_4586, n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593;
  wire n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601;
  wire n_4602, n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609;
  wire n_4610, n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617;
  wire n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625;
  wire n_4626, n_4627, n_4628, n_4629, n_4630, n_4631, n_4632, n_4633;
  wire n_4634, n_4635, n_4636, n_4637, n_4638, n_4639, n_4640, n_4641;
  wire n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649;
  wire n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657;
  wire n_4658, n_4659, n_4660, n_4661, n_4662, n_4663, n_4664, n_4665;
  wire n_4666, n_4667, n_4668, n_4669, n_4670, n_4671, n_4672, n_4673;
  wire n_4674, n_4675, n_4676, n_4677, n_4678, n_4679, n_4680, n_4681;
  wire n_4682, n_4683, n_4684, n_4685, n_4686, n_4687, n_4688, n_4689;
  wire n_4690, n_4691, n_4692, n_4693, n_4694, n_4695, n_4696, n_4697;
  wire n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705;
  wire n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713;
  wire n_4714, n_4715, n_4716, n_4717, n_4718, n_4719, n_4720, n_4721;
  wire n_4722, n_4723, n_4724, n_4725, n_4726, n_4727, n_4729, n_4730;
  wire n_4731, n_4732, n_4733, n_4734, n_4735, n_4736, n_4737, n_4742;
  wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
  wire n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758;
  wire n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766;
  wire n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774;
  wire n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782;
  wire n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790;
  wire n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798;
  wire n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806;
  wire n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814;
  wire n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822;
  wire n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830;
  wire n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838;
  wire n_4839, n_4840, n_4841, n_4842, n_4843, n_4844, n_4845, n_4846;
  wire n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854;
  wire n_4855, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862;
  wire n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870;
  wire n_4871, n_4872, n_4873, n_4874, n_4875, n_4876, n_4877, n_4878;
  wire n_4879, n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886;
  wire n_4887, n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894;
  wire n_4895, n_4896, n_4897, n_4898, n_4899, n_4900, n_4901, n_4902;
  wire n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4910;
  wire n_4911, n_4912, n_4913, n_4914, n_4915, n_4916, n_4917, n_4918;
  wire n_4919, n_4920, n_4921, n_4922, n_4923, n_4924, n_4925, n_4926;
  wire n_4927, n_4928, n_4929, n_4930, n_4931, n_4932, n_4933, n_4934;
  wire n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942;
  wire n_4943, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950;
  wire n_4951, n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4958;
  wire n_4959, n_4960, n_4961, n_4962, n_4963, n_4964, n_4965, n_4966;
  wire n_4967, n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974;
  wire n_4975, n_4976, n_4977, n_4978, n_4979, n_4980, n_4981, n_4982;
  wire n_4983, n_4984, n_4985, n_4986, n_4987, n_4988, n_4989, n_4990;
  wire n_4991, n_4992, n_4993, n_4994, n_4995, n_4996, n_4997, n_4998;
  wire n_4999, n_5000, n_5001, n_5002, n_5003, n_5004, n_5005, n_5006;
  wire n_5007, n_5009, n_5010, n_5011, n_5012, n_5013, n_5014, n_5015;
  wire n_5016, n_5017, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027;
  wire n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035;
  wire n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043;
  wire n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051;
  wire n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059;
  wire n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067;
  wire n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075;
  wire n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083;
  wire n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091;
  wire n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099;
  wire n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107;
  wire n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115;
  wire n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123;
  wire n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131;
  wire n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139;
  wire n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147;
  wire n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155;
  wire n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163;
  wire n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171;
  wire n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179;
  wire n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187;
  wire n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195;
  wire n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203;
  wire n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211;
  wire n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219;
  wire n_5220, n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227;
  wire n_5228, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235;
  wire n_5236, n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243;
  wire n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251;
  wire n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259;
  wire n_5260, n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267;
  wire n_5268, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275;
  wire n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283;
  wire n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291;
  wire n_5292, n_5293, n_5294, n_5295, n_5297, n_5298, n_5299, n_5300;
  wire n_5301, n_5302, n_5303, n_5304, n_5305, n_5310, n_5311, n_5312;
  wire n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320;
  wire n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328;
  wire n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336;
  wire n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344;
  wire n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352;
  wire n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360;
  wire n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368;
  wire n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376;
  wire n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384;
  wire n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392;
  wire n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400;
  wire n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408;
  wire n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416;
  wire n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424;
  wire n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432;
  wire n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440;
  wire n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448;
  wire n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456;
  wire n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464;
  wire n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472;
  wire n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480;
  wire n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488;
  wire n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496;
  wire n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504;
  wire n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512;
  wire n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520;
  wire n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528;
  wire n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536;
  wire n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544;
  wire n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552;
  wire n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560;
  wire n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
  wire n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576;
  wire n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584;
  wire n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5593;
  wire n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600, n_5601;
  wire n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613;
  wire n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620, n_5621;
  wire n_5622, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629;
  wire n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637;
  wire n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645;
  wire n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653;
  wire n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661;
  wire n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669;
  wire n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677;
  wire n_5678, n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685;
  wire n_5686, n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693;
  wire n_5694, n_5695, n_5696, n_5697, n_5698, n_5699, n_5700, n_5701;
  wire n_5702, n_5703, n_5704, n_5705, n_5706, n_5707, n_5708, n_5709;
  wire n_5710, n_5711, n_5712, n_5713, n_5714, n_5715, n_5716, n_5717;
  wire n_5718, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725;
  wire n_5726, n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733;
  wire n_5734, n_5735, n_5736, n_5737, n_5738, n_5739, n_5740, n_5741;
  wire n_5742, n_5743, n_5744, n_5745, n_5746, n_5747, n_5748, n_5749;
  wire n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756, n_5757;
  wire n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764, n_5765;
  wire n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772, n_5773;
  wire n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780, n_5781;
  wire n_5782, n_5783, n_5784, n_5785, n_5786, n_5787, n_5788, n_5789;
  wire n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797;
  wire n_5798, n_5799, n_5800, n_5801, n_5802, n_5803, n_5804, n_5805;
  wire n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5812, n_5813;
  wire n_5814, n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821;
  wire n_5822, n_5823, n_5824, n_5825, n_5826, n_5827, n_5828, n_5829;
  wire n_5830, n_5831, n_5832, n_5833, n_5834, n_5835, n_5836, n_5837;
  wire n_5838, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845;
  wire n_5846, n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853;
  wire n_5854, n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861;
  wire n_5862, n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869;
  wire n_5870, n_5871, n_5872, n_5873, n_5874, n_5875, n_5876, n_5877;
  wire n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885;
  wire n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893;
  wire n_5894, n_5895, n_5897, n_5898, n_5899, n_5900, n_5901, n_5902;
  wire n_5903, n_5904, n_5905, n_5910, n_5911, n_5912, n_5913, n_5914;
  wire n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922;
  wire n_5923, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930;
  wire n_5931, n_5932, n_5933, n_5934, n_5935, n_5936, n_5937, n_5938;
  wire n_5939, n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946;
  wire n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954;
  wire n_5955, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962;
  wire n_5963, n_5964, n_5965, n_5966, n_5967, n_5968, n_5969, n_5970;
  wire n_5971, n_5972, n_5973, n_5974, n_5975, n_5976, n_5977, n_5978;
  wire n_5979, n_5980, n_5981, n_5982, n_5983, n_5984, n_5985, n_5986;
  wire n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5994;
  wire n_5995, n_5996, n_5997, n_5998, n_5999, n_6000, n_6001, n_6002;
  wire n_6003, n_6004, n_6005, n_6006, n_6007, n_6008, n_6009, n_6010;
  wire n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018;
  wire n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025, n_6026;
  wire n_6027, n_6028, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034;
  wire n_6035, n_6036, n_6037, n_6038, n_6039, n_6040, n_6041, n_6042;
  wire n_6043, n_6044, n_6045, n_6046, n_6047, n_6048, n_6049, n_6050;
  wire n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, n_6057, n_6058;
  wire n_6059, n_6060, n_6061, n_6062, n_6063, n_6064, n_6065, n_6066;
  wire n_6067, n_6068, n_6069, n_6070, n_6071, n_6072, n_6073, n_6074;
  wire n_6075, n_6076, n_6077, n_6078, n_6079, n_6080, n_6081, n_6082;
  wire n_6083, n_6084, n_6085, n_6086, n_6087, n_6088, n_6089, n_6090;
  wire n_6091, n_6092, n_6093, n_6094, n_6095, n_6096, n_6097, n_6098;
  wire n_6099, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105, n_6106;
  wire n_6107, n_6108, n_6109, n_6110, n_6111, n_6112, n_6113, n_6114;
  wire n_6115, n_6116, n_6117, n_6118, n_6119, n_6120, n_6121, n_6122;
  wire n_6123, n_6124, n_6125, n_6126, n_6127, n_6128, n_6129, n_6130;
  wire n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137, n_6138;
  wire n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145, n_6146;
  wire n_6147, n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154;
  wire n_6155, n_6156, n_6157, n_6158, n_6159, n_6160, n_6161, n_6162;
  wire n_6163, n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6170;
  wire n_6171, n_6172, n_6173, n_6174, n_6175, n_6176, n_6177, n_6178;
  wire n_6179, n_6180, n_6181, n_6182, n_6183, n_6184, n_6185, n_6186;
  wire n_6187, n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6194;
  wire n_6195, n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202;
  wire n_6203, n_6204, n_6205, n_6206, n_6207, n_6209, n_6210, n_6211;
  wire n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6222, n_6223;
  wire n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231;
  wire n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239;
  wire n_6240, n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247;
  wire n_6248, n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255;
  wire n_6256, n_6257, n_6258, n_6259, n_6260, n_6261, n_6262, n_6263;
  wire n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270, n_6271;
  wire n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278, n_6279;
  wire n_6280, n_6281, n_6282, n_6283, n_6284, n_6285, n_6286, n_6287;
  wire n_6288, n_6289, n_6290, n_6291, n_6292, n_6293, n_6294, n_6295;
  wire n_6296, n_6297, n_6298, n_6299, n_6300, n_6301, n_6302, n_6303;
  wire n_6304, n_6305, n_6306, n_6307, n_6308, n_6309, n_6310, n_6311;
  wire n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319;
  wire n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327;
  wire n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335;
  wire n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343;
  wire n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351;
  wire n_6352, n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359;
  wire n_6360, n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367;
  wire n_6368, n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375;
  wire n_6376, n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383;
  wire n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391;
  wire n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399;
  wire n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407;
  wire n_6408, n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415;
  wire n_6416, n_6417, n_6418, n_6419, n_6420, n_6421, n_6422, n_6423;
  wire n_6424, n_6425, n_6426, n_6427, n_6428, n_6429, n_6430, n_6431;
  wire n_6432, n_6433, n_6434, n_6435, n_6436, n_6437, n_6438, n_6439;
  wire n_6440, n_6441, n_6442, n_6443, n_6444, n_6445, n_6446, n_6447;
  wire n_6448, n_6449, n_6450, n_6451, n_6452, n_6453, n_6454, n_6455;
  wire n_6456, n_6457, n_6458, n_6459, n_6460, n_6461, n_6462, n_6463;
  wire n_6464, n_6465, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471;
  wire n_6472, n_6473, n_6474, n_6475, n_6476, n_6477, n_6478, n_6479;
  wire n_6480, n_6481, n_6482, n_6483, n_6484, n_6485, n_6486, n_6487;
  wire n_6488, n_6489, n_6490, n_6491, n_6492, n_6493, n_6494, n_6495;
  wire n_6496, n_6497, n_6498, n_6499, n_6500, n_6501, n_6502, n_6503;
  wire n_6504, n_6505, n_6506, n_6507, n_6508, n_6509, n_6510, n_6511;
  wire n_6512, n_6513, n_6514, n_6515, n_6516, n_6517, n_6518, n_6519;
  wire n_6520, n_6521, n_6522, n_6523, n_6524, n_6525, n_6526, n_6527;
  wire n_6529, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6536;
  wire n_6537, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548;
  wire n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556;
  wire n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564;
  wire n_6565, n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572;
  wire n_6573, n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6580;
  wire n_6581, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6588;
  wire n_6589, n_6590, n_6591, n_6592, n_6593, n_6594, n_6595, n_6596;
  wire n_6597, n_6598, n_6599, n_6600, n_6601, n_6602, n_6603, n_6604;
  wire n_6605, n_6606, n_6607, n_6608, n_6609, n_6610, n_6611, n_6612;
  wire n_6613, n_6614, n_6615, n_6616, n_6617, n_6618, n_6619, n_6620;
  wire n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6627, n_6628;
  wire n_6629, n_6630, n_6631, n_6632, n_6633, n_6634, n_6635, n_6636;
  wire n_6637, n_6638, n_6639, n_6640, n_6641, n_6642, n_6643, n_6644;
  wire n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652;
  wire n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660;
  wire n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668;
  wire n_6669, n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676;
  wire n_6677, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684;
  wire n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692;
  wire n_6693, n_6694, n_6695, n_6696, n_6697, n_6698, n_6699, n_6700;
  wire n_6701, n_6702, n_6703, n_6704, n_6705, n_6706, n_6707, n_6708;
  wire n_6709, n_6710, n_6711, n_6712, n_6713, n_6714, n_6715, n_6716;
  wire n_6717, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723, n_6724;
  wire n_6725, n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732;
  wire n_6733, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740;
  wire n_6741, n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748;
  wire n_6749, n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756;
  wire n_6757, n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764;
  wire n_6765, n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772;
  wire n_6773, n_6774, n_6775, n_6776, n_6777, n_6778, n_6779, n_6780;
  wire n_6781, n_6782, n_6783, n_6784, n_6785, n_6786, n_6787, n_6788;
  wire n_6789, n_6790, n_6791, n_6792, n_6793, n_6794, n_6795, n_6796;
  wire n_6797, n_6798, n_6799, n_6800, n_6801, n_6802, n_6803, n_6804;
  wire n_6805, n_6806, n_6807, n_6808, n_6809, n_6810, n_6811, n_6812;
  wire n_6813, n_6814, n_6815, n_6816, n_6817, n_6818, n_6819, n_6820;
  wire n_6821, n_6822, n_6823, n_6824, n_6825, n_6826, n_6827, n_6828;
  wire n_6829, n_6830, n_6831, n_6832, n_6833, n_6834, n_6835, n_6836;
  wire n_6837, n_6838, n_6839, n_6840, n_6841, n_6842, n_6843, n_6844;
  wire n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, n_6851, n_6852;
  wire n_6853, n_6854, n_6855, n_6857, n_6858, n_6859, n_6860, n_6861;
  wire n_6862, n_6863, n_6864, n_6865, n_6870, n_6871, n_6872, n_6873;
  wire n_6874, n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881;
  wire n_6882, n_6883, n_6884, n_6885, n_6886, n_6887, n_6888, n_6889;
  wire n_6890, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897;
  wire n_6898, n_6899, n_6900, n_6901, n_6902, n_6903, n_6904, n_6905;
  wire n_6906, n_6907, n_6908, n_6909, n_6910, n_6911, n_6912, n_6913;
  wire n_6914, n_6915, n_6916, n_6917, n_6918, n_6919, n_6920, n_6921;
  wire n_6922, n_6923, n_6924, n_6925, n_6926, n_6927, n_6928, n_6929;
  wire n_6930, n_6931, n_6932, n_6933, n_6934, n_6935, n_6936, n_6937;
  wire n_6938, n_6939, n_6940, n_6941, n_6942, n_6943, n_6944, n_6945;
  wire n_6946, n_6947, n_6948, n_6949, n_6950, n_6951, n_6952, n_6953;
  wire n_6954, n_6955, n_6956, n_6957, n_6958, n_6959, n_6960, n_6961;
  wire n_6962, n_6963, n_6964, n_6965, n_6966, n_6967, n_6968, n_6969;
  wire n_6970, n_6971, n_6972, n_6973, n_6974, n_6975, n_6976, n_6977;
  wire n_6978, n_6979, n_6980, n_6981, n_6982, n_6983, n_6984, n_6985;
  wire n_6986, n_6987, n_6988, n_6989, n_6990, n_6991, n_6992, n_6993;
  wire n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7000, n_7001;
  wire n_7002, n_7003, n_7004, n_7005, n_7006, n_7007, n_7008, n_7009;
  wire n_7010, n_7011, n_7012, n_7013, n_7014, n_7015, n_7016, n_7017;
  wire n_7018, n_7019, n_7020, n_7021, n_7022, n_7023, n_7024, n_7025;
  wire n_7026, n_7027, n_7028, n_7029, n_7030, n_7031, n_7032, n_7033;
  wire n_7034, n_7035, n_7036, n_7037, n_7038, n_7039, n_7040, n_7041;
  wire n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049;
  wire n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7056, n_7057;
  wire n_7058, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065;
  wire n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073;
  wire n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081;
  wire n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089;
  wire n_7090, n_7091, n_7092, n_7093, n_7094, n_7095, n_7096, n_7097;
  wire n_7098, n_7099, n_7100, n_7101, n_7102, n_7103, n_7104, n_7105;
  wire n_7106, n_7107, n_7108, n_7109, n_7110, n_7111, n_7112, n_7113;
  wire n_7114, n_7115, n_7116, n_7117, n_7118, n_7119, n_7120, n_7121;
  wire n_7122, n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129;
  wire n_7130, n_7131, n_7132, n_7133, n_7134, n_7135, n_7136, n_7137;
  wire n_7138, n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145;
  wire n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153;
  wire n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7160, n_7161;
  wire n_7162, n_7163, n_7164, n_7165, n_7166, n_7167, n_7168, n_7169;
  wire n_7170, n_7171, n_7172, n_7173, n_7174, n_7175, n_7176, n_7177;
  wire n_7178, n_7179, n_7180, n_7181, n_7182, n_7183, n_7184, n_7185;
  wire n_7186, n_7187, n_7188, n_7189, n_7190, n_7191, n_7193, n_7194;
  wire n_7195, n_7196, n_7197, n_7198, n_7199, n_7200, n_7201, n_7206;
  wire n_7207, n_7208, n_7209, n_7210, n_7211, n_7212, n_7213, n_7214;
  wire n_7215, n_7216, n_7217, n_7218, n_7219, n_7220, n_7221, n_7222;
  wire n_7223, n_7224, n_7225, n_7226, n_7227, n_7228, n_7229, n_7230;
  wire n_7231, n_7232, n_7233, n_7234, n_7235, n_7236, n_7237, n_7238;
  wire n_7239, n_7240, n_7241, n_7242, n_7243, n_7244, n_7245, n_7246;
  wire n_7247, n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7254;
  wire n_7255, n_7256, n_7257, n_7258, n_7259, n_7260, n_7261, n_7262;
  wire n_7263, n_7264, n_7265, n_7266, n_7267, n_7268, n_7269, n_7270;
  wire n_7271, n_7272, n_7273, n_7274, n_7275, n_7276, n_7277, n_7278;
  wire n_7279, n_7280, n_7281, n_7282, n_7283, n_7284, n_7285, n_7286;
  wire n_7287, n_7288, n_7289, n_7290, n_7291, n_7292, n_7293, n_7294;
  wire n_7295, n_7296, n_7297, n_7298, n_7299, n_7300, n_7301, n_7302;
  wire n_7303, n_7304, n_7305, n_7306, n_7307, n_7308, n_7309, n_7310;
  wire n_7311, n_7312, n_7313, n_7314, n_7315, n_7316, n_7317, n_7318;
  wire n_7319, n_7320, n_7321, n_7322, n_7323, n_7324, n_7325, n_7326;
  wire n_7327, n_7328, n_7329, n_7330, n_7331, n_7332, n_7333, n_7334;
  wire n_7335, n_7336, n_7337, n_7338, n_7339, n_7340, n_7341, n_7342;
  wire n_7343, n_7344, n_7345, n_7346, n_7347, n_7348, n_7349, n_7350;
  wire n_7351, n_7352, n_7353, n_7354, n_7355, n_7356, n_7357, n_7358;
  wire n_7359, n_7360, n_7361, n_7362, n_7363, n_7364, n_7365, n_7366;
  wire n_7367, n_7368, n_7369, n_7370, n_7371, n_7372, n_7373, n_7374;
  wire n_7375, n_7376, n_7377, n_7378, n_7379, n_7380, n_7381, n_7382;
  wire n_7383, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389, n_7390;
  wire n_7391, n_7392, n_7393, n_7394, n_7395, n_7396, n_7397, n_7398;
  wire n_7399, n_7400, n_7401, n_7402, n_7403, n_7404, n_7405, n_7406;
  wire n_7407, n_7408, n_7409, n_7410, n_7411, n_7412, n_7413, n_7414;
  wire n_7415, n_7416, n_7417, n_7418, n_7419, n_7420, n_7421, n_7422;
  wire n_7423, n_7424, n_7425, n_7426, n_7427, n_7428, n_7429, n_7430;
  wire n_7431, n_7432, n_7433, n_7434, n_7435, n_7436, n_7437, n_7438;
  wire n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7446;
  wire n_7447, n_7448, n_7449, n_7450, n_7451, n_7452, n_7453, n_7454;
  wire n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461, n_7462;
  wire n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469, n_7470;
  wire n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477, n_7478;
  wire n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485, n_7486;
  wire n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494;
  wire n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502;
  wire n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510;
  wire n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518;
  wire n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525, n_7526;
  wire n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533, n_7534;
  wire n_7535, n_7537, n_7538, n_7539, n_7540, n_7541, n_7542, n_7543;
  wire n_7544, n_7545, n_7550, n_7551, n_7552, n_7553, n_7554, n_7555;
  wire n_7556, n_7557, n_7558, n_7559, n_7560, n_7561, n_7562, n_7563;
  wire n_7564, n_7565, n_7566, n_7567, n_7568, n_7569, n_7570, n_7571;
  wire n_7572, n_7573, n_7574, n_7575, n_7576, n_7577, n_7578, n_7579;
  wire n_7580, n_7581, n_7582, n_7583, n_7584, n_7585, n_7586, n_7587;
  wire n_7588, n_7589, n_7590, n_7591, n_7592, n_7593, n_7594, n_7595;
  wire n_7596, n_7597, n_7598, n_7599, n_7600, n_7601, n_7602, n_7603;
  wire n_7604, n_7605, n_7606, n_7607, n_7608, n_7609, n_7610, n_7611;
  wire n_7612, n_7613, n_7614, n_7615, n_7616, n_7617, n_7618, n_7619;
  wire n_7620, n_7621, n_7622, n_7623, n_7624, n_7625, n_7626, n_7627;
  wire n_7628, n_7629, n_7630, n_7631, n_7632, n_7633, n_7634, n_7635;
  wire n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643;
  wire n_7644, n_7645, n_7646, n_7647, n_7648, n_7649, n_7650, n_7651;
  wire n_7652, n_7653, n_7654, n_7655, n_7656, n_7657, n_7658, n_7659;
  wire n_7660, n_7661, n_7662, n_7663, n_7664, n_7665, n_7666, n_7667;
  wire n_7668, n_7669, n_7670, n_7671, n_7672, n_7673, n_7674, n_7675;
  wire n_7676, n_7677, n_7678, n_7679, n_7680, n_7681, n_7682, n_7683;
  wire n_7684, n_7685, n_7686, n_7687, n_7688, n_7689, n_7690, n_7691;
  wire n_7692, n_7693, n_7694, n_7695, n_7696, n_7697, n_7698, n_7699;
  wire n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, n_7706, n_7707;
  wire n_7708, n_7709, n_7710, n_7711, n_7712, n_7713, n_7714, n_7715;
  wire n_7716, n_7717, n_7718, n_7719, n_7720, n_7721, n_7722, n_7723;
  wire n_7724, n_7725, n_7726, n_7727, n_7728, n_7729, n_7730, n_7731;
  wire n_7732, n_7733, n_7734, n_7735, n_7736, n_7737, n_7738, n_7739;
  wire n_7740, n_7741, n_7742, n_7743, n_7744, n_7745, n_7746, n_7747;
  wire n_7748, n_7749, n_7750, n_7751, n_7752, n_7753, n_7754, n_7755;
  wire n_7756, n_7757, n_7758, n_7759, n_7760, n_7761, n_7762, n_7763;
  wire n_7764, n_7765, n_7766, n_7767, n_7768, n_7769, n_7770, n_7771;
  wire n_7772, n_7773, n_7774, n_7775, n_7776, n_7777, n_7778, n_7779;
  wire n_7780, n_7781, n_7782, n_7783, n_7784, n_7785, n_7786, n_7787;
  wire n_7788, n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795;
  wire n_7796, n_7797, n_7798, n_7799, n_7800, n_7801, n_7802, n_7803;
  wire n_7804, n_7805, n_7806, n_7807, n_7808, n_7809, n_7810, n_7811;
  wire n_7812, n_7813, n_7814, n_7815, n_7816, n_7817, n_7818, n_7819;
  wire n_7820, n_7821, n_7822, n_7823, n_7824, n_7825, n_7826, n_7827;
  wire n_7828, n_7829, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835;
  wire n_7836, n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7843;
  wire n_7844, n_7845, n_7846, n_7847, n_7848, n_7849, n_7850, n_7851;
  wire n_7852, n_7853, n_7854, n_7855, n_7856, n_7857, n_7858, n_7859;
  wire n_7860, n_7861, n_7862, n_7863, n_7864, n_7865, n_7866, n_7867;
  wire n_7868, n_7869, n_7870, n_7871, n_7872, n_7873, n_7874, n_7875;
  wire n_7876, n_7877, n_7878, n_7879, n_7880, n_7881, n_7882, n_7883;
  wire n_7884, n_7885, n_7886, n_7887, n_7889, n_7890, n_7891, n_7892;
  wire n_7893, n_7894, n_7895, n_7896, n_7897, n_7902, n_7903, n_7904;
  wire n_7905, n_7906, n_7907, n_7908, n_7909, n_7910, n_7911, n_7912;
  wire n_7913, n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920;
  wire n_7921, n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928;
  wire n_7929, n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936;
  wire n_7937, n_7938, n_7939, n_7940, n_7941, n_7942, n_7943, n_7944;
  wire n_7945, n_7946, n_7947, n_7948, n_7949, n_7950, n_7951, n_7952;
  wire n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960;
  wire n_7961, n_7962, n_7963, n_7964, n_7965, n_7966, n_7967, n_7968;
  wire n_7969, n_7970, n_7971, n_7972, n_7973, n_7974, n_7975, n_7976;
  wire n_7977, n_7978, n_7979, n_7980, n_7981, n_7982, n_7983, n_7984;
  wire n_7985, n_7986, n_7987, n_7988, n_7989, n_7990, n_7991, n_7992;
  wire n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999, n_8000;
  wire n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007, n_8008;
  wire n_8009, n_8010, n_8011, n_8012, n_8013, n_8014, n_8015, n_8016;
  wire n_8017, n_8018, n_8019, n_8020, n_8021, n_8022, n_8023, n_8024;
  wire n_8025, n_8026, n_8027, n_8028, n_8029, n_8030, n_8031, n_8032;
  wire n_8033, n_8034, n_8035, n_8036, n_8037, n_8038, n_8039, n_8040;
  wire n_8041, n_8042, n_8043, n_8044, n_8045, n_8046, n_8047, n_8048;
  wire n_8049, n_8050, n_8051, n_8052, n_8053, n_8054, n_8055, n_8056;
  wire n_8057, n_8058, n_8059, n_8060, n_8061, n_8062, n_8063, n_8064;
  wire n_8065, n_8066, n_8067, n_8068, n_8069, n_8070, n_8071, n_8072;
  wire n_8073, n_8074, n_8075, n_8076, n_8077, n_8078, n_8079, n_8080;
  wire n_8081, n_8082, n_8083, n_8084, n_8085, n_8086, n_8087, n_8088;
  wire n_8089, n_8090, n_8091, n_8092, n_8093, n_8094, n_8095, n_8096;
  wire n_8097, n_8098, n_8099, n_8100, n_8101, n_8102, n_8103, n_8104;
  wire n_8105, n_8106, n_8107, n_8108, n_8109, n_8110, n_8111, n_8112;
  wire n_8113, n_8114, n_8115, n_8116, n_8117, n_8118, n_8119, n_8120;
  wire n_8121, n_8122, n_8123, n_8124, n_8125, n_8126, n_8127, n_8128;
  wire n_8129, n_8130, n_8131, n_8132, n_8133, n_8134, n_8135, n_8136;
  wire n_8137, n_8138, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144;
  wire n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152;
  wire n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160;
  wire n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168;
  wire n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176;
  wire n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184;
  wire n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192;
  wire n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200;
  wire n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208;
  wire n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216;
  wire n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224;
  wire n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232;
  wire n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240;
  wire n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8249;
  wire n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256, n_8257;
  wire n_8262, n_8263, n_8264, n_8265, n_8266, n_8267, n_8268, n_8269;
  wire n_8270, n_8271, n_8272, n_8273, n_8274, n_8275, n_8276, n_8277;
  wire n_8278, n_8279, n_8280, n_8281, n_8282, n_8283, n_8284, n_8285;
  wire n_8286, n_8287, n_8288, n_8289, n_8290, n_8291, n_8292, n_8293;
  wire n_8294, n_8295, n_8296, n_8297, n_8298, n_8299, n_8300, n_8301;
  wire n_8302, n_8303, n_8304, n_8305, n_8306, n_8307, n_8308, n_8309;
  wire n_8310, n_8311, n_8312, n_8313, n_8314, n_8315, n_8316, n_8317;
  wire n_8318, n_8319, n_8320, n_8321, n_8322, n_8323, n_8324, n_8325;
  wire n_8326, n_8327, n_8328, n_8329, n_8330, n_8331, n_8332, n_8333;
  wire n_8334, n_8335, n_8336, n_8337, n_8338, n_8339, n_8340, n_8341;
  wire n_8342, n_8343, n_8344, n_8345, n_8346, n_8347, n_8348, n_8349;
  wire n_8350, n_8351, n_8352, n_8353, n_8354, n_8355, n_8356, n_8357;
  wire n_8358, n_8359, n_8360, n_8361, n_8362, n_8363, n_8364, n_8365;
  wire n_8366, n_8367, n_8368, n_8369, n_8370, n_8371, n_8372, n_8373;
  wire n_8374, n_8375, n_8376, n_8377, n_8378, n_8379, n_8380, n_8381;
  wire n_8382, n_8383, n_8384, n_8385, n_8386, n_8387, n_8388, n_8389;
  wire n_8390, n_8391, n_8392, n_8393, n_8394, n_8395, n_8396, n_8397;
  wire n_8398, n_8399, n_8400, n_8401, n_8402, n_8403, n_8404, n_8405;
  wire n_8406, n_8407, n_8408, n_8409, n_8410, n_8411, n_8412, n_8413;
  wire n_8414, n_8415, n_8416, n_8417, n_8418, n_8419, n_8420, n_8421;
  wire n_8422, n_8423, n_8424, n_8425, n_8426, n_8427, n_8428, n_8429;
  wire n_8430, n_8431, n_8432, n_8433, n_8434, n_8435, n_8436, n_8437;
  wire n_8438, n_8439, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445;
  wire n_8446, n_8447, n_8448, n_8449, n_8450, n_8451, n_8452, n_8453;
  wire n_8454, n_8455, n_8456, n_8457, n_8458, n_8459, n_8460, n_8461;
  wire n_8462, n_8463, n_8464, n_8465, n_8466, n_8467, n_8468, n_8469;
  wire n_8470, n_8471, n_8472, n_8473, n_8474, n_8475, n_8476, n_8477;
  wire n_8478, n_8479, n_8480, n_8481, n_8482, n_8483, n_8484, n_8485;
  wire n_8486, n_8487, n_8488, n_8489, n_8490, n_8491, n_8492, n_8493;
  wire n_8494, n_8495, n_8496, n_8497, n_8498, n_8499, n_8500, n_8501;
  wire n_8502, n_8503, n_8504, n_8505, n_8506, n_8507, n_8508, n_8509;
  wire n_8510, n_8511, n_8512, n_8513, n_8514, n_8515, n_8516, n_8517;
  wire n_8518, n_8519, n_8520, n_8521, n_8522, n_8523, n_8524, n_8525;
  wire n_8526, n_8527, n_8528, n_8529, n_8530, n_8531, n_8532, n_8533;
  wire n_8534, n_8535, n_8536, n_8537, n_8538, n_8539, n_8540, n_8541;
  wire n_8542, n_8543, n_8544, n_8545, n_8546, n_8547, n_8548, n_8549;
  wire n_8550, n_8551, n_8552, n_8553, n_8554, n_8555, n_8556, n_8557;
  wire n_8558, n_8559, n_8560, n_8561, n_8562, n_8563, n_8564, n_8565;
  wire n_8566, n_8567, n_8568, n_8569, n_8570, n_8571, n_8572, n_8573;
  wire n_8574, n_8575, n_8576, n_8577, n_8578, n_8579, n_8580, n_8581;
  wire n_8582, n_8583, n_8584, n_8585, n_8586, n_8587, n_8588, n_8589;
  wire n_8590, n_8591, n_8592, n_8593, n_8594, n_8595, n_8596, n_8597;
  wire n_8598, n_8599, n_8600, n_8601, n_8602, n_8603, n_8604, n_8605;
  wire n_8606, n_8607, n_8608, n_8609, n_8610, n_8611, n_8612, n_8613;
  wire n_8614, n_8615, n_8617, n_8618, n_8619, n_8620, n_8621, n_8622;
  wire n_8623, n_8624, n_8625, n_8630, n_8631, n_8632, n_8633, n_8634;
  wire n_8635, n_8636, n_8637, n_8638, n_8639, n_8640, n_8641, n_8642;
  wire n_8643, n_8644, n_8645, n_8646, n_8647, n_8648, n_8649, n_8650;
  wire n_8651, n_8652, n_8653, n_8654, n_8655, n_8656, n_8657, n_8658;
  wire n_8659, n_8660, n_8661, n_8662, n_8663, n_8664, n_8665, n_8666;
  wire n_8667, n_8668, n_8669, n_8670, n_8671, n_8672, n_8673, n_8674;
  wire n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681, n_8682;
  wire n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689, n_8690;
  wire n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697, n_8698;
  wire n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705, n_8706;
  wire n_8707, n_8708, n_8709, n_8710, n_8711, n_8712, n_8713, n_8714;
  wire n_8715, n_8716, n_8717, n_8718, n_8719, n_8720, n_8721, n_8722;
  wire n_8723, n_8724, n_8725, n_8726, n_8727, n_8728, n_8729, n_8730;
  wire n_8731, n_8732, n_8733, n_8734, n_8735, n_8736, n_8737, n_8738;
  wire n_8739, n_8740, n_8741, n_8742, n_8743, n_8744, n_8745, n_8746;
  wire n_8747, n_8748, n_8749, n_8750, n_8751, n_8752, n_8753, n_8754;
  wire n_8755, n_8756, n_8757, n_8758, n_8759, n_8760, n_8761, n_8762;
  wire n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769, n_8770;
  wire n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777, n_8778;
  wire n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786;
  wire n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793, n_8794;
  wire n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802;
  wire n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8809, n_8810;
  wire n_8811, n_8812, n_8813, n_8814, n_8815, n_8816, n_8817, n_8818;
  wire n_8819, n_8820, n_8821, n_8822, n_8823, n_8824, n_8825, n_8826;
  wire n_8827, n_8828, n_8829, n_8830, n_8831, n_8832, n_8833, n_8834;
  wire n_8835, n_8836, n_8837, n_8838, n_8839, n_8840, n_8841, n_8842;
  wire n_8843, n_8844, n_8845, n_8846, n_8847, n_8848, n_8849, n_8850;
  wire n_8851, n_8852, n_8853, n_8854, n_8855, n_8856, n_8857, n_8858;
  wire n_8859, n_8860, n_8861, n_8862, n_8863, n_8864, n_8865, n_8866;
  wire n_8867, n_8868, n_8869, n_8870, n_8871, n_8872, n_8873, n_8874;
  wire n_8875, n_8876, n_8877, n_8878, n_8879, n_8880, n_8881, n_8882;
  wire n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889, n_8890;
  wire n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897, n_8898;
  wire n_8899, n_8900, n_8901, n_8902, n_8903, n_8904, n_8905, n_8906;
  wire n_8907, n_8908, n_8909, n_8910, n_8911, n_8912, n_8913, n_8914;
  wire n_8915, n_8916, n_8917, n_8918, n_8919, n_8920, n_8921, n_8922;
  wire n_8923, n_8924, n_8925, n_8926, n_8927, n_8928, n_8929, n_8930;
  wire n_8931, n_8932, n_8933, n_8934, n_8935, n_8936, n_8937, n_8938;
  wire n_8939, n_8940, n_8941, n_8942, n_8943, n_8944, n_8945, n_8946;
  wire n_8947, n_8948, n_8949, n_8950, n_8951, n_8952, n_8953, n_8954;
  wire n_8955, n_8956, n_8957, n_8958, n_8959, n_8960, n_8961, n_8962;
  wire n_8963, n_8964, n_8965, n_8966, n_8967, n_8968, n_8969, n_8970;
  wire n_8971, n_8972, n_8973, n_8974, n_8975, n_8976, n_8977, n_8978;
  wire n_8979, n_8980, n_8981, n_8982, n_8983, n_8984, n_8985, n_8986;
  wire n_8987, n_8988, n_8989, n_8990, n_8991, n_8993, n_8994, n_8995;
  wire n_8996, n_8997, n_8998, n_8999, n_9000, n_9001, n_9006, n_9007;
  wire n_9008, n_9009, n_9010, n_9011, n_9012, n_9013, n_9014, n_9015;
  wire n_9016, n_9017, n_9018, n_9019, n_9020, n_9021, n_9022, n_9023;
  wire n_9024, n_9025, n_9026, n_9027, n_9028, n_9029, n_9030, n_9031;
  wire n_9032, n_9033, n_9034, n_9035, n_9036, n_9037, n_9038, n_9039;
  wire n_9040, n_9041, n_9042, n_9043, n_9044, n_9045, n_9046, n_9047;
  wire n_9048, n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055;
  wire n_9056, n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063;
  wire n_9064, n_9065, n_9066, n_9067, n_9068, n_9069, n_9070, n_9071;
  wire n_9072, n_9073, n_9074, n_9075, n_9076, n_9077, n_9078, n_9079;
  wire n_9080, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087;
  wire n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095;
  wire n_9096, n_9097, n_9098, n_9099, n_9100, n_9101, n_9102, n_9103;
  wire n_9104, n_9105, n_9106, n_9107, n_9108, n_9109, n_9110, n_9111;
  wire n_9112, n_9113, n_9114, n_9115, n_9116, n_9117, n_9118, n_9119;
  wire n_9120, n_9121, n_9122, n_9123, n_9124, n_9125, n_9126, n_9127;
  wire n_9128, n_9129, n_9130, n_9131, n_9132, n_9133, n_9134, n_9135;
  wire n_9136, n_9137, n_9138, n_9139, n_9140, n_9141, n_9142, n_9143;
  wire n_9144, n_9145, n_9146, n_9147, n_9148, n_9149, n_9150, n_9151;
  wire n_9152, n_9153, n_9154, n_9155, n_9156, n_9157, n_9158, n_9159;
  wire n_9160, n_9161, n_9162, n_9163, n_9164, n_9165, n_9166, n_9167;
  wire n_9168, n_9169, n_9170, n_9171, n_9172, n_9173, n_9174, n_9175;
  wire n_9176, n_9177, n_9178, n_9179, n_9180, n_9181, n_9182, n_9183;
  wire n_9184, n_9185, n_9186, n_9187, n_9188, n_9189, n_9190, n_9191;
  wire n_9192, n_9193, n_9194, n_9195, n_9196, n_9197, n_9198, n_9199;
  wire n_9200, n_9201, n_9202, n_9203, n_9204, n_9205, n_9206, n_9207;
  wire n_9208, n_9209, n_9210, n_9211, n_9212, n_9213, n_9214, n_9215;
  wire n_9216, n_9217, n_9218, n_9219, n_9220, n_9221, n_9222, n_9223;
  wire n_9224, n_9225, n_9226, n_9227, n_9228, n_9229, n_9230, n_9231;
  wire n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9239;
  wire n_9240, n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9247;
  wire n_9248, n_9249, n_9250, n_9251, n_9252, n_9253, n_9254, n_9255;
  wire n_9256, n_9257, n_9258, n_9259, n_9260, n_9261, n_9262, n_9263;
  wire n_9264, n_9265, n_9266, n_9267, n_9268, n_9269, n_9270, n_9271;
  wire n_9272, n_9273, n_9274, n_9275, n_9276, n_9277, n_9278, n_9279;
  wire n_9280, n_9281, n_9282, n_9283, n_9284, n_9285, n_9286, n_9287;
  wire n_9288, n_9289, n_9290, n_9291, n_9292, n_9293, n_9294, n_9295;
  wire n_9296, n_9297, n_9298, n_9299, n_9300, n_9301, n_9302, n_9303;
  wire n_9304, n_9305, n_9306, n_9307, n_9308, n_9309, n_9310, n_9311;
  wire n_9312, n_9313, n_9314, n_9315, n_9316, n_9317, n_9318, n_9319;
  wire n_9320, n_9321, n_9322, n_9323, n_9324, n_9325, n_9326, n_9327;
  wire n_9328, n_9329, n_9330, n_9331, n_9332, n_9333, n_9334, n_9335;
  wire n_9336, n_9337, n_9338, n_9339, n_9340, n_9341, n_9342, n_9343;
  wire n_9344, n_9345, n_9346, n_9347, n_9348, n_9349, n_9350, n_9351;
  wire n_9352, n_9353, n_9354, n_9355, n_9356, n_9357, n_9358, n_9359;
  wire n_9360, n_9361, n_9362, n_9363, n_9364, n_9365, n_9366, n_9367;
  wire n_9368, n_9369, n_9370, n_9371, n_9372, n_9373, n_9374, n_9375;
  wire n_9377, n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9384;
  wire n_9385, n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396;
  wire n_9397, n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404;
  wire n_9405, n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412;
  wire n_9413, n_9414, n_9415, n_9416, n_9417, n_9418, n_9419, n_9420;
  wire n_9421, n_9422, n_9423, n_9424, n_9425, n_9426, n_9427, n_9428;
  wire n_9429, n_9430, n_9431, n_9432, n_9433, n_9434, n_9435, n_9436;
  wire n_9437, n_9438, n_9439, n_9440, n_9441, n_9442, n_9443, n_9444;
  wire n_9445, n_9446, n_9447, n_9448, n_9449, n_9450, n_9451, n_9452;
  wire n_9453, n_9454, n_9455, n_9456, n_9457, n_9458, n_9459, n_9460;
  wire n_9461, n_9462, n_9463, n_9464, n_9465, n_9466, n_9467, n_9468;
  wire n_9469, n_9470, n_9471, n_9472, n_9473, n_9474, n_9475, n_9476;
  wire n_9477, n_9478, n_9479, n_9480, n_9481, n_9482, n_9483, n_9484;
  wire n_9485, n_9486, n_9487, n_9488, n_9489, n_9490, n_9491, n_9492;
  wire n_9493, n_9494, n_9495, n_9496, n_9497, n_9498, n_9499, n_9500;
  wire n_9501, n_9502, n_9503, n_9504, n_9505, n_9506, n_9507, n_9508;
  wire n_9509, n_9510, n_9511, n_9512, n_9513, n_9514, n_9515, n_9516;
  wire n_9517, n_9518, n_9519, n_9520, n_9521, n_9522, n_9523, n_9524;
  wire n_9525, n_9526, n_9527, n_9528, n_9529, n_9530, n_9531, n_9532;
  wire n_9533, n_9534, n_9535, n_9536, n_9537, n_9538, n_9539, n_9540;
  wire n_9541, n_9542, n_9543, n_9544, n_9545, n_9546, n_9547, n_9548;
  wire n_9549, n_9550, n_9551, n_9552, n_9553, n_9554, n_9555, n_9556;
  wire n_9557, n_9558, n_9559, n_9560, n_9561, n_9562, n_9563, n_9564;
  wire n_9565, n_9566, n_9567, n_9568, n_9569, n_9570, n_9571, n_9572;
  wire n_9573, n_9574, n_9575, n_9576, n_9577, n_9578, n_9579, n_9580;
  wire n_9581, n_9582, n_9583, n_9584, n_9585, n_9586, n_9587, n_9588;
  wire n_9589, n_9590, n_9591, n_9592, n_9593, n_9594, n_9595, n_9596;
  wire n_9597, n_9598, n_9599, n_9600, n_9601, n_9602, n_9603, n_9604;
  wire n_9605, n_9606, n_9607, n_9608, n_9609, n_9610, n_9611, n_9612;
  wire n_9613, n_9614, n_9615, n_9616, n_9617, n_9618, n_9619, n_9620;
  wire n_9621, n_9622, n_9623, n_9624, n_9625, n_9626, n_9627, n_9628;
  wire n_9629, n_9630, n_9631, n_9632, n_9633, n_9634, n_9635, n_9636;
  wire n_9637, n_9638, n_9639, n_9640, n_9641, n_9642, n_9643, n_9644;
  wire n_9645, n_9646, n_9647, n_9648, n_9649, n_9650, n_9651, n_9652;
  wire n_9653, n_9654, n_9655, n_9656, n_9657, n_9658, n_9659, n_9660;
  wire n_9661, n_9662, n_9663, n_9664, n_9665, n_9666, n_9667, n_9668;
  wire n_9669, n_9670, n_9671, n_9672, n_9673, n_9674, n_9675, n_9676;
  wire n_9677, n_9678, n_9679, n_9680, n_9681, n_9682, n_9683, n_9684;
  wire n_9685, n_9686, n_9687, n_9688, n_9689, n_9690, n_9691, n_9692;
  wire n_9693, n_9694, n_9695, n_9696, n_9697, n_9698, n_9699, n_9700;
  wire n_9701, n_9702, n_9703, n_9704, n_9705, n_9706, n_9707, n_9708;
  wire n_9709, n_9710, n_9711, n_9712, n_9713, n_9714, n_9715, n_9716;
  wire n_9717, n_9718, n_9719, n_9720, n_9721, n_9722, n_9723, n_9724;
  wire n_9725, n_9726, n_9727, n_9728, n_9729, n_9730, n_9731, n_9732;
  wire n_9733, n_9734, n_9735, n_9736, n_9737, n_9738, n_9739, n_9740;
  wire n_9741, n_9742, n_9743, n_9744, n_9745, n_9746, n_9747, n_9748;
  wire n_9749, n_9750, n_9751, n_9752, n_9753, n_9754, n_9755, n_9756;
  wire n_9757, n_9758, n_9759, n_9760, n_9761, n_9762, n_9763, n_9764;
  wire n_9765, n_9766, n_9767, n_9769, n_9770, n_9771, n_9772, n_9773;
  wire n_9774, n_9775, n_9776, n_9777, n_9782, n_9783, n_9784, n_9785;
  wire n_9786, n_9787, n_9788, n_9789, n_9790, n_9791, n_9792, n_9793;
  wire n_9794, n_9795, n_9796, n_9797, n_9798, n_9799, n_9800, n_9801;
  wire n_9802, n_9803, n_9804, n_9805, n_9806, n_9807, n_9808, n_9809;
  wire n_9810, n_9811, n_9812, n_9813, n_9814, n_9815, n_9816, n_9817;
  wire n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_9825;
  wire n_9826, n_9827, n_9828, n_9829, n_9830, n_9831, n_9832, n_9833;
  wire n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841;
  wire n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848, n_9849;
  wire n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856, n_9857;
  wire n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864, n_9865;
  wire n_9866, n_9867, n_9868, n_9869, n_9870, n_9871, n_9872, n_9873;
  wire n_9874, n_9875, n_9876, n_9877, n_9878, n_9879, n_9880, n_9881;
  wire n_9882, n_9883, n_9884, n_9885, n_9886, n_9887, n_9888, n_9889;
  wire n_9890, n_9891, n_9892, n_9893, n_9894, n_9895, n_9896, n_9897;
  wire n_9898, n_9899, n_9900, n_9901, n_9902, n_9903, n_9904, n_9905;
  wire n_9906, n_9907, n_9908, n_9909, n_9910, n_9911, n_9912, n_9913;
  wire n_9914, n_9915, n_9916, n_9917, n_9918, n_9919, n_9920, n_9921;
  wire n_9922, n_9923, n_9924, n_9925, n_9926, n_9927, n_9928, n_9929;
  wire n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937;
  wire n_9938, n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945;
  wire n_9946, n_9947, n_9948, n_9949, n_9950, n_9951, n_9952, n_9953;
  wire n_9954, n_9955, n_9956, n_9957, n_9958, n_9959, n_9960, n_9961;
  wire n_9962, n_9963, n_9964, n_9965, n_9966, n_9967, n_9968, n_9969;
  wire n_9970, n_9971, n_9972, n_9973, n_9974, n_9975, n_9976, n_9977;
  wire n_9978, n_9979, n_9980, n_9981, n_9982, n_9983, n_9984, n_9985;
  wire n_9986, n_9987, n_9988, n_9989, n_9990, n_9991, n_9992, n_9993;
  wire n_9994, n_9995, n_9996, n_9997, n_9998, n_9999, n_10000, n_10001;
  wire n_10002, n_10003, n_10004, n_10005, n_10006, n_10007, n_10008,
       n_10009;
  wire n_10010, n_10011, n_10012, n_10013, n_10014, n_10015, n_10016,
       n_10017;
  wire n_10018, n_10019, n_10020, n_10021, n_10022, n_10023, n_10024,
       n_10025;
  wire n_10026, n_10027, n_10028, n_10029, n_10030, n_10031, n_10032,
       n_10033;
  wire n_10034, n_10035, n_10036, n_10037, n_10038, n_10039, n_10040,
       n_10041;
  wire n_10042, n_10043, n_10044, n_10045, n_10046, n_10047, n_10048,
       n_10049;
  wire n_10050, n_10051, n_10052, n_10053, n_10054, n_10055, n_10056,
       n_10057;
  wire n_10058, n_10059, n_10060, n_10061, n_10062, n_10063, n_10064,
       n_10065;
  wire n_10066, n_10067, n_10068, n_10069, n_10070, n_10071, n_10072,
       n_10073;
  wire n_10074, n_10075, n_10076, n_10077, n_10078, n_10079, n_10080,
       n_10081;
  wire n_10082, n_10083, n_10084, n_10085, n_10086, n_10087, n_10088,
       n_10089;
  wire n_10090, n_10091, n_10092, n_10093, n_10094, n_10095, n_10096,
       n_10097;
  wire n_10098, n_10099, n_10100, n_10101, n_10102, n_10103, n_10104,
       n_10105;
  wire n_10106, n_10107, n_10108, n_10109, n_10110, n_10111, n_10112,
       n_10113;
  wire n_10114, n_10115, n_10116, n_10117, n_10118, n_10119, n_10120,
       n_10121;
  wire n_10122, n_10123, n_10124, n_10125, n_10126, n_10127, n_10128,
       n_10129;
  wire n_10130, n_10131, n_10132, n_10133, n_10134, n_10135, n_10136,
       n_10137;
  wire n_10138, n_10139, n_10140, n_10141, n_10142, n_10143, n_10144,
       n_10145;
  wire n_10146, n_10147, n_10148, n_10149, n_10150, n_10151, n_10152,
       n_10153;
  wire n_10154, n_10155, n_10156, n_10157, n_10158, n_10159, n_10160,
       n_10161;
  wire n_10162, n_10163, n_10164, n_10165, n_10166, n_10167, n_10169,
       n_10170;
  wire n_10171, n_10172, n_10173, n_10174, n_10175, n_10176, n_10177,
       n_10182;
  wire n_10183, n_10184, n_10185, n_10186, n_10187, n_10188, n_10189,
       n_10190;
  wire n_10191, n_10192, n_10193, n_10194, n_10195, n_10196, n_10197,
       n_10198;
  wire n_10199, n_10200, n_10201, n_10202, n_10203, n_10204, n_10205,
       n_10206;
  wire n_10207, n_10208, n_10209, n_10210, n_10211, n_10212, n_10213,
       n_10214;
  wire n_10215, n_10216, n_10217, n_10218, n_10219, n_10220, n_10221,
       n_10222;
  wire n_10223, n_10224, n_10225, n_10226, n_10227, n_10228, n_10229,
       n_10230;
  wire n_10231, n_10232, n_10233, n_10234, n_10235, n_10236, n_10237,
       n_10238;
  wire n_10239, n_10240, n_10241, n_10242, n_10243, n_10244, n_10245,
       n_10246;
  wire n_10247, n_10248, n_10249, n_10250, n_10251, n_10252, n_10253,
       n_10254;
  wire n_10255, n_10256, n_10257, n_10258, n_10259, n_10260, n_10261,
       n_10262;
  wire n_10263, n_10264, n_10265, n_10266, n_10267, n_10268, n_10269,
       n_10270;
  wire n_10271, n_10272, n_10273, n_10274, n_10275, n_10276, n_10277,
       n_10278;
  wire n_10279, n_10280, n_10281, n_10282, n_10283, n_10284, n_10285,
       n_10286;
  wire n_10287, n_10288, n_10289, n_10290, n_10291, n_10292, n_10293,
       n_10294;
  wire n_10295, n_10296, n_10297, n_10298, n_10299, n_10300, n_10301,
       n_10302;
  wire n_10303, n_10304, n_10305, n_10306, n_10307, n_10308, n_10309,
       n_10310;
  wire n_10311, n_10312, n_10313, n_10314, n_10315, n_10316, n_10317,
       n_10318;
  wire n_10319, n_10320, n_10321, n_10322, n_10323, n_10324, n_10325,
       n_10326;
  wire n_10327, n_10328, n_10329, n_10330, n_10331, n_10332, n_10333,
       n_10334;
  wire n_10335, n_10336, n_10337, n_10338, n_10339, n_10340, n_10341,
       n_10342;
  wire n_10343, n_10344, n_10345, n_10346, n_10347, n_10348, n_10349,
       n_10350;
  wire n_10351, n_10352, n_10353, n_10354, n_10355, n_10356, n_10357,
       n_10358;
  wire n_10359, n_10360, n_10361, n_10362, n_10363, n_10364, n_10365,
       n_10366;
  wire n_10367, n_10368, n_10369, n_10370, n_10371, n_10372, n_10373,
       n_10374;
  wire n_10375, n_10376, n_10377, n_10378, n_10379, n_10380, n_10381,
       n_10382;
  wire n_10383, n_10384, n_10385, n_10386, n_10387, n_10388, n_10389,
       n_10390;
  wire n_10391, n_10392, n_10393, n_10394, n_10395, n_10396, n_10397,
       n_10398;
  wire n_10399, n_10400, n_10401, n_10402, n_10403, n_10404, n_10405,
       n_10406;
  wire n_10407, n_10408, n_10409, n_10410, n_10411, n_10412, n_10413,
       n_10414;
  wire n_10415, n_10416, n_10417, n_10418, n_10419, n_10420, n_10421,
       n_10422;
  wire n_10423, n_10424, n_10425, n_10426, n_10427, n_10428, n_10429,
       n_10430;
  wire n_10431, n_10432, n_10433, n_10434, n_10435, n_10436, n_10437,
       n_10438;
  wire n_10439, n_10440, n_10441, n_10442, n_10443, n_10444, n_10445,
       n_10446;
  wire n_10447, n_10448, n_10449, n_10450, n_10451, n_10452, n_10453,
       n_10454;
  wire n_10455, n_10456, n_10457, n_10458, n_10459, n_10460, n_10461,
       n_10462;
  wire n_10463, n_10464, n_10465, n_10466, n_10467, n_10468, n_10469,
       n_10470;
  wire n_10471, n_10472, n_10473, n_10474, n_10475, n_10476, n_10477,
       n_10478;
  wire n_10479, n_10480, n_10481, n_10482, n_10483, n_10484, n_10485,
       n_10486;
  wire n_10487, n_10488, n_10489, n_10490, n_10491, n_10492, n_10493,
       n_10494;
  wire n_10495, n_10496, n_10497, n_10498, n_10499, n_10500, n_10501,
       n_10502;
  wire n_10503, n_10504, n_10505, n_10506, n_10507, n_10508, n_10509,
       n_10510;
  wire n_10511, n_10512, n_10513, n_10514, n_10515, n_10516, n_10517,
       n_10518;
  wire n_10519, n_10520, n_10521, n_10522, n_10523, n_10524, n_10525,
       n_10526;
  wire n_10527, n_10528, n_10529, n_10530, n_10531, n_10532, n_10533,
       n_10534;
  wire n_10535, n_10536, n_10537, n_10538, n_10539, n_10540, n_10541,
       n_10542;
  wire n_10543, n_10544, n_10545, n_10546, n_10547, n_10548, n_10549,
       n_10550;
  wire n_10551, n_10552, n_10553, n_10554, n_10555, n_10556, n_10557,
       n_10558;
  wire n_10559, n_10560, n_10561, n_10562, n_10563, n_10564, n_10565,
       n_10566;
  wire n_10567, n_10568, n_10569, n_10570, n_10571, n_10572, n_10573,
       n_10574;
  wire n_10575, n_10577, n_10578, n_10579, n_10580, n_10581, n_10582,
       n_10583;
  wire n_10584, n_10585, n_10590, n_10591, n_10592, n_10593, n_10594,
       n_10595;
  wire n_10596, n_10597, n_10598, n_10599, n_10600, n_10601, n_10602,
       n_10603;
  wire n_10604, n_10605, n_10606, n_10607, n_10608, n_10609, n_10610,
       n_10611;
  wire n_10612, n_10613, n_10614, n_10615, n_10616, n_10617, n_10618,
       n_10619;
  wire n_10620, n_10621, n_10622, n_10623, n_10624, n_10625, n_10626,
       n_10627;
  wire n_10628, n_10629, n_10630, n_10631, n_10632, n_10633, n_10634,
       n_10635;
  wire n_10636, n_10637, n_10638, n_10639, n_10640, n_10641, n_10642,
       n_10643;
  wire n_10644, n_10645, n_10646, n_10647, n_10648, n_10649, n_10650,
       n_10651;
  wire n_10652, n_10653, n_10654, n_10655, n_10656, n_10657, n_10658,
       n_10659;
  wire n_10660, n_10661, n_10662, n_10663, n_10664, n_10665, n_10666,
       n_10667;
  wire n_10668, n_10669, n_10670, n_10671, n_10672, n_10673, n_10674,
       n_10675;
  wire n_10676, n_10677, n_10678, n_10679, n_10680, n_10681, n_10682,
       n_10683;
  wire n_10684, n_10685, n_10686, n_10687, n_10688, n_10689, n_10690,
       n_10691;
  wire n_10692, n_10693, n_10694, n_10695, n_10696, n_10697, n_10698,
       n_10699;
  wire n_10700, n_10701, n_10702, n_10703, n_10704, n_10705, n_10706,
       n_10707;
  wire n_10708, n_10709, n_10710, n_10711, n_10712, n_10713, n_10714,
       n_10715;
  wire n_10716, n_10717, n_10718, n_10719, n_10720, n_10721, n_10722,
       n_10723;
  wire n_10724, n_10725, n_10726, n_10727, n_10728, n_10729, n_10730,
       n_10731;
  wire n_10732, n_10733, n_10734, n_10735, n_10736, n_10737, n_10738,
       n_10739;
  wire n_10740, n_10741, n_10742, n_10743, n_10744, n_10745, n_10746,
       n_10747;
  wire n_10748, n_10749, n_10750, n_10751, n_10752, n_10753, n_10754,
       n_10755;
  wire n_10756, n_10757, n_10758, n_10759, n_10760, n_10761, n_10762,
       n_10763;
  wire n_10764, n_10765, n_10766, n_10767, n_10768, n_10769, n_10770,
       n_10771;
  wire n_10772, n_10773, n_10774, n_10775, n_10776, n_10777, n_10778,
       n_10779;
  wire n_10780, n_10781, n_10782, n_10783, n_10784, n_10785, n_10786,
       n_10787;
  wire n_10788, n_10789, n_10790, n_10791, n_10792, n_10793, n_10794,
       n_10795;
  wire n_10796, n_10797, n_10798, n_10799, n_10800, n_10801, n_10802,
       n_10803;
  wire n_10804, n_10805, n_10806, n_10807, n_10808, n_10809, n_10810,
       n_10811;
  wire n_10812, n_10813, n_10814, n_10815, n_10816, n_10817, n_10818,
       n_10819;
  wire n_10820, n_10821, n_10822, n_10823, n_10824, n_10825, n_10826,
       n_10827;
  wire n_10828, n_10829, n_10830, n_10831, n_10832, n_10833, n_10834,
       n_10835;
  wire n_10836, n_10837, n_10838, n_10839, n_10840, n_10841, n_10842,
       n_10843;
  wire n_10844, n_10845, n_10846, n_10847, n_10848, n_10849, n_10850,
       n_10851;
  wire n_10852, n_10853, n_10854, n_10855, n_10856, n_10857, n_10858,
       n_10859;
  wire n_10860, n_10861, n_10862, n_10863, n_10864, n_10865, n_10866,
       n_10867;
  wire n_10868, n_10869, n_10870, n_10871, n_10872, n_10873, n_10874,
       n_10875;
  wire n_10876, n_10877, n_10878, n_10879, n_10880, n_10881, n_10882,
       n_10883;
  wire n_10884, n_10885, n_10886, n_10887, n_10888, n_10889, n_10890,
       n_10891;
  wire n_10892, n_10893, n_10894, n_10895, n_10896, n_10897, n_10898,
       n_10899;
  wire n_10900, n_10901, n_10902, n_10903, n_10904, n_10905, n_10906,
       n_10907;
  wire n_10908, n_10909, n_10910, n_10911, n_10912, n_10913, n_10914,
       n_10915;
  wire n_10916, n_10917, n_10918, n_10919, n_10920, n_10921, n_10922,
       n_10923;
  wire n_10924, n_10925, n_10926, n_10927, n_10928, n_10929, n_10930,
       n_10931;
  wire n_10932, n_10933, n_10934, n_10935, n_10936, n_10937, n_10938,
       n_10939;
  wire n_10940, n_10941, n_10942, n_10943, n_10944, n_10945, n_10946,
       n_10947;
  wire n_10948, n_10949, n_10950, n_10951, n_10952, n_10953, n_10954,
       n_10955;
  wire n_10956, n_10957, n_10958, n_10959, n_10960, n_10961, n_10962,
       n_10963;
  wire n_10964, n_10965, n_10966, n_10967, n_10968, n_10969, n_10970,
       n_10971;
  wire n_10972, n_10973, n_10974, n_10975, n_10976, n_10977, n_10978,
       n_10979;
  wire n_10980, n_10981, n_10982, n_10983, n_10984, n_10985, n_10986,
       n_10987;
  wire n_10988, n_10989, n_10990, n_10991, n_10993, n_10994, n_10995,
       n_10996;
  wire n_10997, n_10998, n_10999, n_11000, n_11001, n_11006, n_11007,
       n_11008;
  wire n_11009, n_11010, n_11011, n_11012, n_11013, n_11014, n_11015,
       n_11016;
  wire n_11017, n_11018, n_11019, n_11020, n_11021, n_11022, n_11023,
       n_11024;
  wire n_11025, n_11026, n_11027, n_11028, n_11029, n_11030, n_11031,
       n_11032;
  wire n_11033, n_11034, n_11035, n_11036, n_11037, n_11038, n_11039,
       n_11040;
  wire n_11041, n_11042, n_11043, n_11044, n_11045, n_11046, n_11047,
       n_11048;
  wire n_11049, n_11050, n_11051, n_11052, n_11053, n_11054, n_11055,
       n_11056;
  wire n_11057, n_11058, n_11059, n_11060, n_11061, n_11062, n_11063,
       n_11064;
  wire n_11065, n_11066, n_11067, n_11068, n_11069, n_11070, n_11071,
       n_11072;
  wire n_11073, n_11074, n_11075, n_11076, n_11077, n_11078, n_11079,
       n_11080;
  wire n_11081, n_11082, n_11083, n_11084, n_11085, n_11086, n_11087,
       n_11088;
  wire n_11089, n_11090, n_11091, n_11092, n_11093, n_11094, n_11095,
       n_11096;
  wire n_11097, n_11098, n_11099, n_11100, n_11101, n_11102, n_11103,
       n_11104;
  wire n_11105, n_11106, n_11107, n_11108, n_11109, n_11110, n_11111,
       n_11112;
  wire n_11113, n_11114, n_11115, n_11116, n_11117, n_11118, n_11119,
       n_11120;
  wire n_11121, n_11122, n_11123, n_11124, n_11125, n_11126, n_11127,
       n_11128;
  wire n_11129, n_11130, n_11131, n_11132, n_11133, n_11134, n_11135,
       n_11136;
  wire n_11137, n_11138, n_11139, n_11140, n_11141, n_11142, n_11143,
       n_11144;
  wire n_11145, n_11146, n_11147, n_11148, n_11149, n_11150, n_11151,
       n_11152;
  wire n_11153, n_11154, n_11155, n_11156, n_11157, n_11158, n_11159,
       n_11160;
  wire n_11161, n_11162, n_11163, n_11164, n_11165, n_11166, n_11167,
       n_11168;
  wire n_11169, n_11170, n_11171, n_11172, n_11173, n_11174, n_11175,
       n_11176;
  wire n_11177, n_11178, n_11179, n_11180, n_11181, n_11182, n_11183,
       n_11184;
  wire n_11185, n_11186, n_11187, n_11188, n_11189, n_11190, n_11191,
       n_11192;
  wire n_11193, n_11194, n_11195, n_11196, n_11197, n_11198, n_11199,
       n_11200;
  wire n_11201, n_11202, n_11203, n_11204, n_11205, n_11206, n_11207,
       n_11208;
  wire n_11209, n_11210, n_11211, n_11212, n_11213, n_11214, n_11215,
       n_11216;
  wire n_11217, n_11218, n_11219, n_11220, n_11221, n_11222, n_11223,
       n_11224;
  wire n_11225, n_11226, n_11227, n_11228, n_11229, n_11230, n_11231,
       n_11232;
  wire n_11233, n_11234, n_11235, n_11236, n_11237, n_11238, n_11239,
       n_11240;
  wire n_11241, n_11242, n_11243, n_11244, n_11245, n_11246, n_11247,
       n_11248;
  wire n_11249, n_11250, n_11251, n_11252, n_11253, n_11254, n_11255,
       n_11256;
  wire n_11257, n_11258, n_11259, n_11260, n_11261, n_11262, n_11263,
       n_11264;
  wire n_11265, n_11266, n_11267, n_11268, n_11269, n_11270, n_11271,
       n_11272;
  wire n_11273, n_11274, n_11275, n_11276, n_11277, n_11278, n_11279,
       n_11280;
  wire n_11281, n_11282, n_11283, n_11284, n_11285, n_11286, n_11287,
       n_11288;
  wire n_11289, n_11290, n_11291, n_11292, n_11293, n_11294, n_11295,
       n_11296;
  wire n_11297, n_11298, n_11299, n_11300, n_11301, n_11302, n_11303,
       n_11304;
  wire n_11305, n_11306, n_11307, n_11308, n_11309, n_11310, n_11311,
       n_11312;
  wire n_11313, n_11314, n_11315, n_11316, n_11317, n_11318, n_11319,
       n_11320;
  wire n_11321, n_11322, n_11323, n_11324, n_11325, n_11326, n_11327,
       n_11328;
  wire n_11329, n_11330, n_11331, n_11332, n_11333, n_11334, n_11335,
       n_11336;
  wire n_11337, n_11338, n_11339, n_11340, n_11341, n_11342, n_11343,
       n_11344;
  wire n_11345, n_11346, n_11347, n_11348, n_11349, n_11350, n_11351,
       n_11352;
  wire n_11353, n_11354, n_11355, n_11356, n_11357, n_11358, n_11359,
       n_11360;
  wire n_11361, n_11362, n_11363, n_11364, n_11365, n_11366, n_11367,
       n_11368;
  wire n_11369, n_11370, n_11371, n_11372, n_11373, n_11374, n_11375,
       n_11376;
  wire n_11377, n_11378, n_11379, n_11380, n_11381, n_11382, n_11383,
       n_11384;
  wire n_11385, n_11386, n_11387, n_11388, n_11389, n_11390, n_11391,
       n_11392;
  wire n_11393, n_11394, n_11395, n_11396, n_11397, n_11398, n_11399,
       n_11400;
  wire n_11401, n_11402, n_11403, n_11404, n_11405, n_11406, n_11407,
       n_11408;
  wire n_11409, n_11410, n_11411, n_11412, n_11413, n_11414, n_11415,
       n_11417;
  wire n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424,
       n_11425;
  wire n_11430, n_11431, n_11432, n_11433, n_11434, n_11435, n_11436,
       n_11437;
  wire n_11438, n_11439, n_11440, n_11441, n_11442, n_11443, n_11444,
       n_11445;
  wire n_11446, n_11447, n_11448, n_11449, n_11450, n_11451, n_11452,
       n_11453;
  wire n_11454, n_11455, n_11456, n_11457, n_11458, n_11459, n_11460,
       n_11461;
  wire n_11462, n_11463, n_11464, n_11465, n_11466, n_11467, n_11468,
       n_11469;
  wire n_11470, n_11471, n_11472, n_11473, n_11474, n_11475, n_11476,
       n_11477;
  wire n_11478, n_11479, n_11480, n_11481, n_11482, n_11483, n_11484,
       n_11485;
  wire n_11486, n_11487, n_11488, n_11489, n_11490, n_11491, n_11492,
       n_11493;
  wire n_11494, n_11495, n_11496, n_11497, n_11498, n_11499, n_11500,
       n_11501;
  wire n_11502, n_11503, n_11504, n_11505, n_11506, n_11507, n_11508,
       n_11509;
  wire n_11510, n_11511, n_11512, n_11513, n_11514, n_11515, n_11516,
       n_11517;
  wire n_11518, n_11519, n_11520, n_11521, n_11522, n_11523, n_11524,
       n_11525;
  wire n_11526, n_11527, n_11528, n_11529, n_11530, n_11531, n_11532,
       n_11533;
  wire n_11534, n_11535, n_11536, n_11537, n_11538, n_11539, n_11540,
       n_11541;
  wire n_11542, n_11543, n_11544, n_11545, n_11546, n_11547, n_11548,
       n_11549;
  wire n_11550, n_11551, n_11552, n_11553, n_11554, n_11555, n_11556,
       n_11557;
  wire n_11558, n_11559, n_11560, n_11561, n_11562, n_11563, n_11564,
       n_11565;
  wire n_11566, n_11567, n_11568, n_11569, n_11570, n_11571, n_11572,
       n_11573;
  wire n_11574, n_11575, n_11576, n_11577, n_11578, n_11579, n_11580,
       n_11581;
  wire n_11582, n_11583, n_11584, n_11585, n_11586, n_11587, n_11588,
       n_11589;
  wire n_11590, n_11591, n_11592, n_11593, n_11594, n_11595, n_11596,
       n_11597;
  wire n_11598, n_11599, n_11600, n_11601, n_11602, n_11603, n_11604,
       n_11605;
  wire n_11606, n_11607, n_11608, n_11609, n_11610, n_11611, n_11612,
       n_11613;
  wire n_11614, n_11615, n_11616, n_11617, n_11618, n_11619, n_11620,
       n_11621;
  wire n_11622, n_11623, n_11624, n_11625, n_11626, n_11627, n_11628,
       n_11629;
  wire n_11630, n_11631, n_11632, n_11633, n_11634, n_11635, n_11636,
       n_11637;
  wire n_11638, n_11639, n_11640, n_11641, n_11642, n_11643, n_11644,
       n_11645;
  wire n_11646, n_11647, n_11648, n_11649, n_11650, n_11651, n_11652,
       n_11653;
  wire n_11654, n_11655, n_11656, n_11657, n_11658, n_11659, n_11660,
       n_11661;
  wire n_11662, n_11663, n_11664, n_11665, n_11666, n_11667, n_11668,
       n_11669;
  wire n_11670, n_11671, n_11672, n_11673, n_11674, n_11675, n_11676,
       n_11677;
  wire n_11678, n_11679, n_11680, n_11681, n_11682, n_11683, n_11684,
       n_11685;
  wire n_11686, n_11687, n_11688, n_11689, n_11690, n_11691, n_11692,
       n_11693;
  wire n_11694, n_11695, n_11696, n_11697, n_11698, n_11699, n_11700,
       n_11701;
  wire n_11702, n_11703, n_11704, n_11705, n_11706, n_11707, n_11708,
       n_11709;
  wire n_11710, n_11711, n_11712, n_11713, n_11714, n_11715, n_11716,
       n_11717;
  wire n_11718, n_11719, n_11720, n_11721, n_11722, n_11723, n_11724,
       n_11725;
  wire n_11726, n_11727, n_11728, n_11729, n_11730, n_11731, n_11732,
       n_11733;
  wire n_11734, n_11735, n_11736, n_11737, n_11738, n_11739, n_11740,
       n_11741;
  wire n_11742, n_11743, n_11744, n_11745, n_11746, n_11747, n_11748,
       n_11749;
  wire n_11750, n_11751, n_11752, n_11753, n_11754, n_11755, n_11756,
       n_11757;
  wire n_11758, n_11759, n_11760, n_11761, n_11762, n_11763, n_11764,
       n_11765;
  wire n_11766, n_11767, n_11768, n_11769, n_11770, n_11771, n_11772,
       n_11773;
  wire n_11774, n_11775, n_11776, n_11777, n_11778, n_11779, n_11780,
       n_11781;
  wire n_11782, n_11783, n_11784, n_11785, n_11786, n_11787, n_11788,
       n_11789;
  wire n_11790, n_11791, n_11792, n_11793, n_11794, n_11795, n_11796,
       n_11797;
  wire n_11798, n_11799, n_11800, n_11801, n_11802, n_11803, n_11804,
       n_11805;
  wire n_11806, n_11807, n_11808, n_11809, n_11810, n_11811, n_11812,
       n_11813;
  wire n_11814, n_11815, n_11816, n_11817, n_11818, n_11819, n_11820,
       n_11821;
  wire n_11822, n_11823, n_11824, n_11825, n_11826, n_11827, n_11828,
       n_11829;
  wire n_11830, n_11831, n_11832, n_11833, n_11834, n_11835, n_11836,
       n_11837;
  wire n_11838, n_11839, n_11840, n_11841, n_11842, n_11843, n_11844,
       n_11845;
  wire n_11846, n_11847, n_11849, n_11850, n_11851, n_11852, n_11853,
       n_11854;
  wire n_11855, n_11856, n_11857, n_11862, n_11863, n_11864, n_11865,
       n_11866;
  wire n_11867, n_11868, n_11869, n_11870, n_11871, n_11872, n_11873,
       n_11874;
  wire n_11875, n_11876, n_11877, n_11878, n_11879, n_11880, n_11881,
       n_11882;
  wire n_11883, n_11884, n_11885, n_11886, n_11887, n_11888, n_11889,
       n_11890;
  wire n_11891, n_11892, n_11893, n_11894, n_11895, n_11896, n_11897,
       n_11898;
  wire n_11899, n_11900, n_11901, n_11902, n_11903, n_11904, n_11905,
       n_11906;
  wire n_11907, n_11908, n_11909, n_11910, n_11911, n_11912, n_11913,
       n_11914;
  wire n_11915, n_11916, n_11917, n_11918, n_11919, n_11920, n_11921,
       n_11922;
  wire n_11923, n_11924, n_11925, n_11926, n_11927, n_11928, n_11929,
       n_11930;
  wire n_11931, n_11932, n_11933, n_11934, n_11935, n_11936, n_11937,
       n_11938;
  wire n_11939, n_11940, n_11941, n_11942, n_11943, n_11944, n_11945,
       n_11946;
  wire n_11947, n_11948, n_11949, n_11950, n_11951, n_11952, n_11953,
       n_11954;
  wire n_11955, n_11956, n_11957, n_11958, n_11959, n_11960, n_11961,
       n_11962;
  wire n_11963, n_11964, n_11965, n_11966, n_11967, n_11968, n_11969,
       n_11970;
  wire n_11971, n_11972, n_11973, n_11974, n_11975, n_11976, n_11977,
       n_11978;
  wire n_11979, n_11980, n_11981, n_11982, n_11983, n_11984, n_11985,
       n_11986;
  wire n_11987, n_11988, n_11989, n_11990, n_11991, n_11992, n_11993,
       n_11994;
  wire n_11995, n_11996, n_11997, n_11998, n_11999, n_12000, n_12001,
       n_12002;
  wire n_12003, n_12004, n_12005, n_12006, n_12007, n_12008, n_12009,
       n_12010;
  wire n_12011, n_12012, n_12013, n_12014, n_12015, n_12016, n_12017,
       n_12018;
  wire n_12019, n_12020, n_12021, n_12022, n_12023, n_12024, n_12025,
       n_12026;
  wire n_12027, n_12028, n_12029, n_12030, n_12031, n_12032, n_12033,
       n_12034;
  wire n_12035, n_12036, n_12037, n_12038, n_12039, n_12040, n_12041,
       n_12042;
  wire n_12043, n_12044, n_12045, n_12046, n_12047, n_12048, n_12049,
       n_12050;
  wire n_12051, n_12052, n_12053, n_12054, n_12055, n_12056, n_12057,
       n_12058;
  wire n_12059, n_12060, n_12061, n_12062, n_12063, n_12064, n_12065,
       n_12066;
  wire n_12067, n_12068, n_12069, n_12070, n_12071, n_12072, n_12073,
       n_12074;
  wire n_12075, n_12076, n_12077, n_12078, n_12079, n_12080, n_12081,
       n_12082;
  wire n_12083, n_12084, n_12085, n_12086, n_12087, n_12088, n_12089,
       n_12090;
  wire n_12091, n_12092, n_12093, n_12094, n_12095, n_12096, n_12097,
       n_12098;
  wire n_12099, n_12100, n_12101, n_12102, n_12103, n_12104, n_12105,
       n_12106;
  wire n_12107, n_12108, n_12109, n_12110, n_12111, n_12112, n_12113,
       n_12114;
  wire n_12115, n_12116, n_12117, n_12118, n_12119, n_12120, n_12121,
       n_12122;
  wire n_12123, n_12124, n_12125, n_12126, n_12127, n_12128, n_12129,
       n_12130;
  wire n_12131, n_12132, n_12133, n_12134, n_12135, n_12136, n_12137,
       n_12138;
  wire n_12139, n_12140, n_12141, n_12142, n_12143, n_12144, n_12145,
       n_12146;
  wire n_12147, n_12148, n_12149, n_12150, n_12151, n_12152, n_12153,
       n_12154;
  wire n_12155, n_12156, n_12157, n_12158, n_12159, n_12160, n_12161,
       n_12162;
  wire n_12163, n_12164, n_12165, n_12166, n_12167, n_12168, n_12169,
       n_12170;
  wire n_12171, n_12172, n_12173, n_12174, n_12175, n_12176, n_12177,
       n_12178;
  wire n_12179, n_12180, n_12181, n_12182, n_12183, n_12184, n_12185,
       n_12186;
  wire n_12187, n_12188, n_12189, n_12190, n_12191, n_12192, n_12193,
       n_12194;
  wire n_12195, n_12196, n_12197, n_12198, n_12199, n_12200, n_12201,
       n_12202;
  wire n_12203, n_12204, n_12205, n_12206, n_12207, n_12208, n_12209,
       n_12210;
  wire n_12211, n_12212, n_12213, n_12214, n_12215, n_12216, n_12217,
       n_12218;
  wire n_12219, n_12220, n_12221, n_12222, n_12223, n_12224, n_12225,
       n_12226;
  wire n_12227, n_12228, n_12229, n_12230, n_12231, n_12232, n_12233,
       n_12234;
  wire n_12235, n_12236, n_12237, n_12238, n_12239, n_12240, n_12241,
       n_12242;
  wire n_12243, n_12244, n_12245, n_12246, n_12247, n_12248, n_12249,
       n_12250;
  wire n_12251, n_12252, n_12253, n_12254, n_12255, n_12256, n_12257,
       n_12258;
  wire n_12259, n_12260, n_12261, n_12262, n_12263, n_12264, n_12265,
       n_12266;
  wire n_12267, n_12268, n_12269, n_12270, n_12271, n_12272, n_12273,
       n_12274;
  wire n_12275, n_12276, n_12277, n_12278, n_12279, n_12280, n_12281,
       n_12282;
  wire n_12283, n_12284, n_12285, n_12286, n_12287, n_12289, n_12290,
       n_12291;
  wire n_12292, n_12293, n_12294, n_12295, n_12296, n_12297, n_12302,
       n_12303;
  wire n_12304, n_12305, n_12306, n_12307, n_12308, n_12309, n_12310,
       n_12311;
  wire n_12312, n_12313, n_12314, n_12315, n_12316, n_12317, n_12318,
       n_12319;
  wire n_12320, n_12321, n_12322, n_12323, n_12324, n_12325, n_12326,
       n_12327;
  wire n_12328, n_12329, n_12330, n_12331, n_12332, n_12333, n_12334,
       n_12335;
  wire n_12336, n_12337, n_12338, n_12339, n_12340, n_12341, n_12342,
       n_12343;
  wire n_12344, n_12345, n_12346, n_12347, n_12348, n_12349, n_12350,
       n_12351;
  wire n_12352, n_12353, n_12354, n_12355, n_12356, n_12357, n_12358,
       n_12359;
  wire n_12360, n_12361, n_12362, n_12363, n_12364, n_12365, n_12366,
       n_12367;
  wire n_12368, n_12369, n_12370, n_12371, n_12372, n_12373, n_12374,
       n_12375;
  wire n_12376, n_12377, n_12378, n_12379, n_12380, n_12381, n_12382,
       n_12383;
  wire n_12384, n_12385, n_12386, n_12387, n_12388, n_12389, n_12390,
       n_12391;
  wire n_12392, n_12393, n_12394, n_12395, n_12396, n_12397, n_12398,
       n_12399;
  wire n_12400, n_12401, n_12402, n_12403, n_12404, n_12405, n_12406,
       n_12407;
  wire n_12408, n_12409, n_12410, n_12411, n_12412, n_12413, n_12414,
       n_12415;
  wire n_12416, n_12417, n_12418, n_12419, n_12420, n_12421, n_12422,
       n_12423;
  wire n_12424, n_12425, n_12426, n_12427, n_12428, n_12429, n_12430,
       n_12431;
  wire n_12432, n_12433, n_12434, n_12435, n_12436, n_12437, n_12438,
       n_12439;
  wire n_12440, n_12441, n_12442, n_12443, n_12444, n_12445, n_12446,
       n_12447;
  wire n_12448, n_12449, n_12450, n_12451, n_12452, n_12453, n_12454,
       n_12455;
  wire n_12456, n_12457, n_12458, n_12459, n_12460, n_12461, n_12462,
       n_12463;
  wire n_12464, n_12465, n_12466, n_12467, n_12468, n_12469, n_12470,
       n_12471;
  wire n_12472, n_12473, n_12474, n_12475, n_12476, n_12477, n_12478,
       n_12479;
  wire n_12480, n_12481, n_12482, n_12483, n_12484, n_12485, n_12486,
       n_12487;
  wire n_12488, n_12489, n_12490, n_12491, n_12492, n_12493, n_12494,
       n_12495;
  wire n_12496, n_12497, n_12498, n_12499, n_12500, n_12501, n_12502,
       n_12503;
  wire n_12504, n_12505, n_12506, n_12507, n_12508, n_12509, n_12510,
       n_12511;
  wire n_12512, n_12513, n_12514, n_12515, n_12516, n_12517, n_12518,
       n_12519;
  wire n_12520, n_12521, n_12522, n_12523, n_12524, n_12525, n_12526,
       n_12527;
  wire n_12528, n_12529, n_12530, n_12531, n_12532, n_12533, n_12534,
       n_12535;
  wire n_12536, n_12537, n_12538, n_12539, n_12540, n_12541, n_12542,
       n_12543;
  wire n_12544, n_12545, n_12546, n_12547, n_12548, n_12549, n_12550,
       n_12551;
  wire n_12552, n_12553, n_12554, n_12555, n_12556, n_12557, n_12558,
       n_12559;
  wire n_12560, n_12561, n_12562, n_12563, n_12564, n_12565, n_12566,
       n_12567;
  wire n_12568, n_12569, n_12570, n_12571, n_12572, n_12573, n_12574,
       n_12575;
  wire n_12576, n_12577, n_12578, n_12579, n_12580, n_12581, n_12582,
       n_12583;
  wire n_12584, n_12585, n_12586, n_12587, n_12588, n_12589, n_12590,
       n_12591;
  wire n_12592, n_12593, n_12594, n_12595, n_12596, n_12597, n_12598,
       n_12599;
  wire n_12600, n_12601, n_12602, n_12603, n_12604, n_12605, n_12606,
       n_12607;
  wire n_12608, n_12609, n_12610, n_12611, n_12612, n_12613, n_12614,
       n_12615;
  wire n_12616, n_12617, n_12618, n_12619, n_12620, n_12621, n_12622,
       n_12623;
  wire n_12624, n_12625, n_12626, n_12627, n_12628, n_12629, n_12630,
       n_12631;
  wire n_12632, n_12633, n_12634, n_12635, n_12636, n_12637, n_12638,
       n_12639;
  wire n_12640, n_12641, n_12642, n_12643, n_12644, n_12645, n_12646,
       n_12647;
  wire n_12648, n_12649, n_12650, n_12651, n_12652, n_12653, n_12654,
       n_12655;
  wire n_12656, n_12657, n_12658, n_12659, n_12660, n_12661, n_12662,
       n_12663;
  wire n_12664, n_12665, n_12666, n_12667, n_12668, n_12669, n_12670,
       n_12671;
  wire n_12672, n_12673, n_12674, n_12675, n_12676, n_12677, n_12678,
       n_12679;
  wire n_12680, n_12681, n_12682, n_12683, n_12684, n_12685, n_12686,
       n_12687;
  wire n_12688, n_12689, n_12690, n_12691, n_12692, n_12693, n_12694,
       n_12695;
  wire n_12696, n_12697, n_12698, n_12699, n_12700, n_12701, n_12702,
       n_12703;
  wire n_12704, n_12705, n_12706, n_12707, n_12708, n_12709, n_12710,
       n_12711;
  wire n_12712, n_12713, n_12714, n_12715, n_12716, n_12717, n_12718,
       n_12719;
  wire n_12720, n_12721, n_12722, n_12723, n_12724, n_12725, n_12726,
       n_12727;
  wire n_12728, n_12729, n_12730, n_12731, n_12732, n_12733, n_12734,
       n_12735;
  wire n_12737, n_12738, n_12739, n_12740, n_12741, n_12742, n_12743,
       n_12744;
  wire n_12745, n_12750, n_12751, n_12752, n_12753, n_12754, n_12755,
       n_12756;
  wire n_12757, n_12758, n_12759, n_12760, n_12761, n_12762, n_12763,
       n_12764;
  wire n_12765, n_12766, n_12767, n_12768, n_12769, n_12770, n_12771,
       n_12772;
  wire n_12773, n_12774, n_12775, n_12776, n_12777, n_12778, n_12779,
       n_12780;
  wire n_12781, n_12782, n_12783, n_12784, n_12785, n_12786, n_12787,
       n_12788;
  wire n_12789, n_12790, n_12791, n_12792, n_12793, n_12794, n_12795,
       n_12796;
  wire n_12797, n_12798, n_12799, n_12800, n_12801, n_12802, n_12803,
       n_12804;
  wire n_12805, n_12806, n_12807, n_12808, n_12809, n_12810, n_12811,
       n_12812;
  wire n_12813, n_12814, n_12815, n_12816, n_12817, n_12818, n_12819,
       n_12820;
  wire n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827,
       n_12828;
  wire n_12829, n_12830, n_12831, n_12832, n_12833, n_12834, n_12835,
       n_12836;
  wire n_12837, n_12838, n_12839, n_12840, n_12841, n_12842, n_12843,
       n_12844;
  wire n_12845, n_12846, n_12847, n_12848, n_12849, n_12850, n_12851,
       n_12852;
  wire n_12853, n_12854, n_12855, n_12856, n_12857, n_12858, n_12859,
       n_12860;
  wire n_12861, n_12862, n_12863, n_12864, n_12865, n_12866, n_12867,
       n_12868;
  wire n_12869, n_12870, n_12871, n_12872, n_12873, n_12874, n_12875,
       n_12876;
  wire n_12877, n_12878, n_12879, n_12880, n_12881, n_12882, n_12883,
       n_12884;
  wire n_12885, n_12886, n_12887, n_12888, n_12889, n_12890, n_12891,
       n_12892;
  wire n_12893, n_12894, n_12895, n_12896, n_12897, n_12898, n_12899,
       n_12900;
  wire n_12901, n_12902, n_12903, n_12904, n_12905, n_12906, n_12907,
       n_12908;
  wire n_12909, n_12910, n_12911, n_12912, n_12913, n_12914, n_12915,
       n_12916;
  wire n_12917, n_12918, n_12919, n_12920, n_12921, n_12922, n_12923,
       n_12924;
  wire n_12925, n_12926, n_12927, n_12928, n_12929, n_12930, n_12931,
       n_12932;
  wire n_12933, n_12934, n_12935, n_12936, n_12937, n_12938, n_12939,
       n_12940;
  wire n_12941, n_12942, n_12943, n_12944, n_12945, n_12946, n_12947,
       n_12948;
  wire n_12949, n_12950, n_12951, n_12952, n_12953, n_12954, n_12955,
       n_12956;
  wire n_12957, n_12958, n_12959, n_12960, n_12961, n_12962, n_12963,
       n_12964;
  wire n_12965, n_12966, n_12967, n_12968, n_12969, n_12970, n_12971,
       n_12972;
  wire n_12973, n_12974, n_12975, n_12976, n_12977, n_12978, n_12979,
       n_12980;
  wire n_12981, n_12982, n_12983, n_12984, n_12985, n_12986, n_12987,
       n_12988;
  wire n_12989, n_12990, n_12991, n_12992, n_12993, n_12994, n_12995,
       n_12996;
  wire n_12997, n_12998, n_12999, n_13000, n_13001, n_13002, n_13003,
       n_13004;
  wire n_13005, n_13006, n_13007, n_13008, n_13009, n_13010, n_13011,
       n_13012;
  wire n_13013, n_13014, n_13015, n_13016, n_13017, n_13018, n_13019,
       n_13020;
  wire n_13021, n_13022, n_13023, n_13024, n_13025, n_13026, n_13027,
       n_13028;
  wire n_13029, n_13030, n_13031, n_13032, n_13033, n_13034, n_13035,
       n_13036;
  wire n_13037, n_13038, n_13039, n_13040, n_13041, n_13042, n_13043,
       n_13044;
  wire n_13045, n_13046, n_13047, n_13048, n_13049, n_13050, n_13051,
       n_13052;
  wire n_13053, n_13054, n_13055, n_13056, n_13057, n_13058, n_13059,
       n_13060;
  wire n_13061, n_13062, n_13063, n_13064, n_13065, n_13066, n_13067,
       n_13068;
  wire n_13069, n_13070, n_13071, n_13072, n_13073, n_13074, n_13075,
       n_13076;
  wire n_13077, n_13078, n_13079, n_13080, n_13081, n_13082, n_13083,
       n_13084;
  wire n_13085, n_13086, n_13087, n_13088, n_13089, n_13090, n_13091,
       n_13092;
  wire n_13093, n_13094, n_13095, n_13096, n_13097, n_13098, n_13099,
       n_13100;
  wire n_13101, n_13102, n_13103, n_13104, n_13105, n_13106, n_13107,
       n_13108;
  wire n_13109, n_13110, n_13111, n_13112, n_13113, n_13114, n_13115,
       n_13116;
  wire n_13117, n_13118, n_13119, n_13120, n_13121, n_13122, n_13123,
       n_13124;
  wire n_13125, n_13126, n_13127, n_13128, n_13129, n_13130, n_13131,
       n_13132;
  wire n_13133, n_13134, n_13135, n_13136, n_13137, n_13138, n_13139,
       n_13140;
  wire n_13141, n_13142, n_13143, n_13144, n_13145, n_13146, n_13147,
       n_13148;
  wire n_13149, n_13150, n_13151, n_13152, n_13153, n_13154, n_13155,
       n_13156;
  wire n_13157, n_13158, n_13159, n_13160, n_13161, n_13162, n_13163,
       n_13164;
  wire n_13165, n_13166, n_13167, n_13168, n_13169, n_13170, n_13171,
       n_13172;
  wire n_13173, n_13174, n_13175, n_13176, n_13177, n_13178, n_13179,
       n_13180;
  wire n_13181, n_13182, n_13183, n_13184, n_13185, n_13186, n_13187,
       n_13188;
  wire n_13189, n_13190, n_13191, n_13193, n_13194, n_13195, n_13196,
       n_13197;
  wire n_13198, n_13199, n_13200, n_13201, n_13206, n_13207, n_13208,
       n_13209;
  wire n_13210, n_13211, n_13212, n_13213, n_13214, n_13215, n_13216,
       n_13217;
  wire n_13218, n_13219, n_13220, n_13221, n_13222, n_13223, n_13224,
       n_13225;
  wire n_13226, n_13227, n_13228, n_13229, n_13230, n_13231, n_13232,
       n_13233;
  wire n_13234, n_13235, n_13236, n_13237, n_13238, n_13239, n_13240,
       n_13241;
  wire n_13242, n_13243, n_13244, n_13245, n_13246, n_13247, n_13248,
       n_13249;
  wire n_13250, n_13251, n_13252, n_13253, n_13254, n_13255, n_13256,
       n_13257;
  wire n_13258, n_13259, n_13260, n_13261, n_13262, n_13263, n_13264,
       n_13265;
  wire n_13266, n_13267, n_13268, n_13269, n_13270, n_13271, n_13272,
       n_13273;
  wire n_13274, n_13275, n_13276, n_13277, n_13278, n_13279, n_13280,
       n_13281;
  wire n_13282, n_13283, n_13284, n_13285, n_13286, n_13287, n_13288,
       n_13289;
  wire n_13290, n_13291, n_13292, n_13293, n_13294, n_13295, n_13296,
       n_13297;
  wire n_13298, n_13299, n_13300, n_13301, n_13302, n_13303, n_13304,
       n_13305;
  wire n_13306, n_13307, n_13308, n_13309, n_13310, n_13311, n_13312,
       n_13313;
  wire n_13314, n_13315, n_13316, n_13317, n_13318, n_13319, n_13320,
       n_13321;
  wire n_13322, n_13323, n_13324, n_13325, n_13326, n_13327, n_13328,
       n_13329;
  wire n_13330, n_13331, n_13332, n_13333, n_13334, n_13335, n_13336,
       n_13337;
  wire n_13338, n_13339, n_13340, n_13341, n_13342, n_13343, n_13344,
       n_13345;
  wire n_13346, n_13347, n_13348, n_13349, n_13350, n_13351, n_13352,
       n_13353;
  wire n_13354, n_13355, n_13356, n_13357, n_13358, n_13359, n_13360,
       n_13361;
  wire n_13362, n_13363, n_13364, n_13365, n_13366, n_13367, n_13368,
       n_13369;
  wire n_13370, n_13371, n_13372, n_13373, n_13374, n_13375, n_13376,
       n_13377;
  wire n_13378, n_13379, n_13380, n_13381, n_13382, n_13383, n_13384,
       n_13385;
  wire n_13386, n_13387, n_13388, n_13389, n_13390, n_13391, n_13392,
       n_13393;
  wire n_13394, n_13395, n_13396, n_13397, n_13398, n_13399, n_13400,
       n_13401;
  wire n_13402, n_13403, n_13404, n_13405, n_13406, n_13407, n_13408,
       n_13409;
  wire n_13410, n_13411, n_13412, n_13413, n_13414, n_13415, n_13416,
       n_13417;
  wire n_13418, n_13419, n_13420, n_13421, n_13422, n_13423, n_13424,
       n_13425;
  wire n_13426, n_13427, n_13428, n_13429, n_13430, n_13431, n_13432,
       n_13433;
  wire n_13434, n_13435, n_13436, n_13437, n_13438, n_13439, n_13440,
       n_13441;
  wire n_13442, n_13443, n_13444, n_13445, n_13446, n_13447, n_13448,
       n_13449;
  wire n_13450, n_13451, n_13452, n_13453, n_13454, n_13455, n_13456,
       n_13457;
  wire n_13458, n_13459, n_13460, n_13461, n_13462, n_13463, n_13464,
       n_13465;
  wire n_13466, n_13467, n_13468, n_13469, n_13470, n_13471, n_13472,
       n_13473;
  wire n_13474, n_13475, n_13476, n_13477, n_13478, n_13479, n_13480,
       n_13481;
  wire n_13482, n_13483, n_13484, n_13485, n_13486, n_13487, n_13488,
       n_13489;
  wire n_13490, n_13491, n_13492, n_13493, n_13494, n_13495, n_13496,
       n_13497;
  wire n_13498, n_13499, n_13500, n_13501, n_13502, n_13503, n_13504,
       n_13505;
  wire n_13506, n_13507, n_13508, n_13509, n_13510, n_13511, n_13512,
       n_13513;
  wire n_13514, n_13515, n_13516, n_13517, n_13518, n_13519, n_13520,
       n_13521;
  wire n_13522, n_13523, n_13524, n_13525, n_13526, n_13527, n_13528,
       n_13529;
  wire n_13530, n_13531, n_13532, n_13533, n_13534, n_13535, n_13536,
       n_13537;
  wire n_13538, n_13539, n_13540, n_13541, n_13542, n_13543, n_13544,
       n_13545;
  wire n_13546, n_13547, n_13548, n_13549, n_13550, n_13551, n_13552,
       n_13553;
  wire n_13554, n_13555, n_13556, n_13557, n_13558, n_13559, n_13560,
       n_13561;
  wire n_13562, n_13563, n_13564, n_13565, n_13566, n_13567, n_13568,
       n_13569;
  wire n_13570, n_13571, n_13572, n_13573, n_13574, n_13575, n_13576,
       n_13577;
  wire n_13578, n_13579, n_13580, n_13581, n_13582, n_13583, n_13584,
       n_13585;
  wire n_13586, n_13587, n_13588, n_13589, n_13590, n_13591, n_13592,
       n_13593;
  wire n_13594, n_13595, n_13596, n_13597, n_13598, n_13599, n_13600,
       n_13601;
  wire n_13602, n_13603, n_13604, n_13605, n_13606, n_13607, n_13608,
       n_13609;
  wire n_13610, n_13611, n_13612, n_13613, n_13614, n_13615, n_13616,
       n_13617;
  wire n_13618, n_13619, n_13620, n_13621, n_13622, n_13623, n_13624,
       n_13625;
  wire n_13626, n_13627, n_13628, n_13629, n_13630, n_13631, n_13632,
       n_13633;
  wire n_13634, n_13635, n_13636, n_13637, n_13638, n_13639, n_13640,
       n_13641;
  wire n_13642, n_13643, n_13644, n_13645, n_13646, n_13647, n_13648,
       n_13649;
  wire n_13650, n_13651, n_13652, n_13653, n_13654, n_13655, n_13657,
       n_13658;
  wire n_13659, n_13660, n_13661, n_13662, n_13663, n_13664, n_13665,
       n_13670;
  wire n_13671, n_13672, n_13673, n_13674, n_13675, n_13676, n_13677,
       n_13678;
  wire n_13679, n_13680, n_13681, n_13682, n_13683, n_13684, n_13685,
       n_13686;
  wire n_13687, n_13688, n_13689, n_13690, n_13691, n_13692, n_13693,
       n_13694;
  wire n_13695, n_13696, n_13697, n_13698, n_13699, n_13700, n_13701,
       n_13702;
  wire n_13703, n_13704, n_13705, n_13706, n_13707, n_13708, n_13709,
       n_13710;
  wire n_13711, n_13712, n_13713, n_13714, n_13715, n_13716, n_13717,
       n_13718;
  wire n_13719, n_13720, n_13721, n_13722, n_13723, n_13724, n_13725,
       n_13726;
  wire n_13727, n_13728, n_13729, n_13730, n_13731, n_13732, n_13733,
       n_13734;
  wire n_13735, n_13736, n_13737, n_13738, n_13739, n_13740, n_13741,
       n_13742;
  wire n_13743, n_13744, n_13745, n_13746, n_13747, n_13748, n_13749,
       n_13750;
  wire n_13751, n_13752, n_13753, n_13754, n_13755, n_13756, n_13757,
       n_13758;
  wire n_13759, n_13760, n_13761, n_13762, n_13763, n_13764, n_13765,
       n_13766;
  wire n_13767, n_13768, n_13769, n_13770, n_13771, n_13772, n_13773,
       n_13774;
  wire n_13775, n_13776, n_13777, n_13778, n_13779, n_13780, n_13781,
       n_13782;
  wire n_13783, n_13784, n_13785, n_13786, n_13787, n_13788, n_13789,
       n_13790;
  wire n_13791, n_13792, n_13793, n_13794, n_13795, n_13796, n_13797,
       n_13798;
  wire n_13799, n_13800, n_13801, n_13802, n_13803, n_13804, n_13805,
       n_13806;
  wire n_13807, n_13808, n_13809, n_13810, n_13811, n_13812, n_13813,
       n_13814;
  wire n_13815, n_13816, n_13817, n_13818, n_13819, n_13820, n_13821,
       n_13822;
  wire n_13823, n_13824, n_13825, n_13826, n_13827, n_13828, n_13829,
       n_13830;
  wire n_13831, n_13832, n_13833, n_13834, n_13835, n_13836, n_13837,
       n_13838;
  wire n_13839, n_13840, n_13841, n_13842, n_13843, n_13844, n_13845,
       n_13846;
  wire n_13847, n_13848, n_13849, n_13850, n_13851, n_13852, n_13853,
       n_13854;
  wire n_13855, n_13856, n_13857, n_13858, n_13859, n_13860, n_13861,
       n_13862;
  wire n_13863, n_13864, n_13865, n_13866, n_13867, n_13868, n_13869,
       n_13870;
  wire n_13871, n_13872, n_13873, n_13874, n_13875, n_13876, n_13877,
       n_13878;
  wire n_13879, n_13880, n_13881, n_13882, n_13883, n_13884, n_13885,
       n_13886;
  wire n_13887, n_13888, n_13889, n_13890, n_13891, n_13892, n_13893,
       n_13894;
  wire n_13895, n_13896, n_13897, n_13898, n_13899, n_13900, n_13901,
       n_13902;
  wire n_13903, n_13904, n_13905, n_13906, n_13907, n_13908, n_13909,
       n_13910;
  wire n_13911, n_13912, n_13913, n_13914, n_13915, n_13916, n_13917,
       n_13918;
  wire n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925,
       n_13926;
  wire n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933,
       n_13934;
  wire n_13935, n_13936, n_13937, n_13938, n_13939, n_13940, n_13941,
       n_13942;
  wire n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949,
       n_13950;
  wire n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957,
       n_13958;
  wire n_13959, n_13960, n_13961, n_13962, n_13963, n_13964, n_13965,
       n_13966;
  wire n_13967, n_13968, n_13969, n_13970, n_13971, n_13972, n_13973,
       n_13974;
  wire n_13975, n_13976, n_13977, n_13978, n_13979, n_13980, n_13981,
       n_13982;
  wire n_13983, n_13984, n_13985, n_13986, n_13987, n_13988, n_13989,
       n_13990;
  wire n_13991, n_13992, n_13993, n_13994, n_13995, n_13996, n_13997,
       n_13998;
  wire n_13999, n_14000, n_14001, n_14002, n_14003, n_14004, n_14005,
       n_14006;
  wire n_14007, n_14008, n_14009, n_14010, n_14011, n_14012, n_14013,
       n_14014;
  wire n_14015, n_14016, n_14017, n_14018, n_14019, n_14020, n_14021,
       n_14022;
  wire n_14023, n_14024, n_14025, n_14026, n_14027, n_14028, n_14029,
       n_14030;
  wire n_14031, n_14032, n_14033, n_14034, n_14035, n_14036, n_14037,
       n_14038;
  wire n_14039, n_14040, n_14041, n_14042, n_14043, n_14044, n_14045,
       n_14046;
  wire n_14047, n_14048, n_14049, n_14050, n_14051, n_14052, n_14053,
       n_14054;
  wire n_14055, n_14056, n_14057, n_14058, n_14059, n_14060, n_14061,
       n_14062;
  wire n_14063, n_14064, n_14065, n_14066, n_14067, n_14068, n_14069,
       n_14070;
  wire n_14071, n_14072, n_14073, n_14074, n_14075, n_14076, n_14077,
       n_14078;
  wire n_14079, n_14080, n_14081, n_14082, n_14083, n_14084, n_14085,
       n_14086;
  wire n_14087, n_14088, n_14089, n_14090, n_14091, n_14092, n_14093,
       n_14094;
  wire n_14095, n_14096, n_14097, n_14098, n_14099, n_14100, n_14101,
       n_14102;
  wire n_14103, n_14104, n_14105, n_14106, n_14107, n_14108, n_14109,
       n_14110;
  wire n_14111, n_14112, n_14113, n_14114, n_14115, n_14116, n_14117,
       n_14118;
  wire n_14119, n_14120, n_14121, n_14122, n_14123, n_14124, n_14125,
       n_14126;
  wire n_14127, n_14129, n_14130, n_14131, n_14132, n_14133, n_14134,
       n_14135;
  wire n_14136, n_14137, n_14141, n_14142, n_14143, n_14144, n_14145,
       n_14146;
  wire n_14147, n_14148, n_14149, n_14150, n_14151, n_14152, n_14153,
       n_14154;
  wire n_14155, n_14156, n_14157, n_14158, n_14159, n_14160, n_14161,
       n_14162;
  wire n_14163, n_14164, n_14165, n_14166, n_14167, n_14168, n_14169,
       n_14170;
  wire n_14171, n_14172, n_14173, n_14174, n_14175, n_14176, n_14177,
       n_14178;
  wire n_14179, n_14180, n_14181, n_14182, n_14183, n_14184, n_14185,
       n_14186;
  wire n_14187, n_14188, n_14189, n_14190, n_14191, n_14192, n_14193,
       n_14194;
  wire n_14195, n_14196, n_14197, n_14198, n_14199, n_14200, n_14201,
       n_14202;
  wire n_14203, n_14204, n_14205, n_14206, n_14207, n_14208, n_14209,
       n_14210;
  wire n_14211, n_14212, n_14213, n_14214, n_14215, n_14216, n_14217,
       n_14218;
  wire n_14219, n_14220, n_14221, n_14222, n_14223, n_14224, n_14225,
       n_14226;
  wire n_14227, n_14228, n_14229, n_14230, n_14231, n_14232, n_14233,
       n_14234;
  wire n_14235, n_14236, n_14237, n_14238, n_14239, n_14240, n_14241,
       n_14242;
  wire n_14243, n_14244, n_14245, n_14246, n_14247, n_14248, n_14249,
       n_14250;
  wire n_14251, n_14252, n_14253, n_14254, n_14255, n_14256, n_14257,
       n_14258;
  wire n_14259, n_14260, n_14261, n_14262, n_14263, n_14264, n_14265,
       n_14266;
  wire n_14267, n_14268, n_14269, n_14270, n_14271, n_14272, n_14273,
       n_14274;
  wire n_14275, n_14276, n_14277, n_14278, n_14279, n_14280, n_14281,
       n_14282;
  wire n_14283, n_14284, n_14285, n_14286, n_14287, n_14288, n_14289,
       n_14290;
  wire n_14291, n_14292, n_14293, n_14294, n_14295, n_14296, n_14297,
       n_14298;
  wire n_14299, n_14300, n_14301, n_14302, n_14303, n_14304, n_14305,
       n_14306;
  wire n_14307, n_14308, n_14309, n_14310, n_14311, n_14312, n_14313,
       n_14314;
  wire n_14315, n_14316, n_14317, n_14318, n_14319, n_14320, n_14321,
       n_14322;
  wire n_14323, n_14324, n_14325, n_14326, n_14327, n_14328, n_14329,
       n_14330;
  wire n_14331, n_14332, n_14333, n_14334, n_14335, n_14336, n_14337,
       n_14338;
  wire n_14339, n_14340, n_14341, n_14342, n_14343, n_14344, n_14345,
       n_14346;
  wire n_14347, n_14348, n_14349, n_14350, n_14351, n_14352, n_14353,
       n_14354;
  wire n_14355, n_14356, n_14357, n_14358, n_14359, n_14360, n_14361,
       n_14362;
  wire n_14363, n_14364, n_14365, n_14366, n_14367, n_14368, n_14369,
       n_14370;
  wire n_14371, n_14372, n_14373, n_14374, n_14375, n_14376, n_14377,
       n_14378;
  wire n_14379, n_14380, n_14381, n_14382, n_14383, n_14384, n_14385,
       n_14386;
  wire n_14387, n_14388, n_14389, n_14390, n_14391, n_14392, n_14393,
       n_14394;
  wire n_14395, n_14396, n_14397, n_14398, n_14399, n_14400, n_14401,
       n_14402;
  wire n_14403, n_14404, n_14405, n_14406, n_14407, n_14408, n_14409,
       n_14410;
  wire n_14411, n_14412, n_14413, n_14414, n_14415, n_14416, n_14417,
       n_14418;
  wire n_14419, n_14420, n_14421, n_14422, n_14423, n_14424, n_14425,
       n_14426;
  wire n_14427, n_14428, n_14429, n_14430, n_14431, n_14432, n_14433,
       n_14434;
  wire n_14435, n_14436, n_14437, n_14438, n_14439, n_14440, n_14441,
       n_14442;
  wire n_14443, n_14444, n_14445, n_14446, n_14447, n_14448, n_14449,
       n_14450;
  wire n_14451, n_14452, n_14453, n_14454, n_14455, n_14456, n_14457,
       n_14458;
  wire n_14459, n_14460, n_14461, n_14462, n_14463, n_14464, n_14465,
       n_14466;
  wire n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, n_14473,
       n_14474;
  wire n_14475, n_14476, n_14477, n_14478, n_14479, n_14480, n_14481,
       n_14482;
  wire n_14483, n_14484, n_14485, n_14486, n_14487, n_14488, n_14489,
       n_14490;
  wire n_14491, n_14492, n_14493, n_14494, n_14495, n_14496, n_14497,
       n_14498;
  wire n_14499, n_14500, n_14501, n_14502, n_14503, n_14504, n_14505,
       n_14506;
  wire n_14507, n_14508, n_14509, n_14510, n_14511, n_14512, n_14513,
       n_14514;
  wire n_14515, n_14516, n_14517, n_14518, n_14519, n_14520, n_14521,
       n_14522;
  wire n_14523, n_14524, n_14525, n_14526, n_14527, n_14528, n_14529,
       n_14530;
  wire n_14531, n_14532, n_14533, n_14534, n_14535, n_14536, n_14537,
       n_14538;
  wire n_14539, n_14540, n_14541, n_14542, n_14543, n_14544, n_14545,
       n_14546;
  wire n_14547, n_14548, n_14549, n_14550, n_14551, n_14552, n_14553,
       n_14554;
  wire n_14555, n_14556, n_14557, n_14558, n_14559, n_14560, n_14561,
       n_14562;
  wire n_14563, n_14564, n_14565, n_14566, n_14567, n_14568, n_14569,
       n_14570;
  wire n_14571, n_14572, n_14573, n_14574, n_14575, n_14576, n_14577,
       n_14578;
  wire n_14579, n_14580, n_14581, n_14582, n_14583, n_14584, n_14585,
       n_14586;
  wire n_14587, n_14588, n_14589, n_14590, n_14591, n_14592, n_14593,
       n_14594;
  wire n_14595, n_14596, n_14597, n_14598, n_14599, n_14600, n_14601,
       n_14602;
  wire n_14603, n_14604, n_14605, n_14606, n_14608, n_14609, n_14610,
       n_14611;
  wire n_14612, n_14613, n_14614, n_14615, n_14616, n_14620, n_14621,
       n_14622;
  wire n_14623, n_14624, n_14625, n_14626, n_14627, n_14628, n_14629,
       n_14630;
  wire n_14631, n_14632, n_14633, n_14634, n_14635, n_14636, n_14637,
       n_14638;
  wire n_14639, n_14640, n_14641, n_14642, n_14643, n_14644, n_14645,
       n_14646;
  wire n_14647, n_14648, n_14649, n_14650, n_14651, n_14652, n_14653,
       n_14654;
  wire n_14655, n_14656, n_14657, n_14658, n_14659, n_14660, n_14661,
       n_14662;
  wire n_14663, n_14664, n_14665, n_14666, n_14667, n_14668, n_14669,
       n_14670;
  wire n_14671, n_14672, n_14673, n_14674, n_14675, n_14676, n_14677,
       n_14678;
  wire n_14679, n_14680, n_14681, n_14682, n_14683, n_14684, n_14685,
       n_14686;
  wire n_14687, n_14688, n_14689, n_14690, n_14691, n_14692, n_14693,
       n_14694;
  wire n_14695, n_14696, n_14697, n_14698, n_14699, n_14700, n_14701,
       n_14702;
  wire n_14703, n_14704, n_14705, n_14706, n_14707, n_14708, n_14709,
       n_14710;
  wire n_14711, n_14712, n_14713, n_14714, n_14715, n_14716, n_14717,
       n_14718;
  wire n_14719, n_14720, n_14721, n_14722, n_14723, n_14724, n_14725,
       n_14726;
  wire n_14727, n_14728, n_14729, n_14730, n_14731, n_14732, n_14733,
       n_14734;
  wire n_14735, n_14736, n_14737, n_14738, n_14739, n_14740, n_14741,
       n_14742;
  wire n_14743, n_14744, n_14745, n_14746, n_14747, n_14748, n_14749,
       n_14750;
  wire n_14751, n_14752, n_14753, n_14754, n_14755, n_14756, n_14757,
       n_14758;
  wire n_14759, n_14760, n_14761, n_14762, n_14763, n_14764, n_14765,
       n_14766;
  wire n_14767, n_14768, n_14769, n_14770, n_14771, n_14772, n_14773,
       n_14774;
  wire n_14775, n_14776, n_14777, n_14778, n_14779, n_14780, n_14781,
       n_14782;
  wire n_14783, n_14784, n_14785, n_14786, n_14787, n_14788, n_14789,
       n_14790;
  wire n_14791, n_14792, n_14793, n_14794, n_14795, n_14796, n_14797,
       n_14798;
  wire n_14799, n_14800, n_14801, n_14802, n_14803, n_14804, n_14805,
       n_14806;
  wire n_14807, n_14808, n_14809, n_14810, n_14811, n_14812, n_14813,
       n_14814;
  wire n_14815, n_14816, n_14817, n_14818, n_14819, n_14820, n_14821,
       n_14822;
  wire n_14823, n_14824, n_14825, n_14826, n_14827, n_14828, n_14829,
       n_14830;
  wire n_14831, n_14832, n_14833, n_14834, n_14835, n_14836, n_14837,
       n_14838;
  wire n_14839, n_14840, n_14841, n_14842, n_14843, n_14844, n_14845,
       n_14846;
  wire n_14847, n_14848, n_14849, n_14850, n_14851, n_14852, n_14853,
       n_14854;
  wire n_14855, n_14856, n_14857, n_14858, n_14859, n_14860, n_14861,
       n_14862;
  wire n_14863, n_14864, n_14865, n_14866, n_14867, n_14868, n_14869,
       n_14870;
  wire n_14871, n_14872, n_14873, n_14874, n_14875, n_14876, n_14877,
       n_14878;
  wire n_14879, n_14880, n_14881, n_14882, n_14883, n_14884, n_14885,
       n_14886;
  wire n_14887, n_14888, n_14889, n_14890, n_14891, n_14892, n_14893,
       n_14894;
  wire n_14895, n_14896, n_14897, n_14898, n_14899, n_14900, n_14901,
       n_14902;
  wire n_14903, n_14904, n_14905, n_14906, n_14907, n_14908, n_14909,
       n_14910;
  wire n_14911, n_14912, n_14913, n_14914, n_14915, n_14916, n_14917,
       n_14918;
  wire n_14919, n_14920, n_14921, n_14922, n_14923, n_14924, n_14925,
       n_14926;
  wire n_14927, n_14928, n_14929, n_14930, n_14931, n_14932, n_14933,
       n_14934;
  wire n_14935, n_14936, n_14937, n_14938, n_14939, n_14940, n_14941,
       n_14942;
  wire n_14943, n_14944, n_14945, n_14946, n_14947, n_14948, n_14949,
       n_14950;
  wire n_14951, n_14952, n_14953, n_14954, n_14955, n_14956, n_14957,
       n_14958;
  wire n_14959, n_14960, n_14961, n_14962, n_14963, n_14964, n_14965,
       n_14966;
  wire n_14967, n_14968, n_14969, n_14970, n_14971, n_14972, n_14973,
       n_14974;
  wire n_14975, n_14976, n_14977, n_14978, n_14979, n_14980, n_14981,
       n_14982;
  wire n_14983, n_14984, n_14985, n_14986, n_14987, n_14988, n_14989,
       n_14990;
  wire n_14991, n_14992, n_14993, n_14994, n_14995, n_14996, n_14997,
       n_14998;
  wire n_14999, n_15000, n_15001, n_15002, n_15003, n_15004, n_15005,
       n_15006;
  wire n_15007, n_15008, n_15009, n_15010, n_15011, n_15012, n_15013,
       n_15014;
  wire n_15015, n_15016, n_15017, n_15018, n_15019, n_15020, n_15021,
       n_15022;
  wire n_15023, n_15024, n_15025, n_15026, n_15027, n_15028, n_15029,
       n_15030;
  wire n_15031, n_15032, n_15033, n_15034, n_15035, n_15036, n_15037,
       n_15038;
  wire n_15039, n_15040, n_15041, n_15042, n_15043, n_15044, n_15045,
       n_15046;
  wire n_15047, n_15048, n_15049, n_15050, n_15051, n_15052, n_15053,
       n_15054;
  wire n_15055, n_15056, n_15057, n_15058, n_15059, n_15060, n_15061,
       n_15062;
  wire n_15063, n_15064, n_15065, n_15066, n_15067, n_15068, n_15069,
       n_15070;
  wire n_15071, n_15072, n_15073, n_15074, n_15075, n_15076, n_15077,
       n_15078;
  wire n_15079, n_15080, n_15081, n_15082, n_15083, n_15084, n_15085,
       n_15086;
  wire n_15087, n_15088, n_15089, n_15090, n_15091, n_15092, n_15093,
       n_15095;
  wire n_15096, n_15097, n_15098, n_15099, n_15100, n_15101, n_15102,
       n_15103;
  wire n_15107, n_15108, n_15109, n_15110, n_15111, n_15112, n_15113,
       n_15114;
  wire n_15115, n_15116, n_15117, n_15118, n_15119, n_15120, n_15121,
       n_15122;
  wire n_15123, n_15124, n_15125, n_15126, n_15127, n_15128, n_15129,
       n_15130;
  wire n_15131, n_15132, n_15133, n_15134, n_15135, n_15136, n_15137,
       n_15138;
  wire n_15139, n_15140, n_15141, n_15142, n_15143, n_15144, n_15145,
       n_15146;
  wire n_15147, n_15148, n_15149, n_15150, n_15151, n_15152, n_15153,
       n_15154;
  wire n_15155, n_15156, n_15157, n_15158, n_15159, n_15160, n_15161,
       n_15162;
  wire n_15163, n_15164, n_15165, n_15166, n_15167, n_15168, n_15169,
       n_15170;
  wire n_15171, n_15172, n_15173, n_15174, n_15175, n_15176, n_15177,
       n_15178;
  wire n_15179, n_15180, n_15181, n_15182, n_15183, n_15184, n_15185,
       n_15186;
  wire n_15187, n_15188, n_15189, n_15190, n_15191, n_15192, n_15193,
       n_15194;
  wire n_15195, n_15196, n_15197, n_15198, n_15199, n_15200, n_15201,
       n_15202;
  wire n_15203, n_15204, n_15205, n_15206, n_15207, n_15208, n_15209,
       n_15210;
  wire n_15211, n_15212, n_15213, n_15214, n_15215, n_15216, n_15217,
       n_15218;
  wire n_15219, n_15220, n_15221, n_15222, n_15223, n_15224, n_15225,
       n_15226;
  wire n_15227, n_15228, n_15229, n_15230, n_15231, n_15232, n_15233,
       n_15234;
  wire n_15235, n_15236, n_15237, n_15238, n_15239, n_15240, n_15241,
       n_15242;
  wire n_15243, n_15244, n_15245, n_15246, n_15247, n_15248, n_15249,
       n_15250;
  wire n_15251, n_15252, n_15253, n_15254, n_15255, n_15256, n_15257,
       n_15258;
  wire n_15259, n_15260, n_15261, n_15262, n_15263, n_15264, n_15265,
       n_15266;
  wire n_15267, n_15268, n_15269, n_15270, n_15271, n_15272, n_15273,
       n_15274;
  wire n_15275, n_15276, n_15277, n_15278, n_15279, n_15280, n_15281,
       n_15282;
  wire n_15283, n_15284, n_15285, n_15286, n_15287, n_15288, n_15289,
       n_15290;
  wire n_15291, n_15292, n_15293, n_15294, n_15295, n_15296, n_15297,
       n_15298;
  wire n_15299, n_15300, n_15301, n_15302, n_15303, n_15304, n_15305,
       n_15306;
  wire n_15307, n_15308, n_15309, n_15310, n_15311, n_15312, n_15313,
       n_15314;
  wire n_15315, n_15316, n_15317, n_15318, n_15319, n_15320, n_15321,
       n_15322;
  wire n_15323, n_15324, n_15325, n_15326, n_15327, n_15328, n_15329,
       n_15330;
  wire n_15331, n_15332, n_15333, n_15334, n_15335, n_15336, n_15337,
       n_15338;
  wire n_15339, n_15340, n_15341, n_15342, n_15343, n_15344, n_15345,
       n_15346;
  wire n_15347, n_15348, n_15349, n_15350, n_15351, n_15352, n_15353,
       n_15354;
  wire n_15355, n_15356, n_15357, n_15358, n_15359, n_15360, n_15361,
       n_15362;
  wire n_15363, n_15364, n_15365, n_15366, n_15367, n_15368, n_15369,
       n_15370;
  wire n_15371, n_15372, n_15373, n_15374, n_15375, n_15376, n_15377,
       n_15378;
  wire n_15379, n_15380, n_15381, n_15382, n_15383, n_15384, n_15385,
       n_15386;
  wire n_15387, n_15388, n_15389, n_15390, n_15391, n_15392, n_15393,
       n_15394;
  wire n_15395, n_15396, n_15397, n_15398, n_15399, n_15400, n_15401,
       n_15402;
  wire n_15403, n_15404, n_15405, n_15406, n_15407, n_15408, n_15409,
       n_15410;
  wire n_15411, n_15412, n_15413, n_15414, n_15415, n_15416, n_15417,
       n_15418;
  wire n_15419, n_15420, n_15421, n_15422, n_15423, n_15424, n_15425,
       n_15426;
  wire n_15427, n_15428, n_15429, n_15430, n_15431, n_15432, n_15433,
       n_15434;
  wire n_15435, n_15436, n_15437, n_15438, n_15439, n_15440, n_15441,
       n_15442;
  wire n_15443, n_15444, n_15445, n_15446, n_15447, n_15448, n_15449,
       n_15450;
  wire n_15451, n_15452, n_15453, n_15454, n_15455, n_15456, n_15457,
       n_15458;
  wire n_15459, n_15460, n_15461, n_15462, n_15463, n_15464, n_15465,
       n_15466;
  wire n_15467, n_15468, n_15469, n_15470, n_15471, n_15472, n_15473,
       n_15474;
  wire n_15475, n_15476, n_15477, n_15478, n_15479, n_15480, n_15481,
       n_15482;
  wire n_15483, n_15484, n_15485, n_15486, n_15487, n_15488, n_15489,
       n_15490;
  wire n_15491, n_15492, n_15493, n_15494, n_15495, n_15496, n_15497,
       n_15498;
  wire n_15499, n_15500, n_15501, n_15502, n_15503, n_15504, n_15505,
       n_15506;
  wire n_15507, n_15508, n_15509, n_15510, n_15511, n_15512, n_15513,
       n_15514;
  wire n_15515, n_15516, n_15517, n_15518, n_15519, n_15520, n_15521,
       n_15522;
  wire n_15523, n_15524, n_15525, n_15526, n_15527, n_15528, n_15529,
       n_15530;
  wire n_15531, n_15532, n_15533, n_15534, n_15535, n_15536, n_15537,
       n_15538;
  wire n_15539, n_15540, n_15541, n_15542, n_15543, n_15544, n_15545,
       n_15546;
  wire n_15547, n_15548, n_15549, n_15550, n_15551, n_15552, n_15553,
       n_15554;
  wire n_15555, n_15556, n_15557, n_15558, n_15559, n_15560, n_15561,
       n_15562;
  wire n_15563, n_15564, n_15565, n_15566, n_15567, n_15568, n_15569,
       n_15570;
  wire n_15571, n_15572, n_15573, n_15574, n_15575, n_15576, n_15577,
       n_15578;
  wire n_15579, n_15580, n_15581, n_15582, n_15583, n_15584, n_15585,
       n_15586;
  wire n_15587, n_15588, n_15590, n_15591, n_15592, n_15593, n_15594,
       n_15595;
  wire n_15596, n_15597, n_15598, n_15600, n_15601, n_15602, n_15605,
       n_15606;
  wire n_15607, n_15608, n_15609, n_15610, n_15611, n_15612, n_15613,
       n_15614;
  wire n_15615, n_15616, n_15617, n_15619, n_15620, n_15621, n_15622,
       n_15623;
  wire n_15624, n_15625, n_15626, n_15627, n_15628, n_15629, n_15630,
       n_15631;
  wire n_15632, n_15633, n_15634, n_15635, n_15636, n_15637, n_15638,
       n_15639;
  wire n_15640, n_15641, n_15642, n_15643, n_15644, n_15645, n_15646,
       n_15647;
  wire n_15648, n_15649, n_15650, n_15651, n_15652, n_15653, n_15654,
       n_15655;
  wire n_15656, n_15657, n_15658, n_15659, n_15660, n_15661, n_15662,
       n_15663;
  wire n_15664, n_15665, n_15666, n_15667, n_15668, n_15669, n_15670,
       n_15671;
  wire n_15672, n_15673, n_15674, n_15675, n_15676, n_15677, n_15678,
       n_15679;
  wire n_15680, n_15681, n_15682, n_15683, n_15684, n_15685, n_15686,
       n_15687;
  wire n_15688, n_15689, n_15690, n_15691, n_15692, n_15693, n_15694,
       n_15695;
  wire n_15696, n_15697, n_15698, n_15699, n_15700, n_15701, n_15702,
       n_15703;
  wire n_15704, n_15705, n_15706, n_15707, n_15708, n_15709, n_15710,
       n_15711;
  wire n_15712, n_15713, n_15714, n_15715, n_15716, n_15717, n_15718,
       n_15719;
  wire n_15720, n_15721, n_15722, n_15723, n_15724, n_15725, n_15726,
       n_15727;
  wire n_15728, n_15729, n_15730, n_15731, n_15732, n_15733, n_15734,
       n_15735;
  wire n_15736, n_15737, n_15738, n_15739, n_15740, n_15741, n_15742,
       n_15743;
  wire n_15744, n_15745, n_15746, n_15747, n_15748, n_15749, n_15750,
       n_15751;
  wire n_15752, n_15753, n_15754, n_15755, n_15756, n_15757, n_15758,
       n_15759;
  wire n_15760, n_15761, n_15762, n_15763, n_15764, n_15765, n_15766,
       n_15767;
  wire n_15768, n_15769, n_15770, n_15771, n_15772, n_15773, n_15774,
       n_15775;
  wire n_15776, n_15777, n_15778, n_15779, n_15780, n_15781, n_15782,
       n_15783;
  wire n_15784, n_15785, n_15786, n_15787, n_15788, n_15789, n_15790,
       n_15791;
  wire n_15792, n_15793, n_15794, n_15795, n_15796, n_15797, n_15798,
       n_15799;
  wire n_15800, n_15801, n_15802, n_15803, n_15804, n_15805, n_15806,
       n_15807;
  wire n_15808, n_15809, n_15810, n_15811, n_15812, n_15813, n_15814,
       n_15815;
  wire n_15816, n_15817, n_15818, n_15819, n_15820, n_15821, n_15822,
       n_15823;
  wire n_15824, n_15825, n_15826, n_15827, n_15828, n_15829, n_15830,
       n_15831;
  wire n_15832, n_15833, n_15834, n_15835, n_15836, n_15837, n_15838,
       n_15839;
  wire n_15840, n_15841, n_15842, n_15843, n_15844, n_15845, n_15846,
       n_15847;
  wire n_15848, n_15849, n_15850, n_15851, n_15852, n_15853, n_15854,
       n_15855;
  wire n_15856, n_15857, n_15858, n_15859, n_15860, n_15861, n_15862,
       n_15863;
  wire n_15864, n_15865, n_15866, n_15867, n_15868, n_15869, n_15870,
       n_15871;
  wire n_15872, n_15873, n_15874, n_15875, n_15876, n_15877, n_15878,
       n_15879;
  wire n_15880, n_15881, n_15882, n_15883, n_15884, n_15885, n_15886,
       n_15887;
  wire n_15888, n_15889, n_15890, n_15891, n_15892, n_15893, n_15894,
       n_15895;
  wire n_15896, n_15897, n_15898, n_15899, n_15900, n_15901, n_15902,
       n_15903;
  wire n_15904, n_15905, n_15906, n_15907, n_15908, n_15909, n_15910,
       n_15911;
  wire n_15912, n_15913, n_15914, n_15915, n_15916, n_15917, n_15918,
       n_15919;
  wire n_15920, n_15921, n_15922, n_15923, n_15924, n_15925, n_15926,
       n_15927;
  wire n_15928, n_15929, n_15930, n_15931, n_15932, n_15933, n_15934,
       n_15935;
  wire n_15936, n_15937, n_15938, n_15939, n_15940, n_15941, n_15942,
       n_15943;
  wire n_15944, n_15945, n_15946, n_15947, n_15948, n_15949, n_15950,
       n_15951;
  wire n_15952, n_15953, n_15954, n_15955, n_15956, n_15957, n_15958,
       n_15959;
  wire n_15960, n_15961, n_15962, n_15963, n_15964, n_15965, n_15966,
       n_15967;
  wire n_15968, n_15969, n_15970, n_15971, n_15972, n_15973, n_15974,
       n_15975;
  wire n_15976, n_15977, n_15978, n_15979, n_15980, n_15981, n_15982,
       n_15983;
  wire n_15984, n_15985, n_15986, n_15987, n_15988, n_15989, n_15990,
       n_15991;
  wire n_15992, n_15993, n_15994, n_15995, n_15996, n_15997, n_15998,
       n_15999;
  wire n_16000, n_16001, n_16002, n_16003, n_16004, n_16005, n_16006,
       n_16007;
  wire n_16008, n_16009, n_16010, n_16011, n_16012, n_16013, n_16014,
       n_16015;
  wire n_16016, n_16017, n_16018, n_16019, n_16020, n_16021, n_16022,
       n_16023;
  wire n_16024, n_16025, n_16026, n_16027, n_16028, n_16029, n_16030,
       n_16031;
  wire n_16032, n_16033, n_16034, n_16035, n_16036, n_16037, n_16038,
       n_16039;
  wire n_16040, n_16041, n_16042, n_16043, n_16044, n_16045, n_16046,
       n_16047;
  wire n_16048, n_16049, n_16050, n_16051, n_16052, n_16053, n_16054,
       n_16055;
  wire n_16056, n_16057, n_16058, n_16059, n_16060, n_16061, n_16062,
       n_16063;
  wire n_16064, n_16065, n_16066, n_16067, n_16068, n_16069, n_16070,
       n_16071;
  wire n_16072, n_16073, n_16074, n_16075, n_16076, n_16077, n_16078,
       n_16079;
  wire n_16080, n_16081, n_16082, n_16083, n_16084, n_16085, n_16086,
       n_16087;
  wire n_16088, n_16089, n_16090, n_16091, n_16093, n_16094, n_16095,
       n_16096;
  wire n_16097, n_16098, n_16099, n_16100, n_16101, n_16103, n_16104,
       n_16105;
  wire n_16106, n_16107, n_16108, n_16109, n_16110, n_16111, n_16112,
       n_16113;
  wire n_16114, n_16115, n_16116, n_16117, n_16118, n_16119, n_16120,
       n_16121;
  wire n_16122, n_16123, n_16124, n_16125, n_16126, n_16127, n_16128,
       n_16129;
  wire n_16130, n_16131, n_16132, n_16133, n_16134, n_16135, n_16136,
       n_16137;
  wire n_16138, n_16139, n_16140, n_16141, n_16142, n_16143, n_16144,
       n_16145;
  wire n_16146, n_16147, n_16148, n_16149, n_16150, n_16151, n_16152,
       n_16153;
  wire n_16154, n_16155, n_16156, n_16157, n_16158, n_16159, n_16160,
       n_16161;
  wire n_16162, n_16163, n_16164, n_16165, n_16166, n_16167, n_16168,
       n_16169;
  wire n_16170, n_16171, n_16172, n_16173, n_16174, n_16175, n_16176,
       n_16177;
  wire n_16178, n_16179, n_16180, n_16181, n_16182, n_16183, n_16184,
       n_16185;
  wire n_16186, n_16187, n_16188, n_16189, n_16190, n_16191, n_16192,
       n_16193;
  wire n_16194, n_16195, n_16196, n_16197, n_16198, n_16199, n_16200,
       n_16203;
  wire n_16204, n_16205, n_16206, n_16207, n_16208, n_16209, n_16210,
       n_16211;
  wire n_16212, n_16213, n_16214, n_16215, n_16216, n_16217, n_16218,
       n_16219;
  wire n_16220, n_16221, n_16222, n_16223, n_16224, n_16225, n_16226,
       n_16227;
  wire n_16228, n_16229, n_16230, n_16231, n_16232, n_16233, n_16234,
       n_16235;
  wire n_16236, n_16237, n_16238, n_16239, n_16240, n_16241, n_16242,
       n_16243;
  wire n_16244, n_16245, n_16246, n_16247, n_16248, n_16249, n_16250,
       n_16251;
  wire n_16252, n_16253, n_16254, n_16255, n_16256, n_16257, n_16258,
       n_16259;
  wire n_16260, n_16261, n_16262, n_16263, n_16264, n_16265, n_16266,
       n_16267;
  wire n_16268, n_16269, n_16270, n_16271, n_16272, n_16273, n_16274,
       n_16275;
  wire n_16276, n_16277, n_16278, n_16279, n_16280, n_16281, n_16282,
       n_16283;
  wire n_16284, n_16285, n_16286, n_16287, n_16288, n_16289, n_16290,
       n_16291;
  wire n_16292, n_16293, n_16294, n_16295, n_16296, n_16297, n_16298,
       n_16299;
  wire n_16300, n_16301, n_16302, n_16303, n_16304, n_16305, n_16306,
       n_16307;
  wire n_16308, n_16309, n_16310, n_16311, n_16312, n_16313, n_16314,
       n_16315;
  wire n_16316, n_16317, n_16318, n_16319, n_16320, n_16321, n_16322,
       n_16323;
  wire n_16324, n_16325, n_16326, n_16327, n_16328, n_16329, n_16330,
       n_16331;
  wire n_16332, n_16333, n_16334, n_16335, n_16336, n_16337, n_16338,
       n_16339;
  wire n_16340, n_16341, n_16342, n_16343, n_16344, n_16345, n_16346,
       n_16347;
  wire n_16348, n_16349, n_16350, n_16351, n_16352, n_16353, n_16354,
       n_16355;
  wire n_16356, n_16357, n_16358, n_16359, n_16360, n_16361, n_16362,
       n_16363;
  wire n_16364, n_16365, n_16366, n_16367, n_16368, n_16369, n_16370,
       n_16371;
  wire n_16372, n_16373, n_16374, n_16375, n_16376, n_16377, n_16378,
       n_16379;
  wire n_16380, n_16381, n_16382, n_16383, n_16384, n_16385, n_16386,
       n_16387;
  wire n_16388, n_16389, n_16390, n_16391, n_16392, n_16393, n_16394,
       n_16395;
  wire n_16396, n_16397, n_16398, n_16399, n_16400, n_16401, n_16402,
       n_16403;
  wire n_16404, n_16405, n_16406, n_16407, n_16408, n_16409, n_16410,
       n_16411;
  wire n_16412, n_16413, n_16414, n_16415, n_16416, n_16417, n_16418,
       n_16419;
  wire n_16420, n_16421, n_16422, n_16423, n_16424, n_16425, n_16426,
       n_16427;
  wire n_16428, n_16429, n_16430, n_16431, n_16432, n_16433, n_16434,
       n_16435;
  wire n_16436, n_16437, n_16438, n_16439, n_16440, n_16441, n_16442,
       n_16443;
  wire n_16444, n_16445, n_16446, n_16447, n_16448, n_16449, n_16450,
       n_16451;
  wire n_16452, n_16453, n_16454, n_16455, n_16456, n_16457, n_16458,
       n_16459;
  wire n_16460, n_16461, n_16462, n_16463, n_16464, n_16465, n_16466,
       n_16467;
  wire n_16468, n_16469, n_16470, n_16471, n_16472, n_16473, n_16474,
       n_16475;
  wire n_16476, n_16477, n_16478, n_16479, n_16480, n_16481, n_16482,
       n_16483;
  wire n_16484, n_16485, n_16486, n_16487, n_16488, n_16489, n_16490,
       n_16491;
  wire n_16492, n_16493, n_16494, n_16495, n_16496, n_16497, n_16498,
       n_16499;
  wire n_16500, n_16501, n_16502, n_16503, n_16504, n_16505, n_16506,
       n_16507;
  wire n_16508, n_16509, n_16510, n_16511, n_16512, n_16513, n_16514,
       n_16515;
  wire n_16516, n_16517, n_16518, n_16519, n_16520, n_16521, n_16522,
       n_16523;
  wire n_16524, n_16525, n_16526, n_16527, n_16528, n_16529, n_16530,
       n_16531;
  wire n_16532, n_16533, n_16534, n_16535, n_16536, n_16537, n_16538,
       n_16539;
  wire n_16540, n_16541, n_16542, n_16543, n_16544, n_16545, n_16546,
       n_16547;
  wire n_16548, n_16549, n_16550, n_16551, n_16552, n_16553, n_16554,
       n_16555;
  wire n_16556, n_16557, n_16558, n_16559, n_16560, n_16561, n_16562,
       n_16563;
  wire n_16564, n_16565, n_16566, n_16567, n_16568, n_16569, n_16570,
       n_16571;
  wire n_16572, n_16573, n_16574, n_16575, n_16576, n_16577, n_16578,
       n_16579;
  wire n_16580, n_16581, n_16582, n_16583, n_16584, n_16585, n_16586,
       n_16587;
  wire n_16588, n_16589, n_16590, n_16591, n_16592, n_16593, n_16594,
       n_16595;
  wire n_16596, n_16597, n_16598, n_16599, n_16600, n_16601, n_16602,
       n_16603;
  wire n_16606, n_16607, n_16608, n_16609, n_16610, n_16611, n_16612,
       n_16613;
  wire n_16614, n_16615, n_16617, n_16618, n_16619, n_16620, n_16624,
       n_16625;
  wire n_16629, n_16630, n_16631, n_16632, n_16639, n_16640, n_16641,
       n_16642;
  wire n_16643, n_16644, n_16645, n_16646, n_16653, n_16654, n_16655,
       n_16656;
  wire n_16657, n_16658, n_16665, n_16666, n_16667, n_16668, n_16669,
       n_16670;
  wire n_16678, n_16679, n_16680, n_16681, n_16682, n_16683, n_16684,
       n_16685;
  wire n_16692, n_16693, n_16694, n_16695, n_16696, n_16697, n_16704,
       n_16705;
  wire n_16707, n_16708, n_16709, n_16710, n_16711, n_16712, n_16719,
       n_16720;
  wire n_16721, n_16722, n_16723, n_16724, n_16731, n_16732, n_16733,
       n_16734;
  wire n_16735, n_16736, n_16743, n_16744, n_16746, n_16747, n_16748,
       n_16749;
  wire n_16750, n_16751, n_16758, n_16759, n_16760, n_16761, n_16762,
       n_16763;
  wire n_16770, n_16771, n_16772, n_16773, n_16775, n_16776, n_16777,
       n_16778;
  wire n_16785, n_16786, n_16787, n_16788, n_16789, n_16790, n_16797,
       n_16798;
  wire n_16799, n_16800, n_16801, n_16802, n_16809, n_16810, n_16812,
       n_16813;
  wire n_16814, n_16815, n_16816, n_16817, n_16818, n_16825, n_16826,
       n_16827;
  wire n_16828, n_16829, n_16830, n_16837, n_16838, n_16839, n_16840,
       n_16842;
  wire n_16843, n_16844, n_16845, n_16852, n_16853, n_16854, n_16855,
       n_16856;
  wire n_16857, n_16864, n_16865, n_16866, n_16867, n_16868, n_16869,
       n_16876;
  wire n_16877, n_16879, n_16880, n_16881, n_16882, n_16883, n_16884,
       n_16891;
  wire n_16892, n_16893, n_16894, n_16895, n_16896, n_16903, n_16904,
       n_16905;
  wire n_16906, n_16908, n_16909, n_16910, n_16911, n_16918, n_16919,
       n_16920;
  wire n_16921, n_16922, n_16923, n_16930, n_16931, n_16932, n_16933,
       n_16934;
  wire n_16935, n_16942, n_16943, n_16945, n_16946, n_16947, n_16948,
       n_16949;
  wire n_16950, n_16957, n_16958, n_16959, n_16960, n_16961, n_16962,
       n_16963;
  wire n_16971, n_16972, n_16973, n_16974, n_16975, n_16976, n_16978,
       n_16979;
  wire n_16980, n_16984, n_16985, n_16986, n_16987, n_16988, n_16989,
       n_16992;
  wire n_16993, n_16994, n_16995, n_16996, n_16997, n_17001, n_17002,
       n_17003;
  wire n_17004, n_17007, n_17008, n_17009, n_17010, n_17012, n_17013,
       n_17016;
  wire n_17017, n_17019, n_17020, n_17021, n_17022, n_17025, n_17026,
       n_17027;
  wire n_17028, n_17030, n_17032, n_17033, n_17034, n_17035, n_17038,
       n_17039;
  wire n_17041, n_17042, n_17044, n_17045, n_17046, n_17047, n_17050,
       n_17051;
  wire n_17053, n_17054, n_17055, n_17056, n_17057, n_17058, n_17062,
       n_17063;
  wire n_17065, n_17066, n_17068, n_17069, n_17071, n_17072, n_17074,
       n_17075;
  wire n_17077, n_17078, n_17080, n_17081, n_17083, n_17084, n_17086,
       n_17087;
  wire n_17089, n_17090, n_17092, n_17093, n_17095, n_17096, n_17098,
       n_17099;
  wire n_17101, n_17102, n_17104, n_17105, n_17107, n_17108, n_17110,
       n_17111;
  wire n_17113, n_17114, n_17116, n_17117, n_17118, n_17119, n_17120,
       n_17121;
  wire n_17122, n_17123, n_17124, n_17125, n_17126;
  or g1 (\asqrt[63] , \a[126] , \a[127] );
  and g2 (n194, \a[126] , \a[127] );
  and g3 (n195, \a[126] , \asqrt[63] );
  not g4 (n_6, \a[124] );
  not g5 (n_7, \a[125] );
  and g6 (n196, n_6, n_7);
  not g7 (n_8, n195);
  not g8 (n_9, n196);
  and g9 (n197, n_8, n_9);
  or g10 (\asqrt[62] , n194, n197);
  and g11 (n199, \a[124] , \asqrt[62] );
  not g12 (n_13, \a[122] );
  not g13 (n_14, \a[123] );
  and g14 (n200, n_13, n_14);
  and g15 (n201, n_6, n200);
  not g16 (n_15, n199);
  not g17 (n_16, n201);
  and g18 (n202, n_15, n_16);
  and g19 (n203, n_6, \asqrt[62] );
  not g20 (n_17, n203);
  and g21 (n204, \a[125] , n_17);
  and g22 (n205, n196, \asqrt[62] );
  not g23 (n_18, n204);
  not g24 (n_19, n205);
  and g25 (n206, n_18, n_19);
  not g26 (n_20, n202);
  and g27 (n207, n_20, n206);
  not g28 (n_21, \asqrt[63] );
  not g29 (n_22, n207);
  and g30 (n208, n_21, n_22);
  not g31 (n_23, n206);
  and g32 (n209, n202, n_23);
  and g33 (n210, \a[126] , n196);
  not g34 (n_24, \a[126] );
  and g35 (n211, n_24, n_9);
  not g36 (n_25, n211);
  and g37 (n212, \a[127] , n_25);
  not g38 (n_26, n210);
  and g39 (n213, n_26, n212);
  not g40 (n_27, n209);
  not g41 (n_28, n213);
  and g42 (n214, n_27, n_28);
  not g43 (n_29, n214);
  or g44 (\asqrt[61] , n208, n_29);
  and g45 (n216, \a[122] , \asqrt[61] );
  not g46 (n_33, \a[120] );
  not g47 (n_34, \a[121] );
  and g48 (n217, n_33, n_34);
  and g49 (n218, n_13, n217);
  not g50 (n_35, n216);
  not g51 (n_36, n218);
  and g52 (n219, n_35, n_36);
  not g53 (n_37, n219);
  and g54 (n220, \asqrt[62] , n_37);
  and g60 (n224, n200, \asqrt[61] );
  and g61 (n225, n_13, \asqrt[61] );
  not g62 (n_40, n225);
  and g63 (n226, \a[123] , n_40);
  not g64 (n_41, n224);
  not g65 (n_42, n226);
  and g66 (n227, n_41, n_42);
  not g67 (n_43, n223);
  and g68 (n228, n_43, n227);
  not g69 (n_44, n220);
  not g70 (n_45, n228);
  and g71 (n229, n_44, n_45);
  not g74 (n_46, n208);
  not g76 (n_47, n232);
  and g77 (n233, n_41, n_47);
  not g78 (n_48, n233);
  and g79 (n234, \a[124] , n_48);
  and g80 (n235, n_6, n_47);
  and g81 (n236, n_41, n235);
  not g82 (n_49, n234);
  not g83 (n_50, n236);
  and g84 (n237, n_49, n_50);
  and g85 (n238, n207, \asqrt[61] );
  not g88 (n_52, n237);
  not g90 (n_53, n229);
  not g92 (n_54, n241);
  and g93 (n242, n_21, n_54);
  and g94 (n243, n229, n237);
  and g95 (n244, n206, \asqrt[61] );
  not g96 (n_55, n244);
  and g97 (n245, n202, n_55);
  and g98 (n246, \asqrt[63] , n_22);
  not g99 (n_56, n245);
  and g100 (n247, n_56, n246);
  not g104 (n_57, n247);
  not g105 (n_58, n250);
  not g107 (n_59, n243);
  and g111 (n254, \a[120] , \asqrt[60] );
  not g112 (n_64, \a[118] );
  not g113 (n_65, \a[119] );
  and g114 (n255, n_64, n_65);
  and g115 (n256, n_33, n255);
  not g116 (n_66, n254);
  not g117 (n_67, n256);
  and g118 (n257, n_66, n_67);
  not g119 (n_68, n257);
  and g120 (n258, \asqrt[61] , n_68);
  and g121 (n259, n_33, \asqrt[60] );
  not g122 (n_69, n259);
  and g123 (n260, \a[121] , n_69);
  and g124 (n261, n217, \asqrt[60] );
  not g125 (n_70, n260);
  not g126 (n_71, n261);
  and g127 (n262, n_70, n_71);
  not g132 (n_72, n266);
  and g133 (n267, n262, n_72);
  not g134 (n_73, n258);
  not g135 (n_74, n267);
  and g136 (n268, n_73, n_74);
  not g137 (n_75, n268);
  and g138 (n269, \asqrt[62] , n_75);
  not g139 (n_76, \asqrt[62] );
  and g140 (n270, n_76, n_73);
  and g141 (n271, n_74, n270);
  not g145 (n_77, n242);
  not g147 (n_78, n275);
  and g148 (n276, n_71, n_78);
  not g149 (n_79, n276);
  and g150 (n277, \a[122] , n_79);
  and g151 (n278, n_13, n_78);
  and g152 (n279, n_71, n278);
  not g153 (n_80, n277);
  not g154 (n_81, n279);
  and g155 (n280, n_80, n_81);
  not g156 (n_82, n271);
  not g157 (n_83, n280);
  and g158 (n281, n_82, n_83);
  not g159 (n_84, n269);
  not g160 (n_85, n281);
  and g161 (n282, n_84, n_85);
  and g162 (n283, n_44, n_43);
  not g163 (n_86, n227);
  and g164 (n284, n_86, n283);
  and g165 (n285, \asqrt[60] , n284);
  and g166 (n286, \asqrt[60] , n283);
  not g167 (n_87, n286);
  and g168 (n287, n227, n_87);
  not g169 (n_88, n285);
  not g170 (n_89, n287);
  and g171 (n288, n_88, n_89);
  and g172 (n289, n_53, n_52);
  and g173 (n290, \asqrt[60] , n289);
  not g176 (n_91, n288);
  not g178 (n_92, n282);
  not g180 (n_93, n293);
  and g181 (n294, n_21, n_93);
  and g182 (n295, n_84, n288);
  and g183 (n296, n_85, n295);
  and g184 (n297, n229, \asqrt[60] );
  not g185 (n_94, n297);
  and g186 (n298, n_52, n_94);
  and g187 (n299, \asqrt[63] , n_59);
  not g188 (n_95, n298);
  and g189 (n300, n_95, n299);
  not g195 (n_96, n300);
  not g196 (n_97, n305);
  not g198 (n_98, n296);
  and g202 (n309, \a[118] , \asqrt[59] );
  not g203 (n_103, \a[116] );
  not g204 (n_104, \a[117] );
  and g205 (n310, n_103, n_104);
  and g206 (n311, n_64, n310);
  not g207 (n_105, n309);
  not g208 (n_106, n311);
  and g209 (n312, n_105, n_106);
  not g210 (n_107, n312);
  and g211 (n313, \asqrt[60] , n_107);
  and g217 (n319, n_64, \asqrt[59] );
  not g218 (n_108, n319);
  and g219 (n320, \a[119] , n_108);
  and g220 (n321, n255, \asqrt[59] );
  not g221 (n_109, n320);
  not g222 (n_110, n321);
  and g223 (n322, n_109, n_110);
  not g224 (n_111, n318);
  and g225 (n323, n_111, n322);
  not g226 (n_112, n313);
  not g227 (n_113, n323);
  and g228 (n324, n_112, n_113);
  not g229 (n_114, n324);
  and g230 (n325, \asqrt[61] , n_114);
  not g231 (n_115, \asqrt[61] );
  and g232 (n326, n_115, n_112);
  and g233 (n327, n_113, n326);
  not g237 (n_116, n294);
  not g239 (n_117, n331);
  and g240 (n332, n_110, n_117);
  not g241 (n_118, n332);
  and g242 (n333, \a[120] , n_118);
  and g243 (n334, n_33, n_117);
  and g244 (n335, n_110, n334);
  not g245 (n_119, n333);
  not g246 (n_120, n335);
  and g247 (n336, n_119, n_120);
  not g248 (n_121, n327);
  not g249 (n_122, n336);
  and g250 (n337, n_121, n_122);
  not g251 (n_123, n325);
  not g252 (n_124, n337);
  and g253 (n338, n_123, n_124);
  not g254 (n_125, n338);
  and g255 (n339, \asqrt[62] , n_125);
  and g256 (n340, n_76, n_123);
  and g257 (n341, n_124, n340);
  and g262 (n345, n_73, n_72);
  and g263 (n346, \asqrt[59] , n345);
  not g264 (n_127, n346);
  and g265 (n347, n262, n_127);
  not g266 (n_128, n344);
  not g267 (n_129, n347);
  and g268 (n348, n_128, n_129);
  not g269 (n_130, n341);
  not g270 (n_131, n348);
  and g271 (n349, n_130, n_131);
  not g272 (n_132, n339);
  not g273 (n_133, n349);
  and g274 (n350, n_132, n_133);
  and g278 (n354, n_84, n_82);
  and g279 (n355, \asqrt[59] , n354);
  not g280 (n_134, n355);
  and g281 (n356, n_83, n_134);
  not g282 (n_135, n353);
  not g283 (n_136, n356);
  and g284 (n357, n_135, n_136);
  and g285 (n358, n_92, n_91);
  and g286 (n359, \asqrt[59] , n358);
  not g289 (n_138, n357);
  not g291 (n_139, n350);
  not g293 (n_140, n362);
  and g294 (n363, n_21, n_140);
  and g295 (n364, n_132, n357);
  and g296 (n365, n_133, n364);
  and g297 (n366, n282, \asqrt[59] );
  not g298 (n_141, n366);
  and g299 (n367, n_91, n_141);
  and g300 (n368, \asqrt[63] , n_98);
  not g301 (n_142, n367);
  and g302 (n369, n_142, n368);
  not g308 (n_143, n369);
  not g309 (n_144, n374);
  not g311 (n_145, n365);
  and g315 (n378, \a[116] , \asqrt[58] );
  not g316 (n_150, \a[114] );
  not g317 (n_151, \a[115] );
  and g318 (n379, n_150, n_151);
  and g319 (n380, n_103, n379);
  not g320 (n_152, n378);
  not g321 (n_153, n380);
  and g322 (n381, n_152, n_153);
  not g323 (n_154, n381);
  and g324 (n382, \asqrt[59] , n_154);
  and g330 (n388, n_103, \asqrt[58] );
  not g331 (n_155, n388);
  and g332 (n389, \a[117] , n_155);
  and g333 (n390, n310, \asqrt[58] );
  not g334 (n_156, n389);
  not g335 (n_157, n390);
  and g336 (n391, n_156, n_157);
  not g337 (n_158, n387);
  and g338 (n392, n_158, n391);
  not g339 (n_159, n382);
  not g340 (n_160, n392);
  and g341 (n393, n_159, n_160);
  not g342 (n_161, n393);
  and g343 (n394, \asqrt[60] , n_161);
  not g344 (n_162, \asqrt[60] );
  and g345 (n395, n_162, n_159);
  and g346 (n396, n_160, n395);
  not g350 (n_163, n363);
  not g352 (n_164, n400);
  and g353 (n401, n_157, n_164);
  not g354 (n_165, n401);
  and g355 (n402, \a[118] , n_165);
  and g356 (n403, n_64, n_164);
  and g357 (n404, n_157, n403);
  not g358 (n_166, n402);
  not g359 (n_167, n404);
  and g360 (n405, n_166, n_167);
  not g361 (n_168, n396);
  not g362 (n_169, n405);
  and g363 (n406, n_168, n_169);
  not g364 (n_170, n394);
  not g365 (n_171, n406);
  and g366 (n407, n_170, n_171);
  not g367 (n_172, n407);
  and g368 (n408, \asqrt[61] , n_172);
  and g369 (n409, n_112, n_111);
  not g370 (n_173, n322);
  and g371 (n410, n_173, n409);
  and g372 (n411, \asqrt[58] , n410);
  and g373 (n412, \asqrt[58] , n409);
  not g374 (n_174, n412);
  and g375 (n413, n322, n_174);
  not g376 (n_175, n411);
  not g377 (n_176, n413);
  and g378 (n414, n_175, n_176);
  and g379 (n415, n_115, n_170);
  and g380 (n416, n_171, n415);
  not g381 (n_177, n414);
  not g382 (n_178, n416);
  and g383 (n417, n_177, n_178);
  not g384 (n_179, n408);
  not g385 (n_180, n417);
  and g386 (n418, n_179, n_180);
  not g387 (n_181, n418);
  and g388 (n419, \asqrt[62] , n_181);
  and g392 (n423, n_123, n_121);
  and g393 (n424, \asqrt[58] , n423);
  not g394 (n_182, n424);
  and g395 (n425, n_122, n_182);
  not g396 (n_183, n422);
  not g397 (n_184, n425);
  and g398 (n426, n_183, n_184);
  and g399 (n427, n_76, n_179);
  and g400 (n428, n_180, n427);
  not g401 (n_185, n426);
  not g402 (n_186, n428);
  and g403 (n429, n_185, n_186);
  not g404 (n_187, n419);
  not g405 (n_188, n429);
  and g406 (n430, n_187, n_188);
  and g410 (n434, n_132, n_130);
  and g411 (n435, \asqrt[58] , n434);
  not g412 (n_189, n435);
  and g413 (n436, n_131, n_189);
  not g414 (n_190, n433);
  not g415 (n_191, n436);
  and g416 (n437, n_190, n_191);
  and g417 (n438, n_139, n_138);
  and g418 (n439, \asqrt[58] , n438);
  not g421 (n_193, n437);
  not g423 (n_194, n430);
  not g425 (n_195, n442);
  and g426 (n443, n_21, n_195);
  and g427 (n444, n_187, n437);
  and g428 (n445, n_188, n444);
  and g429 (n446, n_138, \asqrt[58] );
  not g430 (n_196, n446);
  and g431 (n447, n350, n_196);
  not g432 (n_197, n438);
  and g433 (n448, \asqrt[63] , n_197);
  not g434 (n_198, n447);
  and g435 (n449, n_198, n448);
  not g441 (n_199, n449);
  not g442 (n_200, n454);
  not g444 (n_201, n445);
  and g448 (n458, \a[114] , \asqrt[57] );
  not g449 (n_206, \a[112] );
  not g450 (n_207, \a[113] );
  and g451 (n459, n_206, n_207);
  and g452 (n460, n_150, n459);
  not g453 (n_208, n458);
  not g454 (n_209, n460);
  and g455 (n461, n_208, n_209);
  not g456 (n_210, n461);
  and g457 (n462, \asqrt[58] , n_210);
  and g463 (n468, n_150, \asqrt[57] );
  not g464 (n_211, n468);
  and g465 (n469, \a[115] , n_211);
  and g466 (n470, n379, \asqrt[57] );
  not g467 (n_212, n469);
  not g468 (n_213, n470);
  and g469 (n471, n_212, n_213);
  not g470 (n_214, n467);
  and g471 (n472, n_214, n471);
  not g472 (n_215, n462);
  not g473 (n_216, n472);
  and g474 (n473, n_215, n_216);
  not g475 (n_217, n473);
  and g476 (n474, \asqrt[59] , n_217);
  not g477 (n_218, \asqrt[59] );
  and g478 (n475, n_218, n_215);
  and g479 (n476, n_216, n475);
  not g483 (n_219, n443);
  not g485 (n_220, n480);
  and g486 (n481, n_213, n_220);
  not g487 (n_221, n481);
  and g488 (n482, \a[116] , n_221);
  and g489 (n483, n_103, n_220);
  and g490 (n484, n_213, n483);
  not g491 (n_222, n482);
  not g492 (n_223, n484);
  and g493 (n485, n_222, n_223);
  not g494 (n_224, n476);
  not g495 (n_225, n485);
  and g496 (n486, n_224, n_225);
  not g497 (n_226, n474);
  not g498 (n_227, n486);
  and g499 (n487, n_226, n_227);
  not g500 (n_228, n487);
  and g501 (n488, \asqrt[60] , n_228);
  and g502 (n489, n_159, n_158);
  not g503 (n_229, n391);
  and g504 (n490, n_229, n489);
  and g505 (n491, \asqrt[57] , n490);
  and g506 (n492, \asqrt[57] , n489);
  not g507 (n_230, n492);
  and g508 (n493, n391, n_230);
  not g509 (n_231, n491);
  not g510 (n_232, n493);
  and g511 (n494, n_231, n_232);
  and g512 (n495, n_162, n_226);
  and g513 (n496, n_227, n495);
  not g514 (n_233, n494);
  not g515 (n_234, n496);
  and g516 (n497, n_233, n_234);
  not g517 (n_235, n488);
  not g518 (n_236, n497);
  and g519 (n498, n_235, n_236);
  not g520 (n_237, n498);
  and g521 (n499, \asqrt[61] , n_237);
  and g525 (n503, n_170, n_168);
  and g526 (n504, \asqrt[57] , n503);
  not g527 (n_238, n504);
  and g528 (n505, n_169, n_238);
  not g529 (n_239, n502);
  not g530 (n_240, n505);
  and g531 (n506, n_239, n_240);
  and g532 (n507, n_115, n_235);
  and g533 (n508, n_236, n507);
  not g534 (n_241, n506);
  not g535 (n_242, n508);
  and g536 (n509, n_241, n_242);
  not g537 (n_243, n499);
  not g538 (n_244, n509);
  and g539 (n510, n_243, n_244);
  not g540 (n_245, n510);
  and g541 (n511, \asqrt[62] , n_245);
  and g545 (n515, n_179, n_178);
  and g546 (n516, \asqrt[57] , n515);
  not g547 (n_246, n516);
  and g548 (n517, n_177, n_246);
  not g549 (n_247, n514);
  not g550 (n_248, n517);
  and g551 (n518, n_247, n_248);
  and g552 (n519, n_76, n_243);
  and g553 (n520, n_244, n519);
  not g554 (n_249, n518);
  not g555 (n_250, n520);
  and g556 (n521, n_249, n_250);
  not g557 (n_251, n511);
  not g558 (n_252, n521);
  and g559 (n522, n_251, n_252);
  and g563 (n526, n_187, n_186);
  and g564 (n527, \asqrt[57] , n526);
  not g565 (n_253, n527);
  and g566 (n528, n_185, n_253);
  not g567 (n_254, n525);
  not g568 (n_255, n528);
  and g569 (n529, n_254, n_255);
  and g570 (n530, n_194, n_193);
  and g571 (n531, \asqrt[57] , n530);
  not g574 (n_257, n529);
  not g576 (n_258, n522);
  not g578 (n_259, n534);
  and g579 (n535, n_21, n_259);
  and g580 (n536, n_251, n529);
  and g581 (n537, n_252, n536);
  and g582 (n538, n_193, \asqrt[57] );
  not g583 (n_260, n538);
  and g584 (n539, n430, n_260);
  not g585 (n_261, n530);
  and g586 (n540, \asqrt[63] , n_261);
  not g587 (n_262, n539);
  and g588 (n541, n_262, n540);
  not g594 (n_263, n541);
  not g595 (n_264, n546);
  not g597 (n_265, n537);
  and g601 (n550, \a[112] , \asqrt[56] );
  not g602 (n_270, \a[110] );
  not g603 (n_271, \a[111] );
  and g604 (n551, n_270, n_271);
  and g605 (n552, n_206, n551);
  not g606 (n_272, n550);
  not g607 (n_273, n552);
  and g608 (n553, n_272, n_273);
  not g609 (n_274, n553);
  and g610 (n554, \asqrt[57] , n_274);
  and g611 (n555, n_206, \asqrt[56] );
  not g612 (n_275, n555);
  and g613 (n556, \a[113] , n_275);
  and g614 (n557, n459, \asqrt[56] );
  not g615 (n_276, n556);
  not g616 (n_277, n557);
  and g617 (n558, n_276, n_277);
  not g623 (n_278, n563);
  and g624 (n564, n558, n_278);
  not g625 (n_279, n554);
  not g626 (n_280, n564);
  and g627 (n565, n_279, n_280);
  not g628 (n_281, n565);
  and g629 (n566, \asqrt[58] , n_281);
  not g630 (n_282, \asqrt[58] );
  and g631 (n567, n_282, n_279);
  and g632 (n568, n_280, n567);
  not g636 (n_283, n535);
  not g638 (n_284, n572);
  and g639 (n573, n_277, n_284);
  not g640 (n_285, n573);
  and g641 (n574, \a[114] , n_285);
  and g642 (n575, n_150, n_284);
  and g643 (n576, n_277, n575);
  not g644 (n_286, n574);
  not g645 (n_287, n576);
  and g646 (n577, n_286, n_287);
  not g647 (n_288, n568);
  not g648 (n_289, n577);
  and g649 (n578, n_288, n_289);
  not g650 (n_290, n566);
  not g651 (n_291, n578);
  and g652 (n579, n_290, n_291);
  not g653 (n_292, n579);
  and g654 (n580, \asqrt[59] , n_292);
  and g655 (n581, n_215, n_214);
  not g656 (n_293, n471);
  and g657 (n582, n_293, n581);
  and g658 (n583, \asqrt[56] , n582);
  and g659 (n584, \asqrt[56] , n581);
  not g660 (n_294, n584);
  and g661 (n585, n471, n_294);
  not g662 (n_295, n583);
  not g663 (n_296, n585);
  and g664 (n586, n_295, n_296);
  and g665 (n587, n_218, n_290);
  and g666 (n588, n_291, n587);
  not g667 (n_297, n586);
  not g668 (n_298, n588);
  and g669 (n589, n_297, n_298);
  not g670 (n_299, n580);
  not g671 (n_300, n589);
  and g672 (n590, n_299, n_300);
  not g673 (n_301, n590);
  and g674 (n591, \asqrt[60] , n_301);
  and g678 (n595, n_226, n_224);
  and g679 (n596, \asqrt[56] , n595);
  not g680 (n_302, n596);
  and g681 (n597, n_225, n_302);
  not g682 (n_303, n594);
  not g683 (n_304, n597);
  and g684 (n598, n_303, n_304);
  and g685 (n599, n_162, n_299);
  and g686 (n600, n_300, n599);
  not g687 (n_305, n598);
  not g688 (n_306, n600);
  and g689 (n601, n_305, n_306);
  not g690 (n_307, n591);
  not g691 (n_308, n601);
  and g692 (n602, n_307, n_308);
  not g693 (n_309, n602);
  and g694 (n603, \asqrt[61] , n_309);
  and g698 (n607, n_235, n_234);
  and g699 (n608, \asqrt[56] , n607);
  not g700 (n_310, n608);
  and g701 (n609, n_233, n_310);
  not g702 (n_311, n606);
  not g703 (n_312, n609);
  and g704 (n610, n_311, n_312);
  and g705 (n611, n_115, n_307);
  and g706 (n612, n_308, n611);
  not g707 (n_313, n610);
  not g708 (n_314, n612);
  and g709 (n613, n_313, n_314);
  not g710 (n_315, n603);
  not g711 (n_316, n613);
  and g712 (n614, n_315, n_316);
  not g713 (n_317, n614);
  and g714 (n615, \asqrt[62] , n_317);
  and g718 (n619, n_243, n_242);
  and g719 (n620, \asqrt[56] , n619);
  not g720 (n_318, n620);
  and g721 (n621, n_241, n_318);
  not g722 (n_319, n618);
  not g723 (n_320, n621);
  and g724 (n622, n_319, n_320);
  and g725 (n623, n_76, n_315);
  and g726 (n624, n_316, n623);
  not g727 (n_321, n622);
  not g728 (n_322, n624);
  and g729 (n625, n_321, n_322);
  not g730 (n_323, n615);
  not g731 (n_324, n625);
  and g732 (n626, n_323, n_324);
  and g736 (n630, n_251, n_250);
  and g737 (n631, \asqrt[56] , n630);
  not g738 (n_325, n631);
  and g739 (n632, n_249, n_325);
  not g740 (n_326, n629);
  not g741 (n_327, n632);
  and g742 (n633, n_326, n_327);
  and g743 (n634, n_258, n_257);
  and g744 (n635, \asqrt[56] , n634);
  not g747 (n_329, n633);
  not g749 (n_330, n626);
  not g751 (n_331, n638);
  and g752 (n639, n_21, n_331);
  and g753 (n640, n_323, n633);
  and g754 (n641, n_324, n640);
  and g755 (n642, n_257, \asqrt[56] );
  not g756 (n_332, n642);
  and g757 (n643, n522, n_332);
  not g758 (n_333, n634);
  and g759 (n644, \asqrt[63] , n_333);
  not g760 (n_334, n643);
  and g761 (n645, n_334, n644);
  not g767 (n_335, n645);
  not g768 (n_336, n650);
  not g770 (n_337, n641);
  and g774 (n654, \a[110] , \asqrt[55] );
  not g775 (n_342, \a[108] );
  not g776 (n_343, \a[109] );
  and g777 (n655, n_342, n_343);
  and g778 (n656, n_270, n655);
  not g779 (n_344, n654);
  not g780 (n_345, n656);
  and g781 (n657, n_344, n_345);
  not g782 (n_346, n657);
  and g783 (n658, \asqrt[56] , n_346);
  and g789 (n664, n_270, \asqrt[55] );
  not g790 (n_347, n664);
  and g791 (n665, \a[111] , n_347);
  and g792 (n666, n551, \asqrt[55] );
  not g793 (n_348, n665);
  not g794 (n_349, n666);
  and g795 (n667, n_348, n_349);
  not g796 (n_350, n663);
  and g797 (n668, n_350, n667);
  not g798 (n_351, n658);
  not g799 (n_352, n668);
  and g800 (n669, n_351, n_352);
  not g801 (n_353, n669);
  and g802 (n670, \asqrt[57] , n_353);
  not g803 (n_354, \asqrt[57] );
  and g804 (n671, n_354, n_351);
  and g805 (n672, n_352, n671);
  not g809 (n_355, n639);
  not g811 (n_356, n676);
  and g812 (n677, n_349, n_356);
  not g813 (n_357, n677);
  and g814 (n678, \a[112] , n_357);
  and g815 (n679, n_206, n_356);
  and g816 (n680, n_349, n679);
  not g817 (n_358, n678);
  not g818 (n_359, n680);
  and g819 (n681, n_358, n_359);
  not g820 (n_360, n672);
  not g821 (n_361, n681);
  and g822 (n682, n_360, n_361);
  not g823 (n_362, n670);
  not g824 (n_363, n682);
  and g825 (n683, n_362, n_363);
  not g826 (n_364, n683);
  and g827 (n684, \asqrt[58] , n_364);
  and g828 (n685, n_282, n_362);
  and g829 (n686, n_363, n685);
  and g834 (n690, n_279, n_278);
  and g835 (n691, \asqrt[55] , n690);
  not g836 (n_366, n691);
  and g837 (n692, n558, n_366);
  not g838 (n_367, n689);
  not g839 (n_368, n692);
  and g840 (n693, n_367, n_368);
  not g841 (n_369, n686);
  not g842 (n_370, n693);
  and g843 (n694, n_369, n_370);
  not g844 (n_371, n684);
  not g845 (n_372, n694);
  and g846 (n695, n_371, n_372);
  not g847 (n_373, n695);
  and g848 (n696, \asqrt[59] , n_373);
  and g852 (n700, n_290, n_288);
  and g853 (n701, \asqrt[55] , n700);
  not g854 (n_374, n701);
  and g855 (n702, n_289, n_374);
  not g856 (n_375, n699);
  not g857 (n_376, n702);
  and g858 (n703, n_375, n_376);
  and g859 (n704, n_218, n_371);
  and g860 (n705, n_372, n704);
  not g861 (n_377, n703);
  not g862 (n_378, n705);
  and g863 (n706, n_377, n_378);
  not g864 (n_379, n696);
  not g865 (n_380, n706);
  and g866 (n707, n_379, n_380);
  not g867 (n_381, n707);
  and g868 (n708, \asqrt[60] , n_381);
  and g872 (n712, n_299, n_298);
  and g873 (n713, \asqrt[55] , n712);
  not g874 (n_382, n713);
  and g875 (n714, n_297, n_382);
  not g876 (n_383, n711);
  not g877 (n_384, n714);
  and g878 (n715, n_383, n_384);
  and g879 (n716, n_162, n_379);
  and g880 (n717, n_380, n716);
  not g881 (n_385, n715);
  not g882 (n_386, n717);
  and g883 (n718, n_385, n_386);
  not g884 (n_387, n708);
  not g885 (n_388, n718);
  and g886 (n719, n_387, n_388);
  not g887 (n_389, n719);
  and g888 (n720, \asqrt[61] , n_389);
  and g892 (n724, n_307, n_306);
  and g893 (n725, \asqrt[55] , n724);
  not g894 (n_390, n725);
  and g895 (n726, n_305, n_390);
  not g896 (n_391, n723);
  not g897 (n_392, n726);
  and g898 (n727, n_391, n_392);
  and g899 (n728, n_115, n_387);
  and g900 (n729, n_388, n728);
  not g901 (n_393, n727);
  not g902 (n_394, n729);
  and g903 (n730, n_393, n_394);
  not g904 (n_395, n720);
  not g905 (n_396, n730);
  and g906 (n731, n_395, n_396);
  not g907 (n_397, n731);
  and g908 (n732, \asqrt[62] , n_397);
  and g912 (n736, n_315, n_314);
  and g913 (n737, \asqrt[55] , n736);
  not g914 (n_398, n737);
  and g915 (n738, n_313, n_398);
  not g916 (n_399, n735);
  not g917 (n_400, n738);
  and g918 (n739, n_399, n_400);
  and g919 (n740, n_76, n_395);
  and g920 (n741, n_396, n740);
  not g921 (n_401, n739);
  not g922 (n_402, n741);
  and g923 (n742, n_401, n_402);
  not g924 (n_403, n732);
  not g925 (n_404, n742);
  and g926 (n743, n_403, n_404);
  and g930 (n747, n_323, n_322);
  and g931 (n748, \asqrt[55] , n747);
  not g932 (n_405, n748);
  and g933 (n749, n_321, n_405);
  not g934 (n_406, n746);
  not g935 (n_407, n749);
  and g936 (n750, n_406, n_407);
  and g937 (n751, n_330, n_329);
  and g938 (n752, \asqrt[55] , n751);
  not g941 (n_409, n750);
  not g943 (n_410, n743);
  not g945 (n_411, n755);
  and g946 (n756, n_21, n_411);
  and g947 (n757, n_403, n750);
  and g948 (n758, n_404, n757);
  and g949 (n759, n_329, \asqrt[55] );
  not g950 (n_412, n759);
  and g951 (n760, n626, n_412);
  not g952 (n_413, n751);
  and g953 (n761, \asqrt[63] , n_413);
  not g954 (n_414, n760);
  and g955 (n762, n_414, n761);
  not g961 (n_415, n762);
  not g962 (n_416, n767);
  not g964 (n_417, n758);
  and g968 (n771, \a[108] , \asqrt[54] );
  not g969 (n_422, \a[106] );
  not g970 (n_423, \a[107] );
  and g971 (n772, n_422, n_423);
  and g972 (n773, n_342, n772);
  not g973 (n_424, n771);
  not g974 (n_425, n773);
  and g975 (n774, n_424, n_425);
  not g976 (n_426, n774);
  and g977 (n775, \asqrt[55] , n_426);
  and g983 (n781, n_342, \asqrt[54] );
  not g984 (n_427, n781);
  and g985 (n782, \a[109] , n_427);
  and g986 (n783, n655, \asqrt[54] );
  not g987 (n_428, n782);
  not g988 (n_429, n783);
  and g989 (n784, n_428, n_429);
  not g990 (n_430, n780);
  and g991 (n785, n_430, n784);
  not g992 (n_431, n775);
  not g993 (n_432, n785);
  and g994 (n786, n_431, n_432);
  not g995 (n_433, n786);
  and g996 (n787, \asqrt[56] , n_433);
  not g997 (n_434, \asqrt[56] );
  and g998 (n788, n_434, n_431);
  and g999 (n789, n_432, n788);
  not g1003 (n_435, n756);
  not g1005 (n_436, n793);
  and g1006 (n794, n_429, n_436);
  not g1007 (n_437, n794);
  and g1008 (n795, \a[110] , n_437);
  and g1009 (n796, n_270, n_436);
  and g1010 (n797, n_429, n796);
  not g1011 (n_438, n795);
  not g1012 (n_439, n797);
  and g1013 (n798, n_438, n_439);
  not g1014 (n_440, n789);
  not g1015 (n_441, n798);
  and g1016 (n799, n_440, n_441);
  not g1017 (n_442, n787);
  not g1018 (n_443, n799);
  and g1019 (n800, n_442, n_443);
  not g1020 (n_444, n800);
  and g1021 (n801, \asqrt[57] , n_444);
  and g1022 (n802, n_351, n_350);
  not g1023 (n_445, n667);
  and g1024 (n803, n_445, n802);
  and g1025 (n804, \asqrt[54] , n803);
  and g1026 (n805, \asqrt[54] , n802);
  not g1027 (n_446, n805);
  and g1028 (n806, n667, n_446);
  not g1029 (n_447, n804);
  not g1030 (n_448, n806);
  and g1031 (n807, n_447, n_448);
  and g1032 (n808, n_354, n_442);
  and g1033 (n809, n_443, n808);
  not g1034 (n_449, n807);
  not g1035 (n_450, n809);
  and g1036 (n810, n_449, n_450);
  not g1037 (n_451, n801);
  not g1038 (n_452, n810);
  and g1039 (n811, n_451, n_452);
  not g1040 (n_453, n811);
  and g1041 (n812, \asqrt[58] , n_453);
  and g1045 (n816, n_362, n_360);
  and g1046 (n817, \asqrt[54] , n816);
  not g1047 (n_454, n817);
  and g1048 (n818, n_361, n_454);
  not g1049 (n_455, n815);
  not g1050 (n_456, n818);
  and g1051 (n819, n_455, n_456);
  and g1052 (n820, n_282, n_451);
  and g1053 (n821, n_452, n820);
  not g1054 (n_457, n819);
  not g1055 (n_458, n821);
  and g1056 (n822, n_457, n_458);
  not g1057 (n_459, n812);
  not g1058 (n_460, n822);
  and g1059 (n823, n_459, n_460);
  not g1060 (n_461, n823);
  and g1061 (n824, \asqrt[59] , n_461);
  and g1062 (n825, n_218, n_459);
  and g1063 (n826, n_460, n825);
  and g1067 (n830, n_371, n_369);
  and g1068 (n831, \asqrt[54] , n830);
  not g1069 (n_462, n831);
  and g1070 (n832, n_370, n_462);
  not g1071 (n_463, n829);
  not g1072 (n_464, n832);
  and g1073 (n833, n_463, n_464);
  not g1074 (n_465, n826);
  not g1075 (n_466, n833);
  and g1076 (n834, n_465, n_466);
  not g1077 (n_467, n824);
  not g1078 (n_468, n834);
  and g1079 (n835, n_467, n_468);
  not g1080 (n_469, n835);
  and g1081 (n836, \asqrt[60] , n_469);
  and g1085 (n840, n_379, n_378);
  and g1086 (n841, \asqrt[54] , n840);
  not g1087 (n_470, n841);
  and g1088 (n842, n_377, n_470);
  not g1089 (n_471, n839);
  not g1090 (n_472, n842);
  and g1091 (n843, n_471, n_472);
  and g1092 (n844, n_162, n_467);
  and g1093 (n845, n_468, n844);
  not g1094 (n_473, n843);
  not g1095 (n_474, n845);
  and g1096 (n846, n_473, n_474);
  not g1097 (n_475, n836);
  not g1098 (n_476, n846);
  and g1099 (n847, n_475, n_476);
  not g1100 (n_477, n847);
  and g1101 (n848, \asqrt[61] , n_477);
  and g1105 (n852, n_387, n_386);
  and g1106 (n853, \asqrt[54] , n852);
  not g1107 (n_478, n853);
  and g1108 (n854, n_385, n_478);
  not g1109 (n_479, n851);
  not g1110 (n_480, n854);
  and g1111 (n855, n_479, n_480);
  and g1112 (n856, n_115, n_475);
  and g1113 (n857, n_476, n856);
  not g1114 (n_481, n855);
  not g1115 (n_482, n857);
  and g1116 (n858, n_481, n_482);
  not g1117 (n_483, n848);
  not g1118 (n_484, n858);
  and g1119 (n859, n_483, n_484);
  not g1120 (n_485, n859);
  and g1121 (n860, \asqrt[62] , n_485);
  and g1125 (n864, n_395, n_394);
  and g1126 (n865, \asqrt[54] , n864);
  not g1127 (n_486, n865);
  and g1128 (n866, n_393, n_486);
  not g1129 (n_487, n863);
  not g1130 (n_488, n866);
  and g1131 (n867, n_487, n_488);
  and g1132 (n868, n_76, n_483);
  and g1133 (n869, n_484, n868);
  not g1134 (n_489, n867);
  not g1135 (n_490, n869);
  and g1136 (n870, n_489, n_490);
  not g1137 (n_491, n860);
  not g1138 (n_492, n870);
  and g1139 (n871, n_491, n_492);
  and g1143 (n875, n_403, n_402);
  and g1144 (n876, \asqrt[54] , n875);
  not g1145 (n_493, n876);
  and g1146 (n877, n_401, n_493);
  not g1147 (n_494, n874);
  not g1148 (n_495, n877);
  and g1149 (n878, n_494, n_495);
  and g1150 (n879, n_410, n_409);
  and g1151 (n880, \asqrt[54] , n879);
  not g1154 (n_497, n878);
  not g1156 (n_498, n871);
  not g1158 (n_499, n883);
  and g1159 (n884, n_21, n_499);
  and g1160 (n885, n_491, n878);
  and g1161 (n886, n_492, n885);
  and g1162 (n887, n_409, \asqrt[54] );
  not g1163 (n_500, n887);
  and g1164 (n888, n743, n_500);
  not g1165 (n_501, n879);
  and g1166 (n889, \asqrt[63] , n_501);
  not g1167 (n_502, n888);
  and g1168 (n890, n_502, n889);
  not g1174 (n_503, n890);
  not g1175 (n_504, n895);
  not g1177 (n_505, n886);
  and g1181 (n899, \a[106] , \asqrt[53] );
  not g1182 (n_510, \a[104] );
  not g1183 (n_511, \a[105] );
  and g1184 (n900, n_510, n_511);
  and g1185 (n901, n_422, n900);
  not g1186 (n_512, n899);
  not g1187 (n_513, n901);
  and g1188 (n902, n_512, n_513);
  not g1189 (n_514, n902);
  and g1190 (n903, \asqrt[54] , n_514);
  and g1196 (n909, n_422, \asqrt[53] );
  not g1197 (n_515, n909);
  and g1198 (n910, \a[107] , n_515);
  and g1199 (n911, n772, \asqrt[53] );
  not g1200 (n_516, n910);
  not g1201 (n_517, n911);
  and g1202 (n912, n_516, n_517);
  not g1203 (n_518, n908);
  and g1204 (n913, n_518, n912);
  not g1205 (n_519, n903);
  not g1206 (n_520, n913);
  and g1207 (n914, n_519, n_520);
  not g1208 (n_521, n914);
  and g1209 (n915, \asqrt[55] , n_521);
  not g1210 (n_522, \asqrt[55] );
  and g1211 (n916, n_522, n_519);
  and g1212 (n917, n_520, n916);
  not g1216 (n_523, n884);
  not g1218 (n_524, n921);
  and g1219 (n922, n_517, n_524);
  not g1220 (n_525, n922);
  and g1221 (n923, \a[108] , n_525);
  and g1222 (n924, n_342, n_524);
  and g1223 (n925, n_517, n924);
  not g1224 (n_526, n923);
  not g1225 (n_527, n925);
  and g1226 (n926, n_526, n_527);
  not g1227 (n_528, n917);
  not g1228 (n_529, n926);
  and g1229 (n927, n_528, n_529);
  not g1230 (n_530, n915);
  not g1231 (n_531, n927);
  and g1232 (n928, n_530, n_531);
  not g1233 (n_532, n928);
  and g1234 (n929, \asqrt[56] , n_532);
  and g1235 (n930, n_431, n_430);
  not g1236 (n_533, n784);
  and g1237 (n931, n_533, n930);
  and g1238 (n932, \asqrt[53] , n931);
  and g1239 (n933, \asqrt[53] , n930);
  not g1240 (n_534, n933);
  and g1241 (n934, n784, n_534);
  not g1242 (n_535, n932);
  not g1243 (n_536, n934);
  and g1244 (n935, n_535, n_536);
  and g1245 (n936, n_434, n_530);
  and g1246 (n937, n_531, n936);
  not g1247 (n_537, n935);
  not g1248 (n_538, n937);
  and g1249 (n938, n_537, n_538);
  not g1250 (n_539, n929);
  not g1251 (n_540, n938);
  and g1252 (n939, n_539, n_540);
  not g1253 (n_541, n939);
  and g1254 (n940, \asqrt[57] , n_541);
  and g1258 (n944, n_442, n_440);
  and g1259 (n945, \asqrt[53] , n944);
  not g1260 (n_542, n945);
  and g1261 (n946, n_441, n_542);
  not g1262 (n_543, n943);
  not g1263 (n_544, n946);
  and g1264 (n947, n_543, n_544);
  and g1265 (n948, n_354, n_539);
  and g1266 (n949, n_540, n948);
  not g1267 (n_545, n947);
  not g1268 (n_546, n949);
  and g1269 (n950, n_545, n_546);
  not g1270 (n_547, n940);
  not g1271 (n_548, n950);
  and g1272 (n951, n_547, n_548);
  not g1273 (n_549, n951);
  and g1274 (n952, \asqrt[58] , n_549);
  and g1278 (n956, n_451, n_450);
  and g1279 (n957, \asqrt[53] , n956);
  not g1280 (n_550, n957);
  and g1281 (n958, n_449, n_550);
  not g1282 (n_551, n955);
  not g1283 (n_552, n958);
  and g1284 (n959, n_551, n_552);
  and g1285 (n960, n_282, n_547);
  and g1286 (n961, n_548, n960);
  not g1287 (n_553, n959);
  not g1288 (n_554, n961);
  and g1289 (n962, n_553, n_554);
  not g1290 (n_555, n952);
  not g1291 (n_556, n962);
  and g1292 (n963, n_555, n_556);
  not g1293 (n_557, n963);
  and g1294 (n964, \asqrt[59] , n_557);
  and g1298 (n968, n_459, n_458);
  and g1299 (n969, \asqrt[53] , n968);
  not g1300 (n_558, n969);
  and g1301 (n970, n_457, n_558);
  not g1302 (n_559, n967);
  not g1303 (n_560, n970);
  and g1304 (n971, n_559, n_560);
  and g1305 (n972, n_218, n_555);
  and g1306 (n973, n_556, n972);
  not g1307 (n_561, n971);
  not g1308 (n_562, n973);
  and g1309 (n974, n_561, n_562);
  not g1310 (n_563, n964);
  not g1311 (n_564, n974);
  and g1312 (n975, n_563, n_564);
  not g1313 (n_565, n975);
  and g1314 (n976, \asqrt[60] , n_565);
  and g1315 (n977, n_162, n_563);
  and g1316 (n978, n_564, n977);
  and g1320 (n982, n_467, n_465);
  and g1321 (n983, \asqrt[53] , n982);
  not g1322 (n_566, n983);
  and g1323 (n984, n_466, n_566);
  not g1324 (n_567, n981);
  not g1325 (n_568, n984);
  and g1326 (n985, n_567, n_568);
  not g1327 (n_569, n978);
  not g1328 (n_570, n985);
  and g1329 (n986, n_569, n_570);
  not g1330 (n_571, n976);
  not g1331 (n_572, n986);
  and g1332 (n987, n_571, n_572);
  not g1333 (n_573, n987);
  and g1334 (n988, \asqrt[61] , n_573);
  and g1338 (n992, n_475, n_474);
  and g1339 (n993, \asqrt[53] , n992);
  not g1340 (n_574, n993);
  and g1341 (n994, n_473, n_574);
  not g1342 (n_575, n991);
  not g1343 (n_576, n994);
  and g1344 (n995, n_575, n_576);
  and g1345 (n996, n_115, n_571);
  and g1346 (n997, n_572, n996);
  not g1347 (n_577, n995);
  not g1348 (n_578, n997);
  and g1349 (n998, n_577, n_578);
  not g1350 (n_579, n988);
  not g1351 (n_580, n998);
  and g1352 (n999, n_579, n_580);
  not g1353 (n_581, n999);
  and g1354 (n1000, \asqrt[62] , n_581);
  and g1358 (n1004, n_483, n_482);
  and g1359 (n1005, \asqrt[53] , n1004);
  not g1360 (n_582, n1005);
  and g1361 (n1006, n_481, n_582);
  not g1362 (n_583, n1003);
  not g1363 (n_584, n1006);
  and g1364 (n1007, n_583, n_584);
  and g1365 (n1008, n_76, n_579);
  and g1366 (n1009, n_580, n1008);
  not g1367 (n_585, n1007);
  not g1368 (n_586, n1009);
  and g1369 (n1010, n_585, n_586);
  not g1370 (n_587, n1000);
  not g1371 (n_588, n1010);
  and g1372 (n1011, n_587, n_588);
  and g1376 (n1015, n_491, n_490);
  and g1377 (n1016, \asqrt[53] , n1015);
  not g1378 (n_589, n1016);
  and g1379 (n1017, n_489, n_589);
  not g1380 (n_590, n1014);
  not g1381 (n_591, n1017);
  and g1382 (n1018, n_590, n_591);
  and g1383 (n1019, n_498, n_497);
  and g1384 (n1020, \asqrt[53] , n1019);
  not g1387 (n_593, n1018);
  not g1389 (n_594, n1011);
  not g1391 (n_595, n1023);
  and g1392 (n1024, n_21, n_595);
  and g1393 (n1025, n_587, n1018);
  and g1394 (n1026, n_588, n1025);
  and g1395 (n1027, n_497, \asqrt[53] );
  not g1396 (n_596, n1027);
  and g1397 (n1028, n871, n_596);
  not g1398 (n_597, n1019);
  and g1399 (n1029, \asqrt[63] , n_597);
  not g1400 (n_598, n1028);
  and g1401 (n1030, n_598, n1029);
  not g1407 (n_599, n1030);
  not g1408 (n_600, n1035);
  not g1410 (n_601, n1026);
  and g1414 (n1039, \a[104] , \asqrt[52] );
  not g1415 (n_606, \a[102] );
  not g1416 (n_607, \a[103] );
  and g1417 (n1040, n_606, n_607);
  and g1418 (n1041, n_510, n1040);
  not g1419 (n_608, n1039);
  not g1420 (n_609, n1041);
  and g1421 (n1042, n_608, n_609);
  not g1422 (n_610, n1042);
  and g1423 (n1043, \asqrt[53] , n_610);
  and g1429 (n1049, n_510, \asqrt[52] );
  not g1430 (n_611, n1049);
  and g1431 (n1050, \a[105] , n_611);
  and g1432 (n1051, n900, \asqrt[52] );
  not g1433 (n_612, n1050);
  not g1434 (n_613, n1051);
  and g1435 (n1052, n_612, n_613);
  not g1436 (n_614, n1048);
  and g1437 (n1053, n_614, n1052);
  not g1438 (n_615, n1043);
  not g1439 (n_616, n1053);
  and g1440 (n1054, n_615, n_616);
  not g1441 (n_617, n1054);
  and g1442 (n1055, \asqrt[54] , n_617);
  not g1443 (n_618, \asqrt[54] );
  and g1444 (n1056, n_618, n_615);
  and g1445 (n1057, n_616, n1056);
  not g1449 (n_619, n1024);
  not g1451 (n_620, n1061);
  and g1452 (n1062, n_613, n_620);
  not g1453 (n_621, n1062);
  and g1454 (n1063, \a[106] , n_621);
  and g1455 (n1064, n_422, n_620);
  and g1456 (n1065, n_613, n1064);
  not g1457 (n_622, n1063);
  not g1458 (n_623, n1065);
  and g1459 (n1066, n_622, n_623);
  not g1460 (n_624, n1057);
  not g1461 (n_625, n1066);
  and g1462 (n1067, n_624, n_625);
  not g1463 (n_626, n1055);
  not g1464 (n_627, n1067);
  and g1465 (n1068, n_626, n_627);
  not g1466 (n_628, n1068);
  and g1467 (n1069, \asqrt[55] , n_628);
  and g1468 (n1070, n_519, n_518);
  not g1469 (n_629, n912);
  and g1470 (n1071, n_629, n1070);
  and g1471 (n1072, \asqrt[52] , n1071);
  and g1472 (n1073, \asqrt[52] , n1070);
  not g1473 (n_630, n1073);
  and g1474 (n1074, n912, n_630);
  not g1475 (n_631, n1072);
  not g1476 (n_632, n1074);
  and g1477 (n1075, n_631, n_632);
  and g1478 (n1076, n_522, n_626);
  and g1479 (n1077, n_627, n1076);
  not g1480 (n_633, n1075);
  not g1481 (n_634, n1077);
  and g1482 (n1078, n_633, n_634);
  not g1483 (n_635, n1069);
  not g1484 (n_636, n1078);
  and g1485 (n1079, n_635, n_636);
  not g1486 (n_637, n1079);
  and g1487 (n1080, \asqrt[56] , n_637);
  and g1491 (n1084, n_530, n_528);
  and g1492 (n1085, \asqrt[52] , n1084);
  not g1493 (n_638, n1085);
  and g1494 (n1086, n_529, n_638);
  not g1495 (n_639, n1083);
  not g1496 (n_640, n1086);
  and g1497 (n1087, n_639, n_640);
  and g1498 (n1088, n_434, n_635);
  and g1499 (n1089, n_636, n1088);
  not g1500 (n_641, n1087);
  not g1501 (n_642, n1089);
  and g1502 (n1090, n_641, n_642);
  not g1503 (n_643, n1080);
  not g1504 (n_644, n1090);
  and g1505 (n1091, n_643, n_644);
  not g1506 (n_645, n1091);
  and g1507 (n1092, \asqrt[57] , n_645);
  and g1511 (n1096, n_539, n_538);
  and g1512 (n1097, \asqrt[52] , n1096);
  not g1513 (n_646, n1097);
  and g1514 (n1098, n_537, n_646);
  not g1515 (n_647, n1095);
  not g1516 (n_648, n1098);
  and g1517 (n1099, n_647, n_648);
  and g1518 (n1100, n_354, n_643);
  and g1519 (n1101, n_644, n1100);
  not g1520 (n_649, n1099);
  not g1521 (n_650, n1101);
  and g1522 (n1102, n_649, n_650);
  not g1523 (n_651, n1092);
  not g1524 (n_652, n1102);
  and g1525 (n1103, n_651, n_652);
  not g1526 (n_653, n1103);
  and g1527 (n1104, \asqrt[58] , n_653);
  and g1531 (n1108, n_547, n_546);
  and g1532 (n1109, \asqrt[52] , n1108);
  not g1533 (n_654, n1109);
  and g1534 (n1110, n_545, n_654);
  not g1535 (n_655, n1107);
  not g1536 (n_656, n1110);
  and g1537 (n1111, n_655, n_656);
  and g1538 (n1112, n_282, n_651);
  and g1539 (n1113, n_652, n1112);
  not g1540 (n_657, n1111);
  not g1541 (n_658, n1113);
  and g1542 (n1114, n_657, n_658);
  not g1543 (n_659, n1104);
  not g1544 (n_660, n1114);
  and g1545 (n1115, n_659, n_660);
  not g1546 (n_661, n1115);
  and g1547 (n1116, \asqrt[59] , n_661);
  and g1551 (n1120, n_555, n_554);
  and g1552 (n1121, \asqrt[52] , n1120);
  not g1553 (n_662, n1121);
  and g1554 (n1122, n_553, n_662);
  not g1555 (n_663, n1119);
  not g1556 (n_664, n1122);
  and g1557 (n1123, n_663, n_664);
  and g1558 (n1124, n_218, n_659);
  and g1559 (n1125, n_660, n1124);
  not g1560 (n_665, n1123);
  not g1561 (n_666, n1125);
  and g1562 (n1126, n_665, n_666);
  not g1563 (n_667, n1116);
  not g1564 (n_668, n1126);
  and g1565 (n1127, n_667, n_668);
  not g1566 (n_669, n1127);
  and g1567 (n1128, \asqrt[60] , n_669);
  and g1571 (n1132, n_563, n_562);
  and g1572 (n1133, \asqrt[52] , n1132);
  not g1573 (n_670, n1133);
  and g1574 (n1134, n_561, n_670);
  not g1575 (n_671, n1131);
  not g1576 (n_672, n1134);
  and g1577 (n1135, n_671, n_672);
  and g1578 (n1136, n_162, n_667);
  and g1579 (n1137, n_668, n1136);
  not g1580 (n_673, n1135);
  not g1581 (n_674, n1137);
  and g1582 (n1138, n_673, n_674);
  not g1583 (n_675, n1128);
  not g1584 (n_676, n1138);
  and g1585 (n1139, n_675, n_676);
  not g1586 (n_677, n1139);
  and g1587 (n1140, \asqrt[61] , n_677);
  and g1588 (n1141, n_115, n_675);
  and g1589 (n1142, n_676, n1141);
  and g1593 (n1146, n_571, n_569);
  and g1594 (n1147, \asqrt[52] , n1146);
  not g1595 (n_678, n1147);
  and g1596 (n1148, n_570, n_678);
  not g1597 (n_679, n1145);
  not g1598 (n_680, n1148);
  and g1599 (n1149, n_679, n_680);
  not g1600 (n_681, n1142);
  not g1601 (n_682, n1149);
  and g1602 (n1150, n_681, n_682);
  not g1603 (n_683, n1140);
  not g1604 (n_684, n1150);
  and g1605 (n1151, n_683, n_684);
  not g1606 (n_685, n1151);
  and g1607 (n1152, \asqrt[62] , n_685);
  and g1611 (n1156, n_579, n_578);
  and g1612 (n1157, \asqrt[52] , n1156);
  not g1613 (n_686, n1157);
  and g1614 (n1158, n_577, n_686);
  not g1615 (n_687, n1155);
  not g1616 (n_688, n1158);
  and g1617 (n1159, n_687, n_688);
  and g1618 (n1160, n_76, n_683);
  and g1619 (n1161, n_684, n1160);
  not g1620 (n_689, n1159);
  not g1621 (n_690, n1161);
  and g1622 (n1162, n_689, n_690);
  not g1623 (n_691, n1152);
  not g1624 (n_692, n1162);
  and g1625 (n1163, n_691, n_692);
  and g1629 (n1167, n_587, n_586);
  and g1630 (n1168, \asqrt[52] , n1167);
  not g1631 (n_693, n1168);
  and g1632 (n1169, n_585, n_693);
  not g1633 (n_694, n1166);
  not g1634 (n_695, n1169);
  and g1635 (n1170, n_694, n_695);
  and g1636 (n1171, n_594, n_593);
  and g1637 (n1172, \asqrt[52] , n1171);
  not g1640 (n_697, n1170);
  not g1642 (n_698, n1163);
  not g1644 (n_699, n1175);
  and g1645 (n1176, n_21, n_699);
  and g1646 (n1177, n_691, n1170);
  and g1647 (n1178, n_692, n1177);
  and g1648 (n1179, n_593, \asqrt[52] );
  not g1649 (n_700, n1179);
  and g1650 (n1180, n1011, n_700);
  not g1651 (n_701, n1171);
  and g1652 (n1181, \asqrt[63] , n_701);
  not g1653 (n_702, n1180);
  and g1654 (n1182, n_702, n1181);
  not g1660 (n_703, n1182);
  not g1661 (n_704, n1187);
  not g1663 (n_705, n1178);
  and g1667 (n1191, \a[102] , \asqrt[51] );
  not g1668 (n_710, \a[100] );
  not g1669 (n_711, \a[101] );
  and g1670 (n1192, n_710, n_711);
  and g1671 (n1193, n_606, n1192);
  not g1672 (n_712, n1191);
  not g1673 (n_713, n1193);
  and g1674 (n1194, n_712, n_713);
  not g1675 (n_714, n1194);
  and g1676 (n1195, \asqrt[52] , n_714);
  and g1682 (n1201, n_606, \asqrt[51] );
  not g1683 (n_715, n1201);
  and g1684 (n1202, \a[103] , n_715);
  and g1685 (n1203, n1040, \asqrt[51] );
  not g1686 (n_716, n1202);
  not g1687 (n_717, n1203);
  and g1688 (n1204, n_716, n_717);
  not g1689 (n_718, n1200);
  and g1690 (n1205, n_718, n1204);
  not g1691 (n_719, n1195);
  not g1692 (n_720, n1205);
  and g1693 (n1206, n_719, n_720);
  not g1694 (n_721, n1206);
  and g1695 (n1207, \asqrt[53] , n_721);
  not g1696 (n_722, \asqrt[53] );
  and g1697 (n1208, n_722, n_719);
  and g1698 (n1209, n_720, n1208);
  not g1702 (n_723, n1176);
  not g1704 (n_724, n1213);
  and g1705 (n1214, n_717, n_724);
  not g1706 (n_725, n1214);
  and g1707 (n1215, \a[104] , n_725);
  and g1708 (n1216, n_510, n_724);
  and g1709 (n1217, n_717, n1216);
  not g1710 (n_726, n1215);
  not g1711 (n_727, n1217);
  and g1712 (n1218, n_726, n_727);
  not g1713 (n_728, n1209);
  not g1714 (n_729, n1218);
  and g1715 (n1219, n_728, n_729);
  not g1716 (n_730, n1207);
  not g1717 (n_731, n1219);
  and g1718 (n1220, n_730, n_731);
  not g1719 (n_732, n1220);
  and g1720 (n1221, \asqrt[54] , n_732);
  and g1721 (n1222, n_615, n_614);
  not g1722 (n_733, n1052);
  and g1723 (n1223, n_733, n1222);
  and g1724 (n1224, \asqrt[51] , n1223);
  and g1725 (n1225, \asqrt[51] , n1222);
  not g1726 (n_734, n1225);
  and g1727 (n1226, n1052, n_734);
  not g1728 (n_735, n1224);
  not g1729 (n_736, n1226);
  and g1730 (n1227, n_735, n_736);
  and g1731 (n1228, n_618, n_730);
  and g1732 (n1229, n_731, n1228);
  not g1733 (n_737, n1227);
  not g1734 (n_738, n1229);
  and g1735 (n1230, n_737, n_738);
  not g1736 (n_739, n1221);
  not g1737 (n_740, n1230);
  and g1738 (n1231, n_739, n_740);
  not g1739 (n_741, n1231);
  and g1740 (n1232, \asqrt[55] , n_741);
  and g1744 (n1236, n_626, n_624);
  and g1745 (n1237, \asqrt[51] , n1236);
  not g1746 (n_742, n1237);
  and g1747 (n1238, n_625, n_742);
  not g1748 (n_743, n1235);
  not g1749 (n_744, n1238);
  and g1750 (n1239, n_743, n_744);
  and g1751 (n1240, n_522, n_739);
  and g1752 (n1241, n_740, n1240);
  not g1753 (n_745, n1239);
  not g1754 (n_746, n1241);
  and g1755 (n1242, n_745, n_746);
  not g1756 (n_747, n1232);
  not g1757 (n_748, n1242);
  and g1758 (n1243, n_747, n_748);
  not g1759 (n_749, n1243);
  and g1760 (n1244, \asqrt[56] , n_749);
  and g1764 (n1248, n_635, n_634);
  and g1765 (n1249, \asqrt[51] , n1248);
  not g1766 (n_750, n1249);
  and g1767 (n1250, n_633, n_750);
  not g1768 (n_751, n1247);
  not g1769 (n_752, n1250);
  and g1770 (n1251, n_751, n_752);
  and g1771 (n1252, n_434, n_747);
  and g1772 (n1253, n_748, n1252);
  not g1773 (n_753, n1251);
  not g1774 (n_754, n1253);
  and g1775 (n1254, n_753, n_754);
  not g1776 (n_755, n1244);
  not g1777 (n_756, n1254);
  and g1778 (n1255, n_755, n_756);
  not g1779 (n_757, n1255);
  and g1780 (n1256, \asqrt[57] , n_757);
  and g1784 (n1260, n_643, n_642);
  and g1785 (n1261, \asqrt[51] , n1260);
  not g1786 (n_758, n1261);
  and g1787 (n1262, n_641, n_758);
  not g1788 (n_759, n1259);
  not g1789 (n_760, n1262);
  and g1790 (n1263, n_759, n_760);
  and g1791 (n1264, n_354, n_755);
  and g1792 (n1265, n_756, n1264);
  not g1793 (n_761, n1263);
  not g1794 (n_762, n1265);
  and g1795 (n1266, n_761, n_762);
  not g1796 (n_763, n1256);
  not g1797 (n_764, n1266);
  and g1798 (n1267, n_763, n_764);
  not g1799 (n_765, n1267);
  and g1800 (n1268, \asqrt[58] , n_765);
  and g1804 (n1272, n_651, n_650);
  and g1805 (n1273, \asqrt[51] , n1272);
  not g1806 (n_766, n1273);
  and g1807 (n1274, n_649, n_766);
  not g1808 (n_767, n1271);
  not g1809 (n_768, n1274);
  and g1810 (n1275, n_767, n_768);
  and g1811 (n1276, n_282, n_763);
  and g1812 (n1277, n_764, n1276);
  not g1813 (n_769, n1275);
  not g1814 (n_770, n1277);
  and g1815 (n1278, n_769, n_770);
  not g1816 (n_771, n1268);
  not g1817 (n_772, n1278);
  and g1818 (n1279, n_771, n_772);
  not g1819 (n_773, n1279);
  and g1820 (n1280, \asqrt[59] , n_773);
  and g1824 (n1284, n_659, n_658);
  and g1825 (n1285, \asqrt[51] , n1284);
  not g1826 (n_774, n1285);
  and g1827 (n1286, n_657, n_774);
  not g1828 (n_775, n1283);
  not g1829 (n_776, n1286);
  and g1830 (n1287, n_775, n_776);
  and g1831 (n1288, n_218, n_771);
  and g1832 (n1289, n_772, n1288);
  not g1833 (n_777, n1287);
  not g1834 (n_778, n1289);
  and g1835 (n1290, n_777, n_778);
  not g1836 (n_779, n1280);
  not g1837 (n_780, n1290);
  and g1838 (n1291, n_779, n_780);
  not g1839 (n_781, n1291);
  and g1840 (n1292, \asqrt[60] , n_781);
  and g1844 (n1296, n_667, n_666);
  and g1845 (n1297, \asqrt[51] , n1296);
  not g1846 (n_782, n1297);
  and g1847 (n1298, n_665, n_782);
  not g1848 (n_783, n1295);
  not g1849 (n_784, n1298);
  and g1850 (n1299, n_783, n_784);
  and g1851 (n1300, n_162, n_779);
  and g1852 (n1301, n_780, n1300);
  not g1853 (n_785, n1299);
  not g1854 (n_786, n1301);
  and g1855 (n1302, n_785, n_786);
  not g1856 (n_787, n1292);
  not g1857 (n_788, n1302);
  and g1858 (n1303, n_787, n_788);
  not g1859 (n_789, n1303);
  and g1860 (n1304, \asqrt[61] , n_789);
  and g1864 (n1308, n_675, n_674);
  and g1865 (n1309, \asqrt[51] , n1308);
  not g1866 (n_790, n1309);
  and g1867 (n1310, n_673, n_790);
  not g1868 (n_791, n1307);
  not g1869 (n_792, n1310);
  and g1870 (n1311, n_791, n_792);
  and g1871 (n1312, n_115, n_787);
  and g1872 (n1313, n_788, n1312);
  not g1873 (n_793, n1311);
  not g1874 (n_794, n1313);
  and g1875 (n1314, n_793, n_794);
  not g1876 (n_795, n1304);
  not g1877 (n_796, n1314);
  and g1878 (n1315, n_795, n_796);
  not g1879 (n_797, n1315);
  and g1880 (n1316, \asqrt[62] , n_797);
  and g1881 (n1317, n_76, n_795);
  and g1882 (n1318, n_796, n1317);
  and g1886 (n1322, n_683, n_681);
  and g1887 (n1323, \asqrt[51] , n1322);
  not g1888 (n_798, n1323);
  and g1889 (n1324, n_682, n_798);
  not g1890 (n_799, n1321);
  not g1891 (n_800, n1324);
  and g1892 (n1325, n_799, n_800);
  not g1893 (n_801, n1318);
  not g1894 (n_802, n1325);
  and g1895 (n1326, n_801, n_802);
  not g1896 (n_803, n1316);
  not g1897 (n_804, n1326);
  and g1898 (n1327, n_803, n_804);
  and g1902 (n1331, n_691, n_690);
  and g1903 (n1332, \asqrt[51] , n1331);
  not g1904 (n_805, n1332);
  and g1905 (n1333, n_689, n_805);
  not g1906 (n_806, n1330);
  not g1907 (n_807, n1333);
  and g1908 (n1334, n_806, n_807);
  and g1909 (n1335, n_698, n_697);
  and g1910 (n1336, \asqrt[51] , n1335);
  not g1913 (n_809, n1334);
  not g1915 (n_810, n1327);
  not g1917 (n_811, n1339);
  and g1918 (n1340, n_21, n_811);
  and g1919 (n1341, n_803, n1334);
  and g1920 (n1342, n_804, n1341);
  and g1921 (n1343, n_697, \asqrt[51] );
  not g1922 (n_812, n1343);
  and g1923 (n1344, n1163, n_812);
  not g1924 (n_813, n1335);
  and g1925 (n1345, \asqrt[63] , n_813);
  not g1926 (n_814, n1344);
  and g1927 (n1346, n_814, n1345);
  not g1933 (n_815, n1346);
  not g1934 (n_816, n1351);
  not g1936 (n_817, n1342);
  and g1940 (n1355, \a[100] , \asqrt[50] );
  not g1941 (n_822, \a[98] );
  not g1942 (n_823, \a[99] );
  and g1943 (n1356, n_822, n_823);
  and g1944 (n1357, n_710, n1356);
  not g1945 (n_824, n1355);
  not g1946 (n_825, n1357);
  and g1947 (n1358, n_824, n_825);
  not g1948 (n_826, n1358);
  and g1949 (n1359, \asqrt[51] , n_826);
  and g1955 (n1365, n_710, \asqrt[50] );
  not g1956 (n_827, n1365);
  and g1957 (n1366, \a[101] , n_827);
  and g1958 (n1367, n1192, \asqrt[50] );
  not g1959 (n_828, n1366);
  not g1960 (n_829, n1367);
  and g1961 (n1368, n_828, n_829);
  not g1962 (n_830, n1364);
  and g1963 (n1369, n_830, n1368);
  not g1964 (n_831, n1359);
  not g1965 (n_832, n1369);
  and g1966 (n1370, n_831, n_832);
  not g1967 (n_833, n1370);
  and g1968 (n1371, \asqrt[52] , n_833);
  not g1969 (n_834, \asqrt[52] );
  and g1970 (n1372, n_834, n_831);
  and g1971 (n1373, n_832, n1372);
  not g1975 (n_835, n1340);
  not g1977 (n_836, n1377);
  and g1978 (n1378, n_829, n_836);
  not g1979 (n_837, n1378);
  and g1980 (n1379, \a[102] , n_837);
  and g1981 (n1380, n_606, n_836);
  and g1982 (n1381, n_829, n1380);
  not g1983 (n_838, n1379);
  not g1984 (n_839, n1381);
  and g1985 (n1382, n_838, n_839);
  not g1986 (n_840, n1373);
  not g1987 (n_841, n1382);
  and g1988 (n1383, n_840, n_841);
  not g1989 (n_842, n1371);
  not g1990 (n_843, n1383);
  and g1991 (n1384, n_842, n_843);
  not g1992 (n_844, n1384);
  and g1993 (n1385, \asqrt[53] , n_844);
  and g1994 (n1386, n_719, n_718);
  not g1995 (n_845, n1204);
  and g1996 (n1387, n_845, n1386);
  and g1997 (n1388, \asqrt[50] , n1387);
  and g1998 (n1389, \asqrt[50] , n1386);
  not g1999 (n_846, n1389);
  and g2000 (n1390, n1204, n_846);
  not g2001 (n_847, n1388);
  not g2002 (n_848, n1390);
  and g2003 (n1391, n_847, n_848);
  and g2004 (n1392, n_722, n_842);
  and g2005 (n1393, n_843, n1392);
  not g2006 (n_849, n1391);
  not g2007 (n_850, n1393);
  and g2008 (n1394, n_849, n_850);
  not g2009 (n_851, n1385);
  not g2010 (n_852, n1394);
  and g2011 (n1395, n_851, n_852);
  not g2012 (n_853, n1395);
  and g2013 (n1396, \asqrt[54] , n_853);
  and g2017 (n1400, n_730, n_728);
  and g2018 (n1401, \asqrt[50] , n1400);
  not g2019 (n_854, n1401);
  and g2020 (n1402, n_729, n_854);
  not g2021 (n_855, n1399);
  not g2022 (n_856, n1402);
  and g2023 (n1403, n_855, n_856);
  and g2024 (n1404, n_618, n_851);
  and g2025 (n1405, n_852, n1404);
  not g2026 (n_857, n1403);
  not g2027 (n_858, n1405);
  and g2028 (n1406, n_857, n_858);
  not g2029 (n_859, n1396);
  not g2030 (n_860, n1406);
  and g2031 (n1407, n_859, n_860);
  not g2032 (n_861, n1407);
  and g2033 (n1408, \asqrt[55] , n_861);
  and g2037 (n1412, n_739, n_738);
  and g2038 (n1413, \asqrt[50] , n1412);
  not g2039 (n_862, n1413);
  and g2040 (n1414, n_737, n_862);
  not g2041 (n_863, n1411);
  not g2042 (n_864, n1414);
  and g2043 (n1415, n_863, n_864);
  and g2044 (n1416, n_522, n_859);
  and g2045 (n1417, n_860, n1416);
  not g2046 (n_865, n1415);
  not g2047 (n_866, n1417);
  and g2048 (n1418, n_865, n_866);
  not g2049 (n_867, n1408);
  not g2050 (n_868, n1418);
  and g2051 (n1419, n_867, n_868);
  not g2052 (n_869, n1419);
  and g2053 (n1420, \asqrt[56] , n_869);
  and g2057 (n1424, n_747, n_746);
  and g2058 (n1425, \asqrt[50] , n1424);
  not g2059 (n_870, n1425);
  and g2060 (n1426, n_745, n_870);
  not g2061 (n_871, n1423);
  not g2062 (n_872, n1426);
  and g2063 (n1427, n_871, n_872);
  and g2064 (n1428, n_434, n_867);
  and g2065 (n1429, n_868, n1428);
  not g2066 (n_873, n1427);
  not g2067 (n_874, n1429);
  and g2068 (n1430, n_873, n_874);
  not g2069 (n_875, n1420);
  not g2070 (n_876, n1430);
  and g2071 (n1431, n_875, n_876);
  not g2072 (n_877, n1431);
  and g2073 (n1432, \asqrt[57] , n_877);
  and g2077 (n1436, n_755, n_754);
  and g2078 (n1437, \asqrt[50] , n1436);
  not g2079 (n_878, n1437);
  and g2080 (n1438, n_753, n_878);
  not g2081 (n_879, n1435);
  not g2082 (n_880, n1438);
  and g2083 (n1439, n_879, n_880);
  and g2084 (n1440, n_354, n_875);
  and g2085 (n1441, n_876, n1440);
  not g2086 (n_881, n1439);
  not g2087 (n_882, n1441);
  and g2088 (n1442, n_881, n_882);
  not g2089 (n_883, n1432);
  not g2090 (n_884, n1442);
  and g2091 (n1443, n_883, n_884);
  not g2092 (n_885, n1443);
  and g2093 (n1444, \asqrt[58] , n_885);
  and g2097 (n1448, n_763, n_762);
  and g2098 (n1449, \asqrt[50] , n1448);
  not g2099 (n_886, n1449);
  and g2100 (n1450, n_761, n_886);
  not g2101 (n_887, n1447);
  not g2102 (n_888, n1450);
  and g2103 (n1451, n_887, n_888);
  and g2104 (n1452, n_282, n_883);
  and g2105 (n1453, n_884, n1452);
  not g2106 (n_889, n1451);
  not g2107 (n_890, n1453);
  and g2108 (n1454, n_889, n_890);
  not g2109 (n_891, n1444);
  not g2110 (n_892, n1454);
  and g2111 (n1455, n_891, n_892);
  not g2112 (n_893, n1455);
  and g2113 (n1456, \asqrt[59] , n_893);
  and g2117 (n1460, n_771, n_770);
  and g2118 (n1461, \asqrt[50] , n1460);
  not g2119 (n_894, n1461);
  and g2120 (n1462, n_769, n_894);
  not g2121 (n_895, n1459);
  not g2122 (n_896, n1462);
  and g2123 (n1463, n_895, n_896);
  and g2124 (n1464, n_218, n_891);
  and g2125 (n1465, n_892, n1464);
  not g2126 (n_897, n1463);
  not g2127 (n_898, n1465);
  and g2128 (n1466, n_897, n_898);
  not g2129 (n_899, n1456);
  not g2130 (n_900, n1466);
  and g2131 (n1467, n_899, n_900);
  not g2132 (n_901, n1467);
  and g2133 (n1468, \asqrt[60] , n_901);
  and g2137 (n1472, n_779, n_778);
  and g2138 (n1473, \asqrt[50] , n1472);
  not g2139 (n_902, n1473);
  and g2140 (n1474, n_777, n_902);
  not g2141 (n_903, n1471);
  not g2142 (n_904, n1474);
  and g2143 (n1475, n_903, n_904);
  and g2144 (n1476, n_162, n_899);
  and g2145 (n1477, n_900, n1476);
  not g2146 (n_905, n1475);
  not g2147 (n_906, n1477);
  and g2148 (n1478, n_905, n_906);
  not g2149 (n_907, n1468);
  not g2150 (n_908, n1478);
  and g2151 (n1479, n_907, n_908);
  not g2152 (n_909, n1479);
  and g2153 (n1480, \asqrt[61] , n_909);
  and g2157 (n1484, n_787, n_786);
  and g2158 (n1485, \asqrt[50] , n1484);
  not g2159 (n_910, n1485);
  and g2160 (n1486, n_785, n_910);
  not g2161 (n_911, n1483);
  not g2162 (n_912, n1486);
  and g2163 (n1487, n_911, n_912);
  and g2164 (n1488, n_115, n_907);
  and g2165 (n1489, n_908, n1488);
  not g2166 (n_913, n1487);
  not g2167 (n_914, n1489);
  and g2168 (n1490, n_913, n_914);
  not g2169 (n_915, n1480);
  not g2170 (n_916, n1490);
  and g2171 (n1491, n_915, n_916);
  not g2172 (n_917, n1491);
  and g2173 (n1492, \asqrt[62] , n_917);
  and g2177 (n1496, n_795, n_794);
  and g2178 (n1497, \asqrt[50] , n1496);
  not g2179 (n_918, n1497);
  and g2180 (n1498, n_793, n_918);
  not g2181 (n_919, n1495);
  not g2182 (n_920, n1498);
  and g2183 (n1499, n_919, n_920);
  and g2184 (n1500, n_76, n_915);
  and g2185 (n1501, n_916, n1500);
  not g2186 (n_921, n1499);
  not g2187 (n_922, n1501);
  and g2188 (n1502, n_921, n_922);
  not g2189 (n_923, n1492);
  not g2190 (n_924, n1502);
  and g2191 (n1503, n_923, n_924);
  and g2195 (n1507, n_803, n_801);
  and g2196 (n1508, \asqrt[50] , n1507);
  not g2197 (n_925, n1508);
  and g2198 (n1509, n_802, n_925);
  not g2199 (n_926, n1506);
  not g2200 (n_927, n1509);
  and g2201 (n1510, n_926, n_927);
  and g2202 (n1511, n_810, n_809);
  and g2203 (n1512, \asqrt[50] , n1511);
  not g2206 (n_929, n1510);
  not g2208 (n_930, n1503);
  not g2210 (n_931, n1515);
  and g2211 (n1516, n_21, n_931);
  and g2212 (n1517, n_923, n1510);
  and g2213 (n1518, n_924, n1517);
  and g2214 (n1519, n_809, \asqrt[50] );
  not g2215 (n_932, n1519);
  and g2216 (n1520, n1327, n_932);
  not g2217 (n_933, n1511);
  and g2218 (n1521, \asqrt[63] , n_933);
  not g2219 (n_934, n1520);
  and g2220 (n1522, n_934, n1521);
  not g2226 (n_935, n1522);
  not g2227 (n_936, n1527);
  not g2229 (n_937, n1518);
  and g2233 (n1531, \a[98] , \asqrt[49] );
  not g2234 (n_942, \a[96] );
  not g2235 (n_943, \a[97] );
  and g2236 (n1532, n_942, n_943);
  and g2237 (n1533, n_822, n1532);
  not g2238 (n_944, n1531);
  not g2239 (n_945, n1533);
  and g2240 (n1534, n_944, n_945);
  not g2241 (n_946, n1534);
  and g2242 (n1535, \asqrt[50] , n_946);
  and g2248 (n1541, n_822, \asqrt[49] );
  not g2249 (n_947, n1541);
  and g2250 (n1542, \a[99] , n_947);
  and g2251 (n1543, n1356, \asqrt[49] );
  not g2252 (n_948, n1542);
  not g2253 (n_949, n1543);
  and g2254 (n1544, n_948, n_949);
  not g2255 (n_950, n1540);
  and g2256 (n1545, n_950, n1544);
  not g2257 (n_951, n1535);
  not g2258 (n_952, n1545);
  and g2259 (n1546, n_951, n_952);
  not g2260 (n_953, n1546);
  and g2261 (n1547, \asqrt[51] , n_953);
  not g2262 (n_954, \asqrt[51] );
  and g2263 (n1548, n_954, n_951);
  and g2264 (n1549, n_952, n1548);
  not g2268 (n_955, n1516);
  not g2270 (n_956, n1553);
  and g2271 (n1554, n_949, n_956);
  not g2272 (n_957, n1554);
  and g2273 (n1555, \a[100] , n_957);
  and g2274 (n1556, n_710, n_956);
  and g2275 (n1557, n_949, n1556);
  not g2276 (n_958, n1555);
  not g2277 (n_959, n1557);
  and g2278 (n1558, n_958, n_959);
  not g2279 (n_960, n1549);
  not g2280 (n_961, n1558);
  and g2281 (n1559, n_960, n_961);
  not g2282 (n_962, n1547);
  not g2283 (n_963, n1559);
  and g2284 (n1560, n_962, n_963);
  not g2285 (n_964, n1560);
  and g2286 (n1561, \asqrt[52] , n_964);
  and g2287 (n1562, n_831, n_830);
  not g2288 (n_965, n1368);
  and g2289 (n1563, n_965, n1562);
  and g2290 (n1564, \asqrt[49] , n1563);
  and g2291 (n1565, \asqrt[49] , n1562);
  not g2292 (n_966, n1565);
  and g2293 (n1566, n1368, n_966);
  not g2294 (n_967, n1564);
  not g2295 (n_968, n1566);
  and g2296 (n1567, n_967, n_968);
  and g2297 (n1568, n_834, n_962);
  and g2298 (n1569, n_963, n1568);
  not g2299 (n_969, n1567);
  not g2300 (n_970, n1569);
  and g2301 (n1570, n_969, n_970);
  not g2302 (n_971, n1561);
  not g2303 (n_972, n1570);
  and g2304 (n1571, n_971, n_972);
  not g2305 (n_973, n1571);
  and g2306 (n1572, \asqrt[53] , n_973);
  and g2310 (n1576, n_842, n_840);
  and g2311 (n1577, \asqrt[49] , n1576);
  not g2312 (n_974, n1577);
  and g2313 (n1578, n_841, n_974);
  not g2314 (n_975, n1575);
  not g2315 (n_976, n1578);
  and g2316 (n1579, n_975, n_976);
  and g2317 (n1580, n_722, n_971);
  and g2318 (n1581, n_972, n1580);
  not g2319 (n_977, n1579);
  not g2320 (n_978, n1581);
  and g2321 (n1582, n_977, n_978);
  not g2322 (n_979, n1572);
  not g2323 (n_980, n1582);
  and g2324 (n1583, n_979, n_980);
  not g2325 (n_981, n1583);
  and g2326 (n1584, \asqrt[54] , n_981);
  and g2330 (n1588, n_851, n_850);
  and g2331 (n1589, \asqrt[49] , n1588);
  not g2332 (n_982, n1589);
  and g2333 (n1590, n_849, n_982);
  not g2334 (n_983, n1587);
  not g2335 (n_984, n1590);
  and g2336 (n1591, n_983, n_984);
  and g2337 (n1592, n_618, n_979);
  and g2338 (n1593, n_980, n1592);
  not g2339 (n_985, n1591);
  not g2340 (n_986, n1593);
  and g2341 (n1594, n_985, n_986);
  not g2342 (n_987, n1584);
  not g2343 (n_988, n1594);
  and g2344 (n1595, n_987, n_988);
  not g2345 (n_989, n1595);
  and g2346 (n1596, \asqrt[55] , n_989);
  and g2350 (n1600, n_859, n_858);
  and g2351 (n1601, \asqrt[49] , n1600);
  not g2352 (n_990, n1601);
  and g2353 (n1602, n_857, n_990);
  not g2354 (n_991, n1599);
  not g2355 (n_992, n1602);
  and g2356 (n1603, n_991, n_992);
  and g2357 (n1604, n_522, n_987);
  and g2358 (n1605, n_988, n1604);
  not g2359 (n_993, n1603);
  not g2360 (n_994, n1605);
  and g2361 (n1606, n_993, n_994);
  not g2362 (n_995, n1596);
  not g2363 (n_996, n1606);
  and g2364 (n1607, n_995, n_996);
  not g2365 (n_997, n1607);
  and g2366 (n1608, \asqrt[56] , n_997);
  and g2370 (n1612, n_867, n_866);
  and g2371 (n1613, \asqrt[49] , n1612);
  not g2372 (n_998, n1613);
  and g2373 (n1614, n_865, n_998);
  not g2374 (n_999, n1611);
  not g2375 (n_1000, n1614);
  and g2376 (n1615, n_999, n_1000);
  and g2377 (n1616, n_434, n_995);
  and g2378 (n1617, n_996, n1616);
  not g2379 (n_1001, n1615);
  not g2380 (n_1002, n1617);
  and g2381 (n1618, n_1001, n_1002);
  not g2382 (n_1003, n1608);
  not g2383 (n_1004, n1618);
  and g2384 (n1619, n_1003, n_1004);
  not g2385 (n_1005, n1619);
  and g2386 (n1620, \asqrt[57] , n_1005);
  and g2390 (n1624, n_875, n_874);
  and g2391 (n1625, \asqrt[49] , n1624);
  not g2392 (n_1006, n1625);
  and g2393 (n1626, n_873, n_1006);
  not g2394 (n_1007, n1623);
  not g2395 (n_1008, n1626);
  and g2396 (n1627, n_1007, n_1008);
  and g2397 (n1628, n_354, n_1003);
  and g2398 (n1629, n_1004, n1628);
  not g2399 (n_1009, n1627);
  not g2400 (n_1010, n1629);
  and g2401 (n1630, n_1009, n_1010);
  not g2402 (n_1011, n1620);
  not g2403 (n_1012, n1630);
  and g2404 (n1631, n_1011, n_1012);
  not g2405 (n_1013, n1631);
  and g2406 (n1632, \asqrt[58] , n_1013);
  and g2410 (n1636, n_883, n_882);
  and g2411 (n1637, \asqrt[49] , n1636);
  not g2412 (n_1014, n1637);
  and g2413 (n1638, n_881, n_1014);
  not g2414 (n_1015, n1635);
  not g2415 (n_1016, n1638);
  and g2416 (n1639, n_1015, n_1016);
  and g2417 (n1640, n_282, n_1011);
  and g2418 (n1641, n_1012, n1640);
  not g2419 (n_1017, n1639);
  not g2420 (n_1018, n1641);
  and g2421 (n1642, n_1017, n_1018);
  not g2422 (n_1019, n1632);
  not g2423 (n_1020, n1642);
  and g2424 (n1643, n_1019, n_1020);
  not g2425 (n_1021, n1643);
  and g2426 (n1644, \asqrt[59] , n_1021);
  and g2430 (n1648, n_891, n_890);
  and g2431 (n1649, \asqrt[49] , n1648);
  not g2432 (n_1022, n1649);
  and g2433 (n1650, n_889, n_1022);
  not g2434 (n_1023, n1647);
  not g2435 (n_1024, n1650);
  and g2436 (n1651, n_1023, n_1024);
  and g2437 (n1652, n_218, n_1019);
  and g2438 (n1653, n_1020, n1652);
  not g2439 (n_1025, n1651);
  not g2440 (n_1026, n1653);
  and g2441 (n1654, n_1025, n_1026);
  not g2442 (n_1027, n1644);
  not g2443 (n_1028, n1654);
  and g2444 (n1655, n_1027, n_1028);
  not g2445 (n_1029, n1655);
  and g2446 (n1656, \asqrt[60] , n_1029);
  and g2450 (n1660, n_899, n_898);
  and g2451 (n1661, \asqrt[49] , n1660);
  not g2452 (n_1030, n1661);
  and g2453 (n1662, n_897, n_1030);
  not g2454 (n_1031, n1659);
  not g2455 (n_1032, n1662);
  and g2456 (n1663, n_1031, n_1032);
  and g2457 (n1664, n_162, n_1027);
  and g2458 (n1665, n_1028, n1664);
  not g2459 (n_1033, n1663);
  not g2460 (n_1034, n1665);
  and g2461 (n1666, n_1033, n_1034);
  not g2462 (n_1035, n1656);
  not g2463 (n_1036, n1666);
  and g2464 (n1667, n_1035, n_1036);
  not g2465 (n_1037, n1667);
  and g2466 (n1668, \asqrt[61] , n_1037);
  and g2470 (n1672, n_907, n_906);
  and g2471 (n1673, \asqrt[49] , n1672);
  not g2472 (n_1038, n1673);
  and g2473 (n1674, n_905, n_1038);
  not g2474 (n_1039, n1671);
  not g2475 (n_1040, n1674);
  and g2476 (n1675, n_1039, n_1040);
  and g2477 (n1676, n_115, n_1035);
  and g2478 (n1677, n_1036, n1676);
  not g2479 (n_1041, n1675);
  not g2480 (n_1042, n1677);
  and g2481 (n1678, n_1041, n_1042);
  not g2482 (n_1043, n1668);
  not g2483 (n_1044, n1678);
  and g2484 (n1679, n_1043, n_1044);
  not g2485 (n_1045, n1679);
  and g2486 (n1680, \asqrt[62] , n_1045);
  and g2490 (n1684, n_915, n_914);
  and g2491 (n1685, \asqrt[49] , n1684);
  not g2492 (n_1046, n1685);
  and g2493 (n1686, n_913, n_1046);
  not g2494 (n_1047, n1683);
  not g2495 (n_1048, n1686);
  and g2496 (n1687, n_1047, n_1048);
  and g2497 (n1688, n_76, n_1043);
  and g2498 (n1689, n_1044, n1688);
  not g2499 (n_1049, n1687);
  not g2500 (n_1050, n1689);
  and g2501 (n1690, n_1049, n_1050);
  not g2502 (n_1051, n1680);
  not g2503 (n_1052, n1690);
  and g2504 (n1691, n_1051, n_1052);
  and g2508 (n1695, n_923, n_922);
  and g2509 (n1696, \asqrt[49] , n1695);
  not g2510 (n_1053, n1696);
  and g2511 (n1697, n_921, n_1053);
  not g2512 (n_1054, n1694);
  not g2513 (n_1055, n1697);
  and g2514 (n1698, n_1054, n_1055);
  and g2515 (n1699, n_930, n_929);
  and g2516 (n1700, \asqrt[49] , n1699);
  not g2519 (n_1057, n1698);
  not g2521 (n_1058, n1691);
  not g2523 (n_1059, n1703);
  and g2524 (n1704, n_21, n_1059);
  and g2525 (n1705, n_1051, n1698);
  and g2526 (n1706, n_1052, n1705);
  and g2527 (n1707, n_929, \asqrt[49] );
  not g2528 (n_1060, n1707);
  and g2529 (n1708, n1503, n_1060);
  not g2530 (n_1061, n1699);
  and g2531 (n1709, \asqrt[63] , n_1061);
  not g2532 (n_1062, n1708);
  and g2533 (n1710, n_1062, n1709);
  not g2539 (n_1063, n1710);
  not g2540 (n_1064, n1715);
  not g2542 (n_1065, n1706);
  and g2546 (n1719, \a[96] , \asqrt[48] );
  not g2547 (n_1070, \a[94] );
  not g2548 (n_1071, \a[95] );
  and g2549 (n1720, n_1070, n_1071);
  and g2550 (n1721, n_942, n1720);
  not g2551 (n_1072, n1719);
  not g2552 (n_1073, n1721);
  and g2553 (n1722, n_1072, n_1073);
  not g2554 (n_1074, n1722);
  and g2555 (n1723, \asqrt[49] , n_1074);
  and g2556 (n1724, n_942, \asqrt[48] );
  not g2557 (n_1075, n1724);
  and g2558 (n1725, \a[97] , n_1075);
  and g2559 (n1726, n1532, \asqrt[48] );
  not g2560 (n_1076, n1725);
  not g2561 (n_1077, n1726);
  and g2562 (n1727, n_1076, n_1077);
  not g2568 (n_1078, n1732);
  and g2569 (n1733, n1727, n_1078);
  not g2570 (n_1079, n1723);
  not g2571 (n_1080, n1733);
  and g2572 (n1734, n_1079, n_1080);
  not g2573 (n_1081, n1734);
  and g2574 (n1735, \asqrt[50] , n_1081);
  not g2575 (n_1082, \asqrt[50] );
  and g2576 (n1736, n_1082, n_1079);
  and g2577 (n1737, n_1080, n1736);
  not g2581 (n_1083, n1704);
  not g2583 (n_1084, n1741);
  and g2584 (n1742, n_1077, n_1084);
  not g2585 (n_1085, n1742);
  and g2586 (n1743, \a[98] , n_1085);
  and g2587 (n1744, n_822, n_1084);
  and g2588 (n1745, n_1077, n1744);
  not g2589 (n_1086, n1743);
  not g2590 (n_1087, n1745);
  and g2591 (n1746, n_1086, n_1087);
  not g2592 (n_1088, n1737);
  not g2593 (n_1089, n1746);
  and g2594 (n1747, n_1088, n_1089);
  not g2595 (n_1090, n1735);
  not g2596 (n_1091, n1747);
  and g2597 (n1748, n_1090, n_1091);
  not g2598 (n_1092, n1748);
  and g2599 (n1749, \asqrt[51] , n_1092);
  and g2600 (n1750, n_951, n_950);
  not g2601 (n_1093, n1544);
  and g2602 (n1751, n_1093, n1750);
  and g2603 (n1752, \asqrt[48] , n1751);
  and g2604 (n1753, \asqrt[48] , n1750);
  not g2605 (n_1094, n1753);
  and g2606 (n1754, n1544, n_1094);
  not g2607 (n_1095, n1752);
  not g2608 (n_1096, n1754);
  and g2609 (n1755, n_1095, n_1096);
  and g2610 (n1756, n_954, n_1090);
  and g2611 (n1757, n_1091, n1756);
  not g2612 (n_1097, n1755);
  not g2613 (n_1098, n1757);
  and g2614 (n1758, n_1097, n_1098);
  not g2615 (n_1099, n1749);
  not g2616 (n_1100, n1758);
  and g2617 (n1759, n_1099, n_1100);
  not g2618 (n_1101, n1759);
  and g2619 (n1760, \asqrt[52] , n_1101);
  and g2623 (n1764, n_962, n_960);
  and g2624 (n1765, \asqrt[48] , n1764);
  not g2625 (n_1102, n1765);
  and g2626 (n1766, n_961, n_1102);
  not g2627 (n_1103, n1763);
  not g2628 (n_1104, n1766);
  and g2629 (n1767, n_1103, n_1104);
  and g2630 (n1768, n_834, n_1099);
  and g2631 (n1769, n_1100, n1768);
  not g2632 (n_1105, n1767);
  not g2633 (n_1106, n1769);
  and g2634 (n1770, n_1105, n_1106);
  not g2635 (n_1107, n1760);
  not g2636 (n_1108, n1770);
  and g2637 (n1771, n_1107, n_1108);
  not g2638 (n_1109, n1771);
  and g2639 (n1772, \asqrt[53] , n_1109);
  and g2643 (n1776, n_971, n_970);
  and g2644 (n1777, \asqrt[48] , n1776);
  not g2645 (n_1110, n1777);
  and g2646 (n1778, n_969, n_1110);
  not g2647 (n_1111, n1775);
  not g2648 (n_1112, n1778);
  and g2649 (n1779, n_1111, n_1112);
  and g2650 (n1780, n_722, n_1107);
  and g2651 (n1781, n_1108, n1780);
  not g2652 (n_1113, n1779);
  not g2653 (n_1114, n1781);
  and g2654 (n1782, n_1113, n_1114);
  not g2655 (n_1115, n1772);
  not g2656 (n_1116, n1782);
  and g2657 (n1783, n_1115, n_1116);
  not g2658 (n_1117, n1783);
  and g2659 (n1784, \asqrt[54] , n_1117);
  and g2663 (n1788, n_979, n_978);
  and g2664 (n1789, \asqrt[48] , n1788);
  not g2665 (n_1118, n1789);
  and g2666 (n1790, n_977, n_1118);
  not g2667 (n_1119, n1787);
  not g2668 (n_1120, n1790);
  and g2669 (n1791, n_1119, n_1120);
  and g2670 (n1792, n_618, n_1115);
  and g2671 (n1793, n_1116, n1792);
  not g2672 (n_1121, n1791);
  not g2673 (n_1122, n1793);
  and g2674 (n1794, n_1121, n_1122);
  not g2675 (n_1123, n1784);
  not g2676 (n_1124, n1794);
  and g2677 (n1795, n_1123, n_1124);
  not g2678 (n_1125, n1795);
  and g2679 (n1796, \asqrt[55] , n_1125);
  and g2683 (n1800, n_987, n_986);
  and g2684 (n1801, \asqrt[48] , n1800);
  not g2685 (n_1126, n1801);
  and g2686 (n1802, n_985, n_1126);
  not g2687 (n_1127, n1799);
  not g2688 (n_1128, n1802);
  and g2689 (n1803, n_1127, n_1128);
  and g2690 (n1804, n_522, n_1123);
  and g2691 (n1805, n_1124, n1804);
  not g2692 (n_1129, n1803);
  not g2693 (n_1130, n1805);
  and g2694 (n1806, n_1129, n_1130);
  not g2695 (n_1131, n1796);
  not g2696 (n_1132, n1806);
  and g2697 (n1807, n_1131, n_1132);
  not g2698 (n_1133, n1807);
  and g2699 (n1808, \asqrt[56] , n_1133);
  and g2703 (n1812, n_995, n_994);
  and g2704 (n1813, \asqrt[48] , n1812);
  not g2705 (n_1134, n1813);
  and g2706 (n1814, n_993, n_1134);
  not g2707 (n_1135, n1811);
  not g2708 (n_1136, n1814);
  and g2709 (n1815, n_1135, n_1136);
  and g2710 (n1816, n_434, n_1131);
  and g2711 (n1817, n_1132, n1816);
  not g2712 (n_1137, n1815);
  not g2713 (n_1138, n1817);
  and g2714 (n1818, n_1137, n_1138);
  not g2715 (n_1139, n1808);
  not g2716 (n_1140, n1818);
  and g2717 (n1819, n_1139, n_1140);
  not g2718 (n_1141, n1819);
  and g2719 (n1820, \asqrt[57] , n_1141);
  and g2723 (n1824, n_1003, n_1002);
  and g2724 (n1825, \asqrt[48] , n1824);
  not g2725 (n_1142, n1825);
  and g2726 (n1826, n_1001, n_1142);
  not g2727 (n_1143, n1823);
  not g2728 (n_1144, n1826);
  and g2729 (n1827, n_1143, n_1144);
  and g2730 (n1828, n_354, n_1139);
  and g2731 (n1829, n_1140, n1828);
  not g2732 (n_1145, n1827);
  not g2733 (n_1146, n1829);
  and g2734 (n1830, n_1145, n_1146);
  not g2735 (n_1147, n1820);
  not g2736 (n_1148, n1830);
  and g2737 (n1831, n_1147, n_1148);
  not g2738 (n_1149, n1831);
  and g2739 (n1832, \asqrt[58] , n_1149);
  and g2743 (n1836, n_1011, n_1010);
  and g2744 (n1837, \asqrt[48] , n1836);
  not g2745 (n_1150, n1837);
  and g2746 (n1838, n_1009, n_1150);
  not g2747 (n_1151, n1835);
  not g2748 (n_1152, n1838);
  and g2749 (n1839, n_1151, n_1152);
  and g2750 (n1840, n_282, n_1147);
  and g2751 (n1841, n_1148, n1840);
  not g2752 (n_1153, n1839);
  not g2753 (n_1154, n1841);
  and g2754 (n1842, n_1153, n_1154);
  not g2755 (n_1155, n1832);
  not g2756 (n_1156, n1842);
  and g2757 (n1843, n_1155, n_1156);
  not g2758 (n_1157, n1843);
  and g2759 (n1844, \asqrt[59] , n_1157);
  and g2763 (n1848, n_1019, n_1018);
  and g2764 (n1849, \asqrt[48] , n1848);
  not g2765 (n_1158, n1849);
  and g2766 (n1850, n_1017, n_1158);
  not g2767 (n_1159, n1847);
  not g2768 (n_1160, n1850);
  and g2769 (n1851, n_1159, n_1160);
  and g2770 (n1852, n_218, n_1155);
  and g2771 (n1853, n_1156, n1852);
  not g2772 (n_1161, n1851);
  not g2773 (n_1162, n1853);
  and g2774 (n1854, n_1161, n_1162);
  not g2775 (n_1163, n1844);
  not g2776 (n_1164, n1854);
  and g2777 (n1855, n_1163, n_1164);
  not g2778 (n_1165, n1855);
  and g2779 (n1856, \asqrt[60] , n_1165);
  and g2783 (n1860, n_1027, n_1026);
  and g2784 (n1861, \asqrt[48] , n1860);
  not g2785 (n_1166, n1861);
  and g2786 (n1862, n_1025, n_1166);
  not g2787 (n_1167, n1859);
  not g2788 (n_1168, n1862);
  and g2789 (n1863, n_1167, n_1168);
  and g2790 (n1864, n_162, n_1163);
  and g2791 (n1865, n_1164, n1864);
  not g2792 (n_1169, n1863);
  not g2793 (n_1170, n1865);
  and g2794 (n1866, n_1169, n_1170);
  not g2795 (n_1171, n1856);
  not g2796 (n_1172, n1866);
  and g2797 (n1867, n_1171, n_1172);
  not g2798 (n_1173, n1867);
  and g2799 (n1868, \asqrt[61] , n_1173);
  and g2803 (n1872, n_1035, n_1034);
  and g2804 (n1873, \asqrt[48] , n1872);
  not g2805 (n_1174, n1873);
  and g2806 (n1874, n_1033, n_1174);
  not g2807 (n_1175, n1871);
  not g2808 (n_1176, n1874);
  and g2809 (n1875, n_1175, n_1176);
  and g2810 (n1876, n_115, n_1171);
  and g2811 (n1877, n_1172, n1876);
  not g2812 (n_1177, n1875);
  not g2813 (n_1178, n1877);
  and g2814 (n1878, n_1177, n_1178);
  not g2815 (n_1179, n1868);
  not g2816 (n_1180, n1878);
  and g2817 (n1879, n_1179, n_1180);
  not g2818 (n_1181, n1879);
  and g2819 (n1880, \asqrt[62] , n_1181);
  and g2823 (n1884, n_1043, n_1042);
  and g2824 (n1885, \asqrt[48] , n1884);
  not g2825 (n_1182, n1885);
  and g2826 (n1886, n_1041, n_1182);
  not g2827 (n_1183, n1883);
  not g2828 (n_1184, n1886);
  and g2829 (n1887, n_1183, n_1184);
  and g2830 (n1888, n_76, n_1179);
  and g2831 (n1889, n_1180, n1888);
  not g2832 (n_1185, n1887);
  not g2833 (n_1186, n1889);
  and g2834 (n1890, n_1185, n_1186);
  not g2835 (n_1187, n1880);
  not g2836 (n_1188, n1890);
  and g2837 (n1891, n_1187, n_1188);
  and g2841 (n1895, n_1051, n_1050);
  and g2842 (n1896, \asqrt[48] , n1895);
  not g2843 (n_1189, n1896);
  and g2844 (n1897, n_1049, n_1189);
  not g2845 (n_1190, n1894);
  not g2846 (n_1191, n1897);
  and g2847 (n1898, n_1190, n_1191);
  and g2848 (n1899, n_1058, n_1057);
  and g2849 (n1900, \asqrt[48] , n1899);
  not g2852 (n_1193, n1898);
  not g2854 (n_1194, n1891);
  not g2856 (n_1195, n1903);
  and g2857 (n1904, n_21, n_1195);
  and g2858 (n1905, n_1187, n1898);
  and g2859 (n1906, n_1188, n1905);
  and g2860 (n1907, n_1057, \asqrt[48] );
  not g2861 (n_1196, n1907);
  and g2862 (n1908, n1691, n_1196);
  not g2863 (n_1197, n1899);
  and g2864 (n1909, \asqrt[63] , n_1197);
  not g2865 (n_1198, n1908);
  and g2866 (n1910, n_1198, n1909);
  not g2872 (n_1199, n1910);
  not g2873 (n_1200, n1915);
  not g2875 (n_1201, n1906);
  and g2879 (n1919, \a[94] , \asqrt[47] );
  not g2880 (n_1206, \a[92] );
  not g2881 (n_1207, \a[93] );
  and g2882 (n1920, n_1206, n_1207);
  and g2883 (n1921, n_1070, n1920);
  not g2884 (n_1208, n1919);
  not g2885 (n_1209, n1921);
  and g2886 (n1922, n_1208, n_1209);
  not g2887 (n_1210, n1922);
  and g2888 (n1923, \asqrt[48] , n_1210);
  and g2894 (n1929, n_1070, \asqrt[47] );
  not g2895 (n_1211, n1929);
  and g2896 (n1930, \a[95] , n_1211);
  and g2897 (n1931, n1720, \asqrt[47] );
  not g2898 (n_1212, n1930);
  not g2899 (n_1213, n1931);
  and g2900 (n1932, n_1212, n_1213);
  not g2901 (n_1214, n1928);
  and g2902 (n1933, n_1214, n1932);
  not g2903 (n_1215, n1923);
  not g2904 (n_1216, n1933);
  and g2905 (n1934, n_1215, n_1216);
  not g2906 (n_1217, n1934);
  and g2907 (n1935, \asqrt[49] , n_1217);
  not g2908 (n_1218, \asqrt[49] );
  and g2909 (n1936, n_1218, n_1215);
  and g2910 (n1937, n_1216, n1936);
  not g2914 (n_1219, n1904);
  not g2916 (n_1220, n1941);
  and g2917 (n1942, n_1213, n_1220);
  not g2918 (n_1221, n1942);
  and g2919 (n1943, \a[96] , n_1221);
  and g2920 (n1944, n_942, n_1220);
  and g2921 (n1945, n_1213, n1944);
  not g2922 (n_1222, n1943);
  not g2923 (n_1223, n1945);
  and g2924 (n1946, n_1222, n_1223);
  not g2925 (n_1224, n1937);
  not g2926 (n_1225, n1946);
  and g2927 (n1947, n_1224, n_1225);
  not g2928 (n_1226, n1935);
  not g2929 (n_1227, n1947);
  and g2930 (n1948, n_1226, n_1227);
  not g2931 (n_1228, n1948);
  and g2932 (n1949, \asqrt[50] , n_1228);
  and g2933 (n1950, n_1082, n_1226);
  and g2934 (n1951, n_1227, n1950);
  and g2939 (n1955, n_1079, n_1078);
  and g2940 (n1956, \asqrt[47] , n1955);
  not g2941 (n_1230, n1956);
  and g2942 (n1957, n1727, n_1230);
  not g2943 (n_1231, n1954);
  not g2944 (n_1232, n1957);
  and g2945 (n1958, n_1231, n_1232);
  not g2946 (n_1233, n1951);
  not g2947 (n_1234, n1958);
  and g2948 (n1959, n_1233, n_1234);
  not g2949 (n_1235, n1949);
  not g2950 (n_1236, n1959);
  and g2951 (n1960, n_1235, n_1236);
  not g2952 (n_1237, n1960);
  and g2953 (n1961, \asqrt[51] , n_1237);
  and g2957 (n1965, n_1090, n_1088);
  and g2958 (n1966, \asqrt[47] , n1965);
  not g2959 (n_1238, n1966);
  and g2960 (n1967, n_1089, n_1238);
  not g2961 (n_1239, n1964);
  not g2962 (n_1240, n1967);
  and g2963 (n1968, n_1239, n_1240);
  and g2964 (n1969, n_954, n_1235);
  and g2965 (n1970, n_1236, n1969);
  not g2966 (n_1241, n1968);
  not g2967 (n_1242, n1970);
  and g2968 (n1971, n_1241, n_1242);
  not g2969 (n_1243, n1961);
  not g2970 (n_1244, n1971);
  and g2971 (n1972, n_1243, n_1244);
  not g2972 (n_1245, n1972);
  and g2973 (n1973, \asqrt[52] , n_1245);
  and g2977 (n1977, n_1099, n_1098);
  and g2978 (n1978, \asqrt[47] , n1977);
  not g2979 (n_1246, n1978);
  and g2980 (n1979, n_1097, n_1246);
  not g2981 (n_1247, n1976);
  not g2982 (n_1248, n1979);
  and g2983 (n1980, n_1247, n_1248);
  and g2984 (n1981, n_834, n_1243);
  and g2985 (n1982, n_1244, n1981);
  not g2986 (n_1249, n1980);
  not g2987 (n_1250, n1982);
  and g2988 (n1983, n_1249, n_1250);
  not g2989 (n_1251, n1973);
  not g2990 (n_1252, n1983);
  and g2991 (n1984, n_1251, n_1252);
  not g2992 (n_1253, n1984);
  and g2993 (n1985, \asqrt[53] , n_1253);
  and g2997 (n1989, n_1107, n_1106);
  and g2998 (n1990, \asqrt[47] , n1989);
  not g2999 (n_1254, n1990);
  and g3000 (n1991, n_1105, n_1254);
  not g3001 (n_1255, n1988);
  not g3002 (n_1256, n1991);
  and g3003 (n1992, n_1255, n_1256);
  and g3004 (n1993, n_722, n_1251);
  and g3005 (n1994, n_1252, n1993);
  not g3006 (n_1257, n1992);
  not g3007 (n_1258, n1994);
  and g3008 (n1995, n_1257, n_1258);
  not g3009 (n_1259, n1985);
  not g3010 (n_1260, n1995);
  and g3011 (n1996, n_1259, n_1260);
  not g3012 (n_1261, n1996);
  and g3013 (n1997, \asqrt[54] , n_1261);
  and g3017 (n2001, n_1115, n_1114);
  and g3018 (n2002, \asqrt[47] , n2001);
  not g3019 (n_1262, n2002);
  and g3020 (n2003, n_1113, n_1262);
  not g3021 (n_1263, n2000);
  not g3022 (n_1264, n2003);
  and g3023 (n2004, n_1263, n_1264);
  and g3024 (n2005, n_618, n_1259);
  and g3025 (n2006, n_1260, n2005);
  not g3026 (n_1265, n2004);
  not g3027 (n_1266, n2006);
  and g3028 (n2007, n_1265, n_1266);
  not g3029 (n_1267, n1997);
  not g3030 (n_1268, n2007);
  and g3031 (n2008, n_1267, n_1268);
  not g3032 (n_1269, n2008);
  and g3033 (n2009, \asqrt[55] , n_1269);
  and g3037 (n2013, n_1123, n_1122);
  and g3038 (n2014, \asqrt[47] , n2013);
  not g3039 (n_1270, n2014);
  and g3040 (n2015, n_1121, n_1270);
  not g3041 (n_1271, n2012);
  not g3042 (n_1272, n2015);
  and g3043 (n2016, n_1271, n_1272);
  and g3044 (n2017, n_522, n_1267);
  and g3045 (n2018, n_1268, n2017);
  not g3046 (n_1273, n2016);
  not g3047 (n_1274, n2018);
  and g3048 (n2019, n_1273, n_1274);
  not g3049 (n_1275, n2009);
  not g3050 (n_1276, n2019);
  and g3051 (n2020, n_1275, n_1276);
  not g3052 (n_1277, n2020);
  and g3053 (n2021, \asqrt[56] , n_1277);
  and g3057 (n2025, n_1131, n_1130);
  and g3058 (n2026, \asqrt[47] , n2025);
  not g3059 (n_1278, n2026);
  and g3060 (n2027, n_1129, n_1278);
  not g3061 (n_1279, n2024);
  not g3062 (n_1280, n2027);
  and g3063 (n2028, n_1279, n_1280);
  and g3064 (n2029, n_434, n_1275);
  and g3065 (n2030, n_1276, n2029);
  not g3066 (n_1281, n2028);
  not g3067 (n_1282, n2030);
  and g3068 (n2031, n_1281, n_1282);
  not g3069 (n_1283, n2021);
  not g3070 (n_1284, n2031);
  and g3071 (n2032, n_1283, n_1284);
  not g3072 (n_1285, n2032);
  and g3073 (n2033, \asqrt[57] , n_1285);
  and g3077 (n2037, n_1139, n_1138);
  and g3078 (n2038, \asqrt[47] , n2037);
  not g3079 (n_1286, n2038);
  and g3080 (n2039, n_1137, n_1286);
  not g3081 (n_1287, n2036);
  not g3082 (n_1288, n2039);
  and g3083 (n2040, n_1287, n_1288);
  and g3084 (n2041, n_354, n_1283);
  and g3085 (n2042, n_1284, n2041);
  not g3086 (n_1289, n2040);
  not g3087 (n_1290, n2042);
  and g3088 (n2043, n_1289, n_1290);
  not g3089 (n_1291, n2033);
  not g3090 (n_1292, n2043);
  and g3091 (n2044, n_1291, n_1292);
  not g3092 (n_1293, n2044);
  and g3093 (n2045, \asqrt[58] , n_1293);
  and g3097 (n2049, n_1147, n_1146);
  and g3098 (n2050, \asqrt[47] , n2049);
  not g3099 (n_1294, n2050);
  and g3100 (n2051, n_1145, n_1294);
  not g3101 (n_1295, n2048);
  not g3102 (n_1296, n2051);
  and g3103 (n2052, n_1295, n_1296);
  and g3104 (n2053, n_282, n_1291);
  and g3105 (n2054, n_1292, n2053);
  not g3106 (n_1297, n2052);
  not g3107 (n_1298, n2054);
  and g3108 (n2055, n_1297, n_1298);
  not g3109 (n_1299, n2045);
  not g3110 (n_1300, n2055);
  and g3111 (n2056, n_1299, n_1300);
  not g3112 (n_1301, n2056);
  and g3113 (n2057, \asqrt[59] , n_1301);
  and g3117 (n2061, n_1155, n_1154);
  and g3118 (n2062, \asqrt[47] , n2061);
  not g3119 (n_1302, n2062);
  and g3120 (n2063, n_1153, n_1302);
  not g3121 (n_1303, n2060);
  not g3122 (n_1304, n2063);
  and g3123 (n2064, n_1303, n_1304);
  and g3124 (n2065, n_218, n_1299);
  and g3125 (n2066, n_1300, n2065);
  not g3126 (n_1305, n2064);
  not g3127 (n_1306, n2066);
  and g3128 (n2067, n_1305, n_1306);
  not g3129 (n_1307, n2057);
  not g3130 (n_1308, n2067);
  and g3131 (n2068, n_1307, n_1308);
  not g3132 (n_1309, n2068);
  and g3133 (n2069, \asqrt[60] , n_1309);
  and g3137 (n2073, n_1163, n_1162);
  and g3138 (n2074, \asqrt[47] , n2073);
  not g3139 (n_1310, n2074);
  and g3140 (n2075, n_1161, n_1310);
  not g3141 (n_1311, n2072);
  not g3142 (n_1312, n2075);
  and g3143 (n2076, n_1311, n_1312);
  and g3144 (n2077, n_162, n_1307);
  and g3145 (n2078, n_1308, n2077);
  not g3146 (n_1313, n2076);
  not g3147 (n_1314, n2078);
  and g3148 (n2079, n_1313, n_1314);
  not g3149 (n_1315, n2069);
  not g3150 (n_1316, n2079);
  and g3151 (n2080, n_1315, n_1316);
  not g3152 (n_1317, n2080);
  and g3153 (n2081, \asqrt[61] , n_1317);
  and g3157 (n2085, n_1171, n_1170);
  and g3158 (n2086, \asqrt[47] , n2085);
  not g3159 (n_1318, n2086);
  and g3160 (n2087, n_1169, n_1318);
  not g3161 (n_1319, n2084);
  not g3162 (n_1320, n2087);
  and g3163 (n2088, n_1319, n_1320);
  and g3164 (n2089, n_115, n_1315);
  and g3165 (n2090, n_1316, n2089);
  not g3166 (n_1321, n2088);
  not g3167 (n_1322, n2090);
  and g3168 (n2091, n_1321, n_1322);
  not g3169 (n_1323, n2081);
  not g3170 (n_1324, n2091);
  and g3171 (n2092, n_1323, n_1324);
  not g3172 (n_1325, n2092);
  and g3173 (n2093, \asqrt[62] , n_1325);
  and g3177 (n2097, n_1179, n_1178);
  and g3178 (n2098, \asqrt[47] , n2097);
  not g3179 (n_1326, n2098);
  and g3180 (n2099, n_1177, n_1326);
  not g3181 (n_1327, n2096);
  not g3182 (n_1328, n2099);
  and g3183 (n2100, n_1327, n_1328);
  and g3184 (n2101, n_76, n_1323);
  and g3185 (n2102, n_1324, n2101);
  not g3186 (n_1329, n2100);
  not g3187 (n_1330, n2102);
  and g3188 (n2103, n_1329, n_1330);
  not g3189 (n_1331, n2093);
  not g3190 (n_1332, n2103);
  and g3191 (n2104, n_1331, n_1332);
  and g3195 (n2108, n_1187, n_1186);
  and g3196 (n2109, \asqrt[47] , n2108);
  not g3197 (n_1333, n2109);
  and g3198 (n2110, n_1185, n_1333);
  not g3199 (n_1334, n2107);
  not g3200 (n_1335, n2110);
  and g3201 (n2111, n_1334, n_1335);
  and g3202 (n2112, n_1194, n_1193);
  and g3203 (n2113, \asqrt[47] , n2112);
  not g3206 (n_1337, n2111);
  not g3208 (n_1338, n2104);
  not g3210 (n_1339, n2116);
  and g3211 (n2117, n_21, n_1339);
  and g3212 (n2118, n_1331, n2111);
  and g3213 (n2119, n_1332, n2118);
  and g3214 (n2120, n_1193, \asqrt[47] );
  not g3215 (n_1340, n2120);
  and g3216 (n2121, n1891, n_1340);
  not g3217 (n_1341, n2112);
  and g3218 (n2122, \asqrt[63] , n_1341);
  not g3219 (n_1342, n2121);
  and g3220 (n2123, n_1342, n2122);
  not g3226 (n_1343, n2123);
  not g3227 (n_1344, n2128);
  not g3229 (n_1345, n2119);
  and g3233 (n2132, \a[92] , \asqrt[46] );
  not g3234 (n_1350, \a[90] );
  not g3235 (n_1351, \a[91] );
  and g3236 (n2133, n_1350, n_1351);
  and g3237 (n2134, n_1206, n2133);
  not g3238 (n_1352, n2132);
  not g3239 (n_1353, n2134);
  and g3240 (n2135, n_1352, n_1353);
  not g3241 (n_1354, n2135);
  and g3242 (n2136, \asqrt[47] , n_1354);
  and g3248 (n2142, n_1206, \asqrt[46] );
  not g3249 (n_1355, n2142);
  and g3250 (n2143, \a[93] , n_1355);
  and g3251 (n2144, n1920, \asqrt[46] );
  not g3252 (n_1356, n2143);
  not g3253 (n_1357, n2144);
  and g3254 (n2145, n_1356, n_1357);
  not g3255 (n_1358, n2141);
  and g3256 (n2146, n_1358, n2145);
  not g3257 (n_1359, n2136);
  not g3258 (n_1360, n2146);
  and g3259 (n2147, n_1359, n_1360);
  not g3260 (n_1361, n2147);
  and g3261 (n2148, \asqrt[48] , n_1361);
  not g3262 (n_1362, \asqrt[48] );
  and g3263 (n2149, n_1362, n_1359);
  and g3264 (n2150, n_1360, n2149);
  not g3268 (n_1363, n2117);
  not g3270 (n_1364, n2154);
  and g3271 (n2155, n_1357, n_1364);
  not g3272 (n_1365, n2155);
  and g3273 (n2156, \a[94] , n_1365);
  and g3274 (n2157, n_1070, n_1364);
  and g3275 (n2158, n_1357, n2157);
  not g3276 (n_1366, n2156);
  not g3277 (n_1367, n2158);
  and g3278 (n2159, n_1366, n_1367);
  not g3279 (n_1368, n2150);
  not g3280 (n_1369, n2159);
  and g3281 (n2160, n_1368, n_1369);
  not g3282 (n_1370, n2148);
  not g3283 (n_1371, n2160);
  and g3284 (n2161, n_1370, n_1371);
  not g3285 (n_1372, n2161);
  and g3286 (n2162, \asqrt[49] , n_1372);
  and g3287 (n2163, n_1215, n_1214);
  not g3288 (n_1373, n1932);
  and g3289 (n2164, n_1373, n2163);
  and g3290 (n2165, \asqrt[46] , n2164);
  and g3291 (n2166, \asqrt[46] , n2163);
  not g3292 (n_1374, n2166);
  and g3293 (n2167, n1932, n_1374);
  not g3294 (n_1375, n2165);
  not g3295 (n_1376, n2167);
  and g3296 (n2168, n_1375, n_1376);
  and g3297 (n2169, n_1218, n_1370);
  and g3298 (n2170, n_1371, n2169);
  not g3299 (n_1377, n2168);
  not g3300 (n_1378, n2170);
  and g3301 (n2171, n_1377, n_1378);
  not g3302 (n_1379, n2162);
  not g3303 (n_1380, n2171);
  and g3304 (n2172, n_1379, n_1380);
  not g3305 (n_1381, n2172);
  and g3306 (n2173, \asqrt[50] , n_1381);
  and g3310 (n2177, n_1226, n_1224);
  and g3311 (n2178, \asqrt[46] , n2177);
  not g3312 (n_1382, n2178);
  and g3313 (n2179, n_1225, n_1382);
  not g3314 (n_1383, n2176);
  not g3315 (n_1384, n2179);
  and g3316 (n2180, n_1383, n_1384);
  and g3317 (n2181, n_1082, n_1379);
  and g3318 (n2182, n_1380, n2181);
  not g3319 (n_1385, n2180);
  not g3320 (n_1386, n2182);
  and g3321 (n2183, n_1385, n_1386);
  not g3322 (n_1387, n2173);
  not g3323 (n_1388, n2183);
  and g3324 (n2184, n_1387, n_1388);
  not g3325 (n_1389, n2184);
  and g3326 (n2185, \asqrt[51] , n_1389);
  and g3327 (n2186, n_954, n_1387);
  and g3328 (n2187, n_1388, n2186);
  and g3332 (n2191, n_1235, n_1233);
  and g3333 (n2192, \asqrt[46] , n2191);
  not g3334 (n_1390, n2192);
  and g3335 (n2193, n_1234, n_1390);
  not g3336 (n_1391, n2190);
  not g3337 (n_1392, n2193);
  and g3338 (n2194, n_1391, n_1392);
  not g3339 (n_1393, n2187);
  not g3340 (n_1394, n2194);
  and g3341 (n2195, n_1393, n_1394);
  not g3342 (n_1395, n2185);
  not g3343 (n_1396, n2195);
  and g3344 (n2196, n_1395, n_1396);
  not g3345 (n_1397, n2196);
  and g3346 (n2197, \asqrt[52] , n_1397);
  and g3350 (n2201, n_1243, n_1242);
  and g3351 (n2202, \asqrt[46] , n2201);
  not g3352 (n_1398, n2202);
  and g3353 (n2203, n_1241, n_1398);
  not g3354 (n_1399, n2200);
  not g3355 (n_1400, n2203);
  and g3356 (n2204, n_1399, n_1400);
  and g3357 (n2205, n_834, n_1395);
  and g3358 (n2206, n_1396, n2205);
  not g3359 (n_1401, n2204);
  not g3360 (n_1402, n2206);
  and g3361 (n2207, n_1401, n_1402);
  not g3362 (n_1403, n2197);
  not g3363 (n_1404, n2207);
  and g3364 (n2208, n_1403, n_1404);
  not g3365 (n_1405, n2208);
  and g3366 (n2209, \asqrt[53] , n_1405);
  and g3370 (n2213, n_1251, n_1250);
  and g3371 (n2214, \asqrt[46] , n2213);
  not g3372 (n_1406, n2214);
  and g3373 (n2215, n_1249, n_1406);
  not g3374 (n_1407, n2212);
  not g3375 (n_1408, n2215);
  and g3376 (n2216, n_1407, n_1408);
  and g3377 (n2217, n_722, n_1403);
  and g3378 (n2218, n_1404, n2217);
  not g3379 (n_1409, n2216);
  not g3380 (n_1410, n2218);
  and g3381 (n2219, n_1409, n_1410);
  not g3382 (n_1411, n2209);
  not g3383 (n_1412, n2219);
  and g3384 (n2220, n_1411, n_1412);
  not g3385 (n_1413, n2220);
  and g3386 (n2221, \asqrt[54] , n_1413);
  and g3390 (n2225, n_1259, n_1258);
  and g3391 (n2226, \asqrt[46] , n2225);
  not g3392 (n_1414, n2226);
  and g3393 (n2227, n_1257, n_1414);
  not g3394 (n_1415, n2224);
  not g3395 (n_1416, n2227);
  and g3396 (n2228, n_1415, n_1416);
  and g3397 (n2229, n_618, n_1411);
  and g3398 (n2230, n_1412, n2229);
  not g3399 (n_1417, n2228);
  not g3400 (n_1418, n2230);
  and g3401 (n2231, n_1417, n_1418);
  not g3402 (n_1419, n2221);
  not g3403 (n_1420, n2231);
  and g3404 (n2232, n_1419, n_1420);
  not g3405 (n_1421, n2232);
  and g3406 (n2233, \asqrt[55] , n_1421);
  and g3410 (n2237, n_1267, n_1266);
  and g3411 (n2238, \asqrt[46] , n2237);
  not g3412 (n_1422, n2238);
  and g3413 (n2239, n_1265, n_1422);
  not g3414 (n_1423, n2236);
  not g3415 (n_1424, n2239);
  and g3416 (n2240, n_1423, n_1424);
  and g3417 (n2241, n_522, n_1419);
  and g3418 (n2242, n_1420, n2241);
  not g3419 (n_1425, n2240);
  not g3420 (n_1426, n2242);
  and g3421 (n2243, n_1425, n_1426);
  not g3422 (n_1427, n2233);
  not g3423 (n_1428, n2243);
  and g3424 (n2244, n_1427, n_1428);
  not g3425 (n_1429, n2244);
  and g3426 (n2245, \asqrt[56] , n_1429);
  and g3430 (n2249, n_1275, n_1274);
  and g3431 (n2250, \asqrt[46] , n2249);
  not g3432 (n_1430, n2250);
  and g3433 (n2251, n_1273, n_1430);
  not g3434 (n_1431, n2248);
  not g3435 (n_1432, n2251);
  and g3436 (n2252, n_1431, n_1432);
  and g3437 (n2253, n_434, n_1427);
  and g3438 (n2254, n_1428, n2253);
  not g3439 (n_1433, n2252);
  not g3440 (n_1434, n2254);
  and g3441 (n2255, n_1433, n_1434);
  not g3442 (n_1435, n2245);
  not g3443 (n_1436, n2255);
  and g3444 (n2256, n_1435, n_1436);
  not g3445 (n_1437, n2256);
  and g3446 (n2257, \asqrt[57] , n_1437);
  and g3450 (n2261, n_1283, n_1282);
  and g3451 (n2262, \asqrt[46] , n2261);
  not g3452 (n_1438, n2262);
  and g3453 (n2263, n_1281, n_1438);
  not g3454 (n_1439, n2260);
  not g3455 (n_1440, n2263);
  and g3456 (n2264, n_1439, n_1440);
  and g3457 (n2265, n_354, n_1435);
  and g3458 (n2266, n_1436, n2265);
  not g3459 (n_1441, n2264);
  not g3460 (n_1442, n2266);
  and g3461 (n2267, n_1441, n_1442);
  not g3462 (n_1443, n2257);
  not g3463 (n_1444, n2267);
  and g3464 (n2268, n_1443, n_1444);
  not g3465 (n_1445, n2268);
  and g3466 (n2269, \asqrt[58] , n_1445);
  and g3470 (n2273, n_1291, n_1290);
  and g3471 (n2274, \asqrt[46] , n2273);
  not g3472 (n_1446, n2274);
  and g3473 (n2275, n_1289, n_1446);
  not g3474 (n_1447, n2272);
  not g3475 (n_1448, n2275);
  and g3476 (n2276, n_1447, n_1448);
  and g3477 (n2277, n_282, n_1443);
  and g3478 (n2278, n_1444, n2277);
  not g3479 (n_1449, n2276);
  not g3480 (n_1450, n2278);
  and g3481 (n2279, n_1449, n_1450);
  not g3482 (n_1451, n2269);
  not g3483 (n_1452, n2279);
  and g3484 (n2280, n_1451, n_1452);
  not g3485 (n_1453, n2280);
  and g3486 (n2281, \asqrt[59] , n_1453);
  and g3490 (n2285, n_1299, n_1298);
  and g3491 (n2286, \asqrt[46] , n2285);
  not g3492 (n_1454, n2286);
  and g3493 (n2287, n_1297, n_1454);
  not g3494 (n_1455, n2284);
  not g3495 (n_1456, n2287);
  and g3496 (n2288, n_1455, n_1456);
  and g3497 (n2289, n_218, n_1451);
  and g3498 (n2290, n_1452, n2289);
  not g3499 (n_1457, n2288);
  not g3500 (n_1458, n2290);
  and g3501 (n2291, n_1457, n_1458);
  not g3502 (n_1459, n2281);
  not g3503 (n_1460, n2291);
  and g3504 (n2292, n_1459, n_1460);
  not g3505 (n_1461, n2292);
  and g3506 (n2293, \asqrt[60] , n_1461);
  and g3510 (n2297, n_1307, n_1306);
  and g3511 (n2298, \asqrt[46] , n2297);
  not g3512 (n_1462, n2298);
  and g3513 (n2299, n_1305, n_1462);
  not g3514 (n_1463, n2296);
  not g3515 (n_1464, n2299);
  and g3516 (n2300, n_1463, n_1464);
  and g3517 (n2301, n_162, n_1459);
  and g3518 (n2302, n_1460, n2301);
  not g3519 (n_1465, n2300);
  not g3520 (n_1466, n2302);
  and g3521 (n2303, n_1465, n_1466);
  not g3522 (n_1467, n2293);
  not g3523 (n_1468, n2303);
  and g3524 (n2304, n_1467, n_1468);
  not g3525 (n_1469, n2304);
  and g3526 (n2305, \asqrt[61] , n_1469);
  and g3530 (n2309, n_1315, n_1314);
  and g3531 (n2310, \asqrt[46] , n2309);
  not g3532 (n_1470, n2310);
  and g3533 (n2311, n_1313, n_1470);
  not g3534 (n_1471, n2308);
  not g3535 (n_1472, n2311);
  and g3536 (n2312, n_1471, n_1472);
  and g3537 (n2313, n_115, n_1467);
  and g3538 (n2314, n_1468, n2313);
  not g3539 (n_1473, n2312);
  not g3540 (n_1474, n2314);
  and g3541 (n2315, n_1473, n_1474);
  not g3542 (n_1475, n2305);
  not g3543 (n_1476, n2315);
  and g3544 (n2316, n_1475, n_1476);
  not g3545 (n_1477, n2316);
  and g3546 (n2317, \asqrt[62] , n_1477);
  and g3550 (n2321, n_1323, n_1322);
  and g3551 (n2322, \asqrt[46] , n2321);
  not g3552 (n_1478, n2322);
  and g3553 (n2323, n_1321, n_1478);
  not g3554 (n_1479, n2320);
  not g3555 (n_1480, n2323);
  and g3556 (n2324, n_1479, n_1480);
  and g3557 (n2325, n_76, n_1475);
  and g3558 (n2326, n_1476, n2325);
  not g3559 (n_1481, n2324);
  not g3560 (n_1482, n2326);
  and g3561 (n2327, n_1481, n_1482);
  not g3562 (n_1483, n2317);
  not g3563 (n_1484, n2327);
  and g3564 (n2328, n_1483, n_1484);
  and g3568 (n2332, n_1331, n_1330);
  and g3569 (n2333, \asqrt[46] , n2332);
  not g3570 (n_1485, n2333);
  and g3571 (n2334, n_1329, n_1485);
  not g3572 (n_1486, n2331);
  not g3573 (n_1487, n2334);
  and g3574 (n2335, n_1486, n_1487);
  and g3575 (n2336, n_1338, n_1337);
  and g3576 (n2337, \asqrt[46] , n2336);
  not g3579 (n_1489, n2335);
  not g3581 (n_1490, n2328);
  not g3583 (n_1491, n2340);
  and g3584 (n2341, n_21, n_1491);
  and g3585 (n2342, n_1483, n2335);
  and g3586 (n2343, n_1484, n2342);
  and g3587 (n2344, n_1337, \asqrt[46] );
  not g3588 (n_1492, n2344);
  and g3589 (n2345, n2104, n_1492);
  not g3590 (n_1493, n2336);
  and g3591 (n2346, \asqrt[63] , n_1493);
  not g3592 (n_1494, n2345);
  and g3593 (n2347, n_1494, n2346);
  not g3599 (n_1495, n2347);
  not g3600 (n_1496, n2352);
  not g3602 (n_1497, n2343);
  and g3606 (n2356, \a[90] , \asqrt[45] );
  not g3607 (n_1502, \a[88] );
  not g3608 (n_1503, \a[89] );
  and g3609 (n2357, n_1502, n_1503);
  and g3610 (n2358, n_1350, n2357);
  not g3611 (n_1504, n2356);
  not g3612 (n_1505, n2358);
  and g3613 (n2359, n_1504, n_1505);
  not g3614 (n_1506, n2359);
  and g3615 (n2360, \asqrt[46] , n_1506);
  and g3621 (n2366, n_1350, \asqrt[45] );
  not g3622 (n_1507, n2366);
  and g3623 (n2367, \a[91] , n_1507);
  and g3624 (n2368, n2133, \asqrt[45] );
  not g3625 (n_1508, n2367);
  not g3626 (n_1509, n2368);
  and g3627 (n2369, n_1508, n_1509);
  not g3628 (n_1510, n2365);
  and g3629 (n2370, n_1510, n2369);
  not g3630 (n_1511, n2360);
  not g3631 (n_1512, n2370);
  and g3632 (n2371, n_1511, n_1512);
  not g3633 (n_1513, n2371);
  and g3634 (n2372, \asqrt[47] , n_1513);
  not g3635 (n_1514, \asqrt[47] );
  and g3636 (n2373, n_1514, n_1511);
  and g3637 (n2374, n_1512, n2373);
  not g3641 (n_1515, n2341);
  not g3643 (n_1516, n2378);
  and g3644 (n2379, n_1509, n_1516);
  not g3645 (n_1517, n2379);
  and g3646 (n2380, \a[92] , n_1517);
  and g3647 (n2381, n_1206, n_1516);
  and g3648 (n2382, n_1509, n2381);
  not g3649 (n_1518, n2380);
  not g3650 (n_1519, n2382);
  and g3651 (n2383, n_1518, n_1519);
  not g3652 (n_1520, n2374);
  not g3653 (n_1521, n2383);
  and g3654 (n2384, n_1520, n_1521);
  not g3655 (n_1522, n2372);
  not g3656 (n_1523, n2384);
  and g3657 (n2385, n_1522, n_1523);
  not g3658 (n_1524, n2385);
  and g3659 (n2386, \asqrt[48] , n_1524);
  and g3660 (n2387, n_1359, n_1358);
  not g3661 (n_1525, n2145);
  and g3662 (n2388, n_1525, n2387);
  and g3663 (n2389, \asqrt[45] , n2388);
  and g3664 (n2390, \asqrt[45] , n2387);
  not g3665 (n_1526, n2390);
  and g3666 (n2391, n2145, n_1526);
  not g3667 (n_1527, n2389);
  not g3668 (n_1528, n2391);
  and g3669 (n2392, n_1527, n_1528);
  and g3670 (n2393, n_1362, n_1522);
  and g3671 (n2394, n_1523, n2393);
  not g3672 (n_1529, n2392);
  not g3673 (n_1530, n2394);
  and g3674 (n2395, n_1529, n_1530);
  not g3675 (n_1531, n2386);
  not g3676 (n_1532, n2395);
  and g3677 (n2396, n_1531, n_1532);
  not g3678 (n_1533, n2396);
  and g3679 (n2397, \asqrt[49] , n_1533);
  and g3683 (n2401, n_1370, n_1368);
  and g3684 (n2402, \asqrt[45] , n2401);
  not g3685 (n_1534, n2402);
  and g3686 (n2403, n_1369, n_1534);
  not g3687 (n_1535, n2400);
  not g3688 (n_1536, n2403);
  and g3689 (n2404, n_1535, n_1536);
  and g3690 (n2405, n_1218, n_1531);
  and g3691 (n2406, n_1532, n2405);
  not g3692 (n_1537, n2404);
  not g3693 (n_1538, n2406);
  and g3694 (n2407, n_1537, n_1538);
  not g3695 (n_1539, n2397);
  not g3696 (n_1540, n2407);
  and g3697 (n2408, n_1539, n_1540);
  not g3698 (n_1541, n2408);
  and g3699 (n2409, \asqrt[50] , n_1541);
  and g3703 (n2413, n_1379, n_1378);
  and g3704 (n2414, \asqrt[45] , n2413);
  not g3705 (n_1542, n2414);
  and g3706 (n2415, n_1377, n_1542);
  not g3707 (n_1543, n2412);
  not g3708 (n_1544, n2415);
  and g3709 (n2416, n_1543, n_1544);
  and g3710 (n2417, n_1082, n_1539);
  and g3711 (n2418, n_1540, n2417);
  not g3712 (n_1545, n2416);
  not g3713 (n_1546, n2418);
  and g3714 (n2419, n_1545, n_1546);
  not g3715 (n_1547, n2409);
  not g3716 (n_1548, n2419);
  and g3717 (n2420, n_1547, n_1548);
  not g3718 (n_1549, n2420);
  and g3719 (n2421, \asqrt[51] , n_1549);
  and g3723 (n2425, n_1387, n_1386);
  and g3724 (n2426, \asqrt[45] , n2425);
  not g3725 (n_1550, n2426);
  and g3726 (n2427, n_1385, n_1550);
  not g3727 (n_1551, n2424);
  not g3728 (n_1552, n2427);
  and g3729 (n2428, n_1551, n_1552);
  and g3730 (n2429, n_954, n_1547);
  and g3731 (n2430, n_1548, n2429);
  not g3732 (n_1553, n2428);
  not g3733 (n_1554, n2430);
  and g3734 (n2431, n_1553, n_1554);
  not g3735 (n_1555, n2421);
  not g3736 (n_1556, n2431);
  and g3737 (n2432, n_1555, n_1556);
  not g3738 (n_1557, n2432);
  and g3739 (n2433, \asqrt[52] , n_1557);
  and g3740 (n2434, n_834, n_1555);
  and g3741 (n2435, n_1556, n2434);
  and g3745 (n2439, n_1395, n_1393);
  and g3746 (n2440, \asqrt[45] , n2439);
  not g3747 (n_1558, n2440);
  and g3748 (n2441, n_1394, n_1558);
  not g3749 (n_1559, n2438);
  not g3750 (n_1560, n2441);
  and g3751 (n2442, n_1559, n_1560);
  not g3752 (n_1561, n2435);
  not g3753 (n_1562, n2442);
  and g3754 (n2443, n_1561, n_1562);
  not g3755 (n_1563, n2433);
  not g3756 (n_1564, n2443);
  and g3757 (n2444, n_1563, n_1564);
  not g3758 (n_1565, n2444);
  and g3759 (n2445, \asqrt[53] , n_1565);
  and g3763 (n2449, n_1403, n_1402);
  and g3764 (n2450, \asqrt[45] , n2449);
  not g3765 (n_1566, n2450);
  and g3766 (n2451, n_1401, n_1566);
  not g3767 (n_1567, n2448);
  not g3768 (n_1568, n2451);
  and g3769 (n2452, n_1567, n_1568);
  and g3770 (n2453, n_722, n_1563);
  and g3771 (n2454, n_1564, n2453);
  not g3772 (n_1569, n2452);
  not g3773 (n_1570, n2454);
  and g3774 (n2455, n_1569, n_1570);
  not g3775 (n_1571, n2445);
  not g3776 (n_1572, n2455);
  and g3777 (n2456, n_1571, n_1572);
  not g3778 (n_1573, n2456);
  and g3779 (n2457, \asqrt[54] , n_1573);
  and g3783 (n2461, n_1411, n_1410);
  and g3784 (n2462, \asqrt[45] , n2461);
  not g3785 (n_1574, n2462);
  and g3786 (n2463, n_1409, n_1574);
  not g3787 (n_1575, n2460);
  not g3788 (n_1576, n2463);
  and g3789 (n2464, n_1575, n_1576);
  and g3790 (n2465, n_618, n_1571);
  and g3791 (n2466, n_1572, n2465);
  not g3792 (n_1577, n2464);
  not g3793 (n_1578, n2466);
  and g3794 (n2467, n_1577, n_1578);
  not g3795 (n_1579, n2457);
  not g3796 (n_1580, n2467);
  and g3797 (n2468, n_1579, n_1580);
  not g3798 (n_1581, n2468);
  and g3799 (n2469, \asqrt[55] , n_1581);
  and g3803 (n2473, n_1419, n_1418);
  and g3804 (n2474, \asqrt[45] , n2473);
  not g3805 (n_1582, n2474);
  and g3806 (n2475, n_1417, n_1582);
  not g3807 (n_1583, n2472);
  not g3808 (n_1584, n2475);
  and g3809 (n2476, n_1583, n_1584);
  and g3810 (n2477, n_522, n_1579);
  and g3811 (n2478, n_1580, n2477);
  not g3812 (n_1585, n2476);
  not g3813 (n_1586, n2478);
  and g3814 (n2479, n_1585, n_1586);
  not g3815 (n_1587, n2469);
  not g3816 (n_1588, n2479);
  and g3817 (n2480, n_1587, n_1588);
  not g3818 (n_1589, n2480);
  and g3819 (n2481, \asqrt[56] , n_1589);
  and g3823 (n2485, n_1427, n_1426);
  and g3824 (n2486, \asqrt[45] , n2485);
  not g3825 (n_1590, n2486);
  and g3826 (n2487, n_1425, n_1590);
  not g3827 (n_1591, n2484);
  not g3828 (n_1592, n2487);
  and g3829 (n2488, n_1591, n_1592);
  and g3830 (n2489, n_434, n_1587);
  and g3831 (n2490, n_1588, n2489);
  not g3832 (n_1593, n2488);
  not g3833 (n_1594, n2490);
  and g3834 (n2491, n_1593, n_1594);
  not g3835 (n_1595, n2481);
  not g3836 (n_1596, n2491);
  and g3837 (n2492, n_1595, n_1596);
  not g3838 (n_1597, n2492);
  and g3839 (n2493, \asqrt[57] , n_1597);
  and g3843 (n2497, n_1435, n_1434);
  and g3844 (n2498, \asqrt[45] , n2497);
  not g3845 (n_1598, n2498);
  and g3846 (n2499, n_1433, n_1598);
  not g3847 (n_1599, n2496);
  not g3848 (n_1600, n2499);
  and g3849 (n2500, n_1599, n_1600);
  and g3850 (n2501, n_354, n_1595);
  and g3851 (n2502, n_1596, n2501);
  not g3852 (n_1601, n2500);
  not g3853 (n_1602, n2502);
  and g3854 (n2503, n_1601, n_1602);
  not g3855 (n_1603, n2493);
  not g3856 (n_1604, n2503);
  and g3857 (n2504, n_1603, n_1604);
  not g3858 (n_1605, n2504);
  and g3859 (n2505, \asqrt[58] , n_1605);
  and g3863 (n2509, n_1443, n_1442);
  and g3864 (n2510, \asqrt[45] , n2509);
  not g3865 (n_1606, n2510);
  and g3866 (n2511, n_1441, n_1606);
  not g3867 (n_1607, n2508);
  not g3868 (n_1608, n2511);
  and g3869 (n2512, n_1607, n_1608);
  and g3870 (n2513, n_282, n_1603);
  and g3871 (n2514, n_1604, n2513);
  not g3872 (n_1609, n2512);
  not g3873 (n_1610, n2514);
  and g3874 (n2515, n_1609, n_1610);
  not g3875 (n_1611, n2505);
  not g3876 (n_1612, n2515);
  and g3877 (n2516, n_1611, n_1612);
  not g3878 (n_1613, n2516);
  and g3879 (n2517, \asqrt[59] , n_1613);
  and g3883 (n2521, n_1451, n_1450);
  and g3884 (n2522, \asqrt[45] , n2521);
  not g3885 (n_1614, n2522);
  and g3886 (n2523, n_1449, n_1614);
  not g3887 (n_1615, n2520);
  not g3888 (n_1616, n2523);
  and g3889 (n2524, n_1615, n_1616);
  and g3890 (n2525, n_218, n_1611);
  and g3891 (n2526, n_1612, n2525);
  not g3892 (n_1617, n2524);
  not g3893 (n_1618, n2526);
  and g3894 (n2527, n_1617, n_1618);
  not g3895 (n_1619, n2517);
  not g3896 (n_1620, n2527);
  and g3897 (n2528, n_1619, n_1620);
  not g3898 (n_1621, n2528);
  and g3899 (n2529, \asqrt[60] , n_1621);
  and g3903 (n2533, n_1459, n_1458);
  and g3904 (n2534, \asqrt[45] , n2533);
  not g3905 (n_1622, n2534);
  and g3906 (n2535, n_1457, n_1622);
  not g3907 (n_1623, n2532);
  not g3908 (n_1624, n2535);
  and g3909 (n2536, n_1623, n_1624);
  and g3910 (n2537, n_162, n_1619);
  and g3911 (n2538, n_1620, n2537);
  not g3912 (n_1625, n2536);
  not g3913 (n_1626, n2538);
  and g3914 (n2539, n_1625, n_1626);
  not g3915 (n_1627, n2529);
  not g3916 (n_1628, n2539);
  and g3917 (n2540, n_1627, n_1628);
  not g3918 (n_1629, n2540);
  and g3919 (n2541, \asqrt[61] , n_1629);
  and g3923 (n2545, n_1467, n_1466);
  and g3924 (n2546, \asqrt[45] , n2545);
  not g3925 (n_1630, n2546);
  and g3926 (n2547, n_1465, n_1630);
  not g3927 (n_1631, n2544);
  not g3928 (n_1632, n2547);
  and g3929 (n2548, n_1631, n_1632);
  and g3930 (n2549, n_115, n_1627);
  and g3931 (n2550, n_1628, n2549);
  not g3932 (n_1633, n2548);
  not g3933 (n_1634, n2550);
  and g3934 (n2551, n_1633, n_1634);
  not g3935 (n_1635, n2541);
  not g3936 (n_1636, n2551);
  and g3937 (n2552, n_1635, n_1636);
  not g3938 (n_1637, n2552);
  and g3939 (n2553, \asqrt[62] , n_1637);
  and g3943 (n2557, n_1475, n_1474);
  and g3944 (n2558, \asqrt[45] , n2557);
  not g3945 (n_1638, n2558);
  and g3946 (n2559, n_1473, n_1638);
  not g3947 (n_1639, n2556);
  not g3948 (n_1640, n2559);
  and g3949 (n2560, n_1639, n_1640);
  and g3950 (n2561, n_76, n_1635);
  and g3951 (n2562, n_1636, n2561);
  not g3952 (n_1641, n2560);
  not g3953 (n_1642, n2562);
  and g3954 (n2563, n_1641, n_1642);
  not g3955 (n_1643, n2553);
  not g3956 (n_1644, n2563);
  and g3957 (n2564, n_1643, n_1644);
  and g3961 (n2568, n_1483, n_1482);
  and g3962 (n2569, \asqrt[45] , n2568);
  not g3963 (n_1645, n2569);
  and g3964 (n2570, n_1481, n_1645);
  not g3965 (n_1646, n2567);
  not g3966 (n_1647, n2570);
  and g3967 (n2571, n_1646, n_1647);
  and g3968 (n2572, n_1490, n_1489);
  and g3969 (n2573, \asqrt[45] , n2572);
  not g3972 (n_1649, n2571);
  not g3974 (n_1650, n2564);
  not g3976 (n_1651, n2576);
  and g3977 (n2577, n_21, n_1651);
  and g3978 (n2578, n_1643, n2571);
  and g3979 (n2579, n_1644, n2578);
  and g3980 (n2580, n_1489, \asqrt[45] );
  not g3981 (n_1652, n2580);
  and g3982 (n2581, n2328, n_1652);
  not g3983 (n_1653, n2572);
  and g3984 (n2582, \asqrt[63] , n_1653);
  not g3985 (n_1654, n2581);
  and g3986 (n2583, n_1654, n2582);
  not g3992 (n_1655, n2583);
  not g3993 (n_1656, n2588);
  not g3995 (n_1657, n2579);
  and g3999 (n2592, \a[88] , \asqrt[44] );
  not g4000 (n_1662, \a[86] );
  not g4001 (n_1663, \a[87] );
  and g4002 (n2593, n_1662, n_1663);
  and g4003 (n2594, n_1502, n2593);
  not g4004 (n_1664, n2592);
  not g4005 (n_1665, n2594);
  and g4006 (n2595, n_1664, n_1665);
  not g4007 (n_1666, n2595);
  and g4008 (n2596, \asqrt[45] , n_1666);
  and g4014 (n2602, n_1502, \asqrt[44] );
  not g4015 (n_1667, n2602);
  and g4016 (n2603, \a[89] , n_1667);
  and g4017 (n2604, n2357, \asqrt[44] );
  not g4018 (n_1668, n2603);
  not g4019 (n_1669, n2604);
  and g4020 (n2605, n_1668, n_1669);
  not g4021 (n_1670, n2601);
  and g4022 (n2606, n_1670, n2605);
  not g4023 (n_1671, n2596);
  not g4024 (n_1672, n2606);
  and g4025 (n2607, n_1671, n_1672);
  not g4026 (n_1673, n2607);
  and g4027 (n2608, \asqrt[46] , n_1673);
  not g4028 (n_1674, \asqrt[46] );
  and g4029 (n2609, n_1674, n_1671);
  and g4030 (n2610, n_1672, n2609);
  not g4034 (n_1675, n2577);
  not g4036 (n_1676, n2614);
  and g4037 (n2615, n_1669, n_1676);
  not g4038 (n_1677, n2615);
  and g4039 (n2616, \a[90] , n_1677);
  and g4040 (n2617, n_1350, n_1676);
  and g4041 (n2618, n_1669, n2617);
  not g4042 (n_1678, n2616);
  not g4043 (n_1679, n2618);
  and g4044 (n2619, n_1678, n_1679);
  not g4045 (n_1680, n2610);
  not g4046 (n_1681, n2619);
  and g4047 (n2620, n_1680, n_1681);
  not g4048 (n_1682, n2608);
  not g4049 (n_1683, n2620);
  and g4050 (n2621, n_1682, n_1683);
  not g4051 (n_1684, n2621);
  and g4052 (n2622, \asqrt[47] , n_1684);
  and g4053 (n2623, n_1511, n_1510);
  not g4054 (n_1685, n2369);
  and g4055 (n2624, n_1685, n2623);
  and g4056 (n2625, \asqrt[44] , n2624);
  and g4057 (n2626, \asqrt[44] , n2623);
  not g4058 (n_1686, n2626);
  and g4059 (n2627, n2369, n_1686);
  not g4060 (n_1687, n2625);
  not g4061 (n_1688, n2627);
  and g4062 (n2628, n_1687, n_1688);
  and g4063 (n2629, n_1514, n_1682);
  and g4064 (n2630, n_1683, n2629);
  not g4065 (n_1689, n2628);
  not g4066 (n_1690, n2630);
  and g4067 (n2631, n_1689, n_1690);
  not g4068 (n_1691, n2622);
  not g4069 (n_1692, n2631);
  and g4070 (n2632, n_1691, n_1692);
  not g4071 (n_1693, n2632);
  and g4072 (n2633, \asqrt[48] , n_1693);
  and g4076 (n2637, n_1522, n_1520);
  and g4077 (n2638, \asqrt[44] , n2637);
  not g4078 (n_1694, n2638);
  and g4079 (n2639, n_1521, n_1694);
  not g4080 (n_1695, n2636);
  not g4081 (n_1696, n2639);
  and g4082 (n2640, n_1695, n_1696);
  and g4083 (n2641, n_1362, n_1691);
  and g4084 (n2642, n_1692, n2641);
  not g4085 (n_1697, n2640);
  not g4086 (n_1698, n2642);
  and g4087 (n2643, n_1697, n_1698);
  not g4088 (n_1699, n2633);
  not g4089 (n_1700, n2643);
  and g4090 (n2644, n_1699, n_1700);
  not g4091 (n_1701, n2644);
  and g4092 (n2645, \asqrt[49] , n_1701);
  and g4096 (n2649, n_1531, n_1530);
  and g4097 (n2650, \asqrt[44] , n2649);
  not g4098 (n_1702, n2650);
  and g4099 (n2651, n_1529, n_1702);
  not g4100 (n_1703, n2648);
  not g4101 (n_1704, n2651);
  and g4102 (n2652, n_1703, n_1704);
  and g4103 (n2653, n_1218, n_1699);
  and g4104 (n2654, n_1700, n2653);
  not g4105 (n_1705, n2652);
  not g4106 (n_1706, n2654);
  and g4107 (n2655, n_1705, n_1706);
  not g4108 (n_1707, n2645);
  not g4109 (n_1708, n2655);
  and g4110 (n2656, n_1707, n_1708);
  not g4111 (n_1709, n2656);
  and g4112 (n2657, \asqrt[50] , n_1709);
  and g4116 (n2661, n_1539, n_1538);
  and g4117 (n2662, \asqrt[44] , n2661);
  not g4118 (n_1710, n2662);
  and g4119 (n2663, n_1537, n_1710);
  not g4120 (n_1711, n2660);
  not g4121 (n_1712, n2663);
  and g4122 (n2664, n_1711, n_1712);
  and g4123 (n2665, n_1082, n_1707);
  and g4124 (n2666, n_1708, n2665);
  not g4125 (n_1713, n2664);
  not g4126 (n_1714, n2666);
  and g4127 (n2667, n_1713, n_1714);
  not g4128 (n_1715, n2657);
  not g4129 (n_1716, n2667);
  and g4130 (n2668, n_1715, n_1716);
  not g4131 (n_1717, n2668);
  and g4132 (n2669, \asqrt[51] , n_1717);
  and g4136 (n2673, n_1547, n_1546);
  and g4137 (n2674, \asqrt[44] , n2673);
  not g4138 (n_1718, n2674);
  and g4139 (n2675, n_1545, n_1718);
  not g4140 (n_1719, n2672);
  not g4141 (n_1720, n2675);
  and g4142 (n2676, n_1719, n_1720);
  and g4143 (n2677, n_954, n_1715);
  and g4144 (n2678, n_1716, n2677);
  not g4145 (n_1721, n2676);
  not g4146 (n_1722, n2678);
  and g4147 (n2679, n_1721, n_1722);
  not g4148 (n_1723, n2669);
  not g4149 (n_1724, n2679);
  and g4150 (n2680, n_1723, n_1724);
  not g4151 (n_1725, n2680);
  and g4152 (n2681, \asqrt[52] , n_1725);
  and g4156 (n2685, n_1555, n_1554);
  and g4157 (n2686, \asqrt[44] , n2685);
  not g4158 (n_1726, n2686);
  and g4159 (n2687, n_1553, n_1726);
  not g4160 (n_1727, n2684);
  not g4161 (n_1728, n2687);
  and g4162 (n2688, n_1727, n_1728);
  and g4163 (n2689, n_834, n_1723);
  and g4164 (n2690, n_1724, n2689);
  not g4165 (n_1729, n2688);
  not g4166 (n_1730, n2690);
  and g4167 (n2691, n_1729, n_1730);
  not g4168 (n_1731, n2681);
  not g4169 (n_1732, n2691);
  and g4170 (n2692, n_1731, n_1732);
  not g4171 (n_1733, n2692);
  and g4172 (n2693, \asqrt[53] , n_1733);
  and g4173 (n2694, n_722, n_1731);
  and g4174 (n2695, n_1732, n2694);
  and g4178 (n2699, n_1563, n_1561);
  and g4179 (n2700, \asqrt[44] , n2699);
  not g4180 (n_1734, n2700);
  and g4181 (n2701, n_1562, n_1734);
  not g4182 (n_1735, n2698);
  not g4183 (n_1736, n2701);
  and g4184 (n2702, n_1735, n_1736);
  not g4185 (n_1737, n2695);
  not g4186 (n_1738, n2702);
  and g4187 (n2703, n_1737, n_1738);
  not g4188 (n_1739, n2693);
  not g4189 (n_1740, n2703);
  and g4190 (n2704, n_1739, n_1740);
  not g4191 (n_1741, n2704);
  and g4192 (n2705, \asqrt[54] , n_1741);
  and g4196 (n2709, n_1571, n_1570);
  and g4197 (n2710, \asqrt[44] , n2709);
  not g4198 (n_1742, n2710);
  and g4199 (n2711, n_1569, n_1742);
  not g4200 (n_1743, n2708);
  not g4201 (n_1744, n2711);
  and g4202 (n2712, n_1743, n_1744);
  and g4203 (n2713, n_618, n_1739);
  and g4204 (n2714, n_1740, n2713);
  not g4205 (n_1745, n2712);
  not g4206 (n_1746, n2714);
  and g4207 (n2715, n_1745, n_1746);
  not g4208 (n_1747, n2705);
  not g4209 (n_1748, n2715);
  and g4210 (n2716, n_1747, n_1748);
  not g4211 (n_1749, n2716);
  and g4212 (n2717, \asqrt[55] , n_1749);
  and g4216 (n2721, n_1579, n_1578);
  and g4217 (n2722, \asqrt[44] , n2721);
  not g4218 (n_1750, n2722);
  and g4219 (n2723, n_1577, n_1750);
  not g4220 (n_1751, n2720);
  not g4221 (n_1752, n2723);
  and g4222 (n2724, n_1751, n_1752);
  and g4223 (n2725, n_522, n_1747);
  and g4224 (n2726, n_1748, n2725);
  not g4225 (n_1753, n2724);
  not g4226 (n_1754, n2726);
  and g4227 (n2727, n_1753, n_1754);
  not g4228 (n_1755, n2717);
  not g4229 (n_1756, n2727);
  and g4230 (n2728, n_1755, n_1756);
  not g4231 (n_1757, n2728);
  and g4232 (n2729, \asqrt[56] , n_1757);
  and g4236 (n2733, n_1587, n_1586);
  and g4237 (n2734, \asqrt[44] , n2733);
  not g4238 (n_1758, n2734);
  and g4239 (n2735, n_1585, n_1758);
  not g4240 (n_1759, n2732);
  not g4241 (n_1760, n2735);
  and g4242 (n2736, n_1759, n_1760);
  and g4243 (n2737, n_434, n_1755);
  and g4244 (n2738, n_1756, n2737);
  not g4245 (n_1761, n2736);
  not g4246 (n_1762, n2738);
  and g4247 (n2739, n_1761, n_1762);
  not g4248 (n_1763, n2729);
  not g4249 (n_1764, n2739);
  and g4250 (n2740, n_1763, n_1764);
  not g4251 (n_1765, n2740);
  and g4252 (n2741, \asqrt[57] , n_1765);
  and g4256 (n2745, n_1595, n_1594);
  and g4257 (n2746, \asqrt[44] , n2745);
  not g4258 (n_1766, n2746);
  and g4259 (n2747, n_1593, n_1766);
  not g4260 (n_1767, n2744);
  not g4261 (n_1768, n2747);
  and g4262 (n2748, n_1767, n_1768);
  and g4263 (n2749, n_354, n_1763);
  and g4264 (n2750, n_1764, n2749);
  not g4265 (n_1769, n2748);
  not g4266 (n_1770, n2750);
  and g4267 (n2751, n_1769, n_1770);
  not g4268 (n_1771, n2741);
  not g4269 (n_1772, n2751);
  and g4270 (n2752, n_1771, n_1772);
  not g4271 (n_1773, n2752);
  and g4272 (n2753, \asqrt[58] , n_1773);
  and g4276 (n2757, n_1603, n_1602);
  and g4277 (n2758, \asqrt[44] , n2757);
  not g4278 (n_1774, n2758);
  and g4279 (n2759, n_1601, n_1774);
  not g4280 (n_1775, n2756);
  not g4281 (n_1776, n2759);
  and g4282 (n2760, n_1775, n_1776);
  and g4283 (n2761, n_282, n_1771);
  and g4284 (n2762, n_1772, n2761);
  not g4285 (n_1777, n2760);
  not g4286 (n_1778, n2762);
  and g4287 (n2763, n_1777, n_1778);
  not g4288 (n_1779, n2753);
  not g4289 (n_1780, n2763);
  and g4290 (n2764, n_1779, n_1780);
  not g4291 (n_1781, n2764);
  and g4292 (n2765, \asqrt[59] , n_1781);
  and g4296 (n2769, n_1611, n_1610);
  and g4297 (n2770, \asqrt[44] , n2769);
  not g4298 (n_1782, n2770);
  and g4299 (n2771, n_1609, n_1782);
  not g4300 (n_1783, n2768);
  not g4301 (n_1784, n2771);
  and g4302 (n2772, n_1783, n_1784);
  and g4303 (n2773, n_218, n_1779);
  and g4304 (n2774, n_1780, n2773);
  not g4305 (n_1785, n2772);
  not g4306 (n_1786, n2774);
  and g4307 (n2775, n_1785, n_1786);
  not g4308 (n_1787, n2765);
  not g4309 (n_1788, n2775);
  and g4310 (n2776, n_1787, n_1788);
  not g4311 (n_1789, n2776);
  and g4312 (n2777, \asqrt[60] , n_1789);
  and g4316 (n2781, n_1619, n_1618);
  and g4317 (n2782, \asqrt[44] , n2781);
  not g4318 (n_1790, n2782);
  and g4319 (n2783, n_1617, n_1790);
  not g4320 (n_1791, n2780);
  not g4321 (n_1792, n2783);
  and g4322 (n2784, n_1791, n_1792);
  and g4323 (n2785, n_162, n_1787);
  and g4324 (n2786, n_1788, n2785);
  not g4325 (n_1793, n2784);
  not g4326 (n_1794, n2786);
  and g4327 (n2787, n_1793, n_1794);
  not g4328 (n_1795, n2777);
  not g4329 (n_1796, n2787);
  and g4330 (n2788, n_1795, n_1796);
  not g4331 (n_1797, n2788);
  and g4332 (n2789, \asqrt[61] , n_1797);
  and g4336 (n2793, n_1627, n_1626);
  and g4337 (n2794, \asqrt[44] , n2793);
  not g4338 (n_1798, n2794);
  and g4339 (n2795, n_1625, n_1798);
  not g4340 (n_1799, n2792);
  not g4341 (n_1800, n2795);
  and g4342 (n2796, n_1799, n_1800);
  and g4343 (n2797, n_115, n_1795);
  and g4344 (n2798, n_1796, n2797);
  not g4345 (n_1801, n2796);
  not g4346 (n_1802, n2798);
  and g4347 (n2799, n_1801, n_1802);
  not g4348 (n_1803, n2789);
  not g4349 (n_1804, n2799);
  and g4350 (n2800, n_1803, n_1804);
  not g4351 (n_1805, n2800);
  and g4352 (n2801, \asqrt[62] , n_1805);
  and g4356 (n2805, n_1635, n_1634);
  and g4357 (n2806, \asqrt[44] , n2805);
  not g4358 (n_1806, n2806);
  and g4359 (n2807, n_1633, n_1806);
  not g4360 (n_1807, n2804);
  not g4361 (n_1808, n2807);
  and g4362 (n2808, n_1807, n_1808);
  and g4363 (n2809, n_76, n_1803);
  and g4364 (n2810, n_1804, n2809);
  not g4365 (n_1809, n2808);
  not g4366 (n_1810, n2810);
  and g4367 (n2811, n_1809, n_1810);
  not g4368 (n_1811, n2801);
  not g4369 (n_1812, n2811);
  and g4370 (n2812, n_1811, n_1812);
  and g4374 (n2816, n_1643, n_1642);
  and g4375 (n2817, \asqrt[44] , n2816);
  not g4376 (n_1813, n2817);
  and g4377 (n2818, n_1641, n_1813);
  not g4378 (n_1814, n2815);
  not g4379 (n_1815, n2818);
  and g4380 (n2819, n_1814, n_1815);
  and g4381 (n2820, n_1650, n_1649);
  and g4382 (n2821, \asqrt[44] , n2820);
  not g4385 (n_1817, n2819);
  not g4387 (n_1818, n2812);
  not g4389 (n_1819, n2824);
  and g4390 (n2825, n_21, n_1819);
  and g4391 (n2826, n_1811, n2819);
  and g4392 (n2827, n_1812, n2826);
  and g4393 (n2828, n_1649, \asqrt[44] );
  not g4394 (n_1820, n2828);
  and g4395 (n2829, n2564, n_1820);
  not g4396 (n_1821, n2820);
  and g4397 (n2830, \asqrt[63] , n_1821);
  not g4398 (n_1822, n2829);
  and g4399 (n2831, n_1822, n2830);
  not g4405 (n_1823, n2831);
  not g4406 (n_1824, n2836);
  not g4408 (n_1825, n2827);
  and g4412 (n2840, \a[86] , \asqrt[43] );
  not g4413 (n_1830, \a[84] );
  not g4414 (n_1831, \a[85] );
  and g4415 (n2841, n_1830, n_1831);
  and g4416 (n2842, n_1662, n2841);
  not g4417 (n_1832, n2840);
  not g4418 (n_1833, n2842);
  and g4419 (n2843, n_1832, n_1833);
  not g4420 (n_1834, n2843);
  and g4421 (n2844, \asqrt[44] , n_1834);
  and g4427 (n2850, n_1662, \asqrt[43] );
  not g4428 (n_1835, n2850);
  and g4429 (n2851, \a[87] , n_1835);
  and g4430 (n2852, n2593, \asqrt[43] );
  not g4431 (n_1836, n2851);
  not g4432 (n_1837, n2852);
  and g4433 (n2853, n_1836, n_1837);
  not g4434 (n_1838, n2849);
  and g4435 (n2854, n_1838, n2853);
  not g4436 (n_1839, n2844);
  not g4437 (n_1840, n2854);
  and g4438 (n2855, n_1839, n_1840);
  not g4439 (n_1841, n2855);
  and g4440 (n2856, \asqrt[45] , n_1841);
  not g4441 (n_1842, \asqrt[45] );
  and g4442 (n2857, n_1842, n_1839);
  and g4443 (n2858, n_1840, n2857);
  not g4447 (n_1843, n2825);
  not g4449 (n_1844, n2862);
  and g4450 (n2863, n_1837, n_1844);
  not g4451 (n_1845, n2863);
  and g4452 (n2864, \a[88] , n_1845);
  and g4453 (n2865, n_1502, n_1844);
  and g4454 (n2866, n_1837, n2865);
  not g4455 (n_1846, n2864);
  not g4456 (n_1847, n2866);
  and g4457 (n2867, n_1846, n_1847);
  not g4458 (n_1848, n2858);
  not g4459 (n_1849, n2867);
  and g4460 (n2868, n_1848, n_1849);
  not g4461 (n_1850, n2856);
  not g4462 (n_1851, n2868);
  and g4463 (n2869, n_1850, n_1851);
  not g4464 (n_1852, n2869);
  and g4465 (n2870, \asqrt[46] , n_1852);
  and g4466 (n2871, n_1671, n_1670);
  not g4467 (n_1853, n2605);
  and g4468 (n2872, n_1853, n2871);
  and g4469 (n2873, \asqrt[43] , n2872);
  and g4470 (n2874, \asqrt[43] , n2871);
  not g4471 (n_1854, n2874);
  and g4472 (n2875, n2605, n_1854);
  not g4473 (n_1855, n2873);
  not g4474 (n_1856, n2875);
  and g4475 (n2876, n_1855, n_1856);
  and g4476 (n2877, n_1674, n_1850);
  and g4477 (n2878, n_1851, n2877);
  not g4478 (n_1857, n2876);
  not g4479 (n_1858, n2878);
  and g4480 (n2879, n_1857, n_1858);
  not g4481 (n_1859, n2870);
  not g4482 (n_1860, n2879);
  and g4483 (n2880, n_1859, n_1860);
  not g4484 (n_1861, n2880);
  and g4485 (n2881, \asqrt[47] , n_1861);
  and g4489 (n2885, n_1682, n_1680);
  and g4490 (n2886, \asqrt[43] , n2885);
  not g4491 (n_1862, n2886);
  and g4492 (n2887, n_1681, n_1862);
  not g4493 (n_1863, n2884);
  not g4494 (n_1864, n2887);
  and g4495 (n2888, n_1863, n_1864);
  and g4496 (n2889, n_1514, n_1859);
  and g4497 (n2890, n_1860, n2889);
  not g4498 (n_1865, n2888);
  not g4499 (n_1866, n2890);
  and g4500 (n2891, n_1865, n_1866);
  not g4501 (n_1867, n2881);
  not g4502 (n_1868, n2891);
  and g4503 (n2892, n_1867, n_1868);
  not g4504 (n_1869, n2892);
  and g4505 (n2893, \asqrt[48] , n_1869);
  and g4509 (n2897, n_1691, n_1690);
  and g4510 (n2898, \asqrt[43] , n2897);
  not g4511 (n_1870, n2898);
  and g4512 (n2899, n_1689, n_1870);
  not g4513 (n_1871, n2896);
  not g4514 (n_1872, n2899);
  and g4515 (n2900, n_1871, n_1872);
  and g4516 (n2901, n_1362, n_1867);
  and g4517 (n2902, n_1868, n2901);
  not g4518 (n_1873, n2900);
  not g4519 (n_1874, n2902);
  and g4520 (n2903, n_1873, n_1874);
  not g4521 (n_1875, n2893);
  not g4522 (n_1876, n2903);
  and g4523 (n2904, n_1875, n_1876);
  not g4524 (n_1877, n2904);
  and g4525 (n2905, \asqrt[49] , n_1877);
  and g4529 (n2909, n_1699, n_1698);
  and g4530 (n2910, \asqrt[43] , n2909);
  not g4531 (n_1878, n2910);
  and g4532 (n2911, n_1697, n_1878);
  not g4533 (n_1879, n2908);
  not g4534 (n_1880, n2911);
  and g4535 (n2912, n_1879, n_1880);
  and g4536 (n2913, n_1218, n_1875);
  and g4537 (n2914, n_1876, n2913);
  not g4538 (n_1881, n2912);
  not g4539 (n_1882, n2914);
  and g4540 (n2915, n_1881, n_1882);
  not g4541 (n_1883, n2905);
  not g4542 (n_1884, n2915);
  and g4543 (n2916, n_1883, n_1884);
  not g4544 (n_1885, n2916);
  and g4545 (n2917, \asqrt[50] , n_1885);
  and g4549 (n2921, n_1707, n_1706);
  and g4550 (n2922, \asqrt[43] , n2921);
  not g4551 (n_1886, n2922);
  and g4552 (n2923, n_1705, n_1886);
  not g4553 (n_1887, n2920);
  not g4554 (n_1888, n2923);
  and g4555 (n2924, n_1887, n_1888);
  and g4556 (n2925, n_1082, n_1883);
  and g4557 (n2926, n_1884, n2925);
  not g4558 (n_1889, n2924);
  not g4559 (n_1890, n2926);
  and g4560 (n2927, n_1889, n_1890);
  not g4561 (n_1891, n2917);
  not g4562 (n_1892, n2927);
  and g4563 (n2928, n_1891, n_1892);
  not g4564 (n_1893, n2928);
  and g4565 (n2929, \asqrt[51] , n_1893);
  and g4569 (n2933, n_1715, n_1714);
  and g4570 (n2934, \asqrt[43] , n2933);
  not g4571 (n_1894, n2934);
  and g4572 (n2935, n_1713, n_1894);
  not g4573 (n_1895, n2932);
  not g4574 (n_1896, n2935);
  and g4575 (n2936, n_1895, n_1896);
  and g4576 (n2937, n_954, n_1891);
  and g4577 (n2938, n_1892, n2937);
  not g4578 (n_1897, n2936);
  not g4579 (n_1898, n2938);
  and g4580 (n2939, n_1897, n_1898);
  not g4581 (n_1899, n2929);
  not g4582 (n_1900, n2939);
  and g4583 (n2940, n_1899, n_1900);
  not g4584 (n_1901, n2940);
  and g4585 (n2941, \asqrt[52] , n_1901);
  and g4589 (n2945, n_1723, n_1722);
  and g4590 (n2946, \asqrt[43] , n2945);
  not g4591 (n_1902, n2946);
  and g4592 (n2947, n_1721, n_1902);
  not g4593 (n_1903, n2944);
  not g4594 (n_1904, n2947);
  and g4595 (n2948, n_1903, n_1904);
  and g4596 (n2949, n_834, n_1899);
  and g4597 (n2950, n_1900, n2949);
  not g4598 (n_1905, n2948);
  not g4599 (n_1906, n2950);
  and g4600 (n2951, n_1905, n_1906);
  not g4601 (n_1907, n2941);
  not g4602 (n_1908, n2951);
  and g4603 (n2952, n_1907, n_1908);
  not g4604 (n_1909, n2952);
  and g4605 (n2953, \asqrt[53] , n_1909);
  and g4609 (n2957, n_1731, n_1730);
  and g4610 (n2958, \asqrt[43] , n2957);
  not g4611 (n_1910, n2958);
  and g4612 (n2959, n_1729, n_1910);
  not g4613 (n_1911, n2956);
  not g4614 (n_1912, n2959);
  and g4615 (n2960, n_1911, n_1912);
  and g4616 (n2961, n_722, n_1907);
  and g4617 (n2962, n_1908, n2961);
  not g4618 (n_1913, n2960);
  not g4619 (n_1914, n2962);
  and g4620 (n2963, n_1913, n_1914);
  not g4621 (n_1915, n2953);
  not g4622 (n_1916, n2963);
  and g4623 (n2964, n_1915, n_1916);
  not g4624 (n_1917, n2964);
  and g4625 (n2965, \asqrt[54] , n_1917);
  and g4626 (n2966, n_618, n_1915);
  and g4627 (n2967, n_1916, n2966);
  and g4631 (n2971, n_1739, n_1737);
  and g4632 (n2972, \asqrt[43] , n2971);
  not g4633 (n_1918, n2972);
  and g4634 (n2973, n_1738, n_1918);
  not g4635 (n_1919, n2970);
  not g4636 (n_1920, n2973);
  and g4637 (n2974, n_1919, n_1920);
  not g4638 (n_1921, n2967);
  not g4639 (n_1922, n2974);
  and g4640 (n2975, n_1921, n_1922);
  not g4641 (n_1923, n2965);
  not g4642 (n_1924, n2975);
  and g4643 (n2976, n_1923, n_1924);
  not g4644 (n_1925, n2976);
  and g4645 (n2977, \asqrt[55] , n_1925);
  and g4649 (n2981, n_1747, n_1746);
  and g4650 (n2982, \asqrt[43] , n2981);
  not g4651 (n_1926, n2982);
  and g4652 (n2983, n_1745, n_1926);
  not g4653 (n_1927, n2980);
  not g4654 (n_1928, n2983);
  and g4655 (n2984, n_1927, n_1928);
  and g4656 (n2985, n_522, n_1923);
  and g4657 (n2986, n_1924, n2985);
  not g4658 (n_1929, n2984);
  not g4659 (n_1930, n2986);
  and g4660 (n2987, n_1929, n_1930);
  not g4661 (n_1931, n2977);
  not g4662 (n_1932, n2987);
  and g4663 (n2988, n_1931, n_1932);
  not g4664 (n_1933, n2988);
  and g4665 (n2989, \asqrt[56] , n_1933);
  and g4669 (n2993, n_1755, n_1754);
  and g4670 (n2994, \asqrt[43] , n2993);
  not g4671 (n_1934, n2994);
  and g4672 (n2995, n_1753, n_1934);
  not g4673 (n_1935, n2992);
  not g4674 (n_1936, n2995);
  and g4675 (n2996, n_1935, n_1936);
  and g4676 (n2997, n_434, n_1931);
  and g4677 (n2998, n_1932, n2997);
  not g4678 (n_1937, n2996);
  not g4679 (n_1938, n2998);
  and g4680 (n2999, n_1937, n_1938);
  not g4681 (n_1939, n2989);
  not g4682 (n_1940, n2999);
  and g4683 (n3000, n_1939, n_1940);
  not g4684 (n_1941, n3000);
  and g4685 (n3001, \asqrt[57] , n_1941);
  and g4689 (n3005, n_1763, n_1762);
  and g4690 (n3006, \asqrt[43] , n3005);
  not g4691 (n_1942, n3006);
  and g4692 (n3007, n_1761, n_1942);
  not g4693 (n_1943, n3004);
  not g4694 (n_1944, n3007);
  and g4695 (n3008, n_1943, n_1944);
  and g4696 (n3009, n_354, n_1939);
  and g4697 (n3010, n_1940, n3009);
  not g4698 (n_1945, n3008);
  not g4699 (n_1946, n3010);
  and g4700 (n3011, n_1945, n_1946);
  not g4701 (n_1947, n3001);
  not g4702 (n_1948, n3011);
  and g4703 (n3012, n_1947, n_1948);
  not g4704 (n_1949, n3012);
  and g4705 (n3013, \asqrt[58] , n_1949);
  and g4709 (n3017, n_1771, n_1770);
  and g4710 (n3018, \asqrt[43] , n3017);
  not g4711 (n_1950, n3018);
  and g4712 (n3019, n_1769, n_1950);
  not g4713 (n_1951, n3016);
  not g4714 (n_1952, n3019);
  and g4715 (n3020, n_1951, n_1952);
  and g4716 (n3021, n_282, n_1947);
  and g4717 (n3022, n_1948, n3021);
  not g4718 (n_1953, n3020);
  not g4719 (n_1954, n3022);
  and g4720 (n3023, n_1953, n_1954);
  not g4721 (n_1955, n3013);
  not g4722 (n_1956, n3023);
  and g4723 (n3024, n_1955, n_1956);
  not g4724 (n_1957, n3024);
  and g4725 (n3025, \asqrt[59] , n_1957);
  and g4729 (n3029, n_1779, n_1778);
  and g4730 (n3030, \asqrt[43] , n3029);
  not g4731 (n_1958, n3030);
  and g4732 (n3031, n_1777, n_1958);
  not g4733 (n_1959, n3028);
  not g4734 (n_1960, n3031);
  and g4735 (n3032, n_1959, n_1960);
  and g4736 (n3033, n_218, n_1955);
  and g4737 (n3034, n_1956, n3033);
  not g4738 (n_1961, n3032);
  not g4739 (n_1962, n3034);
  and g4740 (n3035, n_1961, n_1962);
  not g4741 (n_1963, n3025);
  not g4742 (n_1964, n3035);
  and g4743 (n3036, n_1963, n_1964);
  not g4744 (n_1965, n3036);
  and g4745 (n3037, \asqrt[60] , n_1965);
  and g4749 (n3041, n_1787, n_1786);
  and g4750 (n3042, \asqrt[43] , n3041);
  not g4751 (n_1966, n3042);
  and g4752 (n3043, n_1785, n_1966);
  not g4753 (n_1967, n3040);
  not g4754 (n_1968, n3043);
  and g4755 (n3044, n_1967, n_1968);
  and g4756 (n3045, n_162, n_1963);
  and g4757 (n3046, n_1964, n3045);
  not g4758 (n_1969, n3044);
  not g4759 (n_1970, n3046);
  and g4760 (n3047, n_1969, n_1970);
  not g4761 (n_1971, n3037);
  not g4762 (n_1972, n3047);
  and g4763 (n3048, n_1971, n_1972);
  not g4764 (n_1973, n3048);
  and g4765 (n3049, \asqrt[61] , n_1973);
  and g4769 (n3053, n_1795, n_1794);
  and g4770 (n3054, \asqrt[43] , n3053);
  not g4771 (n_1974, n3054);
  and g4772 (n3055, n_1793, n_1974);
  not g4773 (n_1975, n3052);
  not g4774 (n_1976, n3055);
  and g4775 (n3056, n_1975, n_1976);
  and g4776 (n3057, n_115, n_1971);
  and g4777 (n3058, n_1972, n3057);
  not g4778 (n_1977, n3056);
  not g4779 (n_1978, n3058);
  and g4780 (n3059, n_1977, n_1978);
  not g4781 (n_1979, n3049);
  not g4782 (n_1980, n3059);
  and g4783 (n3060, n_1979, n_1980);
  not g4784 (n_1981, n3060);
  and g4785 (n3061, \asqrt[62] , n_1981);
  and g4789 (n3065, n_1803, n_1802);
  and g4790 (n3066, \asqrt[43] , n3065);
  not g4791 (n_1982, n3066);
  and g4792 (n3067, n_1801, n_1982);
  not g4793 (n_1983, n3064);
  not g4794 (n_1984, n3067);
  and g4795 (n3068, n_1983, n_1984);
  and g4796 (n3069, n_76, n_1979);
  and g4797 (n3070, n_1980, n3069);
  not g4798 (n_1985, n3068);
  not g4799 (n_1986, n3070);
  and g4800 (n3071, n_1985, n_1986);
  not g4801 (n_1987, n3061);
  not g4802 (n_1988, n3071);
  and g4803 (n3072, n_1987, n_1988);
  and g4807 (n3076, n_1811, n_1810);
  and g4808 (n3077, \asqrt[43] , n3076);
  not g4809 (n_1989, n3077);
  and g4810 (n3078, n_1809, n_1989);
  not g4811 (n_1990, n3075);
  not g4812 (n_1991, n3078);
  and g4813 (n3079, n_1990, n_1991);
  and g4814 (n3080, n_1818, n_1817);
  and g4815 (n3081, \asqrt[43] , n3080);
  not g4818 (n_1993, n3079);
  not g4820 (n_1994, n3072);
  not g4822 (n_1995, n3084);
  and g4823 (n3085, n_21, n_1995);
  and g4824 (n3086, n_1987, n3079);
  and g4825 (n3087, n_1988, n3086);
  and g4826 (n3088, n_1817, \asqrt[43] );
  not g4827 (n_1996, n3088);
  and g4828 (n3089, n2812, n_1996);
  not g4829 (n_1997, n3080);
  and g4830 (n3090, \asqrt[63] , n_1997);
  not g4831 (n_1998, n3089);
  and g4832 (n3091, n_1998, n3090);
  not g4838 (n_1999, n3091);
  not g4839 (n_2000, n3096);
  not g4841 (n_2001, n3087);
  and g4845 (n3100, \a[84] , \asqrt[42] );
  not g4846 (n_2006, \a[82] );
  not g4847 (n_2007, \a[83] );
  and g4848 (n3101, n_2006, n_2007);
  and g4849 (n3102, n_1830, n3101);
  not g4850 (n_2008, n3100);
  not g4851 (n_2009, n3102);
  and g4852 (n3103, n_2008, n_2009);
  not g4853 (n_2010, n3103);
  and g4854 (n3104, \asqrt[43] , n_2010);
  and g4860 (n3110, n_1830, \asqrt[42] );
  not g4861 (n_2011, n3110);
  and g4862 (n3111, \a[85] , n_2011);
  and g4863 (n3112, n2841, \asqrt[42] );
  not g4864 (n_2012, n3111);
  not g4865 (n_2013, n3112);
  and g4866 (n3113, n_2012, n_2013);
  not g4867 (n_2014, n3109);
  and g4868 (n3114, n_2014, n3113);
  not g4869 (n_2015, n3104);
  not g4870 (n_2016, n3114);
  and g4871 (n3115, n_2015, n_2016);
  not g4872 (n_2017, n3115);
  and g4873 (n3116, \asqrt[44] , n_2017);
  not g4874 (n_2018, \asqrt[44] );
  and g4875 (n3117, n_2018, n_2015);
  and g4876 (n3118, n_2016, n3117);
  not g4880 (n_2019, n3085);
  not g4882 (n_2020, n3122);
  and g4883 (n3123, n_2013, n_2020);
  not g4884 (n_2021, n3123);
  and g4885 (n3124, \a[86] , n_2021);
  and g4886 (n3125, n_1662, n_2020);
  and g4887 (n3126, n_2013, n3125);
  not g4888 (n_2022, n3124);
  not g4889 (n_2023, n3126);
  and g4890 (n3127, n_2022, n_2023);
  not g4891 (n_2024, n3118);
  not g4892 (n_2025, n3127);
  and g4893 (n3128, n_2024, n_2025);
  not g4894 (n_2026, n3116);
  not g4895 (n_2027, n3128);
  and g4896 (n3129, n_2026, n_2027);
  not g4897 (n_2028, n3129);
  and g4898 (n3130, \asqrt[45] , n_2028);
  and g4899 (n3131, n_1839, n_1838);
  not g4900 (n_2029, n2853);
  and g4901 (n3132, n_2029, n3131);
  and g4902 (n3133, \asqrt[42] , n3132);
  and g4903 (n3134, \asqrt[42] , n3131);
  not g4904 (n_2030, n3134);
  and g4905 (n3135, n2853, n_2030);
  not g4906 (n_2031, n3133);
  not g4907 (n_2032, n3135);
  and g4908 (n3136, n_2031, n_2032);
  and g4909 (n3137, n_1842, n_2026);
  and g4910 (n3138, n_2027, n3137);
  not g4911 (n_2033, n3136);
  not g4912 (n_2034, n3138);
  and g4913 (n3139, n_2033, n_2034);
  not g4914 (n_2035, n3130);
  not g4915 (n_2036, n3139);
  and g4916 (n3140, n_2035, n_2036);
  not g4917 (n_2037, n3140);
  and g4918 (n3141, \asqrt[46] , n_2037);
  and g4922 (n3145, n_1850, n_1848);
  and g4923 (n3146, \asqrt[42] , n3145);
  not g4924 (n_2038, n3146);
  and g4925 (n3147, n_1849, n_2038);
  not g4926 (n_2039, n3144);
  not g4927 (n_2040, n3147);
  and g4928 (n3148, n_2039, n_2040);
  and g4929 (n3149, n_1674, n_2035);
  and g4930 (n3150, n_2036, n3149);
  not g4931 (n_2041, n3148);
  not g4932 (n_2042, n3150);
  and g4933 (n3151, n_2041, n_2042);
  not g4934 (n_2043, n3141);
  not g4935 (n_2044, n3151);
  and g4936 (n3152, n_2043, n_2044);
  not g4937 (n_2045, n3152);
  and g4938 (n3153, \asqrt[47] , n_2045);
  and g4942 (n3157, n_1859, n_1858);
  and g4943 (n3158, \asqrt[42] , n3157);
  not g4944 (n_2046, n3158);
  and g4945 (n3159, n_1857, n_2046);
  not g4946 (n_2047, n3156);
  not g4947 (n_2048, n3159);
  and g4948 (n3160, n_2047, n_2048);
  and g4949 (n3161, n_1514, n_2043);
  and g4950 (n3162, n_2044, n3161);
  not g4951 (n_2049, n3160);
  not g4952 (n_2050, n3162);
  and g4953 (n3163, n_2049, n_2050);
  not g4954 (n_2051, n3153);
  not g4955 (n_2052, n3163);
  and g4956 (n3164, n_2051, n_2052);
  not g4957 (n_2053, n3164);
  and g4958 (n3165, \asqrt[48] , n_2053);
  and g4962 (n3169, n_1867, n_1866);
  and g4963 (n3170, \asqrt[42] , n3169);
  not g4964 (n_2054, n3170);
  and g4965 (n3171, n_1865, n_2054);
  not g4966 (n_2055, n3168);
  not g4967 (n_2056, n3171);
  and g4968 (n3172, n_2055, n_2056);
  and g4969 (n3173, n_1362, n_2051);
  and g4970 (n3174, n_2052, n3173);
  not g4971 (n_2057, n3172);
  not g4972 (n_2058, n3174);
  and g4973 (n3175, n_2057, n_2058);
  not g4974 (n_2059, n3165);
  not g4975 (n_2060, n3175);
  and g4976 (n3176, n_2059, n_2060);
  not g4977 (n_2061, n3176);
  and g4978 (n3177, \asqrt[49] , n_2061);
  and g4982 (n3181, n_1875, n_1874);
  and g4983 (n3182, \asqrt[42] , n3181);
  not g4984 (n_2062, n3182);
  and g4985 (n3183, n_1873, n_2062);
  not g4986 (n_2063, n3180);
  not g4987 (n_2064, n3183);
  and g4988 (n3184, n_2063, n_2064);
  and g4989 (n3185, n_1218, n_2059);
  and g4990 (n3186, n_2060, n3185);
  not g4991 (n_2065, n3184);
  not g4992 (n_2066, n3186);
  and g4993 (n3187, n_2065, n_2066);
  not g4994 (n_2067, n3177);
  not g4995 (n_2068, n3187);
  and g4996 (n3188, n_2067, n_2068);
  not g4997 (n_2069, n3188);
  and g4998 (n3189, \asqrt[50] , n_2069);
  and g5002 (n3193, n_1883, n_1882);
  and g5003 (n3194, \asqrt[42] , n3193);
  not g5004 (n_2070, n3194);
  and g5005 (n3195, n_1881, n_2070);
  not g5006 (n_2071, n3192);
  not g5007 (n_2072, n3195);
  and g5008 (n3196, n_2071, n_2072);
  and g5009 (n3197, n_1082, n_2067);
  and g5010 (n3198, n_2068, n3197);
  not g5011 (n_2073, n3196);
  not g5012 (n_2074, n3198);
  and g5013 (n3199, n_2073, n_2074);
  not g5014 (n_2075, n3189);
  not g5015 (n_2076, n3199);
  and g5016 (n3200, n_2075, n_2076);
  not g5017 (n_2077, n3200);
  and g5018 (n3201, \asqrt[51] , n_2077);
  and g5022 (n3205, n_1891, n_1890);
  and g5023 (n3206, \asqrt[42] , n3205);
  not g5024 (n_2078, n3206);
  and g5025 (n3207, n_1889, n_2078);
  not g5026 (n_2079, n3204);
  not g5027 (n_2080, n3207);
  and g5028 (n3208, n_2079, n_2080);
  and g5029 (n3209, n_954, n_2075);
  and g5030 (n3210, n_2076, n3209);
  not g5031 (n_2081, n3208);
  not g5032 (n_2082, n3210);
  and g5033 (n3211, n_2081, n_2082);
  not g5034 (n_2083, n3201);
  not g5035 (n_2084, n3211);
  and g5036 (n3212, n_2083, n_2084);
  not g5037 (n_2085, n3212);
  and g5038 (n3213, \asqrt[52] , n_2085);
  and g5042 (n3217, n_1899, n_1898);
  and g5043 (n3218, \asqrt[42] , n3217);
  not g5044 (n_2086, n3218);
  and g5045 (n3219, n_1897, n_2086);
  not g5046 (n_2087, n3216);
  not g5047 (n_2088, n3219);
  and g5048 (n3220, n_2087, n_2088);
  and g5049 (n3221, n_834, n_2083);
  and g5050 (n3222, n_2084, n3221);
  not g5051 (n_2089, n3220);
  not g5052 (n_2090, n3222);
  and g5053 (n3223, n_2089, n_2090);
  not g5054 (n_2091, n3213);
  not g5055 (n_2092, n3223);
  and g5056 (n3224, n_2091, n_2092);
  not g5057 (n_2093, n3224);
  and g5058 (n3225, \asqrt[53] , n_2093);
  and g5062 (n3229, n_1907, n_1906);
  and g5063 (n3230, \asqrt[42] , n3229);
  not g5064 (n_2094, n3230);
  and g5065 (n3231, n_1905, n_2094);
  not g5066 (n_2095, n3228);
  not g5067 (n_2096, n3231);
  and g5068 (n3232, n_2095, n_2096);
  and g5069 (n3233, n_722, n_2091);
  and g5070 (n3234, n_2092, n3233);
  not g5071 (n_2097, n3232);
  not g5072 (n_2098, n3234);
  and g5073 (n3235, n_2097, n_2098);
  not g5074 (n_2099, n3225);
  not g5075 (n_2100, n3235);
  and g5076 (n3236, n_2099, n_2100);
  not g5077 (n_2101, n3236);
  and g5078 (n3237, \asqrt[54] , n_2101);
  and g5082 (n3241, n_1915, n_1914);
  and g5083 (n3242, \asqrt[42] , n3241);
  not g5084 (n_2102, n3242);
  and g5085 (n3243, n_1913, n_2102);
  not g5086 (n_2103, n3240);
  not g5087 (n_2104, n3243);
  and g5088 (n3244, n_2103, n_2104);
  and g5089 (n3245, n_618, n_2099);
  and g5090 (n3246, n_2100, n3245);
  not g5091 (n_2105, n3244);
  not g5092 (n_2106, n3246);
  and g5093 (n3247, n_2105, n_2106);
  not g5094 (n_2107, n3237);
  not g5095 (n_2108, n3247);
  and g5096 (n3248, n_2107, n_2108);
  not g5097 (n_2109, n3248);
  and g5098 (n3249, \asqrt[55] , n_2109);
  and g5099 (n3250, n_522, n_2107);
  and g5100 (n3251, n_2108, n3250);
  and g5104 (n3255, n_1923, n_1921);
  and g5105 (n3256, \asqrt[42] , n3255);
  not g5106 (n_2110, n3256);
  and g5107 (n3257, n_1922, n_2110);
  not g5108 (n_2111, n3254);
  not g5109 (n_2112, n3257);
  and g5110 (n3258, n_2111, n_2112);
  not g5111 (n_2113, n3251);
  not g5112 (n_2114, n3258);
  and g5113 (n3259, n_2113, n_2114);
  not g5114 (n_2115, n3249);
  not g5115 (n_2116, n3259);
  and g5116 (n3260, n_2115, n_2116);
  not g5117 (n_2117, n3260);
  and g5118 (n3261, \asqrt[56] , n_2117);
  and g5122 (n3265, n_1931, n_1930);
  and g5123 (n3266, \asqrt[42] , n3265);
  not g5124 (n_2118, n3266);
  and g5125 (n3267, n_1929, n_2118);
  not g5126 (n_2119, n3264);
  not g5127 (n_2120, n3267);
  and g5128 (n3268, n_2119, n_2120);
  and g5129 (n3269, n_434, n_2115);
  and g5130 (n3270, n_2116, n3269);
  not g5131 (n_2121, n3268);
  not g5132 (n_2122, n3270);
  and g5133 (n3271, n_2121, n_2122);
  not g5134 (n_2123, n3261);
  not g5135 (n_2124, n3271);
  and g5136 (n3272, n_2123, n_2124);
  not g5137 (n_2125, n3272);
  and g5138 (n3273, \asqrt[57] , n_2125);
  and g5142 (n3277, n_1939, n_1938);
  and g5143 (n3278, \asqrt[42] , n3277);
  not g5144 (n_2126, n3278);
  and g5145 (n3279, n_1937, n_2126);
  not g5146 (n_2127, n3276);
  not g5147 (n_2128, n3279);
  and g5148 (n3280, n_2127, n_2128);
  and g5149 (n3281, n_354, n_2123);
  and g5150 (n3282, n_2124, n3281);
  not g5151 (n_2129, n3280);
  not g5152 (n_2130, n3282);
  and g5153 (n3283, n_2129, n_2130);
  not g5154 (n_2131, n3273);
  not g5155 (n_2132, n3283);
  and g5156 (n3284, n_2131, n_2132);
  not g5157 (n_2133, n3284);
  and g5158 (n3285, \asqrt[58] , n_2133);
  and g5162 (n3289, n_1947, n_1946);
  and g5163 (n3290, \asqrt[42] , n3289);
  not g5164 (n_2134, n3290);
  and g5165 (n3291, n_1945, n_2134);
  not g5166 (n_2135, n3288);
  not g5167 (n_2136, n3291);
  and g5168 (n3292, n_2135, n_2136);
  and g5169 (n3293, n_282, n_2131);
  and g5170 (n3294, n_2132, n3293);
  not g5171 (n_2137, n3292);
  not g5172 (n_2138, n3294);
  and g5173 (n3295, n_2137, n_2138);
  not g5174 (n_2139, n3285);
  not g5175 (n_2140, n3295);
  and g5176 (n3296, n_2139, n_2140);
  not g5177 (n_2141, n3296);
  and g5178 (n3297, \asqrt[59] , n_2141);
  and g5182 (n3301, n_1955, n_1954);
  and g5183 (n3302, \asqrt[42] , n3301);
  not g5184 (n_2142, n3302);
  and g5185 (n3303, n_1953, n_2142);
  not g5186 (n_2143, n3300);
  not g5187 (n_2144, n3303);
  and g5188 (n3304, n_2143, n_2144);
  and g5189 (n3305, n_218, n_2139);
  and g5190 (n3306, n_2140, n3305);
  not g5191 (n_2145, n3304);
  not g5192 (n_2146, n3306);
  and g5193 (n3307, n_2145, n_2146);
  not g5194 (n_2147, n3297);
  not g5195 (n_2148, n3307);
  and g5196 (n3308, n_2147, n_2148);
  not g5197 (n_2149, n3308);
  and g5198 (n3309, \asqrt[60] , n_2149);
  and g5202 (n3313, n_1963, n_1962);
  and g5203 (n3314, \asqrt[42] , n3313);
  not g5204 (n_2150, n3314);
  and g5205 (n3315, n_1961, n_2150);
  not g5206 (n_2151, n3312);
  not g5207 (n_2152, n3315);
  and g5208 (n3316, n_2151, n_2152);
  and g5209 (n3317, n_162, n_2147);
  and g5210 (n3318, n_2148, n3317);
  not g5211 (n_2153, n3316);
  not g5212 (n_2154, n3318);
  and g5213 (n3319, n_2153, n_2154);
  not g5214 (n_2155, n3309);
  not g5215 (n_2156, n3319);
  and g5216 (n3320, n_2155, n_2156);
  not g5217 (n_2157, n3320);
  and g5218 (n3321, \asqrt[61] , n_2157);
  and g5222 (n3325, n_1971, n_1970);
  and g5223 (n3326, \asqrt[42] , n3325);
  not g5224 (n_2158, n3326);
  and g5225 (n3327, n_1969, n_2158);
  not g5226 (n_2159, n3324);
  not g5227 (n_2160, n3327);
  and g5228 (n3328, n_2159, n_2160);
  and g5229 (n3329, n_115, n_2155);
  and g5230 (n3330, n_2156, n3329);
  not g5231 (n_2161, n3328);
  not g5232 (n_2162, n3330);
  and g5233 (n3331, n_2161, n_2162);
  not g5234 (n_2163, n3321);
  not g5235 (n_2164, n3331);
  and g5236 (n3332, n_2163, n_2164);
  not g5237 (n_2165, n3332);
  and g5238 (n3333, \asqrt[62] , n_2165);
  and g5242 (n3337, n_1979, n_1978);
  and g5243 (n3338, \asqrt[42] , n3337);
  not g5244 (n_2166, n3338);
  and g5245 (n3339, n_1977, n_2166);
  not g5246 (n_2167, n3336);
  not g5247 (n_2168, n3339);
  and g5248 (n3340, n_2167, n_2168);
  and g5249 (n3341, n_76, n_2163);
  and g5250 (n3342, n_2164, n3341);
  not g5251 (n_2169, n3340);
  not g5252 (n_2170, n3342);
  and g5253 (n3343, n_2169, n_2170);
  not g5254 (n_2171, n3333);
  not g5255 (n_2172, n3343);
  and g5256 (n3344, n_2171, n_2172);
  and g5260 (n3348, n_1987, n_1986);
  and g5261 (n3349, \asqrt[42] , n3348);
  not g5262 (n_2173, n3349);
  and g5263 (n3350, n_1985, n_2173);
  not g5264 (n_2174, n3347);
  not g5265 (n_2175, n3350);
  and g5266 (n3351, n_2174, n_2175);
  and g5267 (n3352, n_1994, n_1993);
  and g5268 (n3353, \asqrt[42] , n3352);
  not g5271 (n_2177, n3351);
  not g5273 (n_2178, n3344);
  not g5275 (n_2179, n3356);
  and g5276 (n3357, n_21, n_2179);
  and g5277 (n3358, n_2171, n3351);
  and g5278 (n3359, n_2172, n3358);
  and g5279 (n3360, n_1993, \asqrt[42] );
  not g5280 (n_2180, n3360);
  and g5281 (n3361, n3072, n_2180);
  not g5282 (n_2181, n3352);
  and g5283 (n3362, \asqrt[63] , n_2181);
  not g5284 (n_2182, n3361);
  and g5285 (n3363, n_2182, n3362);
  not g5291 (n_2183, n3363);
  not g5292 (n_2184, n3368);
  not g5294 (n_2185, n3359);
  and g5298 (n3372, \a[82] , \asqrt[41] );
  not g5299 (n_2190, \a[80] );
  not g5300 (n_2191, \a[81] );
  and g5301 (n3373, n_2190, n_2191);
  and g5302 (n3374, n_2006, n3373);
  not g5303 (n_2192, n3372);
  not g5304 (n_2193, n3374);
  and g5305 (n3375, n_2192, n_2193);
  not g5306 (n_2194, n3375);
  and g5307 (n3376, \asqrt[42] , n_2194);
  and g5313 (n3382, n_2006, \asqrt[41] );
  not g5314 (n_2195, n3382);
  and g5315 (n3383, \a[83] , n_2195);
  and g5316 (n3384, n3101, \asqrt[41] );
  not g5317 (n_2196, n3383);
  not g5318 (n_2197, n3384);
  and g5319 (n3385, n_2196, n_2197);
  not g5320 (n_2198, n3381);
  and g5321 (n3386, n_2198, n3385);
  not g5322 (n_2199, n3376);
  not g5323 (n_2200, n3386);
  and g5324 (n3387, n_2199, n_2200);
  not g5325 (n_2201, n3387);
  and g5326 (n3388, \asqrt[43] , n_2201);
  not g5327 (n_2202, \asqrt[43] );
  and g5328 (n3389, n_2202, n_2199);
  and g5329 (n3390, n_2200, n3389);
  not g5333 (n_2203, n3357);
  not g5335 (n_2204, n3394);
  and g5336 (n3395, n_2197, n_2204);
  not g5337 (n_2205, n3395);
  and g5338 (n3396, \a[84] , n_2205);
  and g5339 (n3397, n_1830, n_2204);
  and g5340 (n3398, n_2197, n3397);
  not g5341 (n_2206, n3396);
  not g5342 (n_2207, n3398);
  and g5343 (n3399, n_2206, n_2207);
  not g5344 (n_2208, n3390);
  not g5345 (n_2209, n3399);
  and g5346 (n3400, n_2208, n_2209);
  not g5347 (n_2210, n3388);
  not g5348 (n_2211, n3400);
  and g5349 (n3401, n_2210, n_2211);
  not g5350 (n_2212, n3401);
  and g5351 (n3402, \asqrt[44] , n_2212);
  and g5352 (n3403, n_2015, n_2014);
  not g5353 (n_2213, n3113);
  and g5354 (n3404, n_2213, n3403);
  and g5355 (n3405, \asqrt[41] , n3404);
  and g5356 (n3406, \asqrt[41] , n3403);
  not g5357 (n_2214, n3406);
  and g5358 (n3407, n3113, n_2214);
  not g5359 (n_2215, n3405);
  not g5360 (n_2216, n3407);
  and g5361 (n3408, n_2215, n_2216);
  and g5362 (n3409, n_2018, n_2210);
  and g5363 (n3410, n_2211, n3409);
  not g5364 (n_2217, n3408);
  not g5365 (n_2218, n3410);
  and g5366 (n3411, n_2217, n_2218);
  not g5367 (n_2219, n3402);
  not g5368 (n_2220, n3411);
  and g5369 (n3412, n_2219, n_2220);
  not g5370 (n_2221, n3412);
  and g5371 (n3413, \asqrt[45] , n_2221);
  and g5375 (n3417, n_2026, n_2024);
  and g5376 (n3418, \asqrt[41] , n3417);
  not g5377 (n_2222, n3418);
  and g5378 (n3419, n_2025, n_2222);
  not g5379 (n_2223, n3416);
  not g5380 (n_2224, n3419);
  and g5381 (n3420, n_2223, n_2224);
  and g5382 (n3421, n_1842, n_2219);
  and g5383 (n3422, n_2220, n3421);
  not g5384 (n_2225, n3420);
  not g5385 (n_2226, n3422);
  and g5386 (n3423, n_2225, n_2226);
  not g5387 (n_2227, n3413);
  not g5388 (n_2228, n3423);
  and g5389 (n3424, n_2227, n_2228);
  not g5390 (n_2229, n3424);
  and g5391 (n3425, \asqrt[46] , n_2229);
  and g5395 (n3429, n_2035, n_2034);
  and g5396 (n3430, \asqrt[41] , n3429);
  not g5397 (n_2230, n3430);
  and g5398 (n3431, n_2033, n_2230);
  not g5399 (n_2231, n3428);
  not g5400 (n_2232, n3431);
  and g5401 (n3432, n_2231, n_2232);
  and g5402 (n3433, n_1674, n_2227);
  and g5403 (n3434, n_2228, n3433);
  not g5404 (n_2233, n3432);
  not g5405 (n_2234, n3434);
  and g5406 (n3435, n_2233, n_2234);
  not g5407 (n_2235, n3425);
  not g5408 (n_2236, n3435);
  and g5409 (n3436, n_2235, n_2236);
  not g5410 (n_2237, n3436);
  and g5411 (n3437, \asqrt[47] , n_2237);
  and g5415 (n3441, n_2043, n_2042);
  and g5416 (n3442, \asqrt[41] , n3441);
  not g5417 (n_2238, n3442);
  and g5418 (n3443, n_2041, n_2238);
  not g5419 (n_2239, n3440);
  not g5420 (n_2240, n3443);
  and g5421 (n3444, n_2239, n_2240);
  and g5422 (n3445, n_1514, n_2235);
  and g5423 (n3446, n_2236, n3445);
  not g5424 (n_2241, n3444);
  not g5425 (n_2242, n3446);
  and g5426 (n3447, n_2241, n_2242);
  not g5427 (n_2243, n3437);
  not g5428 (n_2244, n3447);
  and g5429 (n3448, n_2243, n_2244);
  not g5430 (n_2245, n3448);
  and g5431 (n3449, \asqrt[48] , n_2245);
  and g5435 (n3453, n_2051, n_2050);
  and g5436 (n3454, \asqrt[41] , n3453);
  not g5437 (n_2246, n3454);
  and g5438 (n3455, n_2049, n_2246);
  not g5439 (n_2247, n3452);
  not g5440 (n_2248, n3455);
  and g5441 (n3456, n_2247, n_2248);
  and g5442 (n3457, n_1362, n_2243);
  and g5443 (n3458, n_2244, n3457);
  not g5444 (n_2249, n3456);
  not g5445 (n_2250, n3458);
  and g5446 (n3459, n_2249, n_2250);
  not g5447 (n_2251, n3449);
  not g5448 (n_2252, n3459);
  and g5449 (n3460, n_2251, n_2252);
  not g5450 (n_2253, n3460);
  and g5451 (n3461, \asqrt[49] , n_2253);
  and g5455 (n3465, n_2059, n_2058);
  and g5456 (n3466, \asqrt[41] , n3465);
  not g5457 (n_2254, n3466);
  and g5458 (n3467, n_2057, n_2254);
  not g5459 (n_2255, n3464);
  not g5460 (n_2256, n3467);
  and g5461 (n3468, n_2255, n_2256);
  and g5462 (n3469, n_1218, n_2251);
  and g5463 (n3470, n_2252, n3469);
  not g5464 (n_2257, n3468);
  not g5465 (n_2258, n3470);
  and g5466 (n3471, n_2257, n_2258);
  not g5467 (n_2259, n3461);
  not g5468 (n_2260, n3471);
  and g5469 (n3472, n_2259, n_2260);
  not g5470 (n_2261, n3472);
  and g5471 (n3473, \asqrt[50] , n_2261);
  and g5475 (n3477, n_2067, n_2066);
  and g5476 (n3478, \asqrt[41] , n3477);
  not g5477 (n_2262, n3478);
  and g5478 (n3479, n_2065, n_2262);
  not g5479 (n_2263, n3476);
  not g5480 (n_2264, n3479);
  and g5481 (n3480, n_2263, n_2264);
  and g5482 (n3481, n_1082, n_2259);
  and g5483 (n3482, n_2260, n3481);
  not g5484 (n_2265, n3480);
  not g5485 (n_2266, n3482);
  and g5486 (n3483, n_2265, n_2266);
  not g5487 (n_2267, n3473);
  not g5488 (n_2268, n3483);
  and g5489 (n3484, n_2267, n_2268);
  not g5490 (n_2269, n3484);
  and g5491 (n3485, \asqrt[51] , n_2269);
  and g5495 (n3489, n_2075, n_2074);
  and g5496 (n3490, \asqrt[41] , n3489);
  not g5497 (n_2270, n3490);
  and g5498 (n3491, n_2073, n_2270);
  not g5499 (n_2271, n3488);
  not g5500 (n_2272, n3491);
  and g5501 (n3492, n_2271, n_2272);
  and g5502 (n3493, n_954, n_2267);
  and g5503 (n3494, n_2268, n3493);
  not g5504 (n_2273, n3492);
  not g5505 (n_2274, n3494);
  and g5506 (n3495, n_2273, n_2274);
  not g5507 (n_2275, n3485);
  not g5508 (n_2276, n3495);
  and g5509 (n3496, n_2275, n_2276);
  not g5510 (n_2277, n3496);
  and g5511 (n3497, \asqrt[52] , n_2277);
  and g5515 (n3501, n_2083, n_2082);
  and g5516 (n3502, \asqrt[41] , n3501);
  not g5517 (n_2278, n3502);
  and g5518 (n3503, n_2081, n_2278);
  not g5519 (n_2279, n3500);
  not g5520 (n_2280, n3503);
  and g5521 (n3504, n_2279, n_2280);
  and g5522 (n3505, n_834, n_2275);
  and g5523 (n3506, n_2276, n3505);
  not g5524 (n_2281, n3504);
  not g5525 (n_2282, n3506);
  and g5526 (n3507, n_2281, n_2282);
  not g5527 (n_2283, n3497);
  not g5528 (n_2284, n3507);
  and g5529 (n3508, n_2283, n_2284);
  not g5530 (n_2285, n3508);
  and g5531 (n3509, \asqrt[53] , n_2285);
  and g5535 (n3513, n_2091, n_2090);
  and g5536 (n3514, \asqrt[41] , n3513);
  not g5537 (n_2286, n3514);
  and g5538 (n3515, n_2089, n_2286);
  not g5539 (n_2287, n3512);
  not g5540 (n_2288, n3515);
  and g5541 (n3516, n_2287, n_2288);
  and g5542 (n3517, n_722, n_2283);
  and g5543 (n3518, n_2284, n3517);
  not g5544 (n_2289, n3516);
  not g5545 (n_2290, n3518);
  and g5546 (n3519, n_2289, n_2290);
  not g5547 (n_2291, n3509);
  not g5548 (n_2292, n3519);
  and g5549 (n3520, n_2291, n_2292);
  not g5550 (n_2293, n3520);
  and g5551 (n3521, \asqrt[54] , n_2293);
  and g5555 (n3525, n_2099, n_2098);
  and g5556 (n3526, \asqrt[41] , n3525);
  not g5557 (n_2294, n3526);
  and g5558 (n3527, n_2097, n_2294);
  not g5559 (n_2295, n3524);
  not g5560 (n_2296, n3527);
  and g5561 (n3528, n_2295, n_2296);
  and g5562 (n3529, n_618, n_2291);
  and g5563 (n3530, n_2292, n3529);
  not g5564 (n_2297, n3528);
  not g5565 (n_2298, n3530);
  and g5566 (n3531, n_2297, n_2298);
  not g5567 (n_2299, n3521);
  not g5568 (n_2300, n3531);
  and g5569 (n3532, n_2299, n_2300);
  not g5570 (n_2301, n3532);
  and g5571 (n3533, \asqrt[55] , n_2301);
  and g5575 (n3537, n_2107, n_2106);
  and g5576 (n3538, \asqrt[41] , n3537);
  not g5577 (n_2302, n3538);
  and g5578 (n3539, n_2105, n_2302);
  not g5579 (n_2303, n3536);
  not g5580 (n_2304, n3539);
  and g5581 (n3540, n_2303, n_2304);
  and g5582 (n3541, n_522, n_2299);
  and g5583 (n3542, n_2300, n3541);
  not g5584 (n_2305, n3540);
  not g5585 (n_2306, n3542);
  and g5586 (n3543, n_2305, n_2306);
  not g5587 (n_2307, n3533);
  not g5588 (n_2308, n3543);
  and g5589 (n3544, n_2307, n_2308);
  not g5590 (n_2309, n3544);
  and g5591 (n3545, \asqrt[56] , n_2309);
  and g5592 (n3546, n_434, n_2307);
  and g5593 (n3547, n_2308, n3546);
  and g5597 (n3551, n_2115, n_2113);
  and g5598 (n3552, \asqrt[41] , n3551);
  not g5599 (n_2310, n3552);
  and g5600 (n3553, n_2114, n_2310);
  not g5601 (n_2311, n3550);
  not g5602 (n_2312, n3553);
  and g5603 (n3554, n_2311, n_2312);
  not g5604 (n_2313, n3547);
  not g5605 (n_2314, n3554);
  and g5606 (n3555, n_2313, n_2314);
  not g5607 (n_2315, n3545);
  not g5608 (n_2316, n3555);
  and g5609 (n3556, n_2315, n_2316);
  not g5610 (n_2317, n3556);
  and g5611 (n3557, \asqrt[57] , n_2317);
  and g5615 (n3561, n_2123, n_2122);
  and g5616 (n3562, \asqrt[41] , n3561);
  not g5617 (n_2318, n3562);
  and g5618 (n3563, n_2121, n_2318);
  not g5619 (n_2319, n3560);
  not g5620 (n_2320, n3563);
  and g5621 (n3564, n_2319, n_2320);
  and g5622 (n3565, n_354, n_2315);
  and g5623 (n3566, n_2316, n3565);
  not g5624 (n_2321, n3564);
  not g5625 (n_2322, n3566);
  and g5626 (n3567, n_2321, n_2322);
  not g5627 (n_2323, n3557);
  not g5628 (n_2324, n3567);
  and g5629 (n3568, n_2323, n_2324);
  not g5630 (n_2325, n3568);
  and g5631 (n3569, \asqrt[58] , n_2325);
  and g5635 (n3573, n_2131, n_2130);
  and g5636 (n3574, \asqrt[41] , n3573);
  not g5637 (n_2326, n3574);
  and g5638 (n3575, n_2129, n_2326);
  not g5639 (n_2327, n3572);
  not g5640 (n_2328, n3575);
  and g5641 (n3576, n_2327, n_2328);
  and g5642 (n3577, n_282, n_2323);
  and g5643 (n3578, n_2324, n3577);
  not g5644 (n_2329, n3576);
  not g5645 (n_2330, n3578);
  and g5646 (n3579, n_2329, n_2330);
  not g5647 (n_2331, n3569);
  not g5648 (n_2332, n3579);
  and g5649 (n3580, n_2331, n_2332);
  not g5650 (n_2333, n3580);
  and g5651 (n3581, \asqrt[59] , n_2333);
  and g5655 (n3585, n_2139, n_2138);
  and g5656 (n3586, \asqrt[41] , n3585);
  not g5657 (n_2334, n3586);
  and g5658 (n3587, n_2137, n_2334);
  not g5659 (n_2335, n3584);
  not g5660 (n_2336, n3587);
  and g5661 (n3588, n_2335, n_2336);
  and g5662 (n3589, n_218, n_2331);
  and g5663 (n3590, n_2332, n3589);
  not g5664 (n_2337, n3588);
  not g5665 (n_2338, n3590);
  and g5666 (n3591, n_2337, n_2338);
  not g5667 (n_2339, n3581);
  not g5668 (n_2340, n3591);
  and g5669 (n3592, n_2339, n_2340);
  not g5670 (n_2341, n3592);
  and g5671 (n3593, \asqrt[60] , n_2341);
  and g5675 (n3597, n_2147, n_2146);
  and g5676 (n3598, \asqrt[41] , n3597);
  not g5677 (n_2342, n3598);
  and g5678 (n3599, n_2145, n_2342);
  not g5679 (n_2343, n3596);
  not g5680 (n_2344, n3599);
  and g5681 (n3600, n_2343, n_2344);
  and g5682 (n3601, n_162, n_2339);
  and g5683 (n3602, n_2340, n3601);
  not g5684 (n_2345, n3600);
  not g5685 (n_2346, n3602);
  and g5686 (n3603, n_2345, n_2346);
  not g5687 (n_2347, n3593);
  not g5688 (n_2348, n3603);
  and g5689 (n3604, n_2347, n_2348);
  not g5690 (n_2349, n3604);
  and g5691 (n3605, \asqrt[61] , n_2349);
  and g5695 (n3609, n_2155, n_2154);
  and g5696 (n3610, \asqrt[41] , n3609);
  not g5697 (n_2350, n3610);
  and g5698 (n3611, n_2153, n_2350);
  not g5699 (n_2351, n3608);
  not g5700 (n_2352, n3611);
  and g5701 (n3612, n_2351, n_2352);
  and g5702 (n3613, n_115, n_2347);
  and g5703 (n3614, n_2348, n3613);
  not g5704 (n_2353, n3612);
  not g5705 (n_2354, n3614);
  and g5706 (n3615, n_2353, n_2354);
  not g5707 (n_2355, n3605);
  not g5708 (n_2356, n3615);
  and g5709 (n3616, n_2355, n_2356);
  not g5710 (n_2357, n3616);
  and g5711 (n3617, \asqrt[62] , n_2357);
  and g5715 (n3621, n_2163, n_2162);
  and g5716 (n3622, \asqrt[41] , n3621);
  not g5717 (n_2358, n3622);
  and g5718 (n3623, n_2161, n_2358);
  not g5719 (n_2359, n3620);
  not g5720 (n_2360, n3623);
  and g5721 (n3624, n_2359, n_2360);
  and g5722 (n3625, n_76, n_2355);
  and g5723 (n3626, n_2356, n3625);
  not g5724 (n_2361, n3624);
  not g5725 (n_2362, n3626);
  and g5726 (n3627, n_2361, n_2362);
  not g5727 (n_2363, n3617);
  not g5728 (n_2364, n3627);
  and g5729 (n3628, n_2363, n_2364);
  and g5733 (n3632, n_2171, n_2170);
  and g5734 (n3633, \asqrt[41] , n3632);
  not g5735 (n_2365, n3633);
  and g5736 (n3634, n_2169, n_2365);
  not g5737 (n_2366, n3631);
  not g5738 (n_2367, n3634);
  and g5739 (n3635, n_2366, n_2367);
  and g5740 (n3636, n_2178, n_2177);
  and g5741 (n3637, \asqrt[41] , n3636);
  not g5744 (n_2369, n3635);
  not g5746 (n_2370, n3628);
  not g5748 (n_2371, n3640);
  and g5749 (n3641, n_21, n_2371);
  and g5750 (n3642, n_2363, n3635);
  and g5751 (n3643, n_2364, n3642);
  and g5752 (n3644, n_2177, \asqrt[41] );
  not g5753 (n_2372, n3644);
  and g5754 (n3645, n3344, n_2372);
  not g5755 (n_2373, n3636);
  and g5756 (n3646, \asqrt[63] , n_2373);
  not g5757 (n_2374, n3645);
  and g5758 (n3647, n_2374, n3646);
  not g5764 (n_2375, n3647);
  not g5765 (n_2376, n3652);
  not g5767 (n_2377, n3643);
  and g5771 (n3656, \a[80] , \asqrt[40] );
  not g5772 (n_2382, \a[78] );
  not g5773 (n_2383, \a[79] );
  and g5774 (n3657, n_2382, n_2383);
  and g5775 (n3658, n_2190, n3657);
  not g5776 (n_2384, n3656);
  not g5777 (n_2385, n3658);
  and g5778 (n3659, n_2384, n_2385);
  not g5779 (n_2386, n3659);
  and g5780 (n3660, \asqrt[41] , n_2386);
  and g5786 (n3666, n_2190, \asqrt[40] );
  not g5787 (n_2387, n3666);
  and g5788 (n3667, \a[81] , n_2387);
  and g5789 (n3668, n3373, \asqrt[40] );
  not g5790 (n_2388, n3667);
  not g5791 (n_2389, n3668);
  and g5792 (n3669, n_2388, n_2389);
  not g5793 (n_2390, n3665);
  and g5794 (n3670, n_2390, n3669);
  not g5795 (n_2391, n3660);
  not g5796 (n_2392, n3670);
  and g5797 (n3671, n_2391, n_2392);
  not g5798 (n_2393, n3671);
  and g5799 (n3672, \asqrt[42] , n_2393);
  not g5800 (n_2394, \asqrt[42] );
  and g5801 (n3673, n_2394, n_2391);
  and g5802 (n3674, n_2392, n3673);
  not g5806 (n_2395, n3641);
  not g5808 (n_2396, n3678);
  and g5809 (n3679, n_2389, n_2396);
  not g5810 (n_2397, n3679);
  and g5811 (n3680, \a[82] , n_2397);
  and g5812 (n3681, n_2006, n_2396);
  and g5813 (n3682, n_2389, n3681);
  not g5814 (n_2398, n3680);
  not g5815 (n_2399, n3682);
  and g5816 (n3683, n_2398, n_2399);
  not g5817 (n_2400, n3674);
  not g5818 (n_2401, n3683);
  and g5819 (n3684, n_2400, n_2401);
  not g5820 (n_2402, n3672);
  not g5821 (n_2403, n3684);
  and g5822 (n3685, n_2402, n_2403);
  not g5823 (n_2404, n3685);
  and g5824 (n3686, \asqrt[43] , n_2404);
  and g5825 (n3687, n_2199, n_2198);
  not g5826 (n_2405, n3385);
  and g5827 (n3688, n_2405, n3687);
  and g5828 (n3689, \asqrt[40] , n3688);
  and g5829 (n3690, \asqrt[40] , n3687);
  not g5830 (n_2406, n3690);
  and g5831 (n3691, n3385, n_2406);
  not g5832 (n_2407, n3689);
  not g5833 (n_2408, n3691);
  and g5834 (n3692, n_2407, n_2408);
  and g5835 (n3693, n_2202, n_2402);
  and g5836 (n3694, n_2403, n3693);
  not g5837 (n_2409, n3692);
  not g5838 (n_2410, n3694);
  and g5839 (n3695, n_2409, n_2410);
  not g5840 (n_2411, n3686);
  not g5841 (n_2412, n3695);
  and g5842 (n3696, n_2411, n_2412);
  not g5843 (n_2413, n3696);
  and g5844 (n3697, \asqrt[44] , n_2413);
  and g5848 (n3701, n_2210, n_2208);
  and g5849 (n3702, \asqrt[40] , n3701);
  not g5850 (n_2414, n3702);
  and g5851 (n3703, n_2209, n_2414);
  not g5852 (n_2415, n3700);
  not g5853 (n_2416, n3703);
  and g5854 (n3704, n_2415, n_2416);
  and g5855 (n3705, n_2018, n_2411);
  and g5856 (n3706, n_2412, n3705);
  not g5857 (n_2417, n3704);
  not g5858 (n_2418, n3706);
  and g5859 (n3707, n_2417, n_2418);
  not g5860 (n_2419, n3697);
  not g5861 (n_2420, n3707);
  and g5862 (n3708, n_2419, n_2420);
  not g5863 (n_2421, n3708);
  and g5864 (n3709, \asqrt[45] , n_2421);
  and g5868 (n3713, n_2219, n_2218);
  and g5869 (n3714, \asqrt[40] , n3713);
  not g5870 (n_2422, n3714);
  and g5871 (n3715, n_2217, n_2422);
  not g5872 (n_2423, n3712);
  not g5873 (n_2424, n3715);
  and g5874 (n3716, n_2423, n_2424);
  and g5875 (n3717, n_1842, n_2419);
  and g5876 (n3718, n_2420, n3717);
  not g5877 (n_2425, n3716);
  not g5878 (n_2426, n3718);
  and g5879 (n3719, n_2425, n_2426);
  not g5880 (n_2427, n3709);
  not g5881 (n_2428, n3719);
  and g5882 (n3720, n_2427, n_2428);
  not g5883 (n_2429, n3720);
  and g5884 (n3721, \asqrt[46] , n_2429);
  and g5888 (n3725, n_2227, n_2226);
  and g5889 (n3726, \asqrt[40] , n3725);
  not g5890 (n_2430, n3726);
  and g5891 (n3727, n_2225, n_2430);
  not g5892 (n_2431, n3724);
  not g5893 (n_2432, n3727);
  and g5894 (n3728, n_2431, n_2432);
  and g5895 (n3729, n_1674, n_2427);
  and g5896 (n3730, n_2428, n3729);
  not g5897 (n_2433, n3728);
  not g5898 (n_2434, n3730);
  and g5899 (n3731, n_2433, n_2434);
  not g5900 (n_2435, n3721);
  not g5901 (n_2436, n3731);
  and g5902 (n3732, n_2435, n_2436);
  not g5903 (n_2437, n3732);
  and g5904 (n3733, \asqrt[47] , n_2437);
  and g5908 (n3737, n_2235, n_2234);
  and g5909 (n3738, \asqrt[40] , n3737);
  not g5910 (n_2438, n3738);
  and g5911 (n3739, n_2233, n_2438);
  not g5912 (n_2439, n3736);
  not g5913 (n_2440, n3739);
  and g5914 (n3740, n_2439, n_2440);
  and g5915 (n3741, n_1514, n_2435);
  and g5916 (n3742, n_2436, n3741);
  not g5917 (n_2441, n3740);
  not g5918 (n_2442, n3742);
  and g5919 (n3743, n_2441, n_2442);
  not g5920 (n_2443, n3733);
  not g5921 (n_2444, n3743);
  and g5922 (n3744, n_2443, n_2444);
  not g5923 (n_2445, n3744);
  and g5924 (n3745, \asqrt[48] , n_2445);
  and g5928 (n3749, n_2243, n_2242);
  and g5929 (n3750, \asqrt[40] , n3749);
  not g5930 (n_2446, n3750);
  and g5931 (n3751, n_2241, n_2446);
  not g5932 (n_2447, n3748);
  not g5933 (n_2448, n3751);
  and g5934 (n3752, n_2447, n_2448);
  and g5935 (n3753, n_1362, n_2443);
  and g5936 (n3754, n_2444, n3753);
  not g5937 (n_2449, n3752);
  not g5938 (n_2450, n3754);
  and g5939 (n3755, n_2449, n_2450);
  not g5940 (n_2451, n3745);
  not g5941 (n_2452, n3755);
  and g5942 (n3756, n_2451, n_2452);
  not g5943 (n_2453, n3756);
  and g5944 (n3757, \asqrt[49] , n_2453);
  and g5948 (n3761, n_2251, n_2250);
  and g5949 (n3762, \asqrt[40] , n3761);
  not g5950 (n_2454, n3762);
  and g5951 (n3763, n_2249, n_2454);
  not g5952 (n_2455, n3760);
  not g5953 (n_2456, n3763);
  and g5954 (n3764, n_2455, n_2456);
  and g5955 (n3765, n_1218, n_2451);
  and g5956 (n3766, n_2452, n3765);
  not g5957 (n_2457, n3764);
  not g5958 (n_2458, n3766);
  and g5959 (n3767, n_2457, n_2458);
  not g5960 (n_2459, n3757);
  not g5961 (n_2460, n3767);
  and g5962 (n3768, n_2459, n_2460);
  not g5963 (n_2461, n3768);
  and g5964 (n3769, \asqrt[50] , n_2461);
  and g5968 (n3773, n_2259, n_2258);
  and g5969 (n3774, \asqrt[40] , n3773);
  not g5970 (n_2462, n3774);
  and g5971 (n3775, n_2257, n_2462);
  not g5972 (n_2463, n3772);
  not g5973 (n_2464, n3775);
  and g5974 (n3776, n_2463, n_2464);
  and g5975 (n3777, n_1082, n_2459);
  and g5976 (n3778, n_2460, n3777);
  not g5977 (n_2465, n3776);
  not g5978 (n_2466, n3778);
  and g5979 (n3779, n_2465, n_2466);
  not g5980 (n_2467, n3769);
  not g5981 (n_2468, n3779);
  and g5982 (n3780, n_2467, n_2468);
  not g5983 (n_2469, n3780);
  and g5984 (n3781, \asqrt[51] , n_2469);
  and g5988 (n3785, n_2267, n_2266);
  and g5989 (n3786, \asqrt[40] , n3785);
  not g5990 (n_2470, n3786);
  and g5991 (n3787, n_2265, n_2470);
  not g5992 (n_2471, n3784);
  not g5993 (n_2472, n3787);
  and g5994 (n3788, n_2471, n_2472);
  and g5995 (n3789, n_954, n_2467);
  and g5996 (n3790, n_2468, n3789);
  not g5997 (n_2473, n3788);
  not g5998 (n_2474, n3790);
  and g5999 (n3791, n_2473, n_2474);
  not g6000 (n_2475, n3781);
  not g6001 (n_2476, n3791);
  and g6002 (n3792, n_2475, n_2476);
  not g6003 (n_2477, n3792);
  and g6004 (n3793, \asqrt[52] , n_2477);
  and g6008 (n3797, n_2275, n_2274);
  and g6009 (n3798, \asqrt[40] , n3797);
  not g6010 (n_2478, n3798);
  and g6011 (n3799, n_2273, n_2478);
  not g6012 (n_2479, n3796);
  not g6013 (n_2480, n3799);
  and g6014 (n3800, n_2479, n_2480);
  and g6015 (n3801, n_834, n_2475);
  and g6016 (n3802, n_2476, n3801);
  not g6017 (n_2481, n3800);
  not g6018 (n_2482, n3802);
  and g6019 (n3803, n_2481, n_2482);
  not g6020 (n_2483, n3793);
  not g6021 (n_2484, n3803);
  and g6022 (n3804, n_2483, n_2484);
  not g6023 (n_2485, n3804);
  and g6024 (n3805, \asqrt[53] , n_2485);
  and g6028 (n3809, n_2283, n_2282);
  and g6029 (n3810, \asqrt[40] , n3809);
  not g6030 (n_2486, n3810);
  and g6031 (n3811, n_2281, n_2486);
  not g6032 (n_2487, n3808);
  not g6033 (n_2488, n3811);
  and g6034 (n3812, n_2487, n_2488);
  and g6035 (n3813, n_722, n_2483);
  and g6036 (n3814, n_2484, n3813);
  not g6037 (n_2489, n3812);
  not g6038 (n_2490, n3814);
  and g6039 (n3815, n_2489, n_2490);
  not g6040 (n_2491, n3805);
  not g6041 (n_2492, n3815);
  and g6042 (n3816, n_2491, n_2492);
  not g6043 (n_2493, n3816);
  and g6044 (n3817, \asqrt[54] , n_2493);
  and g6048 (n3821, n_2291, n_2290);
  and g6049 (n3822, \asqrt[40] , n3821);
  not g6050 (n_2494, n3822);
  and g6051 (n3823, n_2289, n_2494);
  not g6052 (n_2495, n3820);
  not g6053 (n_2496, n3823);
  and g6054 (n3824, n_2495, n_2496);
  and g6055 (n3825, n_618, n_2491);
  and g6056 (n3826, n_2492, n3825);
  not g6057 (n_2497, n3824);
  not g6058 (n_2498, n3826);
  and g6059 (n3827, n_2497, n_2498);
  not g6060 (n_2499, n3817);
  not g6061 (n_2500, n3827);
  and g6062 (n3828, n_2499, n_2500);
  not g6063 (n_2501, n3828);
  and g6064 (n3829, \asqrt[55] , n_2501);
  and g6068 (n3833, n_2299, n_2298);
  and g6069 (n3834, \asqrt[40] , n3833);
  not g6070 (n_2502, n3834);
  and g6071 (n3835, n_2297, n_2502);
  not g6072 (n_2503, n3832);
  not g6073 (n_2504, n3835);
  and g6074 (n3836, n_2503, n_2504);
  and g6075 (n3837, n_522, n_2499);
  and g6076 (n3838, n_2500, n3837);
  not g6077 (n_2505, n3836);
  not g6078 (n_2506, n3838);
  and g6079 (n3839, n_2505, n_2506);
  not g6080 (n_2507, n3829);
  not g6081 (n_2508, n3839);
  and g6082 (n3840, n_2507, n_2508);
  not g6083 (n_2509, n3840);
  and g6084 (n3841, \asqrt[56] , n_2509);
  and g6088 (n3845, n_2307, n_2306);
  and g6089 (n3846, \asqrt[40] , n3845);
  not g6090 (n_2510, n3846);
  and g6091 (n3847, n_2305, n_2510);
  not g6092 (n_2511, n3844);
  not g6093 (n_2512, n3847);
  and g6094 (n3848, n_2511, n_2512);
  and g6095 (n3849, n_434, n_2507);
  and g6096 (n3850, n_2508, n3849);
  not g6097 (n_2513, n3848);
  not g6098 (n_2514, n3850);
  and g6099 (n3851, n_2513, n_2514);
  not g6100 (n_2515, n3841);
  not g6101 (n_2516, n3851);
  and g6102 (n3852, n_2515, n_2516);
  not g6103 (n_2517, n3852);
  and g6104 (n3853, \asqrt[57] , n_2517);
  and g6105 (n3854, n_354, n_2515);
  and g6106 (n3855, n_2516, n3854);
  and g6110 (n3859, n_2315, n_2313);
  and g6111 (n3860, \asqrt[40] , n3859);
  not g6112 (n_2518, n3860);
  and g6113 (n3861, n_2314, n_2518);
  not g6114 (n_2519, n3858);
  not g6115 (n_2520, n3861);
  and g6116 (n3862, n_2519, n_2520);
  not g6117 (n_2521, n3855);
  not g6118 (n_2522, n3862);
  and g6119 (n3863, n_2521, n_2522);
  not g6120 (n_2523, n3853);
  not g6121 (n_2524, n3863);
  and g6122 (n3864, n_2523, n_2524);
  not g6123 (n_2525, n3864);
  and g6124 (n3865, \asqrt[58] , n_2525);
  and g6128 (n3869, n_2323, n_2322);
  and g6129 (n3870, \asqrt[40] , n3869);
  not g6130 (n_2526, n3870);
  and g6131 (n3871, n_2321, n_2526);
  not g6132 (n_2527, n3868);
  not g6133 (n_2528, n3871);
  and g6134 (n3872, n_2527, n_2528);
  and g6135 (n3873, n_282, n_2523);
  and g6136 (n3874, n_2524, n3873);
  not g6137 (n_2529, n3872);
  not g6138 (n_2530, n3874);
  and g6139 (n3875, n_2529, n_2530);
  not g6140 (n_2531, n3865);
  not g6141 (n_2532, n3875);
  and g6142 (n3876, n_2531, n_2532);
  not g6143 (n_2533, n3876);
  and g6144 (n3877, \asqrt[59] , n_2533);
  and g6148 (n3881, n_2331, n_2330);
  and g6149 (n3882, \asqrt[40] , n3881);
  not g6150 (n_2534, n3882);
  and g6151 (n3883, n_2329, n_2534);
  not g6152 (n_2535, n3880);
  not g6153 (n_2536, n3883);
  and g6154 (n3884, n_2535, n_2536);
  and g6155 (n3885, n_218, n_2531);
  and g6156 (n3886, n_2532, n3885);
  not g6157 (n_2537, n3884);
  not g6158 (n_2538, n3886);
  and g6159 (n3887, n_2537, n_2538);
  not g6160 (n_2539, n3877);
  not g6161 (n_2540, n3887);
  and g6162 (n3888, n_2539, n_2540);
  not g6163 (n_2541, n3888);
  and g6164 (n3889, \asqrt[60] , n_2541);
  and g6168 (n3893, n_2339, n_2338);
  and g6169 (n3894, \asqrt[40] , n3893);
  not g6170 (n_2542, n3894);
  and g6171 (n3895, n_2337, n_2542);
  not g6172 (n_2543, n3892);
  not g6173 (n_2544, n3895);
  and g6174 (n3896, n_2543, n_2544);
  and g6175 (n3897, n_162, n_2539);
  and g6176 (n3898, n_2540, n3897);
  not g6177 (n_2545, n3896);
  not g6178 (n_2546, n3898);
  and g6179 (n3899, n_2545, n_2546);
  not g6180 (n_2547, n3889);
  not g6181 (n_2548, n3899);
  and g6182 (n3900, n_2547, n_2548);
  not g6183 (n_2549, n3900);
  and g6184 (n3901, \asqrt[61] , n_2549);
  and g6188 (n3905, n_2347, n_2346);
  and g6189 (n3906, \asqrt[40] , n3905);
  not g6190 (n_2550, n3906);
  and g6191 (n3907, n_2345, n_2550);
  not g6192 (n_2551, n3904);
  not g6193 (n_2552, n3907);
  and g6194 (n3908, n_2551, n_2552);
  and g6195 (n3909, n_115, n_2547);
  and g6196 (n3910, n_2548, n3909);
  not g6197 (n_2553, n3908);
  not g6198 (n_2554, n3910);
  and g6199 (n3911, n_2553, n_2554);
  not g6200 (n_2555, n3901);
  not g6201 (n_2556, n3911);
  and g6202 (n3912, n_2555, n_2556);
  not g6203 (n_2557, n3912);
  and g6204 (n3913, \asqrt[62] , n_2557);
  and g6208 (n3917, n_2355, n_2354);
  and g6209 (n3918, \asqrt[40] , n3917);
  not g6210 (n_2558, n3918);
  and g6211 (n3919, n_2353, n_2558);
  not g6212 (n_2559, n3916);
  not g6213 (n_2560, n3919);
  and g6214 (n3920, n_2559, n_2560);
  and g6215 (n3921, n_76, n_2555);
  and g6216 (n3922, n_2556, n3921);
  not g6217 (n_2561, n3920);
  not g6218 (n_2562, n3922);
  and g6219 (n3923, n_2561, n_2562);
  not g6220 (n_2563, n3913);
  not g6221 (n_2564, n3923);
  and g6222 (n3924, n_2563, n_2564);
  and g6226 (n3928, n_2363, n_2362);
  and g6227 (n3929, \asqrt[40] , n3928);
  not g6228 (n_2565, n3929);
  and g6229 (n3930, n_2361, n_2565);
  not g6230 (n_2566, n3927);
  not g6231 (n_2567, n3930);
  and g6232 (n3931, n_2566, n_2567);
  and g6233 (n3932, n_2370, n_2369);
  and g6234 (n3933, \asqrt[40] , n3932);
  not g6237 (n_2569, n3931);
  not g6239 (n_2570, n3924);
  not g6241 (n_2571, n3936);
  and g6242 (n3937, n_21, n_2571);
  and g6243 (n3938, n_2563, n3931);
  and g6244 (n3939, n_2564, n3938);
  and g6245 (n3940, n_2369, \asqrt[40] );
  not g6246 (n_2572, n3940);
  and g6247 (n3941, n3628, n_2572);
  not g6248 (n_2573, n3932);
  and g6249 (n3942, \asqrt[63] , n_2573);
  not g6250 (n_2574, n3941);
  and g6251 (n3943, n_2574, n3942);
  not g6257 (n_2575, n3943);
  not g6258 (n_2576, n3948);
  not g6260 (n_2577, n3939);
  and g6264 (n3952, \a[78] , \asqrt[39] );
  not g6265 (n_2582, \a[76] );
  not g6266 (n_2583, \a[77] );
  and g6267 (n3953, n_2582, n_2583);
  and g6268 (n3954, n_2382, n3953);
  not g6269 (n_2584, n3952);
  not g6270 (n_2585, n3954);
  and g6271 (n3955, n_2584, n_2585);
  not g6272 (n_2586, n3955);
  and g6273 (n3956, \asqrt[40] , n_2586);
  and g6279 (n3962, n_2382, \asqrt[39] );
  not g6280 (n_2587, n3962);
  and g6281 (n3963, \a[79] , n_2587);
  and g6282 (n3964, n3657, \asqrt[39] );
  not g6283 (n_2588, n3963);
  not g6284 (n_2589, n3964);
  and g6285 (n3965, n_2588, n_2589);
  not g6286 (n_2590, n3961);
  and g6287 (n3966, n_2590, n3965);
  not g6288 (n_2591, n3956);
  not g6289 (n_2592, n3966);
  and g6290 (n3967, n_2591, n_2592);
  not g6291 (n_2593, n3967);
  and g6292 (n3968, \asqrt[41] , n_2593);
  not g6293 (n_2594, \asqrt[41] );
  and g6294 (n3969, n_2594, n_2591);
  and g6295 (n3970, n_2592, n3969);
  not g6299 (n_2595, n3937);
  not g6301 (n_2596, n3974);
  and g6302 (n3975, n_2589, n_2596);
  not g6303 (n_2597, n3975);
  and g6304 (n3976, \a[80] , n_2597);
  and g6305 (n3977, n_2190, n_2596);
  and g6306 (n3978, n_2589, n3977);
  not g6307 (n_2598, n3976);
  not g6308 (n_2599, n3978);
  and g6309 (n3979, n_2598, n_2599);
  not g6310 (n_2600, n3970);
  not g6311 (n_2601, n3979);
  and g6312 (n3980, n_2600, n_2601);
  not g6313 (n_2602, n3968);
  not g6314 (n_2603, n3980);
  and g6315 (n3981, n_2602, n_2603);
  not g6316 (n_2604, n3981);
  and g6317 (n3982, \asqrt[42] , n_2604);
  and g6318 (n3983, n_2391, n_2390);
  not g6319 (n_2605, n3669);
  and g6320 (n3984, n_2605, n3983);
  and g6321 (n3985, \asqrt[39] , n3984);
  and g6322 (n3986, \asqrt[39] , n3983);
  not g6323 (n_2606, n3986);
  and g6324 (n3987, n3669, n_2606);
  not g6325 (n_2607, n3985);
  not g6326 (n_2608, n3987);
  and g6327 (n3988, n_2607, n_2608);
  and g6328 (n3989, n_2394, n_2602);
  and g6329 (n3990, n_2603, n3989);
  not g6330 (n_2609, n3988);
  not g6331 (n_2610, n3990);
  and g6332 (n3991, n_2609, n_2610);
  not g6333 (n_2611, n3982);
  not g6334 (n_2612, n3991);
  and g6335 (n3992, n_2611, n_2612);
  not g6336 (n_2613, n3992);
  and g6337 (n3993, \asqrt[43] , n_2613);
  and g6341 (n3997, n_2402, n_2400);
  and g6342 (n3998, \asqrt[39] , n3997);
  not g6343 (n_2614, n3998);
  and g6344 (n3999, n_2401, n_2614);
  not g6345 (n_2615, n3996);
  not g6346 (n_2616, n3999);
  and g6347 (n4000, n_2615, n_2616);
  and g6348 (n4001, n_2202, n_2611);
  and g6349 (n4002, n_2612, n4001);
  not g6350 (n_2617, n4000);
  not g6351 (n_2618, n4002);
  and g6352 (n4003, n_2617, n_2618);
  not g6353 (n_2619, n3993);
  not g6354 (n_2620, n4003);
  and g6355 (n4004, n_2619, n_2620);
  not g6356 (n_2621, n4004);
  and g6357 (n4005, \asqrt[44] , n_2621);
  and g6361 (n4009, n_2411, n_2410);
  and g6362 (n4010, \asqrt[39] , n4009);
  not g6363 (n_2622, n4010);
  and g6364 (n4011, n_2409, n_2622);
  not g6365 (n_2623, n4008);
  not g6366 (n_2624, n4011);
  and g6367 (n4012, n_2623, n_2624);
  and g6368 (n4013, n_2018, n_2619);
  and g6369 (n4014, n_2620, n4013);
  not g6370 (n_2625, n4012);
  not g6371 (n_2626, n4014);
  and g6372 (n4015, n_2625, n_2626);
  not g6373 (n_2627, n4005);
  not g6374 (n_2628, n4015);
  and g6375 (n4016, n_2627, n_2628);
  not g6376 (n_2629, n4016);
  and g6377 (n4017, \asqrt[45] , n_2629);
  and g6381 (n4021, n_2419, n_2418);
  and g6382 (n4022, \asqrt[39] , n4021);
  not g6383 (n_2630, n4022);
  and g6384 (n4023, n_2417, n_2630);
  not g6385 (n_2631, n4020);
  not g6386 (n_2632, n4023);
  and g6387 (n4024, n_2631, n_2632);
  and g6388 (n4025, n_1842, n_2627);
  and g6389 (n4026, n_2628, n4025);
  not g6390 (n_2633, n4024);
  not g6391 (n_2634, n4026);
  and g6392 (n4027, n_2633, n_2634);
  not g6393 (n_2635, n4017);
  not g6394 (n_2636, n4027);
  and g6395 (n4028, n_2635, n_2636);
  not g6396 (n_2637, n4028);
  and g6397 (n4029, \asqrt[46] , n_2637);
  and g6401 (n4033, n_2427, n_2426);
  and g6402 (n4034, \asqrt[39] , n4033);
  not g6403 (n_2638, n4034);
  and g6404 (n4035, n_2425, n_2638);
  not g6405 (n_2639, n4032);
  not g6406 (n_2640, n4035);
  and g6407 (n4036, n_2639, n_2640);
  and g6408 (n4037, n_1674, n_2635);
  and g6409 (n4038, n_2636, n4037);
  not g6410 (n_2641, n4036);
  not g6411 (n_2642, n4038);
  and g6412 (n4039, n_2641, n_2642);
  not g6413 (n_2643, n4029);
  not g6414 (n_2644, n4039);
  and g6415 (n4040, n_2643, n_2644);
  not g6416 (n_2645, n4040);
  and g6417 (n4041, \asqrt[47] , n_2645);
  and g6421 (n4045, n_2435, n_2434);
  and g6422 (n4046, \asqrt[39] , n4045);
  not g6423 (n_2646, n4046);
  and g6424 (n4047, n_2433, n_2646);
  not g6425 (n_2647, n4044);
  not g6426 (n_2648, n4047);
  and g6427 (n4048, n_2647, n_2648);
  and g6428 (n4049, n_1514, n_2643);
  and g6429 (n4050, n_2644, n4049);
  not g6430 (n_2649, n4048);
  not g6431 (n_2650, n4050);
  and g6432 (n4051, n_2649, n_2650);
  not g6433 (n_2651, n4041);
  not g6434 (n_2652, n4051);
  and g6435 (n4052, n_2651, n_2652);
  not g6436 (n_2653, n4052);
  and g6437 (n4053, \asqrt[48] , n_2653);
  and g6441 (n4057, n_2443, n_2442);
  and g6442 (n4058, \asqrt[39] , n4057);
  not g6443 (n_2654, n4058);
  and g6444 (n4059, n_2441, n_2654);
  not g6445 (n_2655, n4056);
  not g6446 (n_2656, n4059);
  and g6447 (n4060, n_2655, n_2656);
  and g6448 (n4061, n_1362, n_2651);
  and g6449 (n4062, n_2652, n4061);
  not g6450 (n_2657, n4060);
  not g6451 (n_2658, n4062);
  and g6452 (n4063, n_2657, n_2658);
  not g6453 (n_2659, n4053);
  not g6454 (n_2660, n4063);
  and g6455 (n4064, n_2659, n_2660);
  not g6456 (n_2661, n4064);
  and g6457 (n4065, \asqrt[49] , n_2661);
  and g6461 (n4069, n_2451, n_2450);
  and g6462 (n4070, \asqrt[39] , n4069);
  not g6463 (n_2662, n4070);
  and g6464 (n4071, n_2449, n_2662);
  not g6465 (n_2663, n4068);
  not g6466 (n_2664, n4071);
  and g6467 (n4072, n_2663, n_2664);
  and g6468 (n4073, n_1218, n_2659);
  and g6469 (n4074, n_2660, n4073);
  not g6470 (n_2665, n4072);
  not g6471 (n_2666, n4074);
  and g6472 (n4075, n_2665, n_2666);
  not g6473 (n_2667, n4065);
  not g6474 (n_2668, n4075);
  and g6475 (n4076, n_2667, n_2668);
  not g6476 (n_2669, n4076);
  and g6477 (n4077, \asqrt[50] , n_2669);
  and g6481 (n4081, n_2459, n_2458);
  and g6482 (n4082, \asqrt[39] , n4081);
  not g6483 (n_2670, n4082);
  and g6484 (n4083, n_2457, n_2670);
  not g6485 (n_2671, n4080);
  not g6486 (n_2672, n4083);
  and g6487 (n4084, n_2671, n_2672);
  and g6488 (n4085, n_1082, n_2667);
  and g6489 (n4086, n_2668, n4085);
  not g6490 (n_2673, n4084);
  not g6491 (n_2674, n4086);
  and g6492 (n4087, n_2673, n_2674);
  not g6493 (n_2675, n4077);
  not g6494 (n_2676, n4087);
  and g6495 (n4088, n_2675, n_2676);
  not g6496 (n_2677, n4088);
  and g6497 (n4089, \asqrt[51] , n_2677);
  and g6501 (n4093, n_2467, n_2466);
  and g6502 (n4094, \asqrt[39] , n4093);
  not g6503 (n_2678, n4094);
  and g6504 (n4095, n_2465, n_2678);
  not g6505 (n_2679, n4092);
  not g6506 (n_2680, n4095);
  and g6507 (n4096, n_2679, n_2680);
  and g6508 (n4097, n_954, n_2675);
  and g6509 (n4098, n_2676, n4097);
  not g6510 (n_2681, n4096);
  not g6511 (n_2682, n4098);
  and g6512 (n4099, n_2681, n_2682);
  not g6513 (n_2683, n4089);
  not g6514 (n_2684, n4099);
  and g6515 (n4100, n_2683, n_2684);
  not g6516 (n_2685, n4100);
  and g6517 (n4101, \asqrt[52] , n_2685);
  and g6521 (n4105, n_2475, n_2474);
  and g6522 (n4106, \asqrt[39] , n4105);
  not g6523 (n_2686, n4106);
  and g6524 (n4107, n_2473, n_2686);
  not g6525 (n_2687, n4104);
  not g6526 (n_2688, n4107);
  and g6527 (n4108, n_2687, n_2688);
  and g6528 (n4109, n_834, n_2683);
  and g6529 (n4110, n_2684, n4109);
  not g6530 (n_2689, n4108);
  not g6531 (n_2690, n4110);
  and g6532 (n4111, n_2689, n_2690);
  not g6533 (n_2691, n4101);
  not g6534 (n_2692, n4111);
  and g6535 (n4112, n_2691, n_2692);
  not g6536 (n_2693, n4112);
  and g6537 (n4113, \asqrt[53] , n_2693);
  and g6541 (n4117, n_2483, n_2482);
  and g6542 (n4118, \asqrt[39] , n4117);
  not g6543 (n_2694, n4118);
  and g6544 (n4119, n_2481, n_2694);
  not g6545 (n_2695, n4116);
  not g6546 (n_2696, n4119);
  and g6547 (n4120, n_2695, n_2696);
  and g6548 (n4121, n_722, n_2691);
  and g6549 (n4122, n_2692, n4121);
  not g6550 (n_2697, n4120);
  not g6551 (n_2698, n4122);
  and g6552 (n4123, n_2697, n_2698);
  not g6553 (n_2699, n4113);
  not g6554 (n_2700, n4123);
  and g6555 (n4124, n_2699, n_2700);
  not g6556 (n_2701, n4124);
  and g6557 (n4125, \asqrt[54] , n_2701);
  and g6561 (n4129, n_2491, n_2490);
  and g6562 (n4130, \asqrt[39] , n4129);
  not g6563 (n_2702, n4130);
  and g6564 (n4131, n_2489, n_2702);
  not g6565 (n_2703, n4128);
  not g6566 (n_2704, n4131);
  and g6567 (n4132, n_2703, n_2704);
  and g6568 (n4133, n_618, n_2699);
  and g6569 (n4134, n_2700, n4133);
  not g6570 (n_2705, n4132);
  not g6571 (n_2706, n4134);
  and g6572 (n4135, n_2705, n_2706);
  not g6573 (n_2707, n4125);
  not g6574 (n_2708, n4135);
  and g6575 (n4136, n_2707, n_2708);
  not g6576 (n_2709, n4136);
  and g6577 (n4137, \asqrt[55] , n_2709);
  and g6581 (n4141, n_2499, n_2498);
  and g6582 (n4142, \asqrt[39] , n4141);
  not g6583 (n_2710, n4142);
  and g6584 (n4143, n_2497, n_2710);
  not g6585 (n_2711, n4140);
  not g6586 (n_2712, n4143);
  and g6587 (n4144, n_2711, n_2712);
  and g6588 (n4145, n_522, n_2707);
  and g6589 (n4146, n_2708, n4145);
  not g6590 (n_2713, n4144);
  not g6591 (n_2714, n4146);
  and g6592 (n4147, n_2713, n_2714);
  not g6593 (n_2715, n4137);
  not g6594 (n_2716, n4147);
  and g6595 (n4148, n_2715, n_2716);
  not g6596 (n_2717, n4148);
  and g6597 (n4149, \asqrt[56] , n_2717);
  and g6601 (n4153, n_2507, n_2506);
  and g6602 (n4154, \asqrt[39] , n4153);
  not g6603 (n_2718, n4154);
  and g6604 (n4155, n_2505, n_2718);
  not g6605 (n_2719, n4152);
  not g6606 (n_2720, n4155);
  and g6607 (n4156, n_2719, n_2720);
  and g6608 (n4157, n_434, n_2715);
  and g6609 (n4158, n_2716, n4157);
  not g6610 (n_2721, n4156);
  not g6611 (n_2722, n4158);
  and g6612 (n4159, n_2721, n_2722);
  not g6613 (n_2723, n4149);
  not g6614 (n_2724, n4159);
  and g6615 (n4160, n_2723, n_2724);
  not g6616 (n_2725, n4160);
  and g6617 (n4161, \asqrt[57] , n_2725);
  and g6621 (n4165, n_2515, n_2514);
  and g6622 (n4166, \asqrt[39] , n4165);
  not g6623 (n_2726, n4166);
  and g6624 (n4167, n_2513, n_2726);
  not g6625 (n_2727, n4164);
  not g6626 (n_2728, n4167);
  and g6627 (n4168, n_2727, n_2728);
  and g6628 (n4169, n_354, n_2723);
  and g6629 (n4170, n_2724, n4169);
  not g6630 (n_2729, n4168);
  not g6631 (n_2730, n4170);
  and g6632 (n4171, n_2729, n_2730);
  not g6633 (n_2731, n4161);
  not g6634 (n_2732, n4171);
  and g6635 (n4172, n_2731, n_2732);
  not g6636 (n_2733, n4172);
  and g6637 (n4173, \asqrt[58] , n_2733);
  and g6638 (n4174, n_282, n_2731);
  and g6639 (n4175, n_2732, n4174);
  and g6643 (n4179, n_2523, n_2521);
  and g6644 (n4180, \asqrt[39] , n4179);
  not g6645 (n_2734, n4180);
  and g6646 (n4181, n_2522, n_2734);
  not g6647 (n_2735, n4178);
  not g6648 (n_2736, n4181);
  and g6649 (n4182, n_2735, n_2736);
  not g6650 (n_2737, n4175);
  not g6651 (n_2738, n4182);
  and g6652 (n4183, n_2737, n_2738);
  not g6653 (n_2739, n4173);
  not g6654 (n_2740, n4183);
  and g6655 (n4184, n_2739, n_2740);
  not g6656 (n_2741, n4184);
  and g6657 (n4185, \asqrt[59] , n_2741);
  and g6661 (n4189, n_2531, n_2530);
  and g6662 (n4190, \asqrt[39] , n4189);
  not g6663 (n_2742, n4190);
  and g6664 (n4191, n_2529, n_2742);
  not g6665 (n_2743, n4188);
  not g6666 (n_2744, n4191);
  and g6667 (n4192, n_2743, n_2744);
  and g6668 (n4193, n_218, n_2739);
  and g6669 (n4194, n_2740, n4193);
  not g6670 (n_2745, n4192);
  not g6671 (n_2746, n4194);
  and g6672 (n4195, n_2745, n_2746);
  not g6673 (n_2747, n4185);
  not g6674 (n_2748, n4195);
  and g6675 (n4196, n_2747, n_2748);
  not g6676 (n_2749, n4196);
  and g6677 (n4197, \asqrt[60] , n_2749);
  and g6681 (n4201, n_2539, n_2538);
  and g6682 (n4202, \asqrt[39] , n4201);
  not g6683 (n_2750, n4202);
  and g6684 (n4203, n_2537, n_2750);
  not g6685 (n_2751, n4200);
  not g6686 (n_2752, n4203);
  and g6687 (n4204, n_2751, n_2752);
  and g6688 (n4205, n_162, n_2747);
  and g6689 (n4206, n_2748, n4205);
  not g6690 (n_2753, n4204);
  not g6691 (n_2754, n4206);
  and g6692 (n4207, n_2753, n_2754);
  not g6693 (n_2755, n4197);
  not g6694 (n_2756, n4207);
  and g6695 (n4208, n_2755, n_2756);
  not g6696 (n_2757, n4208);
  and g6697 (n4209, \asqrt[61] , n_2757);
  and g6701 (n4213, n_2547, n_2546);
  and g6702 (n4214, \asqrt[39] , n4213);
  not g6703 (n_2758, n4214);
  and g6704 (n4215, n_2545, n_2758);
  not g6705 (n_2759, n4212);
  not g6706 (n_2760, n4215);
  and g6707 (n4216, n_2759, n_2760);
  and g6708 (n4217, n_115, n_2755);
  and g6709 (n4218, n_2756, n4217);
  not g6710 (n_2761, n4216);
  not g6711 (n_2762, n4218);
  and g6712 (n4219, n_2761, n_2762);
  not g6713 (n_2763, n4209);
  not g6714 (n_2764, n4219);
  and g6715 (n4220, n_2763, n_2764);
  not g6716 (n_2765, n4220);
  and g6717 (n4221, \asqrt[62] , n_2765);
  and g6721 (n4225, n_2555, n_2554);
  and g6722 (n4226, \asqrt[39] , n4225);
  not g6723 (n_2766, n4226);
  and g6724 (n4227, n_2553, n_2766);
  not g6725 (n_2767, n4224);
  not g6726 (n_2768, n4227);
  and g6727 (n4228, n_2767, n_2768);
  and g6728 (n4229, n_76, n_2763);
  and g6729 (n4230, n_2764, n4229);
  not g6730 (n_2769, n4228);
  not g6731 (n_2770, n4230);
  and g6732 (n4231, n_2769, n_2770);
  not g6733 (n_2771, n4221);
  not g6734 (n_2772, n4231);
  and g6735 (n4232, n_2771, n_2772);
  and g6739 (n4236, n_2563, n_2562);
  and g6740 (n4237, \asqrt[39] , n4236);
  not g6741 (n_2773, n4237);
  and g6742 (n4238, n_2561, n_2773);
  not g6743 (n_2774, n4235);
  not g6744 (n_2775, n4238);
  and g6745 (n4239, n_2774, n_2775);
  and g6746 (n4240, n_2570, n_2569);
  and g6747 (n4241, \asqrt[39] , n4240);
  not g6750 (n_2777, n4239);
  not g6752 (n_2778, n4232);
  not g6754 (n_2779, n4244);
  and g6755 (n4245, n_21, n_2779);
  and g6756 (n4246, n_2771, n4239);
  and g6757 (n4247, n_2772, n4246);
  and g6758 (n4248, n_2569, \asqrt[39] );
  not g6759 (n_2780, n4248);
  and g6760 (n4249, n3924, n_2780);
  not g6761 (n_2781, n4240);
  and g6762 (n4250, \asqrt[63] , n_2781);
  not g6763 (n_2782, n4249);
  and g6764 (n4251, n_2782, n4250);
  not g6770 (n_2783, n4251);
  not g6771 (n_2784, n4256);
  not g6773 (n_2785, n4247);
  and g6777 (n4260, \a[76] , \asqrt[38] );
  not g6778 (n_2790, \a[74] );
  not g6779 (n_2791, \a[75] );
  and g6780 (n4261, n_2790, n_2791);
  and g6781 (n4262, n_2582, n4261);
  not g6782 (n_2792, n4260);
  not g6783 (n_2793, n4262);
  and g6784 (n4263, n_2792, n_2793);
  not g6785 (n_2794, n4263);
  and g6786 (n4264, \asqrt[39] , n_2794);
  and g6792 (n4270, n_2582, \asqrt[38] );
  not g6793 (n_2795, n4270);
  and g6794 (n4271, \a[77] , n_2795);
  and g6795 (n4272, n3953, \asqrt[38] );
  not g6796 (n_2796, n4271);
  not g6797 (n_2797, n4272);
  and g6798 (n4273, n_2796, n_2797);
  not g6799 (n_2798, n4269);
  and g6800 (n4274, n_2798, n4273);
  not g6801 (n_2799, n4264);
  not g6802 (n_2800, n4274);
  and g6803 (n4275, n_2799, n_2800);
  not g6804 (n_2801, n4275);
  and g6805 (n4276, \asqrt[40] , n_2801);
  not g6806 (n_2802, \asqrt[40] );
  and g6807 (n4277, n_2802, n_2799);
  and g6808 (n4278, n_2800, n4277);
  not g6812 (n_2803, n4245);
  not g6814 (n_2804, n4282);
  and g6815 (n4283, n_2797, n_2804);
  not g6816 (n_2805, n4283);
  and g6817 (n4284, \a[78] , n_2805);
  and g6818 (n4285, n_2382, n_2804);
  and g6819 (n4286, n_2797, n4285);
  not g6820 (n_2806, n4284);
  not g6821 (n_2807, n4286);
  and g6822 (n4287, n_2806, n_2807);
  not g6823 (n_2808, n4278);
  not g6824 (n_2809, n4287);
  and g6825 (n4288, n_2808, n_2809);
  not g6826 (n_2810, n4276);
  not g6827 (n_2811, n4288);
  and g6828 (n4289, n_2810, n_2811);
  not g6829 (n_2812, n4289);
  and g6830 (n4290, \asqrt[41] , n_2812);
  and g6831 (n4291, n_2591, n_2590);
  not g6832 (n_2813, n3965);
  and g6833 (n4292, n_2813, n4291);
  and g6834 (n4293, \asqrt[38] , n4292);
  and g6835 (n4294, \asqrt[38] , n4291);
  not g6836 (n_2814, n4294);
  and g6837 (n4295, n3965, n_2814);
  not g6838 (n_2815, n4293);
  not g6839 (n_2816, n4295);
  and g6840 (n4296, n_2815, n_2816);
  and g6841 (n4297, n_2594, n_2810);
  and g6842 (n4298, n_2811, n4297);
  not g6843 (n_2817, n4296);
  not g6844 (n_2818, n4298);
  and g6845 (n4299, n_2817, n_2818);
  not g6846 (n_2819, n4290);
  not g6847 (n_2820, n4299);
  and g6848 (n4300, n_2819, n_2820);
  not g6849 (n_2821, n4300);
  and g6850 (n4301, \asqrt[42] , n_2821);
  and g6854 (n4305, n_2602, n_2600);
  and g6855 (n4306, \asqrt[38] , n4305);
  not g6856 (n_2822, n4306);
  and g6857 (n4307, n_2601, n_2822);
  not g6858 (n_2823, n4304);
  not g6859 (n_2824, n4307);
  and g6860 (n4308, n_2823, n_2824);
  and g6861 (n4309, n_2394, n_2819);
  and g6862 (n4310, n_2820, n4309);
  not g6863 (n_2825, n4308);
  not g6864 (n_2826, n4310);
  and g6865 (n4311, n_2825, n_2826);
  not g6866 (n_2827, n4301);
  not g6867 (n_2828, n4311);
  and g6868 (n4312, n_2827, n_2828);
  not g6869 (n_2829, n4312);
  and g6870 (n4313, \asqrt[43] , n_2829);
  and g6874 (n4317, n_2611, n_2610);
  and g6875 (n4318, \asqrt[38] , n4317);
  not g6876 (n_2830, n4318);
  and g6877 (n4319, n_2609, n_2830);
  not g6878 (n_2831, n4316);
  not g6879 (n_2832, n4319);
  and g6880 (n4320, n_2831, n_2832);
  and g6881 (n4321, n_2202, n_2827);
  and g6882 (n4322, n_2828, n4321);
  not g6883 (n_2833, n4320);
  not g6884 (n_2834, n4322);
  and g6885 (n4323, n_2833, n_2834);
  not g6886 (n_2835, n4313);
  not g6887 (n_2836, n4323);
  and g6888 (n4324, n_2835, n_2836);
  not g6889 (n_2837, n4324);
  and g6890 (n4325, \asqrt[44] , n_2837);
  and g6894 (n4329, n_2619, n_2618);
  and g6895 (n4330, \asqrt[38] , n4329);
  not g6896 (n_2838, n4330);
  and g6897 (n4331, n_2617, n_2838);
  not g6898 (n_2839, n4328);
  not g6899 (n_2840, n4331);
  and g6900 (n4332, n_2839, n_2840);
  and g6901 (n4333, n_2018, n_2835);
  and g6902 (n4334, n_2836, n4333);
  not g6903 (n_2841, n4332);
  not g6904 (n_2842, n4334);
  and g6905 (n4335, n_2841, n_2842);
  not g6906 (n_2843, n4325);
  not g6907 (n_2844, n4335);
  and g6908 (n4336, n_2843, n_2844);
  not g6909 (n_2845, n4336);
  and g6910 (n4337, \asqrt[45] , n_2845);
  and g6914 (n4341, n_2627, n_2626);
  and g6915 (n4342, \asqrt[38] , n4341);
  not g6916 (n_2846, n4342);
  and g6917 (n4343, n_2625, n_2846);
  not g6918 (n_2847, n4340);
  not g6919 (n_2848, n4343);
  and g6920 (n4344, n_2847, n_2848);
  and g6921 (n4345, n_1842, n_2843);
  and g6922 (n4346, n_2844, n4345);
  not g6923 (n_2849, n4344);
  not g6924 (n_2850, n4346);
  and g6925 (n4347, n_2849, n_2850);
  not g6926 (n_2851, n4337);
  not g6927 (n_2852, n4347);
  and g6928 (n4348, n_2851, n_2852);
  not g6929 (n_2853, n4348);
  and g6930 (n4349, \asqrt[46] , n_2853);
  and g6934 (n4353, n_2635, n_2634);
  and g6935 (n4354, \asqrt[38] , n4353);
  not g6936 (n_2854, n4354);
  and g6937 (n4355, n_2633, n_2854);
  not g6938 (n_2855, n4352);
  not g6939 (n_2856, n4355);
  and g6940 (n4356, n_2855, n_2856);
  and g6941 (n4357, n_1674, n_2851);
  and g6942 (n4358, n_2852, n4357);
  not g6943 (n_2857, n4356);
  not g6944 (n_2858, n4358);
  and g6945 (n4359, n_2857, n_2858);
  not g6946 (n_2859, n4349);
  not g6947 (n_2860, n4359);
  and g6948 (n4360, n_2859, n_2860);
  not g6949 (n_2861, n4360);
  and g6950 (n4361, \asqrt[47] , n_2861);
  and g6954 (n4365, n_2643, n_2642);
  and g6955 (n4366, \asqrt[38] , n4365);
  not g6956 (n_2862, n4366);
  and g6957 (n4367, n_2641, n_2862);
  not g6958 (n_2863, n4364);
  not g6959 (n_2864, n4367);
  and g6960 (n4368, n_2863, n_2864);
  and g6961 (n4369, n_1514, n_2859);
  and g6962 (n4370, n_2860, n4369);
  not g6963 (n_2865, n4368);
  not g6964 (n_2866, n4370);
  and g6965 (n4371, n_2865, n_2866);
  not g6966 (n_2867, n4361);
  not g6967 (n_2868, n4371);
  and g6968 (n4372, n_2867, n_2868);
  not g6969 (n_2869, n4372);
  and g6970 (n4373, \asqrt[48] , n_2869);
  and g6974 (n4377, n_2651, n_2650);
  and g6975 (n4378, \asqrt[38] , n4377);
  not g6976 (n_2870, n4378);
  and g6977 (n4379, n_2649, n_2870);
  not g6978 (n_2871, n4376);
  not g6979 (n_2872, n4379);
  and g6980 (n4380, n_2871, n_2872);
  and g6981 (n4381, n_1362, n_2867);
  and g6982 (n4382, n_2868, n4381);
  not g6983 (n_2873, n4380);
  not g6984 (n_2874, n4382);
  and g6985 (n4383, n_2873, n_2874);
  not g6986 (n_2875, n4373);
  not g6987 (n_2876, n4383);
  and g6988 (n4384, n_2875, n_2876);
  not g6989 (n_2877, n4384);
  and g6990 (n4385, \asqrt[49] , n_2877);
  and g6994 (n4389, n_2659, n_2658);
  and g6995 (n4390, \asqrt[38] , n4389);
  not g6996 (n_2878, n4390);
  and g6997 (n4391, n_2657, n_2878);
  not g6998 (n_2879, n4388);
  not g6999 (n_2880, n4391);
  and g7000 (n4392, n_2879, n_2880);
  and g7001 (n4393, n_1218, n_2875);
  and g7002 (n4394, n_2876, n4393);
  not g7003 (n_2881, n4392);
  not g7004 (n_2882, n4394);
  and g7005 (n4395, n_2881, n_2882);
  not g7006 (n_2883, n4385);
  not g7007 (n_2884, n4395);
  and g7008 (n4396, n_2883, n_2884);
  not g7009 (n_2885, n4396);
  and g7010 (n4397, \asqrt[50] , n_2885);
  and g7014 (n4401, n_2667, n_2666);
  and g7015 (n4402, \asqrt[38] , n4401);
  not g7016 (n_2886, n4402);
  and g7017 (n4403, n_2665, n_2886);
  not g7018 (n_2887, n4400);
  not g7019 (n_2888, n4403);
  and g7020 (n4404, n_2887, n_2888);
  and g7021 (n4405, n_1082, n_2883);
  and g7022 (n4406, n_2884, n4405);
  not g7023 (n_2889, n4404);
  not g7024 (n_2890, n4406);
  and g7025 (n4407, n_2889, n_2890);
  not g7026 (n_2891, n4397);
  not g7027 (n_2892, n4407);
  and g7028 (n4408, n_2891, n_2892);
  not g7029 (n_2893, n4408);
  and g7030 (n4409, \asqrt[51] , n_2893);
  and g7034 (n4413, n_2675, n_2674);
  and g7035 (n4414, \asqrt[38] , n4413);
  not g7036 (n_2894, n4414);
  and g7037 (n4415, n_2673, n_2894);
  not g7038 (n_2895, n4412);
  not g7039 (n_2896, n4415);
  and g7040 (n4416, n_2895, n_2896);
  and g7041 (n4417, n_954, n_2891);
  and g7042 (n4418, n_2892, n4417);
  not g7043 (n_2897, n4416);
  not g7044 (n_2898, n4418);
  and g7045 (n4419, n_2897, n_2898);
  not g7046 (n_2899, n4409);
  not g7047 (n_2900, n4419);
  and g7048 (n4420, n_2899, n_2900);
  not g7049 (n_2901, n4420);
  and g7050 (n4421, \asqrt[52] , n_2901);
  and g7054 (n4425, n_2683, n_2682);
  and g7055 (n4426, \asqrt[38] , n4425);
  not g7056 (n_2902, n4426);
  and g7057 (n4427, n_2681, n_2902);
  not g7058 (n_2903, n4424);
  not g7059 (n_2904, n4427);
  and g7060 (n4428, n_2903, n_2904);
  and g7061 (n4429, n_834, n_2899);
  and g7062 (n4430, n_2900, n4429);
  not g7063 (n_2905, n4428);
  not g7064 (n_2906, n4430);
  and g7065 (n4431, n_2905, n_2906);
  not g7066 (n_2907, n4421);
  not g7067 (n_2908, n4431);
  and g7068 (n4432, n_2907, n_2908);
  not g7069 (n_2909, n4432);
  and g7070 (n4433, \asqrt[53] , n_2909);
  and g7074 (n4437, n_2691, n_2690);
  and g7075 (n4438, \asqrt[38] , n4437);
  not g7076 (n_2910, n4438);
  and g7077 (n4439, n_2689, n_2910);
  not g7078 (n_2911, n4436);
  not g7079 (n_2912, n4439);
  and g7080 (n4440, n_2911, n_2912);
  and g7081 (n4441, n_722, n_2907);
  and g7082 (n4442, n_2908, n4441);
  not g7083 (n_2913, n4440);
  not g7084 (n_2914, n4442);
  and g7085 (n4443, n_2913, n_2914);
  not g7086 (n_2915, n4433);
  not g7087 (n_2916, n4443);
  and g7088 (n4444, n_2915, n_2916);
  not g7089 (n_2917, n4444);
  and g7090 (n4445, \asqrt[54] , n_2917);
  and g7094 (n4449, n_2699, n_2698);
  and g7095 (n4450, \asqrt[38] , n4449);
  not g7096 (n_2918, n4450);
  and g7097 (n4451, n_2697, n_2918);
  not g7098 (n_2919, n4448);
  not g7099 (n_2920, n4451);
  and g7100 (n4452, n_2919, n_2920);
  and g7101 (n4453, n_618, n_2915);
  and g7102 (n4454, n_2916, n4453);
  not g7103 (n_2921, n4452);
  not g7104 (n_2922, n4454);
  and g7105 (n4455, n_2921, n_2922);
  not g7106 (n_2923, n4445);
  not g7107 (n_2924, n4455);
  and g7108 (n4456, n_2923, n_2924);
  not g7109 (n_2925, n4456);
  and g7110 (n4457, \asqrt[55] , n_2925);
  and g7114 (n4461, n_2707, n_2706);
  and g7115 (n4462, \asqrt[38] , n4461);
  not g7116 (n_2926, n4462);
  and g7117 (n4463, n_2705, n_2926);
  not g7118 (n_2927, n4460);
  not g7119 (n_2928, n4463);
  and g7120 (n4464, n_2927, n_2928);
  and g7121 (n4465, n_522, n_2923);
  and g7122 (n4466, n_2924, n4465);
  not g7123 (n_2929, n4464);
  not g7124 (n_2930, n4466);
  and g7125 (n4467, n_2929, n_2930);
  not g7126 (n_2931, n4457);
  not g7127 (n_2932, n4467);
  and g7128 (n4468, n_2931, n_2932);
  not g7129 (n_2933, n4468);
  and g7130 (n4469, \asqrt[56] , n_2933);
  and g7134 (n4473, n_2715, n_2714);
  and g7135 (n4474, \asqrt[38] , n4473);
  not g7136 (n_2934, n4474);
  and g7137 (n4475, n_2713, n_2934);
  not g7138 (n_2935, n4472);
  not g7139 (n_2936, n4475);
  and g7140 (n4476, n_2935, n_2936);
  and g7141 (n4477, n_434, n_2931);
  and g7142 (n4478, n_2932, n4477);
  not g7143 (n_2937, n4476);
  not g7144 (n_2938, n4478);
  and g7145 (n4479, n_2937, n_2938);
  not g7146 (n_2939, n4469);
  not g7147 (n_2940, n4479);
  and g7148 (n4480, n_2939, n_2940);
  not g7149 (n_2941, n4480);
  and g7150 (n4481, \asqrt[57] , n_2941);
  and g7154 (n4485, n_2723, n_2722);
  and g7155 (n4486, \asqrt[38] , n4485);
  not g7156 (n_2942, n4486);
  and g7157 (n4487, n_2721, n_2942);
  not g7158 (n_2943, n4484);
  not g7159 (n_2944, n4487);
  and g7160 (n4488, n_2943, n_2944);
  and g7161 (n4489, n_354, n_2939);
  and g7162 (n4490, n_2940, n4489);
  not g7163 (n_2945, n4488);
  not g7164 (n_2946, n4490);
  and g7165 (n4491, n_2945, n_2946);
  not g7166 (n_2947, n4481);
  not g7167 (n_2948, n4491);
  and g7168 (n4492, n_2947, n_2948);
  not g7169 (n_2949, n4492);
  and g7170 (n4493, \asqrt[58] , n_2949);
  and g7174 (n4497, n_2731, n_2730);
  and g7175 (n4498, \asqrt[38] , n4497);
  not g7176 (n_2950, n4498);
  and g7177 (n4499, n_2729, n_2950);
  not g7178 (n_2951, n4496);
  not g7179 (n_2952, n4499);
  and g7180 (n4500, n_2951, n_2952);
  and g7181 (n4501, n_282, n_2947);
  and g7182 (n4502, n_2948, n4501);
  not g7183 (n_2953, n4500);
  not g7184 (n_2954, n4502);
  and g7185 (n4503, n_2953, n_2954);
  not g7186 (n_2955, n4493);
  not g7187 (n_2956, n4503);
  and g7188 (n4504, n_2955, n_2956);
  not g7189 (n_2957, n4504);
  and g7190 (n4505, \asqrt[59] , n_2957);
  and g7191 (n4506, n_218, n_2955);
  and g7192 (n4507, n_2956, n4506);
  and g7196 (n4511, n_2739, n_2737);
  and g7197 (n4512, \asqrt[38] , n4511);
  not g7198 (n_2958, n4512);
  and g7199 (n4513, n_2738, n_2958);
  not g7200 (n_2959, n4510);
  not g7201 (n_2960, n4513);
  and g7202 (n4514, n_2959, n_2960);
  not g7203 (n_2961, n4507);
  not g7204 (n_2962, n4514);
  and g7205 (n4515, n_2961, n_2962);
  not g7206 (n_2963, n4505);
  not g7207 (n_2964, n4515);
  and g7208 (n4516, n_2963, n_2964);
  not g7209 (n_2965, n4516);
  and g7210 (n4517, \asqrt[60] , n_2965);
  and g7214 (n4521, n_2747, n_2746);
  and g7215 (n4522, \asqrt[38] , n4521);
  not g7216 (n_2966, n4522);
  and g7217 (n4523, n_2745, n_2966);
  not g7218 (n_2967, n4520);
  not g7219 (n_2968, n4523);
  and g7220 (n4524, n_2967, n_2968);
  and g7221 (n4525, n_162, n_2963);
  and g7222 (n4526, n_2964, n4525);
  not g7223 (n_2969, n4524);
  not g7224 (n_2970, n4526);
  and g7225 (n4527, n_2969, n_2970);
  not g7226 (n_2971, n4517);
  not g7227 (n_2972, n4527);
  and g7228 (n4528, n_2971, n_2972);
  not g7229 (n_2973, n4528);
  and g7230 (n4529, \asqrt[61] , n_2973);
  and g7234 (n4533, n_2755, n_2754);
  and g7235 (n4534, \asqrt[38] , n4533);
  not g7236 (n_2974, n4534);
  and g7237 (n4535, n_2753, n_2974);
  not g7238 (n_2975, n4532);
  not g7239 (n_2976, n4535);
  and g7240 (n4536, n_2975, n_2976);
  and g7241 (n4537, n_115, n_2971);
  and g7242 (n4538, n_2972, n4537);
  not g7243 (n_2977, n4536);
  not g7244 (n_2978, n4538);
  and g7245 (n4539, n_2977, n_2978);
  not g7246 (n_2979, n4529);
  not g7247 (n_2980, n4539);
  and g7248 (n4540, n_2979, n_2980);
  not g7249 (n_2981, n4540);
  and g7250 (n4541, \asqrt[62] , n_2981);
  and g7254 (n4545, n_2763, n_2762);
  and g7255 (n4546, \asqrt[38] , n4545);
  not g7256 (n_2982, n4546);
  and g7257 (n4547, n_2761, n_2982);
  not g7258 (n_2983, n4544);
  not g7259 (n_2984, n4547);
  and g7260 (n4548, n_2983, n_2984);
  and g7261 (n4549, n_76, n_2979);
  and g7262 (n4550, n_2980, n4549);
  not g7263 (n_2985, n4548);
  not g7264 (n_2986, n4550);
  and g7265 (n4551, n_2985, n_2986);
  not g7266 (n_2987, n4541);
  not g7267 (n_2988, n4551);
  and g7268 (n4552, n_2987, n_2988);
  and g7272 (n4556, n_2771, n_2770);
  and g7273 (n4557, \asqrt[38] , n4556);
  not g7274 (n_2989, n4557);
  and g7275 (n4558, n_2769, n_2989);
  not g7276 (n_2990, n4555);
  not g7277 (n_2991, n4558);
  and g7278 (n4559, n_2990, n_2991);
  and g7279 (n4560, n_2778, n_2777);
  and g7280 (n4561, \asqrt[38] , n4560);
  not g7283 (n_2993, n4559);
  not g7285 (n_2994, n4552);
  not g7287 (n_2995, n4564);
  and g7288 (n4565, n_21, n_2995);
  and g7289 (n4566, n_2987, n4559);
  and g7290 (n4567, n_2988, n4566);
  and g7291 (n4568, n_2777, \asqrt[38] );
  not g7292 (n_2996, n4568);
  and g7293 (n4569, n4232, n_2996);
  not g7294 (n_2997, n4560);
  and g7295 (n4570, \asqrt[63] , n_2997);
  not g7296 (n_2998, n4569);
  and g7297 (n4571, n_2998, n4570);
  not g7303 (n_2999, n4571);
  not g7304 (n_3000, n4576);
  not g7306 (n_3001, n4567);
  and g7310 (n4580, \a[74] , \asqrt[37] );
  not g7311 (n_3006, \a[72] );
  not g7312 (n_3007, \a[73] );
  and g7313 (n4581, n_3006, n_3007);
  and g7314 (n4582, n_2790, n4581);
  not g7315 (n_3008, n4580);
  not g7316 (n_3009, n4582);
  and g7317 (n4583, n_3008, n_3009);
  not g7318 (n_3010, n4583);
  and g7319 (n4584, \asqrt[38] , n_3010);
  and g7325 (n4590, n_2790, \asqrt[37] );
  not g7326 (n_3011, n4590);
  and g7327 (n4591, \a[75] , n_3011);
  and g7328 (n4592, n4261, \asqrt[37] );
  not g7329 (n_3012, n4591);
  not g7330 (n_3013, n4592);
  and g7331 (n4593, n_3012, n_3013);
  not g7332 (n_3014, n4589);
  and g7333 (n4594, n_3014, n4593);
  not g7334 (n_3015, n4584);
  not g7335 (n_3016, n4594);
  and g7336 (n4595, n_3015, n_3016);
  not g7337 (n_3017, n4595);
  and g7338 (n4596, \asqrt[39] , n_3017);
  not g7339 (n_3018, \asqrt[39] );
  and g7340 (n4597, n_3018, n_3015);
  and g7341 (n4598, n_3016, n4597);
  not g7345 (n_3019, n4565);
  not g7347 (n_3020, n4602);
  and g7348 (n4603, n_3013, n_3020);
  not g7349 (n_3021, n4603);
  and g7350 (n4604, \a[76] , n_3021);
  and g7351 (n4605, n_2582, n_3020);
  and g7352 (n4606, n_3013, n4605);
  not g7353 (n_3022, n4604);
  not g7354 (n_3023, n4606);
  and g7355 (n4607, n_3022, n_3023);
  not g7356 (n_3024, n4598);
  not g7357 (n_3025, n4607);
  and g7358 (n4608, n_3024, n_3025);
  not g7359 (n_3026, n4596);
  not g7360 (n_3027, n4608);
  and g7361 (n4609, n_3026, n_3027);
  not g7362 (n_3028, n4609);
  and g7363 (n4610, \asqrt[40] , n_3028);
  and g7364 (n4611, n_2799, n_2798);
  not g7365 (n_3029, n4273);
  and g7366 (n4612, n_3029, n4611);
  and g7367 (n4613, \asqrt[37] , n4612);
  and g7368 (n4614, \asqrt[37] , n4611);
  not g7369 (n_3030, n4614);
  and g7370 (n4615, n4273, n_3030);
  not g7371 (n_3031, n4613);
  not g7372 (n_3032, n4615);
  and g7373 (n4616, n_3031, n_3032);
  and g7374 (n4617, n_2802, n_3026);
  and g7375 (n4618, n_3027, n4617);
  not g7376 (n_3033, n4616);
  not g7377 (n_3034, n4618);
  and g7378 (n4619, n_3033, n_3034);
  not g7379 (n_3035, n4610);
  not g7380 (n_3036, n4619);
  and g7381 (n4620, n_3035, n_3036);
  not g7382 (n_3037, n4620);
  and g7383 (n4621, \asqrt[41] , n_3037);
  and g7387 (n4625, n_2810, n_2808);
  and g7388 (n4626, \asqrt[37] , n4625);
  not g7389 (n_3038, n4626);
  and g7390 (n4627, n_2809, n_3038);
  not g7391 (n_3039, n4624);
  not g7392 (n_3040, n4627);
  and g7393 (n4628, n_3039, n_3040);
  and g7394 (n4629, n_2594, n_3035);
  and g7395 (n4630, n_3036, n4629);
  not g7396 (n_3041, n4628);
  not g7397 (n_3042, n4630);
  and g7398 (n4631, n_3041, n_3042);
  not g7399 (n_3043, n4621);
  not g7400 (n_3044, n4631);
  and g7401 (n4632, n_3043, n_3044);
  not g7402 (n_3045, n4632);
  and g7403 (n4633, \asqrt[42] , n_3045);
  and g7407 (n4637, n_2819, n_2818);
  and g7408 (n4638, \asqrt[37] , n4637);
  not g7409 (n_3046, n4638);
  and g7410 (n4639, n_2817, n_3046);
  not g7411 (n_3047, n4636);
  not g7412 (n_3048, n4639);
  and g7413 (n4640, n_3047, n_3048);
  and g7414 (n4641, n_2394, n_3043);
  and g7415 (n4642, n_3044, n4641);
  not g7416 (n_3049, n4640);
  not g7417 (n_3050, n4642);
  and g7418 (n4643, n_3049, n_3050);
  not g7419 (n_3051, n4633);
  not g7420 (n_3052, n4643);
  and g7421 (n4644, n_3051, n_3052);
  not g7422 (n_3053, n4644);
  and g7423 (n4645, \asqrt[43] , n_3053);
  and g7427 (n4649, n_2827, n_2826);
  and g7428 (n4650, \asqrt[37] , n4649);
  not g7429 (n_3054, n4650);
  and g7430 (n4651, n_2825, n_3054);
  not g7431 (n_3055, n4648);
  not g7432 (n_3056, n4651);
  and g7433 (n4652, n_3055, n_3056);
  and g7434 (n4653, n_2202, n_3051);
  and g7435 (n4654, n_3052, n4653);
  not g7436 (n_3057, n4652);
  not g7437 (n_3058, n4654);
  and g7438 (n4655, n_3057, n_3058);
  not g7439 (n_3059, n4645);
  not g7440 (n_3060, n4655);
  and g7441 (n4656, n_3059, n_3060);
  not g7442 (n_3061, n4656);
  and g7443 (n4657, \asqrt[44] , n_3061);
  and g7447 (n4661, n_2835, n_2834);
  and g7448 (n4662, \asqrt[37] , n4661);
  not g7449 (n_3062, n4662);
  and g7450 (n4663, n_2833, n_3062);
  not g7451 (n_3063, n4660);
  not g7452 (n_3064, n4663);
  and g7453 (n4664, n_3063, n_3064);
  and g7454 (n4665, n_2018, n_3059);
  and g7455 (n4666, n_3060, n4665);
  not g7456 (n_3065, n4664);
  not g7457 (n_3066, n4666);
  and g7458 (n4667, n_3065, n_3066);
  not g7459 (n_3067, n4657);
  not g7460 (n_3068, n4667);
  and g7461 (n4668, n_3067, n_3068);
  not g7462 (n_3069, n4668);
  and g7463 (n4669, \asqrt[45] , n_3069);
  and g7467 (n4673, n_2843, n_2842);
  and g7468 (n4674, \asqrt[37] , n4673);
  not g7469 (n_3070, n4674);
  and g7470 (n4675, n_2841, n_3070);
  not g7471 (n_3071, n4672);
  not g7472 (n_3072, n4675);
  and g7473 (n4676, n_3071, n_3072);
  and g7474 (n4677, n_1842, n_3067);
  and g7475 (n4678, n_3068, n4677);
  not g7476 (n_3073, n4676);
  not g7477 (n_3074, n4678);
  and g7478 (n4679, n_3073, n_3074);
  not g7479 (n_3075, n4669);
  not g7480 (n_3076, n4679);
  and g7481 (n4680, n_3075, n_3076);
  not g7482 (n_3077, n4680);
  and g7483 (n4681, \asqrt[46] , n_3077);
  and g7487 (n4685, n_2851, n_2850);
  and g7488 (n4686, \asqrt[37] , n4685);
  not g7489 (n_3078, n4686);
  and g7490 (n4687, n_2849, n_3078);
  not g7491 (n_3079, n4684);
  not g7492 (n_3080, n4687);
  and g7493 (n4688, n_3079, n_3080);
  and g7494 (n4689, n_1674, n_3075);
  and g7495 (n4690, n_3076, n4689);
  not g7496 (n_3081, n4688);
  not g7497 (n_3082, n4690);
  and g7498 (n4691, n_3081, n_3082);
  not g7499 (n_3083, n4681);
  not g7500 (n_3084, n4691);
  and g7501 (n4692, n_3083, n_3084);
  not g7502 (n_3085, n4692);
  and g7503 (n4693, \asqrt[47] , n_3085);
  and g7507 (n4697, n_2859, n_2858);
  and g7508 (n4698, \asqrt[37] , n4697);
  not g7509 (n_3086, n4698);
  and g7510 (n4699, n_2857, n_3086);
  not g7511 (n_3087, n4696);
  not g7512 (n_3088, n4699);
  and g7513 (n4700, n_3087, n_3088);
  and g7514 (n4701, n_1514, n_3083);
  and g7515 (n4702, n_3084, n4701);
  not g7516 (n_3089, n4700);
  not g7517 (n_3090, n4702);
  and g7518 (n4703, n_3089, n_3090);
  not g7519 (n_3091, n4693);
  not g7520 (n_3092, n4703);
  and g7521 (n4704, n_3091, n_3092);
  not g7522 (n_3093, n4704);
  and g7523 (n4705, \asqrt[48] , n_3093);
  and g7527 (n4709, n_2867, n_2866);
  and g7528 (n4710, \asqrt[37] , n4709);
  not g7529 (n_3094, n4710);
  and g7530 (n4711, n_2865, n_3094);
  not g7531 (n_3095, n4708);
  not g7532 (n_3096, n4711);
  and g7533 (n4712, n_3095, n_3096);
  and g7534 (n4713, n_1362, n_3091);
  and g7535 (n4714, n_3092, n4713);
  not g7536 (n_3097, n4712);
  not g7537 (n_3098, n4714);
  and g7538 (n4715, n_3097, n_3098);
  not g7539 (n_3099, n4705);
  not g7540 (n_3100, n4715);
  and g7541 (n4716, n_3099, n_3100);
  not g7542 (n_3101, n4716);
  and g7543 (n4717, \asqrt[49] , n_3101);
  and g7547 (n4721, n_2875, n_2874);
  and g7548 (n4722, \asqrt[37] , n4721);
  not g7549 (n_3102, n4722);
  and g7550 (n4723, n_2873, n_3102);
  not g7551 (n_3103, n4720);
  not g7552 (n_3104, n4723);
  and g7553 (n4724, n_3103, n_3104);
  and g7554 (n4725, n_1218, n_3099);
  and g7555 (n4726, n_3100, n4725);
  not g7556 (n_3105, n4724);
  not g7557 (n_3106, n4726);
  and g7558 (n4727, n_3105, n_3106);
  not g7559 (n_3107, n4717);
  not g7560 (n_3108, n4727);
  and g7561 (n4728, n_3107, n_3108);
  not g7562 (n_3109, n4728);
  and g7563 (n4729, \asqrt[50] , n_3109);
  and g7567 (n4733, n_2883, n_2882);
  and g7568 (n4734, \asqrt[37] , n4733);
  not g7569 (n_3110, n4734);
  and g7570 (n4735, n_2881, n_3110);
  not g7571 (n_3111, n4732);
  not g7572 (n_3112, n4735);
  and g7573 (n4736, n_3111, n_3112);
  and g7574 (n4737, n_1082, n_3107);
  and g7575 (n4738, n_3108, n4737);
  not g7576 (n_3113, n4736);
  not g7577 (n_3114, n4738);
  and g7578 (n4739, n_3113, n_3114);
  not g7579 (n_3115, n4729);
  not g7580 (n_3116, n4739);
  and g7581 (n4740, n_3115, n_3116);
  not g7582 (n_3117, n4740);
  and g7583 (n4741, \asqrt[51] , n_3117);
  and g7587 (n4745, n_2891, n_2890);
  and g7588 (n4746, \asqrt[37] , n4745);
  not g7589 (n_3118, n4746);
  and g7590 (n4747, n_2889, n_3118);
  not g7591 (n_3119, n4744);
  not g7592 (n_3120, n4747);
  and g7593 (n4748, n_3119, n_3120);
  and g7594 (n4749, n_954, n_3115);
  and g7595 (n4750, n_3116, n4749);
  not g7596 (n_3121, n4748);
  not g7597 (n_3122, n4750);
  and g7598 (n4751, n_3121, n_3122);
  not g7599 (n_3123, n4741);
  not g7600 (n_3124, n4751);
  and g7601 (n4752, n_3123, n_3124);
  not g7602 (n_3125, n4752);
  and g7603 (n4753, \asqrt[52] , n_3125);
  and g7607 (n4757, n_2899, n_2898);
  and g7608 (n4758, \asqrt[37] , n4757);
  not g7609 (n_3126, n4758);
  and g7610 (n4759, n_2897, n_3126);
  not g7611 (n_3127, n4756);
  not g7612 (n_3128, n4759);
  and g7613 (n4760, n_3127, n_3128);
  and g7614 (n4761, n_834, n_3123);
  and g7615 (n4762, n_3124, n4761);
  not g7616 (n_3129, n4760);
  not g7617 (n_3130, n4762);
  and g7618 (n4763, n_3129, n_3130);
  not g7619 (n_3131, n4753);
  not g7620 (n_3132, n4763);
  and g7621 (n4764, n_3131, n_3132);
  not g7622 (n_3133, n4764);
  and g7623 (n4765, \asqrt[53] , n_3133);
  and g7627 (n4769, n_2907, n_2906);
  and g7628 (n4770, \asqrt[37] , n4769);
  not g7629 (n_3134, n4770);
  and g7630 (n4771, n_2905, n_3134);
  not g7631 (n_3135, n4768);
  not g7632 (n_3136, n4771);
  and g7633 (n4772, n_3135, n_3136);
  and g7634 (n4773, n_722, n_3131);
  and g7635 (n4774, n_3132, n4773);
  not g7636 (n_3137, n4772);
  not g7637 (n_3138, n4774);
  and g7638 (n4775, n_3137, n_3138);
  not g7639 (n_3139, n4765);
  not g7640 (n_3140, n4775);
  and g7641 (n4776, n_3139, n_3140);
  not g7642 (n_3141, n4776);
  and g7643 (n4777, \asqrt[54] , n_3141);
  and g7647 (n4781, n_2915, n_2914);
  and g7648 (n4782, \asqrt[37] , n4781);
  not g7649 (n_3142, n4782);
  and g7650 (n4783, n_2913, n_3142);
  not g7651 (n_3143, n4780);
  not g7652 (n_3144, n4783);
  and g7653 (n4784, n_3143, n_3144);
  and g7654 (n4785, n_618, n_3139);
  and g7655 (n4786, n_3140, n4785);
  not g7656 (n_3145, n4784);
  not g7657 (n_3146, n4786);
  and g7658 (n4787, n_3145, n_3146);
  not g7659 (n_3147, n4777);
  not g7660 (n_3148, n4787);
  and g7661 (n4788, n_3147, n_3148);
  not g7662 (n_3149, n4788);
  and g7663 (n4789, \asqrt[55] , n_3149);
  and g7667 (n4793, n_2923, n_2922);
  and g7668 (n4794, \asqrt[37] , n4793);
  not g7669 (n_3150, n4794);
  and g7670 (n4795, n_2921, n_3150);
  not g7671 (n_3151, n4792);
  not g7672 (n_3152, n4795);
  and g7673 (n4796, n_3151, n_3152);
  and g7674 (n4797, n_522, n_3147);
  and g7675 (n4798, n_3148, n4797);
  not g7676 (n_3153, n4796);
  not g7677 (n_3154, n4798);
  and g7678 (n4799, n_3153, n_3154);
  not g7679 (n_3155, n4789);
  not g7680 (n_3156, n4799);
  and g7681 (n4800, n_3155, n_3156);
  not g7682 (n_3157, n4800);
  and g7683 (n4801, \asqrt[56] , n_3157);
  and g7687 (n4805, n_2931, n_2930);
  and g7688 (n4806, \asqrt[37] , n4805);
  not g7689 (n_3158, n4806);
  and g7690 (n4807, n_2929, n_3158);
  not g7691 (n_3159, n4804);
  not g7692 (n_3160, n4807);
  and g7693 (n4808, n_3159, n_3160);
  and g7694 (n4809, n_434, n_3155);
  and g7695 (n4810, n_3156, n4809);
  not g7696 (n_3161, n4808);
  not g7697 (n_3162, n4810);
  and g7698 (n4811, n_3161, n_3162);
  not g7699 (n_3163, n4801);
  not g7700 (n_3164, n4811);
  and g7701 (n4812, n_3163, n_3164);
  not g7702 (n_3165, n4812);
  and g7703 (n4813, \asqrt[57] , n_3165);
  and g7707 (n4817, n_2939, n_2938);
  and g7708 (n4818, \asqrt[37] , n4817);
  not g7709 (n_3166, n4818);
  and g7710 (n4819, n_2937, n_3166);
  not g7711 (n_3167, n4816);
  not g7712 (n_3168, n4819);
  and g7713 (n4820, n_3167, n_3168);
  and g7714 (n4821, n_354, n_3163);
  and g7715 (n4822, n_3164, n4821);
  not g7716 (n_3169, n4820);
  not g7717 (n_3170, n4822);
  and g7718 (n4823, n_3169, n_3170);
  not g7719 (n_3171, n4813);
  not g7720 (n_3172, n4823);
  and g7721 (n4824, n_3171, n_3172);
  not g7722 (n_3173, n4824);
  and g7723 (n4825, \asqrt[58] , n_3173);
  and g7727 (n4829, n_2947, n_2946);
  and g7728 (n4830, \asqrt[37] , n4829);
  not g7729 (n_3174, n4830);
  and g7730 (n4831, n_2945, n_3174);
  not g7731 (n_3175, n4828);
  not g7732 (n_3176, n4831);
  and g7733 (n4832, n_3175, n_3176);
  and g7734 (n4833, n_282, n_3171);
  and g7735 (n4834, n_3172, n4833);
  not g7736 (n_3177, n4832);
  not g7737 (n_3178, n4834);
  and g7738 (n4835, n_3177, n_3178);
  not g7739 (n_3179, n4825);
  not g7740 (n_3180, n4835);
  and g7741 (n4836, n_3179, n_3180);
  not g7742 (n_3181, n4836);
  and g7743 (n4837, \asqrt[59] , n_3181);
  and g7747 (n4841, n_2955, n_2954);
  and g7748 (n4842, \asqrt[37] , n4841);
  not g7749 (n_3182, n4842);
  and g7750 (n4843, n_2953, n_3182);
  not g7751 (n_3183, n4840);
  not g7752 (n_3184, n4843);
  and g7753 (n4844, n_3183, n_3184);
  and g7754 (n4845, n_218, n_3179);
  and g7755 (n4846, n_3180, n4845);
  not g7756 (n_3185, n4844);
  not g7757 (n_3186, n4846);
  and g7758 (n4847, n_3185, n_3186);
  not g7759 (n_3187, n4837);
  not g7760 (n_3188, n4847);
  and g7761 (n4848, n_3187, n_3188);
  not g7762 (n_3189, n4848);
  and g7763 (n4849, \asqrt[60] , n_3189);
  and g7764 (n4850, n_162, n_3187);
  and g7765 (n4851, n_3188, n4850);
  and g7769 (n4855, n_2963, n_2961);
  and g7770 (n4856, \asqrt[37] , n4855);
  not g7771 (n_3190, n4856);
  and g7772 (n4857, n_2962, n_3190);
  not g7773 (n_3191, n4854);
  not g7774 (n_3192, n4857);
  and g7775 (n4858, n_3191, n_3192);
  not g7776 (n_3193, n4851);
  not g7777 (n_3194, n4858);
  and g7778 (n4859, n_3193, n_3194);
  not g7779 (n_3195, n4849);
  not g7780 (n_3196, n4859);
  and g7781 (n4860, n_3195, n_3196);
  not g7782 (n_3197, n4860);
  and g7783 (n4861, \asqrt[61] , n_3197);
  and g7787 (n4865, n_2971, n_2970);
  and g7788 (n4866, \asqrt[37] , n4865);
  not g7789 (n_3198, n4866);
  and g7790 (n4867, n_2969, n_3198);
  not g7791 (n_3199, n4864);
  not g7792 (n_3200, n4867);
  and g7793 (n4868, n_3199, n_3200);
  and g7794 (n4869, n_115, n_3195);
  and g7795 (n4870, n_3196, n4869);
  not g7796 (n_3201, n4868);
  not g7797 (n_3202, n4870);
  and g7798 (n4871, n_3201, n_3202);
  not g7799 (n_3203, n4861);
  not g7800 (n_3204, n4871);
  and g7801 (n4872, n_3203, n_3204);
  not g7802 (n_3205, n4872);
  and g7803 (n4873, \asqrt[62] , n_3205);
  and g7807 (n4877, n_2979, n_2978);
  and g7808 (n4878, \asqrt[37] , n4877);
  not g7809 (n_3206, n4878);
  and g7810 (n4879, n_2977, n_3206);
  not g7811 (n_3207, n4876);
  not g7812 (n_3208, n4879);
  and g7813 (n4880, n_3207, n_3208);
  and g7814 (n4881, n_76, n_3203);
  and g7815 (n4882, n_3204, n4881);
  not g7816 (n_3209, n4880);
  not g7817 (n_3210, n4882);
  and g7818 (n4883, n_3209, n_3210);
  not g7819 (n_3211, n4873);
  not g7820 (n_3212, n4883);
  and g7821 (n4884, n_3211, n_3212);
  and g7825 (n4888, n_2987, n_2986);
  and g7826 (n4889, \asqrt[37] , n4888);
  not g7827 (n_3213, n4889);
  and g7828 (n4890, n_2985, n_3213);
  not g7829 (n_3214, n4887);
  not g7830 (n_3215, n4890);
  and g7831 (n4891, n_3214, n_3215);
  and g7832 (n4892, n_2994, n_2993);
  and g7833 (n4893, \asqrt[37] , n4892);
  not g7836 (n_3217, n4891);
  not g7838 (n_3218, n4884);
  not g7840 (n_3219, n4896);
  and g7841 (n4897, n_21, n_3219);
  and g7842 (n4898, n_3211, n4891);
  and g7843 (n4899, n_3212, n4898);
  and g7844 (n4900, n_2993, \asqrt[37] );
  not g7845 (n_3220, n4900);
  and g7846 (n4901, n4552, n_3220);
  not g7847 (n_3221, n4892);
  and g7848 (n4902, \asqrt[63] , n_3221);
  not g7849 (n_3222, n4901);
  and g7850 (n4903, n_3222, n4902);
  not g7856 (n_3223, n4903);
  not g7857 (n_3224, n4908);
  not g7859 (n_3225, n4899);
  and g7863 (n4912, \a[72] , \asqrt[36] );
  not g7864 (n_3230, \a[70] );
  not g7865 (n_3231, \a[71] );
  and g7866 (n4913, n_3230, n_3231);
  and g7867 (n4914, n_3006, n4913);
  not g7868 (n_3232, n4912);
  not g7869 (n_3233, n4914);
  and g7870 (n4915, n_3232, n_3233);
  not g7871 (n_3234, n4915);
  and g7872 (n4916, \asqrt[37] , n_3234);
  and g7878 (n4922, n_3006, \asqrt[36] );
  not g7879 (n_3235, n4922);
  and g7880 (n4923, \a[73] , n_3235);
  and g7881 (n4924, n4581, \asqrt[36] );
  not g7882 (n_3236, n4923);
  not g7883 (n_3237, n4924);
  and g7884 (n4925, n_3236, n_3237);
  not g7885 (n_3238, n4921);
  and g7886 (n4926, n_3238, n4925);
  not g7887 (n_3239, n4916);
  not g7888 (n_3240, n4926);
  and g7889 (n4927, n_3239, n_3240);
  not g7890 (n_3241, n4927);
  and g7891 (n4928, \asqrt[38] , n_3241);
  not g7892 (n_3242, \asqrt[38] );
  and g7893 (n4929, n_3242, n_3239);
  and g7894 (n4930, n_3240, n4929);
  not g7898 (n_3243, n4897);
  not g7900 (n_3244, n4934);
  and g7901 (n4935, n_3237, n_3244);
  not g7902 (n_3245, n4935);
  and g7903 (n4936, \a[74] , n_3245);
  and g7904 (n4937, n_2790, n_3244);
  and g7905 (n4938, n_3237, n4937);
  not g7906 (n_3246, n4936);
  not g7907 (n_3247, n4938);
  and g7908 (n4939, n_3246, n_3247);
  not g7909 (n_3248, n4930);
  not g7910 (n_3249, n4939);
  and g7911 (n4940, n_3248, n_3249);
  not g7912 (n_3250, n4928);
  not g7913 (n_3251, n4940);
  and g7914 (n4941, n_3250, n_3251);
  not g7915 (n_3252, n4941);
  and g7916 (n4942, \asqrt[39] , n_3252);
  and g7917 (n4943, n_3015, n_3014);
  not g7918 (n_3253, n4593);
  and g7919 (n4944, n_3253, n4943);
  and g7920 (n4945, \asqrt[36] , n4944);
  and g7921 (n4946, \asqrt[36] , n4943);
  not g7922 (n_3254, n4946);
  and g7923 (n4947, n4593, n_3254);
  not g7924 (n_3255, n4945);
  not g7925 (n_3256, n4947);
  and g7926 (n4948, n_3255, n_3256);
  and g7927 (n4949, n_3018, n_3250);
  and g7928 (n4950, n_3251, n4949);
  not g7929 (n_3257, n4948);
  not g7930 (n_3258, n4950);
  and g7931 (n4951, n_3257, n_3258);
  not g7932 (n_3259, n4942);
  not g7933 (n_3260, n4951);
  and g7934 (n4952, n_3259, n_3260);
  not g7935 (n_3261, n4952);
  and g7936 (n4953, \asqrt[40] , n_3261);
  and g7940 (n4957, n_3026, n_3024);
  and g7941 (n4958, \asqrt[36] , n4957);
  not g7942 (n_3262, n4958);
  and g7943 (n4959, n_3025, n_3262);
  not g7944 (n_3263, n4956);
  not g7945 (n_3264, n4959);
  and g7946 (n4960, n_3263, n_3264);
  and g7947 (n4961, n_2802, n_3259);
  and g7948 (n4962, n_3260, n4961);
  not g7949 (n_3265, n4960);
  not g7950 (n_3266, n4962);
  and g7951 (n4963, n_3265, n_3266);
  not g7952 (n_3267, n4953);
  not g7953 (n_3268, n4963);
  and g7954 (n4964, n_3267, n_3268);
  not g7955 (n_3269, n4964);
  and g7956 (n4965, \asqrt[41] , n_3269);
  and g7960 (n4969, n_3035, n_3034);
  and g7961 (n4970, \asqrt[36] , n4969);
  not g7962 (n_3270, n4970);
  and g7963 (n4971, n_3033, n_3270);
  not g7964 (n_3271, n4968);
  not g7965 (n_3272, n4971);
  and g7966 (n4972, n_3271, n_3272);
  and g7967 (n4973, n_2594, n_3267);
  and g7968 (n4974, n_3268, n4973);
  not g7969 (n_3273, n4972);
  not g7970 (n_3274, n4974);
  and g7971 (n4975, n_3273, n_3274);
  not g7972 (n_3275, n4965);
  not g7973 (n_3276, n4975);
  and g7974 (n4976, n_3275, n_3276);
  not g7975 (n_3277, n4976);
  and g7976 (n4977, \asqrt[42] , n_3277);
  and g7980 (n4981, n_3043, n_3042);
  and g7981 (n4982, \asqrt[36] , n4981);
  not g7982 (n_3278, n4982);
  and g7983 (n4983, n_3041, n_3278);
  not g7984 (n_3279, n4980);
  not g7985 (n_3280, n4983);
  and g7986 (n4984, n_3279, n_3280);
  and g7987 (n4985, n_2394, n_3275);
  and g7988 (n4986, n_3276, n4985);
  not g7989 (n_3281, n4984);
  not g7990 (n_3282, n4986);
  and g7991 (n4987, n_3281, n_3282);
  not g7992 (n_3283, n4977);
  not g7993 (n_3284, n4987);
  and g7994 (n4988, n_3283, n_3284);
  not g7995 (n_3285, n4988);
  and g7996 (n4989, \asqrt[43] , n_3285);
  and g8000 (n4993, n_3051, n_3050);
  and g8001 (n4994, \asqrt[36] , n4993);
  not g8002 (n_3286, n4994);
  and g8003 (n4995, n_3049, n_3286);
  not g8004 (n_3287, n4992);
  not g8005 (n_3288, n4995);
  and g8006 (n4996, n_3287, n_3288);
  and g8007 (n4997, n_2202, n_3283);
  and g8008 (n4998, n_3284, n4997);
  not g8009 (n_3289, n4996);
  not g8010 (n_3290, n4998);
  and g8011 (n4999, n_3289, n_3290);
  not g8012 (n_3291, n4989);
  not g8013 (n_3292, n4999);
  and g8014 (n5000, n_3291, n_3292);
  not g8015 (n_3293, n5000);
  and g8016 (n5001, \asqrt[44] , n_3293);
  and g8020 (n5005, n_3059, n_3058);
  and g8021 (n5006, \asqrt[36] , n5005);
  not g8022 (n_3294, n5006);
  and g8023 (n5007, n_3057, n_3294);
  not g8024 (n_3295, n5004);
  not g8025 (n_3296, n5007);
  and g8026 (n5008, n_3295, n_3296);
  and g8027 (n5009, n_2018, n_3291);
  and g8028 (n5010, n_3292, n5009);
  not g8029 (n_3297, n5008);
  not g8030 (n_3298, n5010);
  and g8031 (n5011, n_3297, n_3298);
  not g8032 (n_3299, n5001);
  not g8033 (n_3300, n5011);
  and g8034 (n5012, n_3299, n_3300);
  not g8035 (n_3301, n5012);
  and g8036 (n5013, \asqrt[45] , n_3301);
  and g8040 (n5017, n_3067, n_3066);
  and g8041 (n5018, \asqrt[36] , n5017);
  not g8042 (n_3302, n5018);
  and g8043 (n5019, n_3065, n_3302);
  not g8044 (n_3303, n5016);
  not g8045 (n_3304, n5019);
  and g8046 (n5020, n_3303, n_3304);
  and g8047 (n5021, n_1842, n_3299);
  and g8048 (n5022, n_3300, n5021);
  not g8049 (n_3305, n5020);
  not g8050 (n_3306, n5022);
  and g8051 (n5023, n_3305, n_3306);
  not g8052 (n_3307, n5013);
  not g8053 (n_3308, n5023);
  and g8054 (n5024, n_3307, n_3308);
  not g8055 (n_3309, n5024);
  and g8056 (n5025, \asqrt[46] , n_3309);
  and g8060 (n5029, n_3075, n_3074);
  and g8061 (n5030, \asqrt[36] , n5029);
  not g8062 (n_3310, n5030);
  and g8063 (n5031, n_3073, n_3310);
  not g8064 (n_3311, n5028);
  not g8065 (n_3312, n5031);
  and g8066 (n5032, n_3311, n_3312);
  and g8067 (n5033, n_1674, n_3307);
  and g8068 (n5034, n_3308, n5033);
  not g8069 (n_3313, n5032);
  not g8070 (n_3314, n5034);
  and g8071 (n5035, n_3313, n_3314);
  not g8072 (n_3315, n5025);
  not g8073 (n_3316, n5035);
  and g8074 (n5036, n_3315, n_3316);
  not g8075 (n_3317, n5036);
  and g8076 (n5037, \asqrt[47] , n_3317);
  and g8080 (n5041, n_3083, n_3082);
  and g8081 (n5042, \asqrt[36] , n5041);
  not g8082 (n_3318, n5042);
  and g8083 (n5043, n_3081, n_3318);
  not g8084 (n_3319, n5040);
  not g8085 (n_3320, n5043);
  and g8086 (n5044, n_3319, n_3320);
  and g8087 (n5045, n_1514, n_3315);
  and g8088 (n5046, n_3316, n5045);
  not g8089 (n_3321, n5044);
  not g8090 (n_3322, n5046);
  and g8091 (n5047, n_3321, n_3322);
  not g8092 (n_3323, n5037);
  not g8093 (n_3324, n5047);
  and g8094 (n5048, n_3323, n_3324);
  not g8095 (n_3325, n5048);
  and g8096 (n5049, \asqrt[48] , n_3325);
  and g8100 (n5053, n_3091, n_3090);
  and g8101 (n5054, \asqrt[36] , n5053);
  not g8102 (n_3326, n5054);
  and g8103 (n5055, n_3089, n_3326);
  not g8104 (n_3327, n5052);
  not g8105 (n_3328, n5055);
  and g8106 (n5056, n_3327, n_3328);
  and g8107 (n5057, n_1362, n_3323);
  and g8108 (n5058, n_3324, n5057);
  not g8109 (n_3329, n5056);
  not g8110 (n_3330, n5058);
  and g8111 (n5059, n_3329, n_3330);
  not g8112 (n_3331, n5049);
  not g8113 (n_3332, n5059);
  and g8114 (n5060, n_3331, n_3332);
  not g8115 (n_3333, n5060);
  and g8116 (n5061, \asqrt[49] , n_3333);
  and g8120 (n5065, n_3099, n_3098);
  and g8121 (n5066, \asqrt[36] , n5065);
  not g8122 (n_3334, n5066);
  and g8123 (n5067, n_3097, n_3334);
  not g8124 (n_3335, n5064);
  not g8125 (n_3336, n5067);
  and g8126 (n5068, n_3335, n_3336);
  and g8127 (n5069, n_1218, n_3331);
  and g8128 (n5070, n_3332, n5069);
  not g8129 (n_3337, n5068);
  not g8130 (n_3338, n5070);
  and g8131 (n5071, n_3337, n_3338);
  not g8132 (n_3339, n5061);
  not g8133 (n_3340, n5071);
  and g8134 (n5072, n_3339, n_3340);
  not g8135 (n_3341, n5072);
  and g8136 (n5073, \asqrt[50] , n_3341);
  and g8140 (n5077, n_3107, n_3106);
  and g8141 (n5078, \asqrt[36] , n5077);
  not g8142 (n_3342, n5078);
  and g8143 (n5079, n_3105, n_3342);
  not g8144 (n_3343, n5076);
  not g8145 (n_3344, n5079);
  and g8146 (n5080, n_3343, n_3344);
  and g8147 (n5081, n_1082, n_3339);
  and g8148 (n5082, n_3340, n5081);
  not g8149 (n_3345, n5080);
  not g8150 (n_3346, n5082);
  and g8151 (n5083, n_3345, n_3346);
  not g8152 (n_3347, n5073);
  not g8153 (n_3348, n5083);
  and g8154 (n5084, n_3347, n_3348);
  not g8155 (n_3349, n5084);
  and g8156 (n5085, \asqrt[51] , n_3349);
  and g8160 (n5089, n_3115, n_3114);
  and g8161 (n5090, \asqrt[36] , n5089);
  not g8162 (n_3350, n5090);
  and g8163 (n5091, n_3113, n_3350);
  not g8164 (n_3351, n5088);
  not g8165 (n_3352, n5091);
  and g8166 (n5092, n_3351, n_3352);
  and g8167 (n5093, n_954, n_3347);
  and g8168 (n5094, n_3348, n5093);
  not g8169 (n_3353, n5092);
  not g8170 (n_3354, n5094);
  and g8171 (n5095, n_3353, n_3354);
  not g8172 (n_3355, n5085);
  not g8173 (n_3356, n5095);
  and g8174 (n5096, n_3355, n_3356);
  not g8175 (n_3357, n5096);
  and g8176 (n5097, \asqrt[52] , n_3357);
  and g8180 (n5101, n_3123, n_3122);
  and g8181 (n5102, \asqrt[36] , n5101);
  not g8182 (n_3358, n5102);
  and g8183 (n5103, n_3121, n_3358);
  not g8184 (n_3359, n5100);
  not g8185 (n_3360, n5103);
  and g8186 (n5104, n_3359, n_3360);
  and g8187 (n5105, n_834, n_3355);
  and g8188 (n5106, n_3356, n5105);
  not g8189 (n_3361, n5104);
  not g8190 (n_3362, n5106);
  and g8191 (n5107, n_3361, n_3362);
  not g8192 (n_3363, n5097);
  not g8193 (n_3364, n5107);
  and g8194 (n5108, n_3363, n_3364);
  not g8195 (n_3365, n5108);
  and g8196 (n5109, \asqrt[53] , n_3365);
  and g8200 (n5113, n_3131, n_3130);
  and g8201 (n5114, \asqrt[36] , n5113);
  not g8202 (n_3366, n5114);
  and g8203 (n5115, n_3129, n_3366);
  not g8204 (n_3367, n5112);
  not g8205 (n_3368, n5115);
  and g8206 (n5116, n_3367, n_3368);
  and g8207 (n5117, n_722, n_3363);
  and g8208 (n5118, n_3364, n5117);
  not g8209 (n_3369, n5116);
  not g8210 (n_3370, n5118);
  and g8211 (n5119, n_3369, n_3370);
  not g8212 (n_3371, n5109);
  not g8213 (n_3372, n5119);
  and g8214 (n5120, n_3371, n_3372);
  not g8215 (n_3373, n5120);
  and g8216 (n5121, \asqrt[54] , n_3373);
  and g8220 (n5125, n_3139, n_3138);
  and g8221 (n5126, \asqrt[36] , n5125);
  not g8222 (n_3374, n5126);
  and g8223 (n5127, n_3137, n_3374);
  not g8224 (n_3375, n5124);
  not g8225 (n_3376, n5127);
  and g8226 (n5128, n_3375, n_3376);
  and g8227 (n5129, n_618, n_3371);
  and g8228 (n5130, n_3372, n5129);
  not g8229 (n_3377, n5128);
  not g8230 (n_3378, n5130);
  and g8231 (n5131, n_3377, n_3378);
  not g8232 (n_3379, n5121);
  not g8233 (n_3380, n5131);
  and g8234 (n5132, n_3379, n_3380);
  not g8235 (n_3381, n5132);
  and g8236 (n5133, \asqrt[55] , n_3381);
  and g8240 (n5137, n_3147, n_3146);
  and g8241 (n5138, \asqrt[36] , n5137);
  not g8242 (n_3382, n5138);
  and g8243 (n5139, n_3145, n_3382);
  not g8244 (n_3383, n5136);
  not g8245 (n_3384, n5139);
  and g8246 (n5140, n_3383, n_3384);
  and g8247 (n5141, n_522, n_3379);
  and g8248 (n5142, n_3380, n5141);
  not g8249 (n_3385, n5140);
  not g8250 (n_3386, n5142);
  and g8251 (n5143, n_3385, n_3386);
  not g8252 (n_3387, n5133);
  not g8253 (n_3388, n5143);
  and g8254 (n5144, n_3387, n_3388);
  not g8255 (n_3389, n5144);
  and g8256 (n5145, \asqrt[56] , n_3389);
  and g8260 (n5149, n_3155, n_3154);
  and g8261 (n5150, \asqrt[36] , n5149);
  not g8262 (n_3390, n5150);
  and g8263 (n5151, n_3153, n_3390);
  not g8264 (n_3391, n5148);
  not g8265 (n_3392, n5151);
  and g8266 (n5152, n_3391, n_3392);
  and g8267 (n5153, n_434, n_3387);
  and g8268 (n5154, n_3388, n5153);
  not g8269 (n_3393, n5152);
  not g8270 (n_3394, n5154);
  and g8271 (n5155, n_3393, n_3394);
  not g8272 (n_3395, n5145);
  not g8273 (n_3396, n5155);
  and g8274 (n5156, n_3395, n_3396);
  not g8275 (n_3397, n5156);
  and g8276 (n5157, \asqrt[57] , n_3397);
  and g8280 (n5161, n_3163, n_3162);
  and g8281 (n5162, \asqrt[36] , n5161);
  not g8282 (n_3398, n5162);
  and g8283 (n5163, n_3161, n_3398);
  not g8284 (n_3399, n5160);
  not g8285 (n_3400, n5163);
  and g8286 (n5164, n_3399, n_3400);
  and g8287 (n5165, n_354, n_3395);
  and g8288 (n5166, n_3396, n5165);
  not g8289 (n_3401, n5164);
  not g8290 (n_3402, n5166);
  and g8291 (n5167, n_3401, n_3402);
  not g8292 (n_3403, n5157);
  not g8293 (n_3404, n5167);
  and g8294 (n5168, n_3403, n_3404);
  not g8295 (n_3405, n5168);
  and g8296 (n5169, \asqrt[58] , n_3405);
  and g8300 (n5173, n_3171, n_3170);
  and g8301 (n5174, \asqrt[36] , n5173);
  not g8302 (n_3406, n5174);
  and g8303 (n5175, n_3169, n_3406);
  not g8304 (n_3407, n5172);
  not g8305 (n_3408, n5175);
  and g8306 (n5176, n_3407, n_3408);
  and g8307 (n5177, n_282, n_3403);
  and g8308 (n5178, n_3404, n5177);
  not g8309 (n_3409, n5176);
  not g8310 (n_3410, n5178);
  and g8311 (n5179, n_3409, n_3410);
  not g8312 (n_3411, n5169);
  not g8313 (n_3412, n5179);
  and g8314 (n5180, n_3411, n_3412);
  not g8315 (n_3413, n5180);
  and g8316 (n5181, \asqrt[59] , n_3413);
  and g8320 (n5185, n_3179, n_3178);
  and g8321 (n5186, \asqrt[36] , n5185);
  not g8322 (n_3414, n5186);
  and g8323 (n5187, n_3177, n_3414);
  not g8324 (n_3415, n5184);
  not g8325 (n_3416, n5187);
  and g8326 (n5188, n_3415, n_3416);
  and g8327 (n5189, n_218, n_3411);
  and g8328 (n5190, n_3412, n5189);
  not g8329 (n_3417, n5188);
  not g8330 (n_3418, n5190);
  and g8331 (n5191, n_3417, n_3418);
  not g8332 (n_3419, n5181);
  not g8333 (n_3420, n5191);
  and g8334 (n5192, n_3419, n_3420);
  not g8335 (n_3421, n5192);
  and g8336 (n5193, \asqrt[60] , n_3421);
  and g8340 (n5197, n_3187, n_3186);
  and g8341 (n5198, \asqrt[36] , n5197);
  not g8342 (n_3422, n5198);
  and g8343 (n5199, n_3185, n_3422);
  not g8344 (n_3423, n5196);
  not g8345 (n_3424, n5199);
  and g8346 (n5200, n_3423, n_3424);
  and g8347 (n5201, n_162, n_3419);
  and g8348 (n5202, n_3420, n5201);
  not g8349 (n_3425, n5200);
  not g8350 (n_3426, n5202);
  and g8351 (n5203, n_3425, n_3426);
  not g8352 (n_3427, n5193);
  not g8353 (n_3428, n5203);
  and g8354 (n5204, n_3427, n_3428);
  not g8355 (n_3429, n5204);
  and g8356 (n5205, \asqrt[61] , n_3429);
  and g8357 (n5206, n_115, n_3427);
  and g8358 (n5207, n_3428, n5206);
  and g8362 (n5211, n_3195, n_3193);
  and g8363 (n5212, \asqrt[36] , n5211);
  not g8364 (n_3430, n5212);
  and g8365 (n5213, n_3194, n_3430);
  not g8366 (n_3431, n5210);
  not g8367 (n_3432, n5213);
  and g8368 (n5214, n_3431, n_3432);
  not g8369 (n_3433, n5207);
  not g8370 (n_3434, n5214);
  and g8371 (n5215, n_3433, n_3434);
  not g8372 (n_3435, n5205);
  not g8373 (n_3436, n5215);
  and g8374 (n5216, n_3435, n_3436);
  not g8375 (n_3437, n5216);
  and g8376 (n5217, \asqrt[62] , n_3437);
  and g8380 (n5221, n_3203, n_3202);
  and g8381 (n5222, \asqrt[36] , n5221);
  not g8382 (n_3438, n5222);
  and g8383 (n5223, n_3201, n_3438);
  not g8384 (n_3439, n5220);
  not g8385 (n_3440, n5223);
  and g8386 (n5224, n_3439, n_3440);
  and g8387 (n5225, n_76, n_3435);
  and g8388 (n5226, n_3436, n5225);
  not g8389 (n_3441, n5224);
  not g8390 (n_3442, n5226);
  and g8391 (n5227, n_3441, n_3442);
  not g8392 (n_3443, n5217);
  not g8393 (n_3444, n5227);
  and g8394 (n5228, n_3443, n_3444);
  and g8398 (n5232, n_3211, n_3210);
  and g8399 (n5233, \asqrt[36] , n5232);
  not g8400 (n_3445, n5233);
  and g8401 (n5234, n_3209, n_3445);
  not g8402 (n_3446, n5231);
  not g8403 (n_3447, n5234);
  and g8404 (n5235, n_3446, n_3447);
  and g8405 (n5236, n_3218, n_3217);
  and g8406 (n5237, \asqrt[36] , n5236);
  not g8409 (n_3449, n5235);
  not g8411 (n_3450, n5228);
  not g8413 (n_3451, n5240);
  and g8414 (n5241, n_21, n_3451);
  and g8415 (n5242, n_3443, n5235);
  and g8416 (n5243, n_3444, n5242);
  and g8417 (n5244, n_3217, \asqrt[36] );
  not g8418 (n_3452, n5244);
  and g8419 (n5245, n4884, n_3452);
  not g8420 (n_3453, n5236);
  and g8421 (n5246, \asqrt[63] , n_3453);
  not g8422 (n_3454, n5245);
  and g8423 (n5247, n_3454, n5246);
  not g8429 (n_3455, n5247);
  not g8430 (n_3456, n5252);
  not g8432 (n_3457, n5243);
  and g8436 (n5256, \a[70] , \asqrt[35] );
  not g8437 (n_3462, \a[68] );
  not g8438 (n_3463, \a[69] );
  and g8439 (n5257, n_3462, n_3463);
  and g8440 (n5258, n_3230, n5257);
  not g8441 (n_3464, n5256);
  not g8442 (n_3465, n5258);
  and g8443 (n5259, n_3464, n_3465);
  not g8444 (n_3466, n5259);
  and g8445 (n5260, \asqrt[36] , n_3466);
  and g8451 (n5266, n_3230, \asqrt[35] );
  not g8452 (n_3467, n5266);
  and g8453 (n5267, \a[71] , n_3467);
  and g8454 (n5268, n4913, \asqrt[35] );
  not g8455 (n_3468, n5267);
  not g8456 (n_3469, n5268);
  and g8457 (n5269, n_3468, n_3469);
  not g8458 (n_3470, n5265);
  and g8459 (n5270, n_3470, n5269);
  not g8460 (n_3471, n5260);
  not g8461 (n_3472, n5270);
  and g8462 (n5271, n_3471, n_3472);
  not g8463 (n_3473, n5271);
  and g8464 (n5272, \asqrt[37] , n_3473);
  not g8465 (n_3474, \asqrt[37] );
  and g8466 (n5273, n_3474, n_3471);
  and g8467 (n5274, n_3472, n5273);
  not g8471 (n_3475, n5241);
  not g8473 (n_3476, n5278);
  and g8474 (n5279, n_3469, n_3476);
  not g8475 (n_3477, n5279);
  and g8476 (n5280, \a[72] , n_3477);
  and g8477 (n5281, n_3006, n_3476);
  and g8478 (n5282, n_3469, n5281);
  not g8479 (n_3478, n5280);
  not g8480 (n_3479, n5282);
  and g8481 (n5283, n_3478, n_3479);
  not g8482 (n_3480, n5274);
  not g8483 (n_3481, n5283);
  and g8484 (n5284, n_3480, n_3481);
  not g8485 (n_3482, n5272);
  not g8486 (n_3483, n5284);
  and g8487 (n5285, n_3482, n_3483);
  not g8488 (n_3484, n5285);
  and g8489 (n5286, \asqrt[38] , n_3484);
  and g8490 (n5287, n_3239, n_3238);
  not g8491 (n_3485, n4925);
  and g8492 (n5288, n_3485, n5287);
  and g8493 (n5289, \asqrt[35] , n5288);
  and g8494 (n5290, \asqrt[35] , n5287);
  not g8495 (n_3486, n5290);
  and g8496 (n5291, n4925, n_3486);
  not g8497 (n_3487, n5289);
  not g8498 (n_3488, n5291);
  and g8499 (n5292, n_3487, n_3488);
  and g8500 (n5293, n_3242, n_3482);
  and g8501 (n5294, n_3483, n5293);
  not g8502 (n_3489, n5292);
  not g8503 (n_3490, n5294);
  and g8504 (n5295, n_3489, n_3490);
  not g8505 (n_3491, n5286);
  not g8506 (n_3492, n5295);
  and g8507 (n5296, n_3491, n_3492);
  not g8508 (n_3493, n5296);
  and g8509 (n5297, \asqrt[39] , n_3493);
  and g8513 (n5301, n_3250, n_3248);
  and g8514 (n5302, \asqrt[35] , n5301);
  not g8515 (n_3494, n5302);
  and g8516 (n5303, n_3249, n_3494);
  not g8517 (n_3495, n5300);
  not g8518 (n_3496, n5303);
  and g8519 (n5304, n_3495, n_3496);
  and g8520 (n5305, n_3018, n_3491);
  and g8521 (n5306, n_3492, n5305);
  not g8522 (n_3497, n5304);
  not g8523 (n_3498, n5306);
  and g8524 (n5307, n_3497, n_3498);
  not g8525 (n_3499, n5297);
  not g8526 (n_3500, n5307);
  and g8527 (n5308, n_3499, n_3500);
  not g8528 (n_3501, n5308);
  and g8529 (n5309, \asqrt[40] , n_3501);
  and g8533 (n5313, n_3259, n_3258);
  and g8534 (n5314, \asqrt[35] , n5313);
  not g8535 (n_3502, n5314);
  and g8536 (n5315, n_3257, n_3502);
  not g8537 (n_3503, n5312);
  not g8538 (n_3504, n5315);
  and g8539 (n5316, n_3503, n_3504);
  and g8540 (n5317, n_2802, n_3499);
  and g8541 (n5318, n_3500, n5317);
  not g8542 (n_3505, n5316);
  not g8543 (n_3506, n5318);
  and g8544 (n5319, n_3505, n_3506);
  not g8545 (n_3507, n5309);
  not g8546 (n_3508, n5319);
  and g8547 (n5320, n_3507, n_3508);
  not g8548 (n_3509, n5320);
  and g8549 (n5321, \asqrt[41] , n_3509);
  and g8553 (n5325, n_3267, n_3266);
  and g8554 (n5326, \asqrt[35] , n5325);
  not g8555 (n_3510, n5326);
  and g8556 (n5327, n_3265, n_3510);
  not g8557 (n_3511, n5324);
  not g8558 (n_3512, n5327);
  and g8559 (n5328, n_3511, n_3512);
  and g8560 (n5329, n_2594, n_3507);
  and g8561 (n5330, n_3508, n5329);
  not g8562 (n_3513, n5328);
  not g8563 (n_3514, n5330);
  and g8564 (n5331, n_3513, n_3514);
  not g8565 (n_3515, n5321);
  not g8566 (n_3516, n5331);
  and g8567 (n5332, n_3515, n_3516);
  not g8568 (n_3517, n5332);
  and g8569 (n5333, \asqrt[42] , n_3517);
  and g8573 (n5337, n_3275, n_3274);
  and g8574 (n5338, \asqrt[35] , n5337);
  not g8575 (n_3518, n5338);
  and g8576 (n5339, n_3273, n_3518);
  not g8577 (n_3519, n5336);
  not g8578 (n_3520, n5339);
  and g8579 (n5340, n_3519, n_3520);
  and g8580 (n5341, n_2394, n_3515);
  and g8581 (n5342, n_3516, n5341);
  not g8582 (n_3521, n5340);
  not g8583 (n_3522, n5342);
  and g8584 (n5343, n_3521, n_3522);
  not g8585 (n_3523, n5333);
  not g8586 (n_3524, n5343);
  and g8587 (n5344, n_3523, n_3524);
  not g8588 (n_3525, n5344);
  and g8589 (n5345, \asqrt[43] , n_3525);
  and g8593 (n5349, n_3283, n_3282);
  and g8594 (n5350, \asqrt[35] , n5349);
  not g8595 (n_3526, n5350);
  and g8596 (n5351, n_3281, n_3526);
  not g8597 (n_3527, n5348);
  not g8598 (n_3528, n5351);
  and g8599 (n5352, n_3527, n_3528);
  and g8600 (n5353, n_2202, n_3523);
  and g8601 (n5354, n_3524, n5353);
  not g8602 (n_3529, n5352);
  not g8603 (n_3530, n5354);
  and g8604 (n5355, n_3529, n_3530);
  not g8605 (n_3531, n5345);
  not g8606 (n_3532, n5355);
  and g8607 (n5356, n_3531, n_3532);
  not g8608 (n_3533, n5356);
  and g8609 (n5357, \asqrt[44] , n_3533);
  and g8613 (n5361, n_3291, n_3290);
  and g8614 (n5362, \asqrt[35] , n5361);
  not g8615 (n_3534, n5362);
  and g8616 (n5363, n_3289, n_3534);
  not g8617 (n_3535, n5360);
  not g8618 (n_3536, n5363);
  and g8619 (n5364, n_3535, n_3536);
  and g8620 (n5365, n_2018, n_3531);
  and g8621 (n5366, n_3532, n5365);
  not g8622 (n_3537, n5364);
  not g8623 (n_3538, n5366);
  and g8624 (n5367, n_3537, n_3538);
  not g8625 (n_3539, n5357);
  not g8626 (n_3540, n5367);
  and g8627 (n5368, n_3539, n_3540);
  not g8628 (n_3541, n5368);
  and g8629 (n5369, \asqrt[45] , n_3541);
  and g8633 (n5373, n_3299, n_3298);
  and g8634 (n5374, \asqrt[35] , n5373);
  not g8635 (n_3542, n5374);
  and g8636 (n5375, n_3297, n_3542);
  not g8637 (n_3543, n5372);
  not g8638 (n_3544, n5375);
  and g8639 (n5376, n_3543, n_3544);
  and g8640 (n5377, n_1842, n_3539);
  and g8641 (n5378, n_3540, n5377);
  not g8642 (n_3545, n5376);
  not g8643 (n_3546, n5378);
  and g8644 (n5379, n_3545, n_3546);
  not g8645 (n_3547, n5369);
  not g8646 (n_3548, n5379);
  and g8647 (n5380, n_3547, n_3548);
  not g8648 (n_3549, n5380);
  and g8649 (n5381, \asqrt[46] , n_3549);
  and g8653 (n5385, n_3307, n_3306);
  and g8654 (n5386, \asqrt[35] , n5385);
  not g8655 (n_3550, n5386);
  and g8656 (n5387, n_3305, n_3550);
  not g8657 (n_3551, n5384);
  not g8658 (n_3552, n5387);
  and g8659 (n5388, n_3551, n_3552);
  and g8660 (n5389, n_1674, n_3547);
  and g8661 (n5390, n_3548, n5389);
  not g8662 (n_3553, n5388);
  not g8663 (n_3554, n5390);
  and g8664 (n5391, n_3553, n_3554);
  not g8665 (n_3555, n5381);
  not g8666 (n_3556, n5391);
  and g8667 (n5392, n_3555, n_3556);
  not g8668 (n_3557, n5392);
  and g8669 (n5393, \asqrt[47] , n_3557);
  and g8673 (n5397, n_3315, n_3314);
  and g8674 (n5398, \asqrt[35] , n5397);
  not g8675 (n_3558, n5398);
  and g8676 (n5399, n_3313, n_3558);
  not g8677 (n_3559, n5396);
  not g8678 (n_3560, n5399);
  and g8679 (n5400, n_3559, n_3560);
  and g8680 (n5401, n_1514, n_3555);
  and g8681 (n5402, n_3556, n5401);
  not g8682 (n_3561, n5400);
  not g8683 (n_3562, n5402);
  and g8684 (n5403, n_3561, n_3562);
  not g8685 (n_3563, n5393);
  not g8686 (n_3564, n5403);
  and g8687 (n5404, n_3563, n_3564);
  not g8688 (n_3565, n5404);
  and g8689 (n5405, \asqrt[48] , n_3565);
  and g8693 (n5409, n_3323, n_3322);
  and g8694 (n5410, \asqrt[35] , n5409);
  not g8695 (n_3566, n5410);
  and g8696 (n5411, n_3321, n_3566);
  not g8697 (n_3567, n5408);
  not g8698 (n_3568, n5411);
  and g8699 (n5412, n_3567, n_3568);
  and g8700 (n5413, n_1362, n_3563);
  and g8701 (n5414, n_3564, n5413);
  not g8702 (n_3569, n5412);
  not g8703 (n_3570, n5414);
  and g8704 (n5415, n_3569, n_3570);
  not g8705 (n_3571, n5405);
  not g8706 (n_3572, n5415);
  and g8707 (n5416, n_3571, n_3572);
  not g8708 (n_3573, n5416);
  and g8709 (n5417, \asqrt[49] , n_3573);
  and g8713 (n5421, n_3331, n_3330);
  and g8714 (n5422, \asqrt[35] , n5421);
  not g8715 (n_3574, n5422);
  and g8716 (n5423, n_3329, n_3574);
  not g8717 (n_3575, n5420);
  not g8718 (n_3576, n5423);
  and g8719 (n5424, n_3575, n_3576);
  and g8720 (n5425, n_1218, n_3571);
  and g8721 (n5426, n_3572, n5425);
  not g8722 (n_3577, n5424);
  not g8723 (n_3578, n5426);
  and g8724 (n5427, n_3577, n_3578);
  not g8725 (n_3579, n5417);
  not g8726 (n_3580, n5427);
  and g8727 (n5428, n_3579, n_3580);
  not g8728 (n_3581, n5428);
  and g8729 (n5429, \asqrt[50] , n_3581);
  and g8733 (n5433, n_3339, n_3338);
  and g8734 (n5434, \asqrt[35] , n5433);
  not g8735 (n_3582, n5434);
  and g8736 (n5435, n_3337, n_3582);
  not g8737 (n_3583, n5432);
  not g8738 (n_3584, n5435);
  and g8739 (n5436, n_3583, n_3584);
  and g8740 (n5437, n_1082, n_3579);
  and g8741 (n5438, n_3580, n5437);
  not g8742 (n_3585, n5436);
  not g8743 (n_3586, n5438);
  and g8744 (n5439, n_3585, n_3586);
  not g8745 (n_3587, n5429);
  not g8746 (n_3588, n5439);
  and g8747 (n5440, n_3587, n_3588);
  not g8748 (n_3589, n5440);
  and g8749 (n5441, \asqrt[51] , n_3589);
  and g8753 (n5445, n_3347, n_3346);
  and g8754 (n5446, \asqrt[35] , n5445);
  not g8755 (n_3590, n5446);
  and g8756 (n5447, n_3345, n_3590);
  not g8757 (n_3591, n5444);
  not g8758 (n_3592, n5447);
  and g8759 (n5448, n_3591, n_3592);
  and g8760 (n5449, n_954, n_3587);
  and g8761 (n5450, n_3588, n5449);
  not g8762 (n_3593, n5448);
  not g8763 (n_3594, n5450);
  and g8764 (n5451, n_3593, n_3594);
  not g8765 (n_3595, n5441);
  not g8766 (n_3596, n5451);
  and g8767 (n5452, n_3595, n_3596);
  not g8768 (n_3597, n5452);
  and g8769 (n5453, \asqrt[52] , n_3597);
  and g8773 (n5457, n_3355, n_3354);
  and g8774 (n5458, \asqrt[35] , n5457);
  not g8775 (n_3598, n5458);
  and g8776 (n5459, n_3353, n_3598);
  not g8777 (n_3599, n5456);
  not g8778 (n_3600, n5459);
  and g8779 (n5460, n_3599, n_3600);
  and g8780 (n5461, n_834, n_3595);
  and g8781 (n5462, n_3596, n5461);
  not g8782 (n_3601, n5460);
  not g8783 (n_3602, n5462);
  and g8784 (n5463, n_3601, n_3602);
  not g8785 (n_3603, n5453);
  not g8786 (n_3604, n5463);
  and g8787 (n5464, n_3603, n_3604);
  not g8788 (n_3605, n5464);
  and g8789 (n5465, \asqrt[53] , n_3605);
  and g8793 (n5469, n_3363, n_3362);
  and g8794 (n5470, \asqrt[35] , n5469);
  not g8795 (n_3606, n5470);
  and g8796 (n5471, n_3361, n_3606);
  not g8797 (n_3607, n5468);
  not g8798 (n_3608, n5471);
  and g8799 (n5472, n_3607, n_3608);
  and g8800 (n5473, n_722, n_3603);
  and g8801 (n5474, n_3604, n5473);
  not g8802 (n_3609, n5472);
  not g8803 (n_3610, n5474);
  and g8804 (n5475, n_3609, n_3610);
  not g8805 (n_3611, n5465);
  not g8806 (n_3612, n5475);
  and g8807 (n5476, n_3611, n_3612);
  not g8808 (n_3613, n5476);
  and g8809 (n5477, \asqrt[54] , n_3613);
  and g8813 (n5481, n_3371, n_3370);
  and g8814 (n5482, \asqrt[35] , n5481);
  not g8815 (n_3614, n5482);
  and g8816 (n5483, n_3369, n_3614);
  not g8817 (n_3615, n5480);
  not g8818 (n_3616, n5483);
  and g8819 (n5484, n_3615, n_3616);
  and g8820 (n5485, n_618, n_3611);
  and g8821 (n5486, n_3612, n5485);
  not g8822 (n_3617, n5484);
  not g8823 (n_3618, n5486);
  and g8824 (n5487, n_3617, n_3618);
  not g8825 (n_3619, n5477);
  not g8826 (n_3620, n5487);
  and g8827 (n5488, n_3619, n_3620);
  not g8828 (n_3621, n5488);
  and g8829 (n5489, \asqrt[55] , n_3621);
  and g8833 (n5493, n_3379, n_3378);
  and g8834 (n5494, \asqrt[35] , n5493);
  not g8835 (n_3622, n5494);
  and g8836 (n5495, n_3377, n_3622);
  not g8837 (n_3623, n5492);
  not g8838 (n_3624, n5495);
  and g8839 (n5496, n_3623, n_3624);
  and g8840 (n5497, n_522, n_3619);
  and g8841 (n5498, n_3620, n5497);
  not g8842 (n_3625, n5496);
  not g8843 (n_3626, n5498);
  and g8844 (n5499, n_3625, n_3626);
  not g8845 (n_3627, n5489);
  not g8846 (n_3628, n5499);
  and g8847 (n5500, n_3627, n_3628);
  not g8848 (n_3629, n5500);
  and g8849 (n5501, \asqrt[56] , n_3629);
  and g8853 (n5505, n_3387, n_3386);
  and g8854 (n5506, \asqrt[35] , n5505);
  not g8855 (n_3630, n5506);
  and g8856 (n5507, n_3385, n_3630);
  not g8857 (n_3631, n5504);
  not g8858 (n_3632, n5507);
  and g8859 (n5508, n_3631, n_3632);
  and g8860 (n5509, n_434, n_3627);
  and g8861 (n5510, n_3628, n5509);
  not g8862 (n_3633, n5508);
  not g8863 (n_3634, n5510);
  and g8864 (n5511, n_3633, n_3634);
  not g8865 (n_3635, n5501);
  not g8866 (n_3636, n5511);
  and g8867 (n5512, n_3635, n_3636);
  not g8868 (n_3637, n5512);
  and g8869 (n5513, \asqrt[57] , n_3637);
  and g8873 (n5517, n_3395, n_3394);
  and g8874 (n5518, \asqrt[35] , n5517);
  not g8875 (n_3638, n5518);
  and g8876 (n5519, n_3393, n_3638);
  not g8877 (n_3639, n5516);
  not g8878 (n_3640, n5519);
  and g8879 (n5520, n_3639, n_3640);
  and g8880 (n5521, n_354, n_3635);
  and g8881 (n5522, n_3636, n5521);
  not g8882 (n_3641, n5520);
  not g8883 (n_3642, n5522);
  and g8884 (n5523, n_3641, n_3642);
  not g8885 (n_3643, n5513);
  not g8886 (n_3644, n5523);
  and g8887 (n5524, n_3643, n_3644);
  not g8888 (n_3645, n5524);
  and g8889 (n5525, \asqrt[58] , n_3645);
  and g8893 (n5529, n_3403, n_3402);
  and g8894 (n5530, \asqrt[35] , n5529);
  not g8895 (n_3646, n5530);
  and g8896 (n5531, n_3401, n_3646);
  not g8897 (n_3647, n5528);
  not g8898 (n_3648, n5531);
  and g8899 (n5532, n_3647, n_3648);
  and g8900 (n5533, n_282, n_3643);
  and g8901 (n5534, n_3644, n5533);
  not g8902 (n_3649, n5532);
  not g8903 (n_3650, n5534);
  and g8904 (n5535, n_3649, n_3650);
  not g8905 (n_3651, n5525);
  not g8906 (n_3652, n5535);
  and g8907 (n5536, n_3651, n_3652);
  not g8908 (n_3653, n5536);
  and g8909 (n5537, \asqrt[59] , n_3653);
  and g8913 (n5541, n_3411, n_3410);
  and g8914 (n5542, \asqrt[35] , n5541);
  not g8915 (n_3654, n5542);
  and g8916 (n5543, n_3409, n_3654);
  not g8917 (n_3655, n5540);
  not g8918 (n_3656, n5543);
  and g8919 (n5544, n_3655, n_3656);
  and g8920 (n5545, n_218, n_3651);
  and g8921 (n5546, n_3652, n5545);
  not g8922 (n_3657, n5544);
  not g8923 (n_3658, n5546);
  and g8924 (n5547, n_3657, n_3658);
  not g8925 (n_3659, n5537);
  not g8926 (n_3660, n5547);
  and g8927 (n5548, n_3659, n_3660);
  not g8928 (n_3661, n5548);
  and g8929 (n5549, \asqrt[60] , n_3661);
  and g8933 (n5553, n_3419, n_3418);
  and g8934 (n5554, \asqrt[35] , n5553);
  not g8935 (n_3662, n5554);
  and g8936 (n5555, n_3417, n_3662);
  not g8937 (n_3663, n5552);
  not g8938 (n_3664, n5555);
  and g8939 (n5556, n_3663, n_3664);
  and g8940 (n5557, n_162, n_3659);
  and g8941 (n5558, n_3660, n5557);
  not g8942 (n_3665, n5556);
  not g8943 (n_3666, n5558);
  and g8944 (n5559, n_3665, n_3666);
  not g8945 (n_3667, n5549);
  not g8946 (n_3668, n5559);
  and g8947 (n5560, n_3667, n_3668);
  not g8948 (n_3669, n5560);
  and g8949 (n5561, \asqrt[61] , n_3669);
  and g8953 (n5565, n_3427, n_3426);
  and g8954 (n5566, \asqrt[35] , n5565);
  not g8955 (n_3670, n5566);
  and g8956 (n5567, n_3425, n_3670);
  not g8957 (n_3671, n5564);
  not g8958 (n_3672, n5567);
  and g8959 (n5568, n_3671, n_3672);
  and g8960 (n5569, n_115, n_3667);
  and g8961 (n5570, n_3668, n5569);
  not g8962 (n_3673, n5568);
  not g8963 (n_3674, n5570);
  and g8964 (n5571, n_3673, n_3674);
  not g8965 (n_3675, n5561);
  not g8966 (n_3676, n5571);
  and g8967 (n5572, n_3675, n_3676);
  not g8968 (n_3677, n5572);
  and g8969 (n5573, \asqrt[62] , n_3677);
  and g8970 (n5574, n_76, n_3675);
  and g8971 (n5575, n_3676, n5574);
  and g8975 (n5579, n_3435, n_3433);
  and g8976 (n5580, \asqrt[35] , n5579);
  not g8977 (n_3678, n5580);
  and g8978 (n5581, n_3434, n_3678);
  not g8979 (n_3679, n5578);
  not g8980 (n_3680, n5581);
  and g8981 (n5582, n_3679, n_3680);
  not g8982 (n_3681, n5575);
  not g8983 (n_3682, n5582);
  and g8984 (n5583, n_3681, n_3682);
  not g8985 (n_3683, n5573);
  not g8986 (n_3684, n5583);
  and g8987 (n5584, n_3683, n_3684);
  and g8991 (n5588, n_3443, n_3442);
  and g8992 (n5589, \asqrt[35] , n5588);
  not g8993 (n_3685, n5589);
  and g8994 (n5590, n_3441, n_3685);
  not g8995 (n_3686, n5587);
  not g8996 (n_3687, n5590);
  and g8997 (n5591, n_3686, n_3687);
  and g8998 (n5592, n_3450, n_3449);
  and g8999 (n5593, \asqrt[35] , n5592);
  not g9002 (n_3689, n5591);
  not g9004 (n_3690, n5584);
  not g9006 (n_3691, n5596);
  and g9007 (n5597, n_21, n_3691);
  and g9008 (n5598, n_3683, n5591);
  and g9009 (n5599, n_3684, n5598);
  and g9010 (n5600, n_3449, \asqrt[35] );
  not g9011 (n_3692, n5600);
  and g9012 (n5601, n5228, n_3692);
  not g9013 (n_3693, n5592);
  and g9014 (n5602, \asqrt[63] , n_3693);
  not g9015 (n_3694, n5601);
  and g9016 (n5603, n_3694, n5602);
  not g9022 (n_3695, n5603);
  not g9023 (n_3696, n5608);
  not g9025 (n_3697, n5599);
  and g9029 (n5612, \a[68] , \asqrt[34] );
  not g9030 (n_3702, \a[66] );
  not g9031 (n_3703, \a[67] );
  and g9032 (n5613, n_3702, n_3703);
  and g9033 (n5614, n_3462, n5613);
  not g9034 (n_3704, n5612);
  not g9035 (n_3705, n5614);
  and g9036 (n5615, n_3704, n_3705);
  not g9037 (n_3706, n5615);
  and g9038 (n5616, \asqrt[35] , n_3706);
  and g9044 (n5622, n_3462, \asqrt[34] );
  not g9045 (n_3707, n5622);
  and g9046 (n5623, \a[69] , n_3707);
  and g9047 (n5624, n5257, \asqrt[34] );
  not g9048 (n_3708, n5623);
  not g9049 (n_3709, n5624);
  and g9050 (n5625, n_3708, n_3709);
  not g9051 (n_3710, n5621);
  and g9052 (n5626, n_3710, n5625);
  not g9053 (n_3711, n5616);
  not g9054 (n_3712, n5626);
  and g9055 (n5627, n_3711, n_3712);
  not g9056 (n_3713, n5627);
  and g9057 (n5628, \asqrt[36] , n_3713);
  not g9058 (n_3714, \asqrt[36] );
  and g9059 (n5629, n_3714, n_3711);
  and g9060 (n5630, n_3712, n5629);
  not g9064 (n_3715, n5597);
  not g9066 (n_3716, n5634);
  and g9067 (n5635, n_3709, n_3716);
  not g9068 (n_3717, n5635);
  and g9069 (n5636, \a[70] , n_3717);
  and g9070 (n5637, n_3230, n_3716);
  and g9071 (n5638, n_3709, n5637);
  not g9072 (n_3718, n5636);
  not g9073 (n_3719, n5638);
  and g9074 (n5639, n_3718, n_3719);
  not g9075 (n_3720, n5630);
  not g9076 (n_3721, n5639);
  and g9077 (n5640, n_3720, n_3721);
  not g9078 (n_3722, n5628);
  not g9079 (n_3723, n5640);
  and g9080 (n5641, n_3722, n_3723);
  not g9081 (n_3724, n5641);
  and g9082 (n5642, \asqrt[37] , n_3724);
  and g9083 (n5643, n_3471, n_3470);
  not g9084 (n_3725, n5269);
  and g9085 (n5644, n_3725, n5643);
  and g9086 (n5645, \asqrt[34] , n5644);
  and g9087 (n5646, \asqrt[34] , n5643);
  not g9088 (n_3726, n5646);
  and g9089 (n5647, n5269, n_3726);
  not g9090 (n_3727, n5645);
  not g9091 (n_3728, n5647);
  and g9092 (n5648, n_3727, n_3728);
  and g9093 (n5649, n_3474, n_3722);
  and g9094 (n5650, n_3723, n5649);
  not g9095 (n_3729, n5648);
  not g9096 (n_3730, n5650);
  and g9097 (n5651, n_3729, n_3730);
  not g9098 (n_3731, n5642);
  not g9099 (n_3732, n5651);
  and g9100 (n5652, n_3731, n_3732);
  not g9101 (n_3733, n5652);
  and g9102 (n5653, \asqrt[38] , n_3733);
  and g9106 (n5657, n_3482, n_3480);
  and g9107 (n5658, \asqrt[34] , n5657);
  not g9108 (n_3734, n5658);
  and g9109 (n5659, n_3481, n_3734);
  not g9110 (n_3735, n5656);
  not g9111 (n_3736, n5659);
  and g9112 (n5660, n_3735, n_3736);
  and g9113 (n5661, n_3242, n_3731);
  and g9114 (n5662, n_3732, n5661);
  not g9115 (n_3737, n5660);
  not g9116 (n_3738, n5662);
  and g9117 (n5663, n_3737, n_3738);
  not g9118 (n_3739, n5653);
  not g9119 (n_3740, n5663);
  and g9120 (n5664, n_3739, n_3740);
  not g9121 (n_3741, n5664);
  and g9122 (n5665, \asqrt[39] , n_3741);
  and g9126 (n5669, n_3491, n_3490);
  and g9127 (n5670, \asqrt[34] , n5669);
  not g9128 (n_3742, n5670);
  and g9129 (n5671, n_3489, n_3742);
  not g9130 (n_3743, n5668);
  not g9131 (n_3744, n5671);
  and g9132 (n5672, n_3743, n_3744);
  and g9133 (n5673, n_3018, n_3739);
  and g9134 (n5674, n_3740, n5673);
  not g9135 (n_3745, n5672);
  not g9136 (n_3746, n5674);
  and g9137 (n5675, n_3745, n_3746);
  not g9138 (n_3747, n5665);
  not g9139 (n_3748, n5675);
  and g9140 (n5676, n_3747, n_3748);
  not g9141 (n_3749, n5676);
  and g9142 (n5677, \asqrt[40] , n_3749);
  and g9146 (n5681, n_3499, n_3498);
  and g9147 (n5682, \asqrt[34] , n5681);
  not g9148 (n_3750, n5682);
  and g9149 (n5683, n_3497, n_3750);
  not g9150 (n_3751, n5680);
  not g9151 (n_3752, n5683);
  and g9152 (n5684, n_3751, n_3752);
  and g9153 (n5685, n_2802, n_3747);
  and g9154 (n5686, n_3748, n5685);
  not g9155 (n_3753, n5684);
  not g9156 (n_3754, n5686);
  and g9157 (n5687, n_3753, n_3754);
  not g9158 (n_3755, n5677);
  not g9159 (n_3756, n5687);
  and g9160 (n5688, n_3755, n_3756);
  not g9161 (n_3757, n5688);
  and g9162 (n5689, \asqrt[41] , n_3757);
  and g9166 (n5693, n_3507, n_3506);
  and g9167 (n5694, \asqrt[34] , n5693);
  not g9168 (n_3758, n5694);
  and g9169 (n5695, n_3505, n_3758);
  not g9170 (n_3759, n5692);
  not g9171 (n_3760, n5695);
  and g9172 (n5696, n_3759, n_3760);
  and g9173 (n5697, n_2594, n_3755);
  and g9174 (n5698, n_3756, n5697);
  not g9175 (n_3761, n5696);
  not g9176 (n_3762, n5698);
  and g9177 (n5699, n_3761, n_3762);
  not g9178 (n_3763, n5689);
  not g9179 (n_3764, n5699);
  and g9180 (n5700, n_3763, n_3764);
  not g9181 (n_3765, n5700);
  and g9182 (n5701, \asqrt[42] , n_3765);
  and g9186 (n5705, n_3515, n_3514);
  and g9187 (n5706, \asqrt[34] , n5705);
  not g9188 (n_3766, n5706);
  and g9189 (n5707, n_3513, n_3766);
  not g9190 (n_3767, n5704);
  not g9191 (n_3768, n5707);
  and g9192 (n5708, n_3767, n_3768);
  and g9193 (n5709, n_2394, n_3763);
  and g9194 (n5710, n_3764, n5709);
  not g9195 (n_3769, n5708);
  not g9196 (n_3770, n5710);
  and g9197 (n5711, n_3769, n_3770);
  not g9198 (n_3771, n5701);
  not g9199 (n_3772, n5711);
  and g9200 (n5712, n_3771, n_3772);
  not g9201 (n_3773, n5712);
  and g9202 (n5713, \asqrt[43] , n_3773);
  and g9206 (n5717, n_3523, n_3522);
  and g9207 (n5718, \asqrt[34] , n5717);
  not g9208 (n_3774, n5718);
  and g9209 (n5719, n_3521, n_3774);
  not g9210 (n_3775, n5716);
  not g9211 (n_3776, n5719);
  and g9212 (n5720, n_3775, n_3776);
  and g9213 (n5721, n_2202, n_3771);
  and g9214 (n5722, n_3772, n5721);
  not g9215 (n_3777, n5720);
  not g9216 (n_3778, n5722);
  and g9217 (n5723, n_3777, n_3778);
  not g9218 (n_3779, n5713);
  not g9219 (n_3780, n5723);
  and g9220 (n5724, n_3779, n_3780);
  not g9221 (n_3781, n5724);
  and g9222 (n5725, \asqrt[44] , n_3781);
  and g9226 (n5729, n_3531, n_3530);
  and g9227 (n5730, \asqrt[34] , n5729);
  not g9228 (n_3782, n5730);
  and g9229 (n5731, n_3529, n_3782);
  not g9230 (n_3783, n5728);
  not g9231 (n_3784, n5731);
  and g9232 (n5732, n_3783, n_3784);
  and g9233 (n5733, n_2018, n_3779);
  and g9234 (n5734, n_3780, n5733);
  not g9235 (n_3785, n5732);
  not g9236 (n_3786, n5734);
  and g9237 (n5735, n_3785, n_3786);
  not g9238 (n_3787, n5725);
  not g9239 (n_3788, n5735);
  and g9240 (n5736, n_3787, n_3788);
  not g9241 (n_3789, n5736);
  and g9242 (n5737, \asqrt[45] , n_3789);
  and g9246 (n5741, n_3539, n_3538);
  and g9247 (n5742, \asqrt[34] , n5741);
  not g9248 (n_3790, n5742);
  and g9249 (n5743, n_3537, n_3790);
  not g9250 (n_3791, n5740);
  not g9251 (n_3792, n5743);
  and g9252 (n5744, n_3791, n_3792);
  and g9253 (n5745, n_1842, n_3787);
  and g9254 (n5746, n_3788, n5745);
  not g9255 (n_3793, n5744);
  not g9256 (n_3794, n5746);
  and g9257 (n5747, n_3793, n_3794);
  not g9258 (n_3795, n5737);
  not g9259 (n_3796, n5747);
  and g9260 (n5748, n_3795, n_3796);
  not g9261 (n_3797, n5748);
  and g9262 (n5749, \asqrt[46] , n_3797);
  and g9266 (n5753, n_3547, n_3546);
  and g9267 (n5754, \asqrt[34] , n5753);
  not g9268 (n_3798, n5754);
  and g9269 (n5755, n_3545, n_3798);
  not g9270 (n_3799, n5752);
  not g9271 (n_3800, n5755);
  and g9272 (n5756, n_3799, n_3800);
  and g9273 (n5757, n_1674, n_3795);
  and g9274 (n5758, n_3796, n5757);
  not g9275 (n_3801, n5756);
  not g9276 (n_3802, n5758);
  and g9277 (n5759, n_3801, n_3802);
  not g9278 (n_3803, n5749);
  not g9279 (n_3804, n5759);
  and g9280 (n5760, n_3803, n_3804);
  not g9281 (n_3805, n5760);
  and g9282 (n5761, \asqrt[47] , n_3805);
  and g9286 (n5765, n_3555, n_3554);
  and g9287 (n5766, \asqrt[34] , n5765);
  not g9288 (n_3806, n5766);
  and g9289 (n5767, n_3553, n_3806);
  not g9290 (n_3807, n5764);
  not g9291 (n_3808, n5767);
  and g9292 (n5768, n_3807, n_3808);
  and g9293 (n5769, n_1514, n_3803);
  and g9294 (n5770, n_3804, n5769);
  not g9295 (n_3809, n5768);
  not g9296 (n_3810, n5770);
  and g9297 (n5771, n_3809, n_3810);
  not g9298 (n_3811, n5761);
  not g9299 (n_3812, n5771);
  and g9300 (n5772, n_3811, n_3812);
  not g9301 (n_3813, n5772);
  and g9302 (n5773, \asqrt[48] , n_3813);
  and g9306 (n5777, n_3563, n_3562);
  and g9307 (n5778, \asqrt[34] , n5777);
  not g9308 (n_3814, n5778);
  and g9309 (n5779, n_3561, n_3814);
  not g9310 (n_3815, n5776);
  not g9311 (n_3816, n5779);
  and g9312 (n5780, n_3815, n_3816);
  and g9313 (n5781, n_1362, n_3811);
  and g9314 (n5782, n_3812, n5781);
  not g9315 (n_3817, n5780);
  not g9316 (n_3818, n5782);
  and g9317 (n5783, n_3817, n_3818);
  not g9318 (n_3819, n5773);
  not g9319 (n_3820, n5783);
  and g9320 (n5784, n_3819, n_3820);
  not g9321 (n_3821, n5784);
  and g9322 (n5785, \asqrt[49] , n_3821);
  and g9326 (n5789, n_3571, n_3570);
  and g9327 (n5790, \asqrt[34] , n5789);
  not g9328 (n_3822, n5790);
  and g9329 (n5791, n_3569, n_3822);
  not g9330 (n_3823, n5788);
  not g9331 (n_3824, n5791);
  and g9332 (n5792, n_3823, n_3824);
  and g9333 (n5793, n_1218, n_3819);
  and g9334 (n5794, n_3820, n5793);
  not g9335 (n_3825, n5792);
  not g9336 (n_3826, n5794);
  and g9337 (n5795, n_3825, n_3826);
  not g9338 (n_3827, n5785);
  not g9339 (n_3828, n5795);
  and g9340 (n5796, n_3827, n_3828);
  not g9341 (n_3829, n5796);
  and g9342 (n5797, \asqrt[50] , n_3829);
  and g9346 (n5801, n_3579, n_3578);
  and g9347 (n5802, \asqrt[34] , n5801);
  not g9348 (n_3830, n5802);
  and g9349 (n5803, n_3577, n_3830);
  not g9350 (n_3831, n5800);
  not g9351 (n_3832, n5803);
  and g9352 (n5804, n_3831, n_3832);
  and g9353 (n5805, n_1082, n_3827);
  and g9354 (n5806, n_3828, n5805);
  not g9355 (n_3833, n5804);
  not g9356 (n_3834, n5806);
  and g9357 (n5807, n_3833, n_3834);
  not g9358 (n_3835, n5797);
  not g9359 (n_3836, n5807);
  and g9360 (n5808, n_3835, n_3836);
  not g9361 (n_3837, n5808);
  and g9362 (n5809, \asqrt[51] , n_3837);
  and g9366 (n5813, n_3587, n_3586);
  and g9367 (n5814, \asqrt[34] , n5813);
  not g9368 (n_3838, n5814);
  and g9369 (n5815, n_3585, n_3838);
  not g9370 (n_3839, n5812);
  not g9371 (n_3840, n5815);
  and g9372 (n5816, n_3839, n_3840);
  and g9373 (n5817, n_954, n_3835);
  and g9374 (n5818, n_3836, n5817);
  not g9375 (n_3841, n5816);
  not g9376 (n_3842, n5818);
  and g9377 (n5819, n_3841, n_3842);
  not g9378 (n_3843, n5809);
  not g9379 (n_3844, n5819);
  and g9380 (n5820, n_3843, n_3844);
  not g9381 (n_3845, n5820);
  and g9382 (n5821, \asqrt[52] , n_3845);
  and g9386 (n5825, n_3595, n_3594);
  and g9387 (n5826, \asqrt[34] , n5825);
  not g9388 (n_3846, n5826);
  and g9389 (n5827, n_3593, n_3846);
  not g9390 (n_3847, n5824);
  not g9391 (n_3848, n5827);
  and g9392 (n5828, n_3847, n_3848);
  and g9393 (n5829, n_834, n_3843);
  and g9394 (n5830, n_3844, n5829);
  not g9395 (n_3849, n5828);
  not g9396 (n_3850, n5830);
  and g9397 (n5831, n_3849, n_3850);
  not g9398 (n_3851, n5821);
  not g9399 (n_3852, n5831);
  and g9400 (n5832, n_3851, n_3852);
  not g9401 (n_3853, n5832);
  and g9402 (n5833, \asqrt[53] , n_3853);
  and g9406 (n5837, n_3603, n_3602);
  and g9407 (n5838, \asqrt[34] , n5837);
  not g9408 (n_3854, n5838);
  and g9409 (n5839, n_3601, n_3854);
  not g9410 (n_3855, n5836);
  not g9411 (n_3856, n5839);
  and g9412 (n5840, n_3855, n_3856);
  and g9413 (n5841, n_722, n_3851);
  and g9414 (n5842, n_3852, n5841);
  not g9415 (n_3857, n5840);
  not g9416 (n_3858, n5842);
  and g9417 (n5843, n_3857, n_3858);
  not g9418 (n_3859, n5833);
  not g9419 (n_3860, n5843);
  and g9420 (n5844, n_3859, n_3860);
  not g9421 (n_3861, n5844);
  and g9422 (n5845, \asqrt[54] , n_3861);
  and g9426 (n5849, n_3611, n_3610);
  and g9427 (n5850, \asqrt[34] , n5849);
  not g9428 (n_3862, n5850);
  and g9429 (n5851, n_3609, n_3862);
  not g9430 (n_3863, n5848);
  not g9431 (n_3864, n5851);
  and g9432 (n5852, n_3863, n_3864);
  and g9433 (n5853, n_618, n_3859);
  and g9434 (n5854, n_3860, n5853);
  not g9435 (n_3865, n5852);
  not g9436 (n_3866, n5854);
  and g9437 (n5855, n_3865, n_3866);
  not g9438 (n_3867, n5845);
  not g9439 (n_3868, n5855);
  and g9440 (n5856, n_3867, n_3868);
  not g9441 (n_3869, n5856);
  and g9442 (n5857, \asqrt[55] , n_3869);
  and g9446 (n5861, n_3619, n_3618);
  and g9447 (n5862, \asqrt[34] , n5861);
  not g9448 (n_3870, n5862);
  and g9449 (n5863, n_3617, n_3870);
  not g9450 (n_3871, n5860);
  not g9451 (n_3872, n5863);
  and g9452 (n5864, n_3871, n_3872);
  and g9453 (n5865, n_522, n_3867);
  and g9454 (n5866, n_3868, n5865);
  not g9455 (n_3873, n5864);
  not g9456 (n_3874, n5866);
  and g9457 (n5867, n_3873, n_3874);
  not g9458 (n_3875, n5857);
  not g9459 (n_3876, n5867);
  and g9460 (n5868, n_3875, n_3876);
  not g9461 (n_3877, n5868);
  and g9462 (n5869, \asqrt[56] , n_3877);
  and g9466 (n5873, n_3627, n_3626);
  and g9467 (n5874, \asqrt[34] , n5873);
  not g9468 (n_3878, n5874);
  and g9469 (n5875, n_3625, n_3878);
  not g9470 (n_3879, n5872);
  not g9471 (n_3880, n5875);
  and g9472 (n5876, n_3879, n_3880);
  and g9473 (n5877, n_434, n_3875);
  and g9474 (n5878, n_3876, n5877);
  not g9475 (n_3881, n5876);
  not g9476 (n_3882, n5878);
  and g9477 (n5879, n_3881, n_3882);
  not g9478 (n_3883, n5869);
  not g9479 (n_3884, n5879);
  and g9480 (n5880, n_3883, n_3884);
  not g9481 (n_3885, n5880);
  and g9482 (n5881, \asqrt[57] , n_3885);
  and g9486 (n5885, n_3635, n_3634);
  and g9487 (n5886, \asqrt[34] , n5885);
  not g9488 (n_3886, n5886);
  and g9489 (n5887, n_3633, n_3886);
  not g9490 (n_3887, n5884);
  not g9491 (n_3888, n5887);
  and g9492 (n5888, n_3887, n_3888);
  and g9493 (n5889, n_354, n_3883);
  and g9494 (n5890, n_3884, n5889);
  not g9495 (n_3889, n5888);
  not g9496 (n_3890, n5890);
  and g9497 (n5891, n_3889, n_3890);
  not g9498 (n_3891, n5881);
  not g9499 (n_3892, n5891);
  and g9500 (n5892, n_3891, n_3892);
  not g9501 (n_3893, n5892);
  and g9502 (n5893, \asqrt[58] , n_3893);
  and g9506 (n5897, n_3643, n_3642);
  and g9507 (n5898, \asqrt[34] , n5897);
  not g9508 (n_3894, n5898);
  and g9509 (n5899, n_3641, n_3894);
  not g9510 (n_3895, n5896);
  not g9511 (n_3896, n5899);
  and g9512 (n5900, n_3895, n_3896);
  and g9513 (n5901, n_282, n_3891);
  and g9514 (n5902, n_3892, n5901);
  not g9515 (n_3897, n5900);
  not g9516 (n_3898, n5902);
  and g9517 (n5903, n_3897, n_3898);
  not g9518 (n_3899, n5893);
  not g9519 (n_3900, n5903);
  and g9520 (n5904, n_3899, n_3900);
  not g9521 (n_3901, n5904);
  and g9522 (n5905, \asqrt[59] , n_3901);
  and g9526 (n5909, n_3651, n_3650);
  and g9527 (n5910, \asqrt[34] , n5909);
  not g9528 (n_3902, n5910);
  and g9529 (n5911, n_3649, n_3902);
  not g9530 (n_3903, n5908);
  not g9531 (n_3904, n5911);
  and g9532 (n5912, n_3903, n_3904);
  and g9533 (n5913, n_218, n_3899);
  and g9534 (n5914, n_3900, n5913);
  not g9535 (n_3905, n5912);
  not g9536 (n_3906, n5914);
  and g9537 (n5915, n_3905, n_3906);
  not g9538 (n_3907, n5905);
  not g9539 (n_3908, n5915);
  and g9540 (n5916, n_3907, n_3908);
  not g9541 (n_3909, n5916);
  and g9542 (n5917, \asqrt[60] , n_3909);
  and g9546 (n5921, n_3659, n_3658);
  and g9547 (n5922, \asqrt[34] , n5921);
  not g9548 (n_3910, n5922);
  and g9549 (n5923, n_3657, n_3910);
  not g9550 (n_3911, n5920);
  not g9551 (n_3912, n5923);
  and g9552 (n5924, n_3911, n_3912);
  and g9553 (n5925, n_162, n_3907);
  and g9554 (n5926, n_3908, n5925);
  not g9555 (n_3913, n5924);
  not g9556 (n_3914, n5926);
  and g9557 (n5927, n_3913, n_3914);
  not g9558 (n_3915, n5917);
  not g9559 (n_3916, n5927);
  and g9560 (n5928, n_3915, n_3916);
  not g9561 (n_3917, n5928);
  and g9562 (n5929, \asqrt[61] , n_3917);
  and g9566 (n5933, n_3667, n_3666);
  and g9567 (n5934, \asqrt[34] , n5933);
  not g9568 (n_3918, n5934);
  and g9569 (n5935, n_3665, n_3918);
  not g9570 (n_3919, n5932);
  not g9571 (n_3920, n5935);
  and g9572 (n5936, n_3919, n_3920);
  and g9573 (n5937, n_115, n_3915);
  and g9574 (n5938, n_3916, n5937);
  not g9575 (n_3921, n5936);
  not g9576 (n_3922, n5938);
  and g9577 (n5939, n_3921, n_3922);
  not g9578 (n_3923, n5929);
  not g9579 (n_3924, n5939);
  and g9580 (n5940, n_3923, n_3924);
  not g9581 (n_3925, n5940);
  and g9582 (n5941, \asqrt[62] , n_3925);
  and g9586 (n5945, n_3675, n_3674);
  and g9587 (n5946, \asqrt[34] , n5945);
  not g9588 (n_3926, n5946);
  and g9589 (n5947, n_3673, n_3926);
  not g9590 (n_3927, n5944);
  not g9591 (n_3928, n5947);
  and g9592 (n5948, n_3927, n_3928);
  and g9593 (n5949, n_76, n_3923);
  and g9594 (n5950, n_3924, n5949);
  not g9595 (n_3929, n5948);
  not g9596 (n_3930, n5950);
  and g9597 (n5951, n_3929, n_3930);
  not g9598 (n_3931, n5941);
  not g9599 (n_3932, n5951);
  and g9600 (n5952, n_3931, n_3932);
  and g9604 (n5956, n_3683, n_3681);
  and g9605 (n5957, \asqrt[34] , n5956);
  not g9606 (n_3933, n5957);
  and g9607 (n5958, n_3682, n_3933);
  not g9608 (n_3934, n5955);
  not g9609 (n_3935, n5958);
  and g9610 (n5959, n_3934, n_3935);
  and g9611 (n5960, n_3690, n_3689);
  and g9612 (n5961, \asqrt[34] , n5960);
  not g9615 (n_3937, n5959);
  not g9617 (n_3938, n5952);
  not g9619 (n_3939, n5964);
  and g9620 (n5965, n_21, n_3939);
  and g9621 (n5966, n_3931, n5959);
  and g9622 (n5967, n_3932, n5966);
  and g9623 (n5968, n_3689, \asqrt[34] );
  not g9624 (n_3940, n5968);
  and g9625 (n5969, n5584, n_3940);
  not g9626 (n_3941, n5960);
  and g9627 (n5970, \asqrt[63] , n_3941);
  not g9628 (n_3942, n5969);
  and g9629 (n5971, n_3942, n5970);
  not g9635 (n_3943, n5971);
  not g9636 (n_3944, n5976);
  not g9638 (n_3945, n5967);
  and g9642 (n5980, \a[66] , \asqrt[33] );
  not g9643 (n_3950, \a[64] );
  not g9644 (n_3951, \a[65] );
  and g9645 (n5981, n_3950, n_3951);
  and g9646 (n5982, n_3702, n5981);
  not g9647 (n_3952, n5980);
  not g9648 (n_3953, n5982);
  and g9649 (n5983, n_3952, n_3953);
  not g9650 (n_3954, n5983);
  and g9651 (n5984, \asqrt[34] , n_3954);
  and g9657 (n5990, n_3702, \asqrt[33] );
  not g9658 (n_3955, n5990);
  and g9659 (n5991, \a[67] , n_3955);
  and g9660 (n5992, n5613, \asqrt[33] );
  not g9661 (n_3956, n5991);
  not g9662 (n_3957, n5992);
  and g9663 (n5993, n_3956, n_3957);
  not g9664 (n_3958, n5989);
  and g9665 (n5994, n_3958, n5993);
  not g9666 (n_3959, n5984);
  not g9667 (n_3960, n5994);
  and g9668 (n5995, n_3959, n_3960);
  not g9669 (n_3961, n5995);
  and g9670 (n5996, \asqrt[35] , n_3961);
  not g9671 (n_3962, \asqrt[35] );
  and g9672 (n5997, n_3962, n_3959);
  and g9673 (n5998, n_3960, n5997);
  not g9677 (n_3963, n5965);
  not g9679 (n_3964, n6002);
  and g9680 (n6003, n_3957, n_3964);
  not g9681 (n_3965, n6003);
  and g9682 (n6004, \a[68] , n_3965);
  and g9683 (n6005, n_3462, n_3964);
  and g9684 (n6006, n_3957, n6005);
  not g9685 (n_3966, n6004);
  not g9686 (n_3967, n6006);
  and g9687 (n6007, n_3966, n_3967);
  not g9688 (n_3968, n5998);
  not g9689 (n_3969, n6007);
  and g9690 (n6008, n_3968, n_3969);
  not g9691 (n_3970, n5996);
  not g9692 (n_3971, n6008);
  and g9693 (n6009, n_3970, n_3971);
  not g9694 (n_3972, n6009);
  and g9695 (n6010, \asqrt[36] , n_3972);
  and g9696 (n6011, n_3711, n_3710);
  not g9697 (n_3973, n5625);
  and g9698 (n6012, n_3973, n6011);
  and g9699 (n6013, \asqrt[33] , n6012);
  and g9700 (n6014, \asqrt[33] , n6011);
  not g9701 (n_3974, n6014);
  and g9702 (n6015, n5625, n_3974);
  not g9703 (n_3975, n6013);
  not g9704 (n_3976, n6015);
  and g9705 (n6016, n_3975, n_3976);
  and g9706 (n6017, n_3714, n_3970);
  and g9707 (n6018, n_3971, n6017);
  not g9708 (n_3977, n6016);
  not g9709 (n_3978, n6018);
  and g9710 (n6019, n_3977, n_3978);
  not g9711 (n_3979, n6010);
  not g9712 (n_3980, n6019);
  and g9713 (n6020, n_3979, n_3980);
  not g9714 (n_3981, n6020);
  and g9715 (n6021, \asqrt[37] , n_3981);
  and g9719 (n6025, n_3722, n_3720);
  and g9720 (n6026, \asqrt[33] , n6025);
  not g9721 (n_3982, n6026);
  and g9722 (n6027, n_3721, n_3982);
  not g9723 (n_3983, n6024);
  not g9724 (n_3984, n6027);
  and g9725 (n6028, n_3983, n_3984);
  and g9726 (n6029, n_3474, n_3979);
  and g9727 (n6030, n_3980, n6029);
  not g9728 (n_3985, n6028);
  not g9729 (n_3986, n6030);
  and g9730 (n6031, n_3985, n_3986);
  not g9731 (n_3987, n6021);
  not g9732 (n_3988, n6031);
  and g9733 (n6032, n_3987, n_3988);
  not g9734 (n_3989, n6032);
  and g9735 (n6033, \asqrt[38] , n_3989);
  and g9739 (n6037, n_3731, n_3730);
  and g9740 (n6038, \asqrt[33] , n6037);
  not g9741 (n_3990, n6038);
  and g9742 (n6039, n_3729, n_3990);
  not g9743 (n_3991, n6036);
  not g9744 (n_3992, n6039);
  and g9745 (n6040, n_3991, n_3992);
  and g9746 (n6041, n_3242, n_3987);
  and g9747 (n6042, n_3988, n6041);
  not g9748 (n_3993, n6040);
  not g9749 (n_3994, n6042);
  and g9750 (n6043, n_3993, n_3994);
  not g9751 (n_3995, n6033);
  not g9752 (n_3996, n6043);
  and g9753 (n6044, n_3995, n_3996);
  not g9754 (n_3997, n6044);
  and g9755 (n6045, \asqrt[39] , n_3997);
  and g9759 (n6049, n_3739, n_3738);
  and g9760 (n6050, \asqrt[33] , n6049);
  not g9761 (n_3998, n6050);
  and g9762 (n6051, n_3737, n_3998);
  not g9763 (n_3999, n6048);
  not g9764 (n_4000, n6051);
  and g9765 (n6052, n_3999, n_4000);
  and g9766 (n6053, n_3018, n_3995);
  and g9767 (n6054, n_3996, n6053);
  not g9768 (n_4001, n6052);
  not g9769 (n_4002, n6054);
  and g9770 (n6055, n_4001, n_4002);
  not g9771 (n_4003, n6045);
  not g9772 (n_4004, n6055);
  and g9773 (n6056, n_4003, n_4004);
  not g9774 (n_4005, n6056);
  and g9775 (n6057, \asqrt[40] , n_4005);
  and g9779 (n6061, n_3747, n_3746);
  and g9780 (n6062, \asqrt[33] , n6061);
  not g9781 (n_4006, n6062);
  and g9782 (n6063, n_3745, n_4006);
  not g9783 (n_4007, n6060);
  not g9784 (n_4008, n6063);
  and g9785 (n6064, n_4007, n_4008);
  and g9786 (n6065, n_2802, n_4003);
  and g9787 (n6066, n_4004, n6065);
  not g9788 (n_4009, n6064);
  not g9789 (n_4010, n6066);
  and g9790 (n6067, n_4009, n_4010);
  not g9791 (n_4011, n6057);
  not g9792 (n_4012, n6067);
  and g9793 (n6068, n_4011, n_4012);
  not g9794 (n_4013, n6068);
  and g9795 (n6069, \asqrt[41] , n_4013);
  and g9799 (n6073, n_3755, n_3754);
  and g9800 (n6074, \asqrt[33] , n6073);
  not g9801 (n_4014, n6074);
  and g9802 (n6075, n_3753, n_4014);
  not g9803 (n_4015, n6072);
  not g9804 (n_4016, n6075);
  and g9805 (n6076, n_4015, n_4016);
  and g9806 (n6077, n_2594, n_4011);
  and g9807 (n6078, n_4012, n6077);
  not g9808 (n_4017, n6076);
  not g9809 (n_4018, n6078);
  and g9810 (n6079, n_4017, n_4018);
  not g9811 (n_4019, n6069);
  not g9812 (n_4020, n6079);
  and g9813 (n6080, n_4019, n_4020);
  not g9814 (n_4021, n6080);
  and g9815 (n6081, \asqrt[42] , n_4021);
  and g9819 (n6085, n_3763, n_3762);
  and g9820 (n6086, \asqrt[33] , n6085);
  not g9821 (n_4022, n6086);
  and g9822 (n6087, n_3761, n_4022);
  not g9823 (n_4023, n6084);
  not g9824 (n_4024, n6087);
  and g9825 (n6088, n_4023, n_4024);
  and g9826 (n6089, n_2394, n_4019);
  and g9827 (n6090, n_4020, n6089);
  not g9828 (n_4025, n6088);
  not g9829 (n_4026, n6090);
  and g9830 (n6091, n_4025, n_4026);
  not g9831 (n_4027, n6081);
  not g9832 (n_4028, n6091);
  and g9833 (n6092, n_4027, n_4028);
  not g9834 (n_4029, n6092);
  and g9835 (n6093, \asqrt[43] , n_4029);
  and g9839 (n6097, n_3771, n_3770);
  and g9840 (n6098, \asqrt[33] , n6097);
  not g9841 (n_4030, n6098);
  and g9842 (n6099, n_3769, n_4030);
  not g9843 (n_4031, n6096);
  not g9844 (n_4032, n6099);
  and g9845 (n6100, n_4031, n_4032);
  and g9846 (n6101, n_2202, n_4027);
  and g9847 (n6102, n_4028, n6101);
  not g9848 (n_4033, n6100);
  not g9849 (n_4034, n6102);
  and g9850 (n6103, n_4033, n_4034);
  not g9851 (n_4035, n6093);
  not g9852 (n_4036, n6103);
  and g9853 (n6104, n_4035, n_4036);
  not g9854 (n_4037, n6104);
  and g9855 (n6105, \asqrt[44] , n_4037);
  and g9859 (n6109, n_3779, n_3778);
  and g9860 (n6110, \asqrt[33] , n6109);
  not g9861 (n_4038, n6110);
  and g9862 (n6111, n_3777, n_4038);
  not g9863 (n_4039, n6108);
  not g9864 (n_4040, n6111);
  and g9865 (n6112, n_4039, n_4040);
  and g9866 (n6113, n_2018, n_4035);
  and g9867 (n6114, n_4036, n6113);
  not g9868 (n_4041, n6112);
  not g9869 (n_4042, n6114);
  and g9870 (n6115, n_4041, n_4042);
  not g9871 (n_4043, n6105);
  not g9872 (n_4044, n6115);
  and g9873 (n6116, n_4043, n_4044);
  not g9874 (n_4045, n6116);
  and g9875 (n6117, \asqrt[45] , n_4045);
  and g9879 (n6121, n_3787, n_3786);
  and g9880 (n6122, \asqrt[33] , n6121);
  not g9881 (n_4046, n6122);
  and g9882 (n6123, n_3785, n_4046);
  not g9883 (n_4047, n6120);
  not g9884 (n_4048, n6123);
  and g9885 (n6124, n_4047, n_4048);
  and g9886 (n6125, n_1842, n_4043);
  and g9887 (n6126, n_4044, n6125);
  not g9888 (n_4049, n6124);
  not g9889 (n_4050, n6126);
  and g9890 (n6127, n_4049, n_4050);
  not g9891 (n_4051, n6117);
  not g9892 (n_4052, n6127);
  and g9893 (n6128, n_4051, n_4052);
  not g9894 (n_4053, n6128);
  and g9895 (n6129, \asqrt[46] , n_4053);
  and g9899 (n6133, n_3795, n_3794);
  and g9900 (n6134, \asqrt[33] , n6133);
  not g9901 (n_4054, n6134);
  and g9902 (n6135, n_3793, n_4054);
  not g9903 (n_4055, n6132);
  not g9904 (n_4056, n6135);
  and g9905 (n6136, n_4055, n_4056);
  and g9906 (n6137, n_1674, n_4051);
  and g9907 (n6138, n_4052, n6137);
  not g9908 (n_4057, n6136);
  not g9909 (n_4058, n6138);
  and g9910 (n6139, n_4057, n_4058);
  not g9911 (n_4059, n6129);
  not g9912 (n_4060, n6139);
  and g9913 (n6140, n_4059, n_4060);
  not g9914 (n_4061, n6140);
  and g9915 (n6141, \asqrt[47] , n_4061);
  and g9919 (n6145, n_3803, n_3802);
  and g9920 (n6146, \asqrt[33] , n6145);
  not g9921 (n_4062, n6146);
  and g9922 (n6147, n_3801, n_4062);
  not g9923 (n_4063, n6144);
  not g9924 (n_4064, n6147);
  and g9925 (n6148, n_4063, n_4064);
  and g9926 (n6149, n_1514, n_4059);
  and g9927 (n6150, n_4060, n6149);
  not g9928 (n_4065, n6148);
  not g9929 (n_4066, n6150);
  and g9930 (n6151, n_4065, n_4066);
  not g9931 (n_4067, n6141);
  not g9932 (n_4068, n6151);
  and g9933 (n6152, n_4067, n_4068);
  not g9934 (n_4069, n6152);
  and g9935 (n6153, \asqrt[48] , n_4069);
  and g9939 (n6157, n_3811, n_3810);
  and g9940 (n6158, \asqrt[33] , n6157);
  not g9941 (n_4070, n6158);
  and g9942 (n6159, n_3809, n_4070);
  not g9943 (n_4071, n6156);
  not g9944 (n_4072, n6159);
  and g9945 (n6160, n_4071, n_4072);
  and g9946 (n6161, n_1362, n_4067);
  and g9947 (n6162, n_4068, n6161);
  not g9948 (n_4073, n6160);
  not g9949 (n_4074, n6162);
  and g9950 (n6163, n_4073, n_4074);
  not g9951 (n_4075, n6153);
  not g9952 (n_4076, n6163);
  and g9953 (n6164, n_4075, n_4076);
  not g9954 (n_4077, n6164);
  and g9955 (n6165, \asqrt[49] , n_4077);
  and g9959 (n6169, n_3819, n_3818);
  and g9960 (n6170, \asqrt[33] , n6169);
  not g9961 (n_4078, n6170);
  and g9962 (n6171, n_3817, n_4078);
  not g9963 (n_4079, n6168);
  not g9964 (n_4080, n6171);
  and g9965 (n6172, n_4079, n_4080);
  and g9966 (n6173, n_1218, n_4075);
  and g9967 (n6174, n_4076, n6173);
  not g9968 (n_4081, n6172);
  not g9969 (n_4082, n6174);
  and g9970 (n6175, n_4081, n_4082);
  not g9971 (n_4083, n6165);
  not g9972 (n_4084, n6175);
  and g9973 (n6176, n_4083, n_4084);
  not g9974 (n_4085, n6176);
  and g9975 (n6177, \asqrt[50] , n_4085);
  and g9979 (n6181, n_3827, n_3826);
  and g9980 (n6182, \asqrt[33] , n6181);
  not g9981 (n_4086, n6182);
  and g9982 (n6183, n_3825, n_4086);
  not g9983 (n_4087, n6180);
  not g9984 (n_4088, n6183);
  and g9985 (n6184, n_4087, n_4088);
  and g9986 (n6185, n_1082, n_4083);
  and g9987 (n6186, n_4084, n6185);
  not g9988 (n_4089, n6184);
  not g9989 (n_4090, n6186);
  and g9990 (n6187, n_4089, n_4090);
  not g9991 (n_4091, n6177);
  not g9992 (n_4092, n6187);
  and g9993 (n6188, n_4091, n_4092);
  not g9994 (n_4093, n6188);
  and g9995 (n6189, \asqrt[51] , n_4093);
  and g9999 (n6193, n_3835, n_3834);
  and g10000 (n6194, \asqrt[33] , n6193);
  not g10001 (n_4094, n6194);
  and g10002 (n6195, n_3833, n_4094);
  not g10003 (n_4095, n6192);
  not g10004 (n_4096, n6195);
  and g10005 (n6196, n_4095, n_4096);
  and g10006 (n6197, n_954, n_4091);
  and g10007 (n6198, n_4092, n6197);
  not g10008 (n_4097, n6196);
  not g10009 (n_4098, n6198);
  and g10010 (n6199, n_4097, n_4098);
  not g10011 (n_4099, n6189);
  not g10012 (n_4100, n6199);
  and g10013 (n6200, n_4099, n_4100);
  not g10014 (n_4101, n6200);
  and g10015 (n6201, \asqrt[52] , n_4101);
  and g10019 (n6205, n_3843, n_3842);
  and g10020 (n6206, \asqrt[33] , n6205);
  not g10021 (n_4102, n6206);
  and g10022 (n6207, n_3841, n_4102);
  not g10023 (n_4103, n6204);
  not g10024 (n_4104, n6207);
  and g10025 (n6208, n_4103, n_4104);
  and g10026 (n6209, n_834, n_4099);
  and g10027 (n6210, n_4100, n6209);
  not g10028 (n_4105, n6208);
  not g10029 (n_4106, n6210);
  and g10030 (n6211, n_4105, n_4106);
  not g10031 (n_4107, n6201);
  not g10032 (n_4108, n6211);
  and g10033 (n6212, n_4107, n_4108);
  not g10034 (n_4109, n6212);
  and g10035 (n6213, \asqrt[53] , n_4109);
  and g10039 (n6217, n_3851, n_3850);
  and g10040 (n6218, \asqrt[33] , n6217);
  not g10041 (n_4110, n6218);
  and g10042 (n6219, n_3849, n_4110);
  not g10043 (n_4111, n6216);
  not g10044 (n_4112, n6219);
  and g10045 (n6220, n_4111, n_4112);
  and g10046 (n6221, n_722, n_4107);
  and g10047 (n6222, n_4108, n6221);
  not g10048 (n_4113, n6220);
  not g10049 (n_4114, n6222);
  and g10050 (n6223, n_4113, n_4114);
  not g10051 (n_4115, n6213);
  not g10052 (n_4116, n6223);
  and g10053 (n6224, n_4115, n_4116);
  not g10054 (n_4117, n6224);
  and g10055 (n6225, \asqrt[54] , n_4117);
  and g10059 (n6229, n_3859, n_3858);
  and g10060 (n6230, \asqrt[33] , n6229);
  not g10061 (n_4118, n6230);
  and g10062 (n6231, n_3857, n_4118);
  not g10063 (n_4119, n6228);
  not g10064 (n_4120, n6231);
  and g10065 (n6232, n_4119, n_4120);
  and g10066 (n6233, n_618, n_4115);
  and g10067 (n6234, n_4116, n6233);
  not g10068 (n_4121, n6232);
  not g10069 (n_4122, n6234);
  and g10070 (n6235, n_4121, n_4122);
  not g10071 (n_4123, n6225);
  not g10072 (n_4124, n6235);
  and g10073 (n6236, n_4123, n_4124);
  not g10074 (n_4125, n6236);
  and g10075 (n6237, \asqrt[55] , n_4125);
  and g10079 (n6241, n_3867, n_3866);
  and g10080 (n6242, \asqrt[33] , n6241);
  not g10081 (n_4126, n6242);
  and g10082 (n6243, n_3865, n_4126);
  not g10083 (n_4127, n6240);
  not g10084 (n_4128, n6243);
  and g10085 (n6244, n_4127, n_4128);
  and g10086 (n6245, n_522, n_4123);
  and g10087 (n6246, n_4124, n6245);
  not g10088 (n_4129, n6244);
  not g10089 (n_4130, n6246);
  and g10090 (n6247, n_4129, n_4130);
  not g10091 (n_4131, n6237);
  not g10092 (n_4132, n6247);
  and g10093 (n6248, n_4131, n_4132);
  not g10094 (n_4133, n6248);
  and g10095 (n6249, \asqrt[56] , n_4133);
  and g10099 (n6253, n_3875, n_3874);
  and g10100 (n6254, \asqrt[33] , n6253);
  not g10101 (n_4134, n6254);
  and g10102 (n6255, n_3873, n_4134);
  not g10103 (n_4135, n6252);
  not g10104 (n_4136, n6255);
  and g10105 (n6256, n_4135, n_4136);
  and g10106 (n6257, n_434, n_4131);
  and g10107 (n6258, n_4132, n6257);
  not g10108 (n_4137, n6256);
  not g10109 (n_4138, n6258);
  and g10110 (n6259, n_4137, n_4138);
  not g10111 (n_4139, n6249);
  not g10112 (n_4140, n6259);
  and g10113 (n6260, n_4139, n_4140);
  not g10114 (n_4141, n6260);
  and g10115 (n6261, \asqrt[57] , n_4141);
  and g10119 (n6265, n_3883, n_3882);
  and g10120 (n6266, \asqrt[33] , n6265);
  not g10121 (n_4142, n6266);
  and g10122 (n6267, n_3881, n_4142);
  not g10123 (n_4143, n6264);
  not g10124 (n_4144, n6267);
  and g10125 (n6268, n_4143, n_4144);
  and g10126 (n6269, n_354, n_4139);
  and g10127 (n6270, n_4140, n6269);
  not g10128 (n_4145, n6268);
  not g10129 (n_4146, n6270);
  and g10130 (n6271, n_4145, n_4146);
  not g10131 (n_4147, n6261);
  not g10132 (n_4148, n6271);
  and g10133 (n6272, n_4147, n_4148);
  not g10134 (n_4149, n6272);
  and g10135 (n6273, \asqrt[58] , n_4149);
  and g10139 (n6277, n_3891, n_3890);
  and g10140 (n6278, \asqrt[33] , n6277);
  not g10141 (n_4150, n6278);
  and g10142 (n6279, n_3889, n_4150);
  not g10143 (n_4151, n6276);
  not g10144 (n_4152, n6279);
  and g10145 (n6280, n_4151, n_4152);
  and g10146 (n6281, n_282, n_4147);
  and g10147 (n6282, n_4148, n6281);
  not g10148 (n_4153, n6280);
  not g10149 (n_4154, n6282);
  and g10150 (n6283, n_4153, n_4154);
  not g10151 (n_4155, n6273);
  not g10152 (n_4156, n6283);
  and g10153 (n6284, n_4155, n_4156);
  not g10154 (n_4157, n6284);
  and g10155 (n6285, \asqrt[59] , n_4157);
  and g10159 (n6289, n_3899, n_3898);
  and g10160 (n6290, \asqrt[33] , n6289);
  not g10161 (n_4158, n6290);
  and g10162 (n6291, n_3897, n_4158);
  not g10163 (n_4159, n6288);
  not g10164 (n_4160, n6291);
  and g10165 (n6292, n_4159, n_4160);
  and g10166 (n6293, n_218, n_4155);
  and g10167 (n6294, n_4156, n6293);
  not g10168 (n_4161, n6292);
  not g10169 (n_4162, n6294);
  and g10170 (n6295, n_4161, n_4162);
  not g10171 (n_4163, n6285);
  not g10172 (n_4164, n6295);
  and g10173 (n6296, n_4163, n_4164);
  not g10174 (n_4165, n6296);
  and g10175 (n6297, \asqrt[60] , n_4165);
  and g10179 (n6301, n_3907, n_3906);
  and g10180 (n6302, \asqrt[33] , n6301);
  not g10181 (n_4166, n6302);
  and g10182 (n6303, n_3905, n_4166);
  not g10183 (n_4167, n6300);
  not g10184 (n_4168, n6303);
  and g10185 (n6304, n_4167, n_4168);
  and g10186 (n6305, n_162, n_4163);
  and g10187 (n6306, n_4164, n6305);
  not g10188 (n_4169, n6304);
  not g10189 (n_4170, n6306);
  and g10190 (n6307, n_4169, n_4170);
  not g10191 (n_4171, n6297);
  not g10192 (n_4172, n6307);
  and g10193 (n6308, n_4171, n_4172);
  not g10194 (n_4173, n6308);
  and g10195 (n6309, \asqrt[61] , n_4173);
  and g10199 (n6313, n_3915, n_3914);
  and g10200 (n6314, \asqrt[33] , n6313);
  not g10201 (n_4174, n6314);
  and g10202 (n6315, n_3913, n_4174);
  not g10203 (n_4175, n6312);
  not g10204 (n_4176, n6315);
  and g10205 (n6316, n_4175, n_4176);
  and g10206 (n6317, n_115, n_4171);
  and g10207 (n6318, n_4172, n6317);
  not g10208 (n_4177, n6316);
  not g10209 (n_4178, n6318);
  and g10210 (n6319, n_4177, n_4178);
  not g10211 (n_4179, n6309);
  not g10212 (n_4180, n6319);
  and g10213 (n6320, n_4179, n_4180);
  not g10214 (n_4181, n6320);
  and g10215 (n6321, \asqrt[62] , n_4181);
  and g10219 (n6325, n_3923, n_3922);
  and g10220 (n6326, \asqrt[33] , n6325);
  not g10221 (n_4182, n6326);
  and g10222 (n6327, n_3921, n_4182);
  not g10223 (n_4183, n6324);
  not g10224 (n_4184, n6327);
  and g10225 (n6328, n_4183, n_4184);
  and g10226 (n6329, n_76, n_4179);
  and g10227 (n6330, n_4180, n6329);
  not g10228 (n_4185, n6328);
  not g10229 (n_4186, n6330);
  and g10230 (n6331, n_4185, n_4186);
  not g10231 (n_4187, n6321);
  not g10232 (n_4188, n6331);
  and g10233 (n6332, n_4187, n_4188);
  and g10237 (n6336, n_3931, n_3930);
  and g10238 (n6337, \asqrt[33] , n6336);
  not g10239 (n_4189, n6337);
  and g10240 (n6338, n_3929, n_4189);
  not g10241 (n_4190, n6335);
  not g10242 (n_4191, n6338);
  and g10243 (n6339, n_4190, n_4191);
  and g10244 (n6340, n_3938, n_3937);
  and g10245 (n6341, \asqrt[33] , n6340);
  not g10248 (n_4193, n6339);
  not g10250 (n_4194, n6332);
  not g10252 (n_4195, n6344);
  and g10253 (n6345, n_21, n_4195);
  and g10254 (n6346, n_4187, n6339);
  and g10255 (n6347, n_4188, n6346);
  and g10256 (n6348, n_3937, \asqrt[33] );
  not g10257 (n_4196, n6348);
  and g10258 (n6349, n5952, n_4196);
  not g10259 (n_4197, n6340);
  and g10260 (n6350, \asqrt[63] , n_4197);
  not g10261 (n_4198, n6349);
  and g10262 (n6351, n_4198, n6350);
  not g10268 (n_4199, n6351);
  not g10269 (n_4200, n6356);
  not g10271 (n_4201, n6347);
  and g10275 (n6360, \a[64] , \asqrt[32] );
  not g10276 (n_4206, \a[62] );
  not g10277 (n_4207, \a[63] );
  and g10278 (n6361, n_4206, n_4207);
  and g10279 (n6362, n_3950, n6361);
  not g10280 (n_4208, n6360);
  not g10281 (n_4209, n6362);
  and g10282 (n6363, n_4208, n_4209);
  not g10283 (n_4210, n6363);
  and g10284 (n6364, \asqrt[33] , n_4210);
  and g10285 (n6365, n_3950, \asqrt[32] );
  not g10286 (n_4211, n6365);
  and g10287 (n6366, \a[65] , n_4211);
  and g10288 (n6367, n5981, \asqrt[32] );
  not g10289 (n_4212, n6366);
  not g10290 (n_4213, n6367);
  and g10291 (n6368, n_4212, n_4213);
  not g10297 (n_4214, n6373);
  and g10298 (n6374, n6368, n_4214);
  not g10299 (n_4215, n6364);
  not g10300 (n_4216, n6374);
  and g10301 (n6375, n_4215, n_4216);
  not g10302 (n_4217, n6375);
  and g10303 (n6376, \asqrt[34] , n_4217);
  not g10304 (n_4218, \asqrt[34] );
  and g10305 (n6377, n_4218, n_4215);
  and g10306 (n6378, n_4216, n6377);
  not g10310 (n_4219, n6345);
  not g10312 (n_4220, n6382);
  and g10313 (n6383, n_4213, n_4220);
  not g10314 (n_4221, n6383);
  and g10315 (n6384, \a[66] , n_4221);
  and g10316 (n6385, n_3702, n_4220);
  and g10317 (n6386, n_4213, n6385);
  not g10318 (n_4222, n6384);
  not g10319 (n_4223, n6386);
  and g10320 (n6387, n_4222, n_4223);
  not g10321 (n_4224, n6378);
  not g10322 (n_4225, n6387);
  and g10323 (n6388, n_4224, n_4225);
  not g10324 (n_4226, n6376);
  not g10325 (n_4227, n6388);
  and g10326 (n6389, n_4226, n_4227);
  not g10327 (n_4228, n6389);
  and g10328 (n6390, \asqrt[35] , n_4228);
  and g10329 (n6391, n_3959, n_3958);
  not g10330 (n_4229, n5993);
  and g10331 (n6392, n_4229, n6391);
  and g10332 (n6393, \asqrt[32] , n6392);
  and g10333 (n6394, \asqrt[32] , n6391);
  not g10334 (n_4230, n6394);
  and g10335 (n6395, n5993, n_4230);
  not g10336 (n_4231, n6393);
  not g10337 (n_4232, n6395);
  and g10338 (n6396, n_4231, n_4232);
  and g10339 (n6397, n_3962, n_4226);
  and g10340 (n6398, n_4227, n6397);
  not g10341 (n_4233, n6396);
  not g10342 (n_4234, n6398);
  and g10343 (n6399, n_4233, n_4234);
  not g10344 (n_4235, n6390);
  not g10345 (n_4236, n6399);
  and g10346 (n6400, n_4235, n_4236);
  not g10347 (n_4237, n6400);
  and g10348 (n6401, \asqrt[36] , n_4237);
  and g10352 (n6405, n_3970, n_3968);
  and g10353 (n6406, \asqrt[32] , n6405);
  not g10354 (n_4238, n6406);
  and g10355 (n6407, n_3969, n_4238);
  not g10356 (n_4239, n6404);
  not g10357 (n_4240, n6407);
  and g10358 (n6408, n_4239, n_4240);
  and g10359 (n6409, n_3714, n_4235);
  and g10360 (n6410, n_4236, n6409);
  not g10361 (n_4241, n6408);
  not g10362 (n_4242, n6410);
  and g10363 (n6411, n_4241, n_4242);
  not g10364 (n_4243, n6401);
  not g10365 (n_4244, n6411);
  and g10366 (n6412, n_4243, n_4244);
  not g10367 (n_4245, n6412);
  and g10368 (n6413, \asqrt[37] , n_4245);
  and g10372 (n6417, n_3979, n_3978);
  and g10373 (n6418, \asqrt[32] , n6417);
  not g10374 (n_4246, n6418);
  and g10375 (n6419, n_3977, n_4246);
  not g10376 (n_4247, n6416);
  not g10377 (n_4248, n6419);
  and g10378 (n6420, n_4247, n_4248);
  and g10379 (n6421, n_3474, n_4243);
  and g10380 (n6422, n_4244, n6421);
  not g10381 (n_4249, n6420);
  not g10382 (n_4250, n6422);
  and g10383 (n6423, n_4249, n_4250);
  not g10384 (n_4251, n6413);
  not g10385 (n_4252, n6423);
  and g10386 (n6424, n_4251, n_4252);
  not g10387 (n_4253, n6424);
  and g10388 (n6425, \asqrt[38] , n_4253);
  and g10392 (n6429, n_3987, n_3986);
  and g10393 (n6430, \asqrt[32] , n6429);
  not g10394 (n_4254, n6430);
  and g10395 (n6431, n_3985, n_4254);
  not g10396 (n_4255, n6428);
  not g10397 (n_4256, n6431);
  and g10398 (n6432, n_4255, n_4256);
  and g10399 (n6433, n_3242, n_4251);
  and g10400 (n6434, n_4252, n6433);
  not g10401 (n_4257, n6432);
  not g10402 (n_4258, n6434);
  and g10403 (n6435, n_4257, n_4258);
  not g10404 (n_4259, n6425);
  not g10405 (n_4260, n6435);
  and g10406 (n6436, n_4259, n_4260);
  not g10407 (n_4261, n6436);
  and g10408 (n6437, \asqrt[39] , n_4261);
  and g10412 (n6441, n_3995, n_3994);
  and g10413 (n6442, \asqrt[32] , n6441);
  not g10414 (n_4262, n6442);
  and g10415 (n6443, n_3993, n_4262);
  not g10416 (n_4263, n6440);
  not g10417 (n_4264, n6443);
  and g10418 (n6444, n_4263, n_4264);
  and g10419 (n6445, n_3018, n_4259);
  and g10420 (n6446, n_4260, n6445);
  not g10421 (n_4265, n6444);
  not g10422 (n_4266, n6446);
  and g10423 (n6447, n_4265, n_4266);
  not g10424 (n_4267, n6437);
  not g10425 (n_4268, n6447);
  and g10426 (n6448, n_4267, n_4268);
  not g10427 (n_4269, n6448);
  and g10428 (n6449, \asqrt[40] , n_4269);
  and g10432 (n6453, n_4003, n_4002);
  and g10433 (n6454, \asqrt[32] , n6453);
  not g10434 (n_4270, n6454);
  and g10435 (n6455, n_4001, n_4270);
  not g10436 (n_4271, n6452);
  not g10437 (n_4272, n6455);
  and g10438 (n6456, n_4271, n_4272);
  and g10439 (n6457, n_2802, n_4267);
  and g10440 (n6458, n_4268, n6457);
  not g10441 (n_4273, n6456);
  not g10442 (n_4274, n6458);
  and g10443 (n6459, n_4273, n_4274);
  not g10444 (n_4275, n6449);
  not g10445 (n_4276, n6459);
  and g10446 (n6460, n_4275, n_4276);
  not g10447 (n_4277, n6460);
  and g10448 (n6461, \asqrt[41] , n_4277);
  and g10452 (n6465, n_4011, n_4010);
  and g10453 (n6466, \asqrt[32] , n6465);
  not g10454 (n_4278, n6466);
  and g10455 (n6467, n_4009, n_4278);
  not g10456 (n_4279, n6464);
  not g10457 (n_4280, n6467);
  and g10458 (n6468, n_4279, n_4280);
  and g10459 (n6469, n_2594, n_4275);
  and g10460 (n6470, n_4276, n6469);
  not g10461 (n_4281, n6468);
  not g10462 (n_4282, n6470);
  and g10463 (n6471, n_4281, n_4282);
  not g10464 (n_4283, n6461);
  not g10465 (n_4284, n6471);
  and g10466 (n6472, n_4283, n_4284);
  not g10467 (n_4285, n6472);
  and g10468 (n6473, \asqrt[42] , n_4285);
  and g10472 (n6477, n_4019, n_4018);
  and g10473 (n6478, \asqrt[32] , n6477);
  not g10474 (n_4286, n6478);
  and g10475 (n6479, n_4017, n_4286);
  not g10476 (n_4287, n6476);
  not g10477 (n_4288, n6479);
  and g10478 (n6480, n_4287, n_4288);
  and g10479 (n6481, n_2394, n_4283);
  and g10480 (n6482, n_4284, n6481);
  not g10481 (n_4289, n6480);
  not g10482 (n_4290, n6482);
  and g10483 (n6483, n_4289, n_4290);
  not g10484 (n_4291, n6473);
  not g10485 (n_4292, n6483);
  and g10486 (n6484, n_4291, n_4292);
  not g10487 (n_4293, n6484);
  and g10488 (n6485, \asqrt[43] , n_4293);
  and g10492 (n6489, n_4027, n_4026);
  and g10493 (n6490, \asqrt[32] , n6489);
  not g10494 (n_4294, n6490);
  and g10495 (n6491, n_4025, n_4294);
  not g10496 (n_4295, n6488);
  not g10497 (n_4296, n6491);
  and g10498 (n6492, n_4295, n_4296);
  and g10499 (n6493, n_2202, n_4291);
  and g10500 (n6494, n_4292, n6493);
  not g10501 (n_4297, n6492);
  not g10502 (n_4298, n6494);
  and g10503 (n6495, n_4297, n_4298);
  not g10504 (n_4299, n6485);
  not g10505 (n_4300, n6495);
  and g10506 (n6496, n_4299, n_4300);
  not g10507 (n_4301, n6496);
  and g10508 (n6497, \asqrt[44] , n_4301);
  and g10512 (n6501, n_4035, n_4034);
  and g10513 (n6502, \asqrt[32] , n6501);
  not g10514 (n_4302, n6502);
  and g10515 (n6503, n_4033, n_4302);
  not g10516 (n_4303, n6500);
  not g10517 (n_4304, n6503);
  and g10518 (n6504, n_4303, n_4304);
  and g10519 (n6505, n_2018, n_4299);
  and g10520 (n6506, n_4300, n6505);
  not g10521 (n_4305, n6504);
  not g10522 (n_4306, n6506);
  and g10523 (n6507, n_4305, n_4306);
  not g10524 (n_4307, n6497);
  not g10525 (n_4308, n6507);
  and g10526 (n6508, n_4307, n_4308);
  not g10527 (n_4309, n6508);
  and g10528 (n6509, \asqrt[45] , n_4309);
  and g10532 (n6513, n_4043, n_4042);
  and g10533 (n6514, \asqrt[32] , n6513);
  not g10534 (n_4310, n6514);
  and g10535 (n6515, n_4041, n_4310);
  not g10536 (n_4311, n6512);
  not g10537 (n_4312, n6515);
  and g10538 (n6516, n_4311, n_4312);
  and g10539 (n6517, n_1842, n_4307);
  and g10540 (n6518, n_4308, n6517);
  not g10541 (n_4313, n6516);
  not g10542 (n_4314, n6518);
  and g10543 (n6519, n_4313, n_4314);
  not g10544 (n_4315, n6509);
  not g10545 (n_4316, n6519);
  and g10546 (n6520, n_4315, n_4316);
  not g10547 (n_4317, n6520);
  and g10548 (n6521, \asqrt[46] , n_4317);
  and g10552 (n6525, n_4051, n_4050);
  and g10553 (n6526, \asqrt[32] , n6525);
  not g10554 (n_4318, n6526);
  and g10555 (n6527, n_4049, n_4318);
  not g10556 (n_4319, n6524);
  not g10557 (n_4320, n6527);
  and g10558 (n6528, n_4319, n_4320);
  and g10559 (n6529, n_1674, n_4315);
  and g10560 (n6530, n_4316, n6529);
  not g10561 (n_4321, n6528);
  not g10562 (n_4322, n6530);
  and g10563 (n6531, n_4321, n_4322);
  not g10564 (n_4323, n6521);
  not g10565 (n_4324, n6531);
  and g10566 (n6532, n_4323, n_4324);
  not g10567 (n_4325, n6532);
  and g10568 (n6533, \asqrt[47] , n_4325);
  and g10572 (n6537, n_4059, n_4058);
  and g10573 (n6538, \asqrt[32] , n6537);
  not g10574 (n_4326, n6538);
  and g10575 (n6539, n_4057, n_4326);
  not g10576 (n_4327, n6536);
  not g10577 (n_4328, n6539);
  and g10578 (n6540, n_4327, n_4328);
  and g10579 (n6541, n_1514, n_4323);
  and g10580 (n6542, n_4324, n6541);
  not g10581 (n_4329, n6540);
  not g10582 (n_4330, n6542);
  and g10583 (n6543, n_4329, n_4330);
  not g10584 (n_4331, n6533);
  not g10585 (n_4332, n6543);
  and g10586 (n6544, n_4331, n_4332);
  not g10587 (n_4333, n6544);
  and g10588 (n6545, \asqrt[48] , n_4333);
  and g10592 (n6549, n_4067, n_4066);
  and g10593 (n6550, \asqrt[32] , n6549);
  not g10594 (n_4334, n6550);
  and g10595 (n6551, n_4065, n_4334);
  not g10596 (n_4335, n6548);
  not g10597 (n_4336, n6551);
  and g10598 (n6552, n_4335, n_4336);
  and g10599 (n6553, n_1362, n_4331);
  and g10600 (n6554, n_4332, n6553);
  not g10601 (n_4337, n6552);
  not g10602 (n_4338, n6554);
  and g10603 (n6555, n_4337, n_4338);
  not g10604 (n_4339, n6545);
  not g10605 (n_4340, n6555);
  and g10606 (n6556, n_4339, n_4340);
  not g10607 (n_4341, n6556);
  and g10608 (n6557, \asqrt[49] , n_4341);
  and g10612 (n6561, n_4075, n_4074);
  and g10613 (n6562, \asqrt[32] , n6561);
  not g10614 (n_4342, n6562);
  and g10615 (n6563, n_4073, n_4342);
  not g10616 (n_4343, n6560);
  not g10617 (n_4344, n6563);
  and g10618 (n6564, n_4343, n_4344);
  and g10619 (n6565, n_1218, n_4339);
  and g10620 (n6566, n_4340, n6565);
  not g10621 (n_4345, n6564);
  not g10622 (n_4346, n6566);
  and g10623 (n6567, n_4345, n_4346);
  not g10624 (n_4347, n6557);
  not g10625 (n_4348, n6567);
  and g10626 (n6568, n_4347, n_4348);
  not g10627 (n_4349, n6568);
  and g10628 (n6569, \asqrt[50] , n_4349);
  and g10632 (n6573, n_4083, n_4082);
  and g10633 (n6574, \asqrt[32] , n6573);
  not g10634 (n_4350, n6574);
  and g10635 (n6575, n_4081, n_4350);
  not g10636 (n_4351, n6572);
  not g10637 (n_4352, n6575);
  and g10638 (n6576, n_4351, n_4352);
  and g10639 (n6577, n_1082, n_4347);
  and g10640 (n6578, n_4348, n6577);
  not g10641 (n_4353, n6576);
  not g10642 (n_4354, n6578);
  and g10643 (n6579, n_4353, n_4354);
  not g10644 (n_4355, n6569);
  not g10645 (n_4356, n6579);
  and g10646 (n6580, n_4355, n_4356);
  not g10647 (n_4357, n6580);
  and g10648 (n6581, \asqrt[51] , n_4357);
  and g10652 (n6585, n_4091, n_4090);
  and g10653 (n6586, \asqrt[32] , n6585);
  not g10654 (n_4358, n6586);
  and g10655 (n6587, n_4089, n_4358);
  not g10656 (n_4359, n6584);
  not g10657 (n_4360, n6587);
  and g10658 (n6588, n_4359, n_4360);
  and g10659 (n6589, n_954, n_4355);
  and g10660 (n6590, n_4356, n6589);
  not g10661 (n_4361, n6588);
  not g10662 (n_4362, n6590);
  and g10663 (n6591, n_4361, n_4362);
  not g10664 (n_4363, n6581);
  not g10665 (n_4364, n6591);
  and g10666 (n6592, n_4363, n_4364);
  not g10667 (n_4365, n6592);
  and g10668 (n6593, \asqrt[52] , n_4365);
  and g10672 (n6597, n_4099, n_4098);
  and g10673 (n6598, \asqrt[32] , n6597);
  not g10674 (n_4366, n6598);
  and g10675 (n6599, n_4097, n_4366);
  not g10676 (n_4367, n6596);
  not g10677 (n_4368, n6599);
  and g10678 (n6600, n_4367, n_4368);
  and g10679 (n6601, n_834, n_4363);
  and g10680 (n6602, n_4364, n6601);
  not g10681 (n_4369, n6600);
  not g10682 (n_4370, n6602);
  and g10683 (n6603, n_4369, n_4370);
  not g10684 (n_4371, n6593);
  not g10685 (n_4372, n6603);
  and g10686 (n6604, n_4371, n_4372);
  not g10687 (n_4373, n6604);
  and g10688 (n6605, \asqrt[53] , n_4373);
  and g10692 (n6609, n_4107, n_4106);
  and g10693 (n6610, \asqrt[32] , n6609);
  not g10694 (n_4374, n6610);
  and g10695 (n6611, n_4105, n_4374);
  not g10696 (n_4375, n6608);
  not g10697 (n_4376, n6611);
  and g10698 (n6612, n_4375, n_4376);
  and g10699 (n6613, n_722, n_4371);
  and g10700 (n6614, n_4372, n6613);
  not g10701 (n_4377, n6612);
  not g10702 (n_4378, n6614);
  and g10703 (n6615, n_4377, n_4378);
  not g10704 (n_4379, n6605);
  not g10705 (n_4380, n6615);
  and g10706 (n6616, n_4379, n_4380);
  not g10707 (n_4381, n6616);
  and g10708 (n6617, \asqrt[54] , n_4381);
  and g10712 (n6621, n_4115, n_4114);
  and g10713 (n6622, \asqrt[32] , n6621);
  not g10714 (n_4382, n6622);
  and g10715 (n6623, n_4113, n_4382);
  not g10716 (n_4383, n6620);
  not g10717 (n_4384, n6623);
  and g10718 (n6624, n_4383, n_4384);
  and g10719 (n6625, n_618, n_4379);
  and g10720 (n6626, n_4380, n6625);
  not g10721 (n_4385, n6624);
  not g10722 (n_4386, n6626);
  and g10723 (n6627, n_4385, n_4386);
  not g10724 (n_4387, n6617);
  not g10725 (n_4388, n6627);
  and g10726 (n6628, n_4387, n_4388);
  not g10727 (n_4389, n6628);
  and g10728 (n6629, \asqrt[55] , n_4389);
  and g10732 (n6633, n_4123, n_4122);
  and g10733 (n6634, \asqrt[32] , n6633);
  not g10734 (n_4390, n6634);
  and g10735 (n6635, n_4121, n_4390);
  not g10736 (n_4391, n6632);
  not g10737 (n_4392, n6635);
  and g10738 (n6636, n_4391, n_4392);
  and g10739 (n6637, n_522, n_4387);
  and g10740 (n6638, n_4388, n6637);
  not g10741 (n_4393, n6636);
  not g10742 (n_4394, n6638);
  and g10743 (n6639, n_4393, n_4394);
  not g10744 (n_4395, n6629);
  not g10745 (n_4396, n6639);
  and g10746 (n6640, n_4395, n_4396);
  not g10747 (n_4397, n6640);
  and g10748 (n6641, \asqrt[56] , n_4397);
  and g10752 (n6645, n_4131, n_4130);
  and g10753 (n6646, \asqrt[32] , n6645);
  not g10754 (n_4398, n6646);
  and g10755 (n6647, n_4129, n_4398);
  not g10756 (n_4399, n6644);
  not g10757 (n_4400, n6647);
  and g10758 (n6648, n_4399, n_4400);
  and g10759 (n6649, n_434, n_4395);
  and g10760 (n6650, n_4396, n6649);
  not g10761 (n_4401, n6648);
  not g10762 (n_4402, n6650);
  and g10763 (n6651, n_4401, n_4402);
  not g10764 (n_4403, n6641);
  not g10765 (n_4404, n6651);
  and g10766 (n6652, n_4403, n_4404);
  not g10767 (n_4405, n6652);
  and g10768 (n6653, \asqrt[57] , n_4405);
  and g10772 (n6657, n_4139, n_4138);
  and g10773 (n6658, \asqrt[32] , n6657);
  not g10774 (n_4406, n6658);
  and g10775 (n6659, n_4137, n_4406);
  not g10776 (n_4407, n6656);
  not g10777 (n_4408, n6659);
  and g10778 (n6660, n_4407, n_4408);
  and g10779 (n6661, n_354, n_4403);
  and g10780 (n6662, n_4404, n6661);
  not g10781 (n_4409, n6660);
  not g10782 (n_4410, n6662);
  and g10783 (n6663, n_4409, n_4410);
  not g10784 (n_4411, n6653);
  not g10785 (n_4412, n6663);
  and g10786 (n6664, n_4411, n_4412);
  not g10787 (n_4413, n6664);
  and g10788 (n6665, \asqrt[58] , n_4413);
  and g10792 (n6669, n_4147, n_4146);
  and g10793 (n6670, \asqrt[32] , n6669);
  not g10794 (n_4414, n6670);
  and g10795 (n6671, n_4145, n_4414);
  not g10796 (n_4415, n6668);
  not g10797 (n_4416, n6671);
  and g10798 (n6672, n_4415, n_4416);
  and g10799 (n6673, n_282, n_4411);
  and g10800 (n6674, n_4412, n6673);
  not g10801 (n_4417, n6672);
  not g10802 (n_4418, n6674);
  and g10803 (n6675, n_4417, n_4418);
  not g10804 (n_4419, n6665);
  not g10805 (n_4420, n6675);
  and g10806 (n6676, n_4419, n_4420);
  not g10807 (n_4421, n6676);
  and g10808 (n6677, \asqrt[59] , n_4421);
  and g10812 (n6681, n_4155, n_4154);
  and g10813 (n6682, \asqrt[32] , n6681);
  not g10814 (n_4422, n6682);
  and g10815 (n6683, n_4153, n_4422);
  not g10816 (n_4423, n6680);
  not g10817 (n_4424, n6683);
  and g10818 (n6684, n_4423, n_4424);
  and g10819 (n6685, n_218, n_4419);
  and g10820 (n6686, n_4420, n6685);
  not g10821 (n_4425, n6684);
  not g10822 (n_4426, n6686);
  and g10823 (n6687, n_4425, n_4426);
  not g10824 (n_4427, n6677);
  not g10825 (n_4428, n6687);
  and g10826 (n6688, n_4427, n_4428);
  not g10827 (n_4429, n6688);
  and g10828 (n6689, \asqrt[60] , n_4429);
  and g10832 (n6693, n_4163, n_4162);
  and g10833 (n6694, \asqrt[32] , n6693);
  not g10834 (n_4430, n6694);
  and g10835 (n6695, n_4161, n_4430);
  not g10836 (n_4431, n6692);
  not g10837 (n_4432, n6695);
  and g10838 (n6696, n_4431, n_4432);
  and g10839 (n6697, n_162, n_4427);
  and g10840 (n6698, n_4428, n6697);
  not g10841 (n_4433, n6696);
  not g10842 (n_4434, n6698);
  and g10843 (n6699, n_4433, n_4434);
  not g10844 (n_4435, n6689);
  not g10845 (n_4436, n6699);
  and g10846 (n6700, n_4435, n_4436);
  not g10847 (n_4437, n6700);
  and g10848 (n6701, \asqrt[61] , n_4437);
  and g10852 (n6705, n_4171, n_4170);
  and g10853 (n6706, \asqrt[32] , n6705);
  not g10854 (n_4438, n6706);
  and g10855 (n6707, n_4169, n_4438);
  not g10856 (n_4439, n6704);
  not g10857 (n_4440, n6707);
  and g10858 (n6708, n_4439, n_4440);
  and g10859 (n6709, n_115, n_4435);
  and g10860 (n6710, n_4436, n6709);
  not g10861 (n_4441, n6708);
  not g10862 (n_4442, n6710);
  and g10863 (n6711, n_4441, n_4442);
  not g10864 (n_4443, n6701);
  not g10865 (n_4444, n6711);
  and g10866 (n6712, n_4443, n_4444);
  not g10867 (n_4445, n6712);
  and g10868 (n6713, \asqrt[62] , n_4445);
  and g10872 (n6717, n_4179, n_4178);
  and g10873 (n6718, \asqrt[32] , n6717);
  not g10874 (n_4446, n6718);
  and g10875 (n6719, n_4177, n_4446);
  not g10876 (n_4447, n6716);
  not g10877 (n_4448, n6719);
  and g10878 (n6720, n_4447, n_4448);
  and g10879 (n6721, n_76, n_4443);
  and g10880 (n6722, n_4444, n6721);
  not g10881 (n_4449, n6720);
  not g10882 (n_4450, n6722);
  and g10883 (n6723, n_4449, n_4450);
  not g10884 (n_4451, n6713);
  not g10885 (n_4452, n6723);
  and g10886 (n6724, n_4451, n_4452);
  and g10890 (n6728, n_4187, n_4186);
  and g10891 (n6729, \asqrt[32] , n6728);
  not g10892 (n_4453, n6729);
  and g10893 (n6730, n_4185, n_4453);
  not g10894 (n_4454, n6727);
  not g10895 (n_4455, n6730);
  and g10896 (n6731, n_4454, n_4455);
  and g10897 (n6732, n_4194, n_4193);
  and g10898 (n6733, \asqrt[32] , n6732);
  not g10901 (n_4457, n6731);
  not g10903 (n_4458, n6724);
  not g10905 (n_4459, n6736);
  and g10906 (n6737, n_21, n_4459);
  and g10907 (n6738, n_4451, n6731);
  and g10908 (n6739, n_4452, n6738);
  and g10909 (n6740, n_4193, \asqrt[32] );
  not g10910 (n_4460, n6740);
  and g10911 (n6741, n6332, n_4460);
  not g10912 (n_4461, n6732);
  and g10913 (n6742, \asqrt[63] , n_4461);
  not g10914 (n_4462, n6741);
  and g10915 (n6743, n_4462, n6742);
  not g10921 (n_4463, n6743);
  not g10922 (n_4464, n6748);
  not g10924 (n_4465, n6739);
  and g10928 (n6752, \a[62] , \asqrt[31] );
  not g10929 (n_4470, \a[60] );
  not g10930 (n_4471, \a[61] );
  and g10931 (n6753, n_4470, n_4471);
  and g10932 (n6754, n_4206, n6753);
  not g10933 (n_4472, n6752);
  not g10934 (n_4473, n6754);
  and g10935 (n6755, n_4472, n_4473);
  not g10936 (n_4474, n6755);
  and g10937 (n6756, \asqrt[32] , n_4474);
  and g10943 (n6762, n_4206, \asqrt[31] );
  not g10944 (n_4475, n6762);
  and g10945 (n6763, \a[63] , n_4475);
  and g10946 (n6764, n6361, \asqrt[31] );
  not g10947 (n_4476, n6763);
  not g10948 (n_4477, n6764);
  and g10949 (n6765, n_4476, n_4477);
  not g10950 (n_4478, n6761);
  and g10951 (n6766, n_4478, n6765);
  not g10952 (n_4479, n6756);
  not g10953 (n_4480, n6766);
  and g10954 (n6767, n_4479, n_4480);
  not g10955 (n_4481, n6767);
  and g10956 (n6768, \asqrt[33] , n_4481);
  not g10957 (n_4482, \asqrt[33] );
  and g10958 (n6769, n_4482, n_4479);
  and g10959 (n6770, n_4480, n6769);
  not g10963 (n_4483, n6737);
  not g10965 (n_4484, n6774);
  and g10966 (n6775, n_4477, n_4484);
  not g10967 (n_4485, n6775);
  and g10968 (n6776, \a[64] , n_4485);
  and g10969 (n6777, n_3950, n_4484);
  and g10970 (n6778, n_4477, n6777);
  not g10971 (n_4486, n6776);
  not g10972 (n_4487, n6778);
  and g10973 (n6779, n_4486, n_4487);
  not g10974 (n_4488, n6770);
  not g10975 (n_4489, n6779);
  and g10976 (n6780, n_4488, n_4489);
  not g10977 (n_4490, n6768);
  not g10978 (n_4491, n6780);
  and g10979 (n6781, n_4490, n_4491);
  not g10980 (n_4492, n6781);
  and g10981 (n6782, \asqrt[34] , n_4492);
  and g10982 (n6783, n_4218, n_4490);
  and g10983 (n6784, n_4491, n6783);
  and g10988 (n6788, n_4215, n_4214);
  and g10989 (n6789, \asqrt[31] , n6788);
  not g10990 (n_4494, n6789);
  and g10991 (n6790, n6368, n_4494);
  not g10992 (n_4495, n6787);
  not g10993 (n_4496, n6790);
  and g10994 (n6791, n_4495, n_4496);
  not g10995 (n_4497, n6784);
  not g10996 (n_4498, n6791);
  and g10997 (n6792, n_4497, n_4498);
  not g10998 (n_4499, n6782);
  not g10999 (n_4500, n6792);
  and g11000 (n6793, n_4499, n_4500);
  not g11001 (n_4501, n6793);
  and g11002 (n6794, \asqrt[35] , n_4501);
  and g11006 (n6798, n_4226, n_4224);
  and g11007 (n6799, \asqrt[31] , n6798);
  not g11008 (n_4502, n6799);
  and g11009 (n6800, n_4225, n_4502);
  not g11010 (n_4503, n6797);
  not g11011 (n_4504, n6800);
  and g11012 (n6801, n_4503, n_4504);
  and g11013 (n6802, n_3962, n_4499);
  and g11014 (n6803, n_4500, n6802);
  not g11015 (n_4505, n6801);
  not g11016 (n_4506, n6803);
  and g11017 (n6804, n_4505, n_4506);
  not g11018 (n_4507, n6794);
  not g11019 (n_4508, n6804);
  and g11020 (n6805, n_4507, n_4508);
  not g11021 (n_4509, n6805);
  and g11022 (n6806, \asqrt[36] , n_4509);
  and g11026 (n6810, n_4235, n_4234);
  and g11027 (n6811, \asqrt[31] , n6810);
  not g11028 (n_4510, n6811);
  and g11029 (n6812, n_4233, n_4510);
  not g11030 (n_4511, n6809);
  not g11031 (n_4512, n6812);
  and g11032 (n6813, n_4511, n_4512);
  and g11033 (n6814, n_3714, n_4507);
  and g11034 (n6815, n_4508, n6814);
  not g11035 (n_4513, n6813);
  not g11036 (n_4514, n6815);
  and g11037 (n6816, n_4513, n_4514);
  not g11038 (n_4515, n6806);
  not g11039 (n_4516, n6816);
  and g11040 (n6817, n_4515, n_4516);
  not g11041 (n_4517, n6817);
  and g11042 (n6818, \asqrt[37] , n_4517);
  and g11046 (n6822, n_4243, n_4242);
  and g11047 (n6823, \asqrt[31] , n6822);
  not g11048 (n_4518, n6823);
  and g11049 (n6824, n_4241, n_4518);
  not g11050 (n_4519, n6821);
  not g11051 (n_4520, n6824);
  and g11052 (n6825, n_4519, n_4520);
  and g11053 (n6826, n_3474, n_4515);
  and g11054 (n6827, n_4516, n6826);
  not g11055 (n_4521, n6825);
  not g11056 (n_4522, n6827);
  and g11057 (n6828, n_4521, n_4522);
  not g11058 (n_4523, n6818);
  not g11059 (n_4524, n6828);
  and g11060 (n6829, n_4523, n_4524);
  not g11061 (n_4525, n6829);
  and g11062 (n6830, \asqrt[38] , n_4525);
  and g11066 (n6834, n_4251, n_4250);
  and g11067 (n6835, \asqrt[31] , n6834);
  not g11068 (n_4526, n6835);
  and g11069 (n6836, n_4249, n_4526);
  not g11070 (n_4527, n6833);
  not g11071 (n_4528, n6836);
  and g11072 (n6837, n_4527, n_4528);
  and g11073 (n6838, n_3242, n_4523);
  and g11074 (n6839, n_4524, n6838);
  not g11075 (n_4529, n6837);
  not g11076 (n_4530, n6839);
  and g11077 (n6840, n_4529, n_4530);
  not g11078 (n_4531, n6830);
  not g11079 (n_4532, n6840);
  and g11080 (n6841, n_4531, n_4532);
  not g11081 (n_4533, n6841);
  and g11082 (n6842, \asqrt[39] , n_4533);
  and g11086 (n6846, n_4259, n_4258);
  and g11087 (n6847, \asqrt[31] , n6846);
  not g11088 (n_4534, n6847);
  and g11089 (n6848, n_4257, n_4534);
  not g11090 (n_4535, n6845);
  not g11091 (n_4536, n6848);
  and g11092 (n6849, n_4535, n_4536);
  and g11093 (n6850, n_3018, n_4531);
  and g11094 (n6851, n_4532, n6850);
  not g11095 (n_4537, n6849);
  not g11096 (n_4538, n6851);
  and g11097 (n6852, n_4537, n_4538);
  not g11098 (n_4539, n6842);
  not g11099 (n_4540, n6852);
  and g11100 (n6853, n_4539, n_4540);
  not g11101 (n_4541, n6853);
  and g11102 (n6854, \asqrt[40] , n_4541);
  and g11106 (n6858, n_4267, n_4266);
  and g11107 (n6859, \asqrt[31] , n6858);
  not g11108 (n_4542, n6859);
  and g11109 (n6860, n_4265, n_4542);
  not g11110 (n_4543, n6857);
  not g11111 (n_4544, n6860);
  and g11112 (n6861, n_4543, n_4544);
  and g11113 (n6862, n_2802, n_4539);
  and g11114 (n6863, n_4540, n6862);
  not g11115 (n_4545, n6861);
  not g11116 (n_4546, n6863);
  and g11117 (n6864, n_4545, n_4546);
  not g11118 (n_4547, n6854);
  not g11119 (n_4548, n6864);
  and g11120 (n6865, n_4547, n_4548);
  not g11121 (n_4549, n6865);
  and g11122 (n6866, \asqrt[41] , n_4549);
  and g11126 (n6870, n_4275, n_4274);
  and g11127 (n6871, \asqrt[31] , n6870);
  not g11128 (n_4550, n6871);
  and g11129 (n6872, n_4273, n_4550);
  not g11130 (n_4551, n6869);
  not g11131 (n_4552, n6872);
  and g11132 (n6873, n_4551, n_4552);
  and g11133 (n6874, n_2594, n_4547);
  and g11134 (n6875, n_4548, n6874);
  not g11135 (n_4553, n6873);
  not g11136 (n_4554, n6875);
  and g11137 (n6876, n_4553, n_4554);
  not g11138 (n_4555, n6866);
  not g11139 (n_4556, n6876);
  and g11140 (n6877, n_4555, n_4556);
  not g11141 (n_4557, n6877);
  and g11142 (n6878, \asqrt[42] , n_4557);
  and g11146 (n6882, n_4283, n_4282);
  and g11147 (n6883, \asqrt[31] , n6882);
  not g11148 (n_4558, n6883);
  and g11149 (n6884, n_4281, n_4558);
  not g11150 (n_4559, n6881);
  not g11151 (n_4560, n6884);
  and g11152 (n6885, n_4559, n_4560);
  and g11153 (n6886, n_2394, n_4555);
  and g11154 (n6887, n_4556, n6886);
  not g11155 (n_4561, n6885);
  not g11156 (n_4562, n6887);
  and g11157 (n6888, n_4561, n_4562);
  not g11158 (n_4563, n6878);
  not g11159 (n_4564, n6888);
  and g11160 (n6889, n_4563, n_4564);
  not g11161 (n_4565, n6889);
  and g11162 (n6890, \asqrt[43] , n_4565);
  and g11166 (n6894, n_4291, n_4290);
  and g11167 (n6895, \asqrt[31] , n6894);
  not g11168 (n_4566, n6895);
  and g11169 (n6896, n_4289, n_4566);
  not g11170 (n_4567, n6893);
  not g11171 (n_4568, n6896);
  and g11172 (n6897, n_4567, n_4568);
  and g11173 (n6898, n_2202, n_4563);
  and g11174 (n6899, n_4564, n6898);
  not g11175 (n_4569, n6897);
  not g11176 (n_4570, n6899);
  and g11177 (n6900, n_4569, n_4570);
  not g11178 (n_4571, n6890);
  not g11179 (n_4572, n6900);
  and g11180 (n6901, n_4571, n_4572);
  not g11181 (n_4573, n6901);
  and g11182 (n6902, \asqrt[44] , n_4573);
  and g11186 (n6906, n_4299, n_4298);
  and g11187 (n6907, \asqrt[31] , n6906);
  not g11188 (n_4574, n6907);
  and g11189 (n6908, n_4297, n_4574);
  not g11190 (n_4575, n6905);
  not g11191 (n_4576, n6908);
  and g11192 (n6909, n_4575, n_4576);
  and g11193 (n6910, n_2018, n_4571);
  and g11194 (n6911, n_4572, n6910);
  not g11195 (n_4577, n6909);
  not g11196 (n_4578, n6911);
  and g11197 (n6912, n_4577, n_4578);
  not g11198 (n_4579, n6902);
  not g11199 (n_4580, n6912);
  and g11200 (n6913, n_4579, n_4580);
  not g11201 (n_4581, n6913);
  and g11202 (n6914, \asqrt[45] , n_4581);
  and g11206 (n6918, n_4307, n_4306);
  and g11207 (n6919, \asqrt[31] , n6918);
  not g11208 (n_4582, n6919);
  and g11209 (n6920, n_4305, n_4582);
  not g11210 (n_4583, n6917);
  not g11211 (n_4584, n6920);
  and g11212 (n6921, n_4583, n_4584);
  and g11213 (n6922, n_1842, n_4579);
  and g11214 (n6923, n_4580, n6922);
  not g11215 (n_4585, n6921);
  not g11216 (n_4586, n6923);
  and g11217 (n6924, n_4585, n_4586);
  not g11218 (n_4587, n6914);
  not g11219 (n_4588, n6924);
  and g11220 (n6925, n_4587, n_4588);
  not g11221 (n_4589, n6925);
  and g11222 (n6926, \asqrt[46] , n_4589);
  and g11226 (n6930, n_4315, n_4314);
  and g11227 (n6931, \asqrt[31] , n6930);
  not g11228 (n_4590, n6931);
  and g11229 (n6932, n_4313, n_4590);
  not g11230 (n_4591, n6929);
  not g11231 (n_4592, n6932);
  and g11232 (n6933, n_4591, n_4592);
  and g11233 (n6934, n_1674, n_4587);
  and g11234 (n6935, n_4588, n6934);
  not g11235 (n_4593, n6933);
  not g11236 (n_4594, n6935);
  and g11237 (n6936, n_4593, n_4594);
  not g11238 (n_4595, n6926);
  not g11239 (n_4596, n6936);
  and g11240 (n6937, n_4595, n_4596);
  not g11241 (n_4597, n6937);
  and g11242 (n6938, \asqrt[47] , n_4597);
  and g11246 (n6942, n_4323, n_4322);
  and g11247 (n6943, \asqrt[31] , n6942);
  not g11248 (n_4598, n6943);
  and g11249 (n6944, n_4321, n_4598);
  not g11250 (n_4599, n6941);
  not g11251 (n_4600, n6944);
  and g11252 (n6945, n_4599, n_4600);
  and g11253 (n6946, n_1514, n_4595);
  and g11254 (n6947, n_4596, n6946);
  not g11255 (n_4601, n6945);
  not g11256 (n_4602, n6947);
  and g11257 (n6948, n_4601, n_4602);
  not g11258 (n_4603, n6938);
  not g11259 (n_4604, n6948);
  and g11260 (n6949, n_4603, n_4604);
  not g11261 (n_4605, n6949);
  and g11262 (n6950, \asqrt[48] , n_4605);
  and g11266 (n6954, n_4331, n_4330);
  and g11267 (n6955, \asqrt[31] , n6954);
  not g11268 (n_4606, n6955);
  and g11269 (n6956, n_4329, n_4606);
  not g11270 (n_4607, n6953);
  not g11271 (n_4608, n6956);
  and g11272 (n6957, n_4607, n_4608);
  and g11273 (n6958, n_1362, n_4603);
  and g11274 (n6959, n_4604, n6958);
  not g11275 (n_4609, n6957);
  not g11276 (n_4610, n6959);
  and g11277 (n6960, n_4609, n_4610);
  not g11278 (n_4611, n6950);
  not g11279 (n_4612, n6960);
  and g11280 (n6961, n_4611, n_4612);
  not g11281 (n_4613, n6961);
  and g11282 (n6962, \asqrt[49] , n_4613);
  and g11286 (n6966, n_4339, n_4338);
  and g11287 (n6967, \asqrt[31] , n6966);
  not g11288 (n_4614, n6967);
  and g11289 (n6968, n_4337, n_4614);
  not g11290 (n_4615, n6965);
  not g11291 (n_4616, n6968);
  and g11292 (n6969, n_4615, n_4616);
  and g11293 (n6970, n_1218, n_4611);
  and g11294 (n6971, n_4612, n6970);
  not g11295 (n_4617, n6969);
  not g11296 (n_4618, n6971);
  and g11297 (n6972, n_4617, n_4618);
  not g11298 (n_4619, n6962);
  not g11299 (n_4620, n6972);
  and g11300 (n6973, n_4619, n_4620);
  not g11301 (n_4621, n6973);
  and g11302 (n6974, \asqrt[50] , n_4621);
  and g11306 (n6978, n_4347, n_4346);
  and g11307 (n6979, \asqrt[31] , n6978);
  not g11308 (n_4622, n6979);
  and g11309 (n6980, n_4345, n_4622);
  not g11310 (n_4623, n6977);
  not g11311 (n_4624, n6980);
  and g11312 (n6981, n_4623, n_4624);
  and g11313 (n6982, n_1082, n_4619);
  and g11314 (n6983, n_4620, n6982);
  not g11315 (n_4625, n6981);
  not g11316 (n_4626, n6983);
  and g11317 (n6984, n_4625, n_4626);
  not g11318 (n_4627, n6974);
  not g11319 (n_4628, n6984);
  and g11320 (n6985, n_4627, n_4628);
  not g11321 (n_4629, n6985);
  and g11322 (n6986, \asqrt[51] , n_4629);
  and g11326 (n6990, n_4355, n_4354);
  and g11327 (n6991, \asqrt[31] , n6990);
  not g11328 (n_4630, n6991);
  and g11329 (n6992, n_4353, n_4630);
  not g11330 (n_4631, n6989);
  not g11331 (n_4632, n6992);
  and g11332 (n6993, n_4631, n_4632);
  and g11333 (n6994, n_954, n_4627);
  and g11334 (n6995, n_4628, n6994);
  not g11335 (n_4633, n6993);
  not g11336 (n_4634, n6995);
  and g11337 (n6996, n_4633, n_4634);
  not g11338 (n_4635, n6986);
  not g11339 (n_4636, n6996);
  and g11340 (n6997, n_4635, n_4636);
  not g11341 (n_4637, n6997);
  and g11342 (n6998, \asqrt[52] , n_4637);
  and g11346 (n7002, n_4363, n_4362);
  and g11347 (n7003, \asqrt[31] , n7002);
  not g11348 (n_4638, n7003);
  and g11349 (n7004, n_4361, n_4638);
  not g11350 (n_4639, n7001);
  not g11351 (n_4640, n7004);
  and g11352 (n7005, n_4639, n_4640);
  and g11353 (n7006, n_834, n_4635);
  and g11354 (n7007, n_4636, n7006);
  not g11355 (n_4641, n7005);
  not g11356 (n_4642, n7007);
  and g11357 (n7008, n_4641, n_4642);
  not g11358 (n_4643, n6998);
  not g11359 (n_4644, n7008);
  and g11360 (n7009, n_4643, n_4644);
  not g11361 (n_4645, n7009);
  and g11362 (n7010, \asqrt[53] , n_4645);
  and g11366 (n7014, n_4371, n_4370);
  and g11367 (n7015, \asqrt[31] , n7014);
  not g11368 (n_4646, n7015);
  and g11369 (n7016, n_4369, n_4646);
  not g11370 (n_4647, n7013);
  not g11371 (n_4648, n7016);
  and g11372 (n7017, n_4647, n_4648);
  and g11373 (n7018, n_722, n_4643);
  and g11374 (n7019, n_4644, n7018);
  not g11375 (n_4649, n7017);
  not g11376 (n_4650, n7019);
  and g11377 (n7020, n_4649, n_4650);
  not g11378 (n_4651, n7010);
  not g11379 (n_4652, n7020);
  and g11380 (n7021, n_4651, n_4652);
  not g11381 (n_4653, n7021);
  and g11382 (n7022, \asqrt[54] , n_4653);
  and g11386 (n7026, n_4379, n_4378);
  and g11387 (n7027, \asqrt[31] , n7026);
  not g11388 (n_4654, n7027);
  and g11389 (n7028, n_4377, n_4654);
  not g11390 (n_4655, n7025);
  not g11391 (n_4656, n7028);
  and g11392 (n7029, n_4655, n_4656);
  and g11393 (n7030, n_618, n_4651);
  and g11394 (n7031, n_4652, n7030);
  not g11395 (n_4657, n7029);
  not g11396 (n_4658, n7031);
  and g11397 (n7032, n_4657, n_4658);
  not g11398 (n_4659, n7022);
  not g11399 (n_4660, n7032);
  and g11400 (n7033, n_4659, n_4660);
  not g11401 (n_4661, n7033);
  and g11402 (n7034, \asqrt[55] , n_4661);
  and g11406 (n7038, n_4387, n_4386);
  and g11407 (n7039, \asqrt[31] , n7038);
  not g11408 (n_4662, n7039);
  and g11409 (n7040, n_4385, n_4662);
  not g11410 (n_4663, n7037);
  not g11411 (n_4664, n7040);
  and g11412 (n7041, n_4663, n_4664);
  and g11413 (n7042, n_522, n_4659);
  and g11414 (n7043, n_4660, n7042);
  not g11415 (n_4665, n7041);
  not g11416 (n_4666, n7043);
  and g11417 (n7044, n_4665, n_4666);
  not g11418 (n_4667, n7034);
  not g11419 (n_4668, n7044);
  and g11420 (n7045, n_4667, n_4668);
  not g11421 (n_4669, n7045);
  and g11422 (n7046, \asqrt[56] , n_4669);
  and g11426 (n7050, n_4395, n_4394);
  and g11427 (n7051, \asqrt[31] , n7050);
  not g11428 (n_4670, n7051);
  and g11429 (n7052, n_4393, n_4670);
  not g11430 (n_4671, n7049);
  not g11431 (n_4672, n7052);
  and g11432 (n7053, n_4671, n_4672);
  and g11433 (n7054, n_434, n_4667);
  and g11434 (n7055, n_4668, n7054);
  not g11435 (n_4673, n7053);
  not g11436 (n_4674, n7055);
  and g11437 (n7056, n_4673, n_4674);
  not g11438 (n_4675, n7046);
  not g11439 (n_4676, n7056);
  and g11440 (n7057, n_4675, n_4676);
  not g11441 (n_4677, n7057);
  and g11442 (n7058, \asqrt[57] , n_4677);
  and g11446 (n7062, n_4403, n_4402);
  and g11447 (n7063, \asqrt[31] , n7062);
  not g11448 (n_4678, n7063);
  and g11449 (n7064, n_4401, n_4678);
  not g11450 (n_4679, n7061);
  not g11451 (n_4680, n7064);
  and g11452 (n7065, n_4679, n_4680);
  and g11453 (n7066, n_354, n_4675);
  and g11454 (n7067, n_4676, n7066);
  not g11455 (n_4681, n7065);
  not g11456 (n_4682, n7067);
  and g11457 (n7068, n_4681, n_4682);
  not g11458 (n_4683, n7058);
  not g11459 (n_4684, n7068);
  and g11460 (n7069, n_4683, n_4684);
  not g11461 (n_4685, n7069);
  and g11462 (n7070, \asqrt[58] , n_4685);
  and g11466 (n7074, n_4411, n_4410);
  and g11467 (n7075, \asqrt[31] , n7074);
  not g11468 (n_4686, n7075);
  and g11469 (n7076, n_4409, n_4686);
  not g11470 (n_4687, n7073);
  not g11471 (n_4688, n7076);
  and g11472 (n7077, n_4687, n_4688);
  and g11473 (n7078, n_282, n_4683);
  and g11474 (n7079, n_4684, n7078);
  not g11475 (n_4689, n7077);
  not g11476 (n_4690, n7079);
  and g11477 (n7080, n_4689, n_4690);
  not g11478 (n_4691, n7070);
  not g11479 (n_4692, n7080);
  and g11480 (n7081, n_4691, n_4692);
  not g11481 (n_4693, n7081);
  and g11482 (n7082, \asqrt[59] , n_4693);
  and g11486 (n7086, n_4419, n_4418);
  and g11487 (n7087, \asqrt[31] , n7086);
  not g11488 (n_4694, n7087);
  and g11489 (n7088, n_4417, n_4694);
  not g11490 (n_4695, n7085);
  not g11491 (n_4696, n7088);
  and g11492 (n7089, n_4695, n_4696);
  and g11493 (n7090, n_218, n_4691);
  and g11494 (n7091, n_4692, n7090);
  not g11495 (n_4697, n7089);
  not g11496 (n_4698, n7091);
  and g11497 (n7092, n_4697, n_4698);
  not g11498 (n_4699, n7082);
  not g11499 (n_4700, n7092);
  and g11500 (n7093, n_4699, n_4700);
  not g11501 (n_4701, n7093);
  and g11502 (n7094, \asqrt[60] , n_4701);
  and g11506 (n7098, n_4427, n_4426);
  and g11507 (n7099, \asqrt[31] , n7098);
  not g11508 (n_4702, n7099);
  and g11509 (n7100, n_4425, n_4702);
  not g11510 (n_4703, n7097);
  not g11511 (n_4704, n7100);
  and g11512 (n7101, n_4703, n_4704);
  and g11513 (n7102, n_162, n_4699);
  and g11514 (n7103, n_4700, n7102);
  not g11515 (n_4705, n7101);
  not g11516 (n_4706, n7103);
  and g11517 (n7104, n_4705, n_4706);
  not g11518 (n_4707, n7094);
  not g11519 (n_4708, n7104);
  and g11520 (n7105, n_4707, n_4708);
  not g11521 (n_4709, n7105);
  and g11522 (n7106, \asqrt[61] , n_4709);
  and g11526 (n7110, n_4435, n_4434);
  and g11527 (n7111, \asqrt[31] , n7110);
  not g11528 (n_4710, n7111);
  and g11529 (n7112, n_4433, n_4710);
  not g11530 (n_4711, n7109);
  not g11531 (n_4712, n7112);
  and g11532 (n7113, n_4711, n_4712);
  and g11533 (n7114, n_115, n_4707);
  and g11534 (n7115, n_4708, n7114);
  not g11535 (n_4713, n7113);
  not g11536 (n_4714, n7115);
  and g11537 (n7116, n_4713, n_4714);
  not g11538 (n_4715, n7106);
  not g11539 (n_4716, n7116);
  and g11540 (n7117, n_4715, n_4716);
  not g11541 (n_4717, n7117);
  and g11542 (n7118, \asqrt[62] , n_4717);
  and g11546 (n7122, n_4443, n_4442);
  and g11547 (n7123, \asqrt[31] , n7122);
  not g11548 (n_4718, n7123);
  and g11549 (n7124, n_4441, n_4718);
  not g11550 (n_4719, n7121);
  not g11551 (n_4720, n7124);
  and g11552 (n7125, n_4719, n_4720);
  and g11553 (n7126, n_76, n_4715);
  and g11554 (n7127, n_4716, n7126);
  not g11555 (n_4721, n7125);
  not g11556 (n_4722, n7127);
  and g11557 (n7128, n_4721, n_4722);
  not g11558 (n_4723, n7118);
  not g11559 (n_4724, n7128);
  and g11560 (n7129, n_4723, n_4724);
  and g11564 (n7133, n_4451, n_4450);
  and g11565 (n7134, \asqrt[31] , n7133);
  not g11566 (n_4725, n7134);
  and g11567 (n7135, n_4449, n_4725);
  not g11568 (n_4726, n7132);
  not g11569 (n_4727, n7135);
  and g11570 (n7136, n_4726, n_4727);
  and g11571 (n7137, n_4458, n_4457);
  and g11572 (n7138, \asqrt[31] , n7137);
  not g11575 (n_4729, n7136);
  not g11577 (n_4730, n7129);
  not g11579 (n_4731, n7141);
  and g11580 (n7142, n_21, n_4731);
  and g11581 (n7143, n_4723, n7136);
  and g11582 (n7144, n_4724, n7143);
  and g11583 (n7145, n_4457, \asqrt[31] );
  not g11584 (n_4732, n7145);
  and g11585 (n7146, n6724, n_4732);
  not g11586 (n_4733, n7137);
  and g11587 (n7147, \asqrt[63] , n_4733);
  not g11588 (n_4734, n7146);
  and g11589 (n7148, n_4734, n7147);
  not g11595 (n_4735, n7148);
  not g11596 (n_4736, n7153);
  not g11598 (n_4737, n7144);
  and g11602 (n7157, \a[60] , \asqrt[30] );
  not g11603 (n_4742, \a[58] );
  not g11604 (n_4743, \a[59] );
  and g11605 (n7158, n_4742, n_4743);
  and g11606 (n7159, n_4470, n7158);
  not g11607 (n_4744, n7157);
  not g11608 (n_4745, n7159);
  and g11609 (n7160, n_4744, n_4745);
  not g11610 (n_4746, n7160);
  and g11611 (n7161, \asqrt[31] , n_4746);
  and g11617 (n7167, n_4470, \asqrt[30] );
  not g11618 (n_4747, n7167);
  and g11619 (n7168, \a[61] , n_4747);
  and g11620 (n7169, n6753, \asqrt[30] );
  not g11621 (n_4748, n7168);
  not g11622 (n_4749, n7169);
  and g11623 (n7170, n_4748, n_4749);
  not g11624 (n_4750, n7166);
  and g11625 (n7171, n_4750, n7170);
  not g11626 (n_4751, n7161);
  not g11627 (n_4752, n7171);
  and g11628 (n7172, n_4751, n_4752);
  not g11629 (n_4753, n7172);
  and g11630 (n7173, \asqrt[32] , n_4753);
  not g11631 (n_4754, \asqrt[32] );
  and g11632 (n7174, n_4754, n_4751);
  and g11633 (n7175, n_4752, n7174);
  not g11637 (n_4755, n7142);
  not g11639 (n_4756, n7179);
  and g11640 (n7180, n_4749, n_4756);
  not g11641 (n_4757, n7180);
  and g11642 (n7181, \a[62] , n_4757);
  and g11643 (n7182, n_4206, n_4756);
  and g11644 (n7183, n_4749, n7182);
  not g11645 (n_4758, n7181);
  not g11646 (n_4759, n7183);
  and g11647 (n7184, n_4758, n_4759);
  not g11648 (n_4760, n7175);
  not g11649 (n_4761, n7184);
  and g11650 (n7185, n_4760, n_4761);
  not g11651 (n_4762, n7173);
  not g11652 (n_4763, n7185);
  and g11653 (n7186, n_4762, n_4763);
  not g11654 (n_4764, n7186);
  and g11655 (n7187, \asqrt[33] , n_4764);
  and g11656 (n7188, n_4479, n_4478);
  not g11657 (n_4765, n6765);
  and g11658 (n7189, n_4765, n7188);
  and g11659 (n7190, \asqrt[30] , n7189);
  and g11660 (n7191, \asqrt[30] , n7188);
  not g11661 (n_4766, n7191);
  and g11662 (n7192, n6765, n_4766);
  not g11663 (n_4767, n7190);
  not g11664 (n_4768, n7192);
  and g11665 (n7193, n_4767, n_4768);
  and g11666 (n7194, n_4482, n_4762);
  and g11667 (n7195, n_4763, n7194);
  not g11668 (n_4769, n7193);
  not g11669 (n_4770, n7195);
  and g11670 (n7196, n_4769, n_4770);
  not g11671 (n_4771, n7187);
  not g11672 (n_4772, n7196);
  and g11673 (n7197, n_4771, n_4772);
  not g11674 (n_4773, n7197);
  and g11675 (n7198, \asqrt[34] , n_4773);
  and g11679 (n7202, n_4490, n_4488);
  and g11680 (n7203, \asqrt[30] , n7202);
  not g11681 (n_4774, n7203);
  and g11682 (n7204, n_4489, n_4774);
  not g11683 (n_4775, n7201);
  not g11684 (n_4776, n7204);
  and g11685 (n7205, n_4775, n_4776);
  and g11686 (n7206, n_4218, n_4771);
  and g11687 (n7207, n_4772, n7206);
  not g11688 (n_4777, n7205);
  not g11689 (n_4778, n7207);
  and g11690 (n7208, n_4777, n_4778);
  not g11691 (n_4779, n7198);
  not g11692 (n_4780, n7208);
  and g11693 (n7209, n_4779, n_4780);
  not g11694 (n_4781, n7209);
  and g11695 (n7210, \asqrt[35] , n_4781);
  and g11696 (n7211, n_3962, n_4779);
  and g11697 (n7212, n_4780, n7211);
  and g11701 (n7216, n_4499, n_4497);
  and g11702 (n7217, \asqrt[30] , n7216);
  not g11703 (n_4782, n7217);
  and g11704 (n7218, n_4498, n_4782);
  not g11705 (n_4783, n7215);
  not g11706 (n_4784, n7218);
  and g11707 (n7219, n_4783, n_4784);
  not g11708 (n_4785, n7212);
  not g11709 (n_4786, n7219);
  and g11710 (n7220, n_4785, n_4786);
  not g11711 (n_4787, n7210);
  not g11712 (n_4788, n7220);
  and g11713 (n7221, n_4787, n_4788);
  not g11714 (n_4789, n7221);
  and g11715 (n7222, \asqrt[36] , n_4789);
  and g11719 (n7226, n_4507, n_4506);
  and g11720 (n7227, \asqrt[30] , n7226);
  not g11721 (n_4790, n7227);
  and g11722 (n7228, n_4505, n_4790);
  not g11723 (n_4791, n7225);
  not g11724 (n_4792, n7228);
  and g11725 (n7229, n_4791, n_4792);
  and g11726 (n7230, n_3714, n_4787);
  and g11727 (n7231, n_4788, n7230);
  not g11728 (n_4793, n7229);
  not g11729 (n_4794, n7231);
  and g11730 (n7232, n_4793, n_4794);
  not g11731 (n_4795, n7222);
  not g11732 (n_4796, n7232);
  and g11733 (n7233, n_4795, n_4796);
  not g11734 (n_4797, n7233);
  and g11735 (n7234, \asqrt[37] , n_4797);
  and g11739 (n7238, n_4515, n_4514);
  and g11740 (n7239, \asqrt[30] , n7238);
  not g11741 (n_4798, n7239);
  and g11742 (n7240, n_4513, n_4798);
  not g11743 (n_4799, n7237);
  not g11744 (n_4800, n7240);
  and g11745 (n7241, n_4799, n_4800);
  and g11746 (n7242, n_3474, n_4795);
  and g11747 (n7243, n_4796, n7242);
  not g11748 (n_4801, n7241);
  not g11749 (n_4802, n7243);
  and g11750 (n7244, n_4801, n_4802);
  not g11751 (n_4803, n7234);
  not g11752 (n_4804, n7244);
  and g11753 (n7245, n_4803, n_4804);
  not g11754 (n_4805, n7245);
  and g11755 (n7246, \asqrt[38] , n_4805);
  and g11759 (n7250, n_4523, n_4522);
  and g11760 (n7251, \asqrt[30] , n7250);
  not g11761 (n_4806, n7251);
  and g11762 (n7252, n_4521, n_4806);
  not g11763 (n_4807, n7249);
  not g11764 (n_4808, n7252);
  and g11765 (n7253, n_4807, n_4808);
  and g11766 (n7254, n_3242, n_4803);
  and g11767 (n7255, n_4804, n7254);
  not g11768 (n_4809, n7253);
  not g11769 (n_4810, n7255);
  and g11770 (n7256, n_4809, n_4810);
  not g11771 (n_4811, n7246);
  not g11772 (n_4812, n7256);
  and g11773 (n7257, n_4811, n_4812);
  not g11774 (n_4813, n7257);
  and g11775 (n7258, \asqrt[39] , n_4813);
  and g11779 (n7262, n_4531, n_4530);
  and g11780 (n7263, \asqrt[30] , n7262);
  not g11781 (n_4814, n7263);
  and g11782 (n7264, n_4529, n_4814);
  not g11783 (n_4815, n7261);
  not g11784 (n_4816, n7264);
  and g11785 (n7265, n_4815, n_4816);
  and g11786 (n7266, n_3018, n_4811);
  and g11787 (n7267, n_4812, n7266);
  not g11788 (n_4817, n7265);
  not g11789 (n_4818, n7267);
  and g11790 (n7268, n_4817, n_4818);
  not g11791 (n_4819, n7258);
  not g11792 (n_4820, n7268);
  and g11793 (n7269, n_4819, n_4820);
  not g11794 (n_4821, n7269);
  and g11795 (n7270, \asqrt[40] , n_4821);
  and g11799 (n7274, n_4539, n_4538);
  and g11800 (n7275, \asqrt[30] , n7274);
  not g11801 (n_4822, n7275);
  and g11802 (n7276, n_4537, n_4822);
  not g11803 (n_4823, n7273);
  not g11804 (n_4824, n7276);
  and g11805 (n7277, n_4823, n_4824);
  and g11806 (n7278, n_2802, n_4819);
  and g11807 (n7279, n_4820, n7278);
  not g11808 (n_4825, n7277);
  not g11809 (n_4826, n7279);
  and g11810 (n7280, n_4825, n_4826);
  not g11811 (n_4827, n7270);
  not g11812 (n_4828, n7280);
  and g11813 (n7281, n_4827, n_4828);
  not g11814 (n_4829, n7281);
  and g11815 (n7282, \asqrt[41] , n_4829);
  and g11819 (n7286, n_4547, n_4546);
  and g11820 (n7287, \asqrt[30] , n7286);
  not g11821 (n_4830, n7287);
  and g11822 (n7288, n_4545, n_4830);
  not g11823 (n_4831, n7285);
  not g11824 (n_4832, n7288);
  and g11825 (n7289, n_4831, n_4832);
  and g11826 (n7290, n_2594, n_4827);
  and g11827 (n7291, n_4828, n7290);
  not g11828 (n_4833, n7289);
  not g11829 (n_4834, n7291);
  and g11830 (n7292, n_4833, n_4834);
  not g11831 (n_4835, n7282);
  not g11832 (n_4836, n7292);
  and g11833 (n7293, n_4835, n_4836);
  not g11834 (n_4837, n7293);
  and g11835 (n7294, \asqrt[42] , n_4837);
  and g11839 (n7298, n_4555, n_4554);
  and g11840 (n7299, \asqrt[30] , n7298);
  not g11841 (n_4838, n7299);
  and g11842 (n7300, n_4553, n_4838);
  not g11843 (n_4839, n7297);
  not g11844 (n_4840, n7300);
  and g11845 (n7301, n_4839, n_4840);
  and g11846 (n7302, n_2394, n_4835);
  and g11847 (n7303, n_4836, n7302);
  not g11848 (n_4841, n7301);
  not g11849 (n_4842, n7303);
  and g11850 (n7304, n_4841, n_4842);
  not g11851 (n_4843, n7294);
  not g11852 (n_4844, n7304);
  and g11853 (n7305, n_4843, n_4844);
  not g11854 (n_4845, n7305);
  and g11855 (n7306, \asqrt[43] , n_4845);
  and g11859 (n7310, n_4563, n_4562);
  and g11860 (n7311, \asqrt[30] , n7310);
  not g11861 (n_4846, n7311);
  and g11862 (n7312, n_4561, n_4846);
  not g11863 (n_4847, n7309);
  not g11864 (n_4848, n7312);
  and g11865 (n7313, n_4847, n_4848);
  and g11866 (n7314, n_2202, n_4843);
  and g11867 (n7315, n_4844, n7314);
  not g11868 (n_4849, n7313);
  not g11869 (n_4850, n7315);
  and g11870 (n7316, n_4849, n_4850);
  not g11871 (n_4851, n7306);
  not g11872 (n_4852, n7316);
  and g11873 (n7317, n_4851, n_4852);
  not g11874 (n_4853, n7317);
  and g11875 (n7318, \asqrt[44] , n_4853);
  and g11879 (n7322, n_4571, n_4570);
  and g11880 (n7323, \asqrt[30] , n7322);
  not g11881 (n_4854, n7323);
  and g11882 (n7324, n_4569, n_4854);
  not g11883 (n_4855, n7321);
  not g11884 (n_4856, n7324);
  and g11885 (n7325, n_4855, n_4856);
  and g11886 (n7326, n_2018, n_4851);
  and g11887 (n7327, n_4852, n7326);
  not g11888 (n_4857, n7325);
  not g11889 (n_4858, n7327);
  and g11890 (n7328, n_4857, n_4858);
  not g11891 (n_4859, n7318);
  not g11892 (n_4860, n7328);
  and g11893 (n7329, n_4859, n_4860);
  not g11894 (n_4861, n7329);
  and g11895 (n7330, \asqrt[45] , n_4861);
  and g11899 (n7334, n_4579, n_4578);
  and g11900 (n7335, \asqrt[30] , n7334);
  not g11901 (n_4862, n7335);
  and g11902 (n7336, n_4577, n_4862);
  not g11903 (n_4863, n7333);
  not g11904 (n_4864, n7336);
  and g11905 (n7337, n_4863, n_4864);
  and g11906 (n7338, n_1842, n_4859);
  and g11907 (n7339, n_4860, n7338);
  not g11908 (n_4865, n7337);
  not g11909 (n_4866, n7339);
  and g11910 (n7340, n_4865, n_4866);
  not g11911 (n_4867, n7330);
  not g11912 (n_4868, n7340);
  and g11913 (n7341, n_4867, n_4868);
  not g11914 (n_4869, n7341);
  and g11915 (n7342, \asqrt[46] , n_4869);
  and g11919 (n7346, n_4587, n_4586);
  and g11920 (n7347, \asqrt[30] , n7346);
  not g11921 (n_4870, n7347);
  and g11922 (n7348, n_4585, n_4870);
  not g11923 (n_4871, n7345);
  not g11924 (n_4872, n7348);
  and g11925 (n7349, n_4871, n_4872);
  and g11926 (n7350, n_1674, n_4867);
  and g11927 (n7351, n_4868, n7350);
  not g11928 (n_4873, n7349);
  not g11929 (n_4874, n7351);
  and g11930 (n7352, n_4873, n_4874);
  not g11931 (n_4875, n7342);
  not g11932 (n_4876, n7352);
  and g11933 (n7353, n_4875, n_4876);
  not g11934 (n_4877, n7353);
  and g11935 (n7354, \asqrt[47] , n_4877);
  and g11939 (n7358, n_4595, n_4594);
  and g11940 (n7359, \asqrt[30] , n7358);
  not g11941 (n_4878, n7359);
  and g11942 (n7360, n_4593, n_4878);
  not g11943 (n_4879, n7357);
  not g11944 (n_4880, n7360);
  and g11945 (n7361, n_4879, n_4880);
  and g11946 (n7362, n_1514, n_4875);
  and g11947 (n7363, n_4876, n7362);
  not g11948 (n_4881, n7361);
  not g11949 (n_4882, n7363);
  and g11950 (n7364, n_4881, n_4882);
  not g11951 (n_4883, n7354);
  not g11952 (n_4884, n7364);
  and g11953 (n7365, n_4883, n_4884);
  not g11954 (n_4885, n7365);
  and g11955 (n7366, \asqrt[48] , n_4885);
  and g11959 (n7370, n_4603, n_4602);
  and g11960 (n7371, \asqrt[30] , n7370);
  not g11961 (n_4886, n7371);
  and g11962 (n7372, n_4601, n_4886);
  not g11963 (n_4887, n7369);
  not g11964 (n_4888, n7372);
  and g11965 (n7373, n_4887, n_4888);
  and g11966 (n7374, n_1362, n_4883);
  and g11967 (n7375, n_4884, n7374);
  not g11968 (n_4889, n7373);
  not g11969 (n_4890, n7375);
  and g11970 (n7376, n_4889, n_4890);
  not g11971 (n_4891, n7366);
  not g11972 (n_4892, n7376);
  and g11973 (n7377, n_4891, n_4892);
  not g11974 (n_4893, n7377);
  and g11975 (n7378, \asqrt[49] , n_4893);
  and g11979 (n7382, n_4611, n_4610);
  and g11980 (n7383, \asqrt[30] , n7382);
  not g11981 (n_4894, n7383);
  and g11982 (n7384, n_4609, n_4894);
  not g11983 (n_4895, n7381);
  not g11984 (n_4896, n7384);
  and g11985 (n7385, n_4895, n_4896);
  and g11986 (n7386, n_1218, n_4891);
  and g11987 (n7387, n_4892, n7386);
  not g11988 (n_4897, n7385);
  not g11989 (n_4898, n7387);
  and g11990 (n7388, n_4897, n_4898);
  not g11991 (n_4899, n7378);
  not g11992 (n_4900, n7388);
  and g11993 (n7389, n_4899, n_4900);
  not g11994 (n_4901, n7389);
  and g11995 (n7390, \asqrt[50] , n_4901);
  and g11999 (n7394, n_4619, n_4618);
  and g12000 (n7395, \asqrt[30] , n7394);
  not g12001 (n_4902, n7395);
  and g12002 (n7396, n_4617, n_4902);
  not g12003 (n_4903, n7393);
  not g12004 (n_4904, n7396);
  and g12005 (n7397, n_4903, n_4904);
  and g12006 (n7398, n_1082, n_4899);
  and g12007 (n7399, n_4900, n7398);
  not g12008 (n_4905, n7397);
  not g12009 (n_4906, n7399);
  and g12010 (n7400, n_4905, n_4906);
  not g12011 (n_4907, n7390);
  not g12012 (n_4908, n7400);
  and g12013 (n7401, n_4907, n_4908);
  not g12014 (n_4909, n7401);
  and g12015 (n7402, \asqrt[51] , n_4909);
  and g12019 (n7406, n_4627, n_4626);
  and g12020 (n7407, \asqrt[30] , n7406);
  not g12021 (n_4910, n7407);
  and g12022 (n7408, n_4625, n_4910);
  not g12023 (n_4911, n7405);
  not g12024 (n_4912, n7408);
  and g12025 (n7409, n_4911, n_4912);
  and g12026 (n7410, n_954, n_4907);
  and g12027 (n7411, n_4908, n7410);
  not g12028 (n_4913, n7409);
  not g12029 (n_4914, n7411);
  and g12030 (n7412, n_4913, n_4914);
  not g12031 (n_4915, n7402);
  not g12032 (n_4916, n7412);
  and g12033 (n7413, n_4915, n_4916);
  not g12034 (n_4917, n7413);
  and g12035 (n7414, \asqrt[52] , n_4917);
  and g12039 (n7418, n_4635, n_4634);
  and g12040 (n7419, \asqrt[30] , n7418);
  not g12041 (n_4918, n7419);
  and g12042 (n7420, n_4633, n_4918);
  not g12043 (n_4919, n7417);
  not g12044 (n_4920, n7420);
  and g12045 (n7421, n_4919, n_4920);
  and g12046 (n7422, n_834, n_4915);
  and g12047 (n7423, n_4916, n7422);
  not g12048 (n_4921, n7421);
  not g12049 (n_4922, n7423);
  and g12050 (n7424, n_4921, n_4922);
  not g12051 (n_4923, n7414);
  not g12052 (n_4924, n7424);
  and g12053 (n7425, n_4923, n_4924);
  not g12054 (n_4925, n7425);
  and g12055 (n7426, \asqrt[53] , n_4925);
  and g12059 (n7430, n_4643, n_4642);
  and g12060 (n7431, \asqrt[30] , n7430);
  not g12061 (n_4926, n7431);
  and g12062 (n7432, n_4641, n_4926);
  not g12063 (n_4927, n7429);
  not g12064 (n_4928, n7432);
  and g12065 (n7433, n_4927, n_4928);
  and g12066 (n7434, n_722, n_4923);
  and g12067 (n7435, n_4924, n7434);
  not g12068 (n_4929, n7433);
  not g12069 (n_4930, n7435);
  and g12070 (n7436, n_4929, n_4930);
  not g12071 (n_4931, n7426);
  not g12072 (n_4932, n7436);
  and g12073 (n7437, n_4931, n_4932);
  not g12074 (n_4933, n7437);
  and g12075 (n7438, \asqrt[54] , n_4933);
  and g12079 (n7442, n_4651, n_4650);
  and g12080 (n7443, \asqrt[30] , n7442);
  not g12081 (n_4934, n7443);
  and g12082 (n7444, n_4649, n_4934);
  not g12083 (n_4935, n7441);
  not g12084 (n_4936, n7444);
  and g12085 (n7445, n_4935, n_4936);
  and g12086 (n7446, n_618, n_4931);
  and g12087 (n7447, n_4932, n7446);
  not g12088 (n_4937, n7445);
  not g12089 (n_4938, n7447);
  and g12090 (n7448, n_4937, n_4938);
  not g12091 (n_4939, n7438);
  not g12092 (n_4940, n7448);
  and g12093 (n7449, n_4939, n_4940);
  not g12094 (n_4941, n7449);
  and g12095 (n7450, \asqrt[55] , n_4941);
  and g12099 (n7454, n_4659, n_4658);
  and g12100 (n7455, \asqrt[30] , n7454);
  not g12101 (n_4942, n7455);
  and g12102 (n7456, n_4657, n_4942);
  not g12103 (n_4943, n7453);
  not g12104 (n_4944, n7456);
  and g12105 (n7457, n_4943, n_4944);
  and g12106 (n7458, n_522, n_4939);
  and g12107 (n7459, n_4940, n7458);
  not g12108 (n_4945, n7457);
  not g12109 (n_4946, n7459);
  and g12110 (n7460, n_4945, n_4946);
  not g12111 (n_4947, n7450);
  not g12112 (n_4948, n7460);
  and g12113 (n7461, n_4947, n_4948);
  not g12114 (n_4949, n7461);
  and g12115 (n7462, \asqrt[56] , n_4949);
  and g12119 (n7466, n_4667, n_4666);
  and g12120 (n7467, \asqrt[30] , n7466);
  not g12121 (n_4950, n7467);
  and g12122 (n7468, n_4665, n_4950);
  not g12123 (n_4951, n7465);
  not g12124 (n_4952, n7468);
  and g12125 (n7469, n_4951, n_4952);
  and g12126 (n7470, n_434, n_4947);
  and g12127 (n7471, n_4948, n7470);
  not g12128 (n_4953, n7469);
  not g12129 (n_4954, n7471);
  and g12130 (n7472, n_4953, n_4954);
  not g12131 (n_4955, n7462);
  not g12132 (n_4956, n7472);
  and g12133 (n7473, n_4955, n_4956);
  not g12134 (n_4957, n7473);
  and g12135 (n7474, \asqrt[57] , n_4957);
  and g12139 (n7478, n_4675, n_4674);
  and g12140 (n7479, \asqrt[30] , n7478);
  not g12141 (n_4958, n7479);
  and g12142 (n7480, n_4673, n_4958);
  not g12143 (n_4959, n7477);
  not g12144 (n_4960, n7480);
  and g12145 (n7481, n_4959, n_4960);
  and g12146 (n7482, n_354, n_4955);
  and g12147 (n7483, n_4956, n7482);
  not g12148 (n_4961, n7481);
  not g12149 (n_4962, n7483);
  and g12150 (n7484, n_4961, n_4962);
  not g12151 (n_4963, n7474);
  not g12152 (n_4964, n7484);
  and g12153 (n7485, n_4963, n_4964);
  not g12154 (n_4965, n7485);
  and g12155 (n7486, \asqrt[58] , n_4965);
  and g12159 (n7490, n_4683, n_4682);
  and g12160 (n7491, \asqrt[30] , n7490);
  not g12161 (n_4966, n7491);
  and g12162 (n7492, n_4681, n_4966);
  not g12163 (n_4967, n7489);
  not g12164 (n_4968, n7492);
  and g12165 (n7493, n_4967, n_4968);
  and g12166 (n7494, n_282, n_4963);
  and g12167 (n7495, n_4964, n7494);
  not g12168 (n_4969, n7493);
  not g12169 (n_4970, n7495);
  and g12170 (n7496, n_4969, n_4970);
  not g12171 (n_4971, n7486);
  not g12172 (n_4972, n7496);
  and g12173 (n7497, n_4971, n_4972);
  not g12174 (n_4973, n7497);
  and g12175 (n7498, \asqrt[59] , n_4973);
  and g12179 (n7502, n_4691, n_4690);
  and g12180 (n7503, \asqrt[30] , n7502);
  not g12181 (n_4974, n7503);
  and g12182 (n7504, n_4689, n_4974);
  not g12183 (n_4975, n7501);
  not g12184 (n_4976, n7504);
  and g12185 (n7505, n_4975, n_4976);
  and g12186 (n7506, n_218, n_4971);
  and g12187 (n7507, n_4972, n7506);
  not g12188 (n_4977, n7505);
  not g12189 (n_4978, n7507);
  and g12190 (n7508, n_4977, n_4978);
  not g12191 (n_4979, n7498);
  not g12192 (n_4980, n7508);
  and g12193 (n7509, n_4979, n_4980);
  not g12194 (n_4981, n7509);
  and g12195 (n7510, \asqrt[60] , n_4981);
  and g12199 (n7514, n_4699, n_4698);
  and g12200 (n7515, \asqrt[30] , n7514);
  not g12201 (n_4982, n7515);
  and g12202 (n7516, n_4697, n_4982);
  not g12203 (n_4983, n7513);
  not g12204 (n_4984, n7516);
  and g12205 (n7517, n_4983, n_4984);
  and g12206 (n7518, n_162, n_4979);
  and g12207 (n7519, n_4980, n7518);
  not g12208 (n_4985, n7517);
  not g12209 (n_4986, n7519);
  and g12210 (n7520, n_4985, n_4986);
  not g12211 (n_4987, n7510);
  not g12212 (n_4988, n7520);
  and g12213 (n7521, n_4987, n_4988);
  not g12214 (n_4989, n7521);
  and g12215 (n7522, \asqrt[61] , n_4989);
  and g12219 (n7526, n_4707, n_4706);
  and g12220 (n7527, \asqrt[30] , n7526);
  not g12221 (n_4990, n7527);
  and g12222 (n7528, n_4705, n_4990);
  not g12223 (n_4991, n7525);
  not g12224 (n_4992, n7528);
  and g12225 (n7529, n_4991, n_4992);
  and g12226 (n7530, n_115, n_4987);
  and g12227 (n7531, n_4988, n7530);
  not g12228 (n_4993, n7529);
  not g12229 (n_4994, n7531);
  and g12230 (n7532, n_4993, n_4994);
  not g12231 (n_4995, n7522);
  not g12232 (n_4996, n7532);
  and g12233 (n7533, n_4995, n_4996);
  not g12234 (n_4997, n7533);
  and g12235 (n7534, \asqrt[62] , n_4997);
  and g12239 (n7538, n_4715, n_4714);
  and g12240 (n7539, \asqrt[30] , n7538);
  not g12241 (n_4998, n7539);
  and g12242 (n7540, n_4713, n_4998);
  not g12243 (n_4999, n7537);
  not g12244 (n_5000, n7540);
  and g12245 (n7541, n_4999, n_5000);
  and g12246 (n7542, n_76, n_4995);
  and g12247 (n7543, n_4996, n7542);
  not g12248 (n_5001, n7541);
  not g12249 (n_5002, n7543);
  and g12250 (n7544, n_5001, n_5002);
  not g12251 (n_5003, n7534);
  not g12252 (n_5004, n7544);
  and g12253 (n7545, n_5003, n_5004);
  and g12257 (n7549, n_4723, n_4722);
  and g12258 (n7550, \asqrt[30] , n7549);
  not g12259 (n_5005, n7550);
  and g12260 (n7551, n_4721, n_5005);
  not g12261 (n_5006, n7548);
  not g12262 (n_5007, n7551);
  and g12263 (n7552, n_5006, n_5007);
  and g12264 (n7553, n_4730, n_4729);
  and g12265 (n7554, \asqrt[30] , n7553);
  not g12268 (n_5009, n7552);
  not g12270 (n_5010, n7545);
  not g12272 (n_5011, n7557);
  and g12273 (n7558, n_21, n_5011);
  and g12274 (n7559, n_5003, n7552);
  and g12275 (n7560, n_5004, n7559);
  and g12276 (n7561, n_4729, \asqrt[30] );
  not g12277 (n_5012, n7561);
  and g12278 (n7562, n7129, n_5012);
  not g12279 (n_5013, n7553);
  and g12280 (n7563, \asqrt[63] , n_5013);
  not g12281 (n_5014, n7562);
  and g12282 (n7564, n_5014, n7563);
  not g12288 (n_5015, n7564);
  not g12289 (n_5016, n7569);
  not g12291 (n_5017, n7560);
  and g12295 (n7573, \a[58] , \asqrt[29] );
  not g12296 (n_5022, \a[56] );
  not g12297 (n_5023, \a[57] );
  and g12298 (n7574, n_5022, n_5023);
  and g12299 (n7575, n_4742, n7574);
  not g12300 (n_5024, n7573);
  not g12301 (n_5025, n7575);
  and g12302 (n7576, n_5024, n_5025);
  not g12303 (n_5026, n7576);
  and g12304 (n7577, \asqrt[30] , n_5026);
  and g12310 (n7583, n_4742, \asqrt[29] );
  not g12311 (n_5027, n7583);
  and g12312 (n7584, \a[59] , n_5027);
  and g12313 (n7585, n7158, \asqrt[29] );
  not g12314 (n_5028, n7584);
  not g12315 (n_5029, n7585);
  and g12316 (n7586, n_5028, n_5029);
  not g12317 (n_5030, n7582);
  and g12318 (n7587, n_5030, n7586);
  not g12319 (n_5031, n7577);
  not g12320 (n_5032, n7587);
  and g12321 (n7588, n_5031, n_5032);
  not g12322 (n_5033, n7588);
  and g12323 (n7589, \asqrt[31] , n_5033);
  not g12324 (n_5034, \asqrt[31] );
  and g12325 (n7590, n_5034, n_5031);
  and g12326 (n7591, n_5032, n7590);
  not g12330 (n_5035, n7558);
  not g12332 (n_5036, n7595);
  and g12333 (n7596, n_5029, n_5036);
  not g12334 (n_5037, n7596);
  and g12335 (n7597, \a[60] , n_5037);
  and g12336 (n7598, n_4470, n_5036);
  and g12337 (n7599, n_5029, n7598);
  not g12338 (n_5038, n7597);
  not g12339 (n_5039, n7599);
  and g12340 (n7600, n_5038, n_5039);
  not g12341 (n_5040, n7591);
  not g12342 (n_5041, n7600);
  and g12343 (n7601, n_5040, n_5041);
  not g12344 (n_5042, n7589);
  not g12345 (n_5043, n7601);
  and g12346 (n7602, n_5042, n_5043);
  not g12347 (n_5044, n7602);
  and g12348 (n7603, \asqrt[32] , n_5044);
  and g12349 (n7604, n_4751, n_4750);
  not g12350 (n_5045, n7170);
  and g12351 (n7605, n_5045, n7604);
  and g12352 (n7606, \asqrt[29] , n7605);
  and g12353 (n7607, \asqrt[29] , n7604);
  not g12354 (n_5046, n7607);
  and g12355 (n7608, n7170, n_5046);
  not g12356 (n_5047, n7606);
  not g12357 (n_5048, n7608);
  and g12358 (n7609, n_5047, n_5048);
  and g12359 (n7610, n_4754, n_5042);
  and g12360 (n7611, n_5043, n7610);
  not g12361 (n_5049, n7609);
  not g12362 (n_5050, n7611);
  and g12363 (n7612, n_5049, n_5050);
  not g12364 (n_5051, n7603);
  not g12365 (n_5052, n7612);
  and g12366 (n7613, n_5051, n_5052);
  not g12367 (n_5053, n7613);
  and g12368 (n7614, \asqrt[33] , n_5053);
  and g12372 (n7618, n_4762, n_4760);
  and g12373 (n7619, \asqrt[29] , n7618);
  not g12374 (n_5054, n7619);
  and g12375 (n7620, n_4761, n_5054);
  not g12376 (n_5055, n7617);
  not g12377 (n_5056, n7620);
  and g12378 (n7621, n_5055, n_5056);
  and g12379 (n7622, n_4482, n_5051);
  and g12380 (n7623, n_5052, n7622);
  not g12381 (n_5057, n7621);
  not g12382 (n_5058, n7623);
  and g12383 (n7624, n_5057, n_5058);
  not g12384 (n_5059, n7614);
  not g12385 (n_5060, n7624);
  and g12386 (n7625, n_5059, n_5060);
  not g12387 (n_5061, n7625);
  and g12388 (n7626, \asqrt[34] , n_5061);
  and g12392 (n7630, n_4771, n_4770);
  and g12393 (n7631, \asqrt[29] , n7630);
  not g12394 (n_5062, n7631);
  and g12395 (n7632, n_4769, n_5062);
  not g12396 (n_5063, n7629);
  not g12397 (n_5064, n7632);
  and g12398 (n7633, n_5063, n_5064);
  and g12399 (n7634, n_4218, n_5059);
  and g12400 (n7635, n_5060, n7634);
  not g12401 (n_5065, n7633);
  not g12402 (n_5066, n7635);
  and g12403 (n7636, n_5065, n_5066);
  not g12404 (n_5067, n7626);
  not g12405 (n_5068, n7636);
  and g12406 (n7637, n_5067, n_5068);
  not g12407 (n_5069, n7637);
  and g12408 (n7638, \asqrt[35] , n_5069);
  and g12412 (n7642, n_4779, n_4778);
  and g12413 (n7643, \asqrt[29] , n7642);
  not g12414 (n_5070, n7643);
  and g12415 (n7644, n_4777, n_5070);
  not g12416 (n_5071, n7641);
  not g12417 (n_5072, n7644);
  and g12418 (n7645, n_5071, n_5072);
  and g12419 (n7646, n_3962, n_5067);
  and g12420 (n7647, n_5068, n7646);
  not g12421 (n_5073, n7645);
  not g12422 (n_5074, n7647);
  and g12423 (n7648, n_5073, n_5074);
  not g12424 (n_5075, n7638);
  not g12425 (n_5076, n7648);
  and g12426 (n7649, n_5075, n_5076);
  not g12427 (n_5077, n7649);
  and g12428 (n7650, \asqrt[36] , n_5077);
  and g12429 (n7651, n_3714, n_5075);
  and g12430 (n7652, n_5076, n7651);
  and g12434 (n7656, n_4787, n_4785);
  and g12435 (n7657, \asqrt[29] , n7656);
  not g12436 (n_5078, n7657);
  and g12437 (n7658, n_4786, n_5078);
  not g12438 (n_5079, n7655);
  not g12439 (n_5080, n7658);
  and g12440 (n7659, n_5079, n_5080);
  not g12441 (n_5081, n7652);
  not g12442 (n_5082, n7659);
  and g12443 (n7660, n_5081, n_5082);
  not g12444 (n_5083, n7650);
  not g12445 (n_5084, n7660);
  and g12446 (n7661, n_5083, n_5084);
  not g12447 (n_5085, n7661);
  and g12448 (n7662, \asqrt[37] , n_5085);
  and g12452 (n7666, n_4795, n_4794);
  and g12453 (n7667, \asqrt[29] , n7666);
  not g12454 (n_5086, n7667);
  and g12455 (n7668, n_4793, n_5086);
  not g12456 (n_5087, n7665);
  not g12457 (n_5088, n7668);
  and g12458 (n7669, n_5087, n_5088);
  and g12459 (n7670, n_3474, n_5083);
  and g12460 (n7671, n_5084, n7670);
  not g12461 (n_5089, n7669);
  not g12462 (n_5090, n7671);
  and g12463 (n7672, n_5089, n_5090);
  not g12464 (n_5091, n7662);
  not g12465 (n_5092, n7672);
  and g12466 (n7673, n_5091, n_5092);
  not g12467 (n_5093, n7673);
  and g12468 (n7674, \asqrt[38] , n_5093);
  and g12472 (n7678, n_4803, n_4802);
  and g12473 (n7679, \asqrt[29] , n7678);
  not g12474 (n_5094, n7679);
  and g12475 (n7680, n_4801, n_5094);
  not g12476 (n_5095, n7677);
  not g12477 (n_5096, n7680);
  and g12478 (n7681, n_5095, n_5096);
  and g12479 (n7682, n_3242, n_5091);
  and g12480 (n7683, n_5092, n7682);
  not g12481 (n_5097, n7681);
  not g12482 (n_5098, n7683);
  and g12483 (n7684, n_5097, n_5098);
  not g12484 (n_5099, n7674);
  not g12485 (n_5100, n7684);
  and g12486 (n7685, n_5099, n_5100);
  not g12487 (n_5101, n7685);
  and g12488 (n7686, \asqrt[39] , n_5101);
  and g12492 (n7690, n_4811, n_4810);
  and g12493 (n7691, \asqrt[29] , n7690);
  not g12494 (n_5102, n7691);
  and g12495 (n7692, n_4809, n_5102);
  not g12496 (n_5103, n7689);
  not g12497 (n_5104, n7692);
  and g12498 (n7693, n_5103, n_5104);
  and g12499 (n7694, n_3018, n_5099);
  and g12500 (n7695, n_5100, n7694);
  not g12501 (n_5105, n7693);
  not g12502 (n_5106, n7695);
  and g12503 (n7696, n_5105, n_5106);
  not g12504 (n_5107, n7686);
  not g12505 (n_5108, n7696);
  and g12506 (n7697, n_5107, n_5108);
  not g12507 (n_5109, n7697);
  and g12508 (n7698, \asqrt[40] , n_5109);
  and g12512 (n7702, n_4819, n_4818);
  and g12513 (n7703, \asqrt[29] , n7702);
  not g12514 (n_5110, n7703);
  and g12515 (n7704, n_4817, n_5110);
  not g12516 (n_5111, n7701);
  not g12517 (n_5112, n7704);
  and g12518 (n7705, n_5111, n_5112);
  and g12519 (n7706, n_2802, n_5107);
  and g12520 (n7707, n_5108, n7706);
  not g12521 (n_5113, n7705);
  not g12522 (n_5114, n7707);
  and g12523 (n7708, n_5113, n_5114);
  not g12524 (n_5115, n7698);
  not g12525 (n_5116, n7708);
  and g12526 (n7709, n_5115, n_5116);
  not g12527 (n_5117, n7709);
  and g12528 (n7710, \asqrt[41] , n_5117);
  and g12532 (n7714, n_4827, n_4826);
  and g12533 (n7715, \asqrt[29] , n7714);
  not g12534 (n_5118, n7715);
  and g12535 (n7716, n_4825, n_5118);
  not g12536 (n_5119, n7713);
  not g12537 (n_5120, n7716);
  and g12538 (n7717, n_5119, n_5120);
  and g12539 (n7718, n_2594, n_5115);
  and g12540 (n7719, n_5116, n7718);
  not g12541 (n_5121, n7717);
  not g12542 (n_5122, n7719);
  and g12543 (n7720, n_5121, n_5122);
  not g12544 (n_5123, n7710);
  not g12545 (n_5124, n7720);
  and g12546 (n7721, n_5123, n_5124);
  not g12547 (n_5125, n7721);
  and g12548 (n7722, \asqrt[42] , n_5125);
  and g12552 (n7726, n_4835, n_4834);
  and g12553 (n7727, \asqrt[29] , n7726);
  not g12554 (n_5126, n7727);
  and g12555 (n7728, n_4833, n_5126);
  not g12556 (n_5127, n7725);
  not g12557 (n_5128, n7728);
  and g12558 (n7729, n_5127, n_5128);
  and g12559 (n7730, n_2394, n_5123);
  and g12560 (n7731, n_5124, n7730);
  not g12561 (n_5129, n7729);
  not g12562 (n_5130, n7731);
  and g12563 (n7732, n_5129, n_5130);
  not g12564 (n_5131, n7722);
  not g12565 (n_5132, n7732);
  and g12566 (n7733, n_5131, n_5132);
  not g12567 (n_5133, n7733);
  and g12568 (n7734, \asqrt[43] , n_5133);
  and g12572 (n7738, n_4843, n_4842);
  and g12573 (n7739, \asqrt[29] , n7738);
  not g12574 (n_5134, n7739);
  and g12575 (n7740, n_4841, n_5134);
  not g12576 (n_5135, n7737);
  not g12577 (n_5136, n7740);
  and g12578 (n7741, n_5135, n_5136);
  and g12579 (n7742, n_2202, n_5131);
  and g12580 (n7743, n_5132, n7742);
  not g12581 (n_5137, n7741);
  not g12582 (n_5138, n7743);
  and g12583 (n7744, n_5137, n_5138);
  not g12584 (n_5139, n7734);
  not g12585 (n_5140, n7744);
  and g12586 (n7745, n_5139, n_5140);
  not g12587 (n_5141, n7745);
  and g12588 (n7746, \asqrt[44] , n_5141);
  and g12592 (n7750, n_4851, n_4850);
  and g12593 (n7751, \asqrt[29] , n7750);
  not g12594 (n_5142, n7751);
  and g12595 (n7752, n_4849, n_5142);
  not g12596 (n_5143, n7749);
  not g12597 (n_5144, n7752);
  and g12598 (n7753, n_5143, n_5144);
  and g12599 (n7754, n_2018, n_5139);
  and g12600 (n7755, n_5140, n7754);
  not g12601 (n_5145, n7753);
  not g12602 (n_5146, n7755);
  and g12603 (n7756, n_5145, n_5146);
  not g12604 (n_5147, n7746);
  not g12605 (n_5148, n7756);
  and g12606 (n7757, n_5147, n_5148);
  not g12607 (n_5149, n7757);
  and g12608 (n7758, \asqrt[45] , n_5149);
  and g12612 (n7762, n_4859, n_4858);
  and g12613 (n7763, \asqrt[29] , n7762);
  not g12614 (n_5150, n7763);
  and g12615 (n7764, n_4857, n_5150);
  not g12616 (n_5151, n7761);
  not g12617 (n_5152, n7764);
  and g12618 (n7765, n_5151, n_5152);
  and g12619 (n7766, n_1842, n_5147);
  and g12620 (n7767, n_5148, n7766);
  not g12621 (n_5153, n7765);
  not g12622 (n_5154, n7767);
  and g12623 (n7768, n_5153, n_5154);
  not g12624 (n_5155, n7758);
  not g12625 (n_5156, n7768);
  and g12626 (n7769, n_5155, n_5156);
  not g12627 (n_5157, n7769);
  and g12628 (n7770, \asqrt[46] , n_5157);
  and g12632 (n7774, n_4867, n_4866);
  and g12633 (n7775, \asqrt[29] , n7774);
  not g12634 (n_5158, n7775);
  and g12635 (n7776, n_4865, n_5158);
  not g12636 (n_5159, n7773);
  not g12637 (n_5160, n7776);
  and g12638 (n7777, n_5159, n_5160);
  and g12639 (n7778, n_1674, n_5155);
  and g12640 (n7779, n_5156, n7778);
  not g12641 (n_5161, n7777);
  not g12642 (n_5162, n7779);
  and g12643 (n7780, n_5161, n_5162);
  not g12644 (n_5163, n7770);
  not g12645 (n_5164, n7780);
  and g12646 (n7781, n_5163, n_5164);
  not g12647 (n_5165, n7781);
  and g12648 (n7782, \asqrt[47] , n_5165);
  and g12652 (n7786, n_4875, n_4874);
  and g12653 (n7787, \asqrt[29] , n7786);
  not g12654 (n_5166, n7787);
  and g12655 (n7788, n_4873, n_5166);
  not g12656 (n_5167, n7785);
  not g12657 (n_5168, n7788);
  and g12658 (n7789, n_5167, n_5168);
  and g12659 (n7790, n_1514, n_5163);
  and g12660 (n7791, n_5164, n7790);
  not g12661 (n_5169, n7789);
  not g12662 (n_5170, n7791);
  and g12663 (n7792, n_5169, n_5170);
  not g12664 (n_5171, n7782);
  not g12665 (n_5172, n7792);
  and g12666 (n7793, n_5171, n_5172);
  not g12667 (n_5173, n7793);
  and g12668 (n7794, \asqrt[48] , n_5173);
  and g12672 (n7798, n_4883, n_4882);
  and g12673 (n7799, \asqrt[29] , n7798);
  not g12674 (n_5174, n7799);
  and g12675 (n7800, n_4881, n_5174);
  not g12676 (n_5175, n7797);
  not g12677 (n_5176, n7800);
  and g12678 (n7801, n_5175, n_5176);
  and g12679 (n7802, n_1362, n_5171);
  and g12680 (n7803, n_5172, n7802);
  not g12681 (n_5177, n7801);
  not g12682 (n_5178, n7803);
  and g12683 (n7804, n_5177, n_5178);
  not g12684 (n_5179, n7794);
  not g12685 (n_5180, n7804);
  and g12686 (n7805, n_5179, n_5180);
  not g12687 (n_5181, n7805);
  and g12688 (n7806, \asqrt[49] , n_5181);
  and g12692 (n7810, n_4891, n_4890);
  and g12693 (n7811, \asqrt[29] , n7810);
  not g12694 (n_5182, n7811);
  and g12695 (n7812, n_4889, n_5182);
  not g12696 (n_5183, n7809);
  not g12697 (n_5184, n7812);
  and g12698 (n7813, n_5183, n_5184);
  and g12699 (n7814, n_1218, n_5179);
  and g12700 (n7815, n_5180, n7814);
  not g12701 (n_5185, n7813);
  not g12702 (n_5186, n7815);
  and g12703 (n7816, n_5185, n_5186);
  not g12704 (n_5187, n7806);
  not g12705 (n_5188, n7816);
  and g12706 (n7817, n_5187, n_5188);
  not g12707 (n_5189, n7817);
  and g12708 (n7818, \asqrt[50] , n_5189);
  and g12712 (n7822, n_4899, n_4898);
  and g12713 (n7823, \asqrt[29] , n7822);
  not g12714 (n_5190, n7823);
  and g12715 (n7824, n_4897, n_5190);
  not g12716 (n_5191, n7821);
  not g12717 (n_5192, n7824);
  and g12718 (n7825, n_5191, n_5192);
  and g12719 (n7826, n_1082, n_5187);
  and g12720 (n7827, n_5188, n7826);
  not g12721 (n_5193, n7825);
  not g12722 (n_5194, n7827);
  and g12723 (n7828, n_5193, n_5194);
  not g12724 (n_5195, n7818);
  not g12725 (n_5196, n7828);
  and g12726 (n7829, n_5195, n_5196);
  not g12727 (n_5197, n7829);
  and g12728 (n7830, \asqrt[51] , n_5197);
  and g12732 (n7834, n_4907, n_4906);
  and g12733 (n7835, \asqrt[29] , n7834);
  not g12734 (n_5198, n7835);
  and g12735 (n7836, n_4905, n_5198);
  not g12736 (n_5199, n7833);
  not g12737 (n_5200, n7836);
  and g12738 (n7837, n_5199, n_5200);
  and g12739 (n7838, n_954, n_5195);
  and g12740 (n7839, n_5196, n7838);
  not g12741 (n_5201, n7837);
  not g12742 (n_5202, n7839);
  and g12743 (n7840, n_5201, n_5202);
  not g12744 (n_5203, n7830);
  not g12745 (n_5204, n7840);
  and g12746 (n7841, n_5203, n_5204);
  not g12747 (n_5205, n7841);
  and g12748 (n7842, \asqrt[52] , n_5205);
  and g12752 (n7846, n_4915, n_4914);
  and g12753 (n7847, \asqrt[29] , n7846);
  not g12754 (n_5206, n7847);
  and g12755 (n7848, n_4913, n_5206);
  not g12756 (n_5207, n7845);
  not g12757 (n_5208, n7848);
  and g12758 (n7849, n_5207, n_5208);
  and g12759 (n7850, n_834, n_5203);
  and g12760 (n7851, n_5204, n7850);
  not g12761 (n_5209, n7849);
  not g12762 (n_5210, n7851);
  and g12763 (n7852, n_5209, n_5210);
  not g12764 (n_5211, n7842);
  not g12765 (n_5212, n7852);
  and g12766 (n7853, n_5211, n_5212);
  not g12767 (n_5213, n7853);
  and g12768 (n7854, \asqrt[53] , n_5213);
  and g12772 (n7858, n_4923, n_4922);
  and g12773 (n7859, \asqrt[29] , n7858);
  not g12774 (n_5214, n7859);
  and g12775 (n7860, n_4921, n_5214);
  not g12776 (n_5215, n7857);
  not g12777 (n_5216, n7860);
  and g12778 (n7861, n_5215, n_5216);
  and g12779 (n7862, n_722, n_5211);
  and g12780 (n7863, n_5212, n7862);
  not g12781 (n_5217, n7861);
  not g12782 (n_5218, n7863);
  and g12783 (n7864, n_5217, n_5218);
  not g12784 (n_5219, n7854);
  not g12785 (n_5220, n7864);
  and g12786 (n7865, n_5219, n_5220);
  not g12787 (n_5221, n7865);
  and g12788 (n7866, \asqrt[54] , n_5221);
  and g12792 (n7870, n_4931, n_4930);
  and g12793 (n7871, \asqrt[29] , n7870);
  not g12794 (n_5222, n7871);
  and g12795 (n7872, n_4929, n_5222);
  not g12796 (n_5223, n7869);
  not g12797 (n_5224, n7872);
  and g12798 (n7873, n_5223, n_5224);
  and g12799 (n7874, n_618, n_5219);
  and g12800 (n7875, n_5220, n7874);
  not g12801 (n_5225, n7873);
  not g12802 (n_5226, n7875);
  and g12803 (n7876, n_5225, n_5226);
  not g12804 (n_5227, n7866);
  not g12805 (n_5228, n7876);
  and g12806 (n7877, n_5227, n_5228);
  not g12807 (n_5229, n7877);
  and g12808 (n7878, \asqrt[55] , n_5229);
  and g12812 (n7882, n_4939, n_4938);
  and g12813 (n7883, \asqrt[29] , n7882);
  not g12814 (n_5230, n7883);
  and g12815 (n7884, n_4937, n_5230);
  not g12816 (n_5231, n7881);
  not g12817 (n_5232, n7884);
  and g12818 (n7885, n_5231, n_5232);
  and g12819 (n7886, n_522, n_5227);
  and g12820 (n7887, n_5228, n7886);
  not g12821 (n_5233, n7885);
  not g12822 (n_5234, n7887);
  and g12823 (n7888, n_5233, n_5234);
  not g12824 (n_5235, n7878);
  not g12825 (n_5236, n7888);
  and g12826 (n7889, n_5235, n_5236);
  not g12827 (n_5237, n7889);
  and g12828 (n7890, \asqrt[56] , n_5237);
  and g12832 (n7894, n_4947, n_4946);
  and g12833 (n7895, \asqrt[29] , n7894);
  not g12834 (n_5238, n7895);
  and g12835 (n7896, n_4945, n_5238);
  not g12836 (n_5239, n7893);
  not g12837 (n_5240, n7896);
  and g12838 (n7897, n_5239, n_5240);
  and g12839 (n7898, n_434, n_5235);
  and g12840 (n7899, n_5236, n7898);
  not g12841 (n_5241, n7897);
  not g12842 (n_5242, n7899);
  and g12843 (n7900, n_5241, n_5242);
  not g12844 (n_5243, n7890);
  not g12845 (n_5244, n7900);
  and g12846 (n7901, n_5243, n_5244);
  not g12847 (n_5245, n7901);
  and g12848 (n7902, \asqrt[57] , n_5245);
  and g12852 (n7906, n_4955, n_4954);
  and g12853 (n7907, \asqrt[29] , n7906);
  not g12854 (n_5246, n7907);
  and g12855 (n7908, n_4953, n_5246);
  not g12856 (n_5247, n7905);
  not g12857 (n_5248, n7908);
  and g12858 (n7909, n_5247, n_5248);
  and g12859 (n7910, n_354, n_5243);
  and g12860 (n7911, n_5244, n7910);
  not g12861 (n_5249, n7909);
  not g12862 (n_5250, n7911);
  and g12863 (n7912, n_5249, n_5250);
  not g12864 (n_5251, n7902);
  not g12865 (n_5252, n7912);
  and g12866 (n7913, n_5251, n_5252);
  not g12867 (n_5253, n7913);
  and g12868 (n7914, \asqrt[58] , n_5253);
  and g12872 (n7918, n_4963, n_4962);
  and g12873 (n7919, \asqrt[29] , n7918);
  not g12874 (n_5254, n7919);
  and g12875 (n7920, n_4961, n_5254);
  not g12876 (n_5255, n7917);
  not g12877 (n_5256, n7920);
  and g12878 (n7921, n_5255, n_5256);
  and g12879 (n7922, n_282, n_5251);
  and g12880 (n7923, n_5252, n7922);
  not g12881 (n_5257, n7921);
  not g12882 (n_5258, n7923);
  and g12883 (n7924, n_5257, n_5258);
  not g12884 (n_5259, n7914);
  not g12885 (n_5260, n7924);
  and g12886 (n7925, n_5259, n_5260);
  not g12887 (n_5261, n7925);
  and g12888 (n7926, \asqrt[59] , n_5261);
  and g12892 (n7930, n_4971, n_4970);
  and g12893 (n7931, \asqrt[29] , n7930);
  not g12894 (n_5262, n7931);
  and g12895 (n7932, n_4969, n_5262);
  not g12896 (n_5263, n7929);
  not g12897 (n_5264, n7932);
  and g12898 (n7933, n_5263, n_5264);
  and g12899 (n7934, n_218, n_5259);
  and g12900 (n7935, n_5260, n7934);
  not g12901 (n_5265, n7933);
  not g12902 (n_5266, n7935);
  and g12903 (n7936, n_5265, n_5266);
  not g12904 (n_5267, n7926);
  not g12905 (n_5268, n7936);
  and g12906 (n7937, n_5267, n_5268);
  not g12907 (n_5269, n7937);
  and g12908 (n7938, \asqrt[60] , n_5269);
  and g12912 (n7942, n_4979, n_4978);
  and g12913 (n7943, \asqrt[29] , n7942);
  not g12914 (n_5270, n7943);
  and g12915 (n7944, n_4977, n_5270);
  not g12916 (n_5271, n7941);
  not g12917 (n_5272, n7944);
  and g12918 (n7945, n_5271, n_5272);
  and g12919 (n7946, n_162, n_5267);
  and g12920 (n7947, n_5268, n7946);
  not g12921 (n_5273, n7945);
  not g12922 (n_5274, n7947);
  and g12923 (n7948, n_5273, n_5274);
  not g12924 (n_5275, n7938);
  not g12925 (n_5276, n7948);
  and g12926 (n7949, n_5275, n_5276);
  not g12927 (n_5277, n7949);
  and g12928 (n7950, \asqrt[61] , n_5277);
  and g12932 (n7954, n_4987, n_4986);
  and g12933 (n7955, \asqrt[29] , n7954);
  not g12934 (n_5278, n7955);
  and g12935 (n7956, n_4985, n_5278);
  not g12936 (n_5279, n7953);
  not g12937 (n_5280, n7956);
  and g12938 (n7957, n_5279, n_5280);
  and g12939 (n7958, n_115, n_5275);
  and g12940 (n7959, n_5276, n7958);
  not g12941 (n_5281, n7957);
  not g12942 (n_5282, n7959);
  and g12943 (n7960, n_5281, n_5282);
  not g12944 (n_5283, n7950);
  not g12945 (n_5284, n7960);
  and g12946 (n7961, n_5283, n_5284);
  not g12947 (n_5285, n7961);
  and g12948 (n7962, \asqrt[62] , n_5285);
  and g12952 (n7966, n_4995, n_4994);
  and g12953 (n7967, \asqrt[29] , n7966);
  not g12954 (n_5286, n7967);
  and g12955 (n7968, n_4993, n_5286);
  not g12956 (n_5287, n7965);
  not g12957 (n_5288, n7968);
  and g12958 (n7969, n_5287, n_5288);
  and g12959 (n7970, n_76, n_5283);
  and g12960 (n7971, n_5284, n7970);
  not g12961 (n_5289, n7969);
  not g12962 (n_5290, n7971);
  and g12963 (n7972, n_5289, n_5290);
  not g12964 (n_5291, n7962);
  not g12965 (n_5292, n7972);
  and g12966 (n7973, n_5291, n_5292);
  and g12970 (n7977, n_5003, n_5002);
  and g12971 (n7978, \asqrt[29] , n7977);
  not g12972 (n_5293, n7978);
  and g12973 (n7979, n_5001, n_5293);
  not g12974 (n_5294, n7976);
  not g12975 (n_5295, n7979);
  and g12976 (n7980, n_5294, n_5295);
  and g12977 (n7981, n_5010, n_5009);
  and g12978 (n7982, \asqrt[29] , n7981);
  not g12981 (n_5297, n7980);
  not g12983 (n_5298, n7973);
  not g12985 (n_5299, n7985);
  and g12986 (n7986, n_21, n_5299);
  and g12987 (n7987, n_5291, n7980);
  and g12988 (n7988, n_5292, n7987);
  and g12989 (n7989, n_5009, \asqrt[29] );
  not g12990 (n_5300, n7989);
  and g12991 (n7990, n7545, n_5300);
  not g12992 (n_5301, n7981);
  and g12993 (n7991, \asqrt[63] , n_5301);
  not g12994 (n_5302, n7990);
  and g12995 (n7992, n_5302, n7991);
  not g13001 (n_5303, n7992);
  not g13002 (n_5304, n7997);
  not g13004 (n_5305, n7988);
  and g13008 (n8001, \a[56] , \asqrt[28] );
  not g13009 (n_5310, \a[54] );
  not g13010 (n_5311, \a[55] );
  and g13011 (n8002, n_5310, n_5311);
  and g13012 (n8003, n_5022, n8002);
  not g13013 (n_5312, n8001);
  not g13014 (n_5313, n8003);
  and g13015 (n8004, n_5312, n_5313);
  not g13016 (n_5314, n8004);
  and g13017 (n8005, \asqrt[29] , n_5314);
  and g13023 (n8011, n_5022, \asqrt[28] );
  not g13024 (n_5315, n8011);
  and g13025 (n8012, \a[57] , n_5315);
  and g13026 (n8013, n7574, \asqrt[28] );
  not g13027 (n_5316, n8012);
  not g13028 (n_5317, n8013);
  and g13029 (n8014, n_5316, n_5317);
  not g13030 (n_5318, n8010);
  and g13031 (n8015, n_5318, n8014);
  not g13032 (n_5319, n8005);
  not g13033 (n_5320, n8015);
  and g13034 (n8016, n_5319, n_5320);
  not g13035 (n_5321, n8016);
  and g13036 (n8017, \asqrt[30] , n_5321);
  not g13037 (n_5322, \asqrt[30] );
  and g13038 (n8018, n_5322, n_5319);
  and g13039 (n8019, n_5320, n8018);
  not g13043 (n_5323, n7986);
  not g13045 (n_5324, n8023);
  and g13046 (n8024, n_5317, n_5324);
  not g13047 (n_5325, n8024);
  and g13048 (n8025, \a[58] , n_5325);
  and g13049 (n8026, n_4742, n_5324);
  and g13050 (n8027, n_5317, n8026);
  not g13051 (n_5326, n8025);
  not g13052 (n_5327, n8027);
  and g13053 (n8028, n_5326, n_5327);
  not g13054 (n_5328, n8019);
  not g13055 (n_5329, n8028);
  and g13056 (n8029, n_5328, n_5329);
  not g13057 (n_5330, n8017);
  not g13058 (n_5331, n8029);
  and g13059 (n8030, n_5330, n_5331);
  not g13060 (n_5332, n8030);
  and g13061 (n8031, \asqrt[31] , n_5332);
  and g13062 (n8032, n_5031, n_5030);
  not g13063 (n_5333, n7586);
  and g13064 (n8033, n_5333, n8032);
  and g13065 (n8034, \asqrt[28] , n8033);
  and g13066 (n8035, \asqrt[28] , n8032);
  not g13067 (n_5334, n8035);
  and g13068 (n8036, n7586, n_5334);
  not g13069 (n_5335, n8034);
  not g13070 (n_5336, n8036);
  and g13071 (n8037, n_5335, n_5336);
  and g13072 (n8038, n_5034, n_5330);
  and g13073 (n8039, n_5331, n8038);
  not g13074 (n_5337, n8037);
  not g13075 (n_5338, n8039);
  and g13076 (n8040, n_5337, n_5338);
  not g13077 (n_5339, n8031);
  not g13078 (n_5340, n8040);
  and g13079 (n8041, n_5339, n_5340);
  not g13080 (n_5341, n8041);
  and g13081 (n8042, \asqrt[32] , n_5341);
  and g13085 (n8046, n_5042, n_5040);
  and g13086 (n8047, \asqrt[28] , n8046);
  not g13087 (n_5342, n8047);
  and g13088 (n8048, n_5041, n_5342);
  not g13089 (n_5343, n8045);
  not g13090 (n_5344, n8048);
  and g13091 (n8049, n_5343, n_5344);
  and g13092 (n8050, n_4754, n_5339);
  and g13093 (n8051, n_5340, n8050);
  not g13094 (n_5345, n8049);
  not g13095 (n_5346, n8051);
  and g13096 (n8052, n_5345, n_5346);
  not g13097 (n_5347, n8042);
  not g13098 (n_5348, n8052);
  and g13099 (n8053, n_5347, n_5348);
  not g13100 (n_5349, n8053);
  and g13101 (n8054, \asqrt[33] , n_5349);
  and g13105 (n8058, n_5051, n_5050);
  and g13106 (n8059, \asqrt[28] , n8058);
  not g13107 (n_5350, n8059);
  and g13108 (n8060, n_5049, n_5350);
  not g13109 (n_5351, n8057);
  not g13110 (n_5352, n8060);
  and g13111 (n8061, n_5351, n_5352);
  and g13112 (n8062, n_4482, n_5347);
  and g13113 (n8063, n_5348, n8062);
  not g13114 (n_5353, n8061);
  not g13115 (n_5354, n8063);
  and g13116 (n8064, n_5353, n_5354);
  not g13117 (n_5355, n8054);
  not g13118 (n_5356, n8064);
  and g13119 (n8065, n_5355, n_5356);
  not g13120 (n_5357, n8065);
  and g13121 (n8066, \asqrt[34] , n_5357);
  and g13125 (n8070, n_5059, n_5058);
  and g13126 (n8071, \asqrt[28] , n8070);
  not g13127 (n_5358, n8071);
  and g13128 (n8072, n_5057, n_5358);
  not g13129 (n_5359, n8069);
  not g13130 (n_5360, n8072);
  and g13131 (n8073, n_5359, n_5360);
  and g13132 (n8074, n_4218, n_5355);
  and g13133 (n8075, n_5356, n8074);
  not g13134 (n_5361, n8073);
  not g13135 (n_5362, n8075);
  and g13136 (n8076, n_5361, n_5362);
  not g13137 (n_5363, n8066);
  not g13138 (n_5364, n8076);
  and g13139 (n8077, n_5363, n_5364);
  not g13140 (n_5365, n8077);
  and g13141 (n8078, \asqrt[35] , n_5365);
  and g13145 (n8082, n_5067, n_5066);
  and g13146 (n8083, \asqrt[28] , n8082);
  not g13147 (n_5366, n8083);
  and g13148 (n8084, n_5065, n_5366);
  not g13149 (n_5367, n8081);
  not g13150 (n_5368, n8084);
  and g13151 (n8085, n_5367, n_5368);
  and g13152 (n8086, n_3962, n_5363);
  and g13153 (n8087, n_5364, n8086);
  not g13154 (n_5369, n8085);
  not g13155 (n_5370, n8087);
  and g13156 (n8088, n_5369, n_5370);
  not g13157 (n_5371, n8078);
  not g13158 (n_5372, n8088);
  and g13159 (n8089, n_5371, n_5372);
  not g13160 (n_5373, n8089);
  and g13161 (n8090, \asqrt[36] , n_5373);
  and g13165 (n8094, n_5075, n_5074);
  and g13166 (n8095, \asqrt[28] , n8094);
  not g13167 (n_5374, n8095);
  and g13168 (n8096, n_5073, n_5374);
  not g13169 (n_5375, n8093);
  not g13170 (n_5376, n8096);
  and g13171 (n8097, n_5375, n_5376);
  and g13172 (n8098, n_3714, n_5371);
  and g13173 (n8099, n_5372, n8098);
  not g13174 (n_5377, n8097);
  not g13175 (n_5378, n8099);
  and g13176 (n8100, n_5377, n_5378);
  not g13177 (n_5379, n8090);
  not g13178 (n_5380, n8100);
  and g13179 (n8101, n_5379, n_5380);
  not g13180 (n_5381, n8101);
  and g13181 (n8102, \asqrt[37] , n_5381);
  and g13182 (n8103, n_3474, n_5379);
  and g13183 (n8104, n_5380, n8103);
  and g13187 (n8108, n_5083, n_5081);
  and g13188 (n8109, \asqrt[28] , n8108);
  not g13189 (n_5382, n8109);
  and g13190 (n8110, n_5082, n_5382);
  not g13191 (n_5383, n8107);
  not g13192 (n_5384, n8110);
  and g13193 (n8111, n_5383, n_5384);
  not g13194 (n_5385, n8104);
  not g13195 (n_5386, n8111);
  and g13196 (n8112, n_5385, n_5386);
  not g13197 (n_5387, n8102);
  not g13198 (n_5388, n8112);
  and g13199 (n8113, n_5387, n_5388);
  not g13200 (n_5389, n8113);
  and g13201 (n8114, \asqrt[38] , n_5389);
  and g13205 (n8118, n_5091, n_5090);
  and g13206 (n8119, \asqrt[28] , n8118);
  not g13207 (n_5390, n8119);
  and g13208 (n8120, n_5089, n_5390);
  not g13209 (n_5391, n8117);
  not g13210 (n_5392, n8120);
  and g13211 (n8121, n_5391, n_5392);
  and g13212 (n8122, n_3242, n_5387);
  and g13213 (n8123, n_5388, n8122);
  not g13214 (n_5393, n8121);
  not g13215 (n_5394, n8123);
  and g13216 (n8124, n_5393, n_5394);
  not g13217 (n_5395, n8114);
  not g13218 (n_5396, n8124);
  and g13219 (n8125, n_5395, n_5396);
  not g13220 (n_5397, n8125);
  and g13221 (n8126, \asqrt[39] , n_5397);
  and g13225 (n8130, n_5099, n_5098);
  and g13226 (n8131, \asqrt[28] , n8130);
  not g13227 (n_5398, n8131);
  and g13228 (n8132, n_5097, n_5398);
  not g13229 (n_5399, n8129);
  not g13230 (n_5400, n8132);
  and g13231 (n8133, n_5399, n_5400);
  and g13232 (n8134, n_3018, n_5395);
  and g13233 (n8135, n_5396, n8134);
  not g13234 (n_5401, n8133);
  not g13235 (n_5402, n8135);
  and g13236 (n8136, n_5401, n_5402);
  not g13237 (n_5403, n8126);
  not g13238 (n_5404, n8136);
  and g13239 (n8137, n_5403, n_5404);
  not g13240 (n_5405, n8137);
  and g13241 (n8138, \asqrt[40] , n_5405);
  and g13245 (n8142, n_5107, n_5106);
  and g13246 (n8143, \asqrt[28] , n8142);
  not g13247 (n_5406, n8143);
  and g13248 (n8144, n_5105, n_5406);
  not g13249 (n_5407, n8141);
  not g13250 (n_5408, n8144);
  and g13251 (n8145, n_5407, n_5408);
  and g13252 (n8146, n_2802, n_5403);
  and g13253 (n8147, n_5404, n8146);
  not g13254 (n_5409, n8145);
  not g13255 (n_5410, n8147);
  and g13256 (n8148, n_5409, n_5410);
  not g13257 (n_5411, n8138);
  not g13258 (n_5412, n8148);
  and g13259 (n8149, n_5411, n_5412);
  not g13260 (n_5413, n8149);
  and g13261 (n8150, \asqrt[41] , n_5413);
  and g13265 (n8154, n_5115, n_5114);
  and g13266 (n8155, \asqrt[28] , n8154);
  not g13267 (n_5414, n8155);
  and g13268 (n8156, n_5113, n_5414);
  not g13269 (n_5415, n8153);
  not g13270 (n_5416, n8156);
  and g13271 (n8157, n_5415, n_5416);
  and g13272 (n8158, n_2594, n_5411);
  and g13273 (n8159, n_5412, n8158);
  not g13274 (n_5417, n8157);
  not g13275 (n_5418, n8159);
  and g13276 (n8160, n_5417, n_5418);
  not g13277 (n_5419, n8150);
  not g13278 (n_5420, n8160);
  and g13279 (n8161, n_5419, n_5420);
  not g13280 (n_5421, n8161);
  and g13281 (n8162, \asqrt[42] , n_5421);
  and g13285 (n8166, n_5123, n_5122);
  and g13286 (n8167, \asqrt[28] , n8166);
  not g13287 (n_5422, n8167);
  and g13288 (n8168, n_5121, n_5422);
  not g13289 (n_5423, n8165);
  not g13290 (n_5424, n8168);
  and g13291 (n8169, n_5423, n_5424);
  and g13292 (n8170, n_2394, n_5419);
  and g13293 (n8171, n_5420, n8170);
  not g13294 (n_5425, n8169);
  not g13295 (n_5426, n8171);
  and g13296 (n8172, n_5425, n_5426);
  not g13297 (n_5427, n8162);
  not g13298 (n_5428, n8172);
  and g13299 (n8173, n_5427, n_5428);
  not g13300 (n_5429, n8173);
  and g13301 (n8174, \asqrt[43] , n_5429);
  and g13305 (n8178, n_5131, n_5130);
  and g13306 (n8179, \asqrt[28] , n8178);
  not g13307 (n_5430, n8179);
  and g13308 (n8180, n_5129, n_5430);
  not g13309 (n_5431, n8177);
  not g13310 (n_5432, n8180);
  and g13311 (n8181, n_5431, n_5432);
  and g13312 (n8182, n_2202, n_5427);
  and g13313 (n8183, n_5428, n8182);
  not g13314 (n_5433, n8181);
  not g13315 (n_5434, n8183);
  and g13316 (n8184, n_5433, n_5434);
  not g13317 (n_5435, n8174);
  not g13318 (n_5436, n8184);
  and g13319 (n8185, n_5435, n_5436);
  not g13320 (n_5437, n8185);
  and g13321 (n8186, \asqrt[44] , n_5437);
  and g13325 (n8190, n_5139, n_5138);
  and g13326 (n8191, \asqrt[28] , n8190);
  not g13327 (n_5438, n8191);
  and g13328 (n8192, n_5137, n_5438);
  not g13329 (n_5439, n8189);
  not g13330 (n_5440, n8192);
  and g13331 (n8193, n_5439, n_5440);
  and g13332 (n8194, n_2018, n_5435);
  and g13333 (n8195, n_5436, n8194);
  not g13334 (n_5441, n8193);
  not g13335 (n_5442, n8195);
  and g13336 (n8196, n_5441, n_5442);
  not g13337 (n_5443, n8186);
  not g13338 (n_5444, n8196);
  and g13339 (n8197, n_5443, n_5444);
  not g13340 (n_5445, n8197);
  and g13341 (n8198, \asqrt[45] , n_5445);
  and g13345 (n8202, n_5147, n_5146);
  and g13346 (n8203, \asqrt[28] , n8202);
  not g13347 (n_5446, n8203);
  and g13348 (n8204, n_5145, n_5446);
  not g13349 (n_5447, n8201);
  not g13350 (n_5448, n8204);
  and g13351 (n8205, n_5447, n_5448);
  and g13352 (n8206, n_1842, n_5443);
  and g13353 (n8207, n_5444, n8206);
  not g13354 (n_5449, n8205);
  not g13355 (n_5450, n8207);
  and g13356 (n8208, n_5449, n_5450);
  not g13357 (n_5451, n8198);
  not g13358 (n_5452, n8208);
  and g13359 (n8209, n_5451, n_5452);
  not g13360 (n_5453, n8209);
  and g13361 (n8210, \asqrt[46] , n_5453);
  and g13365 (n8214, n_5155, n_5154);
  and g13366 (n8215, \asqrt[28] , n8214);
  not g13367 (n_5454, n8215);
  and g13368 (n8216, n_5153, n_5454);
  not g13369 (n_5455, n8213);
  not g13370 (n_5456, n8216);
  and g13371 (n8217, n_5455, n_5456);
  and g13372 (n8218, n_1674, n_5451);
  and g13373 (n8219, n_5452, n8218);
  not g13374 (n_5457, n8217);
  not g13375 (n_5458, n8219);
  and g13376 (n8220, n_5457, n_5458);
  not g13377 (n_5459, n8210);
  not g13378 (n_5460, n8220);
  and g13379 (n8221, n_5459, n_5460);
  not g13380 (n_5461, n8221);
  and g13381 (n8222, \asqrt[47] , n_5461);
  and g13385 (n8226, n_5163, n_5162);
  and g13386 (n8227, \asqrt[28] , n8226);
  not g13387 (n_5462, n8227);
  and g13388 (n8228, n_5161, n_5462);
  not g13389 (n_5463, n8225);
  not g13390 (n_5464, n8228);
  and g13391 (n8229, n_5463, n_5464);
  and g13392 (n8230, n_1514, n_5459);
  and g13393 (n8231, n_5460, n8230);
  not g13394 (n_5465, n8229);
  not g13395 (n_5466, n8231);
  and g13396 (n8232, n_5465, n_5466);
  not g13397 (n_5467, n8222);
  not g13398 (n_5468, n8232);
  and g13399 (n8233, n_5467, n_5468);
  not g13400 (n_5469, n8233);
  and g13401 (n8234, \asqrt[48] , n_5469);
  and g13405 (n8238, n_5171, n_5170);
  and g13406 (n8239, \asqrt[28] , n8238);
  not g13407 (n_5470, n8239);
  and g13408 (n8240, n_5169, n_5470);
  not g13409 (n_5471, n8237);
  not g13410 (n_5472, n8240);
  and g13411 (n8241, n_5471, n_5472);
  and g13412 (n8242, n_1362, n_5467);
  and g13413 (n8243, n_5468, n8242);
  not g13414 (n_5473, n8241);
  not g13415 (n_5474, n8243);
  and g13416 (n8244, n_5473, n_5474);
  not g13417 (n_5475, n8234);
  not g13418 (n_5476, n8244);
  and g13419 (n8245, n_5475, n_5476);
  not g13420 (n_5477, n8245);
  and g13421 (n8246, \asqrt[49] , n_5477);
  and g13425 (n8250, n_5179, n_5178);
  and g13426 (n8251, \asqrt[28] , n8250);
  not g13427 (n_5478, n8251);
  and g13428 (n8252, n_5177, n_5478);
  not g13429 (n_5479, n8249);
  not g13430 (n_5480, n8252);
  and g13431 (n8253, n_5479, n_5480);
  and g13432 (n8254, n_1218, n_5475);
  and g13433 (n8255, n_5476, n8254);
  not g13434 (n_5481, n8253);
  not g13435 (n_5482, n8255);
  and g13436 (n8256, n_5481, n_5482);
  not g13437 (n_5483, n8246);
  not g13438 (n_5484, n8256);
  and g13439 (n8257, n_5483, n_5484);
  not g13440 (n_5485, n8257);
  and g13441 (n8258, \asqrt[50] , n_5485);
  and g13445 (n8262, n_5187, n_5186);
  and g13446 (n8263, \asqrt[28] , n8262);
  not g13447 (n_5486, n8263);
  and g13448 (n8264, n_5185, n_5486);
  not g13449 (n_5487, n8261);
  not g13450 (n_5488, n8264);
  and g13451 (n8265, n_5487, n_5488);
  and g13452 (n8266, n_1082, n_5483);
  and g13453 (n8267, n_5484, n8266);
  not g13454 (n_5489, n8265);
  not g13455 (n_5490, n8267);
  and g13456 (n8268, n_5489, n_5490);
  not g13457 (n_5491, n8258);
  not g13458 (n_5492, n8268);
  and g13459 (n8269, n_5491, n_5492);
  not g13460 (n_5493, n8269);
  and g13461 (n8270, \asqrt[51] , n_5493);
  and g13465 (n8274, n_5195, n_5194);
  and g13466 (n8275, \asqrt[28] , n8274);
  not g13467 (n_5494, n8275);
  and g13468 (n8276, n_5193, n_5494);
  not g13469 (n_5495, n8273);
  not g13470 (n_5496, n8276);
  and g13471 (n8277, n_5495, n_5496);
  and g13472 (n8278, n_954, n_5491);
  and g13473 (n8279, n_5492, n8278);
  not g13474 (n_5497, n8277);
  not g13475 (n_5498, n8279);
  and g13476 (n8280, n_5497, n_5498);
  not g13477 (n_5499, n8270);
  not g13478 (n_5500, n8280);
  and g13479 (n8281, n_5499, n_5500);
  not g13480 (n_5501, n8281);
  and g13481 (n8282, \asqrt[52] , n_5501);
  and g13485 (n8286, n_5203, n_5202);
  and g13486 (n8287, \asqrt[28] , n8286);
  not g13487 (n_5502, n8287);
  and g13488 (n8288, n_5201, n_5502);
  not g13489 (n_5503, n8285);
  not g13490 (n_5504, n8288);
  and g13491 (n8289, n_5503, n_5504);
  and g13492 (n8290, n_834, n_5499);
  and g13493 (n8291, n_5500, n8290);
  not g13494 (n_5505, n8289);
  not g13495 (n_5506, n8291);
  and g13496 (n8292, n_5505, n_5506);
  not g13497 (n_5507, n8282);
  not g13498 (n_5508, n8292);
  and g13499 (n8293, n_5507, n_5508);
  not g13500 (n_5509, n8293);
  and g13501 (n8294, \asqrt[53] , n_5509);
  and g13505 (n8298, n_5211, n_5210);
  and g13506 (n8299, \asqrt[28] , n8298);
  not g13507 (n_5510, n8299);
  and g13508 (n8300, n_5209, n_5510);
  not g13509 (n_5511, n8297);
  not g13510 (n_5512, n8300);
  and g13511 (n8301, n_5511, n_5512);
  and g13512 (n8302, n_722, n_5507);
  and g13513 (n8303, n_5508, n8302);
  not g13514 (n_5513, n8301);
  not g13515 (n_5514, n8303);
  and g13516 (n8304, n_5513, n_5514);
  not g13517 (n_5515, n8294);
  not g13518 (n_5516, n8304);
  and g13519 (n8305, n_5515, n_5516);
  not g13520 (n_5517, n8305);
  and g13521 (n8306, \asqrt[54] , n_5517);
  and g13525 (n8310, n_5219, n_5218);
  and g13526 (n8311, \asqrt[28] , n8310);
  not g13527 (n_5518, n8311);
  and g13528 (n8312, n_5217, n_5518);
  not g13529 (n_5519, n8309);
  not g13530 (n_5520, n8312);
  and g13531 (n8313, n_5519, n_5520);
  and g13532 (n8314, n_618, n_5515);
  and g13533 (n8315, n_5516, n8314);
  not g13534 (n_5521, n8313);
  not g13535 (n_5522, n8315);
  and g13536 (n8316, n_5521, n_5522);
  not g13537 (n_5523, n8306);
  not g13538 (n_5524, n8316);
  and g13539 (n8317, n_5523, n_5524);
  not g13540 (n_5525, n8317);
  and g13541 (n8318, \asqrt[55] , n_5525);
  and g13545 (n8322, n_5227, n_5226);
  and g13546 (n8323, \asqrt[28] , n8322);
  not g13547 (n_5526, n8323);
  and g13548 (n8324, n_5225, n_5526);
  not g13549 (n_5527, n8321);
  not g13550 (n_5528, n8324);
  and g13551 (n8325, n_5527, n_5528);
  and g13552 (n8326, n_522, n_5523);
  and g13553 (n8327, n_5524, n8326);
  not g13554 (n_5529, n8325);
  not g13555 (n_5530, n8327);
  and g13556 (n8328, n_5529, n_5530);
  not g13557 (n_5531, n8318);
  not g13558 (n_5532, n8328);
  and g13559 (n8329, n_5531, n_5532);
  not g13560 (n_5533, n8329);
  and g13561 (n8330, \asqrt[56] , n_5533);
  and g13565 (n8334, n_5235, n_5234);
  and g13566 (n8335, \asqrt[28] , n8334);
  not g13567 (n_5534, n8335);
  and g13568 (n8336, n_5233, n_5534);
  not g13569 (n_5535, n8333);
  not g13570 (n_5536, n8336);
  and g13571 (n8337, n_5535, n_5536);
  and g13572 (n8338, n_434, n_5531);
  and g13573 (n8339, n_5532, n8338);
  not g13574 (n_5537, n8337);
  not g13575 (n_5538, n8339);
  and g13576 (n8340, n_5537, n_5538);
  not g13577 (n_5539, n8330);
  not g13578 (n_5540, n8340);
  and g13579 (n8341, n_5539, n_5540);
  not g13580 (n_5541, n8341);
  and g13581 (n8342, \asqrt[57] , n_5541);
  and g13585 (n8346, n_5243, n_5242);
  and g13586 (n8347, \asqrt[28] , n8346);
  not g13587 (n_5542, n8347);
  and g13588 (n8348, n_5241, n_5542);
  not g13589 (n_5543, n8345);
  not g13590 (n_5544, n8348);
  and g13591 (n8349, n_5543, n_5544);
  and g13592 (n8350, n_354, n_5539);
  and g13593 (n8351, n_5540, n8350);
  not g13594 (n_5545, n8349);
  not g13595 (n_5546, n8351);
  and g13596 (n8352, n_5545, n_5546);
  not g13597 (n_5547, n8342);
  not g13598 (n_5548, n8352);
  and g13599 (n8353, n_5547, n_5548);
  not g13600 (n_5549, n8353);
  and g13601 (n8354, \asqrt[58] , n_5549);
  and g13605 (n8358, n_5251, n_5250);
  and g13606 (n8359, \asqrt[28] , n8358);
  not g13607 (n_5550, n8359);
  and g13608 (n8360, n_5249, n_5550);
  not g13609 (n_5551, n8357);
  not g13610 (n_5552, n8360);
  and g13611 (n8361, n_5551, n_5552);
  and g13612 (n8362, n_282, n_5547);
  and g13613 (n8363, n_5548, n8362);
  not g13614 (n_5553, n8361);
  not g13615 (n_5554, n8363);
  and g13616 (n8364, n_5553, n_5554);
  not g13617 (n_5555, n8354);
  not g13618 (n_5556, n8364);
  and g13619 (n8365, n_5555, n_5556);
  not g13620 (n_5557, n8365);
  and g13621 (n8366, \asqrt[59] , n_5557);
  and g13625 (n8370, n_5259, n_5258);
  and g13626 (n8371, \asqrt[28] , n8370);
  not g13627 (n_5558, n8371);
  and g13628 (n8372, n_5257, n_5558);
  not g13629 (n_5559, n8369);
  not g13630 (n_5560, n8372);
  and g13631 (n8373, n_5559, n_5560);
  and g13632 (n8374, n_218, n_5555);
  and g13633 (n8375, n_5556, n8374);
  not g13634 (n_5561, n8373);
  not g13635 (n_5562, n8375);
  and g13636 (n8376, n_5561, n_5562);
  not g13637 (n_5563, n8366);
  not g13638 (n_5564, n8376);
  and g13639 (n8377, n_5563, n_5564);
  not g13640 (n_5565, n8377);
  and g13641 (n8378, \asqrt[60] , n_5565);
  and g13645 (n8382, n_5267, n_5266);
  and g13646 (n8383, \asqrt[28] , n8382);
  not g13647 (n_5566, n8383);
  and g13648 (n8384, n_5265, n_5566);
  not g13649 (n_5567, n8381);
  not g13650 (n_5568, n8384);
  and g13651 (n8385, n_5567, n_5568);
  and g13652 (n8386, n_162, n_5563);
  and g13653 (n8387, n_5564, n8386);
  not g13654 (n_5569, n8385);
  not g13655 (n_5570, n8387);
  and g13656 (n8388, n_5569, n_5570);
  not g13657 (n_5571, n8378);
  not g13658 (n_5572, n8388);
  and g13659 (n8389, n_5571, n_5572);
  not g13660 (n_5573, n8389);
  and g13661 (n8390, \asqrt[61] , n_5573);
  and g13665 (n8394, n_5275, n_5274);
  and g13666 (n8395, \asqrt[28] , n8394);
  not g13667 (n_5574, n8395);
  and g13668 (n8396, n_5273, n_5574);
  not g13669 (n_5575, n8393);
  not g13670 (n_5576, n8396);
  and g13671 (n8397, n_5575, n_5576);
  and g13672 (n8398, n_115, n_5571);
  and g13673 (n8399, n_5572, n8398);
  not g13674 (n_5577, n8397);
  not g13675 (n_5578, n8399);
  and g13676 (n8400, n_5577, n_5578);
  not g13677 (n_5579, n8390);
  not g13678 (n_5580, n8400);
  and g13679 (n8401, n_5579, n_5580);
  not g13680 (n_5581, n8401);
  and g13681 (n8402, \asqrt[62] , n_5581);
  and g13685 (n8406, n_5283, n_5282);
  and g13686 (n8407, \asqrt[28] , n8406);
  not g13687 (n_5582, n8407);
  and g13688 (n8408, n_5281, n_5582);
  not g13689 (n_5583, n8405);
  not g13690 (n_5584, n8408);
  and g13691 (n8409, n_5583, n_5584);
  and g13692 (n8410, n_76, n_5579);
  and g13693 (n8411, n_5580, n8410);
  not g13694 (n_5585, n8409);
  not g13695 (n_5586, n8411);
  and g13696 (n8412, n_5585, n_5586);
  not g13697 (n_5587, n8402);
  not g13698 (n_5588, n8412);
  and g13699 (n8413, n_5587, n_5588);
  and g13703 (n8417, n_5291, n_5290);
  and g13704 (n8418, \asqrt[28] , n8417);
  not g13705 (n_5589, n8418);
  and g13706 (n8419, n_5289, n_5589);
  not g13707 (n_5590, n8416);
  not g13708 (n_5591, n8419);
  and g13709 (n8420, n_5590, n_5591);
  and g13710 (n8421, n_5298, n_5297);
  and g13711 (n8422, \asqrt[28] , n8421);
  not g13714 (n_5593, n8420);
  not g13716 (n_5594, n8413);
  not g13718 (n_5595, n8425);
  and g13719 (n8426, n_21, n_5595);
  and g13720 (n8427, n_5587, n8420);
  and g13721 (n8428, n_5588, n8427);
  and g13722 (n8429, n_5297, \asqrt[28] );
  not g13723 (n_5596, n8429);
  and g13724 (n8430, n7973, n_5596);
  not g13725 (n_5597, n8421);
  and g13726 (n8431, \asqrt[63] , n_5597);
  not g13727 (n_5598, n8430);
  and g13728 (n8432, n_5598, n8431);
  not g13734 (n_5599, n8432);
  not g13735 (n_5600, n8437);
  not g13737 (n_5601, n8428);
  and g13741 (n8441, \a[54] , \asqrt[27] );
  not g13742 (n_5606, \a[52] );
  not g13743 (n_5607, \a[53] );
  and g13744 (n8442, n_5606, n_5607);
  and g13745 (n8443, n_5310, n8442);
  not g13746 (n_5608, n8441);
  not g13747 (n_5609, n8443);
  and g13748 (n8444, n_5608, n_5609);
  not g13749 (n_5610, n8444);
  and g13750 (n8445, \asqrt[28] , n_5610);
  and g13756 (n8451, n_5310, \asqrt[27] );
  not g13757 (n_5611, n8451);
  and g13758 (n8452, \a[55] , n_5611);
  and g13759 (n8453, n8002, \asqrt[27] );
  not g13760 (n_5612, n8452);
  not g13761 (n_5613, n8453);
  and g13762 (n8454, n_5612, n_5613);
  not g13763 (n_5614, n8450);
  and g13764 (n8455, n_5614, n8454);
  not g13765 (n_5615, n8445);
  not g13766 (n_5616, n8455);
  and g13767 (n8456, n_5615, n_5616);
  not g13768 (n_5617, n8456);
  and g13769 (n8457, \asqrt[29] , n_5617);
  not g13770 (n_5618, \asqrt[29] );
  and g13771 (n8458, n_5618, n_5615);
  and g13772 (n8459, n_5616, n8458);
  not g13776 (n_5619, n8426);
  not g13778 (n_5620, n8463);
  and g13779 (n8464, n_5613, n_5620);
  not g13780 (n_5621, n8464);
  and g13781 (n8465, \a[56] , n_5621);
  and g13782 (n8466, n_5022, n_5620);
  and g13783 (n8467, n_5613, n8466);
  not g13784 (n_5622, n8465);
  not g13785 (n_5623, n8467);
  and g13786 (n8468, n_5622, n_5623);
  not g13787 (n_5624, n8459);
  not g13788 (n_5625, n8468);
  and g13789 (n8469, n_5624, n_5625);
  not g13790 (n_5626, n8457);
  not g13791 (n_5627, n8469);
  and g13792 (n8470, n_5626, n_5627);
  not g13793 (n_5628, n8470);
  and g13794 (n8471, \asqrt[30] , n_5628);
  and g13795 (n8472, n_5319, n_5318);
  not g13796 (n_5629, n8014);
  and g13797 (n8473, n_5629, n8472);
  and g13798 (n8474, \asqrt[27] , n8473);
  and g13799 (n8475, \asqrt[27] , n8472);
  not g13800 (n_5630, n8475);
  and g13801 (n8476, n8014, n_5630);
  not g13802 (n_5631, n8474);
  not g13803 (n_5632, n8476);
  and g13804 (n8477, n_5631, n_5632);
  and g13805 (n8478, n_5322, n_5626);
  and g13806 (n8479, n_5627, n8478);
  not g13807 (n_5633, n8477);
  not g13808 (n_5634, n8479);
  and g13809 (n8480, n_5633, n_5634);
  not g13810 (n_5635, n8471);
  not g13811 (n_5636, n8480);
  and g13812 (n8481, n_5635, n_5636);
  not g13813 (n_5637, n8481);
  and g13814 (n8482, \asqrt[31] , n_5637);
  and g13818 (n8486, n_5330, n_5328);
  and g13819 (n8487, \asqrt[27] , n8486);
  not g13820 (n_5638, n8487);
  and g13821 (n8488, n_5329, n_5638);
  not g13822 (n_5639, n8485);
  not g13823 (n_5640, n8488);
  and g13824 (n8489, n_5639, n_5640);
  and g13825 (n8490, n_5034, n_5635);
  and g13826 (n8491, n_5636, n8490);
  not g13827 (n_5641, n8489);
  not g13828 (n_5642, n8491);
  and g13829 (n8492, n_5641, n_5642);
  not g13830 (n_5643, n8482);
  not g13831 (n_5644, n8492);
  and g13832 (n8493, n_5643, n_5644);
  not g13833 (n_5645, n8493);
  and g13834 (n8494, \asqrt[32] , n_5645);
  and g13838 (n8498, n_5339, n_5338);
  and g13839 (n8499, \asqrt[27] , n8498);
  not g13840 (n_5646, n8499);
  and g13841 (n8500, n_5337, n_5646);
  not g13842 (n_5647, n8497);
  not g13843 (n_5648, n8500);
  and g13844 (n8501, n_5647, n_5648);
  and g13845 (n8502, n_4754, n_5643);
  and g13846 (n8503, n_5644, n8502);
  not g13847 (n_5649, n8501);
  not g13848 (n_5650, n8503);
  and g13849 (n8504, n_5649, n_5650);
  not g13850 (n_5651, n8494);
  not g13851 (n_5652, n8504);
  and g13852 (n8505, n_5651, n_5652);
  not g13853 (n_5653, n8505);
  and g13854 (n8506, \asqrt[33] , n_5653);
  and g13858 (n8510, n_5347, n_5346);
  and g13859 (n8511, \asqrt[27] , n8510);
  not g13860 (n_5654, n8511);
  and g13861 (n8512, n_5345, n_5654);
  not g13862 (n_5655, n8509);
  not g13863 (n_5656, n8512);
  and g13864 (n8513, n_5655, n_5656);
  and g13865 (n8514, n_4482, n_5651);
  and g13866 (n8515, n_5652, n8514);
  not g13867 (n_5657, n8513);
  not g13868 (n_5658, n8515);
  and g13869 (n8516, n_5657, n_5658);
  not g13870 (n_5659, n8506);
  not g13871 (n_5660, n8516);
  and g13872 (n8517, n_5659, n_5660);
  not g13873 (n_5661, n8517);
  and g13874 (n8518, \asqrt[34] , n_5661);
  and g13878 (n8522, n_5355, n_5354);
  and g13879 (n8523, \asqrt[27] , n8522);
  not g13880 (n_5662, n8523);
  and g13881 (n8524, n_5353, n_5662);
  not g13882 (n_5663, n8521);
  not g13883 (n_5664, n8524);
  and g13884 (n8525, n_5663, n_5664);
  and g13885 (n8526, n_4218, n_5659);
  and g13886 (n8527, n_5660, n8526);
  not g13887 (n_5665, n8525);
  not g13888 (n_5666, n8527);
  and g13889 (n8528, n_5665, n_5666);
  not g13890 (n_5667, n8518);
  not g13891 (n_5668, n8528);
  and g13892 (n8529, n_5667, n_5668);
  not g13893 (n_5669, n8529);
  and g13894 (n8530, \asqrt[35] , n_5669);
  and g13898 (n8534, n_5363, n_5362);
  and g13899 (n8535, \asqrt[27] , n8534);
  not g13900 (n_5670, n8535);
  and g13901 (n8536, n_5361, n_5670);
  not g13902 (n_5671, n8533);
  not g13903 (n_5672, n8536);
  and g13904 (n8537, n_5671, n_5672);
  and g13905 (n8538, n_3962, n_5667);
  and g13906 (n8539, n_5668, n8538);
  not g13907 (n_5673, n8537);
  not g13908 (n_5674, n8539);
  and g13909 (n8540, n_5673, n_5674);
  not g13910 (n_5675, n8530);
  not g13911 (n_5676, n8540);
  and g13912 (n8541, n_5675, n_5676);
  not g13913 (n_5677, n8541);
  and g13914 (n8542, \asqrt[36] , n_5677);
  and g13918 (n8546, n_5371, n_5370);
  and g13919 (n8547, \asqrt[27] , n8546);
  not g13920 (n_5678, n8547);
  and g13921 (n8548, n_5369, n_5678);
  not g13922 (n_5679, n8545);
  not g13923 (n_5680, n8548);
  and g13924 (n8549, n_5679, n_5680);
  and g13925 (n8550, n_3714, n_5675);
  and g13926 (n8551, n_5676, n8550);
  not g13927 (n_5681, n8549);
  not g13928 (n_5682, n8551);
  and g13929 (n8552, n_5681, n_5682);
  not g13930 (n_5683, n8542);
  not g13931 (n_5684, n8552);
  and g13932 (n8553, n_5683, n_5684);
  not g13933 (n_5685, n8553);
  and g13934 (n8554, \asqrt[37] , n_5685);
  and g13938 (n8558, n_5379, n_5378);
  and g13939 (n8559, \asqrt[27] , n8558);
  not g13940 (n_5686, n8559);
  and g13941 (n8560, n_5377, n_5686);
  not g13942 (n_5687, n8557);
  not g13943 (n_5688, n8560);
  and g13944 (n8561, n_5687, n_5688);
  and g13945 (n8562, n_3474, n_5683);
  and g13946 (n8563, n_5684, n8562);
  not g13947 (n_5689, n8561);
  not g13948 (n_5690, n8563);
  and g13949 (n8564, n_5689, n_5690);
  not g13950 (n_5691, n8554);
  not g13951 (n_5692, n8564);
  and g13952 (n8565, n_5691, n_5692);
  not g13953 (n_5693, n8565);
  and g13954 (n8566, \asqrt[38] , n_5693);
  and g13955 (n8567, n_3242, n_5691);
  and g13956 (n8568, n_5692, n8567);
  and g13960 (n8572, n_5387, n_5385);
  and g13961 (n8573, \asqrt[27] , n8572);
  not g13962 (n_5694, n8573);
  and g13963 (n8574, n_5386, n_5694);
  not g13964 (n_5695, n8571);
  not g13965 (n_5696, n8574);
  and g13966 (n8575, n_5695, n_5696);
  not g13967 (n_5697, n8568);
  not g13968 (n_5698, n8575);
  and g13969 (n8576, n_5697, n_5698);
  not g13970 (n_5699, n8566);
  not g13971 (n_5700, n8576);
  and g13972 (n8577, n_5699, n_5700);
  not g13973 (n_5701, n8577);
  and g13974 (n8578, \asqrt[39] , n_5701);
  and g13978 (n8582, n_5395, n_5394);
  and g13979 (n8583, \asqrt[27] , n8582);
  not g13980 (n_5702, n8583);
  and g13981 (n8584, n_5393, n_5702);
  not g13982 (n_5703, n8581);
  not g13983 (n_5704, n8584);
  and g13984 (n8585, n_5703, n_5704);
  and g13985 (n8586, n_3018, n_5699);
  and g13986 (n8587, n_5700, n8586);
  not g13987 (n_5705, n8585);
  not g13988 (n_5706, n8587);
  and g13989 (n8588, n_5705, n_5706);
  not g13990 (n_5707, n8578);
  not g13991 (n_5708, n8588);
  and g13992 (n8589, n_5707, n_5708);
  not g13993 (n_5709, n8589);
  and g13994 (n8590, \asqrt[40] , n_5709);
  and g13998 (n8594, n_5403, n_5402);
  and g13999 (n8595, \asqrt[27] , n8594);
  not g14000 (n_5710, n8595);
  and g14001 (n8596, n_5401, n_5710);
  not g14002 (n_5711, n8593);
  not g14003 (n_5712, n8596);
  and g14004 (n8597, n_5711, n_5712);
  and g14005 (n8598, n_2802, n_5707);
  and g14006 (n8599, n_5708, n8598);
  not g14007 (n_5713, n8597);
  not g14008 (n_5714, n8599);
  and g14009 (n8600, n_5713, n_5714);
  not g14010 (n_5715, n8590);
  not g14011 (n_5716, n8600);
  and g14012 (n8601, n_5715, n_5716);
  not g14013 (n_5717, n8601);
  and g14014 (n8602, \asqrt[41] , n_5717);
  and g14018 (n8606, n_5411, n_5410);
  and g14019 (n8607, \asqrt[27] , n8606);
  not g14020 (n_5718, n8607);
  and g14021 (n8608, n_5409, n_5718);
  not g14022 (n_5719, n8605);
  not g14023 (n_5720, n8608);
  and g14024 (n8609, n_5719, n_5720);
  and g14025 (n8610, n_2594, n_5715);
  and g14026 (n8611, n_5716, n8610);
  not g14027 (n_5721, n8609);
  not g14028 (n_5722, n8611);
  and g14029 (n8612, n_5721, n_5722);
  not g14030 (n_5723, n8602);
  not g14031 (n_5724, n8612);
  and g14032 (n8613, n_5723, n_5724);
  not g14033 (n_5725, n8613);
  and g14034 (n8614, \asqrt[42] , n_5725);
  and g14038 (n8618, n_5419, n_5418);
  and g14039 (n8619, \asqrt[27] , n8618);
  not g14040 (n_5726, n8619);
  and g14041 (n8620, n_5417, n_5726);
  not g14042 (n_5727, n8617);
  not g14043 (n_5728, n8620);
  and g14044 (n8621, n_5727, n_5728);
  and g14045 (n8622, n_2394, n_5723);
  and g14046 (n8623, n_5724, n8622);
  not g14047 (n_5729, n8621);
  not g14048 (n_5730, n8623);
  and g14049 (n8624, n_5729, n_5730);
  not g14050 (n_5731, n8614);
  not g14051 (n_5732, n8624);
  and g14052 (n8625, n_5731, n_5732);
  not g14053 (n_5733, n8625);
  and g14054 (n8626, \asqrt[43] , n_5733);
  and g14058 (n8630, n_5427, n_5426);
  and g14059 (n8631, \asqrt[27] , n8630);
  not g14060 (n_5734, n8631);
  and g14061 (n8632, n_5425, n_5734);
  not g14062 (n_5735, n8629);
  not g14063 (n_5736, n8632);
  and g14064 (n8633, n_5735, n_5736);
  and g14065 (n8634, n_2202, n_5731);
  and g14066 (n8635, n_5732, n8634);
  not g14067 (n_5737, n8633);
  not g14068 (n_5738, n8635);
  and g14069 (n8636, n_5737, n_5738);
  not g14070 (n_5739, n8626);
  not g14071 (n_5740, n8636);
  and g14072 (n8637, n_5739, n_5740);
  not g14073 (n_5741, n8637);
  and g14074 (n8638, \asqrt[44] , n_5741);
  and g14078 (n8642, n_5435, n_5434);
  and g14079 (n8643, \asqrt[27] , n8642);
  not g14080 (n_5742, n8643);
  and g14081 (n8644, n_5433, n_5742);
  not g14082 (n_5743, n8641);
  not g14083 (n_5744, n8644);
  and g14084 (n8645, n_5743, n_5744);
  and g14085 (n8646, n_2018, n_5739);
  and g14086 (n8647, n_5740, n8646);
  not g14087 (n_5745, n8645);
  not g14088 (n_5746, n8647);
  and g14089 (n8648, n_5745, n_5746);
  not g14090 (n_5747, n8638);
  not g14091 (n_5748, n8648);
  and g14092 (n8649, n_5747, n_5748);
  not g14093 (n_5749, n8649);
  and g14094 (n8650, \asqrt[45] , n_5749);
  and g14098 (n8654, n_5443, n_5442);
  and g14099 (n8655, \asqrt[27] , n8654);
  not g14100 (n_5750, n8655);
  and g14101 (n8656, n_5441, n_5750);
  not g14102 (n_5751, n8653);
  not g14103 (n_5752, n8656);
  and g14104 (n8657, n_5751, n_5752);
  and g14105 (n8658, n_1842, n_5747);
  and g14106 (n8659, n_5748, n8658);
  not g14107 (n_5753, n8657);
  not g14108 (n_5754, n8659);
  and g14109 (n8660, n_5753, n_5754);
  not g14110 (n_5755, n8650);
  not g14111 (n_5756, n8660);
  and g14112 (n8661, n_5755, n_5756);
  not g14113 (n_5757, n8661);
  and g14114 (n8662, \asqrt[46] , n_5757);
  and g14118 (n8666, n_5451, n_5450);
  and g14119 (n8667, \asqrt[27] , n8666);
  not g14120 (n_5758, n8667);
  and g14121 (n8668, n_5449, n_5758);
  not g14122 (n_5759, n8665);
  not g14123 (n_5760, n8668);
  and g14124 (n8669, n_5759, n_5760);
  and g14125 (n8670, n_1674, n_5755);
  and g14126 (n8671, n_5756, n8670);
  not g14127 (n_5761, n8669);
  not g14128 (n_5762, n8671);
  and g14129 (n8672, n_5761, n_5762);
  not g14130 (n_5763, n8662);
  not g14131 (n_5764, n8672);
  and g14132 (n8673, n_5763, n_5764);
  not g14133 (n_5765, n8673);
  and g14134 (n8674, \asqrt[47] , n_5765);
  and g14138 (n8678, n_5459, n_5458);
  and g14139 (n8679, \asqrt[27] , n8678);
  not g14140 (n_5766, n8679);
  and g14141 (n8680, n_5457, n_5766);
  not g14142 (n_5767, n8677);
  not g14143 (n_5768, n8680);
  and g14144 (n8681, n_5767, n_5768);
  and g14145 (n8682, n_1514, n_5763);
  and g14146 (n8683, n_5764, n8682);
  not g14147 (n_5769, n8681);
  not g14148 (n_5770, n8683);
  and g14149 (n8684, n_5769, n_5770);
  not g14150 (n_5771, n8674);
  not g14151 (n_5772, n8684);
  and g14152 (n8685, n_5771, n_5772);
  not g14153 (n_5773, n8685);
  and g14154 (n8686, \asqrt[48] , n_5773);
  and g14158 (n8690, n_5467, n_5466);
  and g14159 (n8691, \asqrt[27] , n8690);
  not g14160 (n_5774, n8691);
  and g14161 (n8692, n_5465, n_5774);
  not g14162 (n_5775, n8689);
  not g14163 (n_5776, n8692);
  and g14164 (n8693, n_5775, n_5776);
  and g14165 (n8694, n_1362, n_5771);
  and g14166 (n8695, n_5772, n8694);
  not g14167 (n_5777, n8693);
  not g14168 (n_5778, n8695);
  and g14169 (n8696, n_5777, n_5778);
  not g14170 (n_5779, n8686);
  not g14171 (n_5780, n8696);
  and g14172 (n8697, n_5779, n_5780);
  not g14173 (n_5781, n8697);
  and g14174 (n8698, \asqrt[49] , n_5781);
  and g14178 (n8702, n_5475, n_5474);
  and g14179 (n8703, \asqrt[27] , n8702);
  not g14180 (n_5782, n8703);
  and g14181 (n8704, n_5473, n_5782);
  not g14182 (n_5783, n8701);
  not g14183 (n_5784, n8704);
  and g14184 (n8705, n_5783, n_5784);
  and g14185 (n8706, n_1218, n_5779);
  and g14186 (n8707, n_5780, n8706);
  not g14187 (n_5785, n8705);
  not g14188 (n_5786, n8707);
  and g14189 (n8708, n_5785, n_5786);
  not g14190 (n_5787, n8698);
  not g14191 (n_5788, n8708);
  and g14192 (n8709, n_5787, n_5788);
  not g14193 (n_5789, n8709);
  and g14194 (n8710, \asqrt[50] , n_5789);
  and g14198 (n8714, n_5483, n_5482);
  and g14199 (n8715, \asqrt[27] , n8714);
  not g14200 (n_5790, n8715);
  and g14201 (n8716, n_5481, n_5790);
  not g14202 (n_5791, n8713);
  not g14203 (n_5792, n8716);
  and g14204 (n8717, n_5791, n_5792);
  and g14205 (n8718, n_1082, n_5787);
  and g14206 (n8719, n_5788, n8718);
  not g14207 (n_5793, n8717);
  not g14208 (n_5794, n8719);
  and g14209 (n8720, n_5793, n_5794);
  not g14210 (n_5795, n8710);
  not g14211 (n_5796, n8720);
  and g14212 (n8721, n_5795, n_5796);
  not g14213 (n_5797, n8721);
  and g14214 (n8722, \asqrt[51] , n_5797);
  and g14218 (n8726, n_5491, n_5490);
  and g14219 (n8727, \asqrt[27] , n8726);
  not g14220 (n_5798, n8727);
  and g14221 (n8728, n_5489, n_5798);
  not g14222 (n_5799, n8725);
  not g14223 (n_5800, n8728);
  and g14224 (n8729, n_5799, n_5800);
  and g14225 (n8730, n_954, n_5795);
  and g14226 (n8731, n_5796, n8730);
  not g14227 (n_5801, n8729);
  not g14228 (n_5802, n8731);
  and g14229 (n8732, n_5801, n_5802);
  not g14230 (n_5803, n8722);
  not g14231 (n_5804, n8732);
  and g14232 (n8733, n_5803, n_5804);
  not g14233 (n_5805, n8733);
  and g14234 (n8734, \asqrt[52] , n_5805);
  and g14238 (n8738, n_5499, n_5498);
  and g14239 (n8739, \asqrt[27] , n8738);
  not g14240 (n_5806, n8739);
  and g14241 (n8740, n_5497, n_5806);
  not g14242 (n_5807, n8737);
  not g14243 (n_5808, n8740);
  and g14244 (n8741, n_5807, n_5808);
  and g14245 (n8742, n_834, n_5803);
  and g14246 (n8743, n_5804, n8742);
  not g14247 (n_5809, n8741);
  not g14248 (n_5810, n8743);
  and g14249 (n8744, n_5809, n_5810);
  not g14250 (n_5811, n8734);
  not g14251 (n_5812, n8744);
  and g14252 (n8745, n_5811, n_5812);
  not g14253 (n_5813, n8745);
  and g14254 (n8746, \asqrt[53] , n_5813);
  and g14258 (n8750, n_5507, n_5506);
  and g14259 (n8751, \asqrt[27] , n8750);
  not g14260 (n_5814, n8751);
  and g14261 (n8752, n_5505, n_5814);
  not g14262 (n_5815, n8749);
  not g14263 (n_5816, n8752);
  and g14264 (n8753, n_5815, n_5816);
  and g14265 (n8754, n_722, n_5811);
  and g14266 (n8755, n_5812, n8754);
  not g14267 (n_5817, n8753);
  not g14268 (n_5818, n8755);
  and g14269 (n8756, n_5817, n_5818);
  not g14270 (n_5819, n8746);
  not g14271 (n_5820, n8756);
  and g14272 (n8757, n_5819, n_5820);
  not g14273 (n_5821, n8757);
  and g14274 (n8758, \asqrt[54] , n_5821);
  and g14278 (n8762, n_5515, n_5514);
  and g14279 (n8763, \asqrt[27] , n8762);
  not g14280 (n_5822, n8763);
  and g14281 (n8764, n_5513, n_5822);
  not g14282 (n_5823, n8761);
  not g14283 (n_5824, n8764);
  and g14284 (n8765, n_5823, n_5824);
  and g14285 (n8766, n_618, n_5819);
  and g14286 (n8767, n_5820, n8766);
  not g14287 (n_5825, n8765);
  not g14288 (n_5826, n8767);
  and g14289 (n8768, n_5825, n_5826);
  not g14290 (n_5827, n8758);
  not g14291 (n_5828, n8768);
  and g14292 (n8769, n_5827, n_5828);
  not g14293 (n_5829, n8769);
  and g14294 (n8770, \asqrt[55] , n_5829);
  and g14298 (n8774, n_5523, n_5522);
  and g14299 (n8775, \asqrt[27] , n8774);
  not g14300 (n_5830, n8775);
  and g14301 (n8776, n_5521, n_5830);
  not g14302 (n_5831, n8773);
  not g14303 (n_5832, n8776);
  and g14304 (n8777, n_5831, n_5832);
  and g14305 (n8778, n_522, n_5827);
  and g14306 (n8779, n_5828, n8778);
  not g14307 (n_5833, n8777);
  not g14308 (n_5834, n8779);
  and g14309 (n8780, n_5833, n_5834);
  not g14310 (n_5835, n8770);
  not g14311 (n_5836, n8780);
  and g14312 (n8781, n_5835, n_5836);
  not g14313 (n_5837, n8781);
  and g14314 (n8782, \asqrt[56] , n_5837);
  and g14318 (n8786, n_5531, n_5530);
  and g14319 (n8787, \asqrt[27] , n8786);
  not g14320 (n_5838, n8787);
  and g14321 (n8788, n_5529, n_5838);
  not g14322 (n_5839, n8785);
  not g14323 (n_5840, n8788);
  and g14324 (n8789, n_5839, n_5840);
  and g14325 (n8790, n_434, n_5835);
  and g14326 (n8791, n_5836, n8790);
  not g14327 (n_5841, n8789);
  not g14328 (n_5842, n8791);
  and g14329 (n8792, n_5841, n_5842);
  not g14330 (n_5843, n8782);
  not g14331 (n_5844, n8792);
  and g14332 (n8793, n_5843, n_5844);
  not g14333 (n_5845, n8793);
  and g14334 (n8794, \asqrt[57] , n_5845);
  and g14338 (n8798, n_5539, n_5538);
  and g14339 (n8799, \asqrt[27] , n8798);
  not g14340 (n_5846, n8799);
  and g14341 (n8800, n_5537, n_5846);
  not g14342 (n_5847, n8797);
  not g14343 (n_5848, n8800);
  and g14344 (n8801, n_5847, n_5848);
  and g14345 (n8802, n_354, n_5843);
  and g14346 (n8803, n_5844, n8802);
  not g14347 (n_5849, n8801);
  not g14348 (n_5850, n8803);
  and g14349 (n8804, n_5849, n_5850);
  not g14350 (n_5851, n8794);
  not g14351 (n_5852, n8804);
  and g14352 (n8805, n_5851, n_5852);
  not g14353 (n_5853, n8805);
  and g14354 (n8806, \asqrt[58] , n_5853);
  and g14358 (n8810, n_5547, n_5546);
  and g14359 (n8811, \asqrt[27] , n8810);
  not g14360 (n_5854, n8811);
  and g14361 (n8812, n_5545, n_5854);
  not g14362 (n_5855, n8809);
  not g14363 (n_5856, n8812);
  and g14364 (n8813, n_5855, n_5856);
  and g14365 (n8814, n_282, n_5851);
  and g14366 (n8815, n_5852, n8814);
  not g14367 (n_5857, n8813);
  not g14368 (n_5858, n8815);
  and g14369 (n8816, n_5857, n_5858);
  not g14370 (n_5859, n8806);
  not g14371 (n_5860, n8816);
  and g14372 (n8817, n_5859, n_5860);
  not g14373 (n_5861, n8817);
  and g14374 (n8818, \asqrt[59] , n_5861);
  and g14378 (n8822, n_5555, n_5554);
  and g14379 (n8823, \asqrt[27] , n8822);
  not g14380 (n_5862, n8823);
  and g14381 (n8824, n_5553, n_5862);
  not g14382 (n_5863, n8821);
  not g14383 (n_5864, n8824);
  and g14384 (n8825, n_5863, n_5864);
  and g14385 (n8826, n_218, n_5859);
  and g14386 (n8827, n_5860, n8826);
  not g14387 (n_5865, n8825);
  not g14388 (n_5866, n8827);
  and g14389 (n8828, n_5865, n_5866);
  not g14390 (n_5867, n8818);
  not g14391 (n_5868, n8828);
  and g14392 (n8829, n_5867, n_5868);
  not g14393 (n_5869, n8829);
  and g14394 (n8830, \asqrt[60] , n_5869);
  and g14398 (n8834, n_5563, n_5562);
  and g14399 (n8835, \asqrt[27] , n8834);
  not g14400 (n_5870, n8835);
  and g14401 (n8836, n_5561, n_5870);
  not g14402 (n_5871, n8833);
  not g14403 (n_5872, n8836);
  and g14404 (n8837, n_5871, n_5872);
  and g14405 (n8838, n_162, n_5867);
  and g14406 (n8839, n_5868, n8838);
  not g14407 (n_5873, n8837);
  not g14408 (n_5874, n8839);
  and g14409 (n8840, n_5873, n_5874);
  not g14410 (n_5875, n8830);
  not g14411 (n_5876, n8840);
  and g14412 (n8841, n_5875, n_5876);
  not g14413 (n_5877, n8841);
  and g14414 (n8842, \asqrt[61] , n_5877);
  and g14418 (n8846, n_5571, n_5570);
  and g14419 (n8847, \asqrt[27] , n8846);
  not g14420 (n_5878, n8847);
  and g14421 (n8848, n_5569, n_5878);
  not g14422 (n_5879, n8845);
  not g14423 (n_5880, n8848);
  and g14424 (n8849, n_5879, n_5880);
  and g14425 (n8850, n_115, n_5875);
  and g14426 (n8851, n_5876, n8850);
  not g14427 (n_5881, n8849);
  not g14428 (n_5882, n8851);
  and g14429 (n8852, n_5881, n_5882);
  not g14430 (n_5883, n8842);
  not g14431 (n_5884, n8852);
  and g14432 (n8853, n_5883, n_5884);
  not g14433 (n_5885, n8853);
  and g14434 (n8854, \asqrt[62] , n_5885);
  and g14438 (n8858, n_5579, n_5578);
  and g14439 (n8859, \asqrt[27] , n8858);
  not g14440 (n_5886, n8859);
  and g14441 (n8860, n_5577, n_5886);
  not g14442 (n_5887, n8857);
  not g14443 (n_5888, n8860);
  and g14444 (n8861, n_5887, n_5888);
  and g14445 (n8862, n_76, n_5883);
  and g14446 (n8863, n_5884, n8862);
  not g14447 (n_5889, n8861);
  not g14448 (n_5890, n8863);
  and g14449 (n8864, n_5889, n_5890);
  not g14450 (n_5891, n8854);
  not g14451 (n_5892, n8864);
  and g14452 (n8865, n_5891, n_5892);
  and g14456 (n8869, n_5587, n_5586);
  and g14457 (n8870, \asqrt[27] , n8869);
  not g14458 (n_5893, n8870);
  and g14459 (n8871, n_5585, n_5893);
  not g14460 (n_5894, n8868);
  not g14461 (n_5895, n8871);
  and g14462 (n8872, n_5894, n_5895);
  and g14463 (n8873, n_5594, n_5593);
  and g14464 (n8874, \asqrt[27] , n8873);
  not g14467 (n_5897, n8872);
  not g14469 (n_5898, n8865);
  not g14471 (n_5899, n8877);
  and g14472 (n8878, n_21, n_5899);
  and g14473 (n8879, n_5891, n8872);
  and g14474 (n8880, n_5892, n8879);
  and g14475 (n8881, n_5593, \asqrt[27] );
  not g14476 (n_5900, n8881);
  and g14477 (n8882, n8413, n_5900);
  not g14478 (n_5901, n8873);
  and g14479 (n8883, \asqrt[63] , n_5901);
  not g14480 (n_5902, n8882);
  and g14481 (n8884, n_5902, n8883);
  not g14487 (n_5903, n8884);
  not g14488 (n_5904, n8889);
  not g14490 (n_5905, n8880);
  and g14494 (n8893, \a[52] , \asqrt[26] );
  not g14495 (n_5910, \a[50] );
  not g14496 (n_5911, \a[51] );
  and g14497 (n8894, n_5910, n_5911);
  and g14498 (n8895, n_5606, n8894);
  not g14499 (n_5912, n8893);
  not g14500 (n_5913, n8895);
  and g14501 (n8896, n_5912, n_5913);
  not g14502 (n_5914, n8896);
  and g14503 (n8897, \asqrt[27] , n_5914);
  and g14509 (n8903, n_5606, \asqrt[26] );
  not g14510 (n_5915, n8903);
  and g14511 (n8904, \a[53] , n_5915);
  and g14512 (n8905, n8442, \asqrt[26] );
  not g14513 (n_5916, n8904);
  not g14514 (n_5917, n8905);
  and g14515 (n8906, n_5916, n_5917);
  not g14516 (n_5918, n8902);
  and g14517 (n8907, n_5918, n8906);
  not g14518 (n_5919, n8897);
  not g14519 (n_5920, n8907);
  and g14520 (n8908, n_5919, n_5920);
  not g14521 (n_5921, n8908);
  and g14522 (n8909, \asqrt[28] , n_5921);
  not g14523 (n_5922, \asqrt[28] );
  and g14524 (n8910, n_5922, n_5919);
  and g14525 (n8911, n_5920, n8910);
  not g14529 (n_5923, n8878);
  not g14531 (n_5924, n8915);
  and g14532 (n8916, n_5917, n_5924);
  not g14533 (n_5925, n8916);
  and g14534 (n8917, \a[54] , n_5925);
  and g14535 (n8918, n_5310, n_5924);
  and g14536 (n8919, n_5917, n8918);
  not g14537 (n_5926, n8917);
  not g14538 (n_5927, n8919);
  and g14539 (n8920, n_5926, n_5927);
  not g14540 (n_5928, n8911);
  not g14541 (n_5929, n8920);
  and g14542 (n8921, n_5928, n_5929);
  not g14543 (n_5930, n8909);
  not g14544 (n_5931, n8921);
  and g14545 (n8922, n_5930, n_5931);
  not g14546 (n_5932, n8922);
  and g14547 (n8923, \asqrt[29] , n_5932);
  and g14548 (n8924, n_5615, n_5614);
  not g14549 (n_5933, n8454);
  and g14550 (n8925, n_5933, n8924);
  and g14551 (n8926, \asqrt[26] , n8925);
  and g14552 (n8927, \asqrt[26] , n8924);
  not g14553 (n_5934, n8927);
  and g14554 (n8928, n8454, n_5934);
  not g14555 (n_5935, n8926);
  not g14556 (n_5936, n8928);
  and g14557 (n8929, n_5935, n_5936);
  and g14558 (n8930, n_5618, n_5930);
  and g14559 (n8931, n_5931, n8930);
  not g14560 (n_5937, n8929);
  not g14561 (n_5938, n8931);
  and g14562 (n8932, n_5937, n_5938);
  not g14563 (n_5939, n8923);
  not g14564 (n_5940, n8932);
  and g14565 (n8933, n_5939, n_5940);
  not g14566 (n_5941, n8933);
  and g14567 (n8934, \asqrt[30] , n_5941);
  and g14571 (n8938, n_5626, n_5624);
  and g14572 (n8939, \asqrt[26] , n8938);
  not g14573 (n_5942, n8939);
  and g14574 (n8940, n_5625, n_5942);
  not g14575 (n_5943, n8937);
  not g14576 (n_5944, n8940);
  and g14577 (n8941, n_5943, n_5944);
  and g14578 (n8942, n_5322, n_5939);
  and g14579 (n8943, n_5940, n8942);
  not g14580 (n_5945, n8941);
  not g14581 (n_5946, n8943);
  and g14582 (n8944, n_5945, n_5946);
  not g14583 (n_5947, n8934);
  not g14584 (n_5948, n8944);
  and g14585 (n8945, n_5947, n_5948);
  not g14586 (n_5949, n8945);
  and g14587 (n8946, \asqrt[31] , n_5949);
  and g14591 (n8950, n_5635, n_5634);
  and g14592 (n8951, \asqrt[26] , n8950);
  not g14593 (n_5950, n8951);
  and g14594 (n8952, n_5633, n_5950);
  not g14595 (n_5951, n8949);
  not g14596 (n_5952, n8952);
  and g14597 (n8953, n_5951, n_5952);
  and g14598 (n8954, n_5034, n_5947);
  and g14599 (n8955, n_5948, n8954);
  not g14600 (n_5953, n8953);
  not g14601 (n_5954, n8955);
  and g14602 (n8956, n_5953, n_5954);
  not g14603 (n_5955, n8946);
  not g14604 (n_5956, n8956);
  and g14605 (n8957, n_5955, n_5956);
  not g14606 (n_5957, n8957);
  and g14607 (n8958, \asqrt[32] , n_5957);
  and g14611 (n8962, n_5643, n_5642);
  and g14612 (n8963, \asqrt[26] , n8962);
  not g14613 (n_5958, n8963);
  and g14614 (n8964, n_5641, n_5958);
  not g14615 (n_5959, n8961);
  not g14616 (n_5960, n8964);
  and g14617 (n8965, n_5959, n_5960);
  and g14618 (n8966, n_4754, n_5955);
  and g14619 (n8967, n_5956, n8966);
  not g14620 (n_5961, n8965);
  not g14621 (n_5962, n8967);
  and g14622 (n8968, n_5961, n_5962);
  not g14623 (n_5963, n8958);
  not g14624 (n_5964, n8968);
  and g14625 (n8969, n_5963, n_5964);
  not g14626 (n_5965, n8969);
  and g14627 (n8970, \asqrt[33] , n_5965);
  and g14631 (n8974, n_5651, n_5650);
  and g14632 (n8975, \asqrt[26] , n8974);
  not g14633 (n_5966, n8975);
  and g14634 (n8976, n_5649, n_5966);
  not g14635 (n_5967, n8973);
  not g14636 (n_5968, n8976);
  and g14637 (n8977, n_5967, n_5968);
  and g14638 (n8978, n_4482, n_5963);
  and g14639 (n8979, n_5964, n8978);
  not g14640 (n_5969, n8977);
  not g14641 (n_5970, n8979);
  and g14642 (n8980, n_5969, n_5970);
  not g14643 (n_5971, n8970);
  not g14644 (n_5972, n8980);
  and g14645 (n8981, n_5971, n_5972);
  not g14646 (n_5973, n8981);
  and g14647 (n8982, \asqrt[34] , n_5973);
  and g14651 (n8986, n_5659, n_5658);
  and g14652 (n8987, \asqrt[26] , n8986);
  not g14653 (n_5974, n8987);
  and g14654 (n8988, n_5657, n_5974);
  not g14655 (n_5975, n8985);
  not g14656 (n_5976, n8988);
  and g14657 (n8989, n_5975, n_5976);
  and g14658 (n8990, n_4218, n_5971);
  and g14659 (n8991, n_5972, n8990);
  not g14660 (n_5977, n8989);
  not g14661 (n_5978, n8991);
  and g14662 (n8992, n_5977, n_5978);
  not g14663 (n_5979, n8982);
  not g14664 (n_5980, n8992);
  and g14665 (n8993, n_5979, n_5980);
  not g14666 (n_5981, n8993);
  and g14667 (n8994, \asqrt[35] , n_5981);
  and g14671 (n8998, n_5667, n_5666);
  and g14672 (n8999, \asqrt[26] , n8998);
  not g14673 (n_5982, n8999);
  and g14674 (n9000, n_5665, n_5982);
  not g14675 (n_5983, n8997);
  not g14676 (n_5984, n9000);
  and g14677 (n9001, n_5983, n_5984);
  and g14678 (n9002, n_3962, n_5979);
  and g14679 (n9003, n_5980, n9002);
  not g14680 (n_5985, n9001);
  not g14681 (n_5986, n9003);
  and g14682 (n9004, n_5985, n_5986);
  not g14683 (n_5987, n8994);
  not g14684 (n_5988, n9004);
  and g14685 (n9005, n_5987, n_5988);
  not g14686 (n_5989, n9005);
  and g14687 (n9006, \asqrt[36] , n_5989);
  and g14691 (n9010, n_5675, n_5674);
  and g14692 (n9011, \asqrt[26] , n9010);
  not g14693 (n_5990, n9011);
  and g14694 (n9012, n_5673, n_5990);
  not g14695 (n_5991, n9009);
  not g14696 (n_5992, n9012);
  and g14697 (n9013, n_5991, n_5992);
  and g14698 (n9014, n_3714, n_5987);
  and g14699 (n9015, n_5988, n9014);
  not g14700 (n_5993, n9013);
  not g14701 (n_5994, n9015);
  and g14702 (n9016, n_5993, n_5994);
  not g14703 (n_5995, n9006);
  not g14704 (n_5996, n9016);
  and g14705 (n9017, n_5995, n_5996);
  not g14706 (n_5997, n9017);
  and g14707 (n9018, \asqrt[37] , n_5997);
  and g14711 (n9022, n_5683, n_5682);
  and g14712 (n9023, \asqrt[26] , n9022);
  not g14713 (n_5998, n9023);
  and g14714 (n9024, n_5681, n_5998);
  not g14715 (n_5999, n9021);
  not g14716 (n_6000, n9024);
  and g14717 (n9025, n_5999, n_6000);
  and g14718 (n9026, n_3474, n_5995);
  and g14719 (n9027, n_5996, n9026);
  not g14720 (n_6001, n9025);
  not g14721 (n_6002, n9027);
  and g14722 (n9028, n_6001, n_6002);
  not g14723 (n_6003, n9018);
  not g14724 (n_6004, n9028);
  and g14725 (n9029, n_6003, n_6004);
  not g14726 (n_6005, n9029);
  and g14727 (n9030, \asqrt[38] , n_6005);
  and g14731 (n9034, n_5691, n_5690);
  and g14732 (n9035, \asqrt[26] , n9034);
  not g14733 (n_6006, n9035);
  and g14734 (n9036, n_5689, n_6006);
  not g14735 (n_6007, n9033);
  not g14736 (n_6008, n9036);
  and g14737 (n9037, n_6007, n_6008);
  and g14738 (n9038, n_3242, n_6003);
  and g14739 (n9039, n_6004, n9038);
  not g14740 (n_6009, n9037);
  not g14741 (n_6010, n9039);
  and g14742 (n9040, n_6009, n_6010);
  not g14743 (n_6011, n9030);
  not g14744 (n_6012, n9040);
  and g14745 (n9041, n_6011, n_6012);
  not g14746 (n_6013, n9041);
  and g14747 (n9042, \asqrt[39] , n_6013);
  and g14748 (n9043, n_3018, n_6011);
  and g14749 (n9044, n_6012, n9043);
  and g14753 (n9048, n_5699, n_5697);
  and g14754 (n9049, \asqrt[26] , n9048);
  not g14755 (n_6014, n9049);
  and g14756 (n9050, n_5698, n_6014);
  not g14757 (n_6015, n9047);
  not g14758 (n_6016, n9050);
  and g14759 (n9051, n_6015, n_6016);
  not g14760 (n_6017, n9044);
  not g14761 (n_6018, n9051);
  and g14762 (n9052, n_6017, n_6018);
  not g14763 (n_6019, n9042);
  not g14764 (n_6020, n9052);
  and g14765 (n9053, n_6019, n_6020);
  not g14766 (n_6021, n9053);
  and g14767 (n9054, \asqrt[40] , n_6021);
  and g14771 (n9058, n_5707, n_5706);
  and g14772 (n9059, \asqrt[26] , n9058);
  not g14773 (n_6022, n9059);
  and g14774 (n9060, n_5705, n_6022);
  not g14775 (n_6023, n9057);
  not g14776 (n_6024, n9060);
  and g14777 (n9061, n_6023, n_6024);
  and g14778 (n9062, n_2802, n_6019);
  and g14779 (n9063, n_6020, n9062);
  not g14780 (n_6025, n9061);
  not g14781 (n_6026, n9063);
  and g14782 (n9064, n_6025, n_6026);
  not g14783 (n_6027, n9054);
  not g14784 (n_6028, n9064);
  and g14785 (n9065, n_6027, n_6028);
  not g14786 (n_6029, n9065);
  and g14787 (n9066, \asqrt[41] , n_6029);
  and g14791 (n9070, n_5715, n_5714);
  and g14792 (n9071, \asqrt[26] , n9070);
  not g14793 (n_6030, n9071);
  and g14794 (n9072, n_5713, n_6030);
  not g14795 (n_6031, n9069);
  not g14796 (n_6032, n9072);
  and g14797 (n9073, n_6031, n_6032);
  and g14798 (n9074, n_2594, n_6027);
  and g14799 (n9075, n_6028, n9074);
  not g14800 (n_6033, n9073);
  not g14801 (n_6034, n9075);
  and g14802 (n9076, n_6033, n_6034);
  not g14803 (n_6035, n9066);
  not g14804 (n_6036, n9076);
  and g14805 (n9077, n_6035, n_6036);
  not g14806 (n_6037, n9077);
  and g14807 (n9078, \asqrt[42] , n_6037);
  and g14811 (n9082, n_5723, n_5722);
  and g14812 (n9083, \asqrt[26] , n9082);
  not g14813 (n_6038, n9083);
  and g14814 (n9084, n_5721, n_6038);
  not g14815 (n_6039, n9081);
  not g14816 (n_6040, n9084);
  and g14817 (n9085, n_6039, n_6040);
  and g14818 (n9086, n_2394, n_6035);
  and g14819 (n9087, n_6036, n9086);
  not g14820 (n_6041, n9085);
  not g14821 (n_6042, n9087);
  and g14822 (n9088, n_6041, n_6042);
  not g14823 (n_6043, n9078);
  not g14824 (n_6044, n9088);
  and g14825 (n9089, n_6043, n_6044);
  not g14826 (n_6045, n9089);
  and g14827 (n9090, \asqrt[43] , n_6045);
  and g14831 (n9094, n_5731, n_5730);
  and g14832 (n9095, \asqrt[26] , n9094);
  not g14833 (n_6046, n9095);
  and g14834 (n9096, n_5729, n_6046);
  not g14835 (n_6047, n9093);
  not g14836 (n_6048, n9096);
  and g14837 (n9097, n_6047, n_6048);
  and g14838 (n9098, n_2202, n_6043);
  and g14839 (n9099, n_6044, n9098);
  not g14840 (n_6049, n9097);
  not g14841 (n_6050, n9099);
  and g14842 (n9100, n_6049, n_6050);
  not g14843 (n_6051, n9090);
  not g14844 (n_6052, n9100);
  and g14845 (n9101, n_6051, n_6052);
  not g14846 (n_6053, n9101);
  and g14847 (n9102, \asqrt[44] , n_6053);
  and g14851 (n9106, n_5739, n_5738);
  and g14852 (n9107, \asqrt[26] , n9106);
  not g14853 (n_6054, n9107);
  and g14854 (n9108, n_5737, n_6054);
  not g14855 (n_6055, n9105);
  not g14856 (n_6056, n9108);
  and g14857 (n9109, n_6055, n_6056);
  and g14858 (n9110, n_2018, n_6051);
  and g14859 (n9111, n_6052, n9110);
  not g14860 (n_6057, n9109);
  not g14861 (n_6058, n9111);
  and g14862 (n9112, n_6057, n_6058);
  not g14863 (n_6059, n9102);
  not g14864 (n_6060, n9112);
  and g14865 (n9113, n_6059, n_6060);
  not g14866 (n_6061, n9113);
  and g14867 (n9114, \asqrt[45] , n_6061);
  and g14871 (n9118, n_5747, n_5746);
  and g14872 (n9119, \asqrt[26] , n9118);
  not g14873 (n_6062, n9119);
  and g14874 (n9120, n_5745, n_6062);
  not g14875 (n_6063, n9117);
  not g14876 (n_6064, n9120);
  and g14877 (n9121, n_6063, n_6064);
  and g14878 (n9122, n_1842, n_6059);
  and g14879 (n9123, n_6060, n9122);
  not g14880 (n_6065, n9121);
  not g14881 (n_6066, n9123);
  and g14882 (n9124, n_6065, n_6066);
  not g14883 (n_6067, n9114);
  not g14884 (n_6068, n9124);
  and g14885 (n9125, n_6067, n_6068);
  not g14886 (n_6069, n9125);
  and g14887 (n9126, \asqrt[46] , n_6069);
  and g14891 (n9130, n_5755, n_5754);
  and g14892 (n9131, \asqrt[26] , n9130);
  not g14893 (n_6070, n9131);
  and g14894 (n9132, n_5753, n_6070);
  not g14895 (n_6071, n9129);
  not g14896 (n_6072, n9132);
  and g14897 (n9133, n_6071, n_6072);
  and g14898 (n9134, n_1674, n_6067);
  and g14899 (n9135, n_6068, n9134);
  not g14900 (n_6073, n9133);
  not g14901 (n_6074, n9135);
  and g14902 (n9136, n_6073, n_6074);
  not g14903 (n_6075, n9126);
  not g14904 (n_6076, n9136);
  and g14905 (n9137, n_6075, n_6076);
  not g14906 (n_6077, n9137);
  and g14907 (n9138, \asqrt[47] , n_6077);
  and g14911 (n9142, n_5763, n_5762);
  and g14912 (n9143, \asqrt[26] , n9142);
  not g14913 (n_6078, n9143);
  and g14914 (n9144, n_5761, n_6078);
  not g14915 (n_6079, n9141);
  not g14916 (n_6080, n9144);
  and g14917 (n9145, n_6079, n_6080);
  and g14918 (n9146, n_1514, n_6075);
  and g14919 (n9147, n_6076, n9146);
  not g14920 (n_6081, n9145);
  not g14921 (n_6082, n9147);
  and g14922 (n9148, n_6081, n_6082);
  not g14923 (n_6083, n9138);
  not g14924 (n_6084, n9148);
  and g14925 (n9149, n_6083, n_6084);
  not g14926 (n_6085, n9149);
  and g14927 (n9150, \asqrt[48] , n_6085);
  and g14931 (n9154, n_5771, n_5770);
  and g14932 (n9155, \asqrt[26] , n9154);
  not g14933 (n_6086, n9155);
  and g14934 (n9156, n_5769, n_6086);
  not g14935 (n_6087, n9153);
  not g14936 (n_6088, n9156);
  and g14937 (n9157, n_6087, n_6088);
  and g14938 (n9158, n_1362, n_6083);
  and g14939 (n9159, n_6084, n9158);
  not g14940 (n_6089, n9157);
  not g14941 (n_6090, n9159);
  and g14942 (n9160, n_6089, n_6090);
  not g14943 (n_6091, n9150);
  not g14944 (n_6092, n9160);
  and g14945 (n9161, n_6091, n_6092);
  not g14946 (n_6093, n9161);
  and g14947 (n9162, \asqrt[49] , n_6093);
  and g14951 (n9166, n_5779, n_5778);
  and g14952 (n9167, \asqrt[26] , n9166);
  not g14953 (n_6094, n9167);
  and g14954 (n9168, n_5777, n_6094);
  not g14955 (n_6095, n9165);
  not g14956 (n_6096, n9168);
  and g14957 (n9169, n_6095, n_6096);
  and g14958 (n9170, n_1218, n_6091);
  and g14959 (n9171, n_6092, n9170);
  not g14960 (n_6097, n9169);
  not g14961 (n_6098, n9171);
  and g14962 (n9172, n_6097, n_6098);
  not g14963 (n_6099, n9162);
  not g14964 (n_6100, n9172);
  and g14965 (n9173, n_6099, n_6100);
  not g14966 (n_6101, n9173);
  and g14967 (n9174, \asqrt[50] , n_6101);
  and g14971 (n9178, n_5787, n_5786);
  and g14972 (n9179, \asqrt[26] , n9178);
  not g14973 (n_6102, n9179);
  and g14974 (n9180, n_5785, n_6102);
  not g14975 (n_6103, n9177);
  not g14976 (n_6104, n9180);
  and g14977 (n9181, n_6103, n_6104);
  and g14978 (n9182, n_1082, n_6099);
  and g14979 (n9183, n_6100, n9182);
  not g14980 (n_6105, n9181);
  not g14981 (n_6106, n9183);
  and g14982 (n9184, n_6105, n_6106);
  not g14983 (n_6107, n9174);
  not g14984 (n_6108, n9184);
  and g14985 (n9185, n_6107, n_6108);
  not g14986 (n_6109, n9185);
  and g14987 (n9186, \asqrt[51] , n_6109);
  and g14991 (n9190, n_5795, n_5794);
  and g14992 (n9191, \asqrt[26] , n9190);
  not g14993 (n_6110, n9191);
  and g14994 (n9192, n_5793, n_6110);
  not g14995 (n_6111, n9189);
  not g14996 (n_6112, n9192);
  and g14997 (n9193, n_6111, n_6112);
  and g14998 (n9194, n_954, n_6107);
  and g14999 (n9195, n_6108, n9194);
  not g15000 (n_6113, n9193);
  not g15001 (n_6114, n9195);
  and g15002 (n9196, n_6113, n_6114);
  not g15003 (n_6115, n9186);
  not g15004 (n_6116, n9196);
  and g15005 (n9197, n_6115, n_6116);
  not g15006 (n_6117, n9197);
  and g15007 (n9198, \asqrt[52] , n_6117);
  and g15011 (n9202, n_5803, n_5802);
  and g15012 (n9203, \asqrt[26] , n9202);
  not g15013 (n_6118, n9203);
  and g15014 (n9204, n_5801, n_6118);
  not g15015 (n_6119, n9201);
  not g15016 (n_6120, n9204);
  and g15017 (n9205, n_6119, n_6120);
  and g15018 (n9206, n_834, n_6115);
  and g15019 (n9207, n_6116, n9206);
  not g15020 (n_6121, n9205);
  not g15021 (n_6122, n9207);
  and g15022 (n9208, n_6121, n_6122);
  not g15023 (n_6123, n9198);
  not g15024 (n_6124, n9208);
  and g15025 (n9209, n_6123, n_6124);
  not g15026 (n_6125, n9209);
  and g15027 (n9210, \asqrt[53] , n_6125);
  and g15031 (n9214, n_5811, n_5810);
  and g15032 (n9215, \asqrt[26] , n9214);
  not g15033 (n_6126, n9215);
  and g15034 (n9216, n_5809, n_6126);
  not g15035 (n_6127, n9213);
  not g15036 (n_6128, n9216);
  and g15037 (n9217, n_6127, n_6128);
  and g15038 (n9218, n_722, n_6123);
  and g15039 (n9219, n_6124, n9218);
  not g15040 (n_6129, n9217);
  not g15041 (n_6130, n9219);
  and g15042 (n9220, n_6129, n_6130);
  not g15043 (n_6131, n9210);
  not g15044 (n_6132, n9220);
  and g15045 (n9221, n_6131, n_6132);
  not g15046 (n_6133, n9221);
  and g15047 (n9222, \asqrt[54] , n_6133);
  and g15051 (n9226, n_5819, n_5818);
  and g15052 (n9227, \asqrt[26] , n9226);
  not g15053 (n_6134, n9227);
  and g15054 (n9228, n_5817, n_6134);
  not g15055 (n_6135, n9225);
  not g15056 (n_6136, n9228);
  and g15057 (n9229, n_6135, n_6136);
  and g15058 (n9230, n_618, n_6131);
  and g15059 (n9231, n_6132, n9230);
  not g15060 (n_6137, n9229);
  not g15061 (n_6138, n9231);
  and g15062 (n9232, n_6137, n_6138);
  not g15063 (n_6139, n9222);
  not g15064 (n_6140, n9232);
  and g15065 (n9233, n_6139, n_6140);
  not g15066 (n_6141, n9233);
  and g15067 (n9234, \asqrt[55] , n_6141);
  and g15071 (n9238, n_5827, n_5826);
  and g15072 (n9239, \asqrt[26] , n9238);
  not g15073 (n_6142, n9239);
  and g15074 (n9240, n_5825, n_6142);
  not g15075 (n_6143, n9237);
  not g15076 (n_6144, n9240);
  and g15077 (n9241, n_6143, n_6144);
  and g15078 (n9242, n_522, n_6139);
  and g15079 (n9243, n_6140, n9242);
  not g15080 (n_6145, n9241);
  not g15081 (n_6146, n9243);
  and g15082 (n9244, n_6145, n_6146);
  not g15083 (n_6147, n9234);
  not g15084 (n_6148, n9244);
  and g15085 (n9245, n_6147, n_6148);
  not g15086 (n_6149, n9245);
  and g15087 (n9246, \asqrt[56] , n_6149);
  and g15091 (n9250, n_5835, n_5834);
  and g15092 (n9251, \asqrt[26] , n9250);
  not g15093 (n_6150, n9251);
  and g15094 (n9252, n_5833, n_6150);
  not g15095 (n_6151, n9249);
  not g15096 (n_6152, n9252);
  and g15097 (n9253, n_6151, n_6152);
  and g15098 (n9254, n_434, n_6147);
  and g15099 (n9255, n_6148, n9254);
  not g15100 (n_6153, n9253);
  not g15101 (n_6154, n9255);
  and g15102 (n9256, n_6153, n_6154);
  not g15103 (n_6155, n9246);
  not g15104 (n_6156, n9256);
  and g15105 (n9257, n_6155, n_6156);
  not g15106 (n_6157, n9257);
  and g15107 (n9258, \asqrt[57] , n_6157);
  and g15111 (n9262, n_5843, n_5842);
  and g15112 (n9263, \asqrt[26] , n9262);
  not g15113 (n_6158, n9263);
  and g15114 (n9264, n_5841, n_6158);
  not g15115 (n_6159, n9261);
  not g15116 (n_6160, n9264);
  and g15117 (n9265, n_6159, n_6160);
  and g15118 (n9266, n_354, n_6155);
  and g15119 (n9267, n_6156, n9266);
  not g15120 (n_6161, n9265);
  not g15121 (n_6162, n9267);
  and g15122 (n9268, n_6161, n_6162);
  not g15123 (n_6163, n9258);
  not g15124 (n_6164, n9268);
  and g15125 (n9269, n_6163, n_6164);
  not g15126 (n_6165, n9269);
  and g15127 (n9270, \asqrt[58] , n_6165);
  and g15131 (n9274, n_5851, n_5850);
  and g15132 (n9275, \asqrt[26] , n9274);
  not g15133 (n_6166, n9275);
  and g15134 (n9276, n_5849, n_6166);
  not g15135 (n_6167, n9273);
  not g15136 (n_6168, n9276);
  and g15137 (n9277, n_6167, n_6168);
  and g15138 (n9278, n_282, n_6163);
  and g15139 (n9279, n_6164, n9278);
  not g15140 (n_6169, n9277);
  not g15141 (n_6170, n9279);
  and g15142 (n9280, n_6169, n_6170);
  not g15143 (n_6171, n9270);
  not g15144 (n_6172, n9280);
  and g15145 (n9281, n_6171, n_6172);
  not g15146 (n_6173, n9281);
  and g15147 (n9282, \asqrt[59] , n_6173);
  and g15151 (n9286, n_5859, n_5858);
  and g15152 (n9287, \asqrt[26] , n9286);
  not g15153 (n_6174, n9287);
  and g15154 (n9288, n_5857, n_6174);
  not g15155 (n_6175, n9285);
  not g15156 (n_6176, n9288);
  and g15157 (n9289, n_6175, n_6176);
  and g15158 (n9290, n_218, n_6171);
  and g15159 (n9291, n_6172, n9290);
  not g15160 (n_6177, n9289);
  not g15161 (n_6178, n9291);
  and g15162 (n9292, n_6177, n_6178);
  not g15163 (n_6179, n9282);
  not g15164 (n_6180, n9292);
  and g15165 (n9293, n_6179, n_6180);
  not g15166 (n_6181, n9293);
  and g15167 (n9294, \asqrt[60] , n_6181);
  and g15171 (n9298, n_5867, n_5866);
  and g15172 (n9299, \asqrt[26] , n9298);
  not g15173 (n_6182, n9299);
  and g15174 (n9300, n_5865, n_6182);
  not g15175 (n_6183, n9297);
  not g15176 (n_6184, n9300);
  and g15177 (n9301, n_6183, n_6184);
  and g15178 (n9302, n_162, n_6179);
  and g15179 (n9303, n_6180, n9302);
  not g15180 (n_6185, n9301);
  not g15181 (n_6186, n9303);
  and g15182 (n9304, n_6185, n_6186);
  not g15183 (n_6187, n9294);
  not g15184 (n_6188, n9304);
  and g15185 (n9305, n_6187, n_6188);
  not g15186 (n_6189, n9305);
  and g15187 (n9306, \asqrt[61] , n_6189);
  and g15191 (n9310, n_5875, n_5874);
  and g15192 (n9311, \asqrt[26] , n9310);
  not g15193 (n_6190, n9311);
  and g15194 (n9312, n_5873, n_6190);
  not g15195 (n_6191, n9309);
  not g15196 (n_6192, n9312);
  and g15197 (n9313, n_6191, n_6192);
  and g15198 (n9314, n_115, n_6187);
  and g15199 (n9315, n_6188, n9314);
  not g15200 (n_6193, n9313);
  not g15201 (n_6194, n9315);
  and g15202 (n9316, n_6193, n_6194);
  not g15203 (n_6195, n9306);
  not g15204 (n_6196, n9316);
  and g15205 (n9317, n_6195, n_6196);
  not g15206 (n_6197, n9317);
  and g15207 (n9318, \asqrt[62] , n_6197);
  and g15211 (n9322, n_5883, n_5882);
  and g15212 (n9323, \asqrt[26] , n9322);
  not g15213 (n_6198, n9323);
  and g15214 (n9324, n_5881, n_6198);
  not g15215 (n_6199, n9321);
  not g15216 (n_6200, n9324);
  and g15217 (n9325, n_6199, n_6200);
  and g15218 (n9326, n_76, n_6195);
  and g15219 (n9327, n_6196, n9326);
  not g15220 (n_6201, n9325);
  not g15221 (n_6202, n9327);
  and g15222 (n9328, n_6201, n_6202);
  not g15223 (n_6203, n9318);
  not g15224 (n_6204, n9328);
  and g15225 (n9329, n_6203, n_6204);
  and g15229 (n9333, n_5891, n_5890);
  and g15230 (n9334, \asqrt[26] , n9333);
  not g15231 (n_6205, n9334);
  and g15232 (n9335, n_5889, n_6205);
  not g15233 (n_6206, n9332);
  not g15234 (n_6207, n9335);
  and g15235 (n9336, n_6206, n_6207);
  and g15236 (n9337, n_5898, n_5897);
  and g15237 (n9338, \asqrt[26] , n9337);
  not g15240 (n_6209, n9336);
  not g15242 (n_6210, n9329);
  not g15244 (n_6211, n9341);
  and g15245 (n9342, n_21, n_6211);
  and g15246 (n9343, n_6203, n9336);
  and g15247 (n9344, n_6204, n9343);
  and g15248 (n9345, n_5897, \asqrt[26] );
  not g15249 (n_6212, n9345);
  and g15250 (n9346, n8865, n_6212);
  not g15251 (n_6213, n9337);
  and g15252 (n9347, \asqrt[63] , n_6213);
  not g15253 (n_6214, n9346);
  and g15254 (n9348, n_6214, n9347);
  not g15260 (n_6215, n9348);
  not g15261 (n_6216, n9353);
  not g15263 (n_6217, n9344);
  and g15267 (n9357, \a[50] , \asqrt[25] );
  not g15268 (n_6222, \a[48] );
  not g15269 (n_6223, \a[49] );
  and g15270 (n9358, n_6222, n_6223);
  and g15271 (n9359, n_5910, n9358);
  not g15272 (n_6224, n9357);
  not g15273 (n_6225, n9359);
  and g15274 (n9360, n_6224, n_6225);
  not g15275 (n_6226, n9360);
  and g15276 (n9361, \asqrt[26] , n_6226);
  and g15282 (n9367, n_5910, \asqrt[25] );
  not g15283 (n_6227, n9367);
  and g15284 (n9368, \a[51] , n_6227);
  and g15285 (n9369, n8894, \asqrt[25] );
  not g15286 (n_6228, n9368);
  not g15287 (n_6229, n9369);
  and g15288 (n9370, n_6228, n_6229);
  not g15289 (n_6230, n9366);
  and g15290 (n9371, n_6230, n9370);
  not g15291 (n_6231, n9361);
  not g15292 (n_6232, n9371);
  and g15293 (n9372, n_6231, n_6232);
  not g15294 (n_6233, n9372);
  and g15295 (n9373, \asqrt[27] , n_6233);
  not g15296 (n_6234, \asqrt[27] );
  and g15297 (n9374, n_6234, n_6231);
  and g15298 (n9375, n_6232, n9374);
  not g15302 (n_6235, n9342);
  not g15304 (n_6236, n9379);
  and g15305 (n9380, n_6229, n_6236);
  not g15306 (n_6237, n9380);
  and g15307 (n9381, \a[52] , n_6237);
  and g15308 (n9382, n_5606, n_6236);
  and g15309 (n9383, n_6229, n9382);
  not g15310 (n_6238, n9381);
  not g15311 (n_6239, n9383);
  and g15312 (n9384, n_6238, n_6239);
  not g15313 (n_6240, n9375);
  not g15314 (n_6241, n9384);
  and g15315 (n9385, n_6240, n_6241);
  not g15316 (n_6242, n9373);
  not g15317 (n_6243, n9385);
  and g15318 (n9386, n_6242, n_6243);
  not g15319 (n_6244, n9386);
  and g15320 (n9387, \asqrt[28] , n_6244);
  and g15321 (n9388, n_5919, n_5918);
  not g15322 (n_6245, n8906);
  and g15323 (n9389, n_6245, n9388);
  and g15324 (n9390, \asqrt[25] , n9389);
  and g15325 (n9391, \asqrt[25] , n9388);
  not g15326 (n_6246, n9391);
  and g15327 (n9392, n8906, n_6246);
  not g15328 (n_6247, n9390);
  not g15329 (n_6248, n9392);
  and g15330 (n9393, n_6247, n_6248);
  and g15331 (n9394, n_5922, n_6242);
  and g15332 (n9395, n_6243, n9394);
  not g15333 (n_6249, n9393);
  not g15334 (n_6250, n9395);
  and g15335 (n9396, n_6249, n_6250);
  not g15336 (n_6251, n9387);
  not g15337 (n_6252, n9396);
  and g15338 (n9397, n_6251, n_6252);
  not g15339 (n_6253, n9397);
  and g15340 (n9398, \asqrt[29] , n_6253);
  and g15344 (n9402, n_5930, n_5928);
  and g15345 (n9403, \asqrt[25] , n9402);
  not g15346 (n_6254, n9403);
  and g15347 (n9404, n_5929, n_6254);
  not g15348 (n_6255, n9401);
  not g15349 (n_6256, n9404);
  and g15350 (n9405, n_6255, n_6256);
  and g15351 (n9406, n_5618, n_6251);
  and g15352 (n9407, n_6252, n9406);
  not g15353 (n_6257, n9405);
  not g15354 (n_6258, n9407);
  and g15355 (n9408, n_6257, n_6258);
  not g15356 (n_6259, n9398);
  not g15357 (n_6260, n9408);
  and g15358 (n9409, n_6259, n_6260);
  not g15359 (n_6261, n9409);
  and g15360 (n9410, \asqrt[30] , n_6261);
  and g15364 (n9414, n_5939, n_5938);
  and g15365 (n9415, \asqrt[25] , n9414);
  not g15366 (n_6262, n9415);
  and g15367 (n9416, n_5937, n_6262);
  not g15368 (n_6263, n9413);
  not g15369 (n_6264, n9416);
  and g15370 (n9417, n_6263, n_6264);
  and g15371 (n9418, n_5322, n_6259);
  and g15372 (n9419, n_6260, n9418);
  not g15373 (n_6265, n9417);
  not g15374 (n_6266, n9419);
  and g15375 (n9420, n_6265, n_6266);
  not g15376 (n_6267, n9410);
  not g15377 (n_6268, n9420);
  and g15378 (n9421, n_6267, n_6268);
  not g15379 (n_6269, n9421);
  and g15380 (n9422, \asqrt[31] , n_6269);
  and g15384 (n9426, n_5947, n_5946);
  and g15385 (n9427, \asqrt[25] , n9426);
  not g15386 (n_6270, n9427);
  and g15387 (n9428, n_5945, n_6270);
  not g15388 (n_6271, n9425);
  not g15389 (n_6272, n9428);
  and g15390 (n9429, n_6271, n_6272);
  and g15391 (n9430, n_5034, n_6267);
  and g15392 (n9431, n_6268, n9430);
  not g15393 (n_6273, n9429);
  not g15394 (n_6274, n9431);
  and g15395 (n9432, n_6273, n_6274);
  not g15396 (n_6275, n9422);
  not g15397 (n_6276, n9432);
  and g15398 (n9433, n_6275, n_6276);
  not g15399 (n_6277, n9433);
  and g15400 (n9434, \asqrt[32] , n_6277);
  and g15404 (n9438, n_5955, n_5954);
  and g15405 (n9439, \asqrt[25] , n9438);
  not g15406 (n_6278, n9439);
  and g15407 (n9440, n_5953, n_6278);
  not g15408 (n_6279, n9437);
  not g15409 (n_6280, n9440);
  and g15410 (n9441, n_6279, n_6280);
  and g15411 (n9442, n_4754, n_6275);
  and g15412 (n9443, n_6276, n9442);
  not g15413 (n_6281, n9441);
  not g15414 (n_6282, n9443);
  and g15415 (n9444, n_6281, n_6282);
  not g15416 (n_6283, n9434);
  not g15417 (n_6284, n9444);
  and g15418 (n9445, n_6283, n_6284);
  not g15419 (n_6285, n9445);
  and g15420 (n9446, \asqrt[33] , n_6285);
  and g15424 (n9450, n_5963, n_5962);
  and g15425 (n9451, \asqrt[25] , n9450);
  not g15426 (n_6286, n9451);
  and g15427 (n9452, n_5961, n_6286);
  not g15428 (n_6287, n9449);
  not g15429 (n_6288, n9452);
  and g15430 (n9453, n_6287, n_6288);
  and g15431 (n9454, n_4482, n_6283);
  and g15432 (n9455, n_6284, n9454);
  not g15433 (n_6289, n9453);
  not g15434 (n_6290, n9455);
  and g15435 (n9456, n_6289, n_6290);
  not g15436 (n_6291, n9446);
  not g15437 (n_6292, n9456);
  and g15438 (n9457, n_6291, n_6292);
  not g15439 (n_6293, n9457);
  and g15440 (n9458, \asqrt[34] , n_6293);
  and g15444 (n9462, n_5971, n_5970);
  and g15445 (n9463, \asqrt[25] , n9462);
  not g15446 (n_6294, n9463);
  and g15447 (n9464, n_5969, n_6294);
  not g15448 (n_6295, n9461);
  not g15449 (n_6296, n9464);
  and g15450 (n9465, n_6295, n_6296);
  and g15451 (n9466, n_4218, n_6291);
  and g15452 (n9467, n_6292, n9466);
  not g15453 (n_6297, n9465);
  not g15454 (n_6298, n9467);
  and g15455 (n9468, n_6297, n_6298);
  not g15456 (n_6299, n9458);
  not g15457 (n_6300, n9468);
  and g15458 (n9469, n_6299, n_6300);
  not g15459 (n_6301, n9469);
  and g15460 (n9470, \asqrt[35] , n_6301);
  and g15464 (n9474, n_5979, n_5978);
  and g15465 (n9475, \asqrt[25] , n9474);
  not g15466 (n_6302, n9475);
  and g15467 (n9476, n_5977, n_6302);
  not g15468 (n_6303, n9473);
  not g15469 (n_6304, n9476);
  and g15470 (n9477, n_6303, n_6304);
  and g15471 (n9478, n_3962, n_6299);
  and g15472 (n9479, n_6300, n9478);
  not g15473 (n_6305, n9477);
  not g15474 (n_6306, n9479);
  and g15475 (n9480, n_6305, n_6306);
  not g15476 (n_6307, n9470);
  not g15477 (n_6308, n9480);
  and g15478 (n9481, n_6307, n_6308);
  not g15479 (n_6309, n9481);
  and g15480 (n9482, \asqrt[36] , n_6309);
  and g15484 (n9486, n_5987, n_5986);
  and g15485 (n9487, \asqrt[25] , n9486);
  not g15486 (n_6310, n9487);
  and g15487 (n9488, n_5985, n_6310);
  not g15488 (n_6311, n9485);
  not g15489 (n_6312, n9488);
  and g15490 (n9489, n_6311, n_6312);
  and g15491 (n9490, n_3714, n_6307);
  and g15492 (n9491, n_6308, n9490);
  not g15493 (n_6313, n9489);
  not g15494 (n_6314, n9491);
  and g15495 (n9492, n_6313, n_6314);
  not g15496 (n_6315, n9482);
  not g15497 (n_6316, n9492);
  and g15498 (n9493, n_6315, n_6316);
  not g15499 (n_6317, n9493);
  and g15500 (n9494, \asqrt[37] , n_6317);
  and g15504 (n9498, n_5995, n_5994);
  and g15505 (n9499, \asqrt[25] , n9498);
  not g15506 (n_6318, n9499);
  and g15507 (n9500, n_5993, n_6318);
  not g15508 (n_6319, n9497);
  not g15509 (n_6320, n9500);
  and g15510 (n9501, n_6319, n_6320);
  and g15511 (n9502, n_3474, n_6315);
  and g15512 (n9503, n_6316, n9502);
  not g15513 (n_6321, n9501);
  not g15514 (n_6322, n9503);
  and g15515 (n9504, n_6321, n_6322);
  not g15516 (n_6323, n9494);
  not g15517 (n_6324, n9504);
  and g15518 (n9505, n_6323, n_6324);
  not g15519 (n_6325, n9505);
  and g15520 (n9506, \asqrt[38] , n_6325);
  and g15524 (n9510, n_6003, n_6002);
  and g15525 (n9511, \asqrt[25] , n9510);
  not g15526 (n_6326, n9511);
  and g15527 (n9512, n_6001, n_6326);
  not g15528 (n_6327, n9509);
  not g15529 (n_6328, n9512);
  and g15530 (n9513, n_6327, n_6328);
  and g15531 (n9514, n_3242, n_6323);
  and g15532 (n9515, n_6324, n9514);
  not g15533 (n_6329, n9513);
  not g15534 (n_6330, n9515);
  and g15535 (n9516, n_6329, n_6330);
  not g15536 (n_6331, n9506);
  not g15537 (n_6332, n9516);
  and g15538 (n9517, n_6331, n_6332);
  not g15539 (n_6333, n9517);
  and g15540 (n9518, \asqrt[39] , n_6333);
  and g15544 (n9522, n_6011, n_6010);
  and g15545 (n9523, \asqrt[25] , n9522);
  not g15546 (n_6334, n9523);
  and g15547 (n9524, n_6009, n_6334);
  not g15548 (n_6335, n9521);
  not g15549 (n_6336, n9524);
  and g15550 (n9525, n_6335, n_6336);
  and g15551 (n9526, n_3018, n_6331);
  and g15552 (n9527, n_6332, n9526);
  not g15553 (n_6337, n9525);
  not g15554 (n_6338, n9527);
  and g15555 (n9528, n_6337, n_6338);
  not g15556 (n_6339, n9518);
  not g15557 (n_6340, n9528);
  and g15558 (n9529, n_6339, n_6340);
  not g15559 (n_6341, n9529);
  and g15560 (n9530, \asqrt[40] , n_6341);
  and g15561 (n9531, n_2802, n_6339);
  and g15562 (n9532, n_6340, n9531);
  and g15566 (n9536, n_6019, n_6017);
  and g15567 (n9537, \asqrt[25] , n9536);
  not g15568 (n_6342, n9537);
  and g15569 (n9538, n_6018, n_6342);
  not g15570 (n_6343, n9535);
  not g15571 (n_6344, n9538);
  and g15572 (n9539, n_6343, n_6344);
  not g15573 (n_6345, n9532);
  not g15574 (n_6346, n9539);
  and g15575 (n9540, n_6345, n_6346);
  not g15576 (n_6347, n9530);
  not g15577 (n_6348, n9540);
  and g15578 (n9541, n_6347, n_6348);
  not g15579 (n_6349, n9541);
  and g15580 (n9542, \asqrt[41] , n_6349);
  and g15584 (n9546, n_6027, n_6026);
  and g15585 (n9547, \asqrt[25] , n9546);
  not g15586 (n_6350, n9547);
  and g15587 (n9548, n_6025, n_6350);
  not g15588 (n_6351, n9545);
  not g15589 (n_6352, n9548);
  and g15590 (n9549, n_6351, n_6352);
  and g15591 (n9550, n_2594, n_6347);
  and g15592 (n9551, n_6348, n9550);
  not g15593 (n_6353, n9549);
  not g15594 (n_6354, n9551);
  and g15595 (n9552, n_6353, n_6354);
  not g15596 (n_6355, n9542);
  not g15597 (n_6356, n9552);
  and g15598 (n9553, n_6355, n_6356);
  not g15599 (n_6357, n9553);
  and g15600 (n9554, \asqrt[42] , n_6357);
  and g15604 (n9558, n_6035, n_6034);
  and g15605 (n9559, \asqrt[25] , n9558);
  not g15606 (n_6358, n9559);
  and g15607 (n9560, n_6033, n_6358);
  not g15608 (n_6359, n9557);
  not g15609 (n_6360, n9560);
  and g15610 (n9561, n_6359, n_6360);
  and g15611 (n9562, n_2394, n_6355);
  and g15612 (n9563, n_6356, n9562);
  not g15613 (n_6361, n9561);
  not g15614 (n_6362, n9563);
  and g15615 (n9564, n_6361, n_6362);
  not g15616 (n_6363, n9554);
  not g15617 (n_6364, n9564);
  and g15618 (n9565, n_6363, n_6364);
  not g15619 (n_6365, n9565);
  and g15620 (n9566, \asqrt[43] , n_6365);
  and g15624 (n9570, n_6043, n_6042);
  and g15625 (n9571, \asqrt[25] , n9570);
  not g15626 (n_6366, n9571);
  and g15627 (n9572, n_6041, n_6366);
  not g15628 (n_6367, n9569);
  not g15629 (n_6368, n9572);
  and g15630 (n9573, n_6367, n_6368);
  and g15631 (n9574, n_2202, n_6363);
  and g15632 (n9575, n_6364, n9574);
  not g15633 (n_6369, n9573);
  not g15634 (n_6370, n9575);
  and g15635 (n9576, n_6369, n_6370);
  not g15636 (n_6371, n9566);
  not g15637 (n_6372, n9576);
  and g15638 (n9577, n_6371, n_6372);
  not g15639 (n_6373, n9577);
  and g15640 (n9578, \asqrt[44] , n_6373);
  and g15644 (n9582, n_6051, n_6050);
  and g15645 (n9583, \asqrt[25] , n9582);
  not g15646 (n_6374, n9583);
  and g15647 (n9584, n_6049, n_6374);
  not g15648 (n_6375, n9581);
  not g15649 (n_6376, n9584);
  and g15650 (n9585, n_6375, n_6376);
  and g15651 (n9586, n_2018, n_6371);
  and g15652 (n9587, n_6372, n9586);
  not g15653 (n_6377, n9585);
  not g15654 (n_6378, n9587);
  and g15655 (n9588, n_6377, n_6378);
  not g15656 (n_6379, n9578);
  not g15657 (n_6380, n9588);
  and g15658 (n9589, n_6379, n_6380);
  not g15659 (n_6381, n9589);
  and g15660 (n9590, \asqrt[45] , n_6381);
  and g15664 (n9594, n_6059, n_6058);
  and g15665 (n9595, \asqrt[25] , n9594);
  not g15666 (n_6382, n9595);
  and g15667 (n9596, n_6057, n_6382);
  not g15668 (n_6383, n9593);
  not g15669 (n_6384, n9596);
  and g15670 (n9597, n_6383, n_6384);
  and g15671 (n9598, n_1842, n_6379);
  and g15672 (n9599, n_6380, n9598);
  not g15673 (n_6385, n9597);
  not g15674 (n_6386, n9599);
  and g15675 (n9600, n_6385, n_6386);
  not g15676 (n_6387, n9590);
  not g15677 (n_6388, n9600);
  and g15678 (n9601, n_6387, n_6388);
  not g15679 (n_6389, n9601);
  and g15680 (n9602, \asqrt[46] , n_6389);
  and g15684 (n9606, n_6067, n_6066);
  and g15685 (n9607, \asqrt[25] , n9606);
  not g15686 (n_6390, n9607);
  and g15687 (n9608, n_6065, n_6390);
  not g15688 (n_6391, n9605);
  not g15689 (n_6392, n9608);
  and g15690 (n9609, n_6391, n_6392);
  and g15691 (n9610, n_1674, n_6387);
  and g15692 (n9611, n_6388, n9610);
  not g15693 (n_6393, n9609);
  not g15694 (n_6394, n9611);
  and g15695 (n9612, n_6393, n_6394);
  not g15696 (n_6395, n9602);
  not g15697 (n_6396, n9612);
  and g15698 (n9613, n_6395, n_6396);
  not g15699 (n_6397, n9613);
  and g15700 (n9614, \asqrt[47] , n_6397);
  and g15704 (n9618, n_6075, n_6074);
  and g15705 (n9619, \asqrt[25] , n9618);
  not g15706 (n_6398, n9619);
  and g15707 (n9620, n_6073, n_6398);
  not g15708 (n_6399, n9617);
  not g15709 (n_6400, n9620);
  and g15710 (n9621, n_6399, n_6400);
  and g15711 (n9622, n_1514, n_6395);
  and g15712 (n9623, n_6396, n9622);
  not g15713 (n_6401, n9621);
  not g15714 (n_6402, n9623);
  and g15715 (n9624, n_6401, n_6402);
  not g15716 (n_6403, n9614);
  not g15717 (n_6404, n9624);
  and g15718 (n9625, n_6403, n_6404);
  not g15719 (n_6405, n9625);
  and g15720 (n9626, \asqrt[48] , n_6405);
  and g15724 (n9630, n_6083, n_6082);
  and g15725 (n9631, \asqrt[25] , n9630);
  not g15726 (n_6406, n9631);
  and g15727 (n9632, n_6081, n_6406);
  not g15728 (n_6407, n9629);
  not g15729 (n_6408, n9632);
  and g15730 (n9633, n_6407, n_6408);
  and g15731 (n9634, n_1362, n_6403);
  and g15732 (n9635, n_6404, n9634);
  not g15733 (n_6409, n9633);
  not g15734 (n_6410, n9635);
  and g15735 (n9636, n_6409, n_6410);
  not g15736 (n_6411, n9626);
  not g15737 (n_6412, n9636);
  and g15738 (n9637, n_6411, n_6412);
  not g15739 (n_6413, n9637);
  and g15740 (n9638, \asqrt[49] , n_6413);
  and g15744 (n9642, n_6091, n_6090);
  and g15745 (n9643, \asqrt[25] , n9642);
  not g15746 (n_6414, n9643);
  and g15747 (n9644, n_6089, n_6414);
  not g15748 (n_6415, n9641);
  not g15749 (n_6416, n9644);
  and g15750 (n9645, n_6415, n_6416);
  and g15751 (n9646, n_1218, n_6411);
  and g15752 (n9647, n_6412, n9646);
  not g15753 (n_6417, n9645);
  not g15754 (n_6418, n9647);
  and g15755 (n9648, n_6417, n_6418);
  not g15756 (n_6419, n9638);
  not g15757 (n_6420, n9648);
  and g15758 (n9649, n_6419, n_6420);
  not g15759 (n_6421, n9649);
  and g15760 (n9650, \asqrt[50] , n_6421);
  and g15764 (n9654, n_6099, n_6098);
  and g15765 (n9655, \asqrt[25] , n9654);
  not g15766 (n_6422, n9655);
  and g15767 (n9656, n_6097, n_6422);
  not g15768 (n_6423, n9653);
  not g15769 (n_6424, n9656);
  and g15770 (n9657, n_6423, n_6424);
  and g15771 (n9658, n_1082, n_6419);
  and g15772 (n9659, n_6420, n9658);
  not g15773 (n_6425, n9657);
  not g15774 (n_6426, n9659);
  and g15775 (n9660, n_6425, n_6426);
  not g15776 (n_6427, n9650);
  not g15777 (n_6428, n9660);
  and g15778 (n9661, n_6427, n_6428);
  not g15779 (n_6429, n9661);
  and g15780 (n9662, \asqrt[51] , n_6429);
  and g15784 (n9666, n_6107, n_6106);
  and g15785 (n9667, \asqrt[25] , n9666);
  not g15786 (n_6430, n9667);
  and g15787 (n9668, n_6105, n_6430);
  not g15788 (n_6431, n9665);
  not g15789 (n_6432, n9668);
  and g15790 (n9669, n_6431, n_6432);
  and g15791 (n9670, n_954, n_6427);
  and g15792 (n9671, n_6428, n9670);
  not g15793 (n_6433, n9669);
  not g15794 (n_6434, n9671);
  and g15795 (n9672, n_6433, n_6434);
  not g15796 (n_6435, n9662);
  not g15797 (n_6436, n9672);
  and g15798 (n9673, n_6435, n_6436);
  not g15799 (n_6437, n9673);
  and g15800 (n9674, \asqrt[52] , n_6437);
  and g15804 (n9678, n_6115, n_6114);
  and g15805 (n9679, \asqrt[25] , n9678);
  not g15806 (n_6438, n9679);
  and g15807 (n9680, n_6113, n_6438);
  not g15808 (n_6439, n9677);
  not g15809 (n_6440, n9680);
  and g15810 (n9681, n_6439, n_6440);
  and g15811 (n9682, n_834, n_6435);
  and g15812 (n9683, n_6436, n9682);
  not g15813 (n_6441, n9681);
  not g15814 (n_6442, n9683);
  and g15815 (n9684, n_6441, n_6442);
  not g15816 (n_6443, n9674);
  not g15817 (n_6444, n9684);
  and g15818 (n9685, n_6443, n_6444);
  not g15819 (n_6445, n9685);
  and g15820 (n9686, \asqrt[53] , n_6445);
  and g15824 (n9690, n_6123, n_6122);
  and g15825 (n9691, \asqrt[25] , n9690);
  not g15826 (n_6446, n9691);
  and g15827 (n9692, n_6121, n_6446);
  not g15828 (n_6447, n9689);
  not g15829 (n_6448, n9692);
  and g15830 (n9693, n_6447, n_6448);
  and g15831 (n9694, n_722, n_6443);
  and g15832 (n9695, n_6444, n9694);
  not g15833 (n_6449, n9693);
  not g15834 (n_6450, n9695);
  and g15835 (n9696, n_6449, n_6450);
  not g15836 (n_6451, n9686);
  not g15837 (n_6452, n9696);
  and g15838 (n9697, n_6451, n_6452);
  not g15839 (n_6453, n9697);
  and g15840 (n9698, \asqrt[54] , n_6453);
  and g15844 (n9702, n_6131, n_6130);
  and g15845 (n9703, \asqrt[25] , n9702);
  not g15846 (n_6454, n9703);
  and g15847 (n9704, n_6129, n_6454);
  not g15848 (n_6455, n9701);
  not g15849 (n_6456, n9704);
  and g15850 (n9705, n_6455, n_6456);
  and g15851 (n9706, n_618, n_6451);
  and g15852 (n9707, n_6452, n9706);
  not g15853 (n_6457, n9705);
  not g15854 (n_6458, n9707);
  and g15855 (n9708, n_6457, n_6458);
  not g15856 (n_6459, n9698);
  not g15857 (n_6460, n9708);
  and g15858 (n9709, n_6459, n_6460);
  not g15859 (n_6461, n9709);
  and g15860 (n9710, \asqrt[55] , n_6461);
  and g15864 (n9714, n_6139, n_6138);
  and g15865 (n9715, \asqrt[25] , n9714);
  not g15866 (n_6462, n9715);
  and g15867 (n9716, n_6137, n_6462);
  not g15868 (n_6463, n9713);
  not g15869 (n_6464, n9716);
  and g15870 (n9717, n_6463, n_6464);
  and g15871 (n9718, n_522, n_6459);
  and g15872 (n9719, n_6460, n9718);
  not g15873 (n_6465, n9717);
  not g15874 (n_6466, n9719);
  and g15875 (n9720, n_6465, n_6466);
  not g15876 (n_6467, n9710);
  not g15877 (n_6468, n9720);
  and g15878 (n9721, n_6467, n_6468);
  not g15879 (n_6469, n9721);
  and g15880 (n9722, \asqrt[56] , n_6469);
  and g15884 (n9726, n_6147, n_6146);
  and g15885 (n9727, \asqrt[25] , n9726);
  not g15886 (n_6470, n9727);
  and g15887 (n9728, n_6145, n_6470);
  not g15888 (n_6471, n9725);
  not g15889 (n_6472, n9728);
  and g15890 (n9729, n_6471, n_6472);
  and g15891 (n9730, n_434, n_6467);
  and g15892 (n9731, n_6468, n9730);
  not g15893 (n_6473, n9729);
  not g15894 (n_6474, n9731);
  and g15895 (n9732, n_6473, n_6474);
  not g15896 (n_6475, n9722);
  not g15897 (n_6476, n9732);
  and g15898 (n9733, n_6475, n_6476);
  not g15899 (n_6477, n9733);
  and g15900 (n9734, \asqrt[57] , n_6477);
  and g15904 (n9738, n_6155, n_6154);
  and g15905 (n9739, \asqrt[25] , n9738);
  not g15906 (n_6478, n9739);
  and g15907 (n9740, n_6153, n_6478);
  not g15908 (n_6479, n9737);
  not g15909 (n_6480, n9740);
  and g15910 (n9741, n_6479, n_6480);
  and g15911 (n9742, n_354, n_6475);
  and g15912 (n9743, n_6476, n9742);
  not g15913 (n_6481, n9741);
  not g15914 (n_6482, n9743);
  and g15915 (n9744, n_6481, n_6482);
  not g15916 (n_6483, n9734);
  not g15917 (n_6484, n9744);
  and g15918 (n9745, n_6483, n_6484);
  not g15919 (n_6485, n9745);
  and g15920 (n9746, \asqrt[58] , n_6485);
  and g15924 (n9750, n_6163, n_6162);
  and g15925 (n9751, \asqrt[25] , n9750);
  not g15926 (n_6486, n9751);
  and g15927 (n9752, n_6161, n_6486);
  not g15928 (n_6487, n9749);
  not g15929 (n_6488, n9752);
  and g15930 (n9753, n_6487, n_6488);
  and g15931 (n9754, n_282, n_6483);
  and g15932 (n9755, n_6484, n9754);
  not g15933 (n_6489, n9753);
  not g15934 (n_6490, n9755);
  and g15935 (n9756, n_6489, n_6490);
  not g15936 (n_6491, n9746);
  not g15937 (n_6492, n9756);
  and g15938 (n9757, n_6491, n_6492);
  not g15939 (n_6493, n9757);
  and g15940 (n9758, \asqrt[59] , n_6493);
  and g15944 (n9762, n_6171, n_6170);
  and g15945 (n9763, \asqrt[25] , n9762);
  not g15946 (n_6494, n9763);
  and g15947 (n9764, n_6169, n_6494);
  not g15948 (n_6495, n9761);
  not g15949 (n_6496, n9764);
  and g15950 (n9765, n_6495, n_6496);
  and g15951 (n9766, n_218, n_6491);
  and g15952 (n9767, n_6492, n9766);
  not g15953 (n_6497, n9765);
  not g15954 (n_6498, n9767);
  and g15955 (n9768, n_6497, n_6498);
  not g15956 (n_6499, n9758);
  not g15957 (n_6500, n9768);
  and g15958 (n9769, n_6499, n_6500);
  not g15959 (n_6501, n9769);
  and g15960 (n9770, \asqrt[60] , n_6501);
  and g15964 (n9774, n_6179, n_6178);
  and g15965 (n9775, \asqrt[25] , n9774);
  not g15966 (n_6502, n9775);
  and g15967 (n9776, n_6177, n_6502);
  not g15968 (n_6503, n9773);
  not g15969 (n_6504, n9776);
  and g15970 (n9777, n_6503, n_6504);
  and g15971 (n9778, n_162, n_6499);
  and g15972 (n9779, n_6500, n9778);
  not g15973 (n_6505, n9777);
  not g15974 (n_6506, n9779);
  and g15975 (n9780, n_6505, n_6506);
  not g15976 (n_6507, n9770);
  not g15977 (n_6508, n9780);
  and g15978 (n9781, n_6507, n_6508);
  not g15979 (n_6509, n9781);
  and g15980 (n9782, \asqrt[61] , n_6509);
  and g15984 (n9786, n_6187, n_6186);
  and g15985 (n9787, \asqrt[25] , n9786);
  not g15986 (n_6510, n9787);
  and g15987 (n9788, n_6185, n_6510);
  not g15988 (n_6511, n9785);
  not g15989 (n_6512, n9788);
  and g15990 (n9789, n_6511, n_6512);
  and g15991 (n9790, n_115, n_6507);
  and g15992 (n9791, n_6508, n9790);
  not g15993 (n_6513, n9789);
  not g15994 (n_6514, n9791);
  and g15995 (n9792, n_6513, n_6514);
  not g15996 (n_6515, n9782);
  not g15997 (n_6516, n9792);
  and g15998 (n9793, n_6515, n_6516);
  not g15999 (n_6517, n9793);
  and g16000 (n9794, \asqrt[62] , n_6517);
  and g16004 (n9798, n_6195, n_6194);
  and g16005 (n9799, \asqrt[25] , n9798);
  not g16006 (n_6518, n9799);
  and g16007 (n9800, n_6193, n_6518);
  not g16008 (n_6519, n9797);
  not g16009 (n_6520, n9800);
  and g16010 (n9801, n_6519, n_6520);
  and g16011 (n9802, n_76, n_6515);
  and g16012 (n9803, n_6516, n9802);
  not g16013 (n_6521, n9801);
  not g16014 (n_6522, n9803);
  and g16015 (n9804, n_6521, n_6522);
  not g16016 (n_6523, n9794);
  not g16017 (n_6524, n9804);
  and g16018 (n9805, n_6523, n_6524);
  and g16022 (n9809, n_6203, n_6202);
  and g16023 (n9810, \asqrt[25] , n9809);
  not g16024 (n_6525, n9810);
  and g16025 (n9811, n_6201, n_6525);
  not g16026 (n_6526, n9808);
  not g16027 (n_6527, n9811);
  and g16028 (n9812, n_6526, n_6527);
  and g16029 (n9813, n_6210, n_6209);
  and g16030 (n9814, \asqrt[25] , n9813);
  not g16033 (n_6529, n9812);
  not g16035 (n_6530, n9805);
  not g16037 (n_6531, n9817);
  and g16038 (n9818, n_21, n_6531);
  and g16039 (n9819, n_6523, n9812);
  and g16040 (n9820, n_6524, n9819);
  and g16041 (n9821, n_6209, \asqrt[25] );
  not g16042 (n_6532, n9821);
  and g16043 (n9822, n9329, n_6532);
  not g16044 (n_6533, n9813);
  and g16045 (n9823, \asqrt[63] , n_6533);
  not g16046 (n_6534, n9822);
  and g16047 (n9824, n_6534, n9823);
  not g16053 (n_6535, n9824);
  not g16054 (n_6536, n9829);
  not g16056 (n_6537, n9820);
  and g16060 (n9833, \a[48] , \asqrt[24] );
  not g16061 (n_6542, \a[46] );
  not g16062 (n_6543, \a[47] );
  and g16063 (n9834, n_6542, n_6543);
  and g16064 (n9835, n_6222, n9834);
  not g16065 (n_6544, n9833);
  not g16066 (n_6545, n9835);
  and g16067 (n9836, n_6544, n_6545);
  not g16068 (n_6546, n9836);
  and g16069 (n9837, \asqrt[25] , n_6546);
  and g16075 (n9843, n_6222, \asqrt[24] );
  not g16076 (n_6547, n9843);
  and g16077 (n9844, \a[49] , n_6547);
  and g16078 (n9845, n9358, \asqrt[24] );
  not g16079 (n_6548, n9844);
  not g16080 (n_6549, n9845);
  and g16081 (n9846, n_6548, n_6549);
  not g16082 (n_6550, n9842);
  and g16083 (n9847, n_6550, n9846);
  not g16084 (n_6551, n9837);
  not g16085 (n_6552, n9847);
  and g16086 (n9848, n_6551, n_6552);
  not g16087 (n_6553, n9848);
  and g16088 (n9849, \asqrt[26] , n_6553);
  not g16089 (n_6554, \asqrt[26] );
  and g16090 (n9850, n_6554, n_6551);
  and g16091 (n9851, n_6552, n9850);
  not g16095 (n_6555, n9818);
  not g16097 (n_6556, n9855);
  and g16098 (n9856, n_6549, n_6556);
  not g16099 (n_6557, n9856);
  and g16100 (n9857, \a[50] , n_6557);
  and g16101 (n9858, n_5910, n_6556);
  and g16102 (n9859, n_6549, n9858);
  not g16103 (n_6558, n9857);
  not g16104 (n_6559, n9859);
  and g16105 (n9860, n_6558, n_6559);
  not g16106 (n_6560, n9851);
  not g16107 (n_6561, n9860);
  and g16108 (n9861, n_6560, n_6561);
  not g16109 (n_6562, n9849);
  not g16110 (n_6563, n9861);
  and g16111 (n9862, n_6562, n_6563);
  not g16112 (n_6564, n9862);
  and g16113 (n9863, \asqrt[27] , n_6564);
  and g16114 (n9864, n_6231, n_6230);
  not g16115 (n_6565, n9370);
  and g16116 (n9865, n_6565, n9864);
  and g16117 (n9866, \asqrt[24] , n9865);
  and g16118 (n9867, \asqrt[24] , n9864);
  not g16119 (n_6566, n9867);
  and g16120 (n9868, n9370, n_6566);
  not g16121 (n_6567, n9866);
  not g16122 (n_6568, n9868);
  and g16123 (n9869, n_6567, n_6568);
  and g16124 (n9870, n_6234, n_6562);
  and g16125 (n9871, n_6563, n9870);
  not g16126 (n_6569, n9869);
  not g16127 (n_6570, n9871);
  and g16128 (n9872, n_6569, n_6570);
  not g16129 (n_6571, n9863);
  not g16130 (n_6572, n9872);
  and g16131 (n9873, n_6571, n_6572);
  not g16132 (n_6573, n9873);
  and g16133 (n9874, \asqrt[28] , n_6573);
  and g16137 (n9878, n_6242, n_6240);
  and g16138 (n9879, \asqrt[24] , n9878);
  not g16139 (n_6574, n9879);
  and g16140 (n9880, n_6241, n_6574);
  not g16141 (n_6575, n9877);
  not g16142 (n_6576, n9880);
  and g16143 (n9881, n_6575, n_6576);
  and g16144 (n9882, n_5922, n_6571);
  and g16145 (n9883, n_6572, n9882);
  not g16146 (n_6577, n9881);
  not g16147 (n_6578, n9883);
  and g16148 (n9884, n_6577, n_6578);
  not g16149 (n_6579, n9874);
  not g16150 (n_6580, n9884);
  and g16151 (n9885, n_6579, n_6580);
  not g16152 (n_6581, n9885);
  and g16153 (n9886, \asqrt[29] , n_6581);
  and g16157 (n9890, n_6251, n_6250);
  and g16158 (n9891, \asqrt[24] , n9890);
  not g16159 (n_6582, n9891);
  and g16160 (n9892, n_6249, n_6582);
  not g16161 (n_6583, n9889);
  not g16162 (n_6584, n9892);
  and g16163 (n9893, n_6583, n_6584);
  and g16164 (n9894, n_5618, n_6579);
  and g16165 (n9895, n_6580, n9894);
  not g16166 (n_6585, n9893);
  not g16167 (n_6586, n9895);
  and g16168 (n9896, n_6585, n_6586);
  not g16169 (n_6587, n9886);
  not g16170 (n_6588, n9896);
  and g16171 (n9897, n_6587, n_6588);
  not g16172 (n_6589, n9897);
  and g16173 (n9898, \asqrt[30] , n_6589);
  and g16177 (n9902, n_6259, n_6258);
  and g16178 (n9903, \asqrt[24] , n9902);
  not g16179 (n_6590, n9903);
  and g16180 (n9904, n_6257, n_6590);
  not g16181 (n_6591, n9901);
  not g16182 (n_6592, n9904);
  and g16183 (n9905, n_6591, n_6592);
  and g16184 (n9906, n_5322, n_6587);
  and g16185 (n9907, n_6588, n9906);
  not g16186 (n_6593, n9905);
  not g16187 (n_6594, n9907);
  and g16188 (n9908, n_6593, n_6594);
  not g16189 (n_6595, n9898);
  not g16190 (n_6596, n9908);
  and g16191 (n9909, n_6595, n_6596);
  not g16192 (n_6597, n9909);
  and g16193 (n9910, \asqrt[31] , n_6597);
  and g16197 (n9914, n_6267, n_6266);
  and g16198 (n9915, \asqrt[24] , n9914);
  not g16199 (n_6598, n9915);
  and g16200 (n9916, n_6265, n_6598);
  not g16201 (n_6599, n9913);
  not g16202 (n_6600, n9916);
  and g16203 (n9917, n_6599, n_6600);
  and g16204 (n9918, n_5034, n_6595);
  and g16205 (n9919, n_6596, n9918);
  not g16206 (n_6601, n9917);
  not g16207 (n_6602, n9919);
  and g16208 (n9920, n_6601, n_6602);
  not g16209 (n_6603, n9910);
  not g16210 (n_6604, n9920);
  and g16211 (n9921, n_6603, n_6604);
  not g16212 (n_6605, n9921);
  and g16213 (n9922, \asqrt[32] , n_6605);
  and g16217 (n9926, n_6275, n_6274);
  and g16218 (n9927, \asqrt[24] , n9926);
  not g16219 (n_6606, n9927);
  and g16220 (n9928, n_6273, n_6606);
  not g16221 (n_6607, n9925);
  not g16222 (n_6608, n9928);
  and g16223 (n9929, n_6607, n_6608);
  and g16224 (n9930, n_4754, n_6603);
  and g16225 (n9931, n_6604, n9930);
  not g16226 (n_6609, n9929);
  not g16227 (n_6610, n9931);
  and g16228 (n9932, n_6609, n_6610);
  not g16229 (n_6611, n9922);
  not g16230 (n_6612, n9932);
  and g16231 (n9933, n_6611, n_6612);
  not g16232 (n_6613, n9933);
  and g16233 (n9934, \asqrt[33] , n_6613);
  and g16237 (n9938, n_6283, n_6282);
  and g16238 (n9939, \asqrt[24] , n9938);
  not g16239 (n_6614, n9939);
  and g16240 (n9940, n_6281, n_6614);
  not g16241 (n_6615, n9937);
  not g16242 (n_6616, n9940);
  and g16243 (n9941, n_6615, n_6616);
  and g16244 (n9942, n_4482, n_6611);
  and g16245 (n9943, n_6612, n9942);
  not g16246 (n_6617, n9941);
  not g16247 (n_6618, n9943);
  and g16248 (n9944, n_6617, n_6618);
  not g16249 (n_6619, n9934);
  not g16250 (n_6620, n9944);
  and g16251 (n9945, n_6619, n_6620);
  not g16252 (n_6621, n9945);
  and g16253 (n9946, \asqrt[34] , n_6621);
  and g16257 (n9950, n_6291, n_6290);
  and g16258 (n9951, \asqrt[24] , n9950);
  not g16259 (n_6622, n9951);
  and g16260 (n9952, n_6289, n_6622);
  not g16261 (n_6623, n9949);
  not g16262 (n_6624, n9952);
  and g16263 (n9953, n_6623, n_6624);
  and g16264 (n9954, n_4218, n_6619);
  and g16265 (n9955, n_6620, n9954);
  not g16266 (n_6625, n9953);
  not g16267 (n_6626, n9955);
  and g16268 (n9956, n_6625, n_6626);
  not g16269 (n_6627, n9946);
  not g16270 (n_6628, n9956);
  and g16271 (n9957, n_6627, n_6628);
  not g16272 (n_6629, n9957);
  and g16273 (n9958, \asqrt[35] , n_6629);
  and g16277 (n9962, n_6299, n_6298);
  and g16278 (n9963, \asqrt[24] , n9962);
  not g16279 (n_6630, n9963);
  and g16280 (n9964, n_6297, n_6630);
  not g16281 (n_6631, n9961);
  not g16282 (n_6632, n9964);
  and g16283 (n9965, n_6631, n_6632);
  and g16284 (n9966, n_3962, n_6627);
  and g16285 (n9967, n_6628, n9966);
  not g16286 (n_6633, n9965);
  not g16287 (n_6634, n9967);
  and g16288 (n9968, n_6633, n_6634);
  not g16289 (n_6635, n9958);
  not g16290 (n_6636, n9968);
  and g16291 (n9969, n_6635, n_6636);
  not g16292 (n_6637, n9969);
  and g16293 (n9970, \asqrt[36] , n_6637);
  and g16297 (n9974, n_6307, n_6306);
  and g16298 (n9975, \asqrt[24] , n9974);
  not g16299 (n_6638, n9975);
  and g16300 (n9976, n_6305, n_6638);
  not g16301 (n_6639, n9973);
  not g16302 (n_6640, n9976);
  and g16303 (n9977, n_6639, n_6640);
  and g16304 (n9978, n_3714, n_6635);
  and g16305 (n9979, n_6636, n9978);
  not g16306 (n_6641, n9977);
  not g16307 (n_6642, n9979);
  and g16308 (n9980, n_6641, n_6642);
  not g16309 (n_6643, n9970);
  not g16310 (n_6644, n9980);
  and g16311 (n9981, n_6643, n_6644);
  not g16312 (n_6645, n9981);
  and g16313 (n9982, \asqrt[37] , n_6645);
  and g16317 (n9986, n_6315, n_6314);
  and g16318 (n9987, \asqrt[24] , n9986);
  not g16319 (n_6646, n9987);
  and g16320 (n9988, n_6313, n_6646);
  not g16321 (n_6647, n9985);
  not g16322 (n_6648, n9988);
  and g16323 (n9989, n_6647, n_6648);
  and g16324 (n9990, n_3474, n_6643);
  and g16325 (n9991, n_6644, n9990);
  not g16326 (n_6649, n9989);
  not g16327 (n_6650, n9991);
  and g16328 (n9992, n_6649, n_6650);
  not g16329 (n_6651, n9982);
  not g16330 (n_6652, n9992);
  and g16331 (n9993, n_6651, n_6652);
  not g16332 (n_6653, n9993);
  and g16333 (n9994, \asqrt[38] , n_6653);
  and g16337 (n9998, n_6323, n_6322);
  and g16338 (n9999, \asqrt[24] , n9998);
  not g16339 (n_6654, n9999);
  and g16340 (n10000, n_6321, n_6654);
  not g16341 (n_6655, n9997);
  not g16342 (n_6656, n10000);
  and g16343 (n10001, n_6655, n_6656);
  and g16344 (n10002, n_3242, n_6651);
  and g16345 (n10003, n_6652, n10002);
  not g16346 (n_6657, n10001);
  not g16347 (n_6658, n10003);
  and g16348 (n10004, n_6657, n_6658);
  not g16349 (n_6659, n9994);
  not g16350 (n_6660, n10004);
  and g16351 (n10005, n_6659, n_6660);
  not g16352 (n_6661, n10005);
  and g16353 (n10006, \asqrt[39] , n_6661);
  and g16357 (n10010, n_6331, n_6330);
  and g16358 (n10011, \asqrt[24] , n10010);
  not g16359 (n_6662, n10011);
  and g16360 (n10012, n_6329, n_6662);
  not g16361 (n_6663, n10009);
  not g16362 (n_6664, n10012);
  and g16363 (n10013, n_6663, n_6664);
  and g16364 (n10014, n_3018, n_6659);
  and g16365 (n10015, n_6660, n10014);
  not g16366 (n_6665, n10013);
  not g16367 (n_6666, n10015);
  and g16368 (n10016, n_6665, n_6666);
  not g16369 (n_6667, n10006);
  not g16370 (n_6668, n10016);
  and g16371 (n10017, n_6667, n_6668);
  not g16372 (n_6669, n10017);
  and g16373 (n10018, \asqrt[40] , n_6669);
  and g16377 (n10022, n_6339, n_6338);
  and g16378 (n10023, \asqrt[24] , n10022);
  not g16379 (n_6670, n10023);
  and g16380 (n10024, n_6337, n_6670);
  not g16381 (n_6671, n10021);
  not g16382 (n_6672, n10024);
  and g16383 (n10025, n_6671, n_6672);
  and g16384 (n10026, n_2802, n_6667);
  and g16385 (n10027, n_6668, n10026);
  not g16386 (n_6673, n10025);
  not g16387 (n_6674, n10027);
  and g16388 (n10028, n_6673, n_6674);
  not g16389 (n_6675, n10018);
  not g16390 (n_6676, n10028);
  and g16391 (n10029, n_6675, n_6676);
  not g16392 (n_6677, n10029);
  and g16393 (n10030, \asqrt[41] , n_6677);
  and g16394 (n10031, n_2594, n_6675);
  and g16395 (n10032, n_6676, n10031);
  and g16399 (n10036, n_6347, n_6345);
  and g16400 (n10037, \asqrt[24] , n10036);
  not g16401 (n_6678, n10037);
  and g16402 (n10038, n_6346, n_6678);
  not g16403 (n_6679, n10035);
  not g16404 (n_6680, n10038);
  and g16405 (n10039, n_6679, n_6680);
  not g16406 (n_6681, n10032);
  not g16407 (n_6682, n10039);
  and g16408 (n10040, n_6681, n_6682);
  not g16409 (n_6683, n10030);
  not g16410 (n_6684, n10040);
  and g16411 (n10041, n_6683, n_6684);
  not g16412 (n_6685, n10041);
  and g16413 (n10042, \asqrt[42] , n_6685);
  and g16417 (n10046, n_6355, n_6354);
  and g16418 (n10047, \asqrt[24] , n10046);
  not g16419 (n_6686, n10047);
  and g16420 (n10048, n_6353, n_6686);
  not g16421 (n_6687, n10045);
  not g16422 (n_6688, n10048);
  and g16423 (n10049, n_6687, n_6688);
  and g16424 (n10050, n_2394, n_6683);
  and g16425 (n10051, n_6684, n10050);
  not g16426 (n_6689, n10049);
  not g16427 (n_6690, n10051);
  and g16428 (n10052, n_6689, n_6690);
  not g16429 (n_6691, n10042);
  not g16430 (n_6692, n10052);
  and g16431 (n10053, n_6691, n_6692);
  not g16432 (n_6693, n10053);
  and g16433 (n10054, \asqrt[43] , n_6693);
  and g16437 (n10058, n_6363, n_6362);
  and g16438 (n10059, \asqrt[24] , n10058);
  not g16439 (n_6694, n10059);
  and g16440 (n10060, n_6361, n_6694);
  not g16441 (n_6695, n10057);
  not g16442 (n_6696, n10060);
  and g16443 (n10061, n_6695, n_6696);
  and g16444 (n10062, n_2202, n_6691);
  and g16445 (n10063, n_6692, n10062);
  not g16446 (n_6697, n10061);
  not g16447 (n_6698, n10063);
  and g16448 (n10064, n_6697, n_6698);
  not g16449 (n_6699, n10054);
  not g16450 (n_6700, n10064);
  and g16451 (n10065, n_6699, n_6700);
  not g16452 (n_6701, n10065);
  and g16453 (n10066, \asqrt[44] , n_6701);
  and g16457 (n10070, n_6371, n_6370);
  and g16458 (n10071, \asqrt[24] , n10070);
  not g16459 (n_6702, n10071);
  and g16460 (n10072, n_6369, n_6702);
  not g16461 (n_6703, n10069);
  not g16462 (n_6704, n10072);
  and g16463 (n10073, n_6703, n_6704);
  and g16464 (n10074, n_2018, n_6699);
  and g16465 (n10075, n_6700, n10074);
  not g16466 (n_6705, n10073);
  not g16467 (n_6706, n10075);
  and g16468 (n10076, n_6705, n_6706);
  not g16469 (n_6707, n10066);
  not g16470 (n_6708, n10076);
  and g16471 (n10077, n_6707, n_6708);
  not g16472 (n_6709, n10077);
  and g16473 (n10078, \asqrt[45] , n_6709);
  and g16477 (n10082, n_6379, n_6378);
  and g16478 (n10083, \asqrt[24] , n10082);
  not g16479 (n_6710, n10083);
  and g16480 (n10084, n_6377, n_6710);
  not g16481 (n_6711, n10081);
  not g16482 (n_6712, n10084);
  and g16483 (n10085, n_6711, n_6712);
  and g16484 (n10086, n_1842, n_6707);
  and g16485 (n10087, n_6708, n10086);
  not g16486 (n_6713, n10085);
  not g16487 (n_6714, n10087);
  and g16488 (n10088, n_6713, n_6714);
  not g16489 (n_6715, n10078);
  not g16490 (n_6716, n10088);
  and g16491 (n10089, n_6715, n_6716);
  not g16492 (n_6717, n10089);
  and g16493 (n10090, \asqrt[46] , n_6717);
  and g16497 (n10094, n_6387, n_6386);
  and g16498 (n10095, \asqrt[24] , n10094);
  not g16499 (n_6718, n10095);
  and g16500 (n10096, n_6385, n_6718);
  not g16501 (n_6719, n10093);
  not g16502 (n_6720, n10096);
  and g16503 (n10097, n_6719, n_6720);
  and g16504 (n10098, n_1674, n_6715);
  and g16505 (n10099, n_6716, n10098);
  not g16506 (n_6721, n10097);
  not g16507 (n_6722, n10099);
  and g16508 (n10100, n_6721, n_6722);
  not g16509 (n_6723, n10090);
  not g16510 (n_6724, n10100);
  and g16511 (n10101, n_6723, n_6724);
  not g16512 (n_6725, n10101);
  and g16513 (n10102, \asqrt[47] , n_6725);
  and g16517 (n10106, n_6395, n_6394);
  and g16518 (n10107, \asqrt[24] , n10106);
  not g16519 (n_6726, n10107);
  and g16520 (n10108, n_6393, n_6726);
  not g16521 (n_6727, n10105);
  not g16522 (n_6728, n10108);
  and g16523 (n10109, n_6727, n_6728);
  and g16524 (n10110, n_1514, n_6723);
  and g16525 (n10111, n_6724, n10110);
  not g16526 (n_6729, n10109);
  not g16527 (n_6730, n10111);
  and g16528 (n10112, n_6729, n_6730);
  not g16529 (n_6731, n10102);
  not g16530 (n_6732, n10112);
  and g16531 (n10113, n_6731, n_6732);
  not g16532 (n_6733, n10113);
  and g16533 (n10114, \asqrt[48] , n_6733);
  and g16537 (n10118, n_6403, n_6402);
  and g16538 (n10119, \asqrt[24] , n10118);
  not g16539 (n_6734, n10119);
  and g16540 (n10120, n_6401, n_6734);
  not g16541 (n_6735, n10117);
  not g16542 (n_6736, n10120);
  and g16543 (n10121, n_6735, n_6736);
  and g16544 (n10122, n_1362, n_6731);
  and g16545 (n10123, n_6732, n10122);
  not g16546 (n_6737, n10121);
  not g16547 (n_6738, n10123);
  and g16548 (n10124, n_6737, n_6738);
  not g16549 (n_6739, n10114);
  not g16550 (n_6740, n10124);
  and g16551 (n10125, n_6739, n_6740);
  not g16552 (n_6741, n10125);
  and g16553 (n10126, \asqrt[49] , n_6741);
  and g16557 (n10130, n_6411, n_6410);
  and g16558 (n10131, \asqrt[24] , n10130);
  not g16559 (n_6742, n10131);
  and g16560 (n10132, n_6409, n_6742);
  not g16561 (n_6743, n10129);
  not g16562 (n_6744, n10132);
  and g16563 (n10133, n_6743, n_6744);
  and g16564 (n10134, n_1218, n_6739);
  and g16565 (n10135, n_6740, n10134);
  not g16566 (n_6745, n10133);
  not g16567 (n_6746, n10135);
  and g16568 (n10136, n_6745, n_6746);
  not g16569 (n_6747, n10126);
  not g16570 (n_6748, n10136);
  and g16571 (n10137, n_6747, n_6748);
  not g16572 (n_6749, n10137);
  and g16573 (n10138, \asqrt[50] , n_6749);
  and g16577 (n10142, n_6419, n_6418);
  and g16578 (n10143, \asqrt[24] , n10142);
  not g16579 (n_6750, n10143);
  and g16580 (n10144, n_6417, n_6750);
  not g16581 (n_6751, n10141);
  not g16582 (n_6752, n10144);
  and g16583 (n10145, n_6751, n_6752);
  and g16584 (n10146, n_1082, n_6747);
  and g16585 (n10147, n_6748, n10146);
  not g16586 (n_6753, n10145);
  not g16587 (n_6754, n10147);
  and g16588 (n10148, n_6753, n_6754);
  not g16589 (n_6755, n10138);
  not g16590 (n_6756, n10148);
  and g16591 (n10149, n_6755, n_6756);
  not g16592 (n_6757, n10149);
  and g16593 (n10150, \asqrt[51] , n_6757);
  and g16597 (n10154, n_6427, n_6426);
  and g16598 (n10155, \asqrt[24] , n10154);
  not g16599 (n_6758, n10155);
  and g16600 (n10156, n_6425, n_6758);
  not g16601 (n_6759, n10153);
  not g16602 (n_6760, n10156);
  and g16603 (n10157, n_6759, n_6760);
  and g16604 (n10158, n_954, n_6755);
  and g16605 (n10159, n_6756, n10158);
  not g16606 (n_6761, n10157);
  not g16607 (n_6762, n10159);
  and g16608 (n10160, n_6761, n_6762);
  not g16609 (n_6763, n10150);
  not g16610 (n_6764, n10160);
  and g16611 (n10161, n_6763, n_6764);
  not g16612 (n_6765, n10161);
  and g16613 (n10162, \asqrt[52] , n_6765);
  and g16617 (n10166, n_6435, n_6434);
  and g16618 (n10167, \asqrt[24] , n10166);
  not g16619 (n_6766, n10167);
  and g16620 (n10168, n_6433, n_6766);
  not g16621 (n_6767, n10165);
  not g16622 (n_6768, n10168);
  and g16623 (n10169, n_6767, n_6768);
  and g16624 (n10170, n_834, n_6763);
  and g16625 (n10171, n_6764, n10170);
  not g16626 (n_6769, n10169);
  not g16627 (n_6770, n10171);
  and g16628 (n10172, n_6769, n_6770);
  not g16629 (n_6771, n10162);
  not g16630 (n_6772, n10172);
  and g16631 (n10173, n_6771, n_6772);
  not g16632 (n_6773, n10173);
  and g16633 (n10174, \asqrt[53] , n_6773);
  and g16637 (n10178, n_6443, n_6442);
  and g16638 (n10179, \asqrt[24] , n10178);
  not g16639 (n_6774, n10179);
  and g16640 (n10180, n_6441, n_6774);
  not g16641 (n_6775, n10177);
  not g16642 (n_6776, n10180);
  and g16643 (n10181, n_6775, n_6776);
  and g16644 (n10182, n_722, n_6771);
  and g16645 (n10183, n_6772, n10182);
  not g16646 (n_6777, n10181);
  not g16647 (n_6778, n10183);
  and g16648 (n10184, n_6777, n_6778);
  not g16649 (n_6779, n10174);
  not g16650 (n_6780, n10184);
  and g16651 (n10185, n_6779, n_6780);
  not g16652 (n_6781, n10185);
  and g16653 (n10186, \asqrt[54] , n_6781);
  and g16657 (n10190, n_6451, n_6450);
  and g16658 (n10191, \asqrt[24] , n10190);
  not g16659 (n_6782, n10191);
  and g16660 (n10192, n_6449, n_6782);
  not g16661 (n_6783, n10189);
  not g16662 (n_6784, n10192);
  and g16663 (n10193, n_6783, n_6784);
  and g16664 (n10194, n_618, n_6779);
  and g16665 (n10195, n_6780, n10194);
  not g16666 (n_6785, n10193);
  not g16667 (n_6786, n10195);
  and g16668 (n10196, n_6785, n_6786);
  not g16669 (n_6787, n10186);
  not g16670 (n_6788, n10196);
  and g16671 (n10197, n_6787, n_6788);
  not g16672 (n_6789, n10197);
  and g16673 (n10198, \asqrt[55] , n_6789);
  and g16677 (n10202, n_6459, n_6458);
  and g16678 (n10203, \asqrt[24] , n10202);
  not g16679 (n_6790, n10203);
  and g16680 (n10204, n_6457, n_6790);
  not g16681 (n_6791, n10201);
  not g16682 (n_6792, n10204);
  and g16683 (n10205, n_6791, n_6792);
  and g16684 (n10206, n_522, n_6787);
  and g16685 (n10207, n_6788, n10206);
  not g16686 (n_6793, n10205);
  not g16687 (n_6794, n10207);
  and g16688 (n10208, n_6793, n_6794);
  not g16689 (n_6795, n10198);
  not g16690 (n_6796, n10208);
  and g16691 (n10209, n_6795, n_6796);
  not g16692 (n_6797, n10209);
  and g16693 (n10210, \asqrt[56] , n_6797);
  and g16697 (n10214, n_6467, n_6466);
  and g16698 (n10215, \asqrt[24] , n10214);
  not g16699 (n_6798, n10215);
  and g16700 (n10216, n_6465, n_6798);
  not g16701 (n_6799, n10213);
  not g16702 (n_6800, n10216);
  and g16703 (n10217, n_6799, n_6800);
  and g16704 (n10218, n_434, n_6795);
  and g16705 (n10219, n_6796, n10218);
  not g16706 (n_6801, n10217);
  not g16707 (n_6802, n10219);
  and g16708 (n10220, n_6801, n_6802);
  not g16709 (n_6803, n10210);
  not g16710 (n_6804, n10220);
  and g16711 (n10221, n_6803, n_6804);
  not g16712 (n_6805, n10221);
  and g16713 (n10222, \asqrt[57] , n_6805);
  and g16717 (n10226, n_6475, n_6474);
  and g16718 (n10227, \asqrt[24] , n10226);
  not g16719 (n_6806, n10227);
  and g16720 (n10228, n_6473, n_6806);
  not g16721 (n_6807, n10225);
  not g16722 (n_6808, n10228);
  and g16723 (n10229, n_6807, n_6808);
  and g16724 (n10230, n_354, n_6803);
  and g16725 (n10231, n_6804, n10230);
  not g16726 (n_6809, n10229);
  not g16727 (n_6810, n10231);
  and g16728 (n10232, n_6809, n_6810);
  not g16729 (n_6811, n10222);
  not g16730 (n_6812, n10232);
  and g16731 (n10233, n_6811, n_6812);
  not g16732 (n_6813, n10233);
  and g16733 (n10234, \asqrt[58] , n_6813);
  and g16737 (n10238, n_6483, n_6482);
  and g16738 (n10239, \asqrt[24] , n10238);
  not g16739 (n_6814, n10239);
  and g16740 (n10240, n_6481, n_6814);
  not g16741 (n_6815, n10237);
  not g16742 (n_6816, n10240);
  and g16743 (n10241, n_6815, n_6816);
  and g16744 (n10242, n_282, n_6811);
  and g16745 (n10243, n_6812, n10242);
  not g16746 (n_6817, n10241);
  not g16747 (n_6818, n10243);
  and g16748 (n10244, n_6817, n_6818);
  not g16749 (n_6819, n10234);
  not g16750 (n_6820, n10244);
  and g16751 (n10245, n_6819, n_6820);
  not g16752 (n_6821, n10245);
  and g16753 (n10246, \asqrt[59] , n_6821);
  and g16757 (n10250, n_6491, n_6490);
  and g16758 (n10251, \asqrt[24] , n10250);
  not g16759 (n_6822, n10251);
  and g16760 (n10252, n_6489, n_6822);
  not g16761 (n_6823, n10249);
  not g16762 (n_6824, n10252);
  and g16763 (n10253, n_6823, n_6824);
  and g16764 (n10254, n_218, n_6819);
  and g16765 (n10255, n_6820, n10254);
  not g16766 (n_6825, n10253);
  not g16767 (n_6826, n10255);
  and g16768 (n10256, n_6825, n_6826);
  not g16769 (n_6827, n10246);
  not g16770 (n_6828, n10256);
  and g16771 (n10257, n_6827, n_6828);
  not g16772 (n_6829, n10257);
  and g16773 (n10258, \asqrt[60] , n_6829);
  and g16777 (n10262, n_6499, n_6498);
  and g16778 (n10263, \asqrt[24] , n10262);
  not g16779 (n_6830, n10263);
  and g16780 (n10264, n_6497, n_6830);
  not g16781 (n_6831, n10261);
  not g16782 (n_6832, n10264);
  and g16783 (n10265, n_6831, n_6832);
  and g16784 (n10266, n_162, n_6827);
  and g16785 (n10267, n_6828, n10266);
  not g16786 (n_6833, n10265);
  not g16787 (n_6834, n10267);
  and g16788 (n10268, n_6833, n_6834);
  not g16789 (n_6835, n10258);
  not g16790 (n_6836, n10268);
  and g16791 (n10269, n_6835, n_6836);
  not g16792 (n_6837, n10269);
  and g16793 (n10270, \asqrt[61] , n_6837);
  and g16797 (n10274, n_6507, n_6506);
  and g16798 (n10275, \asqrt[24] , n10274);
  not g16799 (n_6838, n10275);
  and g16800 (n10276, n_6505, n_6838);
  not g16801 (n_6839, n10273);
  not g16802 (n_6840, n10276);
  and g16803 (n10277, n_6839, n_6840);
  and g16804 (n10278, n_115, n_6835);
  and g16805 (n10279, n_6836, n10278);
  not g16806 (n_6841, n10277);
  not g16807 (n_6842, n10279);
  and g16808 (n10280, n_6841, n_6842);
  not g16809 (n_6843, n10270);
  not g16810 (n_6844, n10280);
  and g16811 (n10281, n_6843, n_6844);
  not g16812 (n_6845, n10281);
  and g16813 (n10282, \asqrt[62] , n_6845);
  and g16817 (n10286, n_6515, n_6514);
  and g16818 (n10287, \asqrt[24] , n10286);
  not g16819 (n_6846, n10287);
  and g16820 (n10288, n_6513, n_6846);
  not g16821 (n_6847, n10285);
  not g16822 (n_6848, n10288);
  and g16823 (n10289, n_6847, n_6848);
  and g16824 (n10290, n_76, n_6843);
  and g16825 (n10291, n_6844, n10290);
  not g16826 (n_6849, n10289);
  not g16827 (n_6850, n10291);
  and g16828 (n10292, n_6849, n_6850);
  not g16829 (n_6851, n10282);
  not g16830 (n_6852, n10292);
  and g16831 (n10293, n_6851, n_6852);
  and g16835 (n10297, n_6523, n_6522);
  and g16836 (n10298, \asqrt[24] , n10297);
  not g16837 (n_6853, n10298);
  and g16838 (n10299, n_6521, n_6853);
  not g16839 (n_6854, n10296);
  not g16840 (n_6855, n10299);
  and g16841 (n10300, n_6854, n_6855);
  and g16842 (n10301, n_6530, n_6529);
  and g16843 (n10302, \asqrt[24] , n10301);
  not g16846 (n_6857, n10300);
  not g16848 (n_6858, n10293);
  not g16850 (n_6859, n10305);
  and g16851 (n10306, n_21, n_6859);
  and g16852 (n10307, n_6851, n10300);
  and g16853 (n10308, n_6852, n10307);
  and g16854 (n10309, n_6529, \asqrt[24] );
  not g16855 (n_6860, n10309);
  and g16856 (n10310, n9805, n_6860);
  not g16857 (n_6861, n10301);
  and g16858 (n10311, \asqrt[63] , n_6861);
  not g16859 (n_6862, n10310);
  and g16860 (n10312, n_6862, n10311);
  not g16866 (n_6863, n10312);
  not g16867 (n_6864, n10317);
  not g16869 (n_6865, n10308);
  and g16873 (n10321, \a[46] , \asqrt[23] );
  not g16874 (n_6870, \a[44] );
  not g16875 (n_6871, \a[45] );
  and g16876 (n10322, n_6870, n_6871);
  and g16877 (n10323, n_6542, n10322);
  not g16878 (n_6872, n10321);
  not g16879 (n_6873, n10323);
  and g16880 (n10324, n_6872, n_6873);
  not g16881 (n_6874, n10324);
  and g16882 (n10325, \asqrt[24] , n_6874);
  and g16888 (n10331, n_6542, \asqrt[23] );
  not g16889 (n_6875, n10331);
  and g16890 (n10332, \a[47] , n_6875);
  and g16891 (n10333, n9834, \asqrt[23] );
  not g16892 (n_6876, n10332);
  not g16893 (n_6877, n10333);
  and g16894 (n10334, n_6876, n_6877);
  not g16895 (n_6878, n10330);
  and g16896 (n10335, n_6878, n10334);
  not g16897 (n_6879, n10325);
  not g16898 (n_6880, n10335);
  and g16899 (n10336, n_6879, n_6880);
  not g16900 (n_6881, n10336);
  and g16901 (n10337, \asqrt[25] , n_6881);
  not g16902 (n_6882, \asqrt[25] );
  and g16903 (n10338, n_6882, n_6879);
  and g16904 (n10339, n_6880, n10338);
  not g16908 (n_6883, n10306);
  not g16910 (n_6884, n10343);
  and g16911 (n10344, n_6877, n_6884);
  not g16912 (n_6885, n10344);
  and g16913 (n10345, \a[48] , n_6885);
  and g16914 (n10346, n_6222, n_6884);
  and g16915 (n10347, n_6877, n10346);
  not g16916 (n_6886, n10345);
  not g16917 (n_6887, n10347);
  and g16918 (n10348, n_6886, n_6887);
  not g16919 (n_6888, n10339);
  not g16920 (n_6889, n10348);
  and g16921 (n10349, n_6888, n_6889);
  not g16922 (n_6890, n10337);
  not g16923 (n_6891, n10349);
  and g16924 (n10350, n_6890, n_6891);
  not g16925 (n_6892, n10350);
  and g16926 (n10351, \asqrt[26] , n_6892);
  and g16927 (n10352, n_6551, n_6550);
  not g16928 (n_6893, n9846);
  and g16929 (n10353, n_6893, n10352);
  and g16930 (n10354, \asqrt[23] , n10353);
  and g16931 (n10355, \asqrt[23] , n10352);
  not g16932 (n_6894, n10355);
  and g16933 (n10356, n9846, n_6894);
  not g16934 (n_6895, n10354);
  not g16935 (n_6896, n10356);
  and g16936 (n10357, n_6895, n_6896);
  and g16937 (n10358, n_6554, n_6890);
  and g16938 (n10359, n_6891, n10358);
  not g16939 (n_6897, n10357);
  not g16940 (n_6898, n10359);
  and g16941 (n10360, n_6897, n_6898);
  not g16942 (n_6899, n10351);
  not g16943 (n_6900, n10360);
  and g16944 (n10361, n_6899, n_6900);
  not g16945 (n_6901, n10361);
  and g16946 (n10362, \asqrt[27] , n_6901);
  and g16950 (n10366, n_6562, n_6560);
  and g16951 (n10367, \asqrt[23] , n10366);
  not g16952 (n_6902, n10367);
  and g16953 (n10368, n_6561, n_6902);
  not g16954 (n_6903, n10365);
  not g16955 (n_6904, n10368);
  and g16956 (n10369, n_6903, n_6904);
  and g16957 (n10370, n_6234, n_6899);
  and g16958 (n10371, n_6900, n10370);
  not g16959 (n_6905, n10369);
  not g16960 (n_6906, n10371);
  and g16961 (n10372, n_6905, n_6906);
  not g16962 (n_6907, n10362);
  not g16963 (n_6908, n10372);
  and g16964 (n10373, n_6907, n_6908);
  not g16965 (n_6909, n10373);
  and g16966 (n10374, \asqrt[28] , n_6909);
  and g16970 (n10378, n_6571, n_6570);
  and g16971 (n10379, \asqrt[23] , n10378);
  not g16972 (n_6910, n10379);
  and g16973 (n10380, n_6569, n_6910);
  not g16974 (n_6911, n10377);
  not g16975 (n_6912, n10380);
  and g16976 (n10381, n_6911, n_6912);
  and g16977 (n10382, n_5922, n_6907);
  and g16978 (n10383, n_6908, n10382);
  not g16979 (n_6913, n10381);
  not g16980 (n_6914, n10383);
  and g16981 (n10384, n_6913, n_6914);
  not g16982 (n_6915, n10374);
  not g16983 (n_6916, n10384);
  and g16984 (n10385, n_6915, n_6916);
  not g16985 (n_6917, n10385);
  and g16986 (n10386, \asqrt[29] , n_6917);
  and g16990 (n10390, n_6579, n_6578);
  and g16991 (n10391, \asqrt[23] , n10390);
  not g16992 (n_6918, n10391);
  and g16993 (n10392, n_6577, n_6918);
  not g16994 (n_6919, n10389);
  not g16995 (n_6920, n10392);
  and g16996 (n10393, n_6919, n_6920);
  and g16997 (n10394, n_5618, n_6915);
  and g16998 (n10395, n_6916, n10394);
  not g16999 (n_6921, n10393);
  not g17000 (n_6922, n10395);
  and g17001 (n10396, n_6921, n_6922);
  not g17002 (n_6923, n10386);
  not g17003 (n_6924, n10396);
  and g17004 (n10397, n_6923, n_6924);
  not g17005 (n_6925, n10397);
  and g17006 (n10398, \asqrt[30] , n_6925);
  and g17010 (n10402, n_6587, n_6586);
  and g17011 (n10403, \asqrt[23] , n10402);
  not g17012 (n_6926, n10403);
  and g17013 (n10404, n_6585, n_6926);
  not g17014 (n_6927, n10401);
  not g17015 (n_6928, n10404);
  and g17016 (n10405, n_6927, n_6928);
  and g17017 (n10406, n_5322, n_6923);
  and g17018 (n10407, n_6924, n10406);
  not g17019 (n_6929, n10405);
  not g17020 (n_6930, n10407);
  and g17021 (n10408, n_6929, n_6930);
  not g17022 (n_6931, n10398);
  not g17023 (n_6932, n10408);
  and g17024 (n10409, n_6931, n_6932);
  not g17025 (n_6933, n10409);
  and g17026 (n10410, \asqrt[31] , n_6933);
  and g17030 (n10414, n_6595, n_6594);
  and g17031 (n10415, \asqrt[23] , n10414);
  not g17032 (n_6934, n10415);
  and g17033 (n10416, n_6593, n_6934);
  not g17034 (n_6935, n10413);
  not g17035 (n_6936, n10416);
  and g17036 (n10417, n_6935, n_6936);
  and g17037 (n10418, n_5034, n_6931);
  and g17038 (n10419, n_6932, n10418);
  not g17039 (n_6937, n10417);
  not g17040 (n_6938, n10419);
  and g17041 (n10420, n_6937, n_6938);
  not g17042 (n_6939, n10410);
  not g17043 (n_6940, n10420);
  and g17044 (n10421, n_6939, n_6940);
  not g17045 (n_6941, n10421);
  and g17046 (n10422, \asqrt[32] , n_6941);
  and g17050 (n10426, n_6603, n_6602);
  and g17051 (n10427, \asqrt[23] , n10426);
  not g17052 (n_6942, n10427);
  and g17053 (n10428, n_6601, n_6942);
  not g17054 (n_6943, n10425);
  not g17055 (n_6944, n10428);
  and g17056 (n10429, n_6943, n_6944);
  and g17057 (n10430, n_4754, n_6939);
  and g17058 (n10431, n_6940, n10430);
  not g17059 (n_6945, n10429);
  not g17060 (n_6946, n10431);
  and g17061 (n10432, n_6945, n_6946);
  not g17062 (n_6947, n10422);
  not g17063 (n_6948, n10432);
  and g17064 (n10433, n_6947, n_6948);
  not g17065 (n_6949, n10433);
  and g17066 (n10434, \asqrt[33] , n_6949);
  and g17070 (n10438, n_6611, n_6610);
  and g17071 (n10439, \asqrt[23] , n10438);
  not g17072 (n_6950, n10439);
  and g17073 (n10440, n_6609, n_6950);
  not g17074 (n_6951, n10437);
  not g17075 (n_6952, n10440);
  and g17076 (n10441, n_6951, n_6952);
  and g17077 (n10442, n_4482, n_6947);
  and g17078 (n10443, n_6948, n10442);
  not g17079 (n_6953, n10441);
  not g17080 (n_6954, n10443);
  and g17081 (n10444, n_6953, n_6954);
  not g17082 (n_6955, n10434);
  not g17083 (n_6956, n10444);
  and g17084 (n10445, n_6955, n_6956);
  not g17085 (n_6957, n10445);
  and g17086 (n10446, \asqrt[34] , n_6957);
  and g17090 (n10450, n_6619, n_6618);
  and g17091 (n10451, \asqrt[23] , n10450);
  not g17092 (n_6958, n10451);
  and g17093 (n10452, n_6617, n_6958);
  not g17094 (n_6959, n10449);
  not g17095 (n_6960, n10452);
  and g17096 (n10453, n_6959, n_6960);
  and g17097 (n10454, n_4218, n_6955);
  and g17098 (n10455, n_6956, n10454);
  not g17099 (n_6961, n10453);
  not g17100 (n_6962, n10455);
  and g17101 (n10456, n_6961, n_6962);
  not g17102 (n_6963, n10446);
  not g17103 (n_6964, n10456);
  and g17104 (n10457, n_6963, n_6964);
  not g17105 (n_6965, n10457);
  and g17106 (n10458, \asqrt[35] , n_6965);
  and g17110 (n10462, n_6627, n_6626);
  and g17111 (n10463, \asqrt[23] , n10462);
  not g17112 (n_6966, n10463);
  and g17113 (n10464, n_6625, n_6966);
  not g17114 (n_6967, n10461);
  not g17115 (n_6968, n10464);
  and g17116 (n10465, n_6967, n_6968);
  and g17117 (n10466, n_3962, n_6963);
  and g17118 (n10467, n_6964, n10466);
  not g17119 (n_6969, n10465);
  not g17120 (n_6970, n10467);
  and g17121 (n10468, n_6969, n_6970);
  not g17122 (n_6971, n10458);
  not g17123 (n_6972, n10468);
  and g17124 (n10469, n_6971, n_6972);
  not g17125 (n_6973, n10469);
  and g17126 (n10470, \asqrt[36] , n_6973);
  and g17130 (n10474, n_6635, n_6634);
  and g17131 (n10475, \asqrt[23] , n10474);
  not g17132 (n_6974, n10475);
  and g17133 (n10476, n_6633, n_6974);
  not g17134 (n_6975, n10473);
  not g17135 (n_6976, n10476);
  and g17136 (n10477, n_6975, n_6976);
  and g17137 (n10478, n_3714, n_6971);
  and g17138 (n10479, n_6972, n10478);
  not g17139 (n_6977, n10477);
  not g17140 (n_6978, n10479);
  and g17141 (n10480, n_6977, n_6978);
  not g17142 (n_6979, n10470);
  not g17143 (n_6980, n10480);
  and g17144 (n10481, n_6979, n_6980);
  not g17145 (n_6981, n10481);
  and g17146 (n10482, \asqrt[37] , n_6981);
  and g17150 (n10486, n_6643, n_6642);
  and g17151 (n10487, \asqrt[23] , n10486);
  not g17152 (n_6982, n10487);
  and g17153 (n10488, n_6641, n_6982);
  not g17154 (n_6983, n10485);
  not g17155 (n_6984, n10488);
  and g17156 (n10489, n_6983, n_6984);
  and g17157 (n10490, n_3474, n_6979);
  and g17158 (n10491, n_6980, n10490);
  not g17159 (n_6985, n10489);
  not g17160 (n_6986, n10491);
  and g17161 (n10492, n_6985, n_6986);
  not g17162 (n_6987, n10482);
  not g17163 (n_6988, n10492);
  and g17164 (n10493, n_6987, n_6988);
  not g17165 (n_6989, n10493);
  and g17166 (n10494, \asqrt[38] , n_6989);
  and g17170 (n10498, n_6651, n_6650);
  and g17171 (n10499, \asqrt[23] , n10498);
  not g17172 (n_6990, n10499);
  and g17173 (n10500, n_6649, n_6990);
  not g17174 (n_6991, n10497);
  not g17175 (n_6992, n10500);
  and g17176 (n10501, n_6991, n_6992);
  and g17177 (n10502, n_3242, n_6987);
  and g17178 (n10503, n_6988, n10502);
  not g17179 (n_6993, n10501);
  not g17180 (n_6994, n10503);
  and g17181 (n10504, n_6993, n_6994);
  not g17182 (n_6995, n10494);
  not g17183 (n_6996, n10504);
  and g17184 (n10505, n_6995, n_6996);
  not g17185 (n_6997, n10505);
  and g17186 (n10506, \asqrt[39] , n_6997);
  and g17190 (n10510, n_6659, n_6658);
  and g17191 (n10511, \asqrt[23] , n10510);
  not g17192 (n_6998, n10511);
  and g17193 (n10512, n_6657, n_6998);
  not g17194 (n_6999, n10509);
  not g17195 (n_7000, n10512);
  and g17196 (n10513, n_6999, n_7000);
  and g17197 (n10514, n_3018, n_6995);
  and g17198 (n10515, n_6996, n10514);
  not g17199 (n_7001, n10513);
  not g17200 (n_7002, n10515);
  and g17201 (n10516, n_7001, n_7002);
  not g17202 (n_7003, n10506);
  not g17203 (n_7004, n10516);
  and g17204 (n10517, n_7003, n_7004);
  not g17205 (n_7005, n10517);
  and g17206 (n10518, \asqrt[40] , n_7005);
  and g17210 (n10522, n_6667, n_6666);
  and g17211 (n10523, \asqrt[23] , n10522);
  not g17212 (n_7006, n10523);
  and g17213 (n10524, n_6665, n_7006);
  not g17214 (n_7007, n10521);
  not g17215 (n_7008, n10524);
  and g17216 (n10525, n_7007, n_7008);
  and g17217 (n10526, n_2802, n_7003);
  and g17218 (n10527, n_7004, n10526);
  not g17219 (n_7009, n10525);
  not g17220 (n_7010, n10527);
  and g17221 (n10528, n_7009, n_7010);
  not g17222 (n_7011, n10518);
  not g17223 (n_7012, n10528);
  and g17224 (n10529, n_7011, n_7012);
  not g17225 (n_7013, n10529);
  and g17226 (n10530, \asqrt[41] , n_7013);
  and g17230 (n10534, n_6675, n_6674);
  and g17231 (n10535, \asqrt[23] , n10534);
  not g17232 (n_7014, n10535);
  and g17233 (n10536, n_6673, n_7014);
  not g17234 (n_7015, n10533);
  not g17235 (n_7016, n10536);
  and g17236 (n10537, n_7015, n_7016);
  and g17237 (n10538, n_2594, n_7011);
  and g17238 (n10539, n_7012, n10538);
  not g17239 (n_7017, n10537);
  not g17240 (n_7018, n10539);
  and g17241 (n10540, n_7017, n_7018);
  not g17242 (n_7019, n10530);
  not g17243 (n_7020, n10540);
  and g17244 (n10541, n_7019, n_7020);
  not g17245 (n_7021, n10541);
  and g17246 (n10542, \asqrt[42] , n_7021);
  and g17247 (n10543, n_2394, n_7019);
  and g17248 (n10544, n_7020, n10543);
  and g17252 (n10548, n_6683, n_6681);
  and g17253 (n10549, \asqrt[23] , n10548);
  not g17254 (n_7022, n10549);
  and g17255 (n10550, n_6682, n_7022);
  not g17256 (n_7023, n10547);
  not g17257 (n_7024, n10550);
  and g17258 (n10551, n_7023, n_7024);
  not g17259 (n_7025, n10544);
  not g17260 (n_7026, n10551);
  and g17261 (n10552, n_7025, n_7026);
  not g17262 (n_7027, n10542);
  not g17263 (n_7028, n10552);
  and g17264 (n10553, n_7027, n_7028);
  not g17265 (n_7029, n10553);
  and g17266 (n10554, \asqrt[43] , n_7029);
  and g17270 (n10558, n_6691, n_6690);
  and g17271 (n10559, \asqrt[23] , n10558);
  not g17272 (n_7030, n10559);
  and g17273 (n10560, n_6689, n_7030);
  not g17274 (n_7031, n10557);
  not g17275 (n_7032, n10560);
  and g17276 (n10561, n_7031, n_7032);
  and g17277 (n10562, n_2202, n_7027);
  and g17278 (n10563, n_7028, n10562);
  not g17279 (n_7033, n10561);
  not g17280 (n_7034, n10563);
  and g17281 (n10564, n_7033, n_7034);
  not g17282 (n_7035, n10554);
  not g17283 (n_7036, n10564);
  and g17284 (n10565, n_7035, n_7036);
  not g17285 (n_7037, n10565);
  and g17286 (n10566, \asqrt[44] , n_7037);
  and g17290 (n10570, n_6699, n_6698);
  and g17291 (n10571, \asqrt[23] , n10570);
  not g17292 (n_7038, n10571);
  and g17293 (n10572, n_6697, n_7038);
  not g17294 (n_7039, n10569);
  not g17295 (n_7040, n10572);
  and g17296 (n10573, n_7039, n_7040);
  and g17297 (n10574, n_2018, n_7035);
  and g17298 (n10575, n_7036, n10574);
  not g17299 (n_7041, n10573);
  not g17300 (n_7042, n10575);
  and g17301 (n10576, n_7041, n_7042);
  not g17302 (n_7043, n10566);
  not g17303 (n_7044, n10576);
  and g17304 (n10577, n_7043, n_7044);
  not g17305 (n_7045, n10577);
  and g17306 (n10578, \asqrt[45] , n_7045);
  and g17310 (n10582, n_6707, n_6706);
  and g17311 (n10583, \asqrt[23] , n10582);
  not g17312 (n_7046, n10583);
  and g17313 (n10584, n_6705, n_7046);
  not g17314 (n_7047, n10581);
  not g17315 (n_7048, n10584);
  and g17316 (n10585, n_7047, n_7048);
  and g17317 (n10586, n_1842, n_7043);
  and g17318 (n10587, n_7044, n10586);
  not g17319 (n_7049, n10585);
  not g17320 (n_7050, n10587);
  and g17321 (n10588, n_7049, n_7050);
  not g17322 (n_7051, n10578);
  not g17323 (n_7052, n10588);
  and g17324 (n10589, n_7051, n_7052);
  not g17325 (n_7053, n10589);
  and g17326 (n10590, \asqrt[46] , n_7053);
  and g17330 (n10594, n_6715, n_6714);
  and g17331 (n10595, \asqrt[23] , n10594);
  not g17332 (n_7054, n10595);
  and g17333 (n10596, n_6713, n_7054);
  not g17334 (n_7055, n10593);
  not g17335 (n_7056, n10596);
  and g17336 (n10597, n_7055, n_7056);
  and g17337 (n10598, n_1674, n_7051);
  and g17338 (n10599, n_7052, n10598);
  not g17339 (n_7057, n10597);
  not g17340 (n_7058, n10599);
  and g17341 (n10600, n_7057, n_7058);
  not g17342 (n_7059, n10590);
  not g17343 (n_7060, n10600);
  and g17344 (n10601, n_7059, n_7060);
  not g17345 (n_7061, n10601);
  and g17346 (n10602, \asqrt[47] , n_7061);
  and g17350 (n10606, n_6723, n_6722);
  and g17351 (n10607, \asqrt[23] , n10606);
  not g17352 (n_7062, n10607);
  and g17353 (n10608, n_6721, n_7062);
  not g17354 (n_7063, n10605);
  not g17355 (n_7064, n10608);
  and g17356 (n10609, n_7063, n_7064);
  and g17357 (n10610, n_1514, n_7059);
  and g17358 (n10611, n_7060, n10610);
  not g17359 (n_7065, n10609);
  not g17360 (n_7066, n10611);
  and g17361 (n10612, n_7065, n_7066);
  not g17362 (n_7067, n10602);
  not g17363 (n_7068, n10612);
  and g17364 (n10613, n_7067, n_7068);
  not g17365 (n_7069, n10613);
  and g17366 (n10614, \asqrt[48] , n_7069);
  and g17370 (n10618, n_6731, n_6730);
  and g17371 (n10619, \asqrt[23] , n10618);
  not g17372 (n_7070, n10619);
  and g17373 (n10620, n_6729, n_7070);
  not g17374 (n_7071, n10617);
  not g17375 (n_7072, n10620);
  and g17376 (n10621, n_7071, n_7072);
  and g17377 (n10622, n_1362, n_7067);
  and g17378 (n10623, n_7068, n10622);
  not g17379 (n_7073, n10621);
  not g17380 (n_7074, n10623);
  and g17381 (n10624, n_7073, n_7074);
  not g17382 (n_7075, n10614);
  not g17383 (n_7076, n10624);
  and g17384 (n10625, n_7075, n_7076);
  not g17385 (n_7077, n10625);
  and g17386 (n10626, \asqrt[49] , n_7077);
  and g17390 (n10630, n_6739, n_6738);
  and g17391 (n10631, \asqrt[23] , n10630);
  not g17392 (n_7078, n10631);
  and g17393 (n10632, n_6737, n_7078);
  not g17394 (n_7079, n10629);
  not g17395 (n_7080, n10632);
  and g17396 (n10633, n_7079, n_7080);
  and g17397 (n10634, n_1218, n_7075);
  and g17398 (n10635, n_7076, n10634);
  not g17399 (n_7081, n10633);
  not g17400 (n_7082, n10635);
  and g17401 (n10636, n_7081, n_7082);
  not g17402 (n_7083, n10626);
  not g17403 (n_7084, n10636);
  and g17404 (n10637, n_7083, n_7084);
  not g17405 (n_7085, n10637);
  and g17406 (n10638, \asqrt[50] , n_7085);
  and g17410 (n10642, n_6747, n_6746);
  and g17411 (n10643, \asqrt[23] , n10642);
  not g17412 (n_7086, n10643);
  and g17413 (n10644, n_6745, n_7086);
  not g17414 (n_7087, n10641);
  not g17415 (n_7088, n10644);
  and g17416 (n10645, n_7087, n_7088);
  and g17417 (n10646, n_1082, n_7083);
  and g17418 (n10647, n_7084, n10646);
  not g17419 (n_7089, n10645);
  not g17420 (n_7090, n10647);
  and g17421 (n10648, n_7089, n_7090);
  not g17422 (n_7091, n10638);
  not g17423 (n_7092, n10648);
  and g17424 (n10649, n_7091, n_7092);
  not g17425 (n_7093, n10649);
  and g17426 (n10650, \asqrt[51] , n_7093);
  and g17430 (n10654, n_6755, n_6754);
  and g17431 (n10655, \asqrt[23] , n10654);
  not g17432 (n_7094, n10655);
  and g17433 (n10656, n_6753, n_7094);
  not g17434 (n_7095, n10653);
  not g17435 (n_7096, n10656);
  and g17436 (n10657, n_7095, n_7096);
  and g17437 (n10658, n_954, n_7091);
  and g17438 (n10659, n_7092, n10658);
  not g17439 (n_7097, n10657);
  not g17440 (n_7098, n10659);
  and g17441 (n10660, n_7097, n_7098);
  not g17442 (n_7099, n10650);
  not g17443 (n_7100, n10660);
  and g17444 (n10661, n_7099, n_7100);
  not g17445 (n_7101, n10661);
  and g17446 (n10662, \asqrt[52] , n_7101);
  and g17450 (n10666, n_6763, n_6762);
  and g17451 (n10667, \asqrt[23] , n10666);
  not g17452 (n_7102, n10667);
  and g17453 (n10668, n_6761, n_7102);
  not g17454 (n_7103, n10665);
  not g17455 (n_7104, n10668);
  and g17456 (n10669, n_7103, n_7104);
  and g17457 (n10670, n_834, n_7099);
  and g17458 (n10671, n_7100, n10670);
  not g17459 (n_7105, n10669);
  not g17460 (n_7106, n10671);
  and g17461 (n10672, n_7105, n_7106);
  not g17462 (n_7107, n10662);
  not g17463 (n_7108, n10672);
  and g17464 (n10673, n_7107, n_7108);
  not g17465 (n_7109, n10673);
  and g17466 (n10674, \asqrt[53] , n_7109);
  and g17470 (n10678, n_6771, n_6770);
  and g17471 (n10679, \asqrt[23] , n10678);
  not g17472 (n_7110, n10679);
  and g17473 (n10680, n_6769, n_7110);
  not g17474 (n_7111, n10677);
  not g17475 (n_7112, n10680);
  and g17476 (n10681, n_7111, n_7112);
  and g17477 (n10682, n_722, n_7107);
  and g17478 (n10683, n_7108, n10682);
  not g17479 (n_7113, n10681);
  not g17480 (n_7114, n10683);
  and g17481 (n10684, n_7113, n_7114);
  not g17482 (n_7115, n10674);
  not g17483 (n_7116, n10684);
  and g17484 (n10685, n_7115, n_7116);
  not g17485 (n_7117, n10685);
  and g17486 (n10686, \asqrt[54] , n_7117);
  and g17490 (n10690, n_6779, n_6778);
  and g17491 (n10691, \asqrt[23] , n10690);
  not g17492 (n_7118, n10691);
  and g17493 (n10692, n_6777, n_7118);
  not g17494 (n_7119, n10689);
  not g17495 (n_7120, n10692);
  and g17496 (n10693, n_7119, n_7120);
  and g17497 (n10694, n_618, n_7115);
  and g17498 (n10695, n_7116, n10694);
  not g17499 (n_7121, n10693);
  not g17500 (n_7122, n10695);
  and g17501 (n10696, n_7121, n_7122);
  not g17502 (n_7123, n10686);
  not g17503 (n_7124, n10696);
  and g17504 (n10697, n_7123, n_7124);
  not g17505 (n_7125, n10697);
  and g17506 (n10698, \asqrt[55] , n_7125);
  and g17510 (n10702, n_6787, n_6786);
  and g17511 (n10703, \asqrt[23] , n10702);
  not g17512 (n_7126, n10703);
  and g17513 (n10704, n_6785, n_7126);
  not g17514 (n_7127, n10701);
  not g17515 (n_7128, n10704);
  and g17516 (n10705, n_7127, n_7128);
  and g17517 (n10706, n_522, n_7123);
  and g17518 (n10707, n_7124, n10706);
  not g17519 (n_7129, n10705);
  not g17520 (n_7130, n10707);
  and g17521 (n10708, n_7129, n_7130);
  not g17522 (n_7131, n10698);
  not g17523 (n_7132, n10708);
  and g17524 (n10709, n_7131, n_7132);
  not g17525 (n_7133, n10709);
  and g17526 (n10710, \asqrt[56] , n_7133);
  and g17530 (n10714, n_6795, n_6794);
  and g17531 (n10715, \asqrt[23] , n10714);
  not g17532 (n_7134, n10715);
  and g17533 (n10716, n_6793, n_7134);
  not g17534 (n_7135, n10713);
  not g17535 (n_7136, n10716);
  and g17536 (n10717, n_7135, n_7136);
  and g17537 (n10718, n_434, n_7131);
  and g17538 (n10719, n_7132, n10718);
  not g17539 (n_7137, n10717);
  not g17540 (n_7138, n10719);
  and g17541 (n10720, n_7137, n_7138);
  not g17542 (n_7139, n10710);
  not g17543 (n_7140, n10720);
  and g17544 (n10721, n_7139, n_7140);
  not g17545 (n_7141, n10721);
  and g17546 (n10722, \asqrt[57] , n_7141);
  and g17550 (n10726, n_6803, n_6802);
  and g17551 (n10727, \asqrt[23] , n10726);
  not g17552 (n_7142, n10727);
  and g17553 (n10728, n_6801, n_7142);
  not g17554 (n_7143, n10725);
  not g17555 (n_7144, n10728);
  and g17556 (n10729, n_7143, n_7144);
  and g17557 (n10730, n_354, n_7139);
  and g17558 (n10731, n_7140, n10730);
  not g17559 (n_7145, n10729);
  not g17560 (n_7146, n10731);
  and g17561 (n10732, n_7145, n_7146);
  not g17562 (n_7147, n10722);
  not g17563 (n_7148, n10732);
  and g17564 (n10733, n_7147, n_7148);
  not g17565 (n_7149, n10733);
  and g17566 (n10734, \asqrt[58] , n_7149);
  and g17570 (n10738, n_6811, n_6810);
  and g17571 (n10739, \asqrt[23] , n10738);
  not g17572 (n_7150, n10739);
  and g17573 (n10740, n_6809, n_7150);
  not g17574 (n_7151, n10737);
  not g17575 (n_7152, n10740);
  and g17576 (n10741, n_7151, n_7152);
  and g17577 (n10742, n_282, n_7147);
  and g17578 (n10743, n_7148, n10742);
  not g17579 (n_7153, n10741);
  not g17580 (n_7154, n10743);
  and g17581 (n10744, n_7153, n_7154);
  not g17582 (n_7155, n10734);
  not g17583 (n_7156, n10744);
  and g17584 (n10745, n_7155, n_7156);
  not g17585 (n_7157, n10745);
  and g17586 (n10746, \asqrt[59] , n_7157);
  and g17590 (n10750, n_6819, n_6818);
  and g17591 (n10751, \asqrt[23] , n10750);
  not g17592 (n_7158, n10751);
  and g17593 (n10752, n_6817, n_7158);
  not g17594 (n_7159, n10749);
  not g17595 (n_7160, n10752);
  and g17596 (n10753, n_7159, n_7160);
  and g17597 (n10754, n_218, n_7155);
  and g17598 (n10755, n_7156, n10754);
  not g17599 (n_7161, n10753);
  not g17600 (n_7162, n10755);
  and g17601 (n10756, n_7161, n_7162);
  not g17602 (n_7163, n10746);
  not g17603 (n_7164, n10756);
  and g17604 (n10757, n_7163, n_7164);
  not g17605 (n_7165, n10757);
  and g17606 (n10758, \asqrt[60] , n_7165);
  and g17610 (n10762, n_6827, n_6826);
  and g17611 (n10763, \asqrt[23] , n10762);
  not g17612 (n_7166, n10763);
  and g17613 (n10764, n_6825, n_7166);
  not g17614 (n_7167, n10761);
  not g17615 (n_7168, n10764);
  and g17616 (n10765, n_7167, n_7168);
  and g17617 (n10766, n_162, n_7163);
  and g17618 (n10767, n_7164, n10766);
  not g17619 (n_7169, n10765);
  not g17620 (n_7170, n10767);
  and g17621 (n10768, n_7169, n_7170);
  not g17622 (n_7171, n10758);
  not g17623 (n_7172, n10768);
  and g17624 (n10769, n_7171, n_7172);
  not g17625 (n_7173, n10769);
  and g17626 (n10770, \asqrt[61] , n_7173);
  and g17630 (n10774, n_6835, n_6834);
  and g17631 (n10775, \asqrt[23] , n10774);
  not g17632 (n_7174, n10775);
  and g17633 (n10776, n_6833, n_7174);
  not g17634 (n_7175, n10773);
  not g17635 (n_7176, n10776);
  and g17636 (n10777, n_7175, n_7176);
  and g17637 (n10778, n_115, n_7171);
  and g17638 (n10779, n_7172, n10778);
  not g17639 (n_7177, n10777);
  not g17640 (n_7178, n10779);
  and g17641 (n10780, n_7177, n_7178);
  not g17642 (n_7179, n10770);
  not g17643 (n_7180, n10780);
  and g17644 (n10781, n_7179, n_7180);
  not g17645 (n_7181, n10781);
  and g17646 (n10782, \asqrt[62] , n_7181);
  and g17650 (n10786, n_6843, n_6842);
  and g17651 (n10787, \asqrt[23] , n10786);
  not g17652 (n_7182, n10787);
  and g17653 (n10788, n_6841, n_7182);
  not g17654 (n_7183, n10785);
  not g17655 (n_7184, n10788);
  and g17656 (n10789, n_7183, n_7184);
  and g17657 (n10790, n_76, n_7179);
  and g17658 (n10791, n_7180, n10790);
  not g17659 (n_7185, n10789);
  not g17660 (n_7186, n10791);
  and g17661 (n10792, n_7185, n_7186);
  not g17662 (n_7187, n10782);
  not g17663 (n_7188, n10792);
  and g17664 (n10793, n_7187, n_7188);
  and g17668 (n10797, n_6851, n_6850);
  and g17669 (n10798, \asqrt[23] , n10797);
  not g17670 (n_7189, n10798);
  and g17671 (n10799, n_6849, n_7189);
  not g17672 (n_7190, n10796);
  not g17673 (n_7191, n10799);
  and g17674 (n10800, n_7190, n_7191);
  and g17675 (n10801, n_6858, n_6857);
  and g17676 (n10802, \asqrt[23] , n10801);
  not g17679 (n_7193, n10800);
  not g17681 (n_7194, n10793);
  not g17683 (n_7195, n10805);
  and g17684 (n10806, n_21, n_7195);
  and g17685 (n10807, n_7187, n10800);
  and g17686 (n10808, n_7188, n10807);
  and g17687 (n10809, n_6857, \asqrt[23] );
  not g17688 (n_7196, n10809);
  and g17689 (n10810, n10293, n_7196);
  not g17690 (n_7197, n10801);
  and g17691 (n10811, \asqrt[63] , n_7197);
  not g17692 (n_7198, n10810);
  and g17693 (n10812, n_7198, n10811);
  not g17699 (n_7199, n10812);
  not g17700 (n_7200, n10817);
  not g17702 (n_7201, n10808);
  and g17706 (n10821, \a[44] , \asqrt[22] );
  not g17707 (n_7206, \a[42] );
  not g17708 (n_7207, \a[43] );
  and g17709 (n10822, n_7206, n_7207);
  and g17710 (n10823, n_6870, n10822);
  not g17711 (n_7208, n10821);
  not g17712 (n_7209, n10823);
  and g17713 (n10824, n_7208, n_7209);
  not g17714 (n_7210, n10824);
  and g17715 (n10825, \asqrt[23] , n_7210);
  and g17721 (n10831, n_6870, \asqrt[22] );
  not g17722 (n_7211, n10831);
  and g17723 (n10832, \a[45] , n_7211);
  and g17724 (n10833, n10322, \asqrt[22] );
  not g17725 (n_7212, n10832);
  not g17726 (n_7213, n10833);
  and g17727 (n10834, n_7212, n_7213);
  not g17728 (n_7214, n10830);
  and g17729 (n10835, n_7214, n10834);
  not g17730 (n_7215, n10825);
  not g17731 (n_7216, n10835);
  and g17732 (n10836, n_7215, n_7216);
  not g17733 (n_7217, n10836);
  and g17734 (n10837, \asqrt[24] , n_7217);
  not g17735 (n_7218, \asqrt[24] );
  and g17736 (n10838, n_7218, n_7215);
  and g17737 (n10839, n_7216, n10838);
  not g17741 (n_7219, n10806);
  not g17743 (n_7220, n10843);
  and g17744 (n10844, n_7213, n_7220);
  not g17745 (n_7221, n10844);
  and g17746 (n10845, \a[46] , n_7221);
  and g17747 (n10846, n_6542, n_7220);
  and g17748 (n10847, n_7213, n10846);
  not g17749 (n_7222, n10845);
  not g17750 (n_7223, n10847);
  and g17751 (n10848, n_7222, n_7223);
  not g17752 (n_7224, n10839);
  not g17753 (n_7225, n10848);
  and g17754 (n10849, n_7224, n_7225);
  not g17755 (n_7226, n10837);
  not g17756 (n_7227, n10849);
  and g17757 (n10850, n_7226, n_7227);
  not g17758 (n_7228, n10850);
  and g17759 (n10851, \asqrt[25] , n_7228);
  and g17760 (n10852, n_6879, n_6878);
  not g17761 (n_7229, n10334);
  and g17762 (n10853, n_7229, n10852);
  and g17763 (n10854, \asqrt[22] , n10853);
  and g17764 (n10855, \asqrt[22] , n10852);
  not g17765 (n_7230, n10855);
  and g17766 (n10856, n10334, n_7230);
  not g17767 (n_7231, n10854);
  not g17768 (n_7232, n10856);
  and g17769 (n10857, n_7231, n_7232);
  and g17770 (n10858, n_6882, n_7226);
  and g17771 (n10859, n_7227, n10858);
  not g17772 (n_7233, n10857);
  not g17773 (n_7234, n10859);
  and g17774 (n10860, n_7233, n_7234);
  not g17775 (n_7235, n10851);
  not g17776 (n_7236, n10860);
  and g17777 (n10861, n_7235, n_7236);
  not g17778 (n_7237, n10861);
  and g17779 (n10862, \asqrt[26] , n_7237);
  and g17783 (n10866, n_6890, n_6888);
  and g17784 (n10867, \asqrt[22] , n10866);
  not g17785 (n_7238, n10867);
  and g17786 (n10868, n_6889, n_7238);
  not g17787 (n_7239, n10865);
  not g17788 (n_7240, n10868);
  and g17789 (n10869, n_7239, n_7240);
  and g17790 (n10870, n_6554, n_7235);
  and g17791 (n10871, n_7236, n10870);
  not g17792 (n_7241, n10869);
  not g17793 (n_7242, n10871);
  and g17794 (n10872, n_7241, n_7242);
  not g17795 (n_7243, n10862);
  not g17796 (n_7244, n10872);
  and g17797 (n10873, n_7243, n_7244);
  not g17798 (n_7245, n10873);
  and g17799 (n10874, \asqrt[27] , n_7245);
  and g17803 (n10878, n_6899, n_6898);
  and g17804 (n10879, \asqrt[22] , n10878);
  not g17805 (n_7246, n10879);
  and g17806 (n10880, n_6897, n_7246);
  not g17807 (n_7247, n10877);
  not g17808 (n_7248, n10880);
  and g17809 (n10881, n_7247, n_7248);
  and g17810 (n10882, n_6234, n_7243);
  and g17811 (n10883, n_7244, n10882);
  not g17812 (n_7249, n10881);
  not g17813 (n_7250, n10883);
  and g17814 (n10884, n_7249, n_7250);
  not g17815 (n_7251, n10874);
  not g17816 (n_7252, n10884);
  and g17817 (n10885, n_7251, n_7252);
  not g17818 (n_7253, n10885);
  and g17819 (n10886, \asqrt[28] , n_7253);
  and g17823 (n10890, n_6907, n_6906);
  and g17824 (n10891, \asqrt[22] , n10890);
  not g17825 (n_7254, n10891);
  and g17826 (n10892, n_6905, n_7254);
  not g17827 (n_7255, n10889);
  not g17828 (n_7256, n10892);
  and g17829 (n10893, n_7255, n_7256);
  and g17830 (n10894, n_5922, n_7251);
  and g17831 (n10895, n_7252, n10894);
  not g17832 (n_7257, n10893);
  not g17833 (n_7258, n10895);
  and g17834 (n10896, n_7257, n_7258);
  not g17835 (n_7259, n10886);
  not g17836 (n_7260, n10896);
  and g17837 (n10897, n_7259, n_7260);
  not g17838 (n_7261, n10897);
  and g17839 (n10898, \asqrt[29] , n_7261);
  and g17843 (n10902, n_6915, n_6914);
  and g17844 (n10903, \asqrt[22] , n10902);
  not g17845 (n_7262, n10903);
  and g17846 (n10904, n_6913, n_7262);
  not g17847 (n_7263, n10901);
  not g17848 (n_7264, n10904);
  and g17849 (n10905, n_7263, n_7264);
  and g17850 (n10906, n_5618, n_7259);
  and g17851 (n10907, n_7260, n10906);
  not g17852 (n_7265, n10905);
  not g17853 (n_7266, n10907);
  and g17854 (n10908, n_7265, n_7266);
  not g17855 (n_7267, n10898);
  not g17856 (n_7268, n10908);
  and g17857 (n10909, n_7267, n_7268);
  not g17858 (n_7269, n10909);
  and g17859 (n10910, \asqrt[30] , n_7269);
  and g17863 (n10914, n_6923, n_6922);
  and g17864 (n10915, \asqrt[22] , n10914);
  not g17865 (n_7270, n10915);
  and g17866 (n10916, n_6921, n_7270);
  not g17867 (n_7271, n10913);
  not g17868 (n_7272, n10916);
  and g17869 (n10917, n_7271, n_7272);
  and g17870 (n10918, n_5322, n_7267);
  and g17871 (n10919, n_7268, n10918);
  not g17872 (n_7273, n10917);
  not g17873 (n_7274, n10919);
  and g17874 (n10920, n_7273, n_7274);
  not g17875 (n_7275, n10910);
  not g17876 (n_7276, n10920);
  and g17877 (n10921, n_7275, n_7276);
  not g17878 (n_7277, n10921);
  and g17879 (n10922, \asqrt[31] , n_7277);
  and g17883 (n10926, n_6931, n_6930);
  and g17884 (n10927, \asqrt[22] , n10926);
  not g17885 (n_7278, n10927);
  and g17886 (n10928, n_6929, n_7278);
  not g17887 (n_7279, n10925);
  not g17888 (n_7280, n10928);
  and g17889 (n10929, n_7279, n_7280);
  and g17890 (n10930, n_5034, n_7275);
  and g17891 (n10931, n_7276, n10930);
  not g17892 (n_7281, n10929);
  not g17893 (n_7282, n10931);
  and g17894 (n10932, n_7281, n_7282);
  not g17895 (n_7283, n10922);
  not g17896 (n_7284, n10932);
  and g17897 (n10933, n_7283, n_7284);
  not g17898 (n_7285, n10933);
  and g17899 (n10934, \asqrt[32] , n_7285);
  and g17903 (n10938, n_6939, n_6938);
  and g17904 (n10939, \asqrt[22] , n10938);
  not g17905 (n_7286, n10939);
  and g17906 (n10940, n_6937, n_7286);
  not g17907 (n_7287, n10937);
  not g17908 (n_7288, n10940);
  and g17909 (n10941, n_7287, n_7288);
  and g17910 (n10942, n_4754, n_7283);
  and g17911 (n10943, n_7284, n10942);
  not g17912 (n_7289, n10941);
  not g17913 (n_7290, n10943);
  and g17914 (n10944, n_7289, n_7290);
  not g17915 (n_7291, n10934);
  not g17916 (n_7292, n10944);
  and g17917 (n10945, n_7291, n_7292);
  not g17918 (n_7293, n10945);
  and g17919 (n10946, \asqrt[33] , n_7293);
  and g17923 (n10950, n_6947, n_6946);
  and g17924 (n10951, \asqrt[22] , n10950);
  not g17925 (n_7294, n10951);
  and g17926 (n10952, n_6945, n_7294);
  not g17927 (n_7295, n10949);
  not g17928 (n_7296, n10952);
  and g17929 (n10953, n_7295, n_7296);
  and g17930 (n10954, n_4482, n_7291);
  and g17931 (n10955, n_7292, n10954);
  not g17932 (n_7297, n10953);
  not g17933 (n_7298, n10955);
  and g17934 (n10956, n_7297, n_7298);
  not g17935 (n_7299, n10946);
  not g17936 (n_7300, n10956);
  and g17937 (n10957, n_7299, n_7300);
  not g17938 (n_7301, n10957);
  and g17939 (n10958, \asqrt[34] , n_7301);
  and g17943 (n10962, n_6955, n_6954);
  and g17944 (n10963, \asqrt[22] , n10962);
  not g17945 (n_7302, n10963);
  and g17946 (n10964, n_6953, n_7302);
  not g17947 (n_7303, n10961);
  not g17948 (n_7304, n10964);
  and g17949 (n10965, n_7303, n_7304);
  and g17950 (n10966, n_4218, n_7299);
  and g17951 (n10967, n_7300, n10966);
  not g17952 (n_7305, n10965);
  not g17953 (n_7306, n10967);
  and g17954 (n10968, n_7305, n_7306);
  not g17955 (n_7307, n10958);
  not g17956 (n_7308, n10968);
  and g17957 (n10969, n_7307, n_7308);
  not g17958 (n_7309, n10969);
  and g17959 (n10970, \asqrt[35] , n_7309);
  and g17963 (n10974, n_6963, n_6962);
  and g17964 (n10975, \asqrt[22] , n10974);
  not g17965 (n_7310, n10975);
  and g17966 (n10976, n_6961, n_7310);
  not g17967 (n_7311, n10973);
  not g17968 (n_7312, n10976);
  and g17969 (n10977, n_7311, n_7312);
  and g17970 (n10978, n_3962, n_7307);
  and g17971 (n10979, n_7308, n10978);
  not g17972 (n_7313, n10977);
  not g17973 (n_7314, n10979);
  and g17974 (n10980, n_7313, n_7314);
  not g17975 (n_7315, n10970);
  not g17976 (n_7316, n10980);
  and g17977 (n10981, n_7315, n_7316);
  not g17978 (n_7317, n10981);
  and g17979 (n10982, \asqrt[36] , n_7317);
  and g17983 (n10986, n_6971, n_6970);
  and g17984 (n10987, \asqrt[22] , n10986);
  not g17985 (n_7318, n10987);
  and g17986 (n10988, n_6969, n_7318);
  not g17987 (n_7319, n10985);
  not g17988 (n_7320, n10988);
  and g17989 (n10989, n_7319, n_7320);
  and g17990 (n10990, n_3714, n_7315);
  and g17991 (n10991, n_7316, n10990);
  not g17992 (n_7321, n10989);
  not g17993 (n_7322, n10991);
  and g17994 (n10992, n_7321, n_7322);
  not g17995 (n_7323, n10982);
  not g17996 (n_7324, n10992);
  and g17997 (n10993, n_7323, n_7324);
  not g17998 (n_7325, n10993);
  and g17999 (n10994, \asqrt[37] , n_7325);
  and g18003 (n10998, n_6979, n_6978);
  and g18004 (n10999, \asqrt[22] , n10998);
  not g18005 (n_7326, n10999);
  and g18006 (n11000, n_6977, n_7326);
  not g18007 (n_7327, n10997);
  not g18008 (n_7328, n11000);
  and g18009 (n11001, n_7327, n_7328);
  and g18010 (n11002, n_3474, n_7323);
  and g18011 (n11003, n_7324, n11002);
  not g18012 (n_7329, n11001);
  not g18013 (n_7330, n11003);
  and g18014 (n11004, n_7329, n_7330);
  not g18015 (n_7331, n10994);
  not g18016 (n_7332, n11004);
  and g18017 (n11005, n_7331, n_7332);
  not g18018 (n_7333, n11005);
  and g18019 (n11006, \asqrt[38] , n_7333);
  and g18023 (n11010, n_6987, n_6986);
  and g18024 (n11011, \asqrt[22] , n11010);
  not g18025 (n_7334, n11011);
  and g18026 (n11012, n_6985, n_7334);
  not g18027 (n_7335, n11009);
  not g18028 (n_7336, n11012);
  and g18029 (n11013, n_7335, n_7336);
  and g18030 (n11014, n_3242, n_7331);
  and g18031 (n11015, n_7332, n11014);
  not g18032 (n_7337, n11013);
  not g18033 (n_7338, n11015);
  and g18034 (n11016, n_7337, n_7338);
  not g18035 (n_7339, n11006);
  not g18036 (n_7340, n11016);
  and g18037 (n11017, n_7339, n_7340);
  not g18038 (n_7341, n11017);
  and g18039 (n11018, \asqrt[39] , n_7341);
  and g18043 (n11022, n_6995, n_6994);
  and g18044 (n11023, \asqrt[22] , n11022);
  not g18045 (n_7342, n11023);
  and g18046 (n11024, n_6993, n_7342);
  not g18047 (n_7343, n11021);
  not g18048 (n_7344, n11024);
  and g18049 (n11025, n_7343, n_7344);
  and g18050 (n11026, n_3018, n_7339);
  and g18051 (n11027, n_7340, n11026);
  not g18052 (n_7345, n11025);
  not g18053 (n_7346, n11027);
  and g18054 (n11028, n_7345, n_7346);
  not g18055 (n_7347, n11018);
  not g18056 (n_7348, n11028);
  and g18057 (n11029, n_7347, n_7348);
  not g18058 (n_7349, n11029);
  and g18059 (n11030, \asqrt[40] , n_7349);
  and g18063 (n11034, n_7003, n_7002);
  and g18064 (n11035, \asqrt[22] , n11034);
  not g18065 (n_7350, n11035);
  and g18066 (n11036, n_7001, n_7350);
  not g18067 (n_7351, n11033);
  not g18068 (n_7352, n11036);
  and g18069 (n11037, n_7351, n_7352);
  and g18070 (n11038, n_2802, n_7347);
  and g18071 (n11039, n_7348, n11038);
  not g18072 (n_7353, n11037);
  not g18073 (n_7354, n11039);
  and g18074 (n11040, n_7353, n_7354);
  not g18075 (n_7355, n11030);
  not g18076 (n_7356, n11040);
  and g18077 (n11041, n_7355, n_7356);
  not g18078 (n_7357, n11041);
  and g18079 (n11042, \asqrt[41] , n_7357);
  and g18083 (n11046, n_7011, n_7010);
  and g18084 (n11047, \asqrt[22] , n11046);
  not g18085 (n_7358, n11047);
  and g18086 (n11048, n_7009, n_7358);
  not g18087 (n_7359, n11045);
  not g18088 (n_7360, n11048);
  and g18089 (n11049, n_7359, n_7360);
  and g18090 (n11050, n_2594, n_7355);
  and g18091 (n11051, n_7356, n11050);
  not g18092 (n_7361, n11049);
  not g18093 (n_7362, n11051);
  and g18094 (n11052, n_7361, n_7362);
  not g18095 (n_7363, n11042);
  not g18096 (n_7364, n11052);
  and g18097 (n11053, n_7363, n_7364);
  not g18098 (n_7365, n11053);
  and g18099 (n11054, \asqrt[42] , n_7365);
  and g18103 (n11058, n_7019, n_7018);
  and g18104 (n11059, \asqrt[22] , n11058);
  not g18105 (n_7366, n11059);
  and g18106 (n11060, n_7017, n_7366);
  not g18107 (n_7367, n11057);
  not g18108 (n_7368, n11060);
  and g18109 (n11061, n_7367, n_7368);
  and g18110 (n11062, n_2394, n_7363);
  and g18111 (n11063, n_7364, n11062);
  not g18112 (n_7369, n11061);
  not g18113 (n_7370, n11063);
  and g18114 (n11064, n_7369, n_7370);
  not g18115 (n_7371, n11054);
  not g18116 (n_7372, n11064);
  and g18117 (n11065, n_7371, n_7372);
  not g18118 (n_7373, n11065);
  and g18119 (n11066, \asqrt[43] , n_7373);
  and g18120 (n11067, n_2202, n_7371);
  and g18121 (n11068, n_7372, n11067);
  and g18125 (n11072, n_7027, n_7025);
  and g18126 (n11073, \asqrt[22] , n11072);
  not g18127 (n_7374, n11073);
  and g18128 (n11074, n_7026, n_7374);
  not g18129 (n_7375, n11071);
  not g18130 (n_7376, n11074);
  and g18131 (n11075, n_7375, n_7376);
  not g18132 (n_7377, n11068);
  not g18133 (n_7378, n11075);
  and g18134 (n11076, n_7377, n_7378);
  not g18135 (n_7379, n11066);
  not g18136 (n_7380, n11076);
  and g18137 (n11077, n_7379, n_7380);
  not g18138 (n_7381, n11077);
  and g18139 (n11078, \asqrt[44] , n_7381);
  and g18143 (n11082, n_7035, n_7034);
  and g18144 (n11083, \asqrt[22] , n11082);
  not g18145 (n_7382, n11083);
  and g18146 (n11084, n_7033, n_7382);
  not g18147 (n_7383, n11081);
  not g18148 (n_7384, n11084);
  and g18149 (n11085, n_7383, n_7384);
  and g18150 (n11086, n_2018, n_7379);
  and g18151 (n11087, n_7380, n11086);
  not g18152 (n_7385, n11085);
  not g18153 (n_7386, n11087);
  and g18154 (n11088, n_7385, n_7386);
  not g18155 (n_7387, n11078);
  not g18156 (n_7388, n11088);
  and g18157 (n11089, n_7387, n_7388);
  not g18158 (n_7389, n11089);
  and g18159 (n11090, \asqrt[45] , n_7389);
  and g18163 (n11094, n_7043, n_7042);
  and g18164 (n11095, \asqrt[22] , n11094);
  not g18165 (n_7390, n11095);
  and g18166 (n11096, n_7041, n_7390);
  not g18167 (n_7391, n11093);
  not g18168 (n_7392, n11096);
  and g18169 (n11097, n_7391, n_7392);
  and g18170 (n11098, n_1842, n_7387);
  and g18171 (n11099, n_7388, n11098);
  not g18172 (n_7393, n11097);
  not g18173 (n_7394, n11099);
  and g18174 (n11100, n_7393, n_7394);
  not g18175 (n_7395, n11090);
  not g18176 (n_7396, n11100);
  and g18177 (n11101, n_7395, n_7396);
  not g18178 (n_7397, n11101);
  and g18179 (n11102, \asqrt[46] , n_7397);
  and g18183 (n11106, n_7051, n_7050);
  and g18184 (n11107, \asqrt[22] , n11106);
  not g18185 (n_7398, n11107);
  and g18186 (n11108, n_7049, n_7398);
  not g18187 (n_7399, n11105);
  not g18188 (n_7400, n11108);
  and g18189 (n11109, n_7399, n_7400);
  and g18190 (n11110, n_1674, n_7395);
  and g18191 (n11111, n_7396, n11110);
  not g18192 (n_7401, n11109);
  not g18193 (n_7402, n11111);
  and g18194 (n11112, n_7401, n_7402);
  not g18195 (n_7403, n11102);
  not g18196 (n_7404, n11112);
  and g18197 (n11113, n_7403, n_7404);
  not g18198 (n_7405, n11113);
  and g18199 (n11114, \asqrt[47] , n_7405);
  and g18203 (n11118, n_7059, n_7058);
  and g18204 (n11119, \asqrt[22] , n11118);
  not g18205 (n_7406, n11119);
  and g18206 (n11120, n_7057, n_7406);
  not g18207 (n_7407, n11117);
  not g18208 (n_7408, n11120);
  and g18209 (n11121, n_7407, n_7408);
  and g18210 (n11122, n_1514, n_7403);
  and g18211 (n11123, n_7404, n11122);
  not g18212 (n_7409, n11121);
  not g18213 (n_7410, n11123);
  and g18214 (n11124, n_7409, n_7410);
  not g18215 (n_7411, n11114);
  not g18216 (n_7412, n11124);
  and g18217 (n11125, n_7411, n_7412);
  not g18218 (n_7413, n11125);
  and g18219 (n11126, \asqrt[48] , n_7413);
  and g18223 (n11130, n_7067, n_7066);
  and g18224 (n11131, \asqrt[22] , n11130);
  not g18225 (n_7414, n11131);
  and g18226 (n11132, n_7065, n_7414);
  not g18227 (n_7415, n11129);
  not g18228 (n_7416, n11132);
  and g18229 (n11133, n_7415, n_7416);
  and g18230 (n11134, n_1362, n_7411);
  and g18231 (n11135, n_7412, n11134);
  not g18232 (n_7417, n11133);
  not g18233 (n_7418, n11135);
  and g18234 (n11136, n_7417, n_7418);
  not g18235 (n_7419, n11126);
  not g18236 (n_7420, n11136);
  and g18237 (n11137, n_7419, n_7420);
  not g18238 (n_7421, n11137);
  and g18239 (n11138, \asqrt[49] , n_7421);
  and g18243 (n11142, n_7075, n_7074);
  and g18244 (n11143, \asqrt[22] , n11142);
  not g18245 (n_7422, n11143);
  and g18246 (n11144, n_7073, n_7422);
  not g18247 (n_7423, n11141);
  not g18248 (n_7424, n11144);
  and g18249 (n11145, n_7423, n_7424);
  and g18250 (n11146, n_1218, n_7419);
  and g18251 (n11147, n_7420, n11146);
  not g18252 (n_7425, n11145);
  not g18253 (n_7426, n11147);
  and g18254 (n11148, n_7425, n_7426);
  not g18255 (n_7427, n11138);
  not g18256 (n_7428, n11148);
  and g18257 (n11149, n_7427, n_7428);
  not g18258 (n_7429, n11149);
  and g18259 (n11150, \asqrt[50] , n_7429);
  and g18263 (n11154, n_7083, n_7082);
  and g18264 (n11155, \asqrt[22] , n11154);
  not g18265 (n_7430, n11155);
  and g18266 (n11156, n_7081, n_7430);
  not g18267 (n_7431, n11153);
  not g18268 (n_7432, n11156);
  and g18269 (n11157, n_7431, n_7432);
  and g18270 (n11158, n_1082, n_7427);
  and g18271 (n11159, n_7428, n11158);
  not g18272 (n_7433, n11157);
  not g18273 (n_7434, n11159);
  and g18274 (n11160, n_7433, n_7434);
  not g18275 (n_7435, n11150);
  not g18276 (n_7436, n11160);
  and g18277 (n11161, n_7435, n_7436);
  not g18278 (n_7437, n11161);
  and g18279 (n11162, \asqrt[51] , n_7437);
  and g18283 (n11166, n_7091, n_7090);
  and g18284 (n11167, \asqrt[22] , n11166);
  not g18285 (n_7438, n11167);
  and g18286 (n11168, n_7089, n_7438);
  not g18287 (n_7439, n11165);
  not g18288 (n_7440, n11168);
  and g18289 (n11169, n_7439, n_7440);
  and g18290 (n11170, n_954, n_7435);
  and g18291 (n11171, n_7436, n11170);
  not g18292 (n_7441, n11169);
  not g18293 (n_7442, n11171);
  and g18294 (n11172, n_7441, n_7442);
  not g18295 (n_7443, n11162);
  not g18296 (n_7444, n11172);
  and g18297 (n11173, n_7443, n_7444);
  not g18298 (n_7445, n11173);
  and g18299 (n11174, \asqrt[52] , n_7445);
  and g18303 (n11178, n_7099, n_7098);
  and g18304 (n11179, \asqrt[22] , n11178);
  not g18305 (n_7446, n11179);
  and g18306 (n11180, n_7097, n_7446);
  not g18307 (n_7447, n11177);
  not g18308 (n_7448, n11180);
  and g18309 (n11181, n_7447, n_7448);
  and g18310 (n11182, n_834, n_7443);
  and g18311 (n11183, n_7444, n11182);
  not g18312 (n_7449, n11181);
  not g18313 (n_7450, n11183);
  and g18314 (n11184, n_7449, n_7450);
  not g18315 (n_7451, n11174);
  not g18316 (n_7452, n11184);
  and g18317 (n11185, n_7451, n_7452);
  not g18318 (n_7453, n11185);
  and g18319 (n11186, \asqrt[53] , n_7453);
  and g18323 (n11190, n_7107, n_7106);
  and g18324 (n11191, \asqrt[22] , n11190);
  not g18325 (n_7454, n11191);
  and g18326 (n11192, n_7105, n_7454);
  not g18327 (n_7455, n11189);
  not g18328 (n_7456, n11192);
  and g18329 (n11193, n_7455, n_7456);
  and g18330 (n11194, n_722, n_7451);
  and g18331 (n11195, n_7452, n11194);
  not g18332 (n_7457, n11193);
  not g18333 (n_7458, n11195);
  and g18334 (n11196, n_7457, n_7458);
  not g18335 (n_7459, n11186);
  not g18336 (n_7460, n11196);
  and g18337 (n11197, n_7459, n_7460);
  not g18338 (n_7461, n11197);
  and g18339 (n11198, \asqrt[54] , n_7461);
  and g18343 (n11202, n_7115, n_7114);
  and g18344 (n11203, \asqrt[22] , n11202);
  not g18345 (n_7462, n11203);
  and g18346 (n11204, n_7113, n_7462);
  not g18347 (n_7463, n11201);
  not g18348 (n_7464, n11204);
  and g18349 (n11205, n_7463, n_7464);
  and g18350 (n11206, n_618, n_7459);
  and g18351 (n11207, n_7460, n11206);
  not g18352 (n_7465, n11205);
  not g18353 (n_7466, n11207);
  and g18354 (n11208, n_7465, n_7466);
  not g18355 (n_7467, n11198);
  not g18356 (n_7468, n11208);
  and g18357 (n11209, n_7467, n_7468);
  not g18358 (n_7469, n11209);
  and g18359 (n11210, \asqrt[55] , n_7469);
  and g18363 (n11214, n_7123, n_7122);
  and g18364 (n11215, \asqrt[22] , n11214);
  not g18365 (n_7470, n11215);
  and g18366 (n11216, n_7121, n_7470);
  not g18367 (n_7471, n11213);
  not g18368 (n_7472, n11216);
  and g18369 (n11217, n_7471, n_7472);
  and g18370 (n11218, n_522, n_7467);
  and g18371 (n11219, n_7468, n11218);
  not g18372 (n_7473, n11217);
  not g18373 (n_7474, n11219);
  and g18374 (n11220, n_7473, n_7474);
  not g18375 (n_7475, n11210);
  not g18376 (n_7476, n11220);
  and g18377 (n11221, n_7475, n_7476);
  not g18378 (n_7477, n11221);
  and g18379 (n11222, \asqrt[56] , n_7477);
  and g18383 (n11226, n_7131, n_7130);
  and g18384 (n11227, \asqrt[22] , n11226);
  not g18385 (n_7478, n11227);
  and g18386 (n11228, n_7129, n_7478);
  not g18387 (n_7479, n11225);
  not g18388 (n_7480, n11228);
  and g18389 (n11229, n_7479, n_7480);
  and g18390 (n11230, n_434, n_7475);
  and g18391 (n11231, n_7476, n11230);
  not g18392 (n_7481, n11229);
  not g18393 (n_7482, n11231);
  and g18394 (n11232, n_7481, n_7482);
  not g18395 (n_7483, n11222);
  not g18396 (n_7484, n11232);
  and g18397 (n11233, n_7483, n_7484);
  not g18398 (n_7485, n11233);
  and g18399 (n11234, \asqrt[57] , n_7485);
  and g18403 (n11238, n_7139, n_7138);
  and g18404 (n11239, \asqrt[22] , n11238);
  not g18405 (n_7486, n11239);
  and g18406 (n11240, n_7137, n_7486);
  not g18407 (n_7487, n11237);
  not g18408 (n_7488, n11240);
  and g18409 (n11241, n_7487, n_7488);
  and g18410 (n11242, n_354, n_7483);
  and g18411 (n11243, n_7484, n11242);
  not g18412 (n_7489, n11241);
  not g18413 (n_7490, n11243);
  and g18414 (n11244, n_7489, n_7490);
  not g18415 (n_7491, n11234);
  not g18416 (n_7492, n11244);
  and g18417 (n11245, n_7491, n_7492);
  not g18418 (n_7493, n11245);
  and g18419 (n11246, \asqrt[58] , n_7493);
  and g18423 (n11250, n_7147, n_7146);
  and g18424 (n11251, \asqrt[22] , n11250);
  not g18425 (n_7494, n11251);
  and g18426 (n11252, n_7145, n_7494);
  not g18427 (n_7495, n11249);
  not g18428 (n_7496, n11252);
  and g18429 (n11253, n_7495, n_7496);
  and g18430 (n11254, n_282, n_7491);
  and g18431 (n11255, n_7492, n11254);
  not g18432 (n_7497, n11253);
  not g18433 (n_7498, n11255);
  and g18434 (n11256, n_7497, n_7498);
  not g18435 (n_7499, n11246);
  not g18436 (n_7500, n11256);
  and g18437 (n11257, n_7499, n_7500);
  not g18438 (n_7501, n11257);
  and g18439 (n11258, \asqrt[59] , n_7501);
  and g18443 (n11262, n_7155, n_7154);
  and g18444 (n11263, \asqrt[22] , n11262);
  not g18445 (n_7502, n11263);
  and g18446 (n11264, n_7153, n_7502);
  not g18447 (n_7503, n11261);
  not g18448 (n_7504, n11264);
  and g18449 (n11265, n_7503, n_7504);
  and g18450 (n11266, n_218, n_7499);
  and g18451 (n11267, n_7500, n11266);
  not g18452 (n_7505, n11265);
  not g18453 (n_7506, n11267);
  and g18454 (n11268, n_7505, n_7506);
  not g18455 (n_7507, n11258);
  not g18456 (n_7508, n11268);
  and g18457 (n11269, n_7507, n_7508);
  not g18458 (n_7509, n11269);
  and g18459 (n11270, \asqrt[60] , n_7509);
  and g18463 (n11274, n_7163, n_7162);
  and g18464 (n11275, \asqrt[22] , n11274);
  not g18465 (n_7510, n11275);
  and g18466 (n11276, n_7161, n_7510);
  not g18467 (n_7511, n11273);
  not g18468 (n_7512, n11276);
  and g18469 (n11277, n_7511, n_7512);
  and g18470 (n11278, n_162, n_7507);
  and g18471 (n11279, n_7508, n11278);
  not g18472 (n_7513, n11277);
  not g18473 (n_7514, n11279);
  and g18474 (n11280, n_7513, n_7514);
  not g18475 (n_7515, n11270);
  not g18476 (n_7516, n11280);
  and g18477 (n11281, n_7515, n_7516);
  not g18478 (n_7517, n11281);
  and g18479 (n11282, \asqrt[61] , n_7517);
  and g18483 (n11286, n_7171, n_7170);
  and g18484 (n11287, \asqrt[22] , n11286);
  not g18485 (n_7518, n11287);
  and g18486 (n11288, n_7169, n_7518);
  not g18487 (n_7519, n11285);
  not g18488 (n_7520, n11288);
  and g18489 (n11289, n_7519, n_7520);
  and g18490 (n11290, n_115, n_7515);
  and g18491 (n11291, n_7516, n11290);
  not g18492 (n_7521, n11289);
  not g18493 (n_7522, n11291);
  and g18494 (n11292, n_7521, n_7522);
  not g18495 (n_7523, n11282);
  not g18496 (n_7524, n11292);
  and g18497 (n11293, n_7523, n_7524);
  not g18498 (n_7525, n11293);
  and g18499 (n11294, \asqrt[62] , n_7525);
  and g18503 (n11298, n_7179, n_7178);
  and g18504 (n11299, \asqrt[22] , n11298);
  not g18505 (n_7526, n11299);
  and g18506 (n11300, n_7177, n_7526);
  not g18507 (n_7527, n11297);
  not g18508 (n_7528, n11300);
  and g18509 (n11301, n_7527, n_7528);
  and g18510 (n11302, n_76, n_7523);
  and g18511 (n11303, n_7524, n11302);
  not g18512 (n_7529, n11301);
  not g18513 (n_7530, n11303);
  and g18514 (n11304, n_7529, n_7530);
  not g18515 (n_7531, n11294);
  not g18516 (n_7532, n11304);
  and g18517 (n11305, n_7531, n_7532);
  and g18521 (n11309, n_7187, n_7186);
  and g18522 (n11310, \asqrt[22] , n11309);
  not g18523 (n_7533, n11310);
  and g18524 (n11311, n_7185, n_7533);
  not g18525 (n_7534, n11308);
  not g18526 (n_7535, n11311);
  and g18527 (n11312, n_7534, n_7535);
  and g18528 (n11313, n_7194, n_7193);
  and g18529 (n11314, \asqrt[22] , n11313);
  not g18532 (n_7537, n11312);
  not g18534 (n_7538, n11305);
  not g18536 (n_7539, n11317);
  and g18537 (n11318, n_21, n_7539);
  and g18538 (n11319, n_7531, n11312);
  and g18539 (n11320, n_7532, n11319);
  and g18540 (n11321, n_7193, \asqrt[22] );
  not g18541 (n_7540, n11321);
  and g18542 (n11322, n10793, n_7540);
  not g18543 (n_7541, n11313);
  and g18544 (n11323, \asqrt[63] , n_7541);
  not g18545 (n_7542, n11322);
  and g18546 (n11324, n_7542, n11323);
  not g18552 (n_7543, n11324);
  not g18553 (n_7544, n11329);
  not g18555 (n_7545, n11320);
  and g18559 (n11333, \a[42] , \asqrt[21] );
  not g18560 (n_7550, \a[40] );
  not g18561 (n_7551, \a[41] );
  and g18562 (n11334, n_7550, n_7551);
  and g18563 (n11335, n_7206, n11334);
  not g18564 (n_7552, n11333);
  not g18565 (n_7553, n11335);
  and g18566 (n11336, n_7552, n_7553);
  not g18567 (n_7554, n11336);
  and g18568 (n11337, \asqrt[22] , n_7554);
  and g18574 (n11343, n_7206, \asqrt[21] );
  not g18575 (n_7555, n11343);
  and g18576 (n11344, \a[43] , n_7555);
  and g18577 (n11345, n10822, \asqrt[21] );
  not g18578 (n_7556, n11344);
  not g18579 (n_7557, n11345);
  and g18580 (n11346, n_7556, n_7557);
  not g18581 (n_7558, n11342);
  and g18582 (n11347, n_7558, n11346);
  not g18583 (n_7559, n11337);
  not g18584 (n_7560, n11347);
  and g18585 (n11348, n_7559, n_7560);
  not g18586 (n_7561, n11348);
  and g18587 (n11349, \asqrt[23] , n_7561);
  not g18588 (n_7562, \asqrt[23] );
  and g18589 (n11350, n_7562, n_7559);
  and g18590 (n11351, n_7560, n11350);
  not g18594 (n_7563, n11318);
  not g18596 (n_7564, n11355);
  and g18597 (n11356, n_7557, n_7564);
  not g18598 (n_7565, n11356);
  and g18599 (n11357, \a[44] , n_7565);
  and g18600 (n11358, n_6870, n_7564);
  and g18601 (n11359, n_7557, n11358);
  not g18602 (n_7566, n11357);
  not g18603 (n_7567, n11359);
  and g18604 (n11360, n_7566, n_7567);
  not g18605 (n_7568, n11351);
  not g18606 (n_7569, n11360);
  and g18607 (n11361, n_7568, n_7569);
  not g18608 (n_7570, n11349);
  not g18609 (n_7571, n11361);
  and g18610 (n11362, n_7570, n_7571);
  not g18611 (n_7572, n11362);
  and g18612 (n11363, \asqrt[24] , n_7572);
  and g18613 (n11364, n_7215, n_7214);
  not g18614 (n_7573, n10834);
  and g18615 (n11365, n_7573, n11364);
  and g18616 (n11366, \asqrt[21] , n11365);
  and g18617 (n11367, \asqrt[21] , n11364);
  not g18618 (n_7574, n11367);
  and g18619 (n11368, n10834, n_7574);
  not g18620 (n_7575, n11366);
  not g18621 (n_7576, n11368);
  and g18622 (n11369, n_7575, n_7576);
  and g18623 (n11370, n_7218, n_7570);
  and g18624 (n11371, n_7571, n11370);
  not g18625 (n_7577, n11369);
  not g18626 (n_7578, n11371);
  and g18627 (n11372, n_7577, n_7578);
  not g18628 (n_7579, n11363);
  not g18629 (n_7580, n11372);
  and g18630 (n11373, n_7579, n_7580);
  not g18631 (n_7581, n11373);
  and g18632 (n11374, \asqrt[25] , n_7581);
  and g18636 (n11378, n_7226, n_7224);
  and g18637 (n11379, \asqrt[21] , n11378);
  not g18638 (n_7582, n11379);
  and g18639 (n11380, n_7225, n_7582);
  not g18640 (n_7583, n11377);
  not g18641 (n_7584, n11380);
  and g18642 (n11381, n_7583, n_7584);
  and g18643 (n11382, n_6882, n_7579);
  and g18644 (n11383, n_7580, n11382);
  not g18645 (n_7585, n11381);
  not g18646 (n_7586, n11383);
  and g18647 (n11384, n_7585, n_7586);
  not g18648 (n_7587, n11374);
  not g18649 (n_7588, n11384);
  and g18650 (n11385, n_7587, n_7588);
  not g18651 (n_7589, n11385);
  and g18652 (n11386, \asqrt[26] , n_7589);
  and g18656 (n11390, n_7235, n_7234);
  and g18657 (n11391, \asqrt[21] , n11390);
  not g18658 (n_7590, n11391);
  and g18659 (n11392, n_7233, n_7590);
  not g18660 (n_7591, n11389);
  not g18661 (n_7592, n11392);
  and g18662 (n11393, n_7591, n_7592);
  and g18663 (n11394, n_6554, n_7587);
  and g18664 (n11395, n_7588, n11394);
  not g18665 (n_7593, n11393);
  not g18666 (n_7594, n11395);
  and g18667 (n11396, n_7593, n_7594);
  not g18668 (n_7595, n11386);
  not g18669 (n_7596, n11396);
  and g18670 (n11397, n_7595, n_7596);
  not g18671 (n_7597, n11397);
  and g18672 (n11398, \asqrt[27] , n_7597);
  and g18676 (n11402, n_7243, n_7242);
  and g18677 (n11403, \asqrt[21] , n11402);
  not g18678 (n_7598, n11403);
  and g18679 (n11404, n_7241, n_7598);
  not g18680 (n_7599, n11401);
  not g18681 (n_7600, n11404);
  and g18682 (n11405, n_7599, n_7600);
  and g18683 (n11406, n_6234, n_7595);
  and g18684 (n11407, n_7596, n11406);
  not g18685 (n_7601, n11405);
  not g18686 (n_7602, n11407);
  and g18687 (n11408, n_7601, n_7602);
  not g18688 (n_7603, n11398);
  not g18689 (n_7604, n11408);
  and g18690 (n11409, n_7603, n_7604);
  not g18691 (n_7605, n11409);
  and g18692 (n11410, \asqrt[28] , n_7605);
  and g18696 (n11414, n_7251, n_7250);
  and g18697 (n11415, \asqrt[21] , n11414);
  not g18698 (n_7606, n11415);
  and g18699 (n11416, n_7249, n_7606);
  not g18700 (n_7607, n11413);
  not g18701 (n_7608, n11416);
  and g18702 (n11417, n_7607, n_7608);
  and g18703 (n11418, n_5922, n_7603);
  and g18704 (n11419, n_7604, n11418);
  not g18705 (n_7609, n11417);
  not g18706 (n_7610, n11419);
  and g18707 (n11420, n_7609, n_7610);
  not g18708 (n_7611, n11410);
  not g18709 (n_7612, n11420);
  and g18710 (n11421, n_7611, n_7612);
  not g18711 (n_7613, n11421);
  and g18712 (n11422, \asqrt[29] , n_7613);
  and g18716 (n11426, n_7259, n_7258);
  and g18717 (n11427, \asqrt[21] , n11426);
  not g18718 (n_7614, n11427);
  and g18719 (n11428, n_7257, n_7614);
  not g18720 (n_7615, n11425);
  not g18721 (n_7616, n11428);
  and g18722 (n11429, n_7615, n_7616);
  and g18723 (n11430, n_5618, n_7611);
  and g18724 (n11431, n_7612, n11430);
  not g18725 (n_7617, n11429);
  not g18726 (n_7618, n11431);
  and g18727 (n11432, n_7617, n_7618);
  not g18728 (n_7619, n11422);
  not g18729 (n_7620, n11432);
  and g18730 (n11433, n_7619, n_7620);
  not g18731 (n_7621, n11433);
  and g18732 (n11434, \asqrt[30] , n_7621);
  and g18736 (n11438, n_7267, n_7266);
  and g18737 (n11439, \asqrt[21] , n11438);
  not g18738 (n_7622, n11439);
  and g18739 (n11440, n_7265, n_7622);
  not g18740 (n_7623, n11437);
  not g18741 (n_7624, n11440);
  and g18742 (n11441, n_7623, n_7624);
  and g18743 (n11442, n_5322, n_7619);
  and g18744 (n11443, n_7620, n11442);
  not g18745 (n_7625, n11441);
  not g18746 (n_7626, n11443);
  and g18747 (n11444, n_7625, n_7626);
  not g18748 (n_7627, n11434);
  not g18749 (n_7628, n11444);
  and g18750 (n11445, n_7627, n_7628);
  not g18751 (n_7629, n11445);
  and g18752 (n11446, \asqrt[31] , n_7629);
  and g18756 (n11450, n_7275, n_7274);
  and g18757 (n11451, \asqrt[21] , n11450);
  not g18758 (n_7630, n11451);
  and g18759 (n11452, n_7273, n_7630);
  not g18760 (n_7631, n11449);
  not g18761 (n_7632, n11452);
  and g18762 (n11453, n_7631, n_7632);
  and g18763 (n11454, n_5034, n_7627);
  and g18764 (n11455, n_7628, n11454);
  not g18765 (n_7633, n11453);
  not g18766 (n_7634, n11455);
  and g18767 (n11456, n_7633, n_7634);
  not g18768 (n_7635, n11446);
  not g18769 (n_7636, n11456);
  and g18770 (n11457, n_7635, n_7636);
  not g18771 (n_7637, n11457);
  and g18772 (n11458, \asqrt[32] , n_7637);
  and g18776 (n11462, n_7283, n_7282);
  and g18777 (n11463, \asqrt[21] , n11462);
  not g18778 (n_7638, n11463);
  and g18779 (n11464, n_7281, n_7638);
  not g18780 (n_7639, n11461);
  not g18781 (n_7640, n11464);
  and g18782 (n11465, n_7639, n_7640);
  and g18783 (n11466, n_4754, n_7635);
  and g18784 (n11467, n_7636, n11466);
  not g18785 (n_7641, n11465);
  not g18786 (n_7642, n11467);
  and g18787 (n11468, n_7641, n_7642);
  not g18788 (n_7643, n11458);
  not g18789 (n_7644, n11468);
  and g18790 (n11469, n_7643, n_7644);
  not g18791 (n_7645, n11469);
  and g18792 (n11470, \asqrt[33] , n_7645);
  and g18796 (n11474, n_7291, n_7290);
  and g18797 (n11475, \asqrt[21] , n11474);
  not g18798 (n_7646, n11475);
  and g18799 (n11476, n_7289, n_7646);
  not g18800 (n_7647, n11473);
  not g18801 (n_7648, n11476);
  and g18802 (n11477, n_7647, n_7648);
  and g18803 (n11478, n_4482, n_7643);
  and g18804 (n11479, n_7644, n11478);
  not g18805 (n_7649, n11477);
  not g18806 (n_7650, n11479);
  and g18807 (n11480, n_7649, n_7650);
  not g18808 (n_7651, n11470);
  not g18809 (n_7652, n11480);
  and g18810 (n11481, n_7651, n_7652);
  not g18811 (n_7653, n11481);
  and g18812 (n11482, \asqrt[34] , n_7653);
  and g18816 (n11486, n_7299, n_7298);
  and g18817 (n11487, \asqrt[21] , n11486);
  not g18818 (n_7654, n11487);
  and g18819 (n11488, n_7297, n_7654);
  not g18820 (n_7655, n11485);
  not g18821 (n_7656, n11488);
  and g18822 (n11489, n_7655, n_7656);
  and g18823 (n11490, n_4218, n_7651);
  and g18824 (n11491, n_7652, n11490);
  not g18825 (n_7657, n11489);
  not g18826 (n_7658, n11491);
  and g18827 (n11492, n_7657, n_7658);
  not g18828 (n_7659, n11482);
  not g18829 (n_7660, n11492);
  and g18830 (n11493, n_7659, n_7660);
  not g18831 (n_7661, n11493);
  and g18832 (n11494, \asqrt[35] , n_7661);
  and g18836 (n11498, n_7307, n_7306);
  and g18837 (n11499, \asqrt[21] , n11498);
  not g18838 (n_7662, n11499);
  and g18839 (n11500, n_7305, n_7662);
  not g18840 (n_7663, n11497);
  not g18841 (n_7664, n11500);
  and g18842 (n11501, n_7663, n_7664);
  and g18843 (n11502, n_3962, n_7659);
  and g18844 (n11503, n_7660, n11502);
  not g18845 (n_7665, n11501);
  not g18846 (n_7666, n11503);
  and g18847 (n11504, n_7665, n_7666);
  not g18848 (n_7667, n11494);
  not g18849 (n_7668, n11504);
  and g18850 (n11505, n_7667, n_7668);
  not g18851 (n_7669, n11505);
  and g18852 (n11506, \asqrt[36] , n_7669);
  and g18856 (n11510, n_7315, n_7314);
  and g18857 (n11511, \asqrt[21] , n11510);
  not g18858 (n_7670, n11511);
  and g18859 (n11512, n_7313, n_7670);
  not g18860 (n_7671, n11509);
  not g18861 (n_7672, n11512);
  and g18862 (n11513, n_7671, n_7672);
  and g18863 (n11514, n_3714, n_7667);
  and g18864 (n11515, n_7668, n11514);
  not g18865 (n_7673, n11513);
  not g18866 (n_7674, n11515);
  and g18867 (n11516, n_7673, n_7674);
  not g18868 (n_7675, n11506);
  not g18869 (n_7676, n11516);
  and g18870 (n11517, n_7675, n_7676);
  not g18871 (n_7677, n11517);
  and g18872 (n11518, \asqrt[37] , n_7677);
  and g18876 (n11522, n_7323, n_7322);
  and g18877 (n11523, \asqrt[21] , n11522);
  not g18878 (n_7678, n11523);
  and g18879 (n11524, n_7321, n_7678);
  not g18880 (n_7679, n11521);
  not g18881 (n_7680, n11524);
  and g18882 (n11525, n_7679, n_7680);
  and g18883 (n11526, n_3474, n_7675);
  and g18884 (n11527, n_7676, n11526);
  not g18885 (n_7681, n11525);
  not g18886 (n_7682, n11527);
  and g18887 (n11528, n_7681, n_7682);
  not g18888 (n_7683, n11518);
  not g18889 (n_7684, n11528);
  and g18890 (n11529, n_7683, n_7684);
  not g18891 (n_7685, n11529);
  and g18892 (n11530, \asqrt[38] , n_7685);
  and g18896 (n11534, n_7331, n_7330);
  and g18897 (n11535, \asqrt[21] , n11534);
  not g18898 (n_7686, n11535);
  and g18899 (n11536, n_7329, n_7686);
  not g18900 (n_7687, n11533);
  not g18901 (n_7688, n11536);
  and g18902 (n11537, n_7687, n_7688);
  and g18903 (n11538, n_3242, n_7683);
  and g18904 (n11539, n_7684, n11538);
  not g18905 (n_7689, n11537);
  not g18906 (n_7690, n11539);
  and g18907 (n11540, n_7689, n_7690);
  not g18908 (n_7691, n11530);
  not g18909 (n_7692, n11540);
  and g18910 (n11541, n_7691, n_7692);
  not g18911 (n_7693, n11541);
  and g18912 (n11542, \asqrt[39] , n_7693);
  and g18916 (n11546, n_7339, n_7338);
  and g18917 (n11547, \asqrt[21] , n11546);
  not g18918 (n_7694, n11547);
  and g18919 (n11548, n_7337, n_7694);
  not g18920 (n_7695, n11545);
  not g18921 (n_7696, n11548);
  and g18922 (n11549, n_7695, n_7696);
  and g18923 (n11550, n_3018, n_7691);
  and g18924 (n11551, n_7692, n11550);
  not g18925 (n_7697, n11549);
  not g18926 (n_7698, n11551);
  and g18927 (n11552, n_7697, n_7698);
  not g18928 (n_7699, n11542);
  not g18929 (n_7700, n11552);
  and g18930 (n11553, n_7699, n_7700);
  not g18931 (n_7701, n11553);
  and g18932 (n11554, \asqrt[40] , n_7701);
  and g18936 (n11558, n_7347, n_7346);
  and g18937 (n11559, \asqrt[21] , n11558);
  not g18938 (n_7702, n11559);
  and g18939 (n11560, n_7345, n_7702);
  not g18940 (n_7703, n11557);
  not g18941 (n_7704, n11560);
  and g18942 (n11561, n_7703, n_7704);
  and g18943 (n11562, n_2802, n_7699);
  and g18944 (n11563, n_7700, n11562);
  not g18945 (n_7705, n11561);
  not g18946 (n_7706, n11563);
  and g18947 (n11564, n_7705, n_7706);
  not g18948 (n_7707, n11554);
  not g18949 (n_7708, n11564);
  and g18950 (n11565, n_7707, n_7708);
  not g18951 (n_7709, n11565);
  and g18952 (n11566, \asqrt[41] , n_7709);
  and g18956 (n11570, n_7355, n_7354);
  and g18957 (n11571, \asqrt[21] , n11570);
  not g18958 (n_7710, n11571);
  and g18959 (n11572, n_7353, n_7710);
  not g18960 (n_7711, n11569);
  not g18961 (n_7712, n11572);
  and g18962 (n11573, n_7711, n_7712);
  and g18963 (n11574, n_2594, n_7707);
  and g18964 (n11575, n_7708, n11574);
  not g18965 (n_7713, n11573);
  not g18966 (n_7714, n11575);
  and g18967 (n11576, n_7713, n_7714);
  not g18968 (n_7715, n11566);
  not g18969 (n_7716, n11576);
  and g18970 (n11577, n_7715, n_7716);
  not g18971 (n_7717, n11577);
  and g18972 (n11578, \asqrt[42] , n_7717);
  and g18976 (n11582, n_7363, n_7362);
  and g18977 (n11583, \asqrt[21] , n11582);
  not g18978 (n_7718, n11583);
  and g18979 (n11584, n_7361, n_7718);
  not g18980 (n_7719, n11581);
  not g18981 (n_7720, n11584);
  and g18982 (n11585, n_7719, n_7720);
  and g18983 (n11586, n_2394, n_7715);
  and g18984 (n11587, n_7716, n11586);
  not g18985 (n_7721, n11585);
  not g18986 (n_7722, n11587);
  and g18987 (n11588, n_7721, n_7722);
  not g18988 (n_7723, n11578);
  not g18989 (n_7724, n11588);
  and g18990 (n11589, n_7723, n_7724);
  not g18991 (n_7725, n11589);
  and g18992 (n11590, \asqrt[43] , n_7725);
  and g18996 (n11594, n_7371, n_7370);
  and g18997 (n11595, \asqrt[21] , n11594);
  not g18998 (n_7726, n11595);
  and g18999 (n11596, n_7369, n_7726);
  not g19000 (n_7727, n11593);
  not g19001 (n_7728, n11596);
  and g19002 (n11597, n_7727, n_7728);
  and g19003 (n11598, n_2202, n_7723);
  and g19004 (n11599, n_7724, n11598);
  not g19005 (n_7729, n11597);
  not g19006 (n_7730, n11599);
  and g19007 (n11600, n_7729, n_7730);
  not g19008 (n_7731, n11590);
  not g19009 (n_7732, n11600);
  and g19010 (n11601, n_7731, n_7732);
  not g19011 (n_7733, n11601);
  and g19012 (n11602, \asqrt[44] , n_7733);
  and g19013 (n11603, n_2018, n_7731);
  and g19014 (n11604, n_7732, n11603);
  and g19018 (n11608, n_7379, n_7377);
  and g19019 (n11609, \asqrt[21] , n11608);
  not g19020 (n_7734, n11609);
  and g19021 (n11610, n_7378, n_7734);
  not g19022 (n_7735, n11607);
  not g19023 (n_7736, n11610);
  and g19024 (n11611, n_7735, n_7736);
  not g19025 (n_7737, n11604);
  not g19026 (n_7738, n11611);
  and g19027 (n11612, n_7737, n_7738);
  not g19028 (n_7739, n11602);
  not g19029 (n_7740, n11612);
  and g19030 (n11613, n_7739, n_7740);
  not g19031 (n_7741, n11613);
  and g19032 (n11614, \asqrt[45] , n_7741);
  and g19036 (n11618, n_7387, n_7386);
  and g19037 (n11619, \asqrt[21] , n11618);
  not g19038 (n_7742, n11619);
  and g19039 (n11620, n_7385, n_7742);
  not g19040 (n_7743, n11617);
  not g19041 (n_7744, n11620);
  and g19042 (n11621, n_7743, n_7744);
  and g19043 (n11622, n_1842, n_7739);
  and g19044 (n11623, n_7740, n11622);
  not g19045 (n_7745, n11621);
  not g19046 (n_7746, n11623);
  and g19047 (n11624, n_7745, n_7746);
  not g19048 (n_7747, n11614);
  not g19049 (n_7748, n11624);
  and g19050 (n11625, n_7747, n_7748);
  not g19051 (n_7749, n11625);
  and g19052 (n11626, \asqrt[46] , n_7749);
  and g19056 (n11630, n_7395, n_7394);
  and g19057 (n11631, \asqrt[21] , n11630);
  not g19058 (n_7750, n11631);
  and g19059 (n11632, n_7393, n_7750);
  not g19060 (n_7751, n11629);
  not g19061 (n_7752, n11632);
  and g19062 (n11633, n_7751, n_7752);
  and g19063 (n11634, n_1674, n_7747);
  and g19064 (n11635, n_7748, n11634);
  not g19065 (n_7753, n11633);
  not g19066 (n_7754, n11635);
  and g19067 (n11636, n_7753, n_7754);
  not g19068 (n_7755, n11626);
  not g19069 (n_7756, n11636);
  and g19070 (n11637, n_7755, n_7756);
  not g19071 (n_7757, n11637);
  and g19072 (n11638, \asqrt[47] , n_7757);
  and g19076 (n11642, n_7403, n_7402);
  and g19077 (n11643, \asqrt[21] , n11642);
  not g19078 (n_7758, n11643);
  and g19079 (n11644, n_7401, n_7758);
  not g19080 (n_7759, n11641);
  not g19081 (n_7760, n11644);
  and g19082 (n11645, n_7759, n_7760);
  and g19083 (n11646, n_1514, n_7755);
  and g19084 (n11647, n_7756, n11646);
  not g19085 (n_7761, n11645);
  not g19086 (n_7762, n11647);
  and g19087 (n11648, n_7761, n_7762);
  not g19088 (n_7763, n11638);
  not g19089 (n_7764, n11648);
  and g19090 (n11649, n_7763, n_7764);
  not g19091 (n_7765, n11649);
  and g19092 (n11650, \asqrt[48] , n_7765);
  and g19096 (n11654, n_7411, n_7410);
  and g19097 (n11655, \asqrt[21] , n11654);
  not g19098 (n_7766, n11655);
  and g19099 (n11656, n_7409, n_7766);
  not g19100 (n_7767, n11653);
  not g19101 (n_7768, n11656);
  and g19102 (n11657, n_7767, n_7768);
  and g19103 (n11658, n_1362, n_7763);
  and g19104 (n11659, n_7764, n11658);
  not g19105 (n_7769, n11657);
  not g19106 (n_7770, n11659);
  and g19107 (n11660, n_7769, n_7770);
  not g19108 (n_7771, n11650);
  not g19109 (n_7772, n11660);
  and g19110 (n11661, n_7771, n_7772);
  not g19111 (n_7773, n11661);
  and g19112 (n11662, \asqrt[49] , n_7773);
  and g19116 (n11666, n_7419, n_7418);
  and g19117 (n11667, \asqrt[21] , n11666);
  not g19118 (n_7774, n11667);
  and g19119 (n11668, n_7417, n_7774);
  not g19120 (n_7775, n11665);
  not g19121 (n_7776, n11668);
  and g19122 (n11669, n_7775, n_7776);
  and g19123 (n11670, n_1218, n_7771);
  and g19124 (n11671, n_7772, n11670);
  not g19125 (n_7777, n11669);
  not g19126 (n_7778, n11671);
  and g19127 (n11672, n_7777, n_7778);
  not g19128 (n_7779, n11662);
  not g19129 (n_7780, n11672);
  and g19130 (n11673, n_7779, n_7780);
  not g19131 (n_7781, n11673);
  and g19132 (n11674, \asqrt[50] , n_7781);
  and g19136 (n11678, n_7427, n_7426);
  and g19137 (n11679, \asqrt[21] , n11678);
  not g19138 (n_7782, n11679);
  and g19139 (n11680, n_7425, n_7782);
  not g19140 (n_7783, n11677);
  not g19141 (n_7784, n11680);
  and g19142 (n11681, n_7783, n_7784);
  and g19143 (n11682, n_1082, n_7779);
  and g19144 (n11683, n_7780, n11682);
  not g19145 (n_7785, n11681);
  not g19146 (n_7786, n11683);
  and g19147 (n11684, n_7785, n_7786);
  not g19148 (n_7787, n11674);
  not g19149 (n_7788, n11684);
  and g19150 (n11685, n_7787, n_7788);
  not g19151 (n_7789, n11685);
  and g19152 (n11686, \asqrt[51] , n_7789);
  and g19156 (n11690, n_7435, n_7434);
  and g19157 (n11691, \asqrt[21] , n11690);
  not g19158 (n_7790, n11691);
  and g19159 (n11692, n_7433, n_7790);
  not g19160 (n_7791, n11689);
  not g19161 (n_7792, n11692);
  and g19162 (n11693, n_7791, n_7792);
  and g19163 (n11694, n_954, n_7787);
  and g19164 (n11695, n_7788, n11694);
  not g19165 (n_7793, n11693);
  not g19166 (n_7794, n11695);
  and g19167 (n11696, n_7793, n_7794);
  not g19168 (n_7795, n11686);
  not g19169 (n_7796, n11696);
  and g19170 (n11697, n_7795, n_7796);
  not g19171 (n_7797, n11697);
  and g19172 (n11698, \asqrt[52] , n_7797);
  and g19176 (n11702, n_7443, n_7442);
  and g19177 (n11703, \asqrt[21] , n11702);
  not g19178 (n_7798, n11703);
  and g19179 (n11704, n_7441, n_7798);
  not g19180 (n_7799, n11701);
  not g19181 (n_7800, n11704);
  and g19182 (n11705, n_7799, n_7800);
  and g19183 (n11706, n_834, n_7795);
  and g19184 (n11707, n_7796, n11706);
  not g19185 (n_7801, n11705);
  not g19186 (n_7802, n11707);
  and g19187 (n11708, n_7801, n_7802);
  not g19188 (n_7803, n11698);
  not g19189 (n_7804, n11708);
  and g19190 (n11709, n_7803, n_7804);
  not g19191 (n_7805, n11709);
  and g19192 (n11710, \asqrt[53] , n_7805);
  and g19196 (n11714, n_7451, n_7450);
  and g19197 (n11715, \asqrt[21] , n11714);
  not g19198 (n_7806, n11715);
  and g19199 (n11716, n_7449, n_7806);
  not g19200 (n_7807, n11713);
  not g19201 (n_7808, n11716);
  and g19202 (n11717, n_7807, n_7808);
  and g19203 (n11718, n_722, n_7803);
  and g19204 (n11719, n_7804, n11718);
  not g19205 (n_7809, n11717);
  not g19206 (n_7810, n11719);
  and g19207 (n11720, n_7809, n_7810);
  not g19208 (n_7811, n11710);
  not g19209 (n_7812, n11720);
  and g19210 (n11721, n_7811, n_7812);
  not g19211 (n_7813, n11721);
  and g19212 (n11722, \asqrt[54] , n_7813);
  and g19216 (n11726, n_7459, n_7458);
  and g19217 (n11727, \asqrt[21] , n11726);
  not g19218 (n_7814, n11727);
  and g19219 (n11728, n_7457, n_7814);
  not g19220 (n_7815, n11725);
  not g19221 (n_7816, n11728);
  and g19222 (n11729, n_7815, n_7816);
  and g19223 (n11730, n_618, n_7811);
  and g19224 (n11731, n_7812, n11730);
  not g19225 (n_7817, n11729);
  not g19226 (n_7818, n11731);
  and g19227 (n11732, n_7817, n_7818);
  not g19228 (n_7819, n11722);
  not g19229 (n_7820, n11732);
  and g19230 (n11733, n_7819, n_7820);
  not g19231 (n_7821, n11733);
  and g19232 (n11734, \asqrt[55] , n_7821);
  and g19236 (n11738, n_7467, n_7466);
  and g19237 (n11739, \asqrt[21] , n11738);
  not g19238 (n_7822, n11739);
  and g19239 (n11740, n_7465, n_7822);
  not g19240 (n_7823, n11737);
  not g19241 (n_7824, n11740);
  and g19242 (n11741, n_7823, n_7824);
  and g19243 (n11742, n_522, n_7819);
  and g19244 (n11743, n_7820, n11742);
  not g19245 (n_7825, n11741);
  not g19246 (n_7826, n11743);
  and g19247 (n11744, n_7825, n_7826);
  not g19248 (n_7827, n11734);
  not g19249 (n_7828, n11744);
  and g19250 (n11745, n_7827, n_7828);
  not g19251 (n_7829, n11745);
  and g19252 (n11746, \asqrt[56] , n_7829);
  and g19256 (n11750, n_7475, n_7474);
  and g19257 (n11751, \asqrt[21] , n11750);
  not g19258 (n_7830, n11751);
  and g19259 (n11752, n_7473, n_7830);
  not g19260 (n_7831, n11749);
  not g19261 (n_7832, n11752);
  and g19262 (n11753, n_7831, n_7832);
  and g19263 (n11754, n_434, n_7827);
  and g19264 (n11755, n_7828, n11754);
  not g19265 (n_7833, n11753);
  not g19266 (n_7834, n11755);
  and g19267 (n11756, n_7833, n_7834);
  not g19268 (n_7835, n11746);
  not g19269 (n_7836, n11756);
  and g19270 (n11757, n_7835, n_7836);
  not g19271 (n_7837, n11757);
  and g19272 (n11758, \asqrt[57] , n_7837);
  and g19276 (n11762, n_7483, n_7482);
  and g19277 (n11763, \asqrt[21] , n11762);
  not g19278 (n_7838, n11763);
  and g19279 (n11764, n_7481, n_7838);
  not g19280 (n_7839, n11761);
  not g19281 (n_7840, n11764);
  and g19282 (n11765, n_7839, n_7840);
  and g19283 (n11766, n_354, n_7835);
  and g19284 (n11767, n_7836, n11766);
  not g19285 (n_7841, n11765);
  not g19286 (n_7842, n11767);
  and g19287 (n11768, n_7841, n_7842);
  not g19288 (n_7843, n11758);
  not g19289 (n_7844, n11768);
  and g19290 (n11769, n_7843, n_7844);
  not g19291 (n_7845, n11769);
  and g19292 (n11770, \asqrt[58] , n_7845);
  and g19296 (n11774, n_7491, n_7490);
  and g19297 (n11775, \asqrt[21] , n11774);
  not g19298 (n_7846, n11775);
  and g19299 (n11776, n_7489, n_7846);
  not g19300 (n_7847, n11773);
  not g19301 (n_7848, n11776);
  and g19302 (n11777, n_7847, n_7848);
  and g19303 (n11778, n_282, n_7843);
  and g19304 (n11779, n_7844, n11778);
  not g19305 (n_7849, n11777);
  not g19306 (n_7850, n11779);
  and g19307 (n11780, n_7849, n_7850);
  not g19308 (n_7851, n11770);
  not g19309 (n_7852, n11780);
  and g19310 (n11781, n_7851, n_7852);
  not g19311 (n_7853, n11781);
  and g19312 (n11782, \asqrt[59] , n_7853);
  and g19316 (n11786, n_7499, n_7498);
  and g19317 (n11787, \asqrt[21] , n11786);
  not g19318 (n_7854, n11787);
  and g19319 (n11788, n_7497, n_7854);
  not g19320 (n_7855, n11785);
  not g19321 (n_7856, n11788);
  and g19322 (n11789, n_7855, n_7856);
  and g19323 (n11790, n_218, n_7851);
  and g19324 (n11791, n_7852, n11790);
  not g19325 (n_7857, n11789);
  not g19326 (n_7858, n11791);
  and g19327 (n11792, n_7857, n_7858);
  not g19328 (n_7859, n11782);
  not g19329 (n_7860, n11792);
  and g19330 (n11793, n_7859, n_7860);
  not g19331 (n_7861, n11793);
  and g19332 (n11794, \asqrt[60] , n_7861);
  and g19336 (n11798, n_7507, n_7506);
  and g19337 (n11799, \asqrt[21] , n11798);
  not g19338 (n_7862, n11799);
  and g19339 (n11800, n_7505, n_7862);
  not g19340 (n_7863, n11797);
  not g19341 (n_7864, n11800);
  and g19342 (n11801, n_7863, n_7864);
  and g19343 (n11802, n_162, n_7859);
  and g19344 (n11803, n_7860, n11802);
  not g19345 (n_7865, n11801);
  not g19346 (n_7866, n11803);
  and g19347 (n11804, n_7865, n_7866);
  not g19348 (n_7867, n11794);
  not g19349 (n_7868, n11804);
  and g19350 (n11805, n_7867, n_7868);
  not g19351 (n_7869, n11805);
  and g19352 (n11806, \asqrt[61] , n_7869);
  and g19356 (n11810, n_7515, n_7514);
  and g19357 (n11811, \asqrt[21] , n11810);
  not g19358 (n_7870, n11811);
  and g19359 (n11812, n_7513, n_7870);
  not g19360 (n_7871, n11809);
  not g19361 (n_7872, n11812);
  and g19362 (n11813, n_7871, n_7872);
  and g19363 (n11814, n_115, n_7867);
  and g19364 (n11815, n_7868, n11814);
  not g19365 (n_7873, n11813);
  not g19366 (n_7874, n11815);
  and g19367 (n11816, n_7873, n_7874);
  not g19368 (n_7875, n11806);
  not g19369 (n_7876, n11816);
  and g19370 (n11817, n_7875, n_7876);
  not g19371 (n_7877, n11817);
  and g19372 (n11818, \asqrt[62] , n_7877);
  and g19376 (n11822, n_7523, n_7522);
  and g19377 (n11823, \asqrt[21] , n11822);
  not g19378 (n_7878, n11823);
  and g19379 (n11824, n_7521, n_7878);
  not g19380 (n_7879, n11821);
  not g19381 (n_7880, n11824);
  and g19382 (n11825, n_7879, n_7880);
  and g19383 (n11826, n_76, n_7875);
  and g19384 (n11827, n_7876, n11826);
  not g19385 (n_7881, n11825);
  not g19386 (n_7882, n11827);
  and g19387 (n11828, n_7881, n_7882);
  not g19388 (n_7883, n11818);
  not g19389 (n_7884, n11828);
  and g19390 (n11829, n_7883, n_7884);
  and g19394 (n11833, n_7531, n_7530);
  and g19395 (n11834, \asqrt[21] , n11833);
  not g19396 (n_7885, n11834);
  and g19397 (n11835, n_7529, n_7885);
  not g19398 (n_7886, n11832);
  not g19399 (n_7887, n11835);
  and g19400 (n11836, n_7886, n_7887);
  and g19401 (n11837, n_7538, n_7537);
  and g19402 (n11838, \asqrt[21] , n11837);
  not g19405 (n_7889, n11836);
  not g19407 (n_7890, n11829);
  not g19409 (n_7891, n11841);
  and g19410 (n11842, n_21, n_7891);
  and g19411 (n11843, n_7883, n11836);
  and g19412 (n11844, n_7884, n11843);
  and g19413 (n11845, n_7537, \asqrt[21] );
  not g19414 (n_7892, n11845);
  and g19415 (n11846, n11305, n_7892);
  not g19416 (n_7893, n11837);
  and g19417 (n11847, \asqrt[63] , n_7893);
  not g19418 (n_7894, n11846);
  and g19419 (n11848, n_7894, n11847);
  not g19425 (n_7895, n11848);
  not g19426 (n_7896, n11853);
  not g19428 (n_7897, n11844);
  and g19432 (n11857, \a[40] , \asqrt[20] );
  not g19433 (n_7902, \a[38] );
  not g19434 (n_7903, \a[39] );
  and g19435 (n11858, n_7902, n_7903);
  and g19436 (n11859, n_7550, n11858);
  not g19437 (n_7904, n11857);
  not g19438 (n_7905, n11859);
  and g19439 (n11860, n_7904, n_7905);
  not g19440 (n_7906, n11860);
  and g19441 (n11861, \asqrt[21] , n_7906);
  and g19447 (n11867, n_7550, \asqrt[20] );
  not g19448 (n_7907, n11867);
  and g19449 (n11868, \a[41] , n_7907);
  and g19450 (n11869, n11334, \asqrt[20] );
  not g19451 (n_7908, n11868);
  not g19452 (n_7909, n11869);
  and g19453 (n11870, n_7908, n_7909);
  not g19454 (n_7910, n11866);
  and g19455 (n11871, n_7910, n11870);
  not g19456 (n_7911, n11861);
  not g19457 (n_7912, n11871);
  and g19458 (n11872, n_7911, n_7912);
  not g19459 (n_7913, n11872);
  and g19460 (n11873, \asqrt[22] , n_7913);
  not g19461 (n_7914, \asqrt[22] );
  and g19462 (n11874, n_7914, n_7911);
  and g19463 (n11875, n_7912, n11874);
  not g19467 (n_7915, n11842);
  not g19469 (n_7916, n11879);
  and g19470 (n11880, n_7909, n_7916);
  not g19471 (n_7917, n11880);
  and g19472 (n11881, \a[42] , n_7917);
  and g19473 (n11882, n_7206, n_7916);
  and g19474 (n11883, n_7909, n11882);
  not g19475 (n_7918, n11881);
  not g19476 (n_7919, n11883);
  and g19477 (n11884, n_7918, n_7919);
  not g19478 (n_7920, n11875);
  not g19479 (n_7921, n11884);
  and g19480 (n11885, n_7920, n_7921);
  not g19481 (n_7922, n11873);
  not g19482 (n_7923, n11885);
  and g19483 (n11886, n_7922, n_7923);
  not g19484 (n_7924, n11886);
  and g19485 (n11887, \asqrt[23] , n_7924);
  and g19486 (n11888, n_7559, n_7558);
  not g19487 (n_7925, n11346);
  and g19488 (n11889, n_7925, n11888);
  and g19489 (n11890, \asqrt[20] , n11889);
  and g19490 (n11891, \asqrt[20] , n11888);
  not g19491 (n_7926, n11891);
  and g19492 (n11892, n11346, n_7926);
  not g19493 (n_7927, n11890);
  not g19494 (n_7928, n11892);
  and g19495 (n11893, n_7927, n_7928);
  and g19496 (n11894, n_7562, n_7922);
  and g19497 (n11895, n_7923, n11894);
  not g19498 (n_7929, n11893);
  not g19499 (n_7930, n11895);
  and g19500 (n11896, n_7929, n_7930);
  not g19501 (n_7931, n11887);
  not g19502 (n_7932, n11896);
  and g19503 (n11897, n_7931, n_7932);
  not g19504 (n_7933, n11897);
  and g19505 (n11898, \asqrt[24] , n_7933);
  and g19509 (n11902, n_7570, n_7568);
  and g19510 (n11903, \asqrt[20] , n11902);
  not g19511 (n_7934, n11903);
  and g19512 (n11904, n_7569, n_7934);
  not g19513 (n_7935, n11901);
  not g19514 (n_7936, n11904);
  and g19515 (n11905, n_7935, n_7936);
  and g19516 (n11906, n_7218, n_7931);
  and g19517 (n11907, n_7932, n11906);
  not g19518 (n_7937, n11905);
  not g19519 (n_7938, n11907);
  and g19520 (n11908, n_7937, n_7938);
  not g19521 (n_7939, n11898);
  not g19522 (n_7940, n11908);
  and g19523 (n11909, n_7939, n_7940);
  not g19524 (n_7941, n11909);
  and g19525 (n11910, \asqrt[25] , n_7941);
  and g19529 (n11914, n_7579, n_7578);
  and g19530 (n11915, \asqrt[20] , n11914);
  not g19531 (n_7942, n11915);
  and g19532 (n11916, n_7577, n_7942);
  not g19533 (n_7943, n11913);
  not g19534 (n_7944, n11916);
  and g19535 (n11917, n_7943, n_7944);
  and g19536 (n11918, n_6882, n_7939);
  and g19537 (n11919, n_7940, n11918);
  not g19538 (n_7945, n11917);
  not g19539 (n_7946, n11919);
  and g19540 (n11920, n_7945, n_7946);
  not g19541 (n_7947, n11910);
  not g19542 (n_7948, n11920);
  and g19543 (n11921, n_7947, n_7948);
  not g19544 (n_7949, n11921);
  and g19545 (n11922, \asqrt[26] , n_7949);
  and g19549 (n11926, n_7587, n_7586);
  and g19550 (n11927, \asqrt[20] , n11926);
  not g19551 (n_7950, n11927);
  and g19552 (n11928, n_7585, n_7950);
  not g19553 (n_7951, n11925);
  not g19554 (n_7952, n11928);
  and g19555 (n11929, n_7951, n_7952);
  and g19556 (n11930, n_6554, n_7947);
  and g19557 (n11931, n_7948, n11930);
  not g19558 (n_7953, n11929);
  not g19559 (n_7954, n11931);
  and g19560 (n11932, n_7953, n_7954);
  not g19561 (n_7955, n11922);
  not g19562 (n_7956, n11932);
  and g19563 (n11933, n_7955, n_7956);
  not g19564 (n_7957, n11933);
  and g19565 (n11934, \asqrt[27] , n_7957);
  and g19569 (n11938, n_7595, n_7594);
  and g19570 (n11939, \asqrt[20] , n11938);
  not g19571 (n_7958, n11939);
  and g19572 (n11940, n_7593, n_7958);
  not g19573 (n_7959, n11937);
  not g19574 (n_7960, n11940);
  and g19575 (n11941, n_7959, n_7960);
  and g19576 (n11942, n_6234, n_7955);
  and g19577 (n11943, n_7956, n11942);
  not g19578 (n_7961, n11941);
  not g19579 (n_7962, n11943);
  and g19580 (n11944, n_7961, n_7962);
  not g19581 (n_7963, n11934);
  not g19582 (n_7964, n11944);
  and g19583 (n11945, n_7963, n_7964);
  not g19584 (n_7965, n11945);
  and g19585 (n11946, \asqrt[28] , n_7965);
  and g19589 (n11950, n_7603, n_7602);
  and g19590 (n11951, \asqrt[20] , n11950);
  not g19591 (n_7966, n11951);
  and g19592 (n11952, n_7601, n_7966);
  not g19593 (n_7967, n11949);
  not g19594 (n_7968, n11952);
  and g19595 (n11953, n_7967, n_7968);
  and g19596 (n11954, n_5922, n_7963);
  and g19597 (n11955, n_7964, n11954);
  not g19598 (n_7969, n11953);
  not g19599 (n_7970, n11955);
  and g19600 (n11956, n_7969, n_7970);
  not g19601 (n_7971, n11946);
  not g19602 (n_7972, n11956);
  and g19603 (n11957, n_7971, n_7972);
  not g19604 (n_7973, n11957);
  and g19605 (n11958, \asqrt[29] , n_7973);
  and g19609 (n11962, n_7611, n_7610);
  and g19610 (n11963, \asqrt[20] , n11962);
  not g19611 (n_7974, n11963);
  and g19612 (n11964, n_7609, n_7974);
  not g19613 (n_7975, n11961);
  not g19614 (n_7976, n11964);
  and g19615 (n11965, n_7975, n_7976);
  and g19616 (n11966, n_5618, n_7971);
  and g19617 (n11967, n_7972, n11966);
  not g19618 (n_7977, n11965);
  not g19619 (n_7978, n11967);
  and g19620 (n11968, n_7977, n_7978);
  not g19621 (n_7979, n11958);
  not g19622 (n_7980, n11968);
  and g19623 (n11969, n_7979, n_7980);
  not g19624 (n_7981, n11969);
  and g19625 (n11970, \asqrt[30] , n_7981);
  and g19629 (n11974, n_7619, n_7618);
  and g19630 (n11975, \asqrt[20] , n11974);
  not g19631 (n_7982, n11975);
  and g19632 (n11976, n_7617, n_7982);
  not g19633 (n_7983, n11973);
  not g19634 (n_7984, n11976);
  and g19635 (n11977, n_7983, n_7984);
  and g19636 (n11978, n_5322, n_7979);
  and g19637 (n11979, n_7980, n11978);
  not g19638 (n_7985, n11977);
  not g19639 (n_7986, n11979);
  and g19640 (n11980, n_7985, n_7986);
  not g19641 (n_7987, n11970);
  not g19642 (n_7988, n11980);
  and g19643 (n11981, n_7987, n_7988);
  not g19644 (n_7989, n11981);
  and g19645 (n11982, \asqrt[31] , n_7989);
  and g19649 (n11986, n_7627, n_7626);
  and g19650 (n11987, \asqrt[20] , n11986);
  not g19651 (n_7990, n11987);
  and g19652 (n11988, n_7625, n_7990);
  not g19653 (n_7991, n11985);
  not g19654 (n_7992, n11988);
  and g19655 (n11989, n_7991, n_7992);
  and g19656 (n11990, n_5034, n_7987);
  and g19657 (n11991, n_7988, n11990);
  not g19658 (n_7993, n11989);
  not g19659 (n_7994, n11991);
  and g19660 (n11992, n_7993, n_7994);
  not g19661 (n_7995, n11982);
  not g19662 (n_7996, n11992);
  and g19663 (n11993, n_7995, n_7996);
  not g19664 (n_7997, n11993);
  and g19665 (n11994, \asqrt[32] , n_7997);
  and g19669 (n11998, n_7635, n_7634);
  and g19670 (n11999, \asqrt[20] , n11998);
  not g19671 (n_7998, n11999);
  and g19672 (n12000, n_7633, n_7998);
  not g19673 (n_7999, n11997);
  not g19674 (n_8000, n12000);
  and g19675 (n12001, n_7999, n_8000);
  and g19676 (n12002, n_4754, n_7995);
  and g19677 (n12003, n_7996, n12002);
  not g19678 (n_8001, n12001);
  not g19679 (n_8002, n12003);
  and g19680 (n12004, n_8001, n_8002);
  not g19681 (n_8003, n11994);
  not g19682 (n_8004, n12004);
  and g19683 (n12005, n_8003, n_8004);
  not g19684 (n_8005, n12005);
  and g19685 (n12006, \asqrt[33] , n_8005);
  and g19689 (n12010, n_7643, n_7642);
  and g19690 (n12011, \asqrt[20] , n12010);
  not g19691 (n_8006, n12011);
  and g19692 (n12012, n_7641, n_8006);
  not g19693 (n_8007, n12009);
  not g19694 (n_8008, n12012);
  and g19695 (n12013, n_8007, n_8008);
  and g19696 (n12014, n_4482, n_8003);
  and g19697 (n12015, n_8004, n12014);
  not g19698 (n_8009, n12013);
  not g19699 (n_8010, n12015);
  and g19700 (n12016, n_8009, n_8010);
  not g19701 (n_8011, n12006);
  not g19702 (n_8012, n12016);
  and g19703 (n12017, n_8011, n_8012);
  not g19704 (n_8013, n12017);
  and g19705 (n12018, \asqrt[34] , n_8013);
  and g19709 (n12022, n_7651, n_7650);
  and g19710 (n12023, \asqrt[20] , n12022);
  not g19711 (n_8014, n12023);
  and g19712 (n12024, n_7649, n_8014);
  not g19713 (n_8015, n12021);
  not g19714 (n_8016, n12024);
  and g19715 (n12025, n_8015, n_8016);
  and g19716 (n12026, n_4218, n_8011);
  and g19717 (n12027, n_8012, n12026);
  not g19718 (n_8017, n12025);
  not g19719 (n_8018, n12027);
  and g19720 (n12028, n_8017, n_8018);
  not g19721 (n_8019, n12018);
  not g19722 (n_8020, n12028);
  and g19723 (n12029, n_8019, n_8020);
  not g19724 (n_8021, n12029);
  and g19725 (n12030, \asqrt[35] , n_8021);
  and g19729 (n12034, n_7659, n_7658);
  and g19730 (n12035, \asqrt[20] , n12034);
  not g19731 (n_8022, n12035);
  and g19732 (n12036, n_7657, n_8022);
  not g19733 (n_8023, n12033);
  not g19734 (n_8024, n12036);
  and g19735 (n12037, n_8023, n_8024);
  and g19736 (n12038, n_3962, n_8019);
  and g19737 (n12039, n_8020, n12038);
  not g19738 (n_8025, n12037);
  not g19739 (n_8026, n12039);
  and g19740 (n12040, n_8025, n_8026);
  not g19741 (n_8027, n12030);
  not g19742 (n_8028, n12040);
  and g19743 (n12041, n_8027, n_8028);
  not g19744 (n_8029, n12041);
  and g19745 (n12042, \asqrt[36] , n_8029);
  and g19749 (n12046, n_7667, n_7666);
  and g19750 (n12047, \asqrt[20] , n12046);
  not g19751 (n_8030, n12047);
  and g19752 (n12048, n_7665, n_8030);
  not g19753 (n_8031, n12045);
  not g19754 (n_8032, n12048);
  and g19755 (n12049, n_8031, n_8032);
  and g19756 (n12050, n_3714, n_8027);
  and g19757 (n12051, n_8028, n12050);
  not g19758 (n_8033, n12049);
  not g19759 (n_8034, n12051);
  and g19760 (n12052, n_8033, n_8034);
  not g19761 (n_8035, n12042);
  not g19762 (n_8036, n12052);
  and g19763 (n12053, n_8035, n_8036);
  not g19764 (n_8037, n12053);
  and g19765 (n12054, \asqrt[37] , n_8037);
  and g19769 (n12058, n_7675, n_7674);
  and g19770 (n12059, \asqrt[20] , n12058);
  not g19771 (n_8038, n12059);
  and g19772 (n12060, n_7673, n_8038);
  not g19773 (n_8039, n12057);
  not g19774 (n_8040, n12060);
  and g19775 (n12061, n_8039, n_8040);
  and g19776 (n12062, n_3474, n_8035);
  and g19777 (n12063, n_8036, n12062);
  not g19778 (n_8041, n12061);
  not g19779 (n_8042, n12063);
  and g19780 (n12064, n_8041, n_8042);
  not g19781 (n_8043, n12054);
  not g19782 (n_8044, n12064);
  and g19783 (n12065, n_8043, n_8044);
  not g19784 (n_8045, n12065);
  and g19785 (n12066, \asqrt[38] , n_8045);
  and g19789 (n12070, n_7683, n_7682);
  and g19790 (n12071, \asqrt[20] , n12070);
  not g19791 (n_8046, n12071);
  and g19792 (n12072, n_7681, n_8046);
  not g19793 (n_8047, n12069);
  not g19794 (n_8048, n12072);
  and g19795 (n12073, n_8047, n_8048);
  and g19796 (n12074, n_3242, n_8043);
  and g19797 (n12075, n_8044, n12074);
  not g19798 (n_8049, n12073);
  not g19799 (n_8050, n12075);
  and g19800 (n12076, n_8049, n_8050);
  not g19801 (n_8051, n12066);
  not g19802 (n_8052, n12076);
  and g19803 (n12077, n_8051, n_8052);
  not g19804 (n_8053, n12077);
  and g19805 (n12078, \asqrt[39] , n_8053);
  and g19809 (n12082, n_7691, n_7690);
  and g19810 (n12083, \asqrt[20] , n12082);
  not g19811 (n_8054, n12083);
  and g19812 (n12084, n_7689, n_8054);
  not g19813 (n_8055, n12081);
  not g19814 (n_8056, n12084);
  and g19815 (n12085, n_8055, n_8056);
  and g19816 (n12086, n_3018, n_8051);
  and g19817 (n12087, n_8052, n12086);
  not g19818 (n_8057, n12085);
  not g19819 (n_8058, n12087);
  and g19820 (n12088, n_8057, n_8058);
  not g19821 (n_8059, n12078);
  not g19822 (n_8060, n12088);
  and g19823 (n12089, n_8059, n_8060);
  not g19824 (n_8061, n12089);
  and g19825 (n12090, \asqrt[40] , n_8061);
  and g19829 (n12094, n_7699, n_7698);
  and g19830 (n12095, \asqrt[20] , n12094);
  not g19831 (n_8062, n12095);
  and g19832 (n12096, n_7697, n_8062);
  not g19833 (n_8063, n12093);
  not g19834 (n_8064, n12096);
  and g19835 (n12097, n_8063, n_8064);
  and g19836 (n12098, n_2802, n_8059);
  and g19837 (n12099, n_8060, n12098);
  not g19838 (n_8065, n12097);
  not g19839 (n_8066, n12099);
  and g19840 (n12100, n_8065, n_8066);
  not g19841 (n_8067, n12090);
  not g19842 (n_8068, n12100);
  and g19843 (n12101, n_8067, n_8068);
  not g19844 (n_8069, n12101);
  and g19845 (n12102, \asqrt[41] , n_8069);
  and g19849 (n12106, n_7707, n_7706);
  and g19850 (n12107, \asqrt[20] , n12106);
  not g19851 (n_8070, n12107);
  and g19852 (n12108, n_7705, n_8070);
  not g19853 (n_8071, n12105);
  not g19854 (n_8072, n12108);
  and g19855 (n12109, n_8071, n_8072);
  and g19856 (n12110, n_2594, n_8067);
  and g19857 (n12111, n_8068, n12110);
  not g19858 (n_8073, n12109);
  not g19859 (n_8074, n12111);
  and g19860 (n12112, n_8073, n_8074);
  not g19861 (n_8075, n12102);
  not g19862 (n_8076, n12112);
  and g19863 (n12113, n_8075, n_8076);
  not g19864 (n_8077, n12113);
  and g19865 (n12114, \asqrt[42] , n_8077);
  and g19869 (n12118, n_7715, n_7714);
  and g19870 (n12119, \asqrt[20] , n12118);
  not g19871 (n_8078, n12119);
  and g19872 (n12120, n_7713, n_8078);
  not g19873 (n_8079, n12117);
  not g19874 (n_8080, n12120);
  and g19875 (n12121, n_8079, n_8080);
  and g19876 (n12122, n_2394, n_8075);
  and g19877 (n12123, n_8076, n12122);
  not g19878 (n_8081, n12121);
  not g19879 (n_8082, n12123);
  and g19880 (n12124, n_8081, n_8082);
  not g19881 (n_8083, n12114);
  not g19882 (n_8084, n12124);
  and g19883 (n12125, n_8083, n_8084);
  not g19884 (n_8085, n12125);
  and g19885 (n12126, \asqrt[43] , n_8085);
  and g19889 (n12130, n_7723, n_7722);
  and g19890 (n12131, \asqrt[20] , n12130);
  not g19891 (n_8086, n12131);
  and g19892 (n12132, n_7721, n_8086);
  not g19893 (n_8087, n12129);
  not g19894 (n_8088, n12132);
  and g19895 (n12133, n_8087, n_8088);
  and g19896 (n12134, n_2202, n_8083);
  and g19897 (n12135, n_8084, n12134);
  not g19898 (n_8089, n12133);
  not g19899 (n_8090, n12135);
  and g19900 (n12136, n_8089, n_8090);
  not g19901 (n_8091, n12126);
  not g19902 (n_8092, n12136);
  and g19903 (n12137, n_8091, n_8092);
  not g19904 (n_8093, n12137);
  and g19905 (n12138, \asqrt[44] , n_8093);
  and g19909 (n12142, n_7731, n_7730);
  and g19910 (n12143, \asqrt[20] , n12142);
  not g19911 (n_8094, n12143);
  and g19912 (n12144, n_7729, n_8094);
  not g19913 (n_8095, n12141);
  not g19914 (n_8096, n12144);
  and g19915 (n12145, n_8095, n_8096);
  and g19916 (n12146, n_2018, n_8091);
  and g19917 (n12147, n_8092, n12146);
  not g19918 (n_8097, n12145);
  not g19919 (n_8098, n12147);
  and g19920 (n12148, n_8097, n_8098);
  not g19921 (n_8099, n12138);
  not g19922 (n_8100, n12148);
  and g19923 (n12149, n_8099, n_8100);
  not g19924 (n_8101, n12149);
  and g19925 (n12150, \asqrt[45] , n_8101);
  and g19926 (n12151, n_1842, n_8099);
  and g19927 (n12152, n_8100, n12151);
  and g19931 (n12156, n_7739, n_7737);
  and g19932 (n12157, \asqrt[20] , n12156);
  not g19933 (n_8102, n12157);
  and g19934 (n12158, n_7738, n_8102);
  not g19935 (n_8103, n12155);
  not g19936 (n_8104, n12158);
  and g19937 (n12159, n_8103, n_8104);
  not g19938 (n_8105, n12152);
  not g19939 (n_8106, n12159);
  and g19940 (n12160, n_8105, n_8106);
  not g19941 (n_8107, n12150);
  not g19942 (n_8108, n12160);
  and g19943 (n12161, n_8107, n_8108);
  not g19944 (n_8109, n12161);
  and g19945 (n12162, \asqrt[46] , n_8109);
  and g19949 (n12166, n_7747, n_7746);
  and g19950 (n12167, \asqrt[20] , n12166);
  not g19951 (n_8110, n12167);
  and g19952 (n12168, n_7745, n_8110);
  not g19953 (n_8111, n12165);
  not g19954 (n_8112, n12168);
  and g19955 (n12169, n_8111, n_8112);
  and g19956 (n12170, n_1674, n_8107);
  and g19957 (n12171, n_8108, n12170);
  not g19958 (n_8113, n12169);
  not g19959 (n_8114, n12171);
  and g19960 (n12172, n_8113, n_8114);
  not g19961 (n_8115, n12162);
  not g19962 (n_8116, n12172);
  and g19963 (n12173, n_8115, n_8116);
  not g19964 (n_8117, n12173);
  and g19965 (n12174, \asqrt[47] , n_8117);
  and g19969 (n12178, n_7755, n_7754);
  and g19970 (n12179, \asqrt[20] , n12178);
  not g19971 (n_8118, n12179);
  and g19972 (n12180, n_7753, n_8118);
  not g19973 (n_8119, n12177);
  not g19974 (n_8120, n12180);
  and g19975 (n12181, n_8119, n_8120);
  and g19976 (n12182, n_1514, n_8115);
  and g19977 (n12183, n_8116, n12182);
  not g19978 (n_8121, n12181);
  not g19979 (n_8122, n12183);
  and g19980 (n12184, n_8121, n_8122);
  not g19981 (n_8123, n12174);
  not g19982 (n_8124, n12184);
  and g19983 (n12185, n_8123, n_8124);
  not g19984 (n_8125, n12185);
  and g19985 (n12186, \asqrt[48] , n_8125);
  and g19989 (n12190, n_7763, n_7762);
  and g19990 (n12191, \asqrt[20] , n12190);
  not g19991 (n_8126, n12191);
  and g19992 (n12192, n_7761, n_8126);
  not g19993 (n_8127, n12189);
  not g19994 (n_8128, n12192);
  and g19995 (n12193, n_8127, n_8128);
  and g19996 (n12194, n_1362, n_8123);
  and g19997 (n12195, n_8124, n12194);
  not g19998 (n_8129, n12193);
  not g19999 (n_8130, n12195);
  and g20000 (n12196, n_8129, n_8130);
  not g20001 (n_8131, n12186);
  not g20002 (n_8132, n12196);
  and g20003 (n12197, n_8131, n_8132);
  not g20004 (n_8133, n12197);
  and g20005 (n12198, \asqrt[49] , n_8133);
  and g20009 (n12202, n_7771, n_7770);
  and g20010 (n12203, \asqrt[20] , n12202);
  not g20011 (n_8134, n12203);
  and g20012 (n12204, n_7769, n_8134);
  not g20013 (n_8135, n12201);
  not g20014 (n_8136, n12204);
  and g20015 (n12205, n_8135, n_8136);
  and g20016 (n12206, n_1218, n_8131);
  and g20017 (n12207, n_8132, n12206);
  not g20018 (n_8137, n12205);
  not g20019 (n_8138, n12207);
  and g20020 (n12208, n_8137, n_8138);
  not g20021 (n_8139, n12198);
  not g20022 (n_8140, n12208);
  and g20023 (n12209, n_8139, n_8140);
  not g20024 (n_8141, n12209);
  and g20025 (n12210, \asqrt[50] , n_8141);
  and g20029 (n12214, n_7779, n_7778);
  and g20030 (n12215, \asqrt[20] , n12214);
  not g20031 (n_8142, n12215);
  and g20032 (n12216, n_7777, n_8142);
  not g20033 (n_8143, n12213);
  not g20034 (n_8144, n12216);
  and g20035 (n12217, n_8143, n_8144);
  and g20036 (n12218, n_1082, n_8139);
  and g20037 (n12219, n_8140, n12218);
  not g20038 (n_8145, n12217);
  not g20039 (n_8146, n12219);
  and g20040 (n12220, n_8145, n_8146);
  not g20041 (n_8147, n12210);
  not g20042 (n_8148, n12220);
  and g20043 (n12221, n_8147, n_8148);
  not g20044 (n_8149, n12221);
  and g20045 (n12222, \asqrt[51] , n_8149);
  and g20049 (n12226, n_7787, n_7786);
  and g20050 (n12227, \asqrt[20] , n12226);
  not g20051 (n_8150, n12227);
  and g20052 (n12228, n_7785, n_8150);
  not g20053 (n_8151, n12225);
  not g20054 (n_8152, n12228);
  and g20055 (n12229, n_8151, n_8152);
  and g20056 (n12230, n_954, n_8147);
  and g20057 (n12231, n_8148, n12230);
  not g20058 (n_8153, n12229);
  not g20059 (n_8154, n12231);
  and g20060 (n12232, n_8153, n_8154);
  not g20061 (n_8155, n12222);
  not g20062 (n_8156, n12232);
  and g20063 (n12233, n_8155, n_8156);
  not g20064 (n_8157, n12233);
  and g20065 (n12234, \asqrt[52] , n_8157);
  and g20069 (n12238, n_7795, n_7794);
  and g20070 (n12239, \asqrt[20] , n12238);
  not g20071 (n_8158, n12239);
  and g20072 (n12240, n_7793, n_8158);
  not g20073 (n_8159, n12237);
  not g20074 (n_8160, n12240);
  and g20075 (n12241, n_8159, n_8160);
  and g20076 (n12242, n_834, n_8155);
  and g20077 (n12243, n_8156, n12242);
  not g20078 (n_8161, n12241);
  not g20079 (n_8162, n12243);
  and g20080 (n12244, n_8161, n_8162);
  not g20081 (n_8163, n12234);
  not g20082 (n_8164, n12244);
  and g20083 (n12245, n_8163, n_8164);
  not g20084 (n_8165, n12245);
  and g20085 (n12246, \asqrt[53] , n_8165);
  and g20089 (n12250, n_7803, n_7802);
  and g20090 (n12251, \asqrt[20] , n12250);
  not g20091 (n_8166, n12251);
  and g20092 (n12252, n_7801, n_8166);
  not g20093 (n_8167, n12249);
  not g20094 (n_8168, n12252);
  and g20095 (n12253, n_8167, n_8168);
  and g20096 (n12254, n_722, n_8163);
  and g20097 (n12255, n_8164, n12254);
  not g20098 (n_8169, n12253);
  not g20099 (n_8170, n12255);
  and g20100 (n12256, n_8169, n_8170);
  not g20101 (n_8171, n12246);
  not g20102 (n_8172, n12256);
  and g20103 (n12257, n_8171, n_8172);
  not g20104 (n_8173, n12257);
  and g20105 (n12258, \asqrt[54] , n_8173);
  and g20109 (n12262, n_7811, n_7810);
  and g20110 (n12263, \asqrt[20] , n12262);
  not g20111 (n_8174, n12263);
  and g20112 (n12264, n_7809, n_8174);
  not g20113 (n_8175, n12261);
  not g20114 (n_8176, n12264);
  and g20115 (n12265, n_8175, n_8176);
  and g20116 (n12266, n_618, n_8171);
  and g20117 (n12267, n_8172, n12266);
  not g20118 (n_8177, n12265);
  not g20119 (n_8178, n12267);
  and g20120 (n12268, n_8177, n_8178);
  not g20121 (n_8179, n12258);
  not g20122 (n_8180, n12268);
  and g20123 (n12269, n_8179, n_8180);
  not g20124 (n_8181, n12269);
  and g20125 (n12270, \asqrt[55] , n_8181);
  and g20129 (n12274, n_7819, n_7818);
  and g20130 (n12275, \asqrt[20] , n12274);
  not g20131 (n_8182, n12275);
  and g20132 (n12276, n_7817, n_8182);
  not g20133 (n_8183, n12273);
  not g20134 (n_8184, n12276);
  and g20135 (n12277, n_8183, n_8184);
  and g20136 (n12278, n_522, n_8179);
  and g20137 (n12279, n_8180, n12278);
  not g20138 (n_8185, n12277);
  not g20139 (n_8186, n12279);
  and g20140 (n12280, n_8185, n_8186);
  not g20141 (n_8187, n12270);
  not g20142 (n_8188, n12280);
  and g20143 (n12281, n_8187, n_8188);
  not g20144 (n_8189, n12281);
  and g20145 (n12282, \asqrt[56] , n_8189);
  and g20149 (n12286, n_7827, n_7826);
  and g20150 (n12287, \asqrt[20] , n12286);
  not g20151 (n_8190, n12287);
  and g20152 (n12288, n_7825, n_8190);
  not g20153 (n_8191, n12285);
  not g20154 (n_8192, n12288);
  and g20155 (n12289, n_8191, n_8192);
  and g20156 (n12290, n_434, n_8187);
  and g20157 (n12291, n_8188, n12290);
  not g20158 (n_8193, n12289);
  not g20159 (n_8194, n12291);
  and g20160 (n12292, n_8193, n_8194);
  not g20161 (n_8195, n12282);
  not g20162 (n_8196, n12292);
  and g20163 (n12293, n_8195, n_8196);
  not g20164 (n_8197, n12293);
  and g20165 (n12294, \asqrt[57] , n_8197);
  and g20169 (n12298, n_7835, n_7834);
  and g20170 (n12299, \asqrt[20] , n12298);
  not g20171 (n_8198, n12299);
  and g20172 (n12300, n_7833, n_8198);
  not g20173 (n_8199, n12297);
  not g20174 (n_8200, n12300);
  and g20175 (n12301, n_8199, n_8200);
  and g20176 (n12302, n_354, n_8195);
  and g20177 (n12303, n_8196, n12302);
  not g20178 (n_8201, n12301);
  not g20179 (n_8202, n12303);
  and g20180 (n12304, n_8201, n_8202);
  not g20181 (n_8203, n12294);
  not g20182 (n_8204, n12304);
  and g20183 (n12305, n_8203, n_8204);
  not g20184 (n_8205, n12305);
  and g20185 (n12306, \asqrt[58] , n_8205);
  and g20189 (n12310, n_7843, n_7842);
  and g20190 (n12311, \asqrt[20] , n12310);
  not g20191 (n_8206, n12311);
  and g20192 (n12312, n_7841, n_8206);
  not g20193 (n_8207, n12309);
  not g20194 (n_8208, n12312);
  and g20195 (n12313, n_8207, n_8208);
  and g20196 (n12314, n_282, n_8203);
  and g20197 (n12315, n_8204, n12314);
  not g20198 (n_8209, n12313);
  not g20199 (n_8210, n12315);
  and g20200 (n12316, n_8209, n_8210);
  not g20201 (n_8211, n12306);
  not g20202 (n_8212, n12316);
  and g20203 (n12317, n_8211, n_8212);
  not g20204 (n_8213, n12317);
  and g20205 (n12318, \asqrt[59] , n_8213);
  and g20209 (n12322, n_7851, n_7850);
  and g20210 (n12323, \asqrt[20] , n12322);
  not g20211 (n_8214, n12323);
  and g20212 (n12324, n_7849, n_8214);
  not g20213 (n_8215, n12321);
  not g20214 (n_8216, n12324);
  and g20215 (n12325, n_8215, n_8216);
  and g20216 (n12326, n_218, n_8211);
  and g20217 (n12327, n_8212, n12326);
  not g20218 (n_8217, n12325);
  not g20219 (n_8218, n12327);
  and g20220 (n12328, n_8217, n_8218);
  not g20221 (n_8219, n12318);
  not g20222 (n_8220, n12328);
  and g20223 (n12329, n_8219, n_8220);
  not g20224 (n_8221, n12329);
  and g20225 (n12330, \asqrt[60] , n_8221);
  and g20229 (n12334, n_7859, n_7858);
  and g20230 (n12335, \asqrt[20] , n12334);
  not g20231 (n_8222, n12335);
  and g20232 (n12336, n_7857, n_8222);
  not g20233 (n_8223, n12333);
  not g20234 (n_8224, n12336);
  and g20235 (n12337, n_8223, n_8224);
  and g20236 (n12338, n_162, n_8219);
  and g20237 (n12339, n_8220, n12338);
  not g20238 (n_8225, n12337);
  not g20239 (n_8226, n12339);
  and g20240 (n12340, n_8225, n_8226);
  not g20241 (n_8227, n12330);
  not g20242 (n_8228, n12340);
  and g20243 (n12341, n_8227, n_8228);
  not g20244 (n_8229, n12341);
  and g20245 (n12342, \asqrt[61] , n_8229);
  and g20249 (n12346, n_7867, n_7866);
  and g20250 (n12347, \asqrt[20] , n12346);
  not g20251 (n_8230, n12347);
  and g20252 (n12348, n_7865, n_8230);
  not g20253 (n_8231, n12345);
  not g20254 (n_8232, n12348);
  and g20255 (n12349, n_8231, n_8232);
  and g20256 (n12350, n_115, n_8227);
  and g20257 (n12351, n_8228, n12350);
  not g20258 (n_8233, n12349);
  not g20259 (n_8234, n12351);
  and g20260 (n12352, n_8233, n_8234);
  not g20261 (n_8235, n12342);
  not g20262 (n_8236, n12352);
  and g20263 (n12353, n_8235, n_8236);
  not g20264 (n_8237, n12353);
  and g20265 (n12354, \asqrt[62] , n_8237);
  and g20269 (n12358, n_7875, n_7874);
  and g20270 (n12359, \asqrt[20] , n12358);
  not g20271 (n_8238, n12359);
  and g20272 (n12360, n_7873, n_8238);
  not g20273 (n_8239, n12357);
  not g20274 (n_8240, n12360);
  and g20275 (n12361, n_8239, n_8240);
  and g20276 (n12362, n_76, n_8235);
  and g20277 (n12363, n_8236, n12362);
  not g20278 (n_8241, n12361);
  not g20279 (n_8242, n12363);
  and g20280 (n12364, n_8241, n_8242);
  not g20281 (n_8243, n12354);
  not g20282 (n_8244, n12364);
  and g20283 (n12365, n_8243, n_8244);
  and g20287 (n12369, n_7883, n_7882);
  and g20288 (n12370, \asqrt[20] , n12369);
  not g20289 (n_8245, n12370);
  and g20290 (n12371, n_7881, n_8245);
  not g20291 (n_8246, n12368);
  not g20292 (n_8247, n12371);
  and g20293 (n12372, n_8246, n_8247);
  and g20294 (n12373, n_7890, n_7889);
  and g20295 (n12374, \asqrt[20] , n12373);
  not g20298 (n_8249, n12372);
  not g20300 (n_8250, n12365);
  not g20302 (n_8251, n12377);
  and g20303 (n12378, n_21, n_8251);
  and g20304 (n12379, n_8243, n12372);
  and g20305 (n12380, n_8244, n12379);
  and g20306 (n12381, n_7889, \asqrt[20] );
  not g20307 (n_8252, n12381);
  and g20308 (n12382, n11829, n_8252);
  not g20309 (n_8253, n12373);
  and g20310 (n12383, \asqrt[63] , n_8253);
  not g20311 (n_8254, n12382);
  and g20312 (n12384, n_8254, n12383);
  not g20318 (n_8255, n12384);
  not g20319 (n_8256, n12389);
  not g20321 (n_8257, n12380);
  and g20325 (n12393, \a[38] , \asqrt[19] );
  not g20326 (n_8262, \a[36] );
  not g20327 (n_8263, \a[37] );
  and g20328 (n12394, n_8262, n_8263);
  and g20329 (n12395, n_7902, n12394);
  not g20330 (n_8264, n12393);
  not g20331 (n_8265, n12395);
  and g20332 (n12396, n_8264, n_8265);
  not g20333 (n_8266, n12396);
  and g20334 (n12397, \asqrt[20] , n_8266);
  and g20340 (n12403, n_7902, \asqrt[19] );
  not g20341 (n_8267, n12403);
  and g20342 (n12404, \a[39] , n_8267);
  and g20343 (n12405, n11858, \asqrt[19] );
  not g20344 (n_8268, n12404);
  not g20345 (n_8269, n12405);
  and g20346 (n12406, n_8268, n_8269);
  not g20347 (n_8270, n12402);
  and g20348 (n12407, n_8270, n12406);
  not g20349 (n_8271, n12397);
  not g20350 (n_8272, n12407);
  and g20351 (n12408, n_8271, n_8272);
  not g20352 (n_8273, n12408);
  and g20353 (n12409, \asqrt[21] , n_8273);
  not g20354 (n_8274, \asqrt[21] );
  and g20355 (n12410, n_8274, n_8271);
  and g20356 (n12411, n_8272, n12410);
  not g20360 (n_8275, n12378);
  not g20362 (n_8276, n12415);
  and g20363 (n12416, n_8269, n_8276);
  not g20364 (n_8277, n12416);
  and g20365 (n12417, \a[40] , n_8277);
  and g20366 (n12418, n_7550, n_8276);
  and g20367 (n12419, n_8269, n12418);
  not g20368 (n_8278, n12417);
  not g20369 (n_8279, n12419);
  and g20370 (n12420, n_8278, n_8279);
  not g20371 (n_8280, n12411);
  not g20372 (n_8281, n12420);
  and g20373 (n12421, n_8280, n_8281);
  not g20374 (n_8282, n12409);
  not g20375 (n_8283, n12421);
  and g20376 (n12422, n_8282, n_8283);
  not g20377 (n_8284, n12422);
  and g20378 (n12423, \asqrt[22] , n_8284);
  and g20379 (n12424, n_7911, n_7910);
  not g20380 (n_8285, n11870);
  and g20381 (n12425, n_8285, n12424);
  and g20382 (n12426, \asqrt[19] , n12425);
  and g20383 (n12427, \asqrt[19] , n12424);
  not g20384 (n_8286, n12427);
  and g20385 (n12428, n11870, n_8286);
  not g20386 (n_8287, n12426);
  not g20387 (n_8288, n12428);
  and g20388 (n12429, n_8287, n_8288);
  and g20389 (n12430, n_7914, n_8282);
  and g20390 (n12431, n_8283, n12430);
  not g20391 (n_8289, n12429);
  not g20392 (n_8290, n12431);
  and g20393 (n12432, n_8289, n_8290);
  not g20394 (n_8291, n12423);
  not g20395 (n_8292, n12432);
  and g20396 (n12433, n_8291, n_8292);
  not g20397 (n_8293, n12433);
  and g20398 (n12434, \asqrt[23] , n_8293);
  and g20402 (n12438, n_7922, n_7920);
  and g20403 (n12439, \asqrt[19] , n12438);
  not g20404 (n_8294, n12439);
  and g20405 (n12440, n_7921, n_8294);
  not g20406 (n_8295, n12437);
  not g20407 (n_8296, n12440);
  and g20408 (n12441, n_8295, n_8296);
  and g20409 (n12442, n_7562, n_8291);
  and g20410 (n12443, n_8292, n12442);
  not g20411 (n_8297, n12441);
  not g20412 (n_8298, n12443);
  and g20413 (n12444, n_8297, n_8298);
  not g20414 (n_8299, n12434);
  not g20415 (n_8300, n12444);
  and g20416 (n12445, n_8299, n_8300);
  not g20417 (n_8301, n12445);
  and g20418 (n12446, \asqrt[24] , n_8301);
  and g20422 (n12450, n_7931, n_7930);
  and g20423 (n12451, \asqrt[19] , n12450);
  not g20424 (n_8302, n12451);
  and g20425 (n12452, n_7929, n_8302);
  not g20426 (n_8303, n12449);
  not g20427 (n_8304, n12452);
  and g20428 (n12453, n_8303, n_8304);
  and g20429 (n12454, n_7218, n_8299);
  and g20430 (n12455, n_8300, n12454);
  not g20431 (n_8305, n12453);
  not g20432 (n_8306, n12455);
  and g20433 (n12456, n_8305, n_8306);
  not g20434 (n_8307, n12446);
  not g20435 (n_8308, n12456);
  and g20436 (n12457, n_8307, n_8308);
  not g20437 (n_8309, n12457);
  and g20438 (n12458, \asqrt[25] , n_8309);
  and g20442 (n12462, n_7939, n_7938);
  and g20443 (n12463, \asqrt[19] , n12462);
  not g20444 (n_8310, n12463);
  and g20445 (n12464, n_7937, n_8310);
  not g20446 (n_8311, n12461);
  not g20447 (n_8312, n12464);
  and g20448 (n12465, n_8311, n_8312);
  and g20449 (n12466, n_6882, n_8307);
  and g20450 (n12467, n_8308, n12466);
  not g20451 (n_8313, n12465);
  not g20452 (n_8314, n12467);
  and g20453 (n12468, n_8313, n_8314);
  not g20454 (n_8315, n12458);
  not g20455 (n_8316, n12468);
  and g20456 (n12469, n_8315, n_8316);
  not g20457 (n_8317, n12469);
  and g20458 (n12470, \asqrt[26] , n_8317);
  and g20462 (n12474, n_7947, n_7946);
  and g20463 (n12475, \asqrt[19] , n12474);
  not g20464 (n_8318, n12475);
  and g20465 (n12476, n_7945, n_8318);
  not g20466 (n_8319, n12473);
  not g20467 (n_8320, n12476);
  and g20468 (n12477, n_8319, n_8320);
  and g20469 (n12478, n_6554, n_8315);
  and g20470 (n12479, n_8316, n12478);
  not g20471 (n_8321, n12477);
  not g20472 (n_8322, n12479);
  and g20473 (n12480, n_8321, n_8322);
  not g20474 (n_8323, n12470);
  not g20475 (n_8324, n12480);
  and g20476 (n12481, n_8323, n_8324);
  not g20477 (n_8325, n12481);
  and g20478 (n12482, \asqrt[27] , n_8325);
  and g20482 (n12486, n_7955, n_7954);
  and g20483 (n12487, \asqrt[19] , n12486);
  not g20484 (n_8326, n12487);
  and g20485 (n12488, n_7953, n_8326);
  not g20486 (n_8327, n12485);
  not g20487 (n_8328, n12488);
  and g20488 (n12489, n_8327, n_8328);
  and g20489 (n12490, n_6234, n_8323);
  and g20490 (n12491, n_8324, n12490);
  not g20491 (n_8329, n12489);
  not g20492 (n_8330, n12491);
  and g20493 (n12492, n_8329, n_8330);
  not g20494 (n_8331, n12482);
  not g20495 (n_8332, n12492);
  and g20496 (n12493, n_8331, n_8332);
  not g20497 (n_8333, n12493);
  and g20498 (n12494, \asqrt[28] , n_8333);
  and g20502 (n12498, n_7963, n_7962);
  and g20503 (n12499, \asqrt[19] , n12498);
  not g20504 (n_8334, n12499);
  and g20505 (n12500, n_7961, n_8334);
  not g20506 (n_8335, n12497);
  not g20507 (n_8336, n12500);
  and g20508 (n12501, n_8335, n_8336);
  and g20509 (n12502, n_5922, n_8331);
  and g20510 (n12503, n_8332, n12502);
  not g20511 (n_8337, n12501);
  not g20512 (n_8338, n12503);
  and g20513 (n12504, n_8337, n_8338);
  not g20514 (n_8339, n12494);
  not g20515 (n_8340, n12504);
  and g20516 (n12505, n_8339, n_8340);
  not g20517 (n_8341, n12505);
  and g20518 (n12506, \asqrt[29] , n_8341);
  and g20522 (n12510, n_7971, n_7970);
  and g20523 (n12511, \asqrt[19] , n12510);
  not g20524 (n_8342, n12511);
  and g20525 (n12512, n_7969, n_8342);
  not g20526 (n_8343, n12509);
  not g20527 (n_8344, n12512);
  and g20528 (n12513, n_8343, n_8344);
  and g20529 (n12514, n_5618, n_8339);
  and g20530 (n12515, n_8340, n12514);
  not g20531 (n_8345, n12513);
  not g20532 (n_8346, n12515);
  and g20533 (n12516, n_8345, n_8346);
  not g20534 (n_8347, n12506);
  not g20535 (n_8348, n12516);
  and g20536 (n12517, n_8347, n_8348);
  not g20537 (n_8349, n12517);
  and g20538 (n12518, \asqrt[30] , n_8349);
  and g20542 (n12522, n_7979, n_7978);
  and g20543 (n12523, \asqrt[19] , n12522);
  not g20544 (n_8350, n12523);
  and g20545 (n12524, n_7977, n_8350);
  not g20546 (n_8351, n12521);
  not g20547 (n_8352, n12524);
  and g20548 (n12525, n_8351, n_8352);
  and g20549 (n12526, n_5322, n_8347);
  and g20550 (n12527, n_8348, n12526);
  not g20551 (n_8353, n12525);
  not g20552 (n_8354, n12527);
  and g20553 (n12528, n_8353, n_8354);
  not g20554 (n_8355, n12518);
  not g20555 (n_8356, n12528);
  and g20556 (n12529, n_8355, n_8356);
  not g20557 (n_8357, n12529);
  and g20558 (n12530, \asqrt[31] , n_8357);
  and g20562 (n12534, n_7987, n_7986);
  and g20563 (n12535, \asqrt[19] , n12534);
  not g20564 (n_8358, n12535);
  and g20565 (n12536, n_7985, n_8358);
  not g20566 (n_8359, n12533);
  not g20567 (n_8360, n12536);
  and g20568 (n12537, n_8359, n_8360);
  and g20569 (n12538, n_5034, n_8355);
  and g20570 (n12539, n_8356, n12538);
  not g20571 (n_8361, n12537);
  not g20572 (n_8362, n12539);
  and g20573 (n12540, n_8361, n_8362);
  not g20574 (n_8363, n12530);
  not g20575 (n_8364, n12540);
  and g20576 (n12541, n_8363, n_8364);
  not g20577 (n_8365, n12541);
  and g20578 (n12542, \asqrt[32] , n_8365);
  and g20582 (n12546, n_7995, n_7994);
  and g20583 (n12547, \asqrt[19] , n12546);
  not g20584 (n_8366, n12547);
  and g20585 (n12548, n_7993, n_8366);
  not g20586 (n_8367, n12545);
  not g20587 (n_8368, n12548);
  and g20588 (n12549, n_8367, n_8368);
  and g20589 (n12550, n_4754, n_8363);
  and g20590 (n12551, n_8364, n12550);
  not g20591 (n_8369, n12549);
  not g20592 (n_8370, n12551);
  and g20593 (n12552, n_8369, n_8370);
  not g20594 (n_8371, n12542);
  not g20595 (n_8372, n12552);
  and g20596 (n12553, n_8371, n_8372);
  not g20597 (n_8373, n12553);
  and g20598 (n12554, \asqrt[33] , n_8373);
  and g20602 (n12558, n_8003, n_8002);
  and g20603 (n12559, \asqrt[19] , n12558);
  not g20604 (n_8374, n12559);
  and g20605 (n12560, n_8001, n_8374);
  not g20606 (n_8375, n12557);
  not g20607 (n_8376, n12560);
  and g20608 (n12561, n_8375, n_8376);
  and g20609 (n12562, n_4482, n_8371);
  and g20610 (n12563, n_8372, n12562);
  not g20611 (n_8377, n12561);
  not g20612 (n_8378, n12563);
  and g20613 (n12564, n_8377, n_8378);
  not g20614 (n_8379, n12554);
  not g20615 (n_8380, n12564);
  and g20616 (n12565, n_8379, n_8380);
  not g20617 (n_8381, n12565);
  and g20618 (n12566, \asqrt[34] , n_8381);
  and g20622 (n12570, n_8011, n_8010);
  and g20623 (n12571, \asqrt[19] , n12570);
  not g20624 (n_8382, n12571);
  and g20625 (n12572, n_8009, n_8382);
  not g20626 (n_8383, n12569);
  not g20627 (n_8384, n12572);
  and g20628 (n12573, n_8383, n_8384);
  and g20629 (n12574, n_4218, n_8379);
  and g20630 (n12575, n_8380, n12574);
  not g20631 (n_8385, n12573);
  not g20632 (n_8386, n12575);
  and g20633 (n12576, n_8385, n_8386);
  not g20634 (n_8387, n12566);
  not g20635 (n_8388, n12576);
  and g20636 (n12577, n_8387, n_8388);
  not g20637 (n_8389, n12577);
  and g20638 (n12578, \asqrt[35] , n_8389);
  and g20642 (n12582, n_8019, n_8018);
  and g20643 (n12583, \asqrt[19] , n12582);
  not g20644 (n_8390, n12583);
  and g20645 (n12584, n_8017, n_8390);
  not g20646 (n_8391, n12581);
  not g20647 (n_8392, n12584);
  and g20648 (n12585, n_8391, n_8392);
  and g20649 (n12586, n_3962, n_8387);
  and g20650 (n12587, n_8388, n12586);
  not g20651 (n_8393, n12585);
  not g20652 (n_8394, n12587);
  and g20653 (n12588, n_8393, n_8394);
  not g20654 (n_8395, n12578);
  not g20655 (n_8396, n12588);
  and g20656 (n12589, n_8395, n_8396);
  not g20657 (n_8397, n12589);
  and g20658 (n12590, \asqrt[36] , n_8397);
  and g20662 (n12594, n_8027, n_8026);
  and g20663 (n12595, \asqrt[19] , n12594);
  not g20664 (n_8398, n12595);
  and g20665 (n12596, n_8025, n_8398);
  not g20666 (n_8399, n12593);
  not g20667 (n_8400, n12596);
  and g20668 (n12597, n_8399, n_8400);
  and g20669 (n12598, n_3714, n_8395);
  and g20670 (n12599, n_8396, n12598);
  not g20671 (n_8401, n12597);
  not g20672 (n_8402, n12599);
  and g20673 (n12600, n_8401, n_8402);
  not g20674 (n_8403, n12590);
  not g20675 (n_8404, n12600);
  and g20676 (n12601, n_8403, n_8404);
  not g20677 (n_8405, n12601);
  and g20678 (n12602, \asqrt[37] , n_8405);
  and g20682 (n12606, n_8035, n_8034);
  and g20683 (n12607, \asqrt[19] , n12606);
  not g20684 (n_8406, n12607);
  and g20685 (n12608, n_8033, n_8406);
  not g20686 (n_8407, n12605);
  not g20687 (n_8408, n12608);
  and g20688 (n12609, n_8407, n_8408);
  and g20689 (n12610, n_3474, n_8403);
  and g20690 (n12611, n_8404, n12610);
  not g20691 (n_8409, n12609);
  not g20692 (n_8410, n12611);
  and g20693 (n12612, n_8409, n_8410);
  not g20694 (n_8411, n12602);
  not g20695 (n_8412, n12612);
  and g20696 (n12613, n_8411, n_8412);
  not g20697 (n_8413, n12613);
  and g20698 (n12614, \asqrt[38] , n_8413);
  and g20702 (n12618, n_8043, n_8042);
  and g20703 (n12619, \asqrt[19] , n12618);
  not g20704 (n_8414, n12619);
  and g20705 (n12620, n_8041, n_8414);
  not g20706 (n_8415, n12617);
  not g20707 (n_8416, n12620);
  and g20708 (n12621, n_8415, n_8416);
  and g20709 (n12622, n_3242, n_8411);
  and g20710 (n12623, n_8412, n12622);
  not g20711 (n_8417, n12621);
  not g20712 (n_8418, n12623);
  and g20713 (n12624, n_8417, n_8418);
  not g20714 (n_8419, n12614);
  not g20715 (n_8420, n12624);
  and g20716 (n12625, n_8419, n_8420);
  not g20717 (n_8421, n12625);
  and g20718 (n12626, \asqrt[39] , n_8421);
  and g20722 (n12630, n_8051, n_8050);
  and g20723 (n12631, \asqrt[19] , n12630);
  not g20724 (n_8422, n12631);
  and g20725 (n12632, n_8049, n_8422);
  not g20726 (n_8423, n12629);
  not g20727 (n_8424, n12632);
  and g20728 (n12633, n_8423, n_8424);
  and g20729 (n12634, n_3018, n_8419);
  and g20730 (n12635, n_8420, n12634);
  not g20731 (n_8425, n12633);
  not g20732 (n_8426, n12635);
  and g20733 (n12636, n_8425, n_8426);
  not g20734 (n_8427, n12626);
  not g20735 (n_8428, n12636);
  and g20736 (n12637, n_8427, n_8428);
  not g20737 (n_8429, n12637);
  and g20738 (n12638, \asqrt[40] , n_8429);
  and g20742 (n12642, n_8059, n_8058);
  and g20743 (n12643, \asqrt[19] , n12642);
  not g20744 (n_8430, n12643);
  and g20745 (n12644, n_8057, n_8430);
  not g20746 (n_8431, n12641);
  not g20747 (n_8432, n12644);
  and g20748 (n12645, n_8431, n_8432);
  and g20749 (n12646, n_2802, n_8427);
  and g20750 (n12647, n_8428, n12646);
  not g20751 (n_8433, n12645);
  not g20752 (n_8434, n12647);
  and g20753 (n12648, n_8433, n_8434);
  not g20754 (n_8435, n12638);
  not g20755 (n_8436, n12648);
  and g20756 (n12649, n_8435, n_8436);
  not g20757 (n_8437, n12649);
  and g20758 (n12650, \asqrt[41] , n_8437);
  and g20762 (n12654, n_8067, n_8066);
  and g20763 (n12655, \asqrt[19] , n12654);
  not g20764 (n_8438, n12655);
  and g20765 (n12656, n_8065, n_8438);
  not g20766 (n_8439, n12653);
  not g20767 (n_8440, n12656);
  and g20768 (n12657, n_8439, n_8440);
  and g20769 (n12658, n_2594, n_8435);
  and g20770 (n12659, n_8436, n12658);
  not g20771 (n_8441, n12657);
  not g20772 (n_8442, n12659);
  and g20773 (n12660, n_8441, n_8442);
  not g20774 (n_8443, n12650);
  not g20775 (n_8444, n12660);
  and g20776 (n12661, n_8443, n_8444);
  not g20777 (n_8445, n12661);
  and g20778 (n12662, \asqrt[42] , n_8445);
  and g20782 (n12666, n_8075, n_8074);
  and g20783 (n12667, \asqrt[19] , n12666);
  not g20784 (n_8446, n12667);
  and g20785 (n12668, n_8073, n_8446);
  not g20786 (n_8447, n12665);
  not g20787 (n_8448, n12668);
  and g20788 (n12669, n_8447, n_8448);
  and g20789 (n12670, n_2394, n_8443);
  and g20790 (n12671, n_8444, n12670);
  not g20791 (n_8449, n12669);
  not g20792 (n_8450, n12671);
  and g20793 (n12672, n_8449, n_8450);
  not g20794 (n_8451, n12662);
  not g20795 (n_8452, n12672);
  and g20796 (n12673, n_8451, n_8452);
  not g20797 (n_8453, n12673);
  and g20798 (n12674, \asqrt[43] , n_8453);
  and g20802 (n12678, n_8083, n_8082);
  and g20803 (n12679, \asqrt[19] , n12678);
  not g20804 (n_8454, n12679);
  and g20805 (n12680, n_8081, n_8454);
  not g20806 (n_8455, n12677);
  not g20807 (n_8456, n12680);
  and g20808 (n12681, n_8455, n_8456);
  and g20809 (n12682, n_2202, n_8451);
  and g20810 (n12683, n_8452, n12682);
  not g20811 (n_8457, n12681);
  not g20812 (n_8458, n12683);
  and g20813 (n12684, n_8457, n_8458);
  not g20814 (n_8459, n12674);
  not g20815 (n_8460, n12684);
  and g20816 (n12685, n_8459, n_8460);
  not g20817 (n_8461, n12685);
  and g20818 (n12686, \asqrt[44] , n_8461);
  and g20822 (n12690, n_8091, n_8090);
  and g20823 (n12691, \asqrt[19] , n12690);
  not g20824 (n_8462, n12691);
  and g20825 (n12692, n_8089, n_8462);
  not g20826 (n_8463, n12689);
  not g20827 (n_8464, n12692);
  and g20828 (n12693, n_8463, n_8464);
  and g20829 (n12694, n_2018, n_8459);
  and g20830 (n12695, n_8460, n12694);
  not g20831 (n_8465, n12693);
  not g20832 (n_8466, n12695);
  and g20833 (n12696, n_8465, n_8466);
  not g20834 (n_8467, n12686);
  not g20835 (n_8468, n12696);
  and g20836 (n12697, n_8467, n_8468);
  not g20837 (n_8469, n12697);
  and g20838 (n12698, \asqrt[45] , n_8469);
  and g20842 (n12702, n_8099, n_8098);
  and g20843 (n12703, \asqrt[19] , n12702);
  not g20844 (n_8470, n12703);
  and g20845 (n12704, n_8097, n_8470);
  not g20846 (n_8471, n12701);
  not g20847 (n_8472, n12704);
  and g20848 (n12705, n_8471, n_8472);
  and g20849 (n12706, n_1842, n_8467);
  and g20850 (n12707, n_8468, n12706);
  not g20851 (n_8473, n12705);
  not g20852 (n_8474, n12707);
  and g20853 (n12708, n_8473, n_8474);
  not g20854 (n_8475, n12698);
  not g20855 (n_8476, n12708);
  and g20856 (n12709, n_8475, n_8476);
  not g20857 (n_8477, n12709);
  and g20858 (n12710, \asqrt[46] , n_8477);
  and g20859 (n12711, n_1674, n_8475);
  and g20860 (n12712, n_8476, n12711);
  and g20864 (n12716, n_8107, n_8105);
  and g20865 (n12717, \asqrt[19] , n12716);
  not g20866 (n_8478, n12717);
  and g20867 (n12718, n_8106, n_8478);
  not g20868 (n_8479, n12715);
  not g20869 (n_8480, n12718);
  and g20870 (n12719, n_8479, n_8480);
  not g20871 (n_8481, n12712);
  not g20872 (n_8482, n12719);
  and g20873 (n12720, n_8481, n_8482);
  not g20874 (n_8483, n12710);
  not g20875 (n_8484, n12720);
  and g20876 (n12721, n_8483, n_8484);
  not g20877 (n_8485, n12721);
  and g20878 (n12722, \asqrt[47] , n_8485);
  and g20882 (n12726, n_8115, n_8114);
  and g20883 (n12727, \asqrt[19] , n12726);
  not g20884 (n_8486, n12727);
  and g20885 (n12728, n_8113, n_8486);
  not g20886 (n_8487, n12725);
  not g20887 (n_8488, n12728);
  and g20888 (n12729, n_8487, n_8488);
  and g20889 (n12730, n_1514, n_8483);
  and g20890 (n12731, n_8484, n12730);
  not g20891 (n_8489, n12729);
  not g20892 (n_8490, n12731);
  and g20893 (n12732, n_8489, n_8490);
  not g20894 (n_8491, n12722);
  not g20895 (n_8492, n12732);
  and g20896 (n12733, n_8491, n_8492);
  not g20897 (n_8493, n12733);
  and g20898 (n12734, \asqrt[48] , n_8493);
  and g20902 (n12738, n_8123, n_8122);
  and g20903 (n12739, \asqrt[19] , n12738);
  not g20904 (n_8494, n12739);
  and g20905 (n12740, n_8121, n_8494);
  not g20906 (n_8495, n12737);
  not g20907 (n_8496, n12740);
  and g20908 (n12741, n_8495, n_8496);
  and g20909 (n12742, n_1362, n_8491);
  and g20910 (n12743, n_8492, n12742);
  not g20911 (n_8497, n12741);
  not g20912 (n_8498, n12743);
  and g20913 (n12744, n_8497, n_8498);
  not g20914 (n_8499, n12734);
  not g20915 (n_8500, n12744);
  and g20916 (n12745, n_8499, n_8500);
  not g20917 (n_8501, n12745);
  and g20918 (n12746, \asqrt[49] , n_8501);
  and g20922 (n12750, n_8131, n_8130);
  and g20923 (n12751, \asqrt[19] , n12750);
  not g20924 (n_8502, n12751);
  and g20925 (n12752, n_8129, n_8502);
  not g20926 (n_8503, n12749);
  not g20927 (n_8504, n12752);
  and g20928 (n12753, n_8503, n_8504);
  and g20929 (n12754, n_1218, n_8499);
  and g20930 (n12755, n_8500, n12754);
  not g20931 (n_8505, n12753);
  not g20932 (n_8506, n12755);
  and g20933 (n12756, n_8505, n_8506);
  not g20934 (n_8507, n12746);
  not g20935 (n_8508, n12756);
  and g20936 (n12757, n_8507, n_8508);
  not g20937 (n_8509, n12757);
  and g20938 (n12758, \asqrt[50] , n_8509);
  and g20942 (n12762, n_8139, n_8138);
  and g20943 (n12763, \asqrt[19] , n12762);
  not g20944 (n_8510, n12763);
  and g20945 (n12764, n_8137, n_8510);
  not g20946 (n_8511, n12761);
  not g20947 (n_8512, n12764);
  and g20948 (n12765, n_8511, n_8512);
  and g20949 (n12766, n_1082, n_8507);
  and g20950 (n12767, n_8508, n12766);
  not g20951 (n_8513, n12765);
  not g20952 (n_8514, n12767);
  and g20953 (n12768, n_8513, n_8514);
  not g20954 (n_8515, n12758);
  not g20955 (n_8516, n12768);
  and g20956 (n12769, n_8515, n_8516);
  not g20957 (n_8517, n12769);
  and g20958 (n12770, \asqrt[51] , n_8517);
  and g20962 (n12774, n_8147, n_8146);
  and g20963 (n12775, \asqrt[19] , n12774);
  not g20964 (n_8518, n12775);
  and g20965 (n12776, n_8145, n_8518);
  not g20966 (n_8519, n12773);
  not g20967 (n_8520, n12776);
  and g20968 (n12777, n_8519, n_8520);
  and g20969 (n12778, n_954, n_8515);
  and g20970 (n12779, n_8516, n12778);
  not g20971 (n_8521, n12777);
  not g20972 (n_8522, n12779);
  and g20973 (n12780, n_8521, n_8522);
  not g20974 (n_8523, n12770);
  not g20975 (n_8524, n12780);
  and g20976 (n12781, n_8523, n_8524);
  not g20977 (n_8525, n12781);
  and g20978 (n12782, \asqrt[52] , n_8525);
  and g20982 (n12786, n_8155, n_8154);
  and g20983 (n12787, \asqrt[19] , n12786);
  not g20984 (n_8526, n12787);
  and g20985 (n12788, n_8153, n_8526);
  not g20986 (n_8527, n12785);
  not g20987 (n_8528, n12788);
  and g20988 (n12789, n_8527, n_8528);
  and g20989 (n12790, n_834, n_8523);
  and g20990 (n12791, n_8524, n12790);
  not g20991 (n_8529, n12789);
  not g20992 (n_8530, n12791);
  and g20993 (n12792, n_8529, n_8530);
  not g20994 (n_8531, n12782);
  not g20995 (n_8532, n12792);
  and g20996 (n12793, n_8531, n_8532);
  not g20997 (n_8533, n12793);
  and g20998 (n12794, \asqrt[53] , n_8533);
  and g21002 (n12798, n_8163, n_8162);
  and g21003 (n12799, \asqrt[19] , n12798);
  not g21004 (n_8534, n12799);
  and g21005 (n12800, n_8161, n_8534);
  not g21006 (n_8535, n12797);
  not g21007 (n_8536, n12800);
  and g21008 (n12801, n_8535, n_8536);
  and g21009 (n12802, n_722, n_8531);
  and g21010 (n12803, n_8532, n12802);
  not g21011 (n_8537, n12801);
  not g21012 (n_8538, n12803);
  and g21013 (n12804, n_8537, n_8538);
  not g21014 (n_8539, n12794);
  not g21015 (n_8540, n12804);
  and g21016 (n12805, n_8539, n_8540);
  not g21017 (n_8541, n12805);
  and g21018 (n12806, \asqrt[54] , n_8541);
  and g21022 (n12810, n_8171, n_8170);
  and g21023 (n12811, \asqrt[19] , n12810);
  not g21024 (n_8542, n12811);
  and g21025 (n12812, n_8169, n_8542);
  not g21026 (n_8543, n12809);
  not g21027 (n_8544, n12812);
  and g21028 (n12813, n_8543, n_8544);
  and g21029 (n12814, n_618, n_8539);
  and g21030 (n12815, n_8540, n12814);
  not g21031 (n_8545, n12813);
  not g21032 (n_8546, n12815);
  and g21033 (n12816, n_8545, n_8546);
  not g21034 (n_8547, n12806);
  not g21035 (n_8548, n12816);
  and g21036 (n12817, n_8547, n_8548);
  not g21037 (n_8549, n12817);
  and g21038 (n12818, \asqrt[55] , n_8549);
  and g21042 (n12822, n_8179, n_8178);
  and g21043 (n12823, \asqrt[19] , n12822);
  not g21044 (n_8550, n12823);
  and g21045 (n12824, n_8177, n_8550);
  not g21046 (n_8551, n12821);
  not g21047 (n_8552, n12824);
  and g21048 (n12825, n_8551, n_8552);
  and g21049 (n12826, n_522, n_8547);
  and g21050 (n12827, n_8548, n12826);
  not g21051 (n_8553, n12825);
  not g21052 (n_8554, n12827);
  and g21053 (n12828, n_8553, n_8554);
  not g21054 (n_8555, n12818);
  not g21055 (n_8556, n12828);
  and g21056 (n12829, n_8555, n_8556);
  not g21057 (n_8557, n12829);
  and g21058 (n12830, \asqrt[56] , n_8557);
  and g21062 (n12834, n_8187, n_8186);
  and g21063 (n12835, \asqrt[19] , n12834);
  not g21064 (n_8558, n12835);
  and g21065 (n12836, n_8185, n_8558);
  not g21066 (n_8559, n12833);
  not g21067 (n_8560, n12836);
  and g21068 (n12837, n_8559, n_8560);
  and g21069 (n12838, n_434, n_8555);
  and g21070 (n12839, n_8556, n12838);
  not g21071 (n_8561, n12837);
  not g21072 (n_8562, n12839);
  and g21073 (n12840, n_8561, n_8562);
  not g21074 (n_8563, n12830);
  not g21075 (n_8564, n12840);
  and g21076 (n12841, n_8563, n_8564);
  not g21077 (n_8565, n12841);
  and g21078 (n12842, \asqrt[57] , n_8565);
  and g21082 (n12846, n_8195, n_8194);
  and g21083 (n12847, \asqrt[19] , n12846);
  not g21084 (n_8566, n12847);
  and g21085 (n12848, n_8193, n_8566);
  not g21086 (n_8567, n12845);
  not g21087 (n_8568, n12848);
  and g21088 (n12849, n_8567, n_8568);
  and g21089 (n12850, n_354, n_8563);
  and g21090 (n12851, n_8564, n12850);
  not g21091 (n_8569, n12849);
  not g21092 (n_8570, n12851);
  and g21093 (n12852, n_8569, n_8570);
  not g21094 (n_8571, n12842);
  not g21095 (n_8572, n12852);
  and g21096 (n12853, n_8571, n_8572);
  not g21097 (n_8573, n12853);
  and g21098 (n12854, \asqrt[58] , n_8573);
  and g21102 (n12858, n_8203, n_8202);
  and g21103 (n12859, \asqrt[19] , n12858);
  not g21104 (n_8574, n12859);
  and g21105 (n12860, n_8201, n_8574);
  not g21106 (n_8575, n12857);
  not g21107 (n_8576, n12860);
  and g21108 (n12861, n_8575, n_8576);
  and g21109 (n12862, n_282, n_8571);
  and g21110 (n12863, n_8572, n12862);
  not g21111 (n_8577, n12861);
  not g21112 (n_8578, n12863);
  and g21113 (n12864, n_8577, n_8578);
  not g21114 (n_8579, n12854);
  not g21115 (n_8580, n12864);
  and g21116 (n12865, n_8579, n_8580);
  not g21117 (n_8581, n12865);
  and g21118 (n12866, \asqrt[59] , n_8581);
  and g21122 (n12870, n_8211, n_8210);
  and g21123 (n12871, \asqrt[19] , n12870);
  not g21124 (n_8582, n12871);
  and g21125 (n12872, n_8209, n_8582);
  not g21126 (n_8583, n12869);
  not g21127 (n_8584, n12872);
  and g21128 (n12873, n_8583, n_8584);
  and g21129 (n12874, n_218, n_8579);
  and g21130 (n12875, n_8580, n12874);
  not g21131 (n_8585, n12873);
  not g21132 (n_8586, n12875);
  and g21133 (n12876, n_8585, n_8586);
  not g21134 (n_8587, n12866);
  not g21135 (n_8588, n12876);
  and g21136 (n12877, n_8587, n_8588);
  not g21137 (n_8589, n12877);
  and g21138 (n12878, \asqrt[60] , n_8589);
  and g21142 (n12882, n_8219, n_8218);
  and g21143 (n12883, \asqrt[19] , n12882);
  not g21144 (n_8590, n12883);
  and g21145 (n12884, n_8217, n_8590);
  not g21146 (n_8591, n12881);
  not g21147 (n_8592, n12884);
  and g21148 (n12885, n_8591, n_8592);
  and g21149 (n12886, n_162, n_8587);
  and g21150 (n12887, n_8588, n12886);
  not g21151 (n_8593, n12885);
  not g21152 (n_8594, n12887);
  and g21153 (n12888, n_8593, n_8594);
  not g21154 (n_8595, n12878);
  not g21155 (n_8596, n12888);
  and g21156 (n12889, n_8595, n_8596);
  not g21157 (n_8597, n12889);
  and g21158 (n12890, \asqrt[61] , n_8597);
  and g21162 (n12894, n_8227, n_8226);
  and g21163 (n12895, \asqrt[19] , n12894);
  not g21164 (n_8598, n12895);
  and g21165 (n12896, n_8225, n_8598);
  not g21166 (n_8599, n12893);
  not g21167 (n_8600, n12896);
  and g21168 (n12897, n_8599, n_8600);
  and g21169 (n12898, n_115, n_8595);
  and g21170 (n12899, n_8596, n12898);
  not g21171 (n_8601, n12897);
  not g21172 (n_8602, n12899);
  and g21173 (n12900, n_8601, n_8602);
  not g21174 (n_8603, n12890);
  not g21175 (n_8604, n12900);
  and g21176 (n12901, n_8603, n_8604);
  not g21177 (n_8605, n12901);
  and g21178 (n12902, \asqrt[62] , n_8605);
  and g21182 (n12906, n_8235, n_8234);
  and g21183 (n12907, \asqrt[19] , n12906);
  not g21184 (n_8606, n12907);
  and g21185 (n12908, n_8233, n_8606);
  not g21186 (n_8607, n12905);
  not g21187 (n_8608, n12908);
  and g21188 (n12909, n_8607, n_8608);
  and g21189 (n12910, n_76, n_8603);
  and g21190 (n12911, n_8604, n12910);
  not g21191 (n_8609, n12909);
  not g21192 (n_8610, n12911);
  and g21193 (n12912, n_8609, n_8610);
  not g21194 (n_8611, n12902);
  not g21195 (n_8612, n12912);
  and g21196 (n12913, n_8611, n_8612);
  and g21200 (n12917, n_8243, n_8242);
  and g21201 (n12918, \asqrt[19] , n12917);
  not g21202 (n_8613, n12918);
  and g21203 (n12919, n_8241, n_8613);
  not g21204 (n_8614, n12916);
  not g21205 (n_8615, n12919);
  and g21206 (n12920, n_8614, n_8615);
  and g21207 (n12921, n_8250, n_8249);
  and g21208 (n12922, \asqrt[19] , n12921);
  not g21211 (n_8617, n12920);
  not g21213 (n_8618, n12913);
  not g21215 (n_8619, n12925);
  and g21216 (n12926, n_21, n_8619);
  and g21217 (n12927, n_8611, n12920);
  and g21218 (n12928, n_8612, n12927);
  and g21219 (n12929, n_8249, \asqrt[19] );
  not g21220 (n_8620, n12929);
  and g21221 (n12930, n12365, n_8620);
  not g21222 (n_8621, n12921);
  and g21223 (n12931, \asqrt[63] , n_8621);
  not g21224 (n_8622, n12930);
  and g21225 (n12932, n_8622, n12931);
  not g21231 (n_8623, n12932);
  not g21232 (n_8624, n12937);
  not g21234 (n_8625, n12928);
  and g21238 (n12941, \a[36] , \asqrt[18] );
  not g21239 (n_8630, \a[34] );
  not g21240 (n_8631, \a[35] );
  and g21241 (n12942, n_8630, n_8631);
  and g21242 (n12943, n_8262, n12942);
  not g21243 (n_8632, n12941);
  not g21244 (n_8633, n12943);
  and g21245 (n12944, n_8632, n_8633);
  not g21246 (n_8634, n12944);
  and g21247 (n12945, \asqrt[19] , n_8634);
  and g21253 (n12951, n_8262, \asqrt[18] );
  not g21254 (n_8635, n12951);
  and g21255 (n12952, \a[37] , n_8635);
  and g21256 (n12953, n12394, \asqrt[18] );
  not g21257 (n_8636, n12952);
  not g21258 (n_8637, n12953);
  and g21259 (n12954, n_8636, n_8637);
  not g21260 (n_8638, n12950);
  and g21261 (n12955, n_8638, n12954);
  not g21262 (n_8639, n12945);
  not g21263 (n_8640, n12955);
  and g21264 (n12956, n_8639, n_8640);
  not g21265 (n_8641, n12956);
  and g21266 (n12957, \asqrt[20] , n_8641);
  not g21267 (n_8642, \asqrt[20] );
  and g21268 (n12958, n_8642, n_8639);
  and g21269 (n12959, n_8640, n12958);
  not g21273 (n_8643, n12926);
  not g21275 (n_8644, n12963);
  and g21276 (n12964, n_8637, n_8644);
  not g21277 (n_8645, n12964);
  and g21278 (n12965, \a[38] , n_8645);
  and g21279 (n12966, n_7902, n_8644);
  and g21280 (n12967, n_8637, n12966);
  not g21281 (n_8646, n12965);
  not g21282 (n_8647, n12967);
  and g21283 (n12968, n_8646, n_8647);
  not g21284 (n_8648, n12959);
  not g21285 (n_8649, n12968);
  and g21286 (n12969, n_8648, n_8649);
  not g21287 (n_8650, n12957);
  not g21288 (n_8651, n12969);
  and g21289 (n12970, n_8650, n_8651);
  not g21290 (n_8652, n12970);
  and g21291 (n12971, \asqrt[21] , n_8652);
  and g21292 (n12972, n_8271, n_8270);
  not g21293 (n_8653, n12406);
  and g21294 (n12973, n_8653, n12972);
  and g21295 (n12974, \asqrt[18] , n12973);
  and g21296 (n12975, \asqrt[18] , n12972);
  not g21297 (n_8654, n12975);
  and g21298 (n12976, n12406, n_8654);
  not g21299 (n_8655, n12974);
  not g21300 (n_8656, n12976);
  and g21301 (n12977, n_8655, n_8656);
  and g21302 (n12978, n_8274, n_8650);
  and g21303 (n12979, n_8651, n12978);
  not g21304 (n_8657, n12977);
  not g21305 (n_8658, n12979);
  and g21306 (n12980, n_8657, n_8658);
  not g21307 (n_8659, n12971);
  not g21308 (n_8660, n12980);
  and g21309 (n12981, n_8659, n_8660);
  not g21310 (n_8661, n12981);
  and g21311 (n12982, \asqrt[22] , n_8661);
  and g21315 (n12986, n_8282, n_8280);
  and g21316 (n12987, \asqrt[18] , n12986);
  not g21317 (n_8662, n12987);
  and g21318 (n12988, n_8281, n_8662);
  not g21319 (n_8663, n12985);
  not g21320 (n_8664, n12988);
  and g21321 (n12989, n_8663, n_8664);
  and g21322 (n12990, n_7914, n_8659);
  and g21323 (n12991, n_8660, n12990);
  not g21324 (n_8665, n12989);
  not g21325 (n_8666, n12991);
  and g21326 (n12992, n_8665, n_8666);
  not g21327 (n_8667, n12982);
  not g21328 (n_8668, n12992);
  and g21329 (n12993, n_8667, n_8668);
  not g21330 (n_8669, n12993);
  and g21331 (n12994, \asqrt[23] , n_8669);
  and g21335 (n12998, n_8291, n_8290);
  and g21336 (n12999, \asqrt[18] , n12998);
  not g21337 (n_8670, n12999);
  and g21338 (n13000, n_8289, n_8670);
  not g21339 (n_8671, n12997);
  not g21340 (n_8672, n13000);
  and g21341 (n13001, n_8671, n_8672);
  and g21342 (n13002, n_7562, n_8667);
  and g21343 (n13003, n_8668, n13002);
  not g21344 (n_8673, n13001);
  not g21345 (n_8674, n13003);
  and g21346 (n13004, n_8673, n_8674);
  not g21347 (n_8675, n12994);
  not g21348 (n_8676, n13004);
  and g21349 (n13005, n_8675, n_8676);
  not g21350 (n_8677, n13005);
  and g21351 (n13006, \asqrt[24] , n_8677);
  and g21355 (n13010, n_8299, n_8298);
  and g21356 (n13011, \asqrt[18] , n13010);
  not g21357 (n_8678, n13011);
  and g21358 (n13012, n_8297, n_8678);
  not g21359 (n_8679, n13009);
  not g21360 (n_8680, n13012);
  and g21361 (n13013, n_8679, n_8680);
  and g21362 (n13014, n_7218, n_8675);
  and g21363 (n13015, n_8676, n13014);
  not g21364 (n_8681, n13013);
  not g21365 (n_8682, n13015);
  and g21366 (n13016, n_8681, n_8682);
  not g21367 (n_8683, n13006);
  not g21368 (n_8684, n13016);
  and g21369 (n13017, n_8683, n_8684);
  not g21370 (n_8685, n13017);
  and g21371 (n13018, \asqrt[25] , n_8685);
  and g21375 (n13022, n_8307, n_8306);
  and g21376 (n13023, \asqrt[18] , n13022);
  not g21377 (n_8686, n13023);
  and g21378 (n13024, n_8305, n_8686);
  not g21379 (n_8687, n13021);
  not g21380 (n_8688, n13024);
  and g21381 (n13025, n_8687, n_8688);
  and g21382 (n13026, n_6882, n_8683);
  and g21383 (n13027, n_8684, n13026);
  not g21384 (n_8689, n13025);
  not g21385 (n_8690, n13027);
  and g21386 (n13028, n_8689, n_8690);
  not g21387 (n_8691, n13018);
  not g21388 (n_8692, n13028);
  and g21389 (n13029, n_8691, n_8692);
  not g21390 (n_8693, n13029);
  and g21391 (n13030, \asqrt[26] , n_8693);
  and g21395 (n13034, n_8315, n_8314);
  and g21396 (n13035, \asqrt[18] , n13034);
  not g21397 (n_8694, n13035);
  and g21398 (n13036, n_8313, n_8694);
  not g21399 (n_8695, n13033);
  not g21400 (n_8696, n13036);
  and g21401 (n13037, n_8695, n_8696);
  and g21402 (n13038, n_6554, n_8691);
  and g21403 (n13039, n_8692, n13038);
  not g21404 (n_8697, n13037);
  not g21405 (n_8698, n13039);
  and g21406 (n13040, n_8697, n_8698);
  not g21407 (n_8699, n13030);
  not g21408 (n_8700, n13040);
  and g21409 (n13041, n_8699, n_8700);
  not g21410 (n_8701, n13041);
  and g21411 (n13042, \asqrt[27] , n_8701);
  and g21415 (n13046, n_8323, n_8322);
  and g21416 (n13047, \asqrt[18] , n13046);
  not g21417 (n_8702, n13047);
  and g21418 (n13048, n_8321, n_8702);
  not g21419 (n_8703, n13045);
  not g21420 (n_8704, n13048);
  and g21421 (n13049, n_8703, n_8704);
  and g21422 (n13050, n_6234, n_8699);
  and g21423 (n13051, n_8700, n13050);
  not g21424 (n_8705, n13049);
  not g21425 (n_8706, n13051);
  and g21426 (n13052, n_8705, n_8706);
  not g21427 (n_8707, n13042);
  not g21428 (n_8708, n13052);
  and g21429 (n13053, n_8707, n_8708);
  not g21430 (n_8709, n13053);
  and g21431 (n13054, \asqrt[28] , n_8709);
  and g21435 (n13058, n_8331, n_8330);
  and g21436 (n13059, \asqrt[18] , n13058);
  not g21437 (n_8710, n13059);
  and g21438 (n13060, n_8329, n_8710);
  not g21439 (n_8711, n13057);
  not g21440 (n_8712, n13060);
  and g21441 (n13061, n_8711, n_8712);
  and g21442 (n13062, n_5922, n_8707);
  and g21443 (n13063, n_8708, n13062);
  not g21444 (n_8713, n13061);
  not g21445 (n_8714, n13063);
  and g21446 (n13064, n_8713, n_8714);
  not g21447 (n_8715, n13054);
  not g21448 (n_8716, n13064);
  and g21449 (n13065, n_8715, n_8716);
  not g21450 (n_8717, n13065);
  and g21451 (n13066, \asqrt[29] , n_8717);
  and g21455 (n13070, n_8339, n_8338);
  and g21456 (n13071, \asqrt[18] , n13070);
  not g21457 (n_8718, n13071);
  and g21458 (n13072, n_8337, n_8718);
  not g21459 (n_8719, n13069);
  not g21460 (n_8720, n13072);
  and g21461 (n13073, n_8719, n_8720);
  and g21462 (n13074, n_5618, n_8715);
  and g21463 (n13075, n_8716, n13074);
  not g21464 (n_8721, n13073);
  not g21465 (n_8722, n13075);
  and g21466 (n13076, n_8721, n_8722);
  not g21467 (n_8723, n13066);
  not g21468 (n_8724, n13076);
  and g21469 (n13077, n_8723, n_8724);
  not g21470 (n_8725, n13077);
  and g21471 (n13078, \asqrt[30] , n_8725);
  and g21475 (n13082, n_8347, n_8346);
  and g21476 (n13083, \asqrt[18] , n13082);
  not g21477 (n_8726, n13083);
  and g21478 (n13084, n_8345, n_8726);
  not g21479 (n_8727, n13081);
  not g21480 (n_8728, n13084);
  and g21481 (n13085, n_8727, n_8728);
  and g21482 (n13086, n_5322, n_8723);
  and g21483 (n13087, n_8724, n13086);
  not g21484 (n_8729, n13085);
  not g21485 (n_8730, n13087);
  and g21486 (n13088, n_8729, n_8730);
  not g21487 (n_8731, n13078);
  not g21488 (n_8732, n13088);
  and g21489 (n13089, n_8731, n_8732);
  not g21490 (n_8733, n13089);
  and g21491 (n13090, \asqrt[31] , n_8733);
  and g21495 (n13094, n_8355, n_8354);
  and g21496 (n13095, \asqrt[18] , n13094);
  not g21497 (n_8734, n13095);
  and g21498 (n13096, n_8353, n_8734);
  not g21499 (n_8735, n13093);
  not g21500 (n_8736, n13096);
  and g21501 (n13097, n_8735, n_8736);
  and g21502 (n13098, n_5034, n_8731);
  and g21503 (n13099, n_8732, n13098);
  not g21504 (n_8737, n13097);
  not g21505 (n_8738, n13099);
  and g21506 (n13100, n_8737, n_8738);
  not g21507 (n_8739, n13090);
  not g21508 (n_8740, n13100);
  and g21509 (n13101, n_8739, n_8740);
  not g21510 (n_8741, n13101);
  and g21511 (n13102, \asqrt[32] , n_8741);
  and g21515 (n13106, n_8363, n_8362);
  and g21516 (n13107, \asqrt[18] , n13106);
  not g21517 (n_8742, n13107);
  and g21518 (n13108, n_8361, n_8742);
  not g21519 (n_8743, n13105);
  not g21520 (n_8744, n13108);
  and g21521 (n13109, n_8743, n_8744);
  and g21522 (n13110, n_4754, n_8739);
  and g21523 (n13111, n_8740, n13110);
  not g21524 (n_8745, n13109);
  not g21525 (n_8746, n13111);
  and g21526 (n13112, n_8745, n_8746);
  not g21527 (n_8747, n13102);
  not g21528 (n_8748, n13112);
  and g21529 (n13113, n_8747, n_8748);
  not g21530 (n_8749, n13113);
  and g21531 (n13114, \asqrt[33] , n_8749);
  and g21535 (n13118, n_8371, n_8370);
  and g21536 (n13119, \asqrt[18] , n13118);
  not g21537 (n_8750, n13119);
  and g21538 (n13120, n_8369, n_8750);
  not g21539 (n_8751, n13117);
  not g21540 (n_8752, n13120);
  and g21541 (n13121, n_8751, n_8752);
  and g21542 (n13122, n_4482, n_8747);
  and g21543 (n13123, n_8748, n13122);
  not g21544 (n_8753, n13121);
  not g21545 (n_8754, n13123);
  and g21546 (n13124, n_8753, n_8754);
  not g21547 (n_8755, n13114);
  not g21548 (n_8756, n13124);
  and g21549 (n13125, n_8755, n_8756);
  not g21550 (n_8757, n13125);
  and g21551 (n13126, \asqrt[34] , n_8757);
  and g21555 (n13130, n_8379, n_8378);
  and g21556 (n13131, \asqrt[18] , n13130);
  not g21557 (n_8758, n13131);
  and g21558 (n13132, n_8377, n_8758);
  not g21559 (n_8759, n13129);
  not g21560 (n_8760, n13132);
  and g21561 (n13133, n_8759, n_8760);
  and g21562 (n13134, n_4218, n_8755);
  and g21563 (n13135, n_8756, n13134);
  not g21564 (n_8761, n13133);
  not g21565 (n_8762, n13135);
  and g21566 (n13136, n_8761, n_8762);
  not g21567 (n_8763, n13126);
  not g21568 (n_8764, n13136);
  and g21569 (n13137, n_8763, n_8764);
  not g21570 (n_8765, n13137);
  and g21571 (n13138, \asqrt[35] , n_8765);
  and g21575 (n13142, n_8387, n_8386);
  and g21576 (n13143, \asqrt[18] , n13142);
  not g21577 (n_8766, n13143);
  and g21578 (n13144, n_8385, n_8766);
  not g21579 (n_8767, n13141);
  not g21580 (n_8768, n13144);
  and g21581 (n13145, n_8767, n_8768);
  and g21582 (n13146, n_3962, n_8763);
  and g21583 (n13147, n_8764, n13146);
  not g21584 (n_8769, n13145);
  not g21585 (n_8770, n13147);
  and g21586 (n13148, n_8769, n_8770);
  not g21587 (n_8771, n13138);
  not g21588 (n_8772, n13148);
  and g21589 (n13149, n_8771, n_8772);
  not g21590 (n_8773, n13149);
  and g21591 (n13150, \asqrt[36] , n_8773);
  and g21595 (n13154, n_8395, n_8394);
  and g21596 (n13155, \asqrt[18] , n13154);
  not g21597 (n_8774, n13155);
  and g21598 (n13156, n_8393, n_8774);
  not g21599 (n_8775, n13153);
  not g21600 (n_8776, n13156);
  and g21601 (n13157, n_8775, n_8776);
  and g21602 (n13158, n_3714, n_8771);
  and g21603 (n13159, n_8772, n13158);
  not g21604 (n_8777, n13157);
  not g21605 (n_8778, n13159);
  and g21606 (n13160, n_8777, n_8778);
  not g21607 (n_8779, n13150);
  not g21608 (n_8780, n13160);
  and g21609 (n13161, n_8779, n_8780);
  not g21610 (n_8781, n13161);
  and g21611 (n13162, \asqrt[37] , n_8781);
  and g21615 (n13166, n_8403, n_8402);
  and g21616 (n13167, \asqrt[18] , n13166);
  not g21617 (n_8782, n13167);
  and g21618 (n13168, n_8401, n_8782);
  not g21619 (n_8783, n13165);
  not g21620 (n_8784, n13168);
  and g21621 (n13169, n_8783, n_8784);
  and g21622 (n13170, n_3474, n_8779);
  and g21623 (n13171, n_8780, n13170);
  not g21624 (n_8785, n13169);
  not g21625 (n_8786, n13171);
  and g21626 (n13172, n_8785, n_8786);
  not g21627 (n_8787, n13162);
  not g21628 (n_8788, n13172);
  and g21629 (n13173, n_8787, n_8788);
  not g21630 (n_8789, n13173);
  and g21631 (n13174, \asqrt[38] , n_8789);
  and g21635 (n13178, n_8411, n_8410);
  and g21636 (n13179, \asqrt[18] , n13178);
  not g21637 (n_8790, n13179);
  and g21638 (n13180, n_8409, n_8790);
  not g21639 (n_8791, n13177);
  not g21640 (n_8792, n13180);
  and g21641 (n13181, n_8791, n_8792);
  and g21642 (n13182, n_3242, n_8787);
  and g21643 (n13183, n_8788, n13182);
  not g21644 (n_8793, n13181);
  not g21645 (n_8794, n13183);
  and g21646 (n13184, n_8793, n_8794);
  not g21647 (n_8795, n13174);
  not g21648 (n_8796, n13184);
  and g21649 (n13185, n_8795, n_8796);
  not g21650 (n_8797, n13185);
  and g21651 (n13186, \asqrt[39] , n_8797);
  and g21655 (n13190, n_8419, n_8418);
  and g21656 (n13191, \asqrt[18] , n13190);
  not g21657 (n_8798, n13191);
  and g21658 (n13192, n_8417, n_8798);
  not g21659 (n_8799, n13189);
  not g21660 (n_8800, n13192);
  and g21661 (n13193, n_8799, n_8800);
  and g21662 (n13194, n_3018, n_8795);
  and g21663 (n13195, n_8796, n13194);
  not g21664 (n_8801, n13193);
  not g21665 (n_8802, n13195);
  and g21666 (n13196, n_8801, n_8802);
  not g21667 (n_8803, n13186);
  not g21668 (n_8804, n13196);
  and g21669 (n13197, n_8803, n_8804);
  not g21670 (n_8805, n13197);
  and g21671 (n13198, \asqrt[40] , n_8805);
  and g21675 (n13202, n_8427, n_8426);
  and g21676 (n13203, \asqrt[18] , n13202);
  not g21677 (n_8806, n13203);
  and g21678 (n13204, n_8425, n_8806);
  not g21679 (n_8807, n13201);
  not g21680 (n_8808, n13204);
  and g21681 (n13205, n_8807, n_8808);
  and g21682 (n13206, n_2802, n_8803);
  and g21683 (n13207, n_8804, n13206);
  not g21684 (n_8809, n13205);
  not g21685 (n_8810, n13207);
  and g21686 (n13208, n_8809, n_8810);
  not g21687 (n_8811, n13198);
  not g21688 (n_8812, n13208);
  and g21689 (n13209, n_8811, n_8812);
  not g21690 (n_8813, n13209);
  and g21691 (n13210, \asqrt[41] , n_8813);
  and g21695 (n13214, n_8435, n_8434);
  and g21696 (n13215, \asqrt[18] , n13214);
  not g21697 (n_8814, n13215);
  and g21698 (n13216, n_8433, n_8814);
  not g21699 (n_8815, n13213);
  not g21700 (n_8816, n13216);
  and g21701 (n13217, n_8815, n_8816);
  and g21702 (n13218, n_2594, n_8811);
  and g21703 (n13219, n_8812, n13218);
  not g21704 (n_8817, n13217);
  not g21705 (n_8818, n13219);
  and g21706 (n13220, n_8817, n_8818);
  not g21707 (n_8819, n13210);
  not g21708 (n_8820, n13220);
  and g21709 (n13221, n_8819, n_8820);
  not g21710 (n_8821, n13221);
  and g21711 (n13222, \asqrt[42] , n_8821);
  and g21715 (n13226, n_8443, n_8442);
  and g21716 (n13227, \asqrt[18] , n13226);
  not g21717 (n_8822, n13227);
  and g21718 (n13228, n_8441, n_8822);
  not g21719 (n_8823, n13225);
  not g21720 (n_8824, n13228);
  and g21721 (n13229, n_8823, n_8824);
  and g21722 (n13230, n_2394, n_8819);
  and g21723 (n13231, n_8820, n13230);
  not g21724 (n_8825, n13229);
  not g21725 (n_8826, n13231);
  and g21726 (n13232, n_8825, n_8826);
  not g21727 (n_8827, n13222);
  not g21728 (n_8828, n13232);
  and g21729 (n13233, n_8827, n_8828);
  not g21730 (n_8829, n13233);
  and g21731 (n13234, \asqrt[43] , n_8829);
  and g21735 (n13238, n_8451, n_8450);
  and g21736 (n13239, \asqrt[18] , n13238);
  not g21737 (n_8830, n13239);
  and g21738 (n13240, n_8449, n_8830);
  not g21739 (n_8831, n13237);
  not g21740 (n_8832, n13240);
  and g21741 (n13241, n_8831, n_8832);
  and g21742 (n13242, n_2202, n_8827);
  and g21743 (n13243, n_8828, n13242);
  not g21744 (n_8833, n13241);
  not g21745 (n_8834, n13243);
  and g21746 (n13244, n_8833, n_8834);
  not g21747 (n_8835, n13234);
  not g21748 (n_8836, n13244);
  and g21749 (n13245, n_8835, n_8836);
  not g21750 (n_8837, n13245);
  and g21751 (n13246, \asqrt[44] , n_8837);
  and g21755 (n13250, n_8459, n_8458);
  and g21756 (n13251, \asqrt[18] , n13250);
  not g21757 (n_8838, n13251);
  and g21758 (n13252, n_8457, n_8838);
  not g21759 (n_8839, n13249);
  not g21760 (n_8840, n13252);
  and g21761 (n13253, n_8839, n_8840);
  and g21762 (n13254, n_2018, n_8835);
  and g21763 (n13255, n_8836, n13254);
  not g21764 (n_8841, n13253);
  not g21765 (n_8842, n13255);
  and g21766 (n13256, n_8841, n_8842);
  not g21767 (n_8843, n13246);
  not g21768 (n_8844, n13256);
  and g21769 (n13257, n_8843, n_8844);
  not g21770 (n_8845, n13257);
  and g21771 (n13258, \asqrt[45] , n_8845);
  and g21775 (n13262, n_8467, n_8466);
  and g21776 (n13263, \asqrt[18] , n13262);
  not g21777 (n_8846, n13263);
  and g21778 (n13264, n_8465, n_8846);
  not g21779 (n_8847, n13261);
  not g21780 (n_8848, n13264);
  and g21781 (n13265, n_8847, n_8848);
  and g21782 (n13266, n_1842, n_8843);
  and g21783 (n13267, n_8844, n13266);
  not g21784 (n_8849, n13265);
  not g21785 (n_8850, n13267);
  and g21786 (n13268, n_8849, n_8850);
  not g21787 (n_8851, n13258);
  not g21788 (n_8852, n13268);
  and g21789 (n13269, n_8851, n_8852);
  not g21790 (n_8853, n13269);
  and g21791 (n13270, \asqrt[46] , n_8853);
  and g21795 (n13274, n_8475, n_8474);
  and g21796 (n13275, \asqrt[18] , n13274);
  not g21797 (n_8854, n13275);
  and g21798 (n13276, n_8473, n_8854);
  not g21799 (n_8855, n13273);
  not g21800 (n_8856, n13276);
  and g21801 (n13277, n_8855, n_8856);
  and g21802 (n13278, n_1674, n_8851);
  and g21803 (n13279, n_8852, n13278);
  not g21804 (n_8857, n13277);
  not g21805 (n_8858, n13279);
  and g21806 (n13280, n_8857, n_8858);
  not g21807 (n_8859, n13270);
  not g21808 (n_8860, n13280);
  and g21809 (n13281, n_8859, n_8860);
  not g21810 (n_8861, n13281);
  and g21811 (n13282, \asqrt[47] , n_8861);
  and g21812 (n13283, n_1514, n_8859);
  and g21813 (n13284, n_8860, n13283);
  and g21817 (n13288, n_8483, n_8481);
  and g21818 (n13289, \asqrt[18] , n13288);
  not g21819 (n_8862, n13289);
  and g21820 (n13290, n_8482, n_8862);
  not g21821 (n_8863, n13287);
  not g21822 (n_8864, n13290);
  and g21823 (n13291, n_8863, n_8864);
  not g21824 (n_8865, n13284);
  not g21825 (n_8866, n13291);
  and g21826 (n13292, n_8865, n_8866);
  not g21827 (n_8867, n13282);
  not g21828 (n_8868, n13292);
  and g21829 (n13293, n_8867, n_8868);
  not g21830 (n_8869, n13293);
  and g21831 (n13294, \asqrt[48] , n_8869);
  and g21835 (n13298, n_8491, n_8490);
  and g21836 (n13299, \asqrt[18] , n13298);
  not g21837 (n_8870, n13299);
  and g21838 (n13300, n_8489, n_8870);
  not g21839 (n_8871, n13297);
  not g21840 (n_8872, n13300);
  and g21841 (n13301, n_8871, n_8872);
  and g21842 (n13302, n_1362, n_8867);
  and g21843 (n13303, n_8868, n13302);
  not g21844 (n_8873, n13301);
  not g21845 (n_8874, n13303);
  and g21846 (n13304, n_8873, n_8874);
  not g21847 (n_8875, n13294);
  not g21848 (n_8876, n13304);
  and g21849 (n13305, n_8875, n_8876);
  not g21850 (n_8877, n13305);
  and g21851 (n13306, \asqrt[49] , n_8877);
  and g21855 (n13310, n_8499, n_8498);
  and g21856 (n13311, \asqrt[18] , n13310);
  not g21857 (n_8878, n13311);
  and g21858 (n13312, n_8497, n_8878);
  not g21859 (n_8879, n13309);
  not g21860 (n_8880, n13312);
  and g21861 (n13313, n_8879, n_8880);
  and g21862 (n13314, n_1218, n_8875);
  and g21863 (n13315, n_8876, n13314);
  not g21864 (n_8881, n13313);
  not g21865 (n_8882, n13315);
  and g21866 (n13316, n_8881, n_8882);
  not g21867 (n_8883, n13306);
  not g21868 (n_8884, n13316);
  and g21869 (n13317, n_8883, n_8884);
  not g21870 (n_8885, n13317);
  and g21871 (n13318, \asqrt[50] , n_8885);
  and g21875 (n13322, n_8507, n_8506);
  and g21876 (n13323, \asqrt[18] , n13322);
  not g21877 (n_8886, n13323);
  and g21878 (n13324, n_8505, n_8886);
  not g21879 (n_8887, n13321);
  not g21880 (n_8888, n13324);
  and g21881 (n13325, n_8887, n_8888);
  and g21882 (n13326, n_1082, n_8883);
  and g21883 (n13327, n_8884, n13326);
  not g21884 (n_8889, n13325);
  not g21885 (n_8890, n13327);
  and g21886 (n13328, n_8889, n_8890);
  not g21887 (n_8891, n13318);
  not g21888 (n_8892, n13328);
  and g21889 (n13329, n_8891, n_8892);
  not g21890 (n_8893, n13329);
  and g21891 (n13330, \asqrt[51] , n_8893);
  and g21895 (n13334, n_8515, n_8514);
  and g21896 (n13335, \asqrt[18] , n13334);
  not g21897 (n_8894, n13335);
  and g21898 (n13336, n_8513, n_8894);
  not g21899 (n_8895, n13333);
  not g21900 (n_8896, n13336);
  and g21901 (n13337, n_8895, n_8896);
  and g21902 (n13338, n_954, n_8891);
  and g21903 (n13339, n_8892, n13338);
  not g21904 (n_8897, n13337);
  not g21905 (n_8898, n13339);
  and g21906 (n13340, n_8897, n_8898);
  not g21907 (n_8899, n13330);
  not g21908 (n_8900, n13340);
  and g21909 (n13341, n_8899, n_8900);
  not g21910 (n_8901, n13341);
  and g21911 (n13342, \asqrt[52] , n_8901);
  and g21915 (n13346, n_8523, n_8522);
  and g21916 (n13347, \asqrt[18] , n13346);
  not g21917 (n_8902, n13347);
  and g21918 (n13348, n_8521, n_8902);
  not g21919 (n_8903, n13345);
  not g21920 (n_8904, n13348);
  and g21921 (n13349, n_8903, n_8904);
  and g21922 (n13350, n_834, n_8899);
  and g21923 (n13351, n_8900, n13350);
  not g21924 (n_8905, n13349);
  not g21925 (n_8906, n13351);
  and g21926 (n13352, n_8905, n_8906);
  not g21927 (n_8907, n13342);
  not g21928 (n_8908, n13352);
  and g21929 (n13353, n_8907, n_8908);
  not g21930 (n_8909, n13353);
  and g21931 (n13354, \asqrt[53] , n_8909);
  and g21935 (n13358, n_8531, n_8530);
  and g21936 (n13359, \asqrt[18] , n13358);
  not g21937 (n_8910, n13359);
  and g21938 (n13360, n_8529, n_8910);
  not g21939 (n_8911, n13357);
  not g21940 (n_8912, n13360);
  and g21941 (n13361, n_8911, n_8912);
  and g21942 (n13362, n_722, n_8907);
  and g21943 (n13363, n_8908, n13362);
  not g21944 (n_8913, n13361);
  not g21945 (n_8914, n13363);
  and g21946 (n13364, n_8913, n_8914);
  not g21947 (n_8915, n13354);
  not g21948 (n_8916, n13364);
  and g21949 (n13365, n_8915, n_8916);
  not g21950 (n_8917, n13365);
  and g21951 (n13366, \asqrt[54] , n_8917);
  and g21955 (n13370, n_8539, n_8538);
  and g21956 (n13371, \asqrt[18] , n13370);
  not g21957 (n_8918, n13371);
  and g21958 (n13372, n_8537, n_8918);
  not g21959 (n_8919, n13369);
  not g21960 (n_8920, n13372);
  and g21961 (n13373, n_8919, n_8920);
  and g21962 (n13374, n_618, n_8915);
  and g21963 (n13375, n_8916, n13374);
  not g21964 (n_8921, n13373);
  not g21965 (n_8922, n13375);
  and g21966 (n13376, n_8921, n_8922);
  not g21967 (n_8923, n13366);
  not g21968 (n_8924, n13376);
  and g21969 (n13377, n_8923, n_8924);
  not g21970 (n_8925, n13377);
  and g21971 (n13378, \asqrt[55] , n_8925);
  and g21975 (n13382, n_8547, n_8546);
  and g21976 (n13383, \asqrt[18] , n13382);
  not g21977 (n_8926, n13383);
  and g21978 (n13384, n_8545, n_8926);
  not g21979 (n_8927, n13381);
  not g21980 (n_8928, n13384);
  and g21981 (n13385, n_8927, n_8928);
  and g21982 (n13386, n_522, n_8923);
  and g21983 (n13387, n_8924, n13386);
  not g21984 (n_8929, n13385);
  not g21985 (n_8930, n13387);
  and g21986 (n13388, n_8929, n_8930);
  not g21987 (n_8931, n13378);
  not g21988 (n_8932, n13388);
  and g21989 (n13389, n_8931, n_8932);
  not g21990 (n_8933, n13389);
  and g21991 (n13390, \asqrt[56] , n_8933);
  and g21995 (n13394, n_8555, n_8554);
  and g21996 (n13395, \asqrt[18] , n13394);
  not g21997 (n_8934, n13395);
  and g21998 (n13396, n_8553, n_8934);
  not g21999 (n_8935, n13393);
  not g22000 (n_8936, n13396);
  and g22001 (n13397, n_8935, n_8936);
  and g22002 (n13398, n_434, n_8931);
  and g22003 (n13399, n_8932, n13398);
  not g22004 (n_8937, n13397);
  not g22005 (n_8938, n13399);
  and g22006 (n13400, n_8937, n_8938);
  not g22007 (n_8939, n13390);
  not g22008 (n_8940, n13400);
  and g22009 (n13401, n_8939, n_8940);
  not g22010 (n_8941, n13401);
  and g22011 (n13402, \asqrt[57] , n_8941);
  and g22015 (n13406, n_8563, n_8562);
  and g22016 (n13407, \asqrt[18] , n13406);
  not g22017 (n_8942, n13407);
  and g22018 (n13408, n_8561, n_8942);
  not g22019 (n_8943, n13405);
  not g22020 (n_8944, n13408);
  and g22021 (n13409, n_8943, n_8944);
  and g22022 (n13410, n_354, n_8939);
  and g22023 (n13411, n_8940, n13410);
  not g22024 (n_8945, n13409);
  not g22025 (n_8946, n13411);
  and g22026 (n13412, n_8945, n_8946);
  not g22027 (n_8947, n13402);
  not g22028 (n_8948, n13412);
  and g22029 (n13413, n_8947, n_8948);
  not g22030 (n_8949, n13413);
  and g22031 (n13414, \asqrt[58] , n_8949);
  and g22035 (n13418, n_8571, n_8570);
  and g22036 (n13419, \asqrt[18] , n13418);
  not g22037 (n_8950, n13419);
  and g22038 (n13420, n_8569, n_8950);
  not g22039 (n_8951, n13417);
  not g22040 (n_8952, n13420);
  and g22041 (n13421, n_8951, n_8952);
  and g22042 (n13422, n_282, n_8947);
  and g22043 (n13423, n_8948, n13422);
  not g22044 (n_8953, n13421);
  not g22045 (n_8954, n13423);
  and g22046 (n13424, n_8953, n_8954);
  not g22047 (n_8955, n13414);
  not g22048 (n_8956, n13424);
  and g22049 (n13425, n_8955, n_8956);
  not g22050 (n_8957, n13425);
  and g22051 (n13426, \asqrt[59] , n_8957);
  and g22055 (n13430, n_8579, n_8578);
  and g22056 (n13431, \asqrt[18] , n13430);
  not g22057 (n_8958, n13431);
  and g22058 (n13432, n_8577, n_8958);
  not g22059 (n_8959, n13429);
  not g22060 (n_8960, n13432);
  and g22061 (n13433, n_8959, n_8960);
  and g22062 (n13434, n_218, n_8955);
  and g22063 (n13435, n_8956, n13434);
  not g22064 (n_8961, n13433);
  not g22065 (n_8962, n13435);
  and g22066 (n13436, n_8961, n_8962);
  not g22067 (n_8963, n13426);
  not g22068 (n_8964, n13436);
  and g22069 (n13437, n_8963, n_8964);
  not g22070 (n_8965, n13437);
  and g22071 (n13438, \asqrt[60] , n_8965);
  and g22075 (n13442, n_8587, n_8586);
  and g22076 (n13443, \asqrt[18] , n13442);
  not g22077 (n_8966, n13443);
  and g22078 (n13444, n_8585, n_8966);
  not g22079 (n_8967, n13441);
  not g22080 (n_8968, n13444);
  and g22081 (n13445, n_8967, n_8968);
  and g22082 (n13446, n_162, n_8963);
  and g22083 (n13447, n_8964, n13446);
  not g22084 (n_8969, n13445);
  not g22085 (n_8970, n13447);
  and g22086 (n13448, n_8969, n_8970);
  not g22087 (n_8971, n13438);
  not g22088 (n_8972, n13448);
  and g22089 (n13449, n_8971, n_8972);
  not g22090 (n_8973, n13449);
  and g22091 (n13450, \asqrt[61] , n_8973);
  and g22095 (n13454, n_8595, n_8594);
  and g22096 (n13455, \asqrt[18] , n13454);
  not g22097 (n_8974, n13455);
  and g22098 (n13456, n_8593, n_8974);
  not g22099 (n_8975, n13453);
  not g22100 (n_8976, n13456);
  and g22101 (n13457, n_8975, n_8976);
  and g22102 (n13458, n_115, n_8971);
  and g22103 (n13459, n_8972, n13458);
  not g22104 (n_8977, n13457);
  not g22105 (n_8978, n13459);
  and g22106 (n13460, n_8977, n_8978);
  not g22107 (n_8979, n13450);
  not g22108 (n_8980, n13460);
  and g22109 (n13461, n_8979, n_8980);
  not g22110 (n_8981, n13461);
  and g22111 (n13462, \asqrt[62] , n_8981);
  and g22115 (n13466, n_8603, n_8602);
  and g22116 (n13467, \asqrt[18] , n13466);
  not g22117 (n_8982, n13467);
  and g22118 (n13468, n_8601, n_8982);
  not g22119 (n_8983, n13465);
  not g22120 (n_8984, n13468);
  and g22121 (n13469, n_8983, n_8984);
  and g22122 (n13470, n_76, n_8979);
  and g22123 (n13471, n_8980, n13470);
  not g22124 (n_8985, n13469);
  not g22125 (n_8986, n13471);
  and g22126 (n13472, n_8985, n_8986);
  not g22127 (n_8987, n13462);
  not g22128 (n_8988, n13472);
  and g22129 (n13473, n_8987, n_8988);
  and g22133 (n13477, n_8611, n_8610);
  and g22134 (n13478, \asqrt[18] , n13477);
  not g22135 (n_8989, n13478);
  and g22136 (n13479, n_8609, n_8989);
  not g22137 (n_8990, n13476);
  not g22138 (n_8991, n13479);
  and g22139 (n13480, n_8990, n_8991);
  and g22140 (n13481, n_8618, n_8617);
  and g22141 (n13482, \asqrt[18] , n13481);
  not g22144 (n_8993, n13480);
  not g22146 (n_8994, n13473);
  not g22148 (n_8995, n13485);
  and g22149 (n13486, n_21, n_8995);
  and g22150 (n13487, n_8987, n13480);
  and g22151 (n13488, n_8988, n13487);
  and g22152 (n13489, n_8617, \asqrt[18] );
  not g22153 (n_8996, n13489);
  and g22154 (n13490, n12913, n_8996);
  not g22155 (n_8997, n13481);
  and g22156 (n13491, \asqrt[63] , n_8997);
  not g22157 (n_8998, n13490);
  and g22158 (n13492, n_8998, n13491);
  not g22164 (n_8999, n13492);
  not g22165 (n_9000, n13497);
  not g22167 (n_9001, n13488);
  and g22171 (n13501, \a[34] , \asqrt[17] );
  not g22172 (n_9006, \a[32] );
  not g22173 (n_9007, \a[33] );
  and g22174 (n13502, n_9006, n_9007);
  and g22175 (n13503, n_8630, n13502);
  not g22176 (n_9008, n13501);
  not g22177 (n_9009, n13503);
  and g22178 (n13504, n_9008, n_9009);
  not g22179 (n_9010, n13504);
  and g22180 (n13505, \asqrt[18] , n_9010);
  and g22186 (n13511, n_8630, \asqrt[17] );
  not g22187 (n_9011, n13511);
  and g22188 (n13512, \a[35] , n_9011);
  and g22189 (n13513, n12942, \asqrt[17] );
  not g22190 (n_9012, n13512);
  not g22191 (n_9013, n13513);
  and g22192 (n13514, n_9012, n_9013);
  not g22193 (n_9014, n13510);
  and g22194 (n13515, n_9014, n13514);
  not g22195 (n_9015, n13505);
  not g22196 (n_9016, n13515);
  and g22197 (n13516, n_9015, n_9016);
  not g22198 (n_9017, n13516);
  and g22199 (n13517, \asqrt[19] , n_9017);
  not g22200 (n_9018, \asqrt[19] );
  and g22201 (n13518, n_9018, n_9015);
  and g22202 (n13519, n_9016, n13518);
  not g22206 (n_9019, n13486);
  not g22208 (n_9020, n13523);
  and g22209 (n13524, n_9013, n_9020);
  not g22210 (n_9021, n13524);
  and g22211 (n13525, \a[36] , n_9021);
  and g22212 (n13526, n_8262, n_9020);
  and g22213 (n13527, n_9013, n13526);
  not g22214 (n_9022, n13525);
  not g22215 (n_9023, n13527);
  and g22216 (n13528, n_9022, n_9023);
  not g22217 (n_9024, n13519);
  not g22218 (n_9025, n13528);
  and g22219 (n13529, n_9024, n_9025);
  not g22220 (n_9026, n13517);
  not g22221 (n_9027, n13529);
  and g22222 (n13530, n_9026, n_9027);
  not g22223 (n_9028, n13530);
  and g22224 (n13531, \asqrt[20] , n_9028);
  and g22225 (n13532, n_8639, n_8638);
  not g22226 (n_9029, n12954);
  and g22227 (n13533, n_9029, n13532);
  and g22228 (n13534, \asqrt[17] , n13533);
  and g22229 (n13535, \asqrt[17] , n13532);
  not g22230 (n_9030, n13535);
  and g22231 (n13536, n12954, n_9030);
  not g22232 (n_9031, n13534);
  not g22233 (n_9032, n13536);
  and g22234 (n13537, n_9031, n_9032);
  and g22235 (n13538, n_8642, n_9026);
  and g22236 (n13539, n_9027, n13538);
  not g22237 (n_9033, n13537);
  not g22238 (n_9034, n13539);
  and g22239 (n13540, n_9033, n_9034);
  not g22240 (n_9035, n13531);
  not g22241 (n_9036, n13540);
  and g22242 (n13541, n_9035, n_9036);
  not g22243 (n_9037, n13541);
  and g22244 (n13542, \asqrt[21] , n_9037);
  and g22248 (n13546, n_8650, n_8648);
  and g22249 (n13547, \asqrt[17] , n13546);
  not g22250 (n_9038, n13547);
  and g22251 (n13548, n_8649, n_9038);
  not g22252 (n_9039, n13545);
  not g22253 (n_9040, n13548);
  and g22254 (n13549, n_9039, n_9040);
  and g22255 (n13550, n_8274, n_9035);
  and g22256 (n13551, n_9036, n13550);
  not g22257 (n_9041, n13549);
  not g22258 (n_9042, n13551);
  and g22259 (n13552, n_9041, n_9042);
  not g22260 (n_9043, n13542);
  not g22261 (n_9044, n13552);
  and g22262 (n13553, n_9043, n_9044);
  not g22263 (n_9045, n13553);
  and g22264 (n13554, \asqrt[22] , n_9045);
  and g22268 (n13558, n_8659, n_8658);
  and g22269 (n13559, \asqrt[17] , n13558);
  not g22270 (n_9046, n13559);
  and g22271 (n13560, n_8657, n_9046);
  not g22272 (n_9047, n13557);
  not g22273 (n_9048, n13560);
  and g22274 (n13561, n_9047, n_9048);
  and g22275 (n13562, n_7914, n_9043);
  and g22276 (n13563, n_9044, n13562);
  not g22277 (n_9049, n13561);
  not g22278 (n_9050, n13563);
  and g22279 (n13564, n_9049, n_9050);
  not g22280 (n_9051, n13554);
  not g22281 (n_9052, n13564);
  and g22282 (n13565, n_9051, n_9052);
  not g22283 (n_9053, n13565);
  and g22284 (n13566, \asqrt[23] , n_9053);
  and g22288 (n13570, n_8667, n_8666);
  and g22289 (n13571, \asqrt[17] , n13570);
  not g22290 (n_9054, n13571);
  and g22291 (n13572, n_8665, n_9054);
  not g22292 (n_9055, n13569);
  not g22293 (n_9056, n13572);
  and g22294 (n13573, n_9055, n_9056);
  and g22295 (n13574, n_7562, n_9051);
  and g22296 (n13575, n_9052, n13574);
  not g22297 (n_9057, n13573);
  not g22298 (n_9058, n13575);
  and g22299 (n13576, n_9057, n_9058);
  not g22300 (n_9059, n13566);
  not g22301 (n_9060, n13576);
  and g22302 (n13577, n_9059, n_9060);
  not g22303 (n_9061, n13577);
  and g22304 (n13578, \asqrt[24] , n_9061);
  and g22308 (n13582, n_8675, n_8674);
  and g22309 (n13583, \asqrt[17] , n13582);
  not g22310 (n_9062, n13583);
  and g22311 (n13584, n_8673, n_9062);
  not g22312 (n_9063, n13581);
  not g22313 (n_9064, n13584);
  and g22314 (n13585, n_9063, n_9064);
  and g22315 (n13586, n_7218, n_9059);
  and g22316 (n13587, n_9060, n13586);
  not g22317 (n_9065, n13585);
  not g22318 (n_9066, n13587);
  and g22319 (n13588, n_9065, n_9066);
  not g22320 (n_9067, n13578);
  not g22321 (n_9068, n13588);
  and g22322 (n13589, n_9067, n_9068);
  not g22323 (n_9069, n13589);
  and g22324 (n13590, \asqrt[25] , n_9069);
  and g22328 (n13594, n_8683, n_8682);
  and g22329 (n13595, \asqrt[17] , n13594);
  not g22330 (n_9070, n13595);
  and g22331 (n13596, n_8681, n_9070);
  not g22332 (n_9071, n13593);
  not g22333 (n_9072, n13596);
  and g22334 (n13597, n_9071, n_9072);
  and g22335 (n13598, n_6882, n_9067);
  and g22336 (n13599, n_9068, n13598);
  not g22337 (n_9073, n13597);
  not g22338 (n_9074, n13599);
  and g22339 (n13600, n_9073, n_9074);
  not g22340 (n_9075, n13590);
  not g22341 (n_9076, n13600);
  and g22342 (n13601, n_9075, n_9076);
  not g22343 (n_9077, n13601);
  and g22344 (n13602, \asqrt[26] , n_9077);
  and g22348 (n13606, n_8691, n_8690);
  and g22349 (n13607, \asqrt[17] , n13606);
  not g22350 (n_9078, n13607);
  and g22351 (n13608, n_8689, n_9078);
  not g22352 (n_9079, n13605);
  not g22353 (n_9080, n13608);
  and g22354 (n13609, n_9079, n_9080);
  and g22355 (n13610, n_6554, n_9075);
  and g22356 (n13611, n_9076, n13610);
  not g22357 (n_9081, n13609);
  not g22358 (n_9082, n13611);
  and g22359 (n13612, n_9081, n_9082);
  not g22360 (n_9083, n13602);
  not g22361 (n_9084, n13612);
  and g22362 (n13613, n_9083, n_9084);
  not g22363 (n_9085, n13613);
  and g22364 (n13614, \asqrt[27] , n_9085);
  and g22368 (n13618, n_8699, n_8698);
  and g22369 (n13619, \asqrt[17] , n13618);
  not g22370 (n_9086, n13619);
  and g22371 (n13620, n_8697, n_9086);
  not g22372 (n_9087, n13617);
  not g22373 (n_9088, n13620);
  and g22374 (n13621, n_9087, n_9088);
  and g22375 (n13622, n_6234, n_9083);
  and g22376 (n13623, n_9084, n13622);
  not g22377 (n_9089, n13621);
  not g22378 (n_9090, n13623);
  and g22379 (n13624, n_9089, n_9090);
  not g22380 (n_9091, n13614);
  not g22381 (n_9092, n13624);
  and g22382 (n13625, n_9091, n_9092);
  not g22383 (n_9093, n13625);
  and g22384 (n13626, \asqrt[28] , n_9093);
  and g22388 (n13630, n_8707, n_8706);
  and g22389 (n13631, \asqrt[17] , n13630);
  not g22390 (n_9094, n13631);
  and g22391 (n13632, n_8705, n_9094);
  not g22392 (n_9095, n13629);
  not g22393 (n_9096, n13632);
  and g22394 (n13633, n_9095, n_9096);
  and g22395 (n13634, n_5922, n_9091);
  and g22396 (n13635, n_9092, n13634);
  not g22397 (n_9097, n13633);
  not g22398 (n_9098, n13635);
  and g22399 (n13636, n_9097, n_9098);
  not g22400 (n_9099, n13626);
  not g22401 (n_9100, n13636);
  and g22402 (n13637, n_9099, n_9100);
  not g22403 (n_9101, n13637);
  and g22404 (n13638, \asqrt[29] , n_9101);
  and g22408 (n13642, n_8715, n_8714);
  and g22409 (n13643, \asqrt[17] , n13642);
  not g22410 (n_9102, n13643);
  and g22411 (n13644, n_8713, n_9102);
  not g22412 (n_9103, n13641);
  not g22413 (n_9104, n13644);
  and g22414 (n13645, n_9103, n_9104);
  and g22415 (n13646, n_5618, n_9099);
  and g22416 (n13647, n_9100, n13646);
  not g22417 (n_9105, n13645);
  not g22418 (n_9106, n13647);
  and g22419 (n13648, n_9105, n_9106);
  not g22420 (n_9107, n13638);
  not g22421 (n_9108, n13648);
  and g22422 (n13649, n_9107, n_9108);
  not g22423 (n_9109, n13649);
  and g22424 (n13650, \asqrt[30] , n_9109);
  and g22428 (n13654, n_8723, n_8722);
  and g22429 (n13655, \asqrt[17] , n13654);
  not g22430 (n_9110, n13655);
  and g22431 (n13656, n_8721, n_9110);
  not g22432 (n_9111, n13653);
  not g22433 (n_9112, n13656);
  and g22434 (n13657, n_9111, n_9112);
  and g22435 (n13658, n_5322, n_9107);
  and g22436 (n13659, n_9108, n13658);
  not g22437 (n_9113, n13657);
  not g22438 (n_9114, n13659);
  and g22439 (n13660, n_9113, n_9114);
  not g22440 (n_9115, n13650);
  not g22441 (n_9116, n13660);
  and g22442 (n13661, n_9115, n_9116);
  not g22443 (n_9117, n13661);
  and g22444 (n13662, \asqrt[31] , n_9117);
  and g22448 (n13666, n_8731, n_8730);
  and g22449 (n13667, \asqrt[17] , n13666);
  not g22450 (n_9118, n13667);
  and g22451 (n13668, n_8729, n_9118);
  not g22452 (n_9119, n13665);
  not g22453 (n_9120, n13668);
  and g22454 (n13669, n_9119, n_9120);
  and g22455 (n13670, n_5034, n_9115);
  and g22456 (n13671, n_9116, n13670);
  not g22457 (n_9121, n13669);
  not g22458 (n_9122, n13671);
  and g22459 (n13672, n_9121, n_9122);
  not g22460 (n_9123, n13662);
  not g22461 (n_9124, n13672);
  and g22462 (n13673, n_9123, n_9124);
  not g22463 (n_9125, n13673);
  and g22464 (n13674, \asqrt[32] , n_9125);
  and g22468 (n13678, n_8739, n_8738);
  and g22469 (n13679, \asqrt[17] , n13678);
  not g22470 (n_9126, n13679);
  and g22471 (n13680, n_8737, n_9126);
  not g22472 (n_9127, n13677);
  not g22473 (n_9128, n13680);
  and g22474 (n13681, n_9127, n_9128);
  and g22475 (n13682, n_4754, n_9123);
  and g22476 (n13683, n_9124, n13682);
  not g22477 (n_9129, n13681);
  not g22478 (n_9130, n13683);
  and g22479 (n13684, n_9129, n_9130);
  not g22480 (n_9131, n13674);
  not g22481 (n_9132, n13684);
  and g22482 (n13685, n_9131, n_9132);
  not g22483 (n_9133, n13685);
  and g22484 (n13686, \asqrt[33] , n_9133);
  and g22488 (n13690, n_8747, n_8746);
  and g22489 (n13691, \asqrt[17] , n13690);
  not g22490 (n_9134, n13691);
  and g22491 (n13692, n_8745, n_9134);
  not g22492 (n_9135, n13689);
  not g22493 (n_9136, n13692);
  and g22494 (n13693, n_9135, n_9136);
  and g22495 (n13694, n_4482, n_9131);
  and g22496 (n13695, n_9132, n13694);
  not g22497 (n_9137, n13693);
  not g22498 (n_9138, n13695);
  and g22499 (n13696, n_9137, n_9138);
  not g22500 (n_9139, n13686);
  not g22501 (n_9140, n13696);
  and g22502 (n13697, n_9139, n_9140);
  not g22503 (n_9141, n13697);
  and g22504 (n13698, \asqrt[34] , n_9141);
  and g22508 (n13702, n_8755, n_8754);
  and g22509 (n13703, \asqrt[17] , n13702);
  not g22510 (n_9142, n13703);
  and g22511 (n13704, n_8753, n_9142);
  not g22512 (n_9143, n13701);
  not g22513 (n_9144, n13704);
  and g22514 (n13705, n_9143, n_9144);
  and g22515 (n13706, n_4218, n_9139);
  and g22516 (n13707, n_9140, n13706);
  not g22517 (n_9145, n13705);
  not g22518 (n_9146, n13707);
  and g22519 (n13708, n_9145, n_9146);
  not g22520 (n_9147, n13698);
  not g22521 (n_9148, n13708);
  and g22522 (n13709, n_9147, n_9148);
  not g22523 (n_9149, n13709);
  and g22524 (n13710, \asqrt[35] , n_9149);
  and g22528 (n13714, n_8763, n_8762);
  and g22529 (n13715, \asqrt[17] , n13714);
  not g22530 (n_9150, n13715);
  and g22531 (n13716, n_8761, n_9150);
  not g22532 (n_9151, n13713);
  not g22533 (n_9152, n13716);
  and g22534 (n13717, n_9151, n_9152);
  and g22535 (n13718, n_3962, n_9147);
  and g22536 (n13719, n_9148, n13718);
  not g22537 (n_9153, n13717);
  not g22538 (n_9154, n13719);
  and g22539 (n13720, n_9153, n_9154);
  not g22540 (n_9155, n13710);
  not g22541 (n_9156, n13720);
  and g22542 (n13721, n_9155, n_9156);
  not g22543 (n_9157, n13721);
  and g22544 (n13722, \asqrt[36] , n_9157);
  and g22548 (n13726, n_8771, n_8770);
  and g22549 (n13727, \asqrt[17] , n13726);
  not g22550 (n_9158, n13727);
  and g22551 (n13728, n_8769, n_9158);
  not g22552 (n_9159, n13725);
  not g22553 (n_9160, n13728);
  and g22554 (n13729, n_9159, n_9160);
  and g22555 (n13730, n_3714, n_9155);
  and g22556 (n13731, n_9156, n13730);
  not g22557 (n_9161, n13729);
  not g22558 (n_9162, n13731);
  and g22559 (n13732, n_9161, n_9162);
  not g22560 (n_9163, n13722);
  not g22561 (n_9164, n13732);
  and g22562 (n13733, n_9163, n_9164);
  not g22563 (n_9165, n13733);
  and g22564 (n13734, \asqrt[37] , n_9165);
  and g22568 (n13738, n_8779, n_8778);
  and g22569 (n13739, \asqrt[17] , n13738);
  not g22570 (n_9166, n13739);
  and g22571 (n13740, n_8777, n_9166);
  not g22572 (n_9167, n13737);
  not g22573 (n_9168, n13740);
  and g22574 (n13741, n_9167, n_9168);
  and g22575 (n13742, n_3474, n_9163);
  and g22576 (n13743, n_9164, n13742);
  not g22577 (n_9169, n13741);
  not g22578 (n_9170, n13743);
  and g22579 (n13744, n_9169, n_9170);
  not g22580 (n_9171, n13734);
  not g22581 (n_9172, n13744);
  and g22582 (n13745, n_9171, n_9172);
  not g22583 (n_9173, n13745);
  and g22584 (n13746, \asqrt[38] , n_9173);
  and g22588 (n13750, n_8787, n_8786);
  and g22589 (n13751, \asqrt[17] , n13750);
  not g22590 (n_9174, n13751);
  and g22591 (n13752, n_8785, n_9174);
  not g22592 (n_9175, n13749);
  not g22593 (n_9176, n13752);
  and g22594 (n13753, n_9175, n_9176);
  and g22595 (n13754, n_3242, n_9171);
  and g22596 (n13755, n_9172, n13754);
  not g22597 (n_9177, n13753);
  not g22598 (n_9178, n13755);
  and g22599 (n13756, n_9177, n_9178);
  not g22600 (n_9179, n13746);
  not g22601 (n_9180, n13756);
  and g22602 (n13757, n_9179, n_9180);
  not g22603 (n_9181, n13757);
  and g22604 (n13758, \asqrt[39] , n_9181);
  and g22608 (n13762, n_8795, n_8794);
  and g22609 (n13763, \asqrt[17] , n13762);
  not g22610 (n_9182, n13763);
  and g22611 (n13764, n_8793, n_9182);
  not g22612 (n_9183, n13761);
  not g22613 (n_9184, n13764);
  and g22614 (n13765, n_9183, n_9184);
  and g22615 (n13766, n_3018, n_9179);
  and g22616 (n13767, n_9180, n13766);
  not g22617 (n_9185, n13765);
  not g22618 (n_9186, n13767);
  and g22619 (n13768, n_9185, n_9186);
  not g22620 (n_9187, n13758);
  not g22621 (n_9188, n13768);
  and g22622 (n13769, n_9187, n_9188);
  not g22623 (n_9189, n13769);
  and g22624 (n13770, \asqrt[40] , n_9189);
  and g22628 (n13774, n_8803, n_8802);
  and g22629 (n13775, \asqrt[17] , n13774);
  not g22630 (n_9190, n13775);
  and g22631 (n13776, n_8801, n_9190);
  not g22632 (n_9191, n13773);
  not g22633 (n_9192, n13776);
  and g22634 (n13777, n_9191, n_9192);
  and g22635 (n13778, n_2802, n_9187);
  and g22636 (n13779, n_9188, n13778);
  not g22637 (n_9193, n13777);
  not g22638 (n_9194, n13779);
  and g22639 (n13780, n_9193, n_9194);
  not g22640 (n_9195, n13770);
  not g22641 (n_9196, n13780);
  and g22642 (n13781, n_9195, n_9196);
  not g22643 (n_9197, n13781);
  and g22644 (n13782, \asqrt[41] , n_9197);
  and g22648 (n13786, n_8811, n_8810);
  and g22649 (n13787, \asqrt[17] , n13786);
  not g22650 (n_9198, n13787);
  and g22651 (n13788, n_8809, n_9198);
  not g22652 (n_9199, n13785);
  not g22653 (n_9200, n13788);
  and g22654 (n13789, n_9199, n_9200);
  and g22655 (n13790, n_2594, n_9195);
  and g22656 (n13791, n_9196, n13790);
  not g22657 (n_9201, n13789);
  not g22658 (n_9202, n13791);
  and g22659 (n13792, n_9201, n_9202);
  not g22660 (n_9203, n13782);
  not g22661 (n_9204, n13792);
  and g22662 (n13793, n_9203, n_9204);
  not g22663 (n_9205, n13793);
  and g22664 (n13794, \asqrt[42] , n_9205);
  and g22668 (n13798, n_8819, n_8818);
  and g22669 (n13799, \asqrt[17] , n13798);
  not g22670 (n_9206, n13799);
  and g22671 (n13800, n_8817, n_9206);
  not g22672 (n_9207, n13797);
  not g22673 (n_9208, n13800);
  and g22674 (n13801, n_9207, n_9208);
  and g22675 (n13802, n_2394, n_9203);
  and g22676 (n13803, n_9204, n13802);
  not g22677 (n_9209, n13801);
  not g22678 (n_9210, n13803);
  and g22679 (n13804, n_9209, n_9210);
  not g22680 (n_9211, n13794);
  not g22681 (n_9212, n13804);
  and g22682 (n13805, n_9211, n_9212);
  not g22683 (n_9213, n13805);
  and g22684 (n13806, \asqrt[43] , n_9213);
  and g22688 (n13810, n_8827, n_8826);
  and g22689 (n13811, \asqrt[17] , n13810);
  not g22690 (n_9214, n13811);
  and g22691 (n13812, n_8825, n_9214);
  not g22692 (n_9215, n13809);
  not g22693 (n_9216, n13812);
  and g22694 (n13813, n_9215, n_9216);
  and g22695 (n13814, n_2202, n_9211);
  and g22696 (n13815, n_9212, n13814);
  not g22697 (n_9217, n13813);
  not g22698 (n_9218, n13815);
  and g22699 (n13816, n_9217, n_9218);
  not g22700 (n_9219, n13806);
  not g22701 (n_9220, n13816);
  and g22702 (n13817, n_9219, n_9220);
  not g22703 (n_9221, n13817);
  and g22704 (n13818, \asqrt[44] , n_9221);
  and g22708 (n13822, n_8835, n_8834);
  and g22709 (n13823, \asqrt[17] , n13822);
  not g22710 (n_9222, n13823);
  and g22711 (n13824, n_8833, n_9222);
  not g22712 (n_9223, n13821);
  not g22713 (n_9224, n13824);
  and g22714 (n13825, n_9223, n_9224);
  and g22715 (n13826, n_2018, n_9219);
  and g22716 (n13827, n_9220, n13826);
  not g22717 (n_9225, n13825);
  not g22718 (n_9226, n13827);
  and g22719 (n13828, n_9225, n_9226);
  not g22720 (n_9227, n13818);
  not g22721 (n_9228, n13828);
  and g22722 (n13829, n_9227, n_9228);
  not g22723 (n_9229, n13829);
  and g22724 (n13830, \asqrt[45] , n_9229);
  and g22728 (n13834, n_8843, n_8842);
  and g22729 (n13835, \asqrt[17] , n13834);
  not g22730 (n_9230, n13835);
  and g22731 (n13836, n_8841, n_9230);
  not g22732 (n_9231, n13833);
  not g22733 (n_9232, n13836);
  and g22734 (n13837, n_9231, n_9232);
  and g22735 (n13838, n_1842, n_9227);
  and g22736 (n13839, n_9228, n13838);
  not g22737 (n_9233, n13837);
  not g22738 (n_9234, n13839);
  and g22739 (n13840, n_9233, n_9234);
  not g22740 (n_9235, n13830);
  not g22741 (n_9236, n13840);
  and g22742 (n13841, n_9235, n_9236);
  not g22743 (n_9237, n13841);
  and g22744 (n13842, \asqrt[46] , n_9237);
  and g22748 (n13846, n_8851, n_8850);
  and g22749 (n13847, \asqrt[17] , n13846);
  not g22750 (n_9238, n13847);
  and g22751 (n13848, n_8849, n_9238);
  not g22752 (n_9239, n13845);
  not g22753 (n_9240, n13848);
  and g22754 (n13849, n_9239, n_9240);
  and g22755 (n13850, n_1674, n_9235);
  and g22756 (n13851, n_9236, n13850);
  not g22757 (n_9241, n13849);
  not g22758 (n_9242, n13851);
  and g22759 (n13852, n_9241, n_9242);
  not g22760 (n_9243, n13842);
  not g22761 (n_9244, n13852);
  and g22762 (n13853, n_9243, n_9244);
  not g22763 (n_9245, n13853);
  and g22764 (n13854, \asqrt[47] , n_9245);
  and g22768 (n13858, n_8859, n_8858);
  and g22769 (n13859, \asqrt[17] , n13858);
  not g22770 (n_9246, n13859);
  and g22771 (n13860, n_8857, n_9246);
  not g22772 (n_9247, n13857);
  not g22773 (n_9248, n13860);
  and g22774 (n13861, n_9247, n_9248);
  and g22775 (n13862, n_1514, n_9243);
  and g22776 (n13863, n_9244, n13862);
  not g22777 (n_9249, n13861);
  not g22778 (n_9250, n13863);
  and g22779 (n13864, n_9249, n_9250);
  not g22780 (n_9251, n13854);
  not g22781 (n_9252, n13864);
  and g22782 (n13865, n_9251, n_9252);
  not g22783 (n_9253, n13865);
  and g22784 (n13866, \asqrt[48] , n_9253);
  and g22785 (n13867, n_1362, n_9251);
  and g22786 (n13868, n_9252, n13867);
  and g22790 (n13872, n_8867, n_8865);
  and g22791 (n13873, \asqrt[17] , n13872);
  not g22792 (n_9254, n13873);
  and g22793 (n13874, n_8866, n_9254);
  not g22794 (n_9255, n13871);
  not g22795 (n_9256, n13874);
  and g22796 (n13875, n_9255, n_9256);
  not g22797 (n_9257, n13868);
  not g22798 (n_9258, n13875);
  and g22799 (n13876, n_9257, n_9258);
  not g22800 (n_9259, n13866);
  not g22801 (n_9260, n13876);
  and g22802 (n13877, n_9259, n_9260);
  not g22803 (n_9261, n13877);
  and g22804 (n13878, \asqrt[49] , n_9261);
  and g22808 (n13882, n_8875, n_8874);
  and g22809 (n13883, \asqrt[17] , n13882);
  not g22810 (n_9262, n13883);
  and g22811 (n13884, n_8873, n_9262);
  not g22812 (n_9263, n13881);
  not g22813 (n_9264, n13884);
  and g22814 (n13885, n_9263, n_9264);
  and g22815 (n13886, n_1218, n_9259);
  and g22816 (n13887, n_9260, n13886);
  not g22817 (n_9265, n13885);
  not g22818 (n_9266, n13887);
  and g22819 (n13888, n_9265, n_9266);
  not g22820 (n_9267, n13878);
  not g22821 (n_9268, n13888);
  and g22822 (n13889, n_9267, n_9268);
  not g22823 (n_9269, n13889);
  and g22824 (n13890, \asqrt[50] , n_9269);
  and g22828 (n13894, n_8883, n_8882);
  and g22829 (n13895, \asqrt[17] , n13894);
  not g22830 (n_9270, n13895);
  and g22831 (n13896, n_8881, n_9270);
  not g22832 (n_9271, n13893);
  not g22833 (n_9272, n13896);
  and g22834 (n13897, n_9271, n_9272);
  and g22835 (n13898, n_1082, n_9267);
  and g22836 (n13899, n_9268, n13898);
  not g22837 (n_9273, n13897);
  not g22838 (n_9274, n13899);
  and g22839 (n13900, n_9273, n_9274);
  not g22840 (n_9275, n13890);
  not g22841 (n_9276, n13900);
  and g22842 (n13901, n_9275, n_9276);
  not g22843 (n_9277, n13901);
  and g22844 (n13902, \asqrt[51] , n_9277);
  and g22848 (n13906, n_8891, n_8890);
  and g22849 (n13907, \asqrt[17] , n13906);
  not g22850 (n_9278, n13907);
  and g22851 (n13908, n_8889, n_9278);
  not g22852 (n_9279, n13905);
  not g22853 (n_9280, n13908);
  and g22854 (n13909, n_9279, n_9280);
  and g22855 (n13910, n_954, n_9275);
  and g22856 (n13911, n_9276, n13910);
  not g22857 (n_9281, n13909);
  not g22858 (n_9282, n13911);
  and g22859 (n13912, n_9281, n_9282);
  not g22860 (n_9283, n13902);
  not g22861 (n_9284, n13912);
  and g22862 (n13913, n_9283, n_9284);
  not g22863 (n_9285, n13913);
  and g22864 (n13914, \asqrt[52] , n_9285);
  and g22868 (n13918, n_8899, n_8898);
  and g22869 (n13919, \asqrt[17] , n13918);
  not g22870 (n_9286, n13919);
  and g22871 (n13920, n_8897, n_9286);
  not g22872 (n_9287, n13917);
  not g22873 (n_9288, n13920);
  and g22874 (n13921, n_9287, n_9288);
  and g22875 (n13922, n_834, n_9283);
  and g22876 (n13923, n_9284, n13922);
  not g22877 (n_9289, n13921);
  not g22878 (n_9290, n13923);
  and g22879 (n13924, n_9289, n_9290);
  not g22880 (n_9291, n13914);
  not g22881 (n_9292, n13924);
  and g22882 (n13925, n_9291, n_9292);
  not g22883 (n_9293, n13925);
  and g22884 (n13926, \asqrt[53] , n_9293);
  and g22888 (n13930, n_8907, n_8906);
  and g22889 (n13931, \asqrt[17] , n13930);
  not g22890 (n_9294, n13931);
  and g22891 (n13932, n_8905, n_9294);
  not g22892 (n_9295, n13929);
  not g22893 (n_9296, n13932);
  and g22894 (n13933, n_9295, n_9296);
  and g22895 (n13934, n_722, n_9291);
  and g22896 (n13935, n_9292, n13934);
  not g22897 (n_9297, n13933);
  not g22898 (n_9298, n13935);
  and g22899 (n13936, n_9297, n_9298);
  not g22900 (n_9299, n13926);
  not g22901 (n_9300, n13936);
  and g22902 (n13937, n_9299, n_9300);
  not g22903 (n_9301, n13937);
  and g22904 (n13938, \asqrt[54] , n_9301);
  and g22908 (n13942, n_8915, n_8914);
  and g22909 (n13943, \asqrt[17] , n13942);
  not g22910 (n_9302, n13943);
  and g22911 (n13944, n_8913, n_9302);
  not g22912 (n_9303, n13941);
  not g22913 (n_9304, n13944);
  and g22914 (n13945, n_9303, n_9304);
  and g22915 (n13946, n_618, n_9299);
  and g22916 (n13947, n_9300, n13946);
  not g22917 (n_9305, n13945);
  not g22918 (n_9306, n13947);
  and g22919 (n13948, n_9305, n_9306);
  not g22920 (n_9307, n13938);
  not g22921 (n_9308, n13948);
  and g22922 (n13949, n_9307, n_9308);
  not g22923 (n_9309, n13949);
  and g22924 (n13950, \asqrt[55] , n_9309);
  and g22928 (n13954, n_8923, n_8922);
  and g22929 (n13955, \asqrt[17] , n13954);
  not g22930 (n_9310, n13955);
  and g22931 (n13956, n_8921, n_9310);
  not g22932 (n_9311, n13953);
  not g22933 (n_9312, n13956);
  and g22934 (n13957, n_9311, n_9312);
  and g22935 (n13958, n_522, n_9307);
  and g22936 (n13959, n_9308, n13958);
  not g22937 (n_9313, n13957);
  not g22938 (n_9314, n13959);
  and g22939 (n13960, n_9313, n_9314);
  not g22940 (n_9315, n13950);
  not g22941 (n_9316, n13960);
  and g22942 (n13961, n_9315, n_9316);
  not g22943 (n_9317, n13961);
  and g22944 (n13962, \asqrt[56] , n_9317);
  and g22948 (n13966, n_8931, n_8930);
  and g22949 (n13967, \asqrt[17] , n13966);
  not g22950 (n_9318, n13967);
  and g22951 (n13968, n_8929, n_9318);
  not g22952 (n_9319, n13965);
  not g22953 (n_9320, n13968);
  and g22954 (n13969, n_9319, n_9320);
  and g22955 (n13970, n_434, n_9315);
  and g22956 (n13971, n_9316, n13970);
  not g22957 (n_9321, n13969);
  not g22958 (n_9322, n13971);
  and g22959 (n13972, n_9321, n_9322);
  not g22960 (n_9323, n13962);
  not g22961 (n_9324, n13972);
  and g22962 (n13973, n_9323, n_9324);
  not g22963 (n_9325, n13973);
  and g22964 (n13974, \asqrt[57] , n_9325);
  and g22968 (n13978, n_8939, n_8938);
  and g22969 (n13979, \asqrt[17] , n13978);
  not g22970 (n_9326, n13979);
  and g22971 (n13980, n_8937, n_9326);
  not g22972 (n_9327, n13977);
  not g22973 (n_9328, n13980);
  and g22974 (n13981, n_9327, n_9328);
  and g22975 (n13982, n_354, n_9323);
  and g22976 (n13983, n_9324, n13982);
  not g22977 (n_9329, n13981);
  not g22978 (n_9330, n13983);
  and g22979 (n13984, n_9329, n_9330);
  not g22980 (n_9331, n13974);
  not g22981 (n_9332, n13984);
  and g22982 (n13985, n_9331, n_9332);
  not g22983 (n_9333, n13985);
  and g22984 (n13986, \asqrt[58] , n_9333);
  and g22988 (n13990, n_8947, n_8946);
  and g22989 (n13991, \asqrt[17] , n13990);
  not g22990 (n_9334, n13991);
  and g22991 (n13992, n_8945, n_9334);
  not g22992 (n_9335, n13989);
  not g22993 (n_9336, n13992);
  and g22994 (n13993, n_9335, n_9336);
  and g22995 (n13994, n_282, n_9331);
  and g22996 (n13995, n_9332, n13994);
  not g22997 (n_9337, n13993);
  not g22998 (n_9338, n13995);
  and g22999 (n13996, n_9337, n_9338);
  not g23000 (n_9339, n13986);
  not g23001 (n_9340, n13996);
  and g23002 (n13997, n_9339, n_9340);
  not g23003 (n_9341, n13997);
  and g23004 (n13998, \asqrt[59] , n_9341);
  and g23008 (n14002, n_8955, n_8954);
  and g23009 (n14003, \asqrt[17] , n14002);
  not g23010 (n_9342, n14003);
  and g23011 (n14004, n_8953, n_9342);
  not g23012 (n_9343, n14001);
  not g23013 (n_9344, n14004);
  and g23014 (n14005, n_9343, n_9344);
  and g23015 (n14006, n_218, n_9339);
  and g23016 (n14007, n_9340, n14006);
  not g23017 (n_9345, n14005);
  not g23018 (n_9346, n14007);
  and g23019 (n14008, n_9345, n_9346);
  not g23020 (n_9347, n13998);
  not g23021 (n_9348, n14008);
  and g23022 (n14009, n_9347, n_9348);
  not g23023 (n_9349, n14009);
  and g23024 (n14010, \asqrt[60] , n_9349);
  and g23028 (n14014, n_8963, n_8962);
  and g23029 (n14015, \asqrt[17] , n14014);
  not g23030 (n_9350, n14015);
  and g23031 (n14016, n_8961, n_9350);
  not g23032 (n_9351, n14013);
  not g23033 (n_9352, n14016);
  and g23034 (n14017, n_9351, n_9352);
  and g23035 (n14018, n_162, n_9347);
  and g23036 (n14019, n_9348, n14018);
  not g23037 (n_9353, n14017);
  not g23038 (n_9354, n14019);
  and g23039 (n14020, n_9353, n_9354);
  not g23040 (n_9355, n14010);
  not g23041 (n_9356, n14020);
  and g23042 (n14021, n_9355, n_9356);
  not g23043 (n_9357, n14021);
  and g23044 (n14022, \asqrt[61] , n_9357);
  and g23048 (n14026, n_8971, n_8970);
  and g23049 (n14027, \asqrt[17] , n14026);
  not g23050 (n_9358, n14027);
  and g23051 (n14028, n_8969, n_9358);
  not g23052 (n_9359, n14025);
  not g23053 (n_9360, n14028);
  and g23054 (n14029, n_9359, n_9360);
  and g23055 (n14030, n_115, n_9355);
  and g23056 (n14031, n_9356, n14030);
  not g23057 (n_9361, n14029);
  not g23058 (n_9362, n14031);
  and g23059 (n14032, n_9361, n_9362);
  not g23060 (n_9363, n14022);
  not g23061 (n_9364, n14032);
  and g23062 (n14033, n_9363, n_9364);
  not g23063 (n_9365, n14033);
  and g23064 (n14034, \asqrt[62] , n_9365);
  and g23068 (n14038, n_8979, n_8978);
  and g23069 (n14039, \asqrt[17] , n14038);
  not g23070 (n_9366, n14039);
  and g23071 (n14040, n_8977, n_9366);
  not g23072 (n_9367, n14037);
  not g23073 (n_9368, n14040);
  and g23074 (n14041, n_9367, n_9368);
  and g23075 (n14042, n_76, n_9363);
  and g23076 (n14043, n_9364, n14042);
  not g23077 (n_9369, n14041);
  not g23078 (n_9370, n14043);
  and g23079 (n14044, n_9369, n_9370);
  not g23080 (n_9371, n14034);
  not g23081 (n_9372, n14044);
  and g23082 (n14045, n_9371, n_9372);
  and g23086 (n14049, n_8987, n_8986);
  and g23087 (n14050, \asqrt[17] , n14049);
  not g23088 (n_9373, n14050);
  and g23089 (n14051, n_8985, n_9373);
  not g23090 (n_9374, n14048);
  not g23091 (n_9375, n14051);
  and g23092 (n14052, n_9374, n_9375);
  and g23093 (n14053, n_8994, n_8993);
  and g23094 (n14054, \asqrt[17] , n14053);
  not g23097 (n_9377, n14052);
  not g23099 (n_9378, n14045);
  not g23101 (n_9379, n14057);
  and g23102 (n14058, n_21, n_9379);
  and g23103 (n14059, n_9371, n14052);
  and g23104 (n14060, n_9372, n14059);
  and g23105 (n14061, n_8993, \asqrt[17] );
  not g23106 (n_9380, n14061);
  and g23107 (n14062, n13473, n_9380);
  not g23108 (n_9381, n14053);
  and g23109 (n14063, \asqrt[63] , n_9381);
  not g23110 (n_9382, n14062);
  and g23111 (n14064, n_9382, n14063);
  not g23117 (n_9383, n14064);
  not g23118 (n_9384, n14069);
  not g23120 (n_9385, n14060);
  and g23124 (n14073, \a[32] , \asqrt[16] );
  not g23125 (n_9390, \a[30] );
  not g23126 (n_9391, \a[31] );
  and g23127 (n14074, n_9390, n_9391);
  and g23128 (n14075, n_9006, n14074);
  not g23129 (n_9392, n14073);
  not g23130 (n_9393, n14075);
  and g23131 (n14076, n_9392, n_9393);
  not g23132 (n_9394, n14076);
  and g23133 (n14077, \asqrt[17] , n_9394);
  and g23139 (n14083, n_9006, \asqrt[16] );
  not g23140 (n_9395, n14083);
  and g23141 (n14084, \a[33] , n_9395);
  and g23142 (n14085, n13502, \asqrt[16] );
  not g23143 (n_9396, n14084);
  not g23144 (n_9397, n14085);
  and g23145 (n14086, n_9396, n_9397);
  not g23146 (n_9398, n14082);
  and g23147 (n14087, n_9398, n14086);
  not g23148 (n_9399, n14077);
  not g23149 (n_9400, n14087);
  and g23150 (n14088, n_9399, n_9400);
  not g23151 (n_9401, n14088);
  and g23152 (n14089, \asqrt[18] , n_9401);
  not g23153 (n_9402, \asqrt[18] );
  and g23154 (n14090, n_9402, n_9399);
  and g23155 (n14091, n_9400, n14090);
  not g23159 (n_9403, n14058);
  not g23161 (n_9404, n14095);
  and g23162 (n14096, n_9397, n_9404);
  not g23163 (n_9405, n14096);
  and g23164 (n14097, \a[34] , n_9405);
  and g23165 (n14098, n_8630, n_9404);
  and g23166 (n14099, n_9397, n14098);
  not g23167 (n_9406, n14097);
  not g23168 (n_9407, n14099);
  and g23169 (n14100, n_9406, n_9407);
  not g23170 (n_9408, n14091);
  not g23171 (n_9409, n14100);
  and g23172 (n14101, n_9408, n_9409);
  not g23173 (n_9410, n14089);
  not g23174 (n_9411, n14101);
  and g23175 (n14102, n_9410, n_9411);
  not g23176 (n_9412, n14102);
  and g23177 (n14103, \asqrt[19] , n_9412);
  and g23178 (n14104, n_9015, n_9014);
  not g23179 (n_9413, n13514);
  and g23180 (n14105, n_9413, n14104);
  and g23181 (n14106, \asqrt[16] , n14105);
  and g23182 (n14107, \asqrt[16] , n14104);
  not g23183 (n_9414, n14107);
  and g23184 (n14108, n13514, n_9414);
  not g23185 (n_9415, n14106);
  not g23186 (n_9416, n14108);
  and g23187 (n14109, n_9415, n_9416);
  and g23188 (n14110, n_9018, n_9410);
  and g23189 (n14111, n_9411, n14110);
  not g23190 (n_9417, n14109);
  not g23191 (n_9418, n14111);
  and g23192 (n14112, n_9417, n_9418);
  not g23193 (n_9419, n14103);
  not g23194 (n_9420, n14112);
  and g23195 (n14113, n_9419, n_9420);
  not g23196 (n_9421, n14113);
  and g23197 (n14114, \asqrt[20] , n_9421);
  and g23201 (n14118, n_9026, n_9024);
  and g23202 (n14119, \asqrt[16] , n14118);
  not g23203 (n_9422, n14119);
  and g23204 (n14120, n_9025, n_9422);
  not g23205 (n_9423, n14117);
  not g23206 (n_9424, n14120);
  and g23207 (n14121, n_9423, n_9424);
  and g23208 (n14122, n_8642, n_9419);
  and g23209 (n14123, n_9420, n14122);
  not g23210 (n_9425, n14121);
  not g23211 (n_9426, n14123);
  and g23212 (n14124, n_9425, n_9426);
  not g23213 (n_9427, n14114);
  not g23214 (n_9428, n14124);
  and g23215 (n14125, n_9427, n_9428);
  not g23216 (n_9429, n14125);
  and g23217 (n14126, \asqrt[21] , n_9429);
  and g23221 (n14130, n_9035, n_9034);
  and g23222 (n14131, \asqrt[16] , n14130);
  not g23223 (n_9430, n14131);
  and g23224 (n14132, n_9033, n_9430);
  not g23225 (n_9431, n14129);
  not g23226 (n_9432, n14132);
  and g23227 (n14133, n_9431, n_9432);
  and g23228 (n14134, n_8274, n_9427);
  and g23229 (n14135, n_9428, n14134);
  not g23230 (n_9433, n14133);
  not g23231 (n_9434, n14135);
  and g23232 (n14136, n_9433, n_9434);
  not g23233 (n_9435, n14126);
  not g23234 (n_9436, n14136);
  and g23235 (n14137, n_9435, n_9436);
  not g23236 (n_9437, n14137);
  and g23237 (n14138, \asqrt[22] , n_9437);
  and g23241 (n14142, n_9043, n_9042);
  and g23242 (n14143, \asqrt[16] , n14142);
  not g23243 (n_9438, n14143);
  and g23244 (n14144, n_9041, n_9438);
  not g23245 (n_9439, n14141);
  not g23246 (n_9440, n14144);
  and g23247 (n14145, n_9439, n_9440);
  and g23248 (n14146, n_7914, n_9435);
  and g23249 (n14147, n_9436, n14146);
  not g23250 (n_9441, n14145);
  not g23251 (n_9442, n14147);
  and g23252 (n14148, n_9441, n_9442);
  not g23253 (n_9443, n14138);
  not g23254 (n_9444, n14148);
  and g23255 (n14149, n_9443, n_9444);
  not g23256 (n_9445, n14149);
  and g23257 (n14150, \asqrt[23] , n_9445);
  and g23261 (n14154, n_9051, n_9050);
  and g23262 (n14155, \asqrt[16] , n14154);
  not g23263 (n_9446, n14155);
  and g23264 (n14156, n_9049, n_9446);
  not g23265 (n_9447, n14153);
  not g23266 (n_9448, n14156);
  and g23267 (n14157, n_9447, n_9448);
  and g23268 (n14158, n_7562, n_9443);
  and g23269 (n14159, n_9444, n14158);
  not g23270 (n_9449, n14157);
  not g23271 (n_9450, n14159);
  and g23272 (n14160, n_9449, n_9450);
  not g23273 (n_9451, n14150);
  not g23274 (n_9452, n14160);
  and g23275 (n14161, n_9451, n_9452);
  not g23276 (n_9453, n14161);
  and g23277 (n14162, \asqrt[24] , n_9453);
  and g23281 (n14166, n_9059, n_9058);
  and g23282 (n14167, \asqrt[16] , n14166);
  not g23283 (n_9454, n14167);
  and g23284 (n14168, n_9057, n_9454);
  not g23285 (n_9455, n14165);
  not g23286 (n_9456, n14168);
  and g23287 (n14169, n_9455, n_9456);
  and g23288 (n14170, n_7218, n_9451);
  and g23289 (n14171, n_9452, n14170);
  not g23290 (n_9457, n14169);
  not g23291 (n_9458, n14171);
  and g23292 (n14172, n_9457, n_9458);
  not g23293 (n_9459, n14162);
  not g23294 (n_9460, n14172);
  and g23295 (n14173, n_9459, n_9460);
  not g23296 (n_9461, n14173);
  and g23297 (n14174, \asqrt[25] , n_9461);
  and g23301 (n14178, n_9067, n_9066);
  and g23302 (n14179, \asqrt[16] , n14178);
  not g23303 (n_9462, n14179);
  and g23304 (n14180, n_9065, n_9462);
  not g23305 (n_9463, n14177);
  not g23306 (n_9464, n14180);
  and g23307 (n14181, n_9463, n_9464);
  and g23308 (n14182, n_6882, n_9459);
  and g23309 (n14183, n_9460, n14182);
  not g23310 (n_9465, n14181);
  not g23311 (n_9466, n14183);
  and g23312 (n14184, n_9465, n_9466);
  not g23313 (n_9467, n14174);
  not g23314 (n_9468, n14184);
  and g23315 (n14185, n_9467, n_9468);
  not g23316 (n_9469, n14185);
  and g23317 (n14186, \asqrt[26] , n_9469);
  and g23321 (n14190, n_9075, n_9074);
  and g23322 (n14191, \asqrt[16] , n14190);
  not g23323 (n_9470, n14191);
  and g23324 (n14192, n_9073, n_9470);
  not g23325 (n_9471, n14189);
  not g23326 (n_9472, n14192);
  and g23327 (n14193, n_9471, n_9472);
  and g23328 (n14194, n_6554, n_9467);
  and g23329 (n14195, n_9468, n14194);
  not g23330 (n_9473, n14193);
  not g23331 (n_9474, n14195);
  and g23332 (n14196, n_9473, n_9474);
  not g23333 (n_9475, n14186);
  not g23334 (n_9476, n14196);
  and g23335 (n14197, n_9475, n_9476);
  not g23336 (n_9477, n14197);
  and g23337 (n14198, \asqrt[27] , n_9477);
  and g23341 (n14202, n_9083, n_9082);
  and g23342 (n14203, \asqrt[16] , n14202);
  not g23343 (n_9478, n14203);
  and g23344 (n14204, n_9081, n_9478);
  not g23345 (n_9479, n14201);
  not g23346 (n_9480, n14204);
  and g23347 (n14205, n_9479, n_9480);
  and g23348 (n14206, n_6234, n_9475);
  and g23349 (n14207, n_9476, n14206);
  not g23350 (n_9481, n14205);
  not g23351 (n_9482, n14207);
  and g23352 (n14208, n_9481, n_9482);
  not g23353 (n_9483, n14198);
  not g23354 (n_9484, n14208);
  and g23355 (n14209, n_9483, n_9484);
  not g23356 (n_9485, n14209);
  and g23357 (n14210, \asqrt[28] , n_9485);
  and g23361 (n14214, n_9091, n_9090);
  and g23362 (n14215, \asqrt[16] , n14214);
  not g23363 (n_9486, n14215);
  and g23364 (n14216, n_9089, n_9486);
  not g23365 (n_9487, n14213);
  not g23366 (n_9488, n14216);
  and g23367 (n14217, n_9487, n_9488);
  and g23368 (n14218, n_5922, n_9483);
  and g23369 (n14219, n_9484, n14218);
  not g23370 (n_9489, n14217);
  not g23371 (n_9490, n14219);
  and g23372 (n14220, n_9489, n_9490);
  not g23373 (n_9491, n14210);
  not g23374 (n_9492, n14220);
  and g23375 (n14221, n_9491, n_9492);
  not g23376 (n_9493, n14221);
  and g23377 (n14222, \asqrt[29] , n_9493);
  and g23381 (n14226, n_9099, n_9098);
  and g23382 (n14227, \asqrt[16] , n14226);
  not g23383 (n_9494, n14227);
  and g23384 (n14228, n_9097, n_9494);
  not g23385 (n_9495, n14225);
  not g23386 (n_9496, n14228);
  and g23387 (n14229, n_9495, n_9496);
  and g23388 (n14230, n_5618, n_9491);
  and g23389 (n14231, n_9492, n14230);
  not g23390 (n_9497, n14229);
  not g23391 (n_9498, n14231);
  and g23392 (n14232, n_9497, n_9498);
  not g23393 (n_9499, n14222);
  not g23394 (n_9500, n14232);
  and g23395 (n14233, n_9499, n_9500);
  not g23396 (n_9501, n14233);
  and g23397 (n14234, \asqrt[30] , n_9501);
  and g23401 (n14238, n_9107, n_9106);
  and g23402 (n14239, \asqrt[16] , n14238);
  not g23403 (n_9502, n14239);
  and g23404 (n14240, n_9105, n_9502);
  not g23405 (n_9503, n14237);
  not g23406 (n_9504, n14240);
  and g23407 (n14241, n_9503, n_9504);
  and g23408 (n14242, n_5322, n_9499);
  and g23409 (n14243, n_9500, n14242);
  not g23410 (n_9505, n14241);
  not g23411 (n_9506, n14243);
  and g23412 (n14244, n_9505, n_9506);
  not g23413 (n_9507, n14234);
  not g23414 (n_9508, n14244);
  and g23415 (n14245, n_9507, n_9508);
  not g23416 (n_9509, n14245);
  and g23417 (n14246, \asqrt[31] , n_9509);
  and g23421 (n14250, n_9115, n_9114);
  and g23422 (n14251, \asqrt[16] , n14250);
  not g23423 (n_9510, n14251);
  and g23424 (n14252, n_9113, n_9510);
  not g23425 (n_9511, n14249);
  not g23426 (n_9512, n14252);
  and g23427 (n14253, n_9511, n_9512);
  and g23428 (n14254, n_5034, n_9507);
  and g23429 (n14255, n_9508, n14254);
  not g23430 (n_9513, n14253);
  not g23431 (n_9514, n14255);
  and g23432 (n14256, n_9513, n_9514);
  not g23433 (n_9515, n14246);
  not g23434 (n_9516, n14256);
  and g23435 (n14257, n_9515, n_9516);
  not g23436 (n_9517, n14257);
  and g23437 (n14258, \asqrt[32] , n_9517);
  and g23441 (n14262, n_9123, n_9122);
  and g23442 (n14263, \asqrt[16] , n14262);
  not g23443 (n_9518, n14263);
  and g23444 (n14264, n_9121, n_9518);
  not g23445 (n_9519, n14261);
  not g23446 (n_9520, n14264);
  and g23447 (n14265, n_9519, n_9520);
  and g23448 (n14266, n_4754, n_9515);
  and g23449 (n14267, n_9516, n14266);
  not g23450 (n_9521, n14265);
  not g23451 (n_9522, n14267);
  and g23452 (n14268, n_9521, n_9522);
  not g23453 (n_9523, n14258);
  not g23454 (n_9524, n14268);
  and g23455 (n14269, n_9523, n_9524);
  not g23456 (n_9525, n14269);
  and g23457 (n14270, \asqrt[33] , n_9525);
  and g23461 (n14274, n_9131, n_9130);
  and g23462 (n14275, \asqrt[16] , n14274);
  not g23463 (n_9526, n14275);
  and g23464 (n14276, n_9129, n_9526);
  not g23465 (n_9527, n14273);
  not g23466 (n_9528, n14276);
  and g23467 (n14277, n_9527, n_9528);
  and g23468 (n14278, n_4482, n_9523);
  and g23469 (n14279, n_9524, n14278);
  not g23470 (n_9529, n14277);
  not g23471 (n_9530, n14279);
  and g23472 (n14280, n_9529, n_9530);
  not g23473 (n_9531, n14270);
  not g23474 (n_9532, n14280);
  and g23475 (n14281, n_9531, n_9532);
  not g23476 (n_9533, n14281);
  and g23477 (n14282, \asqrt[34] , n_9533);
  and g23481 (n14286, n_9139, n_9138);
  and g23482 (n14287, \asqrt[16] , n14286);
  not g23483 (n_9534, n14287);
  and g23484 (n14288, n_9137, n_9534);
  not g23485 (n_9535, n14285);
  not g23486 (n_9536, n14288);
  and g23487 (n14289, n_9535, n_9536);
  and g23488 (n14290, n_4218, n_9531);
  and g23489 (n14291, n_9532, n14290);
  not g23490 (n_9537, n14289);
  not g23491 (n_9538, n14291);
  and g23492 (n14292, n_9537, n_9538);
  not g23493 (n_9539, n14282);
  not g23494 (n_9540, n14292);
  and g23495 (n14293, n_9539, n_9540);
  not g23496 (n_9541, n14293);
  and g23497 (n14294, \asqrt[35] , n_9541);
  and g23501 (n14298, n_9147, n_9146);
  and g23502 (n14299, \asqrt[16] , n14298);
  not g23503 (n_9542, n14299);
  and g23504 (n14300, n_9145, n_9542);
  not g23505 (n_9543, n14297);
  not g23506 (n_9544, n14300);
  and g23507 (n14301, n_9543, n_9544);
  and g23508 (n14302, n_3962, n_9539);
  and g23509 (n14303, n_9540, n14302);
  not g23510 (n_9545, n14301);
  not g23511 (n_9546, n14303);
  and g23512 (n14304, n_9545, n_9546);
  not g23513 (n_9547, n14294);
  not g23514 (n_9548, n14304);
  and g23515 (n14305, n_9547, n_9548);
  not g23516 (n_9549, n14305);
  and g23517 (n14306, \asqrt[36] , n_9549);
  and g23521 (n14310, n_9155, n_9154);
  and g23522 (n14311, \asqrt[16] , n14310);
  not g23523 (n_9550, n14311);
  and g23524 (n14312, n_9153, n_9550);
  not g23525 (n_9551, n14309);
  not g23526 (n_9552, n14312);
  and g23527 (n14313, n_9551, n_9552);
  and g23528 (n14314, n_3714, n_9547);
  and g23529 (n14315, n_9548, n14314);
  not g23530 (n_9553, n14313);
  not g23531 (n_9554, n14315);
  and g23532 (n14316, n_9553, n_9554);
  not g23533 (n_9555, n14306);
  not g23534 (n_9556, n14316);
  and g23535 (n14317, n_9555, n_9556);
  not g23536 (n_9557, n14317);
  and g23537 (n14318, \asqrt[37] , n_9557);
  and g23541 (n14322, n_9163, n_9162);
  and g23542 (n14323, \asqrt[16] , n14322);
  not g23543 (n_9558, n14323);
  and g23544 (n14324, n_9161, n_9558);
  not g23545 (n_9559, n14321);
  not g23546 (n_9560, n14324);
  and g23547 (n14325, n_9559, n_9560);
  and g23548 (n14326, n_3474, n_9555);
  and g23549 (n14327, n_9556, n14326);
  not g23550 (n_9561, n14325);
  not g23551 (n_9562, n14327);
  and g23552 (n14328, n_9561, n_9562);
  not g23553 (n_9563, n14318);
  not g23554 (n_9564, n14328);
  and g23555 (n14329, n_9563, n_9564);
  not g23556 (n_9565, n14329);
  and g23557 (n14330, \asqrt[38] , n_9565);
  and g23561 (n14334, n_9171, n_9170);
  and g23562 (n14335, \asqrt[16] , n14334);
  not g23563 (n_9566, n14335);
  and g23564 (n14336, n_9169, n_9566);
  not g23565 (n_9567, n14333);
  not g23566 (n_9568, n14336);
  and g23567 (n14337, n_9567, n_9568);
  and g23568 (n14338, n_3242, n_9563);
  and g23569 (n14339, n_9564, n14338);
  not g23570 (n_9569, n14337);
  not g23571 (n_9570, n14339);
  and g23572 (n14340, n_9569, n_9570);
  not g23573 (n_9571, n14330);
  not g23574 (n_9572, n14340);
  and g23575 (n14341, n_9571, n_9572);
  not g23576 (n_9573, n14341);
  and g23577 (n14342, \asqrt[39] , n_9573);
  and g23581 (n14346, n_9179, n_9178);
  and g23582 (n14347, \asqrt[16] , n14346);
  not g23583 (n_9574, n14347);
  and g23584 (n14348, n_9177, n_9574);
  not g23585 (n_9575, n14345);
  not g23586 (n_9576, n14348);
  and g23587 (n14349, n_9575, n_9576);
  and g23588 (n14350, n_3018, n_9571);
  and g23589 (n14351, n_9572, n14350);
  not g23590 (n_9577, n14349);
  not g23591 (n_9578, n14351);
  and g23592 (n14352, n_9577, n_9578);
  not g23593 (n_9579, n14342);
  not g23594 (n_9580, n14352);
  and g23595 (n14353, n_9579, n_9580);
  not g23596 (n_9581, n14353);
  and g23597 (n14354, \asqrt[40] , n_9581);
  and g23601 (n14358, n_9187, n_9186);
  and g23602 (n14359, \asqrt[16] , n14358);
  not g23603 (n_9582, n14359);
  and g23604 (n14360, n_9185, n_9582);
  not g23605 (n_9583, n14357);
  not g23606 (n_9584, n14360);
  and g23607 (n14361, n_9583, n_9584);
  and g23608 (n14362, n_2802, n_9579);
  and g23609 (n14363, n_9580, n14362);
  not g23610 (n_9585, n14361);
  not g23611 (n_9586, n14363);
  and g23612 (n14364, n_9585, n_9586);
  not g23613 (n_9587, n14354);
  not g23614 (n_9588, n14364);
  and g23615 (n14365, n_9587, n_9588);
  not g23616 (n_9589, n14365);
  and g23617 (n14366, \asqrt[41] , n_9589);
  and g23621 (n14370, n_9195, n_9194);
  and g23622 (n14371, \asqrt[16] , n14370);
  not g23623 (n_9590, n14371);
  and g23624 (n14372, n_9193, n_9590);
  not g23625 (n_9591, n14369);
  not g23626 (n_9592, n14372);
  and g23627 (n14373, n_9591, n_9592);
  and g23628 (n14374, n_2594, n_9587);
  and g23629 (n14375, n_9588, n14374);
  not g23630 (n_9593, n14373);
  not g23631 (n_9594, n14375);
  and g23632 (n14376, n_9593, n_9594);
  not g23633 (n_9595, n14366);
  not g23634 (n_9596, n14376);
  and g23635 (n14377, n_9595, n_9596);
  not g23636 (n_9597, n14377);
  and g23637 (n14378, \asqrt[42] , n_9597);
  and g23641 (n14382, n_9203, n_9202);
  and g23642 (n14383, \asqrt[16] , n14382);
  not g23643 (n_9598, n14383);
  and g23644 (n14384, n_9201, n_9598);
  not g23645 (n_9599, n14381);
  not g23646 (n_9600, n14384);
  and g23647 (n14385, n_9599, n_9600);
  and g23648 (n14386, n_2394, n_9595);
  and g23649 (n14387, n_9596, n14386);
  not g23650 (n_9601, n14385);
  not g23651 (n_9602, n14387);
  and g23652 (n14388, n_9601, n_9602);
  not g23653 (n_9603, n14378);
  not g23654 (n_9604, n14388);
  and g23655 (n14389, n_9603, n_9604);
  not g23656 (n_9605, n14389);
  and g23657 (n14390, \asqrt[43] , n_9605);
  and g23661 (n14394, n_9211, n_9210);
  and g23662 (n14395, \asqrt[16] , n14394);
  not g23663 (n_9606, n14395);
  and g23664 (n14396, n_9209, n_9606);
  not g23665 (n_9607, n14393);
  not g23666 (n_9608, n14396);
  and g23667 (n14397, n_9607, n_9608);
  and g23668 (n14398, n_2202, n_9603);
  and g23669 (n14399, n_9604, n14398);
  not g23670 (n_9609, n14397);
  not g23671 (n_9610, n14399);
  and g23672 (n14400, n_9609, n_9610);
  not g23673 (n_9611, n14390);
  not g23674 (n_9612, n14400);
  and g23675 (n14401, n_9611, n_9612);
  not g23676 (n_9613, n14401);
  and g23677 (n14402, \asqrt[44] , n_9613);
  and g23681 (n14406, n_9219, n_9218);
  and g23682 (n14407, \asqrt[16] , n14406);
  not g23683 (n_9614, n14407);
  and g23684 (n14408, n_9217, n_9614);
  not g23685 (n_9615, n14405);
  not g23686 (n_9616, n14408);
  and g23687 (n14409, n_9615, n_9616);
  and g23688 (n14410, n_2018, n_9611);
  and g23689 (n14411, n_9612, n14410);
  not g23690 (n_9617, n14409);
  not g23691 (n_9618, n14411);
  and g23692 (n14412, n_9617, n_9618);
  not g23693 (n_9619, n14402);
  not g23694 (n_9620, n14412);
  and g23695 (n14413, n_9619, n_9620);
  not g23696 (n_9621, n14413);
  and g23697 (n14414, \asqrt[45] , n_9621);
  and g23701 (n14418, n_9227, n_9226);
  and g23702 (n14419, \asqrt[16] , n14418);
  not g23703 (n_9622, n14419);
  and g23704 (n14420, n_9225, n_9622);
  not g23705 (n_9623, n14417);
  not g23706 (n_9624, n14420);
  and g23707 (n14421, n_9623, n_9624);
  and g23708 (n14422, n_1842, n_9619);
  and g23709 (n14423, n_9620, n14422);
  not g23710 (n_9625, n14421);
  not g23711 (n_9626, n14423);
  and g23712 (n14424, n_9625, n_9626);
  not g23713 (n_9627, n14414);
  not g23714 (n_9628, n14424);
  and g23715 (n14425, n_9627, n_9628);
  not g23716 (n_9629, n14425);
  and g23717 (n14426, \asqrt[46] , n_9629);
  and g23721 (n14430, n_9235, n_9234);
  and g23722 (n14431, \asqrt[16] , n14430);
  not g23723 (n_9630, n14431);
  and g23724 (n14432, n_9233, n_9630);
  not g23725 (n_9631, n14429);
  not g23726 (n_9632, n14432);
  and g23727 (n14433, n_9631, n_9632);
  and g23728 (n14434, n_1674, n_9627);
  and g23729 (n14435, n_9628, n14434);
  not g23730 (n_9633, n14433);
  not g23731 (n_9634, n14435);
  and g23732 (n14436, n_9633, n_9634);
  not g23733 (n_9635, n14426);
  not g23734 (n_9636, n14436);
  and g23735 (n14437, n_9635, n_9636);
  not g23736 (n_9637, n14437);
  and g23737 (n14438, \asqrt[47] , n_9637);
  and g23741 (n14442, n_9243, n_9242);
  and g23742 (n14443, \asqrt[16] , n14442);
  not g23743 (n_9638, n14443);
  and g23744 (n14444, n_9241, n_9638);
  not g23745 (n_9639, n14441);
  not g23746 (n_9640, n14444);
  and g23747 (n14445, n_9639, n_9640);
  and g23748 (n14446, n_1514, n_9635);
  and g23749 (n14447, n_9636, n14446);
  not g23750 (n_9641, n14445);
  not g23751 (n_9642, n14447);
  and g23752 (n14448, n_9641, n_9642);
  not g23753 (n_9643, n14438);
  not g23754 (n_9644, n14448);
  and g23755 (n14449, n_9643, n_9644);
  not g23756 (n_9645, n14449);
  and g23757 (n14450, \asqrt[48] , n_9645);
  and g23761 (n14454, n_9251, n_9250);
  and g23762 (n14455, \asqrt[16] , n14454);
  not g23763 (n_9646, n14455);
  and g23764 (n14456, n_9249, n_9646);
  not g23765 (n_9647, n14453);
  not g23766 (n_9648, n14456);
  and g23767 (n14457, n_9647, n_9648);
  and g23768 (n14458, n_1362, n_9643);
  and g23769 (n14459, n_9644, n14458);
  not g23770 (n_9649, n14457);
  not g23771 (n_9650, n14459);
  and g23772 (n14460, n_9649, n_9650);
  not g23773 (n_9651, n14450);
  not g23774 (n_9652, n14460);
  and g23775 (n14461, n_9651, n_9652);
  not g23776 (n_9653, n14461);
  and g23777 (n14462, \asqrt[49] , n_9653);
  and g23778 (n14463, n_1218, n_9651);
  and g23779 (n14464, n_9652, n14463);
  and g23783 (n14468, n_9259, n_9257);
  and g23784 (n14469, \asqrt[16] , n14468);
  not g23785 (n_9654, n14469);
  and g23786 (n14470, n_9258, n_9654);
  not g23787 (n_9655, n14467);
  not g23788 (n_9656, n14470);
  and g23789 (n14471, n_9655, n_9656);
  not g23790 (n_9657, n14464);
  not g23791 (n_9658, n14471);
  and g23792 (n14472, n_9657, n_9658);
  not g23793 (n_9659, n14462);
  not g23794 (n_9660, n14472);
  and g23795 (n14473, n_9659, n_9660);
  not g23796 (n_9661, n14473);
  and g23797 (n14474, \asqrt[50] , n_9661);
  and g23801 (n14478, n_9267, n_9266);
  and g23802 (n14479, \asqrt[16] , n14478);
  not g23803 (n_9662, n14479);
  and g23804 (n14480, n_9265, n_9662);
  not g23805 (n_9663, n14477);
  not g23806 (n_9664, n14480);
  and g23807 (n14481, n_9663, n_9664);
  and g23808 (n14482, n_1082, n_9659);
  and g23809 (n14483, n_9660, n14482);
  not g23810 (n_9665, n14481);
  not g23811 (n_9666, n14483);
  and g23812 (n14484, n_9665, n_9666);
  not g23813 (n_9667, n14474);
  not g23814 (n_9668, n14484);
  and g23815 (n14485, n_9667, n_9668);
  not g23816 (n_9669, n14485);
  and g23817 (n14486, \asqrt[51] , n_9669);
  and g23821 (n14490, n_9275, n_9274);
  and g23822 (n14491, \asqrt[16] , n14490);
  not g23823 (n_9670, n14491);
  and g23824 (n14492, n_9273, n_9670);
  not g23825 (n_9671, n14489);
  not g23826 (n_9672, n14492);
  and g23827 (n14493, n_9671, n_9672);
  and g23828 (n14494, n_954, n_9667);
  and g23829 (n14495, n_9668, n14494);
  not g23830 (n_9673, n14493);
  not g23831 (n_9674, n14495);
  and g23832 (n14496, n_9673, n_9674);
  not g23833 (n_9675, n14486);
  not g23834 (n_9676, n14496);
  and g23835 (n14497, n_9675, n_9676);
  not g23836 (n_9677, n14497);
  and g23837 (n14498, \asqrt[52] , n_9677);
  and g23841 (n14502, n_9283, n_9282);
  and g23842 (n14503, \asqrt[16] , n14502);
  not g23843 (n_9678, n14503);
  and g23844 (n14504, n_9281, n_9678);
  not g23845 (n_9679, n14501);
  not g23846 (n_9680, n14504);
  and g23847 (n14505, n_9679, n_9680);
  and g23848 (n14506, n_834, n_9675);
  and g23849 (n14507, n_9676, n14506);
  not g23850 (n_9681, n14505);
  not g23851 (n_9682, n14507);
  and g23852 (n14508, n_9681, n_9682);
  not g23853 (n_9683, n14498);
  not g23854 (n_9684, n14508);
  and g23855 (n14509, n_9683, n_9684);
  not g23856 (n_9685, n14509);
  and g23857 (n14510, \asqrt[53] , n_9685);
  and g23861 (n14514, n_9291, n_9290);
  and g23862 (n14515, \asqrt[16] , n14514);
  not g23863 (n_9686, n14515);
  and g23864 (n14516, n_9289, n_9686);
  not g23865 (n_9687, n14513);
  not g23866 (n_9688, n14516);
  and g23867 (n14517, n_9687, n_9688);
  and g23868 (n14518, n_722, n_9683);
  and g23869 (n14519, n_9684, n14518);
  not g23870 (n_9689, n14517);
  not g23871 (n_9690, n14519);
  and g23872 (n14520, n_9689, n_9690);
  not g23873 (n_9691, n14510);
  not g23874 (n_9692, n14520);
  and g23875 (n14521, n_9691, n_9692);
  not g23876 (n_9693, n14521);
  and g23877 (n14522, \asqrt[54] , n_9693);
  and g23881 (n14526, n_9299, n_9298);
  and g23882 (n14527, \asqrt[16] , n14526);
  not g23883 (n_9694, n14527);
  and g23884 (n14528, n_9297, n_9694);
  not g23885 (n_9695, n14525);
  not g23886 (n_9696, n14528);
  and g23887 (n14529, n_9695, n_9696);
  and g23888 (n14530, n_618, n_9691);
  and g23889 (n14531, n_9692, n14530);
  not g23890 (n_9697, n14529);
  not g23891 (n_9698, n14531);
  and g23892 (n14532, n_9697, n_9698);
  not g23893 (n_9699, n14522);
  not g23894 (n_9700, n14532);
  and g23895 (n14533, n_9699, n_9700);
  not g23896 (n_9701, n14533);
  and g23897 (n14534, \asqrt[55] , n_9701);
  and g23901 (n14538, n_9307, n_9306);
  and g23902 (n14539, \asqrt[16] , n14538);
  not g23903 (n_9702, n14539);
  and g23904 (n14540, n_9305, n_9702);
  not g23905 (n_9703, n14537);
  not g23906 (n_9704, n14540);
  and g23907 (n14541, n_9703, n_9704);
  and g23908 (n14542, n_522, n_9699);
  and g23909 (n14543, n_9700, n14542);
  not g23910 (n_9705, n14541);
  not g23911 (n_9706, n14543);
  and g23912 (n14544, n_9705, n_9706);
  not g23913 (n_9707, n14534);
  not g23914 (n_9708, n14544);
  and g23915 (n14545, n_9707, n_9708);
  not g23916 (n_9709, n14545);
  and g23917 (n14546, \asqrt[56] , n_9709);
  and g23921 (n14550, n_9315, n_9314);
  and g23922 (n14551, \asqrt[16] , n14550);
  not g23923 (n_9710, n14551);
  and g23924 (n14552, n_9313, n_9710);
  not g23925 (n_9711, n14549);
  not g23926 (n_9712, n14552);
  and g23927 (n14553, n_9711, n_9712);
  and g23928 (n14554, n_434, n_9707);
  and g23929 (n14555, n_9708, n14554);
  not g23930 (n_9713, n14553);
  not g23931 (n_9714, n14555);
  and g23932 (n14556, n_9713, n_9714);
  not g23933 (n_9715, n14546);
  not g23934 (n_9716, n14556);
  and g23935 (n14557, n_9715, n_9716);
  not g23936 (n_9717, n14557);
  and g23937 (n14558, \asqrt[57] , n_9717);
  and g23941 (n14562, n_9323, n_9322);
  and g23942 (n14563, \asqrt[16] , n14562);
  not g23943 (n_9718, n14563);
  and g23944 (n14564, n_9321, n_9718);
  not g23945 (n_9719, n14561);
  not g23946 (n_9720, n14564);
  and g23947 (n14565, n_9719, n_9720);
  and g23948 (n14566, n_354, n_9715);
  and g23949 (n14567, n_9716, n14566);
  not g23950 (n_9721, n14565);
  not g23951 (n_9722, n14567);
  and g23952 (n14568, n_9721, n_9722);
  not g23953 (n_9723, n14558);
  not g23954 (n_9724, n14568);
  and g23955 (n14569, n_9723, n_9724);
  not g23956 (n_9725, n14569);
  and g23957 (n14570, \asqrt[58] , n_9725);
  and g23961 (n14574, n_9331, n_9330);
  and g23962 (n14575, \asqrt[16] , n14574);
  not g23963 (n_9726, n14575);
  and g23964 (n14576, n_9329, n_9726);
  not g23965 (n_9727, n14573);
  not g23966 (n_9728, n14576);
  and g23967 (n14577, n_9727, n_9728);
  and g23968 (n14578, n_282, n_9723);
  and g23969 (n14579, n_9724, n14578);
  not g23970 (n_9729, n14577);
  not g23971 (n_9730, n14579);
  and g23972 (n14580, n_9729, n_9730);
  not g23973 (n_9731, n14570);
  not g23974 (n_9732, n14580);
  and g23975 (n14581, n_9731, n_9732);
  not g23976 (n_9733, n14581);
  and g23977 (n14582, \asqrt[59] , n_9733);
  and g23981 (n14586, n_9339, n_9338);
  and g23982 (n14587, \asqrt[16] , n14586);
  not g23983 (n_9734, n14587);
  and g23984 (n14588, n_9337, n_9734);
  not g23985 (n_9735, n14585);
  not g23986 (n_9736, n14588);
  and g23987 (n14589, n_9735, n_9736);
  and g23988 (n14590, n_218, n_9731);
  and g23989 (n14591, n_9732, n14590);
  not g23990 (n_9737, n14589);
  not g23991 (n_9738, n14591);
  and g23992 (n14592, n_9737, n_9738);
  not g23993 (n_9739, n14582);
  not g23994 (n_9740, n14592);
  and g23995 (n14593, n_9739, n_9740);
  not g23996 (n_9741, n14593);
  and g23997 (n14594, \asqrt[60] , n_9741);
  and g24001 (n14598, n_9347, n_9346);
  and g24002 (n14599, \asqrt[16] , n14598);
  not g24003 (n_9742, n14599);
  and g24004 (n14600, n_9345, n_9742);
  not g24005 (n_9743, n14597);
  not g24006 (n_9744, n14600);
  and g24007 (n14601, n_9743, n_9744);
  and g24008 (n14602, n_162, n_9739);
  and g24009 (n14603, n_9740, n14602);
  not g24010 (n_9745, n14601);
  not g24011 (n_9746, n14603);
  and g24012 (n14604, n_9745, n_9746);
  not g24013 (n_9747, n14594);
  not g24014 (n_9748, n14604);
  and g24015 (n14605, n_9747, n_9748);
  not g24016 (n_9749, n14605);
  and g24017 (n14606, \asqrt[61] , n_9749);
  and g24021 (n14610, n_9355, n_9354);
  and g24022 (n14611, \asqrt[16] , n14610);
  not g24023 (n_9750, n14611);
  and g24024 (n14612, n_9353, n_9750);
  not g24025 (n_9751, n14609);
  not g24026 (n_9752, n14612);
  and g24027 (n14613, n_9751, n_9752);
  and g24028 (n14614, n_115, n_9747);
  and g24029 (n14615, n_9748, n14614);
  not g24030 (n_9753, n14613);
  not g24031 (n_9754, n14615);
  and g24032 (n14616, n_9753, n_9754);
  not g24033 (n_9755, n14606);
  not g24034 (n_9756, n14616);
  and g24035 (n14617, n_9755, n_9756);
  not g24036 (n_9757, n14617);
  and g24037 (n14618, \asqrt[62] , n_9757);
  and g24041 (n14622, n_9363, n_9362);
  and g24042 (n14623, \asqrt[16] , n14622);
  not g24043 (n_9758, n14623);
  and g24044 (n14624, n_9361, n_9758);
  not g24045 (n_9759, n14621);
  not g24046 (n_9760, n14624);
  and g24047 (n14625, n_9759, n_9760);
  and g24048 (n14626, n_76, n_9755);
  and g24049 (n14627, n_9756, n14626);
  not g24050 (n_9761, n14625);
  not g24051 (n_9762, n14627);
  and g24052 (n14628, n_9761, n_9762);
  not g24053 (n_9763, n14618);
  not g24054 (n_9764, n14628);
  and g24055 (n14629, n_9763, n_9764);
  and g24059 (n14633, n_9371, n_9370);
  and g24060 (n14634, \asqrt[16] , n14633);
  not g24061 (n_9765, n14634);
  and g24062 (n14635, n_9369, n_9765);
  not g24063 (n_9766, n14632);
  not g24064 (n_9767, n14635);
  and g24065 (n14636, n_9766, n_9767);
  and g24066 (n14637, n_9378, n_9377);
  and g24067 (n14638, \asqrt[16] , n14637);
  not g24070 (n_9769, n14636);
  not g24072 (n_9770, n14629);
  not g24074 (n_9771, n14641);
  and g24075 (n14642, n_21, n_9771);
  and g24076 (n14643, n_9763, n14636);
  and g24077 (n14644, n_9764, n14643);
  and g24078 (n14645, n_9377, \asqrt[16] );
  not g24079 (n_9772, n14645);
  and g24080 (n14646, n14045, n_9772);
  not g24081 (n_9773, n14637);
  and g24082 (n14647, \asqrt[63] , n_9773);
  not g24083 (n_9774, n14646);
  and g24084 (n14648, n_9774, n14647);
  not g24090 (n_9775, n14648);
  not g24091 (n_9776, n14653);
  not g24093 (n_9777, n14644);
  and g24097 (n14657, \a[30] , \asqrt[15] );
  not g24098 (n_9782, \a[28] );
  not g24099 (n_9783, \a[29] );
  and g24100 (n14658, n_9782, n_9783);
  and g24101 (n14659, n_9390, n14658);
  not g24102 (n_9784, n14657);
  not g24103 (n_9785, n14659);
  and g24104 (n14660, n_9784, n_9785);
  not g24105 (n_9786, n14660);
  and g24106 (n14661, \asqrt[16] , n_9786);
  and g24112 (n14667, n_9390, \asqrt[15] );
  not g24113 (n_9787, n14667);
  and g24114 (n14668, \a[31] , n_9787);
  and g24115 (n14669, n14074, \asqrt[15] );
  not g24116 (n_9788, n14668);
  not g24117 (n_9789, n14669);
  and g24118 (n14670, n_9788, n_9789);
  not g24119 (n_9790, n14666);
  and g24120 (n14671, n_9790, n14670);
  not g24121 (n_9791, n14661);
  not g24122 (n_9792, n14671);
  and g24123 (n14672, n_9791, n_9792);
  not g24124 (n_9793, n14672);
  and g24125 (n14673, \asqrt[17] , n_9793);
  not g24126 (n_9794, \asqrt[17] );
  and g24127 (n14674, n_9794, n_9791);
  and g24128 (n14675, n_9792, n14674);
  not g24132 (n_9795, n14642);
  not g24134 (n_9796, n14679);
  and g24135 (n14680, n_9789, n_9796);
  not g24136 (n_9797, n14680);
  and g24137 (n14681, \a[32] , n_9797);
  and g24138 (n14682, n_9006, n_9796);
  and g24139 (n14683, n_9789, n14682);
  not g24140 (n_9798, n14681);
  not g24141 (n_9799, n14683);
  and g24142 (n14684, n_9798, n_9799);
  not g24143 (n_9800, n14675);
  not g24144 (n_9801, n14684);
  and g24145 (n14685, n_9800, n_9801);
  not g24146 (n_9802, n14673);
  not g24147 (n_9803, n14685);
  and g24148 (n14686, n_9802, n_9803);
  not g24149 (n_9804, n14686);
  and g24150 (n14687, \asqrt[18] , n_9804);
  and g24151 (n14688, n_9399, n_9398);
  not g24152 (n_9805, n14086);
  and g24153 (n14689, n_9805, n14688);
  and g24154 (n14690, \asqrt[15] , n14689);
  and g24155 (n14691, \asqrt[15] , n14688);
  not g24156 (n_9806, n14691);
  and g24157 (n14692, n14086, n_9806);
  not g24158 (n_9807, n14690);
  not g24159 (n_9808, n14692);
  and g24160 (n14693, n_9807, n_9808);
  and g24161 (n14694, n_9402, n_9802);
  and g24162 (n14695, n_9803, n14694);
  not g24163 (n_9809, n14693);
  not g24164 (n_9810, n14695);
  and g24165 (n14696, n_9809, n_9810);
  not g24166 (n_9811, n14687);
  not g24167 (n_9812, n14696);
  and g24168 (n14697, n_9811, n_9812);
  not g24169 (n_9813, n14697);
  and g24170 (n14698, \asqrt[19] , n_9813);
  and g24174 (n14702, n_9410, n_9408);
  and g24175 (n14703, \asqrt[15] , n14702);
  not g24176 (n_9814, n14703);
  and g24177 (n14704, n_9409, n_9814);
  not g24178 (n_9815, n14701);
  not g24179 (n_9816, n14704);
  and g24180 (n14705, n_9815, n_9816);
  and g24181 (n14706, n_9018, n_9811);
  and g24182 (n14707, n_9812, n14706);
  not g24183 (n_9817, n14705);
  not g24184 (n_9818, n14707);
  and g24185 (n14708, n_9817, n_9818);
  not g24186 (n_9819, n14698);
  not g24187 (n_9820, n14708);
  and g24188 (n14709, n_9819, n_9820);
  not g24189 (n_9821, n14709);
  and g24190 (n14710, \asqrt[20] , n_9821);
  and g24194 (n14714, n_9419, n_9418);
  and g24195 (n14715, \asqrt[15] , n14714);
  not g24196 (n_9822, n14715);
  and g24197 (n14716, n_9417, n_9822);
  not g24198 (n_9823, n14713);
  not g24199 (n_9824, n14716);
  and g24200 (n14717, n_9823, n_9824);
  and g24201 (n14718, n_8642, n_9819);
  and g24202 (n14719, n_9820, n14718);
  not g24203 (n_9825, n14717);
  not g24204 (n_9826, n14719);
  and g24205 (n14720, n_9825, n_9826);
  not g24206 (n_9827, n14710);
  not g24207 (n_9828, n14720);
  and g24208 (n14721, n_9827, n_9828);
  not g24209 (n_9829, n14721);
  and g24210 (n14722, \asqrt[21] , n_9829);
  and g24214 (n14726, n_9427, n_9426);
  and g24215 (n14727, \asqrt[15] , n14726);
  not g24216 (n_9830, n14727);
  and g24217 (n14728, n_9425, n_9830);
  not g24218 (n_9831, n14725);
  not g24219 (n_9832, n14728);
  and g24220 (n14729, n_9831, n_9832);
  and g24221 (n14730, n_8274, n_9827);
  and g24222 (n14731, n_9828, n14730);
  not g24223 (n_9833, n14729);
  not g24224 (n_9834, n14731);
  and g24225 (n14732, n_9833, n_9834);
  not g24226 (n_9835, n14722);
  not g24227 (n_9836, n14732);
  and g24228 (n14733, n_9835, n_9836);
  not g24229 (n_9837, n14733);
  and g24230 (n14734, \asqrt[22] , n_9837);
  and g24234 (n14738, n_9435, n_9434);
  and g24235 (n14739, \asqrt[15] , n14738);
  not g24236 (n_9838, n14739);
  and g24237 (n14740, n_9433, n_9838);
  not g24238 (n_9839, n14737);
  not g24239 (n_9840, n14740);
  and g24240 (n14741, n_9839, n_9840);
  and g24241 (n14742, n_7914, n_9835);
  and g24242 (n14743, n_9836, n14742);
  not g24243 (n_9841, n14741);
  not g24244 (n_9842, n14743);
  and g24245 (n14744, n_9841, n_9842);
  not g24246 (n_9843, n14734);
  not g24247 (n_9844, n14744);
  and g24248 (n14745, n_9843, n_9844);
  not g24249 (n_9845, n14745);
  and g24250 (n14746, \asqrt[23] , n_9845);
  and g24254 (n14750, n_9443, n_9442);
  and g24255 (n14751, \asqrt[15] , n14750);
  not g24256 (n_9846, n14751);
  and g24257 (n14752, n_9441, n_9846);
  not g24258 (n_9847, n14749);
  not g24259 (n_9848, n14752);
  and g24260 (n14753, n_9847, n_9848);
  and g24261 (n14754, n_7562, n_9843);
  and g24262 (n14755, n_9844, n14754);
  not g24263 (n_9849, n14753);
  not g24264 (n_9850, n14755);
  and g24265 (n14756, n_9849, n_9850);
  not g24266 (n_9851, n14746);
  not g24267 (n_9852, n14756);
  and g24268 (n14757, n_9851, n_9852);
  not g24269 (n_9853, n14757);
  and g24270 (n14758, \asqrt[24] , n_9853);
  and g24274 (n14762, n_9451, n_9450);
  and g24275 (n14763, \asqrt[15] , n14762);
  not g24276 (n_9854, n14763);
  and g24277 (n14764, n_9449, n_9854);
  not g24278 (n_9855, n14761);
  not g24279 (n_9856, n14764);
  and g24280 (n14765, n_9855, n_9856);
  and g24281 (n14766, n_7218, n_9851);
  and g24282 (n14767, n_9852, n14766);
  not g24283 (n_9857, n14765);
  not g24284 (n_9858, n14767);
  and g24285 (n14768, n_9857, n_9858);
  not g24286 (n_9859, n14758);
  not g24287 (n_9860, n14768);
  and g24288 (n14769, n_9859, n_9860);
  not g24289 (n_9861, n14769);
  and g24290 (n14770, \asqrt[25] , n_9861);
  and g24294 (n14774, n_9459, n_9458);
  and g24295 (n14775, \asqrt[15] , n14774);
  not g24296 (n_9862, n14775);
  and g24297 (n14776, n_9457, n_9862);
  not g24298 (n_9863, n14773);
  not g24299 (n_9864, n14776);
  and g24300 (n14777, n_9863, n_9864);
  and g24301 (n14778, n_6882, n_9859);
  and g24302 (n14779, n_9860, n14778);
  not g24303 (n_9865, n14777);
  not g24304 (n_9866, n14779);
  and g24305 (n14780, n_9865, n_9866);
  not g24306 (n_9867, n14770);
  not g24307 (n_9868, n14780);
  and g24308 (n14781, n_9867, n_9868);
  not g24309 (n_9869, n14781);
  and g24310 (n14782, \asqrt[26] , n_9869);
  and g24314 (n14786, n_9467, n_9466);
  and g24315 (n14787, \asqrt[15] , n14786);
  not g24316 (n_9870, n14787);
  and g24317 (n14788, n_9465, n_9870);
  not g24318 (n_9871, n14785);
  not g24319 (n_9872, n14788);
  and g24320 (n14789, n_9871, n_9872);
  and g24321 (n14790, n_6554, n_9867);
  and g24322 (n14791, n_9868, n14790);
  not g24323 (n_9873, n14789);
  not g24324 (n_9874, n14791);
  and g24325 (n14792, n_9873, n_9874);
  not g24326 (n_9875, n14782);
  not g24327 (n_9876, n14792);
  and g24328 (n14793, n_9875, n_9876);
  not g24329 (n_9877, n14793);
  and g24330 (n14794, \asqrt[27] , n_9877);
  and g24334 (n14798, n_9475, n_9474);
  and g24335 (n14799, \asqrt[15] , n14798);
  not g24336 (n_9878, n14799);
  and g24337 (n14800, n_9473, n_9878);
  not g24338 (n_9879, n14797);
  not g24339 (n_9880, n14800);
  and g24340 (n14801, n_9879, n_9880);
  and g24341 (n14802, n_6234, n_9875);
  and g24342 (n14803, n_9876, n14802);
  not g24343 (n_9881, n14801);
  not g24344 (n_9882, n14803);
  and g24345 (n14804, n_9881, n_9882);
  not g24346 (n_9883, n14794);
  not g24347 (n_9884, n14804);
  and g24348 (n14805, n_9883, n_9884);
  not g24349 (n_9885, n14805);
  and g24350 (n14806, \asqrt[28] , n_9885);
  and g24354 (n14810, n_9483, n_9482);
  and g24355 (n14811, \asqrt[15] , n14810);
  not g24356 (n_9886, n14811);
  and g24357 (n14812, n_9481, n_9886);
  not g24358 (n_9887, n14809);
  not g24359 (n_9888, n14812);
  and g24360 (n14813, n_9887, n_9888);
  and g24361 (n14814, n_5922, n_9883);
  and g24362 (n14815, n_9884, n14814);
  not g24363 (n_9889, n14813);
  not g24364 (n_9890, n14815);
  and g24365 (n14816, n_9889, n_9890);
  not g24366 (n_9891, n14806);
  not g24367 (n_9892, n14816);
  and g24368 (n14817, n_9891, n_9892);
  not g24369 (n_9893, n14817);
  and g24370 (n14818, \asqrt[29] , n_9893);
  and g24374 (n14822, n_9491, n_9490);
  and g24375 (n14823, \asqrt[15] , n14822);
  not g24376 (n_9894, n14823);
  and g24377 (n14824, n_9489, n_9894);
  not g24378 (n_9895, n14821);
  not g24379 (n_9896, n14824);
  and g24380 (n14825, n_9895, n_9896);
  and g24381 (n14826, n_5618, n_9891);
  and g24382 (n14827, n_9892, n14826);
  not g24383 (n_9897, n14825);
  not g24384 (n_9898, n14827);
  and g24385 (n14828, n_9897, n_9898);
  not g24386 (n_9899, n14818);
  not g24387 (n_9900, n14828);
  and g24388 (n14829, n_9899, n_9900);
  not g24389 (n_9901, n14829);
  and g24390 (n14830, \asqrt[30] , n_9901);
  and g24394 (n14834, n_9499, n_9498);
  and g24395 (n14835, \asqrt[15] , n14834);
  not g24396 (n_9902, n14835);
  and g24397 (n14836, n_9497, n_9902);
  not g24398 (n_9903, n14833);
  not g24399 (n_9904, n14836);
  and g24400 (n14837, n_9903, n_9904);
  and g24401 (n14838, n_5322, n_9899);
  and g24402 (n14839, n_9900, n14838);
  not g24403 (n_9905, n14837);
  not g24404 (n_9906, n14839);
  and g24405 (n14840, n_9905, n_9906);
  not g24406 (n_9907, n14830);
  not g24407 (n_9908, n14840);
  and g24408 (n14841, n_9907, n_9908);
  not g24409 (n_9909, n14841);
  and g24410 (n14842, \asqrt[31] , n_9909);
  and g24414 (n14846, n_9507, n_9506);
  and g24415 (n14847, \asqrt[15] , n14846);
  not g24416 (n_9910, n14847);
  and g24417 (n14848, n_9505, n_9910);
  not g24418 (n_9911, n14845);
  not g24419 (n_9912, n14848);
  and g24420 (n14849, n_9911, n_9912);
  and g24421 (n14850, n_5034, n_9907);
  and g24422 (n14851, n_9908, n14850);
  not g24423 (n_9913, n14849);
  not g24424 (n_9914, n14851);
  and g24425 (n14852, n_9913, n_9914);
  not g24426 (n_9915, n14842);
  not g24427 (n_9916, n14852);
  and g24428 (n14853, n_9915, n_9916);
  not g24429 (n_9917, n14853);
  and g24430 (n14854, \asqrt[32] , n_9917);
  and g24434 (n14858, n_9515, n_9514);
  and g24435 (n14859, \asqrt[15] , n14858);
  not g24436 (n_9918, n14859);
  and g24437 (n14860, n_9513, n_9918);
  not g24438 (n_9919, n14857);
  not g24439 (n_9920, n14860);
  and g24440 (n14861, n_9919, n_9920);
  and g24441 (n14862, n_4754, n_9915);
  and g24442 (n14863, n_9916, n14862);
  not g24443 (n_9921, n14861);
  not g24444 (n_9922, n14863);
  and g24445 (n14864, n_9921, n_9922);
  not g24446 (n_9923, n14854);
  not g24447 (n_9924, n14864);
  and g24448 (n14865, n_9923, n_9924);
  not g24449 (n_9925, n14865);
  and g24450 (n14866, \asqrt[33] , n_9925);
  and g24454 (n14870, n_9523, n_9522);
  and g24455 (n14871, \asqrt[15] , n14870);
  not g24456 (n_9926, n14871);
  and g24457 (n14872, n_9521, n_9926);
  not g24458 (n_9927, n14869);
  not g24459 (n_9928, n14872);
  and g24460 (n14873, n_9927, n_9928);
  and g24461 (n14874, n_4482, n_9923);
  and g24462 (n14875, n_9924, n14874);
  not g24463 (n_9929, n14873);
  not g24464 (n_9930, n14875);
  and g24465 (n14876, n_9929, n_9930);
  not g24466 (n_9931, n14866);
  not g24467 (n_9932, n14876);
  and g24468 (n14877, n_9931, n_9932);
  not g24469 (n_9933, n14877);
  and g24470 (n14878, \asqrt[34] , n_9933);
  and g24474 (n14882, n_9531, n_9530);
  and g24475 (n14883, \asqrt[15] , n14882);
  not g24476 (n_9934, n14883);
  and g24477 (n14884, n_9529, n_9934);
  not g24478 (n_9935, n14881);
  not g24479 (n_9936, n14884);
  and g24480 (n14885, n_9935, n_9936);
  and g24481 (n14886, n_4218, n_9931);
  and g24482 (n14887, n_9932, n14886);
  not g24483 (n_9937, n14885);
  not g24484 (n_9938, n14887);
  and g24485 (n14888, n_9937, n_9938);
  not g24486 (n_9939, n14878);
  not g24487 (n_9940, n14888);
  and g24488 (n14889, n_9939, n_9940);
  not g24489 (n_9941, n14889);
  and g24490 (n14890, \asqrt[35] , n_9941);
  and g24494 (n14894, n_9539, n_9538);
  and g24495 (n14895, \asqrt[15] , n14894);
  not g24496 (n_9942, n14895);
  and g24497 (n14896, n_9537, n_9942);
  not g24498 (n_9943, n14893);
  not g24499 (n_9944, n14896);
  and g24500 (n14897, n_9943, n_9944);
  and g24501 (n14898, n_3962, n_9939);
  and g24502 (n14899, n_9940, n14898);
  not g24503 (n_9945, n14897);
  not g24504 (n_9946, n14899);
  and g24505 (n14900, n_9945, n_9946);
  not g24506 (n_9947, n14890);
  not g24507 (n_9948, n14900);
  and g24508 (n14901, n_9947, n_9948);
  not g24509 (n_9949, n14901);
  and g24510 (n14902, \asqrt[36] , n_9949);
  and g24514 (n14906, n_9547, n_9546);
  and g24515 (n14907, \asqrt[15] , n14906);
  not g24516 (n_9950, n14907);
  and g24517 (n14908, n_9545, n_9950);
  not g24518 (n_9951, n14905);
  not g24519 (n_9952, n14908);
  and g24520 (n14909, n_9951, n_9952);
  and g24521 (n14910, n_3714, n_9947);
  and g24522 (n14911, n_9948, n14910);
  not g24523 (n_9953, n14909);
  not g24524 (n_9954, n14911);
  and g24525 (n14912, n_9953, n_9954);
  not g24526 (n_9955, n14902);
  not g24527 (n_9956, n14912);
  and g24528 (n14913, n_9955, n_9956);
  not g24529 (n_9957, n14913);
  and g24530 (n14914, \asqrt[37] , n_9957);
  and g24534 (n14918, n_9555, n_9554);
  and g24535 (n14919, \asqrt[15] , n14918);
  not g24536 (n_9958, n14919);
  and g24537 (n14920, n_9553, n_9958);
  not g24538 (n_9959, n14917);
  not g24539 (n_9960, n14920);
  and g24540 (n14921, n_9959, n_9960);
  and g24541 (n14922, n_3474, n_9955);
  and g24542 (n14923, n_9956, n14922);
  not g24543 (n_9961, n14921);
  not g24544 (n_9962, n14923);
  and g24545 (n14924, n_9961, n_9962);
  not g24546 (n_9963, n14914);
  not g24547 (n_9964, n14924);
  and g24548 (n14925, n_9963, n_9964);
  not g24549 (n_9965, n14925);
  and g24550 (n14926, \asqrt[38] , n_9965);
  and g24554 (n14930, n_9563, n_9562);
  and g24555 (n14931, \asqrt[15] , n14930);
  not g24556 (n_9966, n14931);
  and g24557 (n14932, n_9561, n_9966);
  not g24558 (n_9967, n14929);
  not g24559 (n_9968, n14932);
  and g24560 (n14933, n_9967, n_9968);
  and g24561 (n14934, n_3242, n_9963);
  and g24562 (n14935, n_9964, n14934);
  not g24563 (n_9969, n14933);
  not g24564 (n_9970, n14935);
  and g24565 (n14936, n_9969, n_9970);
  not g24566 (n_9971, n14926);
  not g24567 (n_9972, n14936);
  and g24568 (n14937, n_9971, n_9972);
  not g24569 (n_9973, n14937);
  and g24570 (n14938, \asqrt[39] , n_9973);
  and g24574 (n14942, n_9571, n_9570);
  and g24575 (n14943, \asqrt[15] , n14942);
  not g24576 (n_9974, n14943);
  and g24577 (n14944, n_9569, n_9974);
  not g24578 (n_9975, n14941);
  not g24579 (n_9976, n14944);
  and g24580 (n14945, n_9975, n_9976);
  and g24581 (n14946, n_3018, n_9971);
  and g24582 (n14947, n_9972, n14946);
  not g24583 (n_9977, n14945);
  not g24584 (n_9978, n14947);
  and g24585 (n14948, n_9977, n_9978);
  not g24586 (n_9979, n14938);
  not g24587 (n_9980, n14948);
  and g24588 (n14949, n_9979, n_9980);
  not g24589 (n_9981, n14949);
  and g24590 (n14950, \asqrt[40] , n_9981);
  and g24594 (n14954, n_9579, n_9578);
  and g24595 (n14955, \asqrt[15] , n14954);
  not g24596 (n_9982, n14955);
  and g24597 (n14956, n_9577, n_9982);
  not g24598 (n_9983, n14953);
  not g24599 (n_9984, n14956);
  and g24600 (n14957, n_9983, n_9984);
  and g24601 (n14958, n_2802, n_9979);
  and g24602 (n14959, n_9980, n14958);
  not g24603 (n_9985, n14957);
  not g24604 (n_9986, n14959);
  and g24605 (n14960, n_9985, n_9986);
  not g24606 (n_9987, n14950);
  not g24607 (n_9988, n14960);
  and g24608 (n14961, n_9987, n_9988);
  not g24609 (n_9989, n14961);
  and g24610 (n14962, \asqrt[41] , n_9989);
  and g24614 (n14966, n_9587, n_9586);
  and g24615 (n14967, \asqrt[15] , n14966);
  not g24616 (n_9990, n14967);
  and g24617 (n14968, n_9585, n_9990);
  not g24618 (n_9991, n14965);
  not g24619 (n_9992, n14968);
  and g24620 (n14969, n_9991, n_9992);
  and g24621 (n14970, n_2594, n_9987);
  and g24622 (n14971, n_9988, n14970);
  not g24623 (n_9993, n14969);
  not g24624 (n_9994, n14971);
  and g24625 (n14972, n_9993, n_9994);
  not g24626 (n_9995, n14962);
  not g24627 (n_9996, n14972);
  and g24628 (n14973, n_9995, n_9996);
  not g24629 (n_9997, n14973);
  and g24630 (n14974, \asqrt[42] , n_9997);
  and g24634 (n14978, n_9595, n_9594);
  and g24635 (n14979, \asqrt[15] , n14978);
  not g24636 (n_9998, n14979);
  and g24637 (n14980, n_9593, n_9998);
  not g24638 (n_9999, n14977);
  not g24639 (n_10000, n14980);
  and g24640 (n14981, n_9999, n_10000);
  and g24641 (n14982, n_2394, n_9995);
  and g24642 (n14983, n_9996, n14982);
  not g24643 (n_10001, n14981);
  not g24644 (n_10002, n14983);
  and g24645 (n14984, n_10001, n_10002);
  not g24646 (n_10003, n14974);
  not g24647 (n_10004, n14984);
  and g24648 (n14985, n_10003, n_10004);
  not g24649 (n_10005, n14985);
  and g24650 (n14986, \asqrt[43] , n_10005);
  and g24654 (n14990, n_9603, n_9602);
  and g24655 (n14991, \asqrt[15] , n14990);
  not g24656 (n_10006, n14991);
  and g24657 (n14992, n_9601, n_10006);
  not g24658 (n_10007, n14989);
  not g24659 (n_10008, n14992);
  and g24660 (n14993, n_10007, n_10008);
  and g24661 (n14994, n_2202, n_10003);
  and g24662 (n14995, n_10004, n14994);
  not g24663 (n_10009, n14993);
  not g24664 (n_10010, n14995);
  and g24665 (n14996, n_10009, n_10010);
  not g24666 (n_10011, n14986);
  not g24667 (n_10012, n14996);
  and g24668 (n14997, n_10011, n_10012);
  not g24669 (n_10013, n14997);
  and g24670 (n14998, \asqrt[44] , n_10013);
  and g24674 (n15002, n_9611, n_9610);
  and g24675 (n15003, \asqrt[15] , n15002);
  not g24676 (n_10014, n15003);
  and g24677 (n15004, n_9609, n_10014);
  not g24678 (n_10015, n15001);
  not g24679 (n_10016, n15004);
  and g24680 (n15005, n_10015, n_10016);
  and g24681 (n15006, n_2018, n_10011);
  and g24682 (n15007, n_10012, n15006);
  not g24683 (n_10017, n15005);
  not g24684 (n_10018, n15007);
  and g24685 (n15008, n_10017, n_10018);
  not g24686 (n_10019, n14998);
  not g24687 (n_10020, n15008);
  and g24688 (n15009, n_10019, n_10020);
  not g24689 (n_10021, n15009);
  and g24690 (n15010, \asqrt[45] , n_10021);
  and g24694 (n15014, n_9619, n_9618);
  and g24695 (n15015, \asqrt[15] , n15014);
  not g24696 (n_10022, n15015);
  and g24697 (n15016, n_9617, n_10022);
  not g24698 (n_10023, n15013);
  not g24699 (n_10024, n15016);
  and g24700 (n15017, n_10023, n_10024);
  and g24701 (n15018, n_1842, n_10019);
  and g24702 (n15019, n_10020, n15018);
  not g24703 (n_10025, n15017);
  not g24704 (n_10026, n15019);
  and g24705 (n15020, n_10025, n_10026);
  not g24706 (n_10027, n15010);
  not g24707 (n_10028, n15020);
  and g24708 (n15021, n_10027, n_10028);
  not g24709 (n_10029, n15021);
  and g24710 (n15022, \asqrt[46] , n_10029);
  and g24714 (n15026, n_9627, n_9626);
  and g24715 (n15027, \asqrt[15] , n15026);
  not g24716 (n_10030, n15027);
  and g24717 (n15028, n_9625, n_10030);
  not g24718 (n_10031, n15025);
  not g24719 (n_10032, n15028);
  and g24720 (n15029, n_10031, n_10032);
  and g24721 (n15030, n_1674, n_10027);
  and g24722 (n15031, n_10028, n15030);
  not g24723 (n_10033, n15029);
  not g24724 (n_10034, n15031);
  and g24725 (n15032, n_10033, n_10034);
  not g24726 (n_10035, n15022);
  not g24727 (n_10036, n15032);
  and g24728 (n15033, n_10035, n_10036);
  not g24729 (n_10037, n15033);
  and g24730 (n15034, \asqrt[47] , n_10037);
  and g24734 (n15038, n_9635, n_9634);
  and g24735 (n15039, \asqrt[15] , n15038);
  not g24736 (n_10038, n15039);
  and g24737 (n15040, n_9633, n_10038);
  not g24738 (n_10039, n15037);
  not g24739 (n_10040, n15040);
  and g24740 (n15041, n_10039, n_10040);
  and g24741 (n15042, n_1514, n_10035);
  and g24742 (n15043, n_10036, n15042);
  not g24743 (n_10041, n15041);
  not g24744 (n_10042, n15043);
  and g24745 (n15044, n_10041, n_10042);
  not g24746 (n_10043, n15034);
  not g24747 (n_10044, n15044);
  and g24748 (n15045, n_10043, n_10044);
  not g24749 (n_10045, n15045);
  and g24750 (n15046, \asqrt[48] , n_10045);
  and g24754 (n15050, n_9643, n_9642);
  and g24755 (n15051, \asqrt[15] , n15050);
  not g24756 (n_10046, n15051);
  and g24757 (n15052, n_9641, n_10046);
  not g24758 (n_10047, n15049);
  not g24759 (n_10048, n15052);
  and g24760 (n15053, n_10047, n_10048);
  and g24761 (n15054, n_1362, n_10043);
  and g24762 (n15055, n_10044, n15054);
  not g24763 (n_10049, n15053);
  not g24764 (n_10050, n15055);
  and g24765 (n15056, n_10049, n_10050);
  not g24766 (n_10051, n15046);
  not g24767 (n_10052, n15056);
  and g24768 (n15057, n_10051, n_10052);
  not g24769 (n_10053, n15057);
  and g24770 (n15058, \asqrt[49] , n_10053);
  and g24774 (n15062, n_9651, n_9650);
  and g24775 (n15063, \asqrt[15] , n15062);
  not g24776 (n_10054, n15063);
  and g24777 (n15064, n_9649, n_10054);
  not g24778 (n_10055, n15061);
  not g24779 (n_10056, n15064);
  and g24780 (n15065, n_10055, n_10056);
  and g24781 (n15066, n_1218, n_10051);
  and g24782 (n15067, n_10052, n15066);
  not g24783 (n_10057, n15065);
  not g24784 (n_10058, n15067);
  and g24785 (n15068, n_10057, n_10058);
  not g24786 (n_10059, n15058);
  not g24787 (n_10060, n15068);
  and g24788 (n15069, n_10059, n_10060);
  not g24789 (n_10061, n15069);
  and g24790 (n15070, \asqrt[50] , n_10061);
  and g24791 (n15071, n_1082, n_10059);
  and g24792 (n15072, n_10060, n15071);
  and g24796 (n15076, n_9659, n_9657);
  and g24797 (n15077, \asqrt[15] , n15076);
  not g24798 (n_10062, n15077);
  and g24799 (n15078, n_9658, n_10062);
  not g24800 (n_10063, n15075);
  not g24801 (n_10064, n15078);
  and g24802 (n15079, n_10063, n_10064);
  not g24803 (n_10065, n15072);
  not g24804 (n_10066, n15079);
  and g24805 (n15080, n_10065, n_10066);
  not g24806 (n_10067, n15070);
  not g24807 (n_10068, n15080);
  and g24808 (n15081, n_10067, n_10068);
  not g24809 (n_10069, n15081);
  and g24810 (n15082, \asqrt[51] , n_10069);
  and g24814 (n15086, n_9667, n_9666);
  and g24815 (n15087, \asqrt[15] , n15086);
  not g24816 (n_10070, n15087);
  and g24817 (n15088, n_9665, n_10070);
  not g24818 (n_10071, n15085);
  not g24819 (n_10072, n15088);
  and g24820 (n15089, n_10071, n_10072);
  and g24821 (n15090, n_954, n_10067);
  and g24822 (n15091, n_10068, n15090);
  not g24823 (n_10073, n15089);
  not g24824 (n_10074, n15091);
  and g24825 (n15092, n_10073, n_10074);
  not g24826 (n_10075, n15082);
  not g24827 (n_10076, n15092);
  and g24828 (n15093, n_10075, n_10076);
  not g24829 (n_10077, n15093);
  and g24830 (n15094, \asqrt[52] , n_10077);
  and g24834 (n15098, n_9675, n_9674);
  and g24835 (n15099, \asqrt[15] , n15098);
  not g24836 (n_10078, n15099);
  and g24837 (n15100, n_9673, n_10078);
  not g24838 (n_10079, n15097);
  not g24839 (n_10080, n15100);
  and g24840 (n15101, n_10079, n_10080);
  and g24841 (n15102, n_834, n_10075);
  and g24842 (n15103, n_10076, n15102);
  not g24843 (n_10081, n15101);
  not g24844 (n_10082, n15103);
  and g24845 (n15104, n_10081, n_10082);
  not g24846 (n_10083, n15094);
  not g24847 (n_10084, n15104);
  and g24848 (n15105, n_10083, n_10084);
  not g24849 (n_10085, n15105);
  and g24850 (n15106, \asqrt[53] , n_10085);
  and g24854 (n15110, n_9683, n_9682);
  and g24855 (n15111, \asqrt[15] , n15110);
  not g24856 (n_10086, n15111);
  and g24857 (n15112, n_9681, n_10086);
  not g24858 (n_10087, n15109);
  not g24859 (n_10088, n15112);
  and g24860 (n15113, n_10087, n_10088);
  and g24861 (n15114, n_722, n_10083);
  and g24862 (n15115, n_10084, n15114);
  not g24863 (n_10089, n15113);
  not g24864 (n_10090, n15115);
  and g24865 (n15116, n_10089, n_10090);
  not g24866 (n_10091, n15106);
  not g24867 (n_10092, n15116);
  and g24868 (n15117, n_10091, n_10092);
  not g24869 (n_10093, n15117);
  and g24870 (n15118, \asqrt[54] , n_10093);
  and g24874 (n15122, n_9691, n_9690);
  and g24875 (n15123, \asqrt[15] , n15122);
  not g24876 (n_10094, n15123);
  and g24877 (n15124, n_9689, n_10094);
  not g24878 (n_10095, n15121);
  not g24879 (n_10096, n15124);
  and g24880 (n15125, n_10095, n_10096);
  and g24881 (n15126, n_618, n_10091);
  and g24882 (n15127, n_10092, n15126);
  not g24883 (n_10097, n15125);
  not g24884 (n_10098, n15127);
  and g24885 (n15128, n_10097, n_10098);
  not g24886 (n_10099, n15118);
  not g24887 (n_10100, n15128);
  and g24888 (n15129, n_10099, n_10100);
  not g24889 (n_10101, n15129);
  and g24890 (n15130, \asqrt[55] , n_10101);
  and g24894 (n15134, n_9699, n_9698);
  and g24895 (n15135, \asqrt[15] , n15134);
  not g24896 (n_10102, n15135);
  and g24897 (n15136, n_9697, n_10102);
  not g24898 (n_10103, n15133);
  not g24899 (n_10104, n15136);
  and g24900 (n15137, n_10103, n_10104);
  and g24901 (n15138, n_522, n_10099);
  and g24902 (n15139, n_10100, n15138);
  not g24903 (n_10105, n15137);
  not g24904 (n_10106, n15139);
  and g24905 (n15140, n_10105, n_10106);
  not g24906 (n_10107, n15130);
  not g24907 (n_10108, n15140);
  and g24908 (n15141, n_10107, n_10108);
  not g24909 (n_10109, n15141);
  and g24910 (n15142, \asqrt[56] , n_10109);
  and g24914 (n15146, n_9707, n_9706);
  and g24915 (n15147, \asqrt[15] , n15146);
  not g24916 (n_10110, n15147);
  and g24917 (n15148, n_9705, n_10110);
  not g24918 (n_10111, n15145);
  not g24919 (n_10112, n15148);
  and g24920 (n15149, n_10111, n_10112);
  and g24921 (n15150, n_434, n_10107);
  and g24922 (n15151, n_10108, n15150);
  not g24923 (n_10113, n15149);
  not g24924 (n_10114, n15151);
  and g24925 (n15152, n_10113, n_10114);
  not g24926 (n_10115, n15142);
  not g24927 (n_10116, n15152);
  and g24928 (n15153, n_10115, n_10116);
  not g24929 (n_10117, n15153);
  and g24930 (n15154, \asqrt[57] , n_10117);
  and g24934 (n15158, n_9715, n_9714);
  and g24935 (n15159, \asqrt[15] , n15158);
  not g24936 (n_10118, n15159);
  and g24937 (n15160, n_9713, n_10118);
  not g24938 (n_10119, n15157);
  not g24939 (n_10120, n15160);
  and g24940 (n15161, n_10119, n_10120);
  and g24941 (n15162, n_354, n_10115);
  and g24942 (n15163, n_10116, n15162);
  not g24943 (n_10121, n15161);
  not g24944 (n_10122, n15163);
  and g24945 (n15164, n_10121, n_10122);
  not g24946 (n_10123, n15154);
  not g24947 (n_10124, n15164);
  and g24948 (n15165, n_10123, n_10124);
  not g24949 (n_10125, n15165);
  and g24950 (n15166, \asqrt[58] , n_10125);
  and g24954 (n15170, n_9723, n_9722);
  and g24955 (n15171, \asqrt[15] , n15170);
  not g24956 (n_10126, n15171);
  and g24957 (n15172, n_9721, n_10126);
  not g24958 (n_10127, n15169);
  not g24959 (n_10128, n15172);
  and g24960 (n15173, n_10127, n_10128);
  and g24961 (n15174, n_282, n_10123);
  and g24962 (n15175, n_10124, n15174);
  not g24963 (n_10129, n15173);
  not g24964 (n_10130, n15175);
  and g24965 (n15176, n_10129, n_10130);
  not g24966 (n_10131, n15166);
  not g24967 (n_10132, n15176);
  and g24968 (n15177, n_10131, n_10132);
  not g24969 (n_10133, n15177);
  and g24970 (n15178, \asqrt[59] , n_10133);
  and g24974 (n15182, n_9731, n_9730);
  and g24975 (n15183, \asqrt[15] , n15182);
  not g24976 (n_10134, n15183);
  and g24977 (n15184, n_9729, n_10134);
  not g24978 (n_10135, n15181);
  not g24979 (n_10136, n15184);
  and g24980 (n15185, n_10135, n_10136);
  and g24981 (n15186, n_218, n_10131);
  and g24982 (n15187, n_10132, n15186);
  not g24983 (n_10137, n15185);
  not g24984 (n_10138, n15187);
  and g24985 (n15188, n_10137, n_10138);
  not g24986 (n_10139, n15178);
  not g24987 (n_10140, n15188);
  and g24988 (n15189, n_10139, n_10140);
  not g24989 (n_10141, n15189);
  and g24990 (n15190, \asqrt[60] , n_10141);
  and g24994 (n15194, n_9739, n_9738);
  and g24995 (n15195, \asqrt[15] , n15194);
  not g24996 (n_10142, n15195);
  and g24997 (n15196, n_9737, n_10142);
  not g24998 (n_10143, n15193);
  not g24999 (n_10144, n15196);
  and g25000 (n15197, n_10143, n_10144);
  and g25001 (n15198, n_162, n_10139);
  and g25002 (n15199, n_10140, n15198);
  not g25003 (n_10145, n15197);
  not g25004 (n_10146, n15199);
  and g25005 (n15200, n_10145, n_10146);
  not g25006 (n_10147, n15190);
  not g25007 (n_10148, n15200);
  and g25008 (n15201, n_10147, n_10148);
  not g25009 (n_10149, n15201);
  and g25010 (n15202, \asqrt[61] , n_10149);
  and g25014 (n15206, n_9747, n_9746);
  and g25015 (n15207, \asqrt[15] , n15206);
  not g25016 (n_10150, n15207);
  and g25017 (n15208, n_9745, n_10150);
  not g25018 (n_10151, n15205);
  not g25019 (n_10152, n15208);
  and g25020 (n15209, n_10151, n_10152);
  and g25021 (n15210, n_115, n_10147);
  and g25022 (n15211, n_10148, n15210);
  not g25023 (n_10153, n15209);
  not g25024 (n_10154, n15211);
  and g25025 (n15212, n_10153, n_10154);
  not g25026 (n_10155, n15202);
  not g25027 (n_10156, n15212);
  and g25028 (n15213, n_10155, n_10156);
  not g25029 (n_10157, n15213);
  and g25030 (n15214, \asqrt[62] , n_10157);
  and g25034 (n15218, n_9755, n_9754);
  and g25035 (n15219, \asqrt[15] , n15218);
  not g25036 (n_10158, n15219);
  and g25037 (n15220, n_9753, n_10158);
  not g25038 (n_10159, n15217);
  not g25039 (n_10160, n15220);
  and g25040 (n15221, n_10159, n_10160);
  and g25041 (n15222, n_76, n_10155);
  and g25042 (n15223, n_10156, n15222);
  not g25043 (n_10161, n15221);
  not g25044 (n_10162, n15223);
  and g25045 (n15224, n_10161, n_10162);
  not g25046 (n_10163, n15214);
  not g25047 (n_10164, n15224);
  and g25048 (n15225, n_10163, n_10164);
  and g25052 (n15229, n_9763, n_9762);
  and g25053 (n15230, \asqrt[15] , n15229);
  not g25054 (n_10165, n15230);
  and g25055 (n15231, n_9761, n_10165);
  not g25056 (n_10166, n15228);
  not g25057 (n_10167, n15231);
  and g25058 (n15232, n_10166, n_10167);
  and g25059 (n15233, n_9770, n_9769);
  and g25060 (n15234, \asqrt[15] , n15233);
  not g25063 (n_10169, n15232);
  not g25065 (n_10170, n15225);
  not g25067 (n_10171, n15237);
  and g25068 (n15238, n_21, n_10171);
  and g25069 (n15239, n_10163, n15232);
  and g25070 (n15240, n_10164, n15239);
  and g25071 (n15241, n_9769, \asqrt[15] );
  not g25072 (n_10172, n15241);
  and g25073 (n15242, n14629, n_10172);
  not g25074 (n_10173, n15233);
  and g25075 (n15243, \asqrt[63] , n_10173);
  not g25076 (n_10174, n15242);
  and g25077 (n15244, n_10174, n15243);
  not g25083 (n_10175, n15244);
  not g25084 (n_10176, n15249);
  not g25086 (n_10177, n15240);
  and g25090 (n15253, \a[28] , \asqrt[14] );
  not g25091 (n_10182, \a[26] );
  not g25092 (n_10183, \a[27] );
  and g25093 (n15254, n_10182, n_10183);
  and g25094 (n15255, n_9782, n15254);
  not g25095 (n_10184, n15253);
  not g25096 (n_10185, n15255);
  and g25097 (n15256, n_10184, n_10185);
  not g25098 (n_10186, n15256);
  and g25099 (n15257, \asqrt[15] , n_10186);
  and g25105 (n15263, n_9782, \asqrt[14] );
  not g25106 (n_10187, n15263);
  and g25107 (n15264, \a[29] , n_10187);
  and g25108 (n15265, n14658, \asqrt[14] );
  not g25109 (n_10188, n15264);
  not g25110 (n_10189, n15265);
  and g25111 (n15266, n_10188, n_10189);
  not g25112 (n_10190, n15262);
  and g25113 (n15267, n_10190, n15266);
  not g25114 (n_10191, n15257);
  not g25115 (n_10192, n15267);
  and g25116 (n15268, n_10191, n_10192);
  not g25117 (n_10193, n15268);
  and g25118 (n15269, \asqrt[16] , n_10193);
  not g25119 (n_10194, \asqrt[16] );
  and g25120 (n15270, n_10194, n_10191);
  and g25121 (n15271, n_10192, n15270);
  not g25125 (n_10195, n15238);
  not g25127 (n_10196, n15275);
  and g25128 (n15276, n_10189, n_10196);
  not g25129 (n_10197, n15276);
  and g25130 (n15277, \a[30] , n_10197);
  and g25131 (n15278, n_9390, n_10196);
  and g25132 (n15279, n_10189, n15278);
  not g25133 (n_10198, n15277);
  not g25134 (n_10199, n15279);
  and g25135 (n15280, n_10198, n_10199);
  not g25136 (n_10200, n15271);
  not g25137 (n_10201, n15280);
  and g25138 (n15281, n_10200, n_10201);
  not g25139 (n_10202, n15269);
  not g25140 (n_10203, n15281);
  and g25141 (n15282, n_10202, n_10203);
  not g25142 (n_10204, n15282);
  and g25143 (n15283, \asqrt[17] , n_10204);
  and g25144 (n15284, n_9791, n_9790);
  not g25145 (n_10205, n14670);
  and g25146 (n15285, n_10205, n15284);
  and g25147 (n15286, \asqrt[14] , n15285);
  and g25148 (n15287, \asqrt[14] , n15284);
  not g25149 (n_10206, n15287);
  and g25150 (n15288, n14670, n_10206);
  not g25151 (n_10207, n15286);
  not g25152 (n_10208, n15288);
  and g25153 (n15289, n_10207, n_10208);
  and g25154 (n15290, n_9794, n_10202);
  and g25155 (n15291, n_10203, n15290);
  not g25156 (n_10209, n15289);
  not g25157 (n_10210, n15291);
  and g25158 (n15292, n_10209, n_10210);
  not g25159 (n_10211, n15283);
  not g25160 (n_10212, n15292);
  and g25161 (n15293, n_10211, n_10212);
  not g25162 (n_10213, n15293);
  and g25163 (n15294, \asqrt[18] , n_10213);
  and g25167 (n15298, n_9802, n_9800);
  and g25168 (n15299, \asqrt[14] , n15298);
  not g25169 (n_10214, n15299);
  and g25170 (n15300, n_9801, n_10214);
  not g25171 (n_10215, n15297);
  not g25172 (n_10216, n15300);
  and g25173 (n15301, n_10215, n_10216);
  and g25174 (n15302, n_9402, n_10211);
  and g25175 (n15303, n_10212, n15302);
  not g25176 (n_10217, n15301);
  not g25177 (n_10218, n15303);
  and g25178 (n15304, n_10217, n_10218);
  not g25179 (n_10219, n15294);
  not g25180 (n_10220, n15304);
  and g25181 (n15305, n_10219, n_10220);
  not g25182 (n_10221, n15305);
  and g25183 (n15306, \asqrt[19] , n_10221);
  and g25187 (n15310, n_9811, n_9810);
  and g25188 (n15311, \asqrt[14] , n15310);
  not g25189 (n_10222, n15311);
  and g25190 (n15312, n_9809, n_10222);
  not g25191 (n_10223, n15309);
  not g25192 (n_10224, n15312);
  and g25193 (n15313, n_10223, n_10224);
  and g25194 (n15314, n_9018, n_10219);
  and g25195 (n15315, n_10220, n15314);
  not g25196 (n_10225, n15313);
  not g25197 (n_10226, n15315);
  and g25198 (n15316, n_10225, n_10226);
  not g25199 (n_10227, n15306);
  not g25200 (n_10228, n15316);
  and g25201 (n15317, n_10227, n_10228);
  not g25202 (n_10229, n15317);
  and g25203 (n15318, \asqrt[20] , n_10229);
  and g25207 (n15322, n_9819, n_9818);
  and g25208 (n15323, \asqrt[14] , n15322);
  not g25209 (n_10230, n15323);
  and g25210 (n15324, n_9817, n_10230);
  not g25211 (n_10231, n15321);
  not g25212 (n_10232, n15324);
  and g25213 (n15325, n_10231, n_10232);
  and g25214 (n15326, n_8642, n_10227);
  and g25215 (n15327, n_10228, n15326);
  not g25216 (n_10233, n15325);
  not g25217 (n_10234, n15327);
  and g25218 (n15328, n_10233, n_10234);
  not g25219 (n_10235, n15318);
  not g25220 (n_10236, n15328);
  and g25221 (n15329, n_10235, n_10236);
  not g25222 (n_10237, n15329);
  and g25223 (n15330, \asqrt[21] , n_10237);
  and g25227 (n15334, n_9827, n_9826);
  and g25228 (n15335, \asqrt[14] , n15334);
  not g25229 (n_10238, n15335);
  and g25230 (n15336, n_9825, n_10238);
  not g25231 (n_10239, n15333);
  not g25232 (n_10240, n15336);
  and g25233 (n15337, n_10239, n_10240);
  and g25234 (n15338, n_8274, n_10235);
  and g25235 (n15339, n_10236, n15338);
  not g25236 (n_10241, n15337);
  not g25237 (n_10242, n15339);
  and g25238 (n15340, n_10241, n_10242);
  not g25239 (n_10243, n15330);
  not g25240 (n_10244, n15340);
  and g25241 (n15341, n_10243, n_10244);
  not g25242 (n_10245, n15341);
  and g25243 (n15342, \asqrt[22] , n_10245);
  and g25247 (n15346, n_9835, n_9834);
  and g25248 (n15347, \asqrt[14] , n15346);
  not g25249 (n_10246, n15347);
  and g25250 (n15348, n_9833, n_10246);
  not g25251 (n_10247, n15345);
  not g25252 (n_10248, n15348);
  and g25253 (n15349, n_10247, n_10248);
  and g25254 (n15350, n_7914, n_10243);
  and g25255 (n15351, n_10244, n15350);
  not g25256 (n_10249, n15349);
  not g25257 (n_10250, n15351);
  and g25258 (n15352, n_10249, n_10250);
  not g25259 (n_10251, n15342);
  not g25260 (n_10252, n15352);
  and g25261 (n15353, n_10251, n_10252);
  not g25262 (n_10253, n15353);
  and g25263 (n15354, \asqrt[23] , n_10253);
  and g25267 (n15358, n_9843, n_9842);
  and g25268 (n15359, \asqrt[14] , n15358);
  not g25269 (n_10254, n15359);
  and g25270 (n15360, n_9841, n_10254);
  not g25271 (n_10255, n15357);
  not g25272 (n_10256, n15360);
  and g25273 (n15361, n_10255, n_10256);
  and g25274 (n15362, n_7562, n_10251);
  and g25275 (n15363, n_10252, n15362);
  not g25276 (n_10257, n15361);
  not g25277 (n_10258, n15363);
  and g25278 (n15364, n_10257, n_10258);
  not g25279 (n_10259, n15354);
  not g25280 (n_10260, n15364);
  and g25281 (n15365, n_10259, n_10260);
  not g25282 (n_10261, n15365);
  and g25283 (n15366, \asqrt[24] , n_10261);
  and g25287 (n15370, n_9851, n_9850);
  and g25288 (n15371, \asqrt[14] , n15370);
  not g25289 (n_10262, n15371);
  and g25290 (n15372, n_9849, n_10262);
  not g25291 (n_10263, n15369);
  not g25292 (n_10264, n15372);
  and g25293 (n15373, n_10263, n_10264);
  and g25294 (n15374, n_7218, n_10259);
  and g25295 (n15375, n_10260, n15374);
  not g25296 (n_10265, n15373);
  not g25297 (n_10266, n15375);
  and g25298 (n15376, n_10265, n_10266);
  not g25299 (n_10267, n15366);
  not g25300 (n_10268, n15376);
  and g25301 (n15377, n_10267, n_10268);
  not g25302 (n_10269, n15377);
  and g25303 (n15378, \asqrt[25] , n_10269);
  and g25307 (n15382, n_9859, n_9858);
  and g25308 (n15383, \asqrt[14] , n15382);
  not g25309 (n_10270, n15383);
  and g25310 (n15384, n_9857, n_10270);
  not g25311 (n_10271, n15381);
  not g25312 (n_10272, n15384);
  and g25313 (n15385, n_10271, n_10272);
  and g25314 (n15386, n_6882, n_10267);
  and g25315 (n15387, n_10268, n15386);
  not g25316 (n_10273, n15385);
  not g25317 (n_10274, n15387);
  and g25318 (n15388, n_10273, n_10274);
  not g25319 (n_10275, n15378);
  not g25320 (n_10276, n15388);
  and g25321 (n15389, n_10275, n_10276);
  not g25322 (n_10277, n15389);
  and g25323 (n15390, \asqrt[26] , n_10277);
  and g25327 (n15394, n_9867, n_9866);
  and g25328 (n15395, \asqrt[14] , n15394);
  not g25329 (n_10278, n15395);
  and g25330 (n15396, n_9865, n_10278);
  not g25331 (n_10279, n15393);
  not g25332 (n_10280, n15396);
  and g25333 (n15397, n_10279, n_10280);
  and g25334 (n15398, n_6554, n_10275);
  and g25335 (n15399, n_10276, n15398);
  not g25336 (n_10281, n15397);
  not g25337 (n_10282, n15399);
  and g25338 (n15400, n_10281, n_10282);
  not g25339 (n_10283, n15390);
  not g25340 (n_10284, n15400);
  and g25341 (n15401, n_10283, n_10284);
  not g25342 (n_10285, n15401);
  and g25343 (n15402, \asqrt[27] , n_10285);
  and g25347 (n15406, n_9875, n_9874);
  and g25348 (n15407, \asqrt[14] , n15406);
  not g25349 (n_10286, n15407);
  and g25350 (n15408, n_9873, n_10286);
  not g25351 (n_10287, n15405);
  not g25352 (n_10288, n15408);
  and g25353 (n15409, n_10287, n_10288);
  and g25354 (n15410, n_6234, n_10283);
  and g25355 (n15411, n_10284, n15410);
  not g25356 (n_10289, n15409);
  not g25357 (n_10290, n15411);
  and g25358 (n15412, n_10289, n_10290);
  not g25359 (n_10291, n15402);
  not g25360 (n_10292, n15412);
  and g25361 (n15413, n_10291, n_10292);
  not g25362 (n_10293, n15413);
  and g25363 (n15414, \asqrt[28] , n_10293);
  and g25367 (n15418, n_9883, n_9882);
  and g25368 (n15419, \asqrt[14] , n15418);
  not g25369 (n_10294, n15419);
  and g25370 (n15420, n_9881, n_10294);
  not g25371 (n_10295, n15417);
  not g25372 (n_10296, n15420);
  and g25373 (n15421, n_10295, n_10296);
  and g25374 (n15422, n_5922, n_10291);
  and g25375 (n15423, n_10292, n15422);
  not g25376 (n_10297, n15421);
  not g25377 (n_10298, n15423);
  and g25378 (n15424, n_10297, n_10298);
  not g25379 (n_10299, n15414);
  not g25380 (n_10300, n15424);
  and g25381 (n15425, n_10299, n_10300);
  not g25382 (n_10301, n15425);
  and g25383 (n15426, \asqrt[29] , n_10301);
  and g25387 (n15430, n_9891, n_9890);
  and g25388 (n15431, \asqrt[14] , n15430);
  not g25389 (n_10302, n15431);
  and g25390 (n15432, n_9889, n_10302);
  not g25391 (n_10303, n15429);
  not g25392 (n_10304, n15432);
  and g25393 (n15433, n_10303, n_10304);
  and g25394 (n15434, n_5618, n_10299);
  and g25395 (n15435, n_10300, n15434);
  not g25396 (n_10305, n15433);
  not g25397 (n_10306, n15435);
  and g25398 (n15436, n_10305, n_10306);
  not g25399 (n_10307, n15426);
  not g25400 (n_10308, n15436);
  and g25401 (n15437, n_10307, n_10308);
  not g25402 (n_10309, n15437);
  and g25403 (n15438, \asqrt[30] , n_10309);
  and g25407 (n15442, n_9899, n_9898);
  and g25408 (n15443, \asqrt[14] , n15442);
  not g25409 (n_10310, n15443);
  and g25410 (n15444, n_9897, n_10310);
  not g25411 (n_10311, n15441);
  not g25412 (n_10312, n15444);
  and g25413 (n15445, n_10311, n_10312);
  and g25414 (n15446, n_5322, n_10307);
  and g25415 (n15447, n_10308, n15446);
  not g25416 (n_10313, n15445);
  not g25417 (n_10314, n15447);
  and g25418 (n15448, n_10313, n_10314);
  not g25419 (n_10315, n15438);
  not g25420 (n_10316, n15448);
  and g25421 (n15449, n_10315, n_10316);
  not g25422 (n_10317, n15449);
  and g25423 (n15450, \asqrt[31] , n_10317);
  and g25427 (n15454, n_9907, n_9906);
  and g25428 (n15455, \asqrt[14] , n15454);
  not g25429 (n_10318, n15455);
  and g25430 (n15456, n_9905, n_10318);
  not g25431 (n_10319, n15453);
  not g25432 (n_10320, n15456);
  and g25433 (n15457, n_10319, n_10320);
  and g25434 (n15458, n_5034, n_10315);
  and g25435 (n15459, n_10316, n15458);
  not g25436 (n_10321, n15457);
  not g25437 (n_10322, n15459);
  and g25438 (n15460, n_10321, n_10322);
  not g25439 (n_10323, n15450);
  not g25440 (n_10324, n15460);
  and g25441 (n15461, n_10323, n_10324);
  not g25442 (n_10325, n15461);
  and g25443 (n15462, \asqrt[32] , n_10325);
  and g25447 (n15466, n_9915, n_9914);
  and g25448 (n15467, \asqrt[14] , n15466);
  not g25449 (n_10326, n15467);
  and g25450 (n15468, n_9913, n_10326);
  not g25451 (n_10327, n15465);
  not g25452 (n_10328, n15468);
  and g25453 (n15469, n_10327, n_10328);
  and g25454 (n15470, n_4754, n_10323);
  and g25455 (n15471, n_10324, n15470);
  not g25456 (n_10329, n15469);
  not g25457 (n_10330, n15471);
  and g25458 (n15472, n_10329, n_10330);
  not g25459 (n_10331, n15462);
  not g25460 (n_10332, n15472);
  and g25461 (n15473, n_10331, n_10332);
  not g25462 (n_10333, n15473);
  and g25463 (n15474, \asqrt[33] , n_10333);
  and g25467 (n15478, n_9923, n_9922);
  and g25468 (n15479, \asqrt[14] , n15478);
  not g25469 (n_10334, n15479);
  and g25470 (n15480, n_9921, n_10334);
  not g25471 (n_10335, n15477);
  not g25472 (n_10336, n15480);
  and g25473 (n15481, n_10335, n_10336);
  and g25474 (n15482, n_4482, n_10331);
  and g25475 (n15483, n_10332, n15482);
  not g25476 (n_10337, n15481);
  not g25477 (n_10338, n15483);
  and g25478 (n15484, n_10337, n_10338);
  not g25479 (n_10339, n15474);
  not g25480 (n_10340, n15484);
  and g25481 (n15485, n_10339, n_10340);
  not g25482 (n_10341, n15485);
  and g25483 (n15486, \asqrt[34] , n_10341);
  and g25487 (n15490, n_9931, n_9930);
  and g25488 (n15491, \asqrt[14] , n15490);
  not g25489 (n_10342, n15491);
  and g25490 (n15492, n_9929, n_10342);
  not g25491 (n_10343, n15489);
  not g25492 (n_10344, n15492);
  and g25493 (n15493, n_10343, n_10344);
  and g25494 (n15494, n_4218, n_10339);
  and g25495 (n15495, n_10340, n15494);
  not g25496 (n_10345, n15493);
  not g25497 (n_10346, n15495);
  and g25498 (n15496, n_10345, n_10346);
  not g25499 (n_10347, n15486);
  not g25500 (n_10348, n15496);
  and g25501 (n15497, n_10347, n_10348);
  not g25502 (n_10349, n15497);
  and g25503 (n15498, \asqrt[35] , n_10349);
  and g25507 (n15502, n_9939, n_9938);
  and g25508 (n15503, \asqrt[14] , n15502);
  not g25509 (n_10350, n15503);
  and g25510 (n15504, n_9937, n_10350);
  not g25511 (n_10351, n15501);
  not g25512 (n_10352, n15504);
  and g25513 (n15505, n_10351, n_10352);
  and g25514 (n15506, n_3962, n_10347);
  and g25515 (n15507, n_10348, n15506);
  not g25516 (n_10353, n15505);
  not g25517 (n_10354, n15507);
  and g25518 (n15508, n_10353, n_10354);
  not g25519 (n_10355, n15498);
  not g25520 (n_10356, n15508);
  and g25521 (n15509, n_10355, n_10356);
  not g25522 (n_10357, n15509);
  and g25523 (n15510, \asqrt[36] , n_10357);
  and g25527 (n15514, n_9947, n_9946);
  and g25528 (n15515, \asqrt[14] , n15514);
  not g25529 (n_10358, n15515);
  and g25530 (n15516, n_9945, n_10358);
  not g25531 (n_10359, n15513);
  not g25532 (n_10360, n15516);
  and g25533 (n15517, n_10359, n_10360);
  and g25534 (n15518, n_3714, n_10355);
  and g25535 (n15519, n_10356, n15518);
  not g25536 (n_10361, n15517);
  not g25537 (n_10362, n15519);
  and g25538 (n15520, n_10361, n_10362);
  not g25539 (n_10363, n15510);
  not g25540 (n_10364, n15520);
  and g25541 (n15521, n_10363, n_10364);
  not g25542 (n_10365, n15521);
  and g25543 (n15522, \asqrt[37] , n_10365);
  and g25547 (n15526, n_9955, n_9954);
  and g25548 (n15527, \asqrt[14] , n15526);
  not g25549 (n_10366, n15527);
  and g25550 (n15528, n_9953, n_10366);
  not g25551 (n_10367, n15525);
  not g25552 (n_10368, n15528);
  and g25553 (n15529, n_10367, n_10368);
  and g25554 (n15530, n_3474, n_10363);
  and g25555 (n15531, n_10364, n15530);
  not g25556 (n_10369, n15529);
  not g25557 (n_10370, n15531);
  and g25558 (n15532, n_10369, n_10370);
  not g25559 (n_10371, n15522);
  not g25560 (n_10372, n15532);
  and g25561 (n15533, n_10371, n_10372);
  not g25562 (n_10373, n15533);
  and g25563 (n15534, \asqrt[38] , n_10373);
  and g25567 (n15538, n_9963, n_9962);
  and g25568 (n15539, \asqrt[14] , n15538);
  not g25569 (n_10374, n15539);
  and g25570 (n15540, n_9961, n_10374);
  not g25571 (n_10375, n15537);
  not g25572 (n_10376, n15540);
  and g25573 (n15541, n_10375, n_10376);
  and g25574 (n15542, n_3242, n_10371);
  and g25575 (n15543, n_10372, n15542);
  not g25576 (n_10377, n15541);
  not g25577 (n_10378, n15543);
  and g25578 (n15544, n_10377, n_10378);
  not g25579 (n_10379, n15534);
  not g25580 (n_10380, n15544);
  and g25581 (n15545, n_10379, n_10380);
  not g25582 (n_10381, n15545);
  and g25583 (n15546, \asqrt[39] , n_10381);
  and g25587 (n15550, n_9971, n_9970);
  and g25588 (n15551, \asqrt[14] , n15550);
  not g25589 (n_10382, n15551);
  and g25590 (n15552, n_9969, n_10382);
  not g25591 (n_10383, n15549);
  not g25592 (n_10384, n15552);
  and g25593 (n15553, n_10383, n_10384);
  and g25594 (n15554, n_3018, n_10379);
  and g25595 (n15555, n_10380, n15554);
  not g25596 (n_10385, n15553);
  not g25597 (n_10386, n15555);
  and g25598 (n15556, n_10385, n_10386);
  not g25599 (n_10387, n15546);
  not g25600 (n_10388, n15556);
  and g25601 (n15557, n_10387, n_10388);
  not g25602 (n_10389, n15557);
  and g25603 (n15558, \asqrt[40] , n_10389);
  and g25607 (n15562, n_9979, n_9978);
  and g25608 (n15563, \asqrt[14] , n15562);
  not g25609 (n_10390, n15563);
  and g25610 (n15564, n_9977, n_10390);
  not g25611 (n_10391, n15561);
  not g25612 (n_10392, n15564);
  and g25613 (n15565, n_10391, n_10392);
  and g25614 (n15566, n_2802, n_10387);
  and g25615 (n15567, n_10388, n15566);
  not g25616 (n_10393, n15565);
  not g25617 (n_10394, n15567);
  and g25618 (n15568, n_10393, n_10394);
  not g25619 (n_10395, n15558);
  not g25620 (n_10396, n15568);
  and g25621 (n15569, n_10395, n_10396);
  not g25622 (n_10397, n15569);
  and g25623 (n15570, \asqrt[41] , n_10397);
  and g25627 (n15574, n_9987, n_9986);
  and g25628 (n15575, \asqrt[14] , n15574);
  not g25629 (n_10398, n15575);
  and g25630 (n15576, n_9985, n_10398);
  not g25631 (n_10399, n15573);
  not g25632 (n_10400, n15576);
  and g25633 (n15577, n_10399, n_10400);
  and g25634 (n15578, n_2594, n_10395);
  and g25635 (n15579, n_10396, n15578);
  not g25636 (n_10401, n15577);
  not g25637 (n_10402, n15579);
  and g25638 (n15580, n_10401, n_10402);
  not g25639 (n_10403, n15570);
  not g25640 (n_10404, n15580);
  and g25641 (n15581, n_10403, n_10404);
  not g25642 (n_10405, n15581);
  and g25643 (n15582, \asqrt[42] , n_10405);
  and g25647 (n15586, n_9995, n_9994);
  and g25648 (n15587, \asqrt[14] , n15586);
  not g25649 (n_10406, n15587);
  and g25650 (n15588, n_9993, n_10406);
  not g25651 (n_10407, n15585);
  not g25652 (n_10408, n15588);
  and g25653 (n15589, n_10407, n_10408);
  and g25654 (n15590, n_2394, n_10403);
  and g25655 (n15591, n_10404, n15590);
  not g25656 (n_10409, n15589);
  not g25657 (n_10410, n15591);
  and g25658 (n15592, n_10409, n_10410);
  not g25659 (n_10411, n15582);
  not g25660 (n_10412, n15592);
  and g25661 (n15593, n_10411, n_10412);
  not g25662 (n_10413, n15593);
  and g25663 (n15594, \asqrt[43] , n_10413);
  and g25667 (n15598, n_10003, n_10002);
  and g25668 (n15599, \asqrt[14] , n15598);
  not g25669 (n_10414, n15599);
  and g25670 (n15600, n_10001, n_10414);
  not g25671 (n_10415, n15597);
  not g25672 (n_10416, n15600);
  and g25673 (n15601, n_10415, n_10416);
  and g25674 (n15602, n_2202, n_10411);
  and g25675 (n15603, n_10412, n15602);
  not g25676 (n_10417, n15601);
  not g25677 (n_10418, n15603);
  and g25678 (n15604, n_10417, n_10418);
  not g25679 (n_10419, n15594);
  not g25680 (n_10420, n15604);
  and g25681 (n15605, n_10419, n_10420);
  not g25682 (n_10421, n15605);
  and g25683 (n15606, \asqrt[44] , n_10421);
  and g25687 (n15610, n_10011, n_10010);
  and g25688 (n15611, \asqrt[14] , n15610);
  not g25689 (n_10422, n15611);
  and g25690 (n15612, n_10009, n_10422);
  not g25691 (n_10423, n15609);
  not g25692 (n_10424, n15612);
  and g25693 (n15613, n_10423, n_10424);
  and g25694 (n15614, n_2018, n_10419);
  and g25695 (n15615, n_10420, n15614);
  not g25696 (n_10425, n15613);
  not g25697 (n_10426, n15615);
  and g25698 (n15616, n_10425, n_10426);
  not g25699 (n_10427, n15606);
  not g25700 (n_10428, n15616);
  and g25701 (n15617, n_10427, n_10428);
  not g25702 (n_10429, n15617);
  and g25703 (n15618, \asqrt[45] , n_10429);
  and g25707 (n15622, n_10019, n_10018);
  and g25708 (n15623, \asqrt[14] , n15622);
  not g25709 (n_10430, n15623);
  and g25710 (n15624, n_10017, n_10430);
  not g25711 (n_10431, n15621);
  not g25712 (n_10432, n15624);
  and g25713 (n15625, n_10431, n_10432);
  and g25714 (n15626, n_1842, n_10427);
  and g25715 (n15627, n_10428, n15626);
  not g25716 (n_10433, n15625);
  not g25717 (n_10434, n15627);
  and g25718 (n15628, n_10433, n_10434);
  not g25719 (n_10435, n15618);
  not g25720 (n_10436, n15628);
  and g25721 (n15629, n_10435, n_10436);
  not g25722 (n_10437, n15629);
  and g25723 (n15630, \asqrt[46] , n_10437);
  and g25727 (n15634, n_10027, n_10026);
  and g25728 (n15635, \asqrt[14] , n15634);
  not g25729 (n_10438, n15635);
  and g25730 (n15636, n_10025, n_10438);
  not g25731 (n_10439, n15633);
  not g25732 (n_10440, n15636);
  and g25733 (n15637, n_10439, n_10440);
  and g25734 (n15638, n_1674, n_10435);
  and g25735 (n15639, n_10436, n15638);
  not g25736 (n_10441, n15637);
  not g25737 (n_10442, n15639);
  and g25738 (n15640, n_10441, n_10442);
  not g25739 (n_10443, n15630);
  not g25740 (n_10444, n15640);
  and g25741 (n15641, n_10443, n_10444);
  not g25742 (n_10445, n15641);
  and g25743 (n15642, \asqrt[47] , n_10445);
  and g25747 (n15646, n_10035, n_10034);
  and g25748 (n15647, \asqrt[14] , n15646);
  not g25749 (n_10446, n15647);
  and g25750 (n15648, n_10033, n_10446);
  not g25751 (n_10447, n15645);
  not g25752 (n_10448, n15648);
  and g25753 (n15649, n_10447, n_10448);
  and g25754 (n15650, n_1514, n_10443);
  and g25755 (n15651, n_10444, n15650);
  not g25756 (n_10449, n15649);
  not g25757 (n_10450, n15651);
  and g25758 (n15652, n_10449, n_10450);
  not g25759 (n_10451, n15642);
  not g25760 (n_10452, n15652);
  and g25761 (n15653, n_10451, n_10452);
  not g25762 (n_10453, n15653);
  and g25763 (n15654, \asqrt[48] , n_10453);
  and g25767 (n15658, n_10043, n_10042);
  and g25768 (n15659, \asqrt[14] , n15658);
  not g25769 (n_10454, n15659);
  and g25770 (n15660, n_10041, n_10454);
  not g25771 (n_10455, n15657);
  not g25772 (n_10456, n15660);
  and g25773 (n15661, n_10455, n_10456);
  and g25774 (n15662, n_1362, n_10451);
  and g25775 (n15663, n_10452, n15662);
  not g25776 (n_10457, n15661);
  not g25777 (n_10458, n15663);
  and g25778 (n15664, n_10457, n_10458);
  not g25779 (n_10459, n15654);
  not g25780 (n_10460, n15664);
  and g25781 (n15665, n_10459, n_10460);
  not g25782 (n_10461, n15665);
  and g25783 (n15666, \asqrt[49] , n_10461);
  and g25787 (n15670, n_10051, n_10050);
  and g25788 (n15671, \asqrt[14] , n15670);
  not g25789 (n_10462, n15671);
  and g25790 (n15672, n_10049, n_10462);
  not g25791 (n_10463, n15669);
  not g25792 (n_10464, n15672);
  and g25793 (n15673, n_10463, n_10464);
  and g25794 (n15674, n_1218, n_10459);
  and g25795 (n15675, n_10460, n15674);
  not g25796 (n_10465, n15673);
  not g25797 (n_10466, n15675);
  and g25798 (n15676, n_10465, n_10466);
  not g25799 (n_10467, n15666);
  not g25800 (n_10468, n15676);
  and g25801 (n15677, n_10467, n_10468);
  not g25802 (n_10469, n15677);
  and g25803 (n15678, \asqrt[50] , n_10469);
  and g25807 (n15682, n_10059, n_10058);
  and g25808 (n15683, \asqrt[14] , n15682);
  not g25809 (n_10470, n15683);
  and g25810 (n15684, n_10057, n_10470);
  not g25811 (n_10471, n15681);
  not g25812 (n_10472, n15684);
  and g25813 (n15685, n_10471, n_10472);
  and g25814 (n15686, n_1082, n_10467);
  and g25815 (n15687, n_10468, n15686);
  not g25816 (n_10473, n15685);
  not g25817 (n_10474, n15687);
  and g25818 (n15688, n_10473, n_10474);
  not g25819 (n_10475, n15678);
  not g25820 (n_10476, n15688);
  and g25821 (n15689, n_10475, n_10476);
  not g25822 (n_10477, n15689);
  and g25823 (n15690, \asqrt[51] , n_10477);
  and g25824 (n15691, n_954, n_10475);
  and g25825 (n15692, n_10476, n15691);
  and g25829 (n15696, n_10067, n_10065);
  and g25830 (n15697, \asqrt[14] , n15696);
  not g25831 (n_10478, n15697);
  and g25832 (n15698, n_10066, n_10478);
  not g25833 (n_10479, n15695);
  not g25834 (n_10480, n15698);
  and g25835 (n15699, n_10479, n_10480);
  not g25836 (n_10481, n15692);
  not g25837 (n_10482, n15699);
  and g25838 (n15700, n_10481, n_10482);
  not g25839 (n_10483, n15690);
  not g25840 (n_10484, n15700);
  and g25841 (n15701, n_10483, n_10484);
  not g25842 (n_10485, n15701);
  and g25843 (n15702, \asqrt[52] , n_10485);
  and g25847 (n15706, n_10075, n_10074);
  and g25848 (n15707, \asqrt[14] , n15706);
  not g25849 (n_10486, n15707);
  and g25850 (n15708, n_10073, n_10486);
  not g25851 (n_10487, n15705);
  not g25852 (n_10488, n15708);
  and g25853 (n15709, n_10487, n_10488);
  and g25854 (n15710, n_834, n_10483);
  and g25855 (n15711, n_10484, n15710);
  not g25856 (n_10489, n15709);
  not g25857 (n_10490, n15711);
  and g25858 (n15712, n_10489, n_10490);
  not g25859 (n_10491, n15702);
  not g25860 (n_10492, n15712);
  and g25861 (n15713, n_10491, n_10492);
  not g25862 (n_10493, n15713);
  and g25863 (n15714, \asqrt[53] , n_10493);
  and g25867 (n15718, n_10083, n_10082);
  and g25868 (n15719, \asqrt[14] , n15718);
  not g25869 (n_10494, n15719);
  and g25870 (n15720, n_10081, n_10494);
  not g25871 (n_10495, n15717);
  not g25872 (n_10496, n15720);
  and g25873 (n15721, n_10495, n_10496);
  and g25874 (n15722, n_722, n_10491);
  and g25875 (n15723, n_10492, n15722);
  not g25876 (n_10497, n15721);
  not g25877 (n_10498, n15723);
  and g25878 (n15724, n_10497, n_10498);
  not g25879 (n_10499, n15714);
  not g25880 (n_10500, n15724);
  and g25881 (n15725, n_10499, n_10500);
  not g25882 (n_10501, n15725);
  and g25883 (n15726, \asqrt[54] , n_10501);
  and g25887 (n15730, n_10091, n_10090);
  and g25888 (n15731, \asqrt[14] , n15730);
  not g25889 (n_10502, n15731);
  and g25890 (n15732, n_10089, n_10502);
  not g25891 (n_10503, n15729);
  not g25892 (n_10504, n15732);
  and g25893 (n15733, n_10503, n_10504);
  and g25894 (n15734, n_618, n_10499);
  and g25895 (n15735, n_10500, n15734);
  not g25896 (n_10505, n15733);
  not g25897 (n_10506, n15735);
  and g25898 (n15736, n_10505, n_10506);
  not g25899 (n_10507, n15726);
  not g25900 (n_10508, n15736);
  and g25901 (n15737, n_10507, n_10508);
  not g25902 (n_10509, n15737);
  and g25903 (n15738, \asqrt[55] , n_10509);
  and g25907 (n15742, n_10099, n_10098);
  and g25908 (n15743, \asqrt[14] , n15742);
  not g25909 (n_10510, n15743);
  and g25910 (n15744, n_10097, n_10510);
  not g25911 (n_10511, n15741);
  not g25912 (n_10512, n15744);
  and g25913 (n15745, n_10511, n_10512);
  and g25914 (n15746, n_522, n_10507);
  and g25915 (n15747, n_10508, n15746);
  not g25916 (n_10513, n15745);
  not g25917 (n_10514, n15747);
  and g25918 (n15748, n_10513, n_10514);
  not g25919 (n_10515, n15738);
  not g25920 (n_10516, n15748);
  and g25921 (n15749, n_10515, n_10516);
  not g25922 (n_10517, n15749);
  and g25923 (n15750, \asqrt[56] , n_10517);
  and g25927 (n15754, n_10107, n_10106);
  and g25928 (n15755, \asqrt[14] , n15754);
  not g25929 (n_10518, n15755);
  and g25930 (n15756, n_10105, n_10518);
  not g25931 (n_10519, n15753);
  not g25932 (n_10520, n15756);
  and g25933 (n15757, n_10519, n_10520);
  and g25934 (n15758, n_434, n_10515);
  and g25935 (n15759, n_10516, n15758);
  not g25936 (n_10521, n15757);
  not g25937 (n_10522, n15759);
  and g25938 (n15760, n_10521, n_10522);
  not g25939 (n_10523, n15750);
  not g25940 (n_10524, n15760);
  and g25941 (n15761, n_10523, n_10524);
  not g25942 (n_10525, n15761);
  and g25943 (n15762, \asqrt[57] , n_10525);
  and g25947 (n15766, n_10115, n_10114);
  and g25948 (n15767, \asqrt[14] , n15766);
  not g25949 (n_10526, n15767);
  and g25950 (n15768, n_10113, n_10526);
  not g25951 (n_10527, n15765);
  not g25952 (n_10528, n15768);
  and g25953 (n15769, n_10527, n_10528);
  and g25954 (n15770, n_354, n_10523);
  and g25955 (n15771, n_10524, n15770);
  not g25956 (n_10529, n15769);
  not g25957 (n_10530, n15771);
  and g25958 (n15772, n_10529, n_10530);
  not g25959 (n_10531, n15762);
  not g25960 (n_10532, n15772);
  and g25961 (n15773, n_10531, n_10532);
  not g25962 (n_10533, n15773);
  and g25963 (n15774, \asqrt[58] , n_10533);
  and g25967 (n15778, n_10123, n_10122);
  and g25968 (n15779, \asqrt[14] , n15778);
  not g25969 (n_10534, n15779);
  and g25970 (n15780, n_10121, n_10534);
  not g25971 (n_10535, n15777);
  not g25972 (n_10536, n15780);
  and g25973 (n15781, n_10535, n_10536);
  and g25974 (n15782, n_282, n_10531);
  and g25975 (n15783, n_10532, n15782);
  not g25976 (n_10537, n15781);
  not g25977 (n_10538, n15783);
  and g25978 (n15784, n_10537, n_10538);
  not g25979 (n_10539, n15774);
  not g25980 (n_10540, n15784);
  and g25981 (n15785, n_10539, n_10540);
  not g25982 (n_10541, n15785);
  and g25983 (n15786, \asqrt[59] , n_10541);
  and g25987 (n15790, n_10131, n_10130);
  and g25988 (n15791, \asqrt[14] , n15790);
  not g25989 (n_10542, n15791);
  and g25990 (n15792, n_10129, n_10542);
  not g25991 (n_10543, n15789);
  not g25992 (n_10544, n15792);
  and g25993 (n15793, n_10543, n_10544);
  and g25994 (n15794, n_218, n_10539);
  and g25995 (n15795, n_10540, n15794);
  not g25996 (n_10545, n15793);
  not g25997 (n_10546, n15795);
  and g25998 (n15796, n_10545, n_10546);
  not g25999 (n_10547, n15786);
  not g26000 (n_10548, n15796);
  and g26001 (n15797, n_10547, n_10548);
  not g26002 (n_10549, n15797);
  and g26003 (n15798, \asqrt[60] , n_10549);
  and g26007 (n15802, n_10139, n_10138);
  and g26008 (n15803, \asqrt[14] , n15802);
  not g26009 (n_10550, n15803);
  and g26010 (n15804, n_10137, n_10550);
  not g26011 (n_10551, n15801);
  not g26012 (n_10552, n15804);
  and g26013 (n15805, n_10551, n_10552);
  and g26014 (n15806, n_162, n_10547);
  and g26015 (n15807, n_10548, n15806);
  not g26016 (n_10553, n15805);
  not g26017 (n_10554, n15807);
  and g26018 (n15808, n_10553, n_10554);
  not g26019 (n_10555, n15798);
  not g26020 (n_10556, n15808);
  and g26021 (n15809, n_10555, n_10556);
  not g26022 (n_10557, n15809);
  and g26023 (n15810, \asqrt[61] , n_10557);
  and g26027 (n15814, n_10147, n_10146);
  and g26028 (n15815, \asqrt[14] , n15814);
  not g26029 (n_10558, n15815);
  and g26030 (n15816, n_10145, n_10558);
  not g26031 (n_10559, n15813);
  not g26032 (n_10560, n15816);
  and g26033 (n15817, n_10559, n_10560);
  and g26034 (n15818, n_115, n_10555);
  and g26035 (n15819, n_10556, n15818);
  not g26036 (n_10561, n15817);
  not g26037 (n_10562, n15819);
  and g26038 (n15820, n_10561, n_10562);
  not g26039 (n_10563, n15810);
  not g26040 (n_10564, n15820);
  and g26041 (n15821, n_10563, n_10564);
  not g26042 (n_10565, n15821);
  and g26043 (n15822, \asqrt[62] , n_10565);
  and g26047 (n15826, n_10155, n_10154);
  and g26048 (n15827, \asqrt[14] , n15826);
  not g26049 (n_10566, n15827);
  and g26050 (n15828, n_10153, n_10566);
  not g26051 (n_10567, n15825);
  not g26052 (n_10568, n15828);
  and g26053 (n15829, n_10567, n_10568);
  and g26054 (n15830, n_76, n_10563);
  and g26055 (n15831, n_10564, n15830);
  not g26056 (n_10569, n15829);
  not g26057 (n_10570, n15831);
  and g26058 (n15832, n_10569, n_10570);
  not g26059 (n_10571, n15822);
  not g26060 (n_10572, n15832);
  and g26061 (n15833, n_10571, n_10572);
  and g26065 (n15837, n_10163, n_10162);
  and g26066 (n15838, \asqrt[14] , n15837);
  not g26067 (n_10573, n15838);
  and g26068 (n15839, n_10161, n_10573);
  not g26069 (n_10574, n15836);
  not g26070 (n_10575, n15839);
  and g26071 (n15840, n_10574, n_10575);
  and g26072 (n15841, n_10170, n_10169);
  and g26073 (n15842, \asqrt[14] , n15841);
  not g26076 (n_10577, n15840);
  not g26078 (n_10578, n15833);
  not g26080 (n_10579, n15845);
  and g26081 (n15846, n_21, n_10579);
  and g26082 (n15847, n_10571, n15840);
  and g26083 (n15848, n_10572, n15847);
  and g26084 (n15849, n_10169, \asqrt[14] );
  not g26085 (n_10580, n15849);
  and g26086 (n15850, n15225, n_10580);
  not g26087 (n_10581, n15841);
  and g26088 (n15851, \asqrt[63] , n_10581);
  not g26089 (n_10582, n15850);
  and g26090 (n15852, n_10582, n15851);
  not g26096 (n_10583, n15852);
  not g26097 (n_10584, n15857);
  not g26099 (n_10585, n15848);
  and g26103 (n15861, \a[26] , \asqrt[13] );
  not g26104 (n_10590, \a[24] );
  not g26105 (n_10591, \a[25] );
  and g26106 (n15862, n_10590, n_10591);
  and g26107 (n15863, n_10182, n15862);
  not g26108 (n_10592, n15861);
  not g26109 (n_10593, n15863);
  and g26110 (n15864, n_10592, n_10593);
  not g26111 (n_10594, n15864);
  and g26112 (n15865, \asqrt[14] , n_10594);
  and g26118 (n15871, n_10182, \asqrt[13] );
  not g26119 (n_10595, n15871);
  and g26120 (n15872, \a[27] , n_10595);
  and g26121 (n15873, n15254, \asqrt[13] );
  not g26122 (n_10596, n15872);
  not g26123 (n_10597, n15873);
  and g26124 (n15874, n_10596, n_10597);
  not g26125 (n_10598, n15870);
  and g26126 (n15875, n_10598, n15874);
  not g26127 (n_10599, n15865);
  not g26128 (n_10600, n15875);
  and g26129 (n15876, n_10599, n_10600);
  not g26130 (n_10601, n15876);
  and g26131 (n15877, \asqrt[15] , n_10601);
  not g26132 (n_10602, \asqrt[15] );
  and g26133 (n15878, n_10602, n_10599);
  and g26134 (n15879, n_10600, n15878);
  not g26138 (n_10603, n15846);
  not g26140 (n_10604, n15883);
  and g26141 (n15884, n_10597, n_10604);
  not g26142 (n_10605, n15884);
  and g26143 (n15885, \a[28] , n_10605);
  and g26144 (n15886, n_9782, n_10604);
  and g26145 (n15887, n_10597, n15886);
  not g26146 (n_10606, n15885);
  not g26147 (n_10607, n15887);
  and g26148 (n15888, n_10606, n_10607);
  not g26149 (n_10608, n15879);
  not g26150 (n_10609, n15888);
  and g26151 (n15889, n_10608, n_10609);
  not g26152 (n_10610, n15877);
  not g26153 (n_10611, n15889);
  and g26154 (n15890, n_10610, n_10611);
  not g26155 (n_10612, n15890);
  and g26156 (n15891, \asqrt[16] , n_10612);
  and g26157 (n15892, n_10191, n_10190);
  not g26158 (n_10613, n15266);
  and g26159 (n15893, n_10613, n15892);
  and g26160 (n15894, \asqrt[13] , n15893);
  and g26161 (n15895, \asqrt[13] , n15892);
  not g26162 (n_10614, n15895);
  and g26163 (n15896, n15266, n_10614);
  not g26164 (n_10615, n15894);
  not g26165 (n_10616, n15896);
  and g26166 (n15897, n_10615, n_10616);
  and g26167 (n15898, n_10194, n_10610);
  and g26168 (n15899, n_10611, n15898);
  not g26169 (n_10617, n15897);
  not g26170 (n_10618, n15899);
  and g26171 (n15900, n_10617, n_10618);
  not g26172 (n_10619, n15891);
  not g26173 (n_10620, n15900);
  and g26174 (n15901, n_10619, n_10620);
  not g26175 (n_10621, n15901);
  and g26176 (n15902, \asqrt[17] , n_10621);
  and g26180 (n15906, n_10202, n_10200);
  and g26181 (n15907, \asqrt[13] , n15906);
  not g26182 (n_10622, n15907);
  and g26183 (n15908, n_10201, n_10622);
  not g26184 (n_10623, n15905);
  not g26185 (n_10624, n15908);
  and g26186 (n15909, n_10623, n_10624);
  and g26187 (n15910, n_9794, n_10619);
  and g26188 (n15911, n_10620, n15910);
  not g26189 (n_10625, n15909);
  not g26190 (n_10626, n15911);
  and g26191 (n15912, n_10625, n_10626);
  not g26192 (n_10627, n15902);
  not g26193 (n_10628, n15912);
  and g26194 (n15913, n_10627, n_10628);
  not g26195 (n_10629, n15913);
  and g26196 (n15914, \asqrt[18] , n_10629);
  and g26200 (n15918, n_10211, n_10210);
  and g26201 (n15919, \asqrt[13] , n15918);
  not g26202 (n_10630, n15919);
  and g26203 (n15920, n_10209, n_10630);
  not g26204 (n_10631, n15917);
  not g26205 (n_10632, n15920);
  and g26206 (n15921, n_10631, n_10632);
  and g26207 (n15922, n_9402, n_10627);
  and g26208 (n15923, n_10628, n15922);
  not g26209 (n_10633, n15921);
  not g26210 (n_10634, n15923);
  and g26211 (n15924, n_10633, n_10634);
  not g26212 (n_10635, n15914);
  not g26213 (n_10636, n15924);
  and g26214 (n15925, n_10635, n_10636);
  not g26215 (n_10637, n15925);
  and g26216 (n15926, \asqrt[19] , n_10637);
  and g26220 (n15930, n_10219, n_10218);
  and g26221 (n15931, \asqrt[13] , n15930);
  not g26222 (n_10638, n15931);
  and g26223 (n15932, n_10217, n_10638);
  not g26224 (n_10639, n15929);
  not g26225 (n_10640, n15932);
  and g26226 (n15933, n_10639, n_10640);
  and g26227 (n15934, n_9018, n_10635);
  and g26228 (n15935, n_10636, n15934);
  not g26229 (n_10641, n15933);
  not g26230 (n_10642, n15935);
  and g26231 (n15936, n_10641, n_10642);
  not g26232 (n_10643, n15926);
  not g26233 (n_10644, n15936);
  and g26234 (n15937, n_10643, n_10644);
  not g26235 (n_10645, n15937);
  and g26236 (n15938, \asqrt[20] , n_10645);
  and g26240 (n15942, n_10227, n_10226);
  and g26241 (n15943, \asqrt[13] , n15942);
  not g26242 (n_10646, n15943);
  and g26243 (n15944, n_10225, n_10646);
  not g26244 (n_10647, n15941);
  not g26245 (n_10648, n15944);
  and g26246 (n15945, n_10647, n_10648);
  and g26247 (n15946, n_8642, n_10643);
  and g26248 (n15947, n_10644, n15946);
  not g26249 (n_10649, n15945);
  not g26250 (n_10650, n15947);
  and g26251 (n15948, n_10649, n_10650);
  not g26252 (n_10651, n15938);
  not g26253 (n_10652, n15948);
  and g26254 (n15949, n_10651, n_10652);
  not g26255 (n_10653, n15949);
  and g26256 (n15950, \asqrt[21] , n_10653);
  and g26260 (n15954, n_10235, n_10234);
  and g26261 (n15955, \asqrt[13] , n15954);
  not g26262 (n_10654, n15955);
  and g26263 (n15956, n_10233, n_10654);
  not g26264 (n_10655, n15953);
  not g26265 (n_10656, n15956);
  and g26266 (n15957, n_10655, n_10656);
  and g26267 (n15958, n_8274, n_10651);
  and g26268 (n15959, n_10652, n15958);
  not g26269 (n_10657, n15957);
  not g26270 (n_10658, n15959);
  and g26271 (n15960, n_10657, n_10658);
  not g26272 (n_10659, n15950);
  not g26273 (n_10660, n15960);
  and g26274 (n15961, n_10659, n_10660);
  not g26275 (n_10661, n15961);
  and g26276 (n15962, \asqrt[22] , n_10661);
  and g26280 (n15966, n_10243, n_10242);
  and g26281 (n15967, \asqrt[13] , n15966);
  not g26282 (n_10662, n15967);
  and g26283 (n15968, n_10241, n_10662);
  not g26284 (n_10663, n15965);
  not g26285 (n_10664, n15968);
  and g26286 (n15969, n_10663, n_10664);
  and g26287 (n15970, n_7914, n_10659);
  and g26288 (n15971, n_10660, n15970);
  not g26289 (n_10665, n15969);
  not g26290 (n_10666, n15971);
  and g26291 (n15972, n_10665, n_10666);
  not g26292 (n_10667, n15962);
  not g26293 (n_10668, n15972);
  and g26294 (n15973, n_10667, n_10668);
  not g26295 (n_10669, n15973);
  and g26296 (n15974, \asqrt[23] , n_10669);
  and g26300 (n15978, n_10251, n_10250);
  and g26301 (n15979, \asqrt[13] , n15978);
  not g26302 (n_10670, n15979);
  and g26303 (n15980, n_10249, n_10670);
  not g26304 (n_10671, n15977);
  not g26305 (n_10672, n15980);
  and g26306 (n15981, n_10671, n_10672);
  and g26307 (n15982, n_7562, n_10667);
  and g26308 (n15983, n_10668, n15982);
  not g26309 (n_10673, n15981);
  not g26310 (n_10674, n15983);
  and g26311 (n15984, n_10673, n_10674);
  not g26312 (n_10675, n15974);
  not g26313 (n_10676, n15984);
  and g26314 (n15985, n_10675, n_10676);
  not g26315 (n_10677, n15985);
  and g26316 (n15986, \asqrt[24] , n_10677);
  and g26320 (n15990, n_10259, n_10258);
  and g26321 (n15991, \asqrt[13] , n15990);
  not g26322 (n_10678, n15991);
  and g26323 (n15992, n_10257, n_10678);
  not g26324 (n_10679, n15989);
  not g26325 (n_10680, n15992);
  and g26326 (n15993, n_10679, n_10680);
  and g26327 (n15994, n_7218, n_10675);
  and g26328 (n15995, n_10676, n15994);
  not g26329 (n_10681, n15993);
  not g26330 (n_10682, n15995);
  and g26331 (n15996, n_10681, n_10682);
  not g26332 (n_10683, n15986);
  not g26333 (n_10684, n15996);
  and g26334 (n15997, n_10683, n_10684);
  not g26335 (n_10685, n15997);
  and g26336 (n15998, \asqrt[25] , n_10685);
  and g26340 (n16002, n_10267, n_10266);
  and g26341 (n16003, \asqrt[13] , n16002);
  not g26342 (n_10686, n16003);
  and g26343 (n16004, n_10265, n_10686);
  not g26344 (n_10687, n16001);
  not g26345 (n_10688, n16004);
  and g26346 (n16005, n_10687, n_10688);
  and g26347 (n16006, n_6882, n_10683);
  and g26348 (n16007, n_10684, n16006);
  not g26349 (n_10689, n16005);
  not g26350 (n_10690, n16007);
  and g26351 (n16008, n_10689, n_10690);
  not g26352 (n_10691, n15998);
  not g26353 (n_10692, n16008);
  and g26354 (n16009, n_10691, n_10692);
  not g26355 (n_10693, n16009);
  and g26356 (n16010, \asqrt[26] , n_10693);
  and g26360 (n16014, n_10275, n_10274);
  and g26361 (n16015, \asqrt[13] , n16014);
  not g26362 (n_10694, n16015);
  and g26363 (n16016, n_10273, n_10694);
  not g26364 (n_10695, n16013);
  not g26365 (n_10696, n16016);
  and g26366 (n16017, n_10695, n_10696);
  and g26367 (n16018, n_6554, n_10691);
  and g26368 (n16019, n_10692, n16018);
  not g26369 (n_10697, n16017);
  not g26370 (n_10698, n16019);
  and g26371 (n16020, n_10697, n_10698);
  not g26372 (n_10699, n16010);
  not g26373 (n_10700, n16020);
  and g26374 (n16021, n_10699, n_10700);
  not g26375 (n_10701, n16021);
  and g26376 (n16022, \asqrt[27] , n_10701);
  and g26380 (n16026, n_10283, n_10282);
  and g26381 (n16027, \asqrt[13] , n16026);
  not g26382 (n_10702, n16027);
  and g26383 (n16028, n_10281, n_10702);
  not g26384 (n_10703, n16025);
  not g26385 (n_10704, n16028);
  and g26386 (n16029, n_10703, n_10704);
  and g26387 (n16030, n_6234, n_10699);
  and g26388 (n16031, n_10700, n16030);
  not g26389 (n_10705, n16029);
  not g26390 (n_10706, n16031);
  and g26391 (n16032, n_10705, n_10706);
  not g26392 (n_10707, n16022);
  not g26393 (n_10708, n16032);
  and g26394 (n16033, n_10707, n_10708);
  not g26395 (n_10709, n16033);
  and g26396 (n16034, \asqrt[28] , n_10709);
  and g26400 (n16038, n_10291, n_10290);
  and g26401 (n16039, \asqrt[13] , n16038);
  not g26402 (n_10710, n16039);
  and g26403 (n16040, n_10289, n_10710);
  not g26404 (n_10711, n16037);
  not g26405 (n_10712, n16040);
  and g26406 (n16041, n_10711, n_10712);
  and g26407 (n16042, n_5922, n_10707);
  and g26408 (n16043, n_10708, n16042);
  not g26409 (n_10713, n16041);
  not g26410 (n_10714, n16043);
  and g26411 (n16044, n_10713, n_10714);
  not g26412 (n_10715, n16034);
  not g26413 (n_10716, n16044);
  and g26414 (n16045, n_10715, n_10716);
  not g26415 (n_10717, n16045);
  and g26416 (n16046, \asqrt[29] , n_10717);
  and g26420 (n16050, n_10299, n_10298);
  and g26421 (n16051, \asqrt[13] , n16050);
  not g26422 (n_10718, n16051);
  and g26423 (n16052, n_10297, n_10718);
  not g26424 (n_10719, n16049);
  not g26425 (n_10720, n16052);
  and g26426 (n16053, n_10719, n_10720);
  and g26427 (n16054, n_5618, n_10715);
  and g26428 (n16055, n_10716, n16054);
  not g26429 (n_10721, n16053);
  not g26430 (n_10722, n16055);
  and g26431 (n16056, n_10721, n_10722);
  not g26432 (n_10723, n16046);
  not g26433 (n_10724, n16056);
  and g26434 (n16057, n_10723, n_10724);
  not g26435 (n_10725, n16057);
  and g26436 (n16058, \asqrt[30] , n_10725);
  and g26440 (n16062, n_10307, n_10306);
  and g26441 (n16063, \asqrt[13] , n16062);
  not g26442 (n_10726, n16063);
  and g26443 (n16064, n_10305, n_10726);
  not g26444 (n_10727, n16061);
  not g26445 (n_10728, n16064);
  and g26446 (n16065, n_10727, n_10728);
  and g26447 (n16066, n_5322, n_10723);
  and g26448 (n16067, n_10724, n16066);
  not g26449 (n_10729, n16065);
  not g26450 (n_10730, n16067);
  and g26451 (n16068, n_10729, n_10730);
  not g26452 (n_10731, n16058);
  not g26453 (n_10732, n16068);
  and g26454 (n16069, n_10731, n_10732);
  not g26455 (n_10733, n16069);
  and g26456 (n16070, \asqrt[31] , n_10733);
  and g26460 (n16074, n_10315, n_10314);
  and g26461 (n16075, \asqrt[13] , n16074);
  not g26462 (n_10734, n16075);
  and g26463 (n16076, n_10313, n_10734);
  not g26464 (n_10735, n16073);
  not g26465 (n_10736, n16076);
  and g26466 (n16077, n_10735, n_10736);
  and g26467 (n16078, n_5034, n_10731);
  and g26468 (n16079, n_10732, n16078);
  not g26469 (n_10737, n16077);
  not g26470 (n_10738, n16079);
  and g26471 (n16080, n_10737, n_10738);
  not g26472 (n_10739, n16070);
  not g26473 (n_10740, n16080);
  and g26474 (n16081, n_10739, n_10740);
  not g26475 (n_10741, n16081);
  and g26476 (n16082, \asqrt[32] , n_10741);
  and g26480 (n16086, n_10323, n_10322);
  and g26481 (n16087, \asqrt[13] , n16086);
  not g26482 (n_10742, n16087);
  and g26483 (n16088, n_10321, n_10742);
  not g26484 (n_10743, n16085);
  not g26485 (n_10744, n16088);
  and g26486 (n16089, n_10743, n_10744);
  and g26487 (n16090, n_4754, n_10739);
  and g26488 (n16091, n_10740, n16090);
  not g26489 (n_10745, n16089);
  not g26490 (n_10746, n16091);
  and g26491 (n16092, n_10745, n_10746);
  not g26492 (n_10747, n16082);
  not g26493 (n_10748, n16092);
  and g26494 (n16093, n_10747, n_10748);
  not g26495 (n_10749, n16093);
  and g26496 (n16094, \asqrt[33] , n_10749);
  and g26500 (n16098, n_10331, n_10330);
  and g26501 (n16099, \asqrt[13] , n16098);
  not g26502 (n_10750, n16099);
  and g26503 (n16100, n_10329, n_10750);
  not g26504 (n_10751, n16097);
  not g26505 (n_10752, n16100);
  and g26506 (n16101, n_10751, n_10752);
  and g26507 (n16102, n_4482, n_10747);
  and g26508 (n16103, n_10748, n16102);
  not g26509 (n_10753, n16101);
  not g26510 (n_10754, n16103);
  and g26511 (n16104, n_10753, n_10754);
  not g26512 (n_10755, n16094);
  not g26513 (n_10756, n16104);
  and g26514 (n16105, n_10755, n_10756);
  not g26515 (n_10757, n16105);
  and g26516 (n16106, \asqrt[34] , n_10757);
  and g26520 (n16110, n_10339, n_10338);
  and g26521 (n16111, \asqrt[13] , n16110);
  not g26522 (n_10758, n16111);
  and g26523 (n16112, n_10337, n_10758);
  not g26524 (n_10759, n16109);
  not g26525 (n_10760, n16112);
  and g26526 (n16113, n_10759, n_10760);
  and g26527 (n16114, n_4218, n_10755);
  and g26528 (n16115, n_10756, n16114);
  not g26529 (n_10761, n16113);
  not g26530 (n_10762, n16115);
  and g26531 (n16116, n_10761, n_10762);
  not g26532 (n_10763, n16106);
  not g26533 (n_10764, n16116);
  and g26534 (n16117, n_10763, n_10764);
  not g26535 (n_10765, n16117);
  and g26536 (n16118, \asqrt[35] , n_10765);
  and g26540 (n16122, n_10347, n_10346);
  and g26541 (n16123, \asqrt[13] , n16122);
  not g26542 (n_10766, n16123);
  and g26543 (n16124, n_10345, n_10766);
  not g26544 (n_10767, n16121);
  not g26545 (n_10768, n16124);
  and g26546 (n16125, n_10767, n_10768);
  and g26547 (n16126, n_3962, n_10763);
  and g26548 (n16127, n_10764, n16126);
  not g26549 (n_10769, n16125);
  not g26550 (n_10770, n16127);
  and g26551 (n16128, n_10769, n_10770);
  not g26552 (n_10771, n16118);
  not g26553 (n_10772, n16128);
  and g26554 (n16129, n_10771, n_10772);
  not g26555 (n_10773, n16129);
  and g26556 (n16130, \asqrt[36] , n_10773);
  and g26560 (n16134, n_10355, n_10354);
  and g26561 (n16135, \asqrt[13] , n16134);
  not g26562 (n_10774, n16135);
  and g26563 (n16136, n_10353, n_10774);
  not g26564 (n_10775, n16133);
  not g26565 (n_10776, n16136);
  and g26566 (n16137, n_10775, n_10776);
  and g26567 (n16138, n_3714, n_10771);
  and g26568 (n16139, n_10772, n16138);
  not g26569 (n_10777, n16137);
  not g26570 (n_10778, n16139);
  and g26571 (n16140, n_10777, n_10778);
  not g26572 (n_10779, n16130);
  not g26573 (n_10780, n16140);
  and g26574 (n16141, n_10779, n_10780);
  not g26575 (n_10781, n16141);
  and g26576 (n16142, \asqrt[37] , n_10781);
  and g26580 (n16146, n_10363, n_10362);
  and g26581 (n16147, \asqrt[13] , n16146);
  not g26582 (n_10782, n16147);
  and g26583 (n16148, n_10361, n_10782);
  not g26584 (n_10783, n16145);
  not g26585 (n_10784, n16148);
  and g26586 (n16149, n_10783, n_10784);
  and g26587 (n16150, n_3474, n_10779);
  and g26588 (n16151, n_10780, n16150);
  not g26589 (n_10785, n16149);
  not g26590 (n_10786, n16151);
  and g26591 (n16152, n_10785, n_10786);
  not g26592 (n_10787, n16142);
  not g26593 (n_10788, n16152);
  and g26594 (n16153, n_10787, n_10788);
  not g26595 (n_10789, n16153);
  and g26596 (n16154, \asqrt[38] , n_10789);
  and g26600 (n16158, n_10371, n_10370);
  and g26601 (n16159, \asqrt[13] , n16158);
  not g26602 (n_10790, n16159);
  and g26603 (n16160, n_10369, n_10790);
  not g26604 (n_10791, n16157);
  not g26605 (n_10792, n16160);
  and g26606 (n16161, n_10791, n_10792);
  and g26607 (n16162, n_3242, n_10787);
  and g26608 (n16163, n_10788, n16162);
  not g26609 (n_10793, n16161);
  not g26610 (n_10794, n16163);
  and g26611 (n16164, n_10793, n_10794);
  not g26612 (n_10795, n16154);
  not g26613 (n_10796, n16164);
  and g26614 (n16165, n_10795, n_10796);
  not g26615 (n_10797, n16165);
  and g26616 (n16166, \asqrt[39] , n_10797);
  and g26620 (n16170, n_10379, n_10378);
  and g26621 (n16171, \asqrt[13] , n16170);
  not g26622 (n_10798, n16171);
  and g26623 (n16172, n_10377, n_10798);
  not g26624 (n_10799, n16169);
  not g26625 (n_10800, n16172);
  and g26626 (n16173, n_10799, n_10800);
  and g26627 (n16174, n_3018, n_10795);
  and g26628 (n16175, n_10796, n16174);
  not g26629 (n_10801, n16173);
  not g26630 (n_10802, n16175);
  and g26631 (n16176, n_10801, n_10802);
  not g26632 (n_10803, n16166);
  not g26633 (n_10804, n16176);
  and g26634 (n16177, n_10803, n_10804);
  not g26635 (n_10805, n16177);
  and g26636 (n16178, \asqrt[40] , n_10805);
  and g26640 (n16182, n_10387, n_10386);
  and g26641 (n16183, \asqrt[13] , n16182);
  not g26642 (n_10806, n16183);
  and g26643 (n16184, n_10385, n_10806);
  not g26644 (n_10807, n16181);
  not g26645 (n_10808, n16184);
  and g26646 (n16185, n_10807, n_10808);
  and g26647 (n16186, n_2802, n_10803);
  and g26648 (n16187, n_10804, n16186);
  not g26649 (n_10809, n16185);
  not g26650 (n_10810, n16187);
  and g26651 (n16188, n_10809, n_10810);
  not g26652 (n_10811, n16178);
  not g26653 (n_10812, n16188);
  and g26654 (n16189, n_10811, n_10812);
  not g26655 (n_10813, n16189);
  and g26656 (n16190, \asqrt[41] , n_10813);
  and g26660 (n16194, n_10395, n_10394);
  and g26661 (n16195, \asqrt[13] , n16194);
  not g26662 (n_10814, n16195);
  and g26663 (n16196, n_10393, n_10814);
  not g26664 (n_10815, n16193);
  not g26665 (n_10816, n16196);
  and g26666 (n16197, n_10815, n_10816);
  and g26667 (n16198, n_2594, n_10811);
  and g26668 (n16199, n_10812, n16198);
  not g26669 (n_10817, n16197);
  not g26670 (n_10818, n16199);
  and g26671 (n16200, n_10817, n_10818);
  not g26672 (n_10819, n16190);
  not g26673 (n_10820, n16200);
  and g26674 (n16201, n_10819, n_10820);
  not g26675 (n_10821, n16201);
  and g26676 (n16202, \asqrt[42] , n_10821);
  and g26680 (n16206, n_10403, n_10402);
  and g26681 (n16207, \asqrt[13] , n16206);
  not g26682 (n_10822, n16207);
  and g26683 (n16208, n_10401, n_10822);
  not g26684 (n_10823, n16205);
  not g26685 (n_10824, n16208);
  and g26686 (n16209, n_10823, n_10824);
  and g26687 (n16210, n_2394, n_10819);
  and g26688 (n16211, n_10820, n16210);
  not g26689 (n_10825, n16209);
  not g26690 (n_10826, n16211);
  and g26691 (n16212, n_10825, n_10826);
  not g26692 (n_10827, n16202);
  not g26693 (n_10828, n16212);
  and g26694 (n16213, n_10827, n_10828);
  not g26695 (n_10829, n16213);
  and g26696 (n16214, \asqrt[43] , n_10829);
  and g26700 (n16218, n_10411, n_10410);
  and g26701 (n16219, \asqrt[13] , n16218);
  not g26702 (n_10830, n16219);
  and g26703 (n16220, n_10409, n_10830);
  not g26704 (n_10831, n16217);
  not g26705 (n_10832, n16220);
  and g26706 (n16221, n_10831, n_10832);
  and g26707 (n16222, n_2202, n_10827);
  and g26708 (n16223, n_10828, n16222);
  not g26709 (n_10833, n16221);
  not g26710 (n_10834, n16223);
  and g26711 (n16224, n_10833, n_10834);
  not g26712 (n_10835, n16214);
  not g26713 (n_10836, n16224);
  and g26714 (n16225, n_10835, n_10836);
  not g26715 (n_10837, n16225);
  and g26716 (n16226, \asqrt[44] , n_10837);
  and g26720 (n16230, n_10419, n_10418);
  and g26721 (n16231, \asqrt[13] , n16230);
  not g26722 (n_10838, n16231);
  and g26723 (n16232, n_10417, n_10838);
  not g26724 (n_10839, n16229);
  not g26725 (n_10840, n16232);
  and g26726 (n16233, n_10839, n_10840);
  and g26727 (n16234, n_2018, n_10835);
  and g26728 (n16235, n_10836, n16234);
  not g26729 (n_10841, n16233);
  not g26730 (n_10842, n16235);
  and g26731 (n16236, n_10841, n_10842);
  not g26732 (n_10843, n16226);
  not g26733 (n_10844, n16236);
  and g26734 (n16237, n_10843, n_10844);
  not g26735 (n_10845, n16237);
  and g26736 (n16238, \asqrt[45] , n_10845);
  and g26740 (n16242, n_10427, n_10426);
  and g26741 (n16243, \asqrt[13] , n16242);
  not g26742 (n_10846, n16243);
  and g26743 (n16244, n_10425, n_10846);
  not g26744 (n_10847, n16241);
  not g26745 (n_10848, n16244);
  and g26746 (n16245, n_10847, n_10848);
  and g26747 (n16246, n_1842, n_10843);
  and g26748 (n16247, n_10844, n16246);
  not g26749 (n_10849, n16245);
  not g26750 (n_10850, n16247);
  and g26751 (n16248, n_10849, n_10850);
  not g26752 (n_10851, n16238);
  not g26753 (n_10852, n16248);
  and g26754 (n16249, n_10851, n_10852);
  not g26755 (n_10853, n16249);
  and g26756 (n16250, \asqrt[46] , n_10853);
  and g26760 (n16254, n_10435, n_10434);
  and g26761 (n16255, \asqrt[13] , n16254);
  not g26762 (n_10854, n16255);
  and g26763 (n16256, n_10433, n_10854);
  not g26764 (n_10855, n16253);
  not g26765 (n_10856, n16256);
  and g26766 (n16257, n_10855, n_10856);
  and g26767 (n16258, n_1674, n_10851);
  and g26768 (n16259, n_10852, n16258);
  not g26769 (n_10857, n16257);
  not g26770 (n_10858, n16259);
  and g26771 (n16260, n_10857, n_10858);
  not g26772 (n_10859, n16250);
  not g26773 (n_10860, n16260);
  and g26774 (n16261, n_10859, n_10860);
  not g26775 (n_10861, n16261);
  and g26776 (n16262, \asqrt[47] , n_10861);
  and g26780 (n16266, n_10443, n_10442);
  and g26781 (n16267, \asqrt[13] , n16266);
  not g26782 (n_10862, n16267);
  and g26783 (n16268, n_10441, n_10862);
  not g26784 (n_10863, n16265);
  not g26785 (n_10864, n16268);
  and g26786 (n16269, n_10863, n_10864);
  and g26787 (n16270, n_1514, n_10859);
  and g26788 (n16271, n_10860, n16270);
  not g26789 (n_10865, n16269);
  not g26790 (n_10866, n16271);
  and g26791 (n16272, n_10865, n_10866);
  not g26792 (n_10867, n16262);
  not g26793 (n_10868, n16272);
  and g26794 (n16273, n_10867, n_10868);
  not g26795 (n_10869, n16273);
  and g26796 (n16274, \asqrt[48] , n_10869);
  and g26800 (n16278, n_10451, n_10450);
  and g26801 (n16279, \asqrt[13] , n16278);
  not g26802 (n_10870, n16279);
  and g26803 (n16280, n_10449, n_10870);
  not g26804 (n_10871, n16277);
  not g26805 (n_10872, n16280);
  and g26806 (n16281, n_10871, n_10872);
  and g26807 (n16282, n_1362, n_10867);
  and g26808 (n16283, n_10868, n16282);
  not g26809 (n_10873, n16281);
  not g26810 (n_10874, n16283);
  and g26811 (n16284, n_10873, n_10874);
  not g26812 (n_10875, n16274);
  not g26813 (n_10876, n16284);
  and g26814 (n16285, n_10875, n_10876);
  not g26815 (n_10877, n16285);
  and g26816 (n16286, \asqrt[49] , n_10877);
  and g26820 (n16290, n_10459, n_10458);
  and g26821 (n16291, \asqrt[13] , n16290);
  not g26822 (n_10878, n16291);
  and g26823 (n16292, n_10457, n_10878);
  not g26824 (n_10879, n16289);
  not g26825 (n_10880, n16292);
  and g26826 (n16293, n_10879, n_10880);
  and g26827 (n16294, n_1218, n_10875);
  and g26828 (n16295, n_10876, n16294);
  not g26829 (n_10881, n16293);
  not g26830 (n_10882, n16295);
  and g26831 (n16296, n_10881, n_10882);
  not g26832 (n_10883, n16286);
  not g26833 (n_10884, n16296);
  and g26834 (n16297, n_10883, n_10884);
  not g26835 (n_10885, n16297);
  and g26836 (n16298, \asqrt[50] , n_10885);
  and g26840 (n16302, n_10467, n_10466);
  and g26841 (n16303, \asqrt[13] , n16302);
  not g26842 (n_10886, n16303);
  and g26843 (n16304, n_10465, n_10886);
  not g26844 (n_10887, n16301);
  not g26845 (n_10888, n16304);
  and g26846 (n16305, n_10887, n_10888);
  and g26847 (n16306, n_1082, n_10883);
  and g26848 (n16307, n_10884, n16306);
  not g26849 (n_10889, n16305);
  not g26850 (n_10890, n16307);
  and g26851 (n16308, n_10889, n_10890);
  not g26852 (n_10891, n16298);
  not g26853 (n_10892, n16308);
  and g26854 (n16309, n_10891, n_10892);
  not g26855 (n_10893, n16309);
  and g26856 (n16310, \asqrt[51] , n_10893);
  and g26860 (n16314, n_10475, n_10474);
  and g26861 (n16315, \asqrt[13] , n16314);
  not g26862 (n_10894, n16315);
  and g26863 (n16316, n_10473, n_10894);
  not g26864 (n_10895, n16313);
  not g26865 (n_10896, n16316);
  and g26866 (n16317, n_10895, n_10896);
  and g26867 (n16318, n_954, n_10891);
  and g26868 (n16319, n_10892, n16318);
  not g26869 (n_10897, n16317);
  not g26870 (n_10898, n16319);
  and g26871 (n16320, n_10897, n_10898);
  not g26872 (n_10899, n16310);
  not g26873 (n_10900, n16320);
  and g26874 (n16321, n_10899, n_10900);
  not g26875 (n_10901, n16321);
  and g26876 (n16322, \asqrt[52] , n_10901);
  and g26877 (n16323, n_834, n_10899);
  and g26878 (n16324, n_10900, n16323);
  and g26882 (n16328, n_10483, n_10481);
  and g26883 (n16329, \asqrt[13] , n16328);
  not g26884 (n_10902, n16329);
  and g26885 (n16330, n_10482, n_10902);
  not g26886 (n_10903, n16327);
  not g26887 (n_10904, n16330);
  and g26888 (n16331, n_10903, n_10904);
  not g26889 (n_10905, n16324);
  not g26890 (n_10906, n16331);
  and g26891 (n16332, n_10905, n_10906);
  not g26892 (n_10907, n16322);
  not g26893 (n_10908, n16332);
  and g26894 (n16333, n_10907, n_10908);
  not g26895 (n_10909, n16333);
  and g26896 (n16334, \asqrt[53] , n_10909);
  and g26900 (n16338, n_10491, n_10490);
  and g26901 (n16339, \asqrt[13] , n16338);
  not g26902 (n_10910, n16339);
  and g26903 (n16340, n_10489, n_10910);
  not g26904 (n_10911, n16337);
  not g26905 (n_10912, n16340);
  and g26906 (n16341, n_10911, n_10912);
  and g26907 (n16342, n_722, n_10907);
  and g26908 (n16343, n_10908, n16342);
  not g26909 (n_10913, n16341);
  not g26910 (n_10914, n16343);
  and g26911 (n16344, n_10913, n_10914);
  not g26912 (n_10915, n16334);
  not g26913 (n_10916, n16344);
  and g26914 (n16345, n_10915, n_10916);
  not g26915 (n_10917, n16345);
  and g26916 (n16346, \asqrt[54] , n_10917);
  and g26920 (n16350, n_10499, n_10498);
  and g26921 (n16351, \asqrt[13] , n16350);
  not g26922 (n_10918, n16351);
  and g26923 (n16352, n_10497, n_10918);
  not g26924 (n_10919, n16349);
  not g26925 (n_10920, n16352);
  and g26926 (n16353, n_10919, n_10920);
  and g26927 (n16354, n_618, n_10915);
  and g26928 (n16355, n_10916, n16354);
  not g26929 (n_10921, n16353);
  not g26930 (n_10922, n16355);
  and g26931 (n16356, n_10921, n_10922);
  not g26932 (n_10923, n16346);
  not g26933 (n_10924, n16356);
  and g26934 (n16357, n_10923, n_10924);
  not g26935 (n_10925, n16357);
  and g26936 (n16358, \asqrt[55] , n_10925);
  and g26940 (n16362, n_10507, n_10506);
  and g26941 (n16363, \asqrt[13] , n16362);
  not g26942 (n_10926, n16363);
  and g26943 (n16364, n_10505, n_10926);
  not g26944 (n_10927, n16361);
  not g26945 (n_10928, n16364);
  and g26946 (n16365, n_10927, n_10928);
  and g26947 (n16366, n_522, n_10923);
  and g26948 (n16367, n_10924, n16366);
  not g26949 (n_10929, n16365);
  not g26950 (n_10930, n16367);
  and g26951 (n16368, n_10929, n_10930);
  not g26952 (n_10931, n16358);
  not g26953 (n_10932, n16368);
  and g26954 (n16369, n_10931, n_10932);
  not g26955 (n_10933, n16369);
  and g26956 (n16370, \asqrt[56] , n_10933);
  and g26960 (n16374, n_10515, n_10514);
  and g26961 (n16375, \asqrt[13] , n16374);
  not g26962 (n_10934, n16375);
  and g26963 (n16376, n_10513, n_10934);
  not g26964 (n_10935, n16373);
  not g26965 (n_10936, n16376);
  and g26966 (n16377, n_10935, n_10936);
  and g26967 (n16378, n_434, n_10931);
  and g26968 (n16379, n_10932, n16378);
  not g26969 (n_10937, n16377);
  not g26970 (n_10938, n16379);
  and g26971 (n16380, n_10937, n_10938);
  not g26972 (n_10939, n16370);
  not g26973 (n_10940, n16380);
  and g26974 (n16381, n_10939, n_10940);
  not g26975 (n_10941, n16381);
  and g26976 (n16382, \asqrt[57] , n_10941);
  and g26980 (n16386, n_10523, n_10522);
  and g26981 (n16387, \asqrt[13] , n16386);
  not g26982 (n_10942, n16387);
  and g26983 (n16388, n_10521, n_10942);
  not g26984 (n_10943, n16385);
  not g26985 (n_10944, n16388);
  and g26986 (n16389, n_10943, n_10944);
  and g26987 (n16390, n_354, n_10939);
  and g26988 (n16391, n_10940, n16390);
  not g26989 (n_10945, n16389);
  not g26990 (n_10946, n16391);
  and g26991 (n16392, n_10945, n_10946);
  not g26992 (n_10947, n16382);
  not g26993 (n_10948, n16392);
  and g26994 (n16393, n_10947, n_10948);
  not g26995 (n_10949, n16393);
  and g26996 (n16394, \asqrt[58] , n_10949);
  and g27000 (n16398, n_10531, n_10530);
  and g27001 (n16399, \asqrt[13] , n16398);
  not g27002 (n_10950, n16399);
  and g27003 (n16400, n_10529, n_10950);
  not g27004 (n_10951, n16397);
  not g27005 (n_10952, n16400);
  and g27006 (n16401, n_10951, n_10952);
  and g27007 (n16402, n_282, n_10947);
  and g27008 (n16403, n_10948, n16402);
  not g27009 (n_10953, n16401);
  not g27010 (n_10954, n16403);
  and g27011 (n16404, n_10953, n_10954);
  not g27012 (n_10955, n16394);
  not g27013 (n_10956, n16404);
  and g27014 (n16405, n_10955, n_10956);
  not g27015 (n_10957, n16405);
  and g27016 (n16406, \asqrt[59] , n_10957);
  and g27020 (n16410, n_10539, n_10538);
  and g27021 (n16411, \asqrt[13] , n16410);
  not g27022 (n_10958, n16411);
  and g27023 (n16412, n_10537, n_10958);
  not g27024 (n_10959, n16409);
  not g27025 (n_10960, n16412);
  and g27026 (n16413, n_10959, n_10960);
  and g27027 (n16414, n_218, n_10955);
  and g27028 (n16415, n_10956, n16414);
  not g27029 (n_10961, n16413);
  not g27030 (n_10962, n16415);
  and g27031 (n16416, n_10961, n_10962);
  not g27032 (n_10963, n16406);
  not g27033 (n_10964, n16416);
  and g27034 (n16417, n_10963, n_10964);
  not g27035 (n_10965, n16417);
  and g27036 (n16418, \asqrt[60] , n_10965);
  and g27040 (n16422, n_10547, n_10546);
  and g27041 (n16423, \asqrt[13] , n16422);
  not g27042 (n_10966, n16423);
  and g27043 (n16424, n_10545, n_10966);
  not g27044 (n_10967, n16421);
  not g27045 (n_10968, n16424);
  and g27046 (n16425, n_10967, n_10968);
  and g27047 (n16426, n_162, n_10963);
  and g27048 (n16427, n_10964, n16426);
  not g27049 (n_10969, n16425);
  not g27050 (n_10970, n16427);
  and g27051 (n16428, n_10969, n_10970);
  not g27052 (n_10971, n16418);
  not g27053 (n_10972, n16428);
  and g27054 (n16429, n_10971, n_10972);
  not g27055 (n_10973, n16429);
  and g27056 (n16430, \asqrt[61] , n_10973);
  and g27060 (n16434, n_10555, n_10554);
  and g27061 (n16435, \asqrt[13] , n16434);
  not g27062 (n_10974, n16435);
  and g27063 (n16436, n_10553, n_10974);
  not g27064 (n_10975, n16433);
  not g27065 (n_10976, n16436);
  and g27066 (n16437, n_10975, n_10976);
  and g27067 (n16438, n_115, n_10971);
  and g27068 (n16439, n_10972, n16438);
  not g27069 (n_10977, n16437);
  not g27070 (n_10978, n16439);
  and g27071 (n16440, n_10977, n_10978);
  not g27072 (n_10979, n16430);
  not g27073 (n_10980, n16440);
  and g27074 (n16441, n_10979, n_10980);
  not g27075 (n_10981, n16441);
  and g27076 (n16442, \asqrt[62] , n_10981);
  and g27080 (n16446, n_10563, n_10562);
  and g27081 (n16447, \asqrt[13] , n16446);
  not g27082 (n_10982, n16447);
  and g27083 (n16448, n_10561, n_10982);
  not g27084 (n_10983, n16445);
  not g27085 (n_10984, n16448);
  and g27086 (n16449, n_10983, n_10984);
  and g27087 (n16450, n_76, n_10979);
  and g27088 (n16451, n_10980, n16450);
  not g27089 (n_10985, n16449);
  not g27090 (n_10986, n16451);
  and g27091 (n16452, n_10985, n_10986);
  not g27092 (n_10987, n16442);
  not g27093 (n_10988, n16452);
  and g27094 (n16453, n_10987, n_10988);
  and g27098 (n16457, n_10571, n_10570);
  and g27099 (n16458, \asqrt[13] , n16457);
  not g27100 (n_10989, n16458);
  and g27101 (n16459, n_10569, n_10989);
  not g27102 (n_10990, n16456);
  not g27103 (n_10991, n16459);
  and g27104 (n16460, n_10990, n_10991);
  and g27105 (n16461, n_10578, n_10577);
  and g27106 (n16462, \asqrt[13] , n16461);
  not g27109 (n_10993, n16460);
  not g27111 (n_10994, n16453);
  not g27113 (n_10995, n16465);
  and g27114 (n16466, n_21, n_10995);
  and g27115 (n16467, n_10987, n16460);
  and g27116 (n16468, n_10988, n16467);
  and g27117 (n16469, n_10577, \asqrt[13] );
  not g27118 (n_10996, n16469);
  and g27119 (n16470, n15833, n_10996);
  not g27120 (n_10997, n16461);
  and g27121 (n16471, \asqrt[63] , n_10997);
  not g27122 (n_10998, n16470);
  and g27123 (n16472, n_10998, n16471);
  not g27129 (n_10999, n16472);
  not g27130 (n_11000, n16477);
  not g27132 (n_11001, n16468);
  and g27136 (n16481, \a[24] , \asqrt[12] );
  not g27137 (n_11006, \a[22] );
  not g27138 (n_11007, \a[23] );
  and g27139 (n16482, n_11006, n_11007);
  and g27140 (n16483, n_10590, n16482);
  not g27141 (n_11008, n16481);
  not g27142 (n_11009, n16483);
  and g27143 (n16484, n_11008, n_11009);
  not g27144 (n_11010, n16484);
  and g27145 (n16485, \asqrt[13] , n_11010);
  and g27151 (n16491, n_10590, \asqrt[12] );
  not g27152 (n_11011, n16491);
  and g27153 (n16492, \a[25] , n_11011);
  and g27154 (n16493, n15862, \asqrt[12] );
  not g27155 (n_11012, n16492);
  not g27156 (n_11013, n16493);
  and g27157 (n16494, n_11012, n_11013);
  not g27158 (n_11014, n16490);
  and g27159 (n16495, n_11014, n16494);
  not g27160 (n_11015, n16485);
  not g27161 (n_11016, n16495);
  and g27162 (n16496, n_11015, n_11016);
  not g27163 (n_11017, n16496);
  and g27164 (n16497, \asqrt[14] , n_11017);
  not g27165 (n_11018, \asqrt[14] );
  and g27166 (n16498, n_11018, n_11015);
  and g27167 (n16499, n_11016, n16498);
  not g27171 (n_11019, n16466);
  not g27173 (n_11020, n16503);
  and g27174 (n16504, n_11013, n_11020);
  not g27175 (n_11021, n16504);
  and g27176 (n16505, \a[26] , n_11021);
  and g27177 (n16506, n_10182, n_11020);
  and g27178 (n16507, n_11013, n16506);
  not g27179 (n_11022, n16505);
  not g27180 (n_11023, n16507);
  and g27181 (n16508, n_11022, n_11023);
  not g27182 (n_11024, n16499);
  not g27183 (n_11025, n16508);
  and g27184 (n16509, n_11024, n_11025);
  not g27185 (n_11026, n16497);
  not g27186 (n_11027, n16509);
  and g27187 (n16510, n_11026, n_11027);
  not g27188 (n_11028, n16510);
  and g27189 (n16511, \asqrt[15] , n_11028);
  and g27190 (n16512, n_10599, n_10598);
  not g27191 (n_11029, n15874);
  and g27192 (n16513, n_11029, n16512);
  and g27193 (n16514, \asqrt[12] , n16513);
  and g27194 (n16515, \asqrt[12] , n16512);
  not g27195 (n_11030, n16515);
  and g27196 (n16516, n15874, n_11030);
  not g27197 (n_11031, n16514);
  not g27198 (n_11032, n16516);
  and g27199 (n16517, n_11031, n_11032);
  and g27200 (n16518, n_10602, n_11026);
  and g27201 (n16519, n_11027, n16518);
  not g27202 (n_11033, n16517);
  not g27203 (n_11034, n16519);
  and g27204 (n16520, n_11033, n_11034);
  not g27205 (n_11035, n16511);
  not g27206 (n_11036, n16520);
  and g27207 (n16521, n_11035, n_11036);
  not g27208 (n_11037, n16521);
  and g27209 (n16522, \asqrt[16] , n_11037);
  and g27213 (n16526, n_10610, n_10608);
  and g27214 (n16527, \asqrt[12] , n16526);
  not g27215 (n_11038, n16527);
  and g27216 (n16528, n_10609, n_11038);
  not g27217 (n_11039, n16525);
  not g27218 (n_11040, n16528);
  and g27219 (n16529, n_11039, n_11040);
  and g27220 (n16530, n_10194, n_11035);
  and g27221 (n16531, n_11036, n16530);
  not g27222 (n_11041, n16529);
  not g27223 (n_11042, n16531);
  and g27224 (n16532, n_11041, n_11042);
  not g27225 (n_11043, n16522);
  not g27226 (n_11044, n16532);
  and g27227 (n16533, n_11043, n_11044);
  not g27228 (n_11045, n16533);
  and g27229 (n16534, \asqrt[17] , n_11045);
  and g27233 (n16538, n_10619, n_10618);
  and g27234 (n16539, \asqrt[12] , n16538);
  not g27235 (n_11046, n16539);
  and g27236 (n16540, n_10617, n_11046);
  not g27237 (n_11047, n16537);
  not g27238 (n_11048, n16540);
  and g27239 (n16541, n_11047, n_11048);
  and g27240 (n16542, n_9794, n_11043);
  and g27241 (n16543, n_11044, n16542);
  not g27242 (n_11049, n16541);
  not g27243 (n_11050, n16543);
  and g27244 (n16544, n_11049, n_11050);
  not g27245 (n_11051, n16534);
  not g27246 (n_11052, n16544);
  and g27247 (n16545, n_11051, n_11052);
  not g27248 (n_11053, n16545);
  and g27249 (n16546, \asqrt[18] , n_11053);
  and g27253 (n16550, n_10627, n_10626);
  and g27254 (n16551, \asqrt[12] , n16550);
  not g27255 (n_11054, n16551);
  and g27256 (n16552, n_10625, n_11054);
  not g27257 (n_11055, n16549);
  not g27258 (n_11056, n16552);
  and g27259 (n16553, n_11055, n_11056);
  and g27260 (n16554, n_9402, n_11051);
  and g27261 (n16555, n_11052, n16554);
  not g27262 (n_11057, n16553);
  not g27263 (n_11058, n16555);
  and g27264 (n16556, n_11057, n_11058);
  not g27265 (n_11059, n16546);
  not g27266 (n_11060, n16556);
  and g27267 (n16557, n_11059, n_11060);
  not g27268 (n_11061, n16557);
  and g27269 (n16558, \asqrt[19] , n_11061);
  and g27273 (n16562, n_10635, n_10634);
  and g27274 (n16563, \asqrt[12] , n16562);
  not g27275 (n_11062, n16563);
  and g27276 (n16564, n_10633, n_11062);
  not g27277 (n_11063, n16561);
  not g27278 (n_11064, n16564);
  and g27279 (n16565, n_11063, n_11064);
  and g27280 (n16566, n_9018, n_11059);
  and g27281 (n16567, n_11060, n16566);
  not g27282 (n_11065, n16565);
  not g27283 (n_11066, n16567);
  and g27284 (n16568, n_11065, n_11066);
  not g27285 (n_11067, n16558);
  not g27286 (n_11068, n16568);
  and g27287 (n16569, n_11067, n_11068);
  not g27288 (n_11069, n16569);
  and g27289 (n16570, \asqrt[20] , n_11069);
  and g27293 (n16574, n_10643, n_10642);
  and g27294 (n16575, \asqrt[12] , n16574);
  not g27295 (n_11070, n16575);
  and g27296 (n16576, n_10641, n_11070);
  not g27297 (n_11071, n16573);
  not g27298 (n_11072, n16576);
  and g27299 (n16577, n_11071, n_11072);
  and g27300 (n16578, n_8642, n_11067);
  and g27301 (n16579, n_11068, n16578);
  not g27302 (n_11073, n16577);
  not g27303 (n_11074, n16579);
  and g27304 (n16580, n_11073, n_11074);
  not g27305 (n_11075, n16570);
  not g27306 (n_11076, n16580);
  and g27307 (n16581, n_11075, n_11076);
  not g27308 (n_11077, n16581);
  and g27309 (n16582, \asqrt[21] , n_11077);
  and g27313 (n16586, n_10651, n_10650);
  and g27314 (n16587, \asqrt[12] , n16586);
  not g27315 (n_11078, n16587);
  and g27316 (n16588, n_10649, n_11078);
  not g27317 (n_11079, n16585);
  not g27318 (n_11080, n16588);
  and g27319 (n16589, n_11079, n_11080);
  and g27320 (n16590, n_8274, n_11075);
  and g27321 (n16591, n_11076, n16590);
  not g27322 (n_11081, n16589);
  not g27323 (n_11082, n16591);
  and g27324 (n16592, n_11081, n_11082);
  not g27325 (n_11083, n16582);
  not g27326 (n_11084, n16592);
  and g27327 (n16593, n_11083, n_11084);
  not g27328 (n_11085, n16593);
  and g27329 (n16594, \asqrt[22] , n_11085);
  and g27333 (n16598, n_10659, n_10658);
  and g27334 (n16599, \asqrt[12] , n16598);
  not g27335 (n_11086, n16599);
  and g27336 (n16600, n_10657, n_11086);
  not g27337 (n_11087, n16597);
  not g27338 (n_11088, n16600);
  and g27339 (n16601, n_11087, n_11088);
  and g27340 (n16602, n_7914, n_11083);
  and g27341 (n16603, n_11084, n16602);
  not g27342 (n_11089, n16601);
  not g27343 (n_11090, n16603);
  and g27344 (n16604, n_11089, n_11090);
  not g27345 (n_11091, n16594);
  not g27346 (n_11092, n16604);
  and g27347 (n16605, n_11091, n_11092);
  not g27348 (n_11093, n16605);
  and g27349 (n16606, \asqrt[23] , n_11093);
  and g27353 (n16610, n_10667, n_10666);
  and g27354 (n16611, \asqrt[12] , n16610);
  not g27355 (n_11094, n16611);
  and g27356 (n16612, n_10665, n_11094);
  not g27357 (n_11095, n16609);
  not g27358 (n_11096, n16612);
  and g27359 (n16613, n_11095, n_11096);
  and g27360 (n16614, n_7562, n_11091);
  and g27361 (n16615, n_11092, n16614);
  not g27362 (n_11097, n16613);
  not g27363 (n_11098, n16615);
  and g27364 (n16616, n_11097, n_11098);
  not g27365 (n_11099, n16606);
  not g27366 (n_11100, n16616);
  and g27367 (n16617, n_11099, n_11100);
  not g27368 (n_11101, n16617);
  and g27369 (n16618, \asqrt[24] , n_11101);
  and g27373 (n16622, n_10675, n_10674);
  and g27374 (n16623, \asqrt[12] , n16622);
  not g27375 (n_11102, n16623);
  and g27376 (n16624, n_10673, n_11102);
  not g27377 (n_11103, n16621);
  not g27378 (n_11104, n16624);
  and g27379 (n16625, n_11103, n_11104);
  and g27380 (n16626, n_7218, n_11099);
  and g27381 (n16627, n_11100, n16626);
  not g27382 (n_11105, n16625);
  not g27383 (n_11106, n16627);
  and g27384 (n16628, n_11105, n_11106);
  not g27385 (n_11107, n16618);
  not g27386 (n_11108, n16628);
  and g27387 (n16629, n_11107, n_11108);
  not g27388 (n_11109, n16629);
  and g27389 (n16630, \asqrt[25] , n_11109);
  and g27393 (n16634, n_10683, n_10682);
  and g27394 (n16635, \asqrt[12] , n16634);
  not g27395 (n_11110, n16635);
  and g27396 (n16636, n_10681, n_11110);
  not g27397 (n_11111, n16633);
  not g27398 (n_11112, n16636);
  and g27399 (n16637, n_11111, n_11112);
  and g27400 (n16638, n_6882, n_11107);
  and g27401 (n16639, n_11108, n16638);
  not g27402 (n_11113, n16637);
  not g27403 (n_11114, n16639);
  and g27404 (n16640, n_11113, n_11114);
  not g27405 (n_11115, n16630);
  not g27406 (n_11116, n16640);
  and g27407 (n16641, n_11115, n_11116);
  not g27408 (n_11117, n16641);
  and g27409 (n16642, \asqrt[26] , n_11117);
  and g27413 (n16646, n_10691, n_10690);
  and g27414 (n16647, \asqrt[12] , n16646);
  not g27415 (n_11118, n16647);
  and g27416 (n16648, n_10689, n_11118);
  not g27417 (n_11119, n16645);
  not g27418 (n_11120, n16648);
  and g27419 (n16649, n_11119, n_11120);
  and g27420 (n16650, n_6554, n_11115);
  and g27421 (n16651, n_11116, n16650);
  not g27422 (n_11121, n16649);
  not g27423 (n_11122, n16651);
  and g27424 (n16652, n_11121, n_11122);
  not g27425 (n_11123, n16642);
  not g27426 (n_11124, n16652);
  and g27427 (n16653, n_11123, n_11124);
  not g27428 (n_11125, n16653);
  and g27429 (n16654, \asqrt[27] , n_11125);
  and g27433 (n16658, n_10699, n_10698);
  and g27434 (n16659, \asqrt[12] , n16658);
  not g27435 (n_11126, n16659);
  and g27436 (n16660, n_10697, n_11126);
  not g27437 (n_11127, n16657);
  not g27438 (n_11128, n16660);
  and g27439 (n16661, n_11127, n_11128);
  and g27440 (n16662, n_6234, n_11123);
  and g27441 (n16663, n_11124, n16662);
  not g27442 (n_11129, n16661);
  not g27443 (n_11130, n16663);
  and g27444 (n16664, n_11129, n_11130);
  not g27445 (n_11131, n16654);
  not g27446 (n_11132, n16664);
  and g27447 (n16665, n_11131, n_11132);
  not g27448 (n_11133, n16665);
  and g27449 (n16666, \asqrt[28] , n_11133);
  and g27453 (n16670, n_10707, n_10706);
  and g27454 (n16671, \asqrt[12] , n16670);
  not g27455 (n_11134, n16671);
  and g27456 (n16672, n_10705, n_11134);
  not g27457 (n_11135, n16669);
  not g27458 (n_11136, n16672);
  and g27459 (n16673, n_11135, n_11136);
  and g27460 (n16674, n_5922, n_11131);
  and g27461 (n16675, n_11132, n16674);
  not g27462 (n_11137, n16673);
  not g27463 (n_11138, n16675);
  and g27464 (n16676, n_11137, n_11138);
  not g27465 (n_11139, n16666);
  not g27466 (n_11140, n16676);
  and g27467 (n16677, n_11139, n_11140);
  not g27468 (n_11141, n16677);
  and g27469 (n16678, \asqrt[29] , n_11141);
  and g27473 (n16682, n_10715, n_10714);
  and g27474 (n16683, \asqrt[12] , n16682);
  not g27475 (n_11142, n16683);
  and g27476 (n16684, n_10713, n_11142);
  not g27477 (n_11143, n16681);
  not g27478 (n_11144, n16684);
  and g27479 (n16685, n_11143, n_11144);
  and g27480 (n16686, n_5618, n_11139);
  and g27481 (n16687, n_11140, n16686);
  not g27482 (n_11145, n16685);
  not g27483 (n_11146, n16687);
  and g27484 (n16688, n_11145, n_11146);
  not g27485 (n_11147, n16678);
  not g27486 (n_11148, n16688);
  and g27487 (n16689, n_11147, n_11148);
  not g27488 (n_11149, n16689);
  and g27489 (n16690, \asqrt[30] , n_11149);
  and g27493 (n16694, n_10723, n_10722);
  and g27494 (n16695, \asqrt[12] , n16694);
  not g27495 (n_11150, n16695);
  and g27496 (n16696, n_10721, n_11150);
  not g27497 (n_11151, n16693);
  not g27498 (n_11152, n16696);
  and g27499 (n16697, n_11151, n_11152);
  and g27500 (n16698, n_5322, n_11147);
  and g27501 (n16699, n_11148, n16698);
  not g27502 (n_11153, n16697);
  not g27503 (n_11154, n16699);
  and g27504 (n16700, n_11153, n_11154);
  not g27505 (n_11155, n16690);
  not g27506 (n_11156, n16700);
  and g27507 (n16701, n_11155, n_11156);
  not g27508 (n_11157, n16701);
  and g27509 (n16702, \asqrt[31] , n_11157);
  and g27513 (n16706, n_10731, n_10730);
  and g27514 (n16707, \asqrt[12] , n16706);
  not g27515 (n_11158, n16707);
  and g27516 (n16708, n_10729, n_11158);
  not g27517 (n_11159, n16705);
  not g27518 (n_11160, n16708);
  and g27519 (n16709, n_11159, n_11160);
  and g27520 (n16710, n_5034, n_11155);
  and g27521 (n16711, n_11156, n16710);
  not g27522 (n_11161, n16709);
  not g27523 (n_11162, n16711);
  and g27524 (n16712, n_11161, n_11162);
  not g27525 (n_11163, n16702);
  not g27526 (n_11164, n16712);
  and g27527 (n16713, n_11163, n_11164);
  not g27528 (n_11165, n16713);
  and g27529 (n16714, \asqrt[32] , n_11165);
  and g27533 (n16718, n_10739, n_10738);
  and g27534 (n16719, \asqrt[12] , n16718);
  not g27535 (n_11166, n16719);
  and g27536 (n16720, n_10737, n_11166);
  not g27537 (n_11167, n16717);
  not g27538 (n_11168, n16720);
  and g27539 (n16721, n_11167, n_11168);
  and g27540 (n16722, n_4754, n_11163);
  and g27541 (n16723, n_11164, n16722);
  not g27542 (n_11169, n16721);
  not g27543 (n_11170, n16723);
  and g27544 (n16724, n_11169, n_11170);
  not g27545 (n_11171, n16714);
  not g27546 (n_11172, n16724);
  and g27547 (n16725, n_11171, n_11172);
  not g27548 (n_11173, n16725);
  and g27549 (n16726, \asqrt[33] , n_11173);
  and g27553 (n16730, n_10747, n_10746);
  and g27554 (n16731, \asqrt[12] , n16730);
  not g27555 (n_11174, n16731);
  and g27556 (n16732, n_10745, n_11174);
  not g27557 (n_11175, n16729);
  not g27558 (n_11176, n16732);
  and g27559 (n16733, n_11175, n_11176);
  and g27560 (n16734, n_4482, n_11171);
  and g27561 (n16735, n_11172, n16734);
  not g27562 (n_11177, n16733);
  not g27563 (n_11178, n16735);
  and g27564 (n16736, n_11177, n_11178);
  not g27565 (n_11179, n16726);
  not g27566 (n_11180, n16736);
  and g27567 (n16737, n_11179, n_11180);
  not g27568 (n_11181, n16737);
  and g27569 (n16738, \asqrt[34] , n_11181);
  and g27573 (n16742, n_10755, n_10754);
  and g27574 (n16743, \asqrt[12] , n16742);
  not g27575 (n_11182, n16743);
  and g27576 (n16744, n_10753, n_11182);
  not g27577 (n_11183, n16741);
  not g27578 (n_11184, n16744);
  and g27579 (n16745, n_11183, n_11184);
  and g27580 (n16746, n_4218, n_11179);
  and g27581 (n16747, n_11180, n16746);
  not g27582 (n_11185, n16745);
  not g27583 (n_11186, n16747);
  and g27584 (n16748, n_11185, n_11186);
  not g27585 (n_11187, n16738);
  not g27586 (n_11188, n16748);
  and g27587 (n16749, n_11187, n_11188);
  not g27588 (n_11189, n16749);
  and g27589 (n16750, \asqrt[35] , n_11189);
  and g27593 (n16754, n_10763, n_10762);
  and g27594 (n16755, \asqrt[12] , n16754);
  not g27595 (n_11190, n16755);
  and g27596 (n16756, n_10761, n_11190);
  not g27597 (n_11191, n16753);
  not g27598 (n_11192, n16756);
  and g27599 (n16757, n_11191, n_11192);
  and g27600 (n16758, n_3962, n_11187);
  and g27601 (n16759, n_11188, n16758);
  not g27602 (n_11193, n16757);
  not g27603 (n_11194, n16759);
  and g27604 (n16760, n_11193, n_11194);
  not g27605 (n_11195, n16750);
  not g27606 (n_11196, n16760);
  and g27607 (n16761, n_11195, n_11196);
  not g27608 (n_11197, n16761);
  and g27609 (n16762, \asqrt[36] , n_11197);
  and g27613 (n16766, n_10771, n_10770);
  and g27614 (n16767, \asqrt[12] , n16766);
  not g27615 (n_11198, n16767);
  and g27616 (n16768, n_10769, n_11198);
  not g27617 (n_11199, n16765);
  not g27618 (n_11200, n16768);
  and g27619 (n16769, n_11199, n_11200);
  and g27620 (n16770, n_3714, n_11195);
  and g27621 (n16771, n_11196, n16770);
  not g27622 (n_11201, n16769);
  not g27623 (n_11202, n16771);
  and g27624 (n16772, n_11201, n_11202);
  not g27625 (n_11203, n16762);
  not g27626 (n_11204, n16772);
  and g27627 (n16773, n_11203, n_11204);
  not g27628 (n_11205, n16773);
  and g27629 (n16774, \asqrt[37] , n_11205);
  and g27633 (n16778, n_10779, n_10778);
  and g27634 (n16779, \asqrt[12] , n16778);
  not g27635 (n_11206, n16779);
  and g27636 (n16780, n_10777, n_11206);
  not g27637 (n_11207, n16777);
  not g27638 (n_11208, n16780);
  and g27639 (n16781, n_11207, n_11208);
  and g27640 (n16782, n_3474, n_11203);
  and g27641 (n16783, n_11204, n16782);
  not g27642 (n_11209, n16781);
  not g27643 (n_11210, n16783);
  and g27644 (n16784, n_11209, n_11210);
  not g27645 (n_11211, n16774);
  not g27646 (n_11212, n16784);
  and g27647 (n16785, n_11211, n_11212);
  not g27648 (n_11213, n16785);
  and g27649 (n16786, \asqrt[38] , n_11213);
  and g27653 (n16790, n_10787, n_10786);
  and g27654 (n16791, \asqrt[12] , n16790);
  not g27655 (n_11214, n16791);
  and g27656 (n16792, n_10785, n_11214);
  not g27657 (n_11215, n16789);
  not g27658 (n_11216, n16792);
  and g27659 (n16793, n_11215, n_11216);
  and g27660 (n16794, n_3242, n_11211);
  and g27661 (n16795, n_11212, n16794);
  not g27662 (n_11217, n16793);
  not g27663 (n_11218, n16795);
  and g27664 (n16796, n_11217, n_11218);
  not g27665 (n_11219, n16786);
  not g27666 (n_11220, n16796);
  and g27667 (n16797, n_11219, n_11220);
  not g27668 (n_11221, n16797);
  and g27669 (n16798, \asqrt[39] , n_11221);
  and g27673 (n16802, n_10795, n_10794);
  and g27674 (n16803, \asqrt[12] , n16802);
  not g27675 (n_11222, n16803);
  and g27676 (n16804, n_10793, n_11222);
  not g27677 (n_11223, n16801);
  not g27678 (n_11224, n16804);
  and g27679 (n16805, n_11223, n_11224);
  and g27680 (n16806, n_3018, n_11219);
  and g27681 (n16807, n_11220, n16806);
  not g27682 (n_11225, n16805);
  not g27683 (n_11226, n16807);
  and g27684 (n16808, n_11225, n_11226);
  not g27685 (n_11227, n16798);
  not g27686 (n_11228, n16808);
  and g27687 (n16809, n_11227, n_11228);
  not g27688 (n_11229, n16809);
  and g27689 (n16810, \asqrt[40] , n_11229);
  and g27693 (n16814, n_10803, n_10802);
  and g27694 (n16815, \asqrt[12] , n16814);
  not g27695 (n_11230, n16815);
  and g27696 (n16816, n_10801, n_11230);
  not g27697 (n_11231, n16813);
  not g27698 (n_11232, n16816);
  and g27699 (n16817, n_11231, n_11232);
  and g27700 (n16818, n_2802, n_11227);
  and g27701 (n16819, n_11228, n16818);
  not g27702 (n_11233, n16817);
  not g27703 (n_11234, n16819);
  and g27704 (n16820, n_11233, n_11234);
  not g27705 (n_11235, n16810);
  not g27706 (n_11236, n16820);
  and g27707 (n16821, n_11235, n_11236);
  not g27708 (n_11237, n16821);
  and g27709 (n16822, \asqrt[41] , n_11237);
  and g27713 (n16826, n_10811, n_10810);
  and g27714 (n16827, \asqrt[12] , n16826);
  not g27715 (n_11238, n16827);
  and g27716 (n16828, n_10809, n_11238);
  not g27717 (n_11239, n16825);
  not g27718 (n_11240, n16828);
  and g27719 (n16829, n_11239, n_11240);
  and g27720 (n16830, n_2594, n_11235);
  and g27721 (n16831, n_11236, n16830);
  not g27722 (n_11241, n16829);
  not g27723 (n_11242, n16831);
  and g27724 (n16832, n_11241, n_11242);
  not g27725 (n_11243, n16822);
  not g27726 (n_11244, n16832);
  and g27727 (n16833, n_11243, n_11244);
  not g27728 (n_11245, n16833);
  and g27729 (n16834, \asqrt[42] , n_11245);
  and g27733 (n16838, n_10819, n_10818);
  and g27734 (n16839, \asqrt[12] , n16838);
  not g27735 (n_11246, n16839);
  and g27736 (n16840, n_10817, n_11246);
  not g27737 (n_11247, n16837);
  not g27738 (n_11248, n16840);
  and g27739 (n16841, n_11247, n_11248);
  and g27740 (n16842, n_2394, n_11243);
  and g27741 (n16843, n_11244, n16842);
  not g27742 (n_11249, n16841);
  not g27743 (n_11250, n16843);
  and g27744 (n16844, n_11249, n_11250);
  not g27745 (n_11251, n16834);
  not g27746 (n_11252, n16844);
  and g27747 (n16845, n_11251, n_11252);
  not g27748 (n_11253, n16845);
  and g27749 (n16846, \asqrt[43] , n_11253);
  and g27753 (n16850, n_10827, n_10826);
  and g27754 (n16851, \asqrt[12] , n16850);
  not g27755 (n_11254, n16851);
  and g27756 (n16852, n_10825, n_11254);
  not g27757 (n_11255, n16849);
  not g27758 (n_11256, n16852);
  and g27759 (n16853, n_11255, n_11256);
  and g27760 (n16854, n_2202, n_11251);
  and g27761 (n16855, n_11252, n16854);
  not g27762 (n_11257, n16853);
  not g27763 (n_11258, n16855);
  and g27764 (n16856, n_11257, n_11258);
  not g27765 (n_11259, n16846);
  not g27766 (n_11260, n16856);
  and g27767 (n16857, n_11259, n_11260);
  not g27768 (n_11261, n16857);
  and g27769 (n16858, \asqrt[44] , n_11261);
  and g27773 (n16862, n_10835, n_10834);
  and g27774 (n16863, \asqrt[12] , n16862);
  not g27775 (n_11262, n16863);
  and g27776 (n16864, n_10833, n_11262);
  not g27777 (n_11263, n16861);
  not g27778 (n_11264, n16864);
  and g27779 (n16865, n_11263, n_11264);
  and g27780 (n16866, n_2018, n_11259);
  and g27781 (n16867, n_11260, n16866);
  not g27782 (n_11265, n16865);
  not g27783 (n_11266, n16867);
  and g27784 (n16868, n_11265, n_11266);
  not g27785 (n_11267, n16858);
  not g27786 (n_11268, n16868);
  and g27787 (n16869, n_11267, n_11268);
  not g27788 (n_11269, n16869);
  and g27789 (n16870, \asqrt[45] , n_11269);
  and g27793 (n16874, n_10843, n_10842);
  and g27794 (n16875, \asqrt[12] , n16874);
  not g27795 (n_11270, n16875);
  and g27796 (n16876, n_10841, n_11270);
  not g27797 (n_11271, n16873);
  not g27798 (n_11272, n16876);
  and g27799 (n16877, n_11271, n_11272);
  and g27800 (n16878, n_1842, n_11267);
  and g27801 (n16879, n_11268, n16878);
  not g27802 (n_11273, n16877);
  not g27803 (n_11274, n16879);
  and g27804 (n16880, n_11273, n_11274);
  not g27805 (n_11275, n16870);
  not g27806 (n_11276, n16880);
  and g27807 (n16881, n_11275, n_11276);
  not g27808 (n_11277, n16881);
  and g27809 (n16882, \asqrt[46] , n_11277);
  and g27813 (n16886, n_10851, n_10850);
  and g27814 (n16887, \asqrt[12] , n16886);
  not g27815 (n_11278, n16887);
  and g27816 (n16888, n_10849, n_11278);
  not g27817 (n_11279, n16885);
  not g27818 (n_11280, n16888);
  and g27819 (n16889, n_11279, n_11280);
  and g27820 (n16890, n_1674, n_11275);
  and g27821 (n16891, n_11276, n16890);
  not g27822 (n_11281, n16889);
  not g27823 (n_11282, n16891);
  and g27824 (n16892, n_11281, n_11282);
  not g27825 (n_11283, n16882);
  not g27826 (n_11284, n16892);
  and g27827 (n16893, n_11283, n_11284);
  not g27828 (n_11285, n16893);
  and g27829 (n16894, \asqrt[47] , n_11285);
  and g27833 (n16898, n_10859, n_10858);
  and g27834 (n16899, \asqrt[12] , n16898);
  not g27835 (n_11286, n16899);
  and g27836 (n16900, n_10857, n_11286);
  not g27837 (n_11287, n16897);
  not g27838 (n_11288, n16900);
  and g27839 (n16901, n_11287, n_11288);
  and g27840 (n16902, n_1514, n_11283);
  and g27841 (n16903, n_11284, n16902);
  not g27842 (n_11289, n16901);
  not g27843 (n_11290, n16903);
  and g27844 (n16904, n_11289, n_11290);
  not g27845 (n_11291, n16894);
  not g27846 (n_11292, n16904);
  and g27847 (n16905, n_11291, n_11292);
  not g27848 (n_11293, n16905);
  and g27849 (n16906, \asqrt[48] , n_11293);
  and g27853 (n16910, n_10867, n_10866);
  and g27854 (n16911, \asqrt[12] , n16910);
  not g27855 (n_11294, n16911);
  and g27856 (n16912, n_10865, n_11294);
  not g27857 (n_11295, n16909);
  not g27858 (n_11296, n16912);
  and g27859 (n16913, n_11295, n_11296);
  and g27860 (n16914, n_1362, n_11291);
  and g27861 (n16915, n_11292, n16914);
  not g27862 (n_11297, n16913);
  not g27863 (n_11298, n16915);
  and g27864 (n16916, n_11297, n_11298);
  not g27865 (n_11299, n16906);
  not g27866 (n_11300, n16916);
  and g27867 (n16917, n_11299, n_11300);
  not g27868 (n_11301, n16917);
  and g27869 (n16918, \asqrt[49] , n_11301);
  and g27873 (n16922, n_10875, n_10874);
  and g27874 (n16923, \asqrt[12] , n16922);
  not g27875 (n_11302, n16923);
  and g27876 (n16924, n_10873, n_11302);
  not g27877 (n_11303, n16921);
  not g27878 (n_11304, n16924);
  and g27879 (n16925, n_11303, n_11304);
  and g27880 (n16926, n_1218, n_11299);
  and g27881 (n16927, n_11300, n16926);
  not g27882 (n_11305, n16925);
  not g27883 (n_11306, n16927);
  and g27884 (n16928, n_11305, n_11306);
  not g27885 (n_11307, n16918);
  not g27886 (n_11308, n16928);
  and g27887 (n16929, n_11307, n_11308);
  not g27888 (n_11309, n16929);
  and g27889 (n16930, \asqrt[50] , n_11309);
  and g27893 (n16934, n_10883, n_10882);
  and g27894 (n16935, \asqrt[12] , n16934);
  not g27895 (n_11310, n16935);
  and g27896 (n16936, n_10881, n_11310);
  not g27897 (n_11311, n16933);
  not g27898 (n_11312, n16936);
  and g27899 (n16937, n_11311, n_11312);
  and g27900 (n16938, n_1082, n_11307);
  and g27901 (n16939, n_11308, n16938);
  not g27902 (n_11313, n16937);
  not g27903 (n_11314, n16939);
  and g27904 (n16940, n_11313, n_11314);
  not g27905 (n_11315, n16930);
  not g27906 (n_11316, n16940);
  and g27907 (n16941, n_11315, n_11316);
  not g27908 (n_11317, n16941);
  and g27909 (n16942, \asqrt[51] , n_11317);
  and g27913 (n16946, n_10891, n_10890);
  and g27914 (n16947, \asqrt[12] , n16946);
  not g27915 (n_11318, n16947);
  and g27916 (n16948, n_10889, n_11318);
  not g27917 (n_11319, n16945);
  not g27918 (n_11320, n16948);
  and g27919 (n16949, n_11319, n_11320);
  and g27920 (n16950, n_954, n_11315);
  and g27921 (n16951, n_11316, n16950);
  not g27922 (n_11321, n16949);
  not g27923 (n_11322, n16951);
  and g27924 (n16952, n_11321, n_11322);
  not g27925 (n_11323, n16942);
  not g27926 (n_11324, n16952);
  and g27927 (n16953, n_11323, n_11324);
  not g27928 (n_11325, n16953);
  and g27929 (n16954, \asqrt[52] , n_11325);
  and g27933 (n16958, n_10899, n_10898);
  and g27934 (n16959, \asqrt[12] , n16958);
  not g27935 (n_11326, n16959);
  and g27936 (n16960, n_10897, n_11326);
  not g27937 (n_11327, n16957);
  not g27938 (n_11328, n16960);
  and g27939 (n16961, n_11327, n_11328);
  and g27940 (n16962, n_834, n_11323);
  and g27941 (n16963, n_11324, n16962);
  not g27942 (n_11329, n16961);
  not g27943 (n_11330, n16963);
  and g27944 (n16964, n_11329, n_11330);
  not g27945 (n_11331, n16954);
  not g27946 (n_11332, n16964);
  and g27947 (n16965, n_11331, n_11332);
  not g27948 (n_11333, n16965);
  and g27949 (n16966, \asqrt[53] , n_11333);
  and g27950 (n16967, n_722, n_11331);
  and g27951 (n16968, n_11332, n16967);
  and g27955 (n16972, n_10907, n_10905);
  and g27956 (n16973, \asqrt[12] , n16972);
  not g27957 (n_11334, n16973);
  and g27958 (n16974, n_10906, n_11334);
  not g27959 (n_11335, n16971);
  not g27960 (n_11336, n16974);
  and g27961 (n16975, n_11335, n_11336);
  not g27962 (n_11337, n16968);
  not g27963 (n_11338, n16975);
  and g27964 (n16976, n_11337, n_11338);
  not g27965 (n_11339, n16966);
  not g27966 (n_11340, n16976);
  and g27967 (n16977, n_11339, n_11340);
  not g27968 (n_11341, n16977);
  and g27969 (n16978, \asqrt[54] , n_11341);
  and g27973 (n16982, n_10915, n_10914);
  and g27974 (n16983, \asqrt[12] , n16982);
  not g27975 (n_11342, n16983);
  and g27976 (n16984, n_10913, n_11342);
  not g27977 (n_11343, n16981);
  not g27978 (n_11344, n16984);
  and g27979 (n16985, n_11343, n_11344);
  and g27980 (n16986, n_618, n_11339);
  and g27981 (n16987, n_11340, n16986);
  not g27982 (n_11345, n16985);
  not g27983 (n_11346, n16987);
  and g27984 (n16988, n_11345, n_11346);
  not g27985 (n_11347, n16978);
  not g27986 (n_11348, n16988);
  and g27987 (n16989, n_11347, n_11348);
  not g27988 (n_11349, n16989);
  and g27989 (n16990, \asqrt[55] , n_11349);
  and g27993 (n16994, n_10923, n_10922);
  and g27994 (n16995, \asqrt[12] , n16994);
  not g27995 (n_11350, n16995);
  and g27996 (n16996, n_10921, n_11350);
  not g27997 (n_11351, n16993);
  not g27998 (n_11352, n16996);
  and g27999 (n16997, n_11351, n_11352);
  and g28000 (n16998, n_522, n_11347);
  and g28001 (n16999, n_11348, n16998);
  not g28002 (n_11353, n16997);
  not g28003 (n_11354, n16999);
  and g28004 (n17000, n_11353, n_11354);
  not g28005 (n_11355, n16990);
  not g28006 (n_11356, n17000);
  and g28007 (n17001, n_11355, n_11356);
  not g28008 (n_11357, n17001);
  and g28009 (n17002, \asqrt[56] , n_11357);
  and g28013 (n17006, n_10931, n_10930);
  and g28014 (n17007, \asqrt[12] , n17006);
  not g28015 (n_11358, n17007);
  and g28016 (n17008, n_10929, n_11358);
  not g28017 (n_11359, n17005);
  not g28018 (n_11360, n17008);
  and g28019 (n17009, n_11359, n_11360);
  and g28020 (n17010, n_434, n_11355);
  and g28021 (n17011, n_11356, n17010);
  not g28022 (n_11361, n17009);
  not g28023 (n_11362, n17011);
  and g28024 (n17012, n_11361, n_11362);
  not g28025 (n_11363, n17002);
  not g28026 (n_11364, n17012);
  and g28027 (n17013, n_11363, n_11364);
  not g28028 (n_11365, n17013);
  and g28029 (n17014, \asqrt[57] , n_11365);
  and g28033 (n17018, n_10939, n_10938);
  and g28034 (n17019, \asqrt[12] , n17018);
  not g28035 (n_11366, n17019);
  and g28036 (n17020, n_10937, n_11366);
  not g28037 (n_11367, n17017);
  not g28038 (n_11368, n17020);
  and g28039 (n17021, n_11367, n_11368);
  and g28040 (n17022, n_354, n_11363);
  and g28041 (n17023, n_11364, n17022);
  not g28042 (n_11369, n17021);
  not g28043 (n_11370, n17023);
  and g28044 (n17024, n_11369, n_11370);
  not g28045 (n_11371, n17014);
  not g28046 (n_11372, n17024);
  and g28047 (n17025, n_11371, n_11372);
  not g28048 (n_11373, n17025);
  and g28049 (n17026, \asqrt[58] , n_11373);
  and g28053 (n17030, n_10947, n_10946);
  and g28054 (n17031, \asqrt[12] , n17030);
  not g28055 (n_11374, n17031);
  and g28056 (n17032, n_10945, n_11374);
  not g28057 (n_11375, n17029);
  not g28058 (n_11376, n17032);
  and g28059 (n17033, n_11375, n_11376);
  and g28060 (n17034, n_282, n_11371);
  and g28061 (n17035, n_11372, n17034);
  not g28062 (n_11377, n17033);
  not g28063 (n_11378, n17035);
  and g28064 (n17036, n_11377, n_11378);
  not g28065 (n_11379, n17026);
  not g28066 (n_11380, n17036);
  and g28067 (n17037, n_11379, n_11380);
  not g28068 (n_11381, n17037);
  and g28069 (n17038, \asqrt[59] , n_11381);
  and g28073 (n17042, n_10955, n_10954);
  and g28074 (n17043, \asqrt[12] , n17042);
  not g28075 (n_11382, n17043);
  and g28076 (n17044, n_10953, n_11382);
  not g28077 (n_11383, n17041);
  not g28078 (n_11384, n17044);
  and g28079 (n17045, n_11383, n_11384);
  and g28080 (n17046, n_218, n_11379);
  and g28081 (n17047, n_11380, n17046);
  not g28082 (n_11385, n17045);
  not g28083 (n_11386, n17047);
  and g28084 (n17048, n_11385, n_11386);
  not g28085 (n_11387, n17038);
  not g28086 (n_11388, n17048);
  and g28087 (n17049, n_11387, n_11388);
  not g28088 (n_11389, n17049);
  and g28089 (n17050, \asqrt[60] , n_11389);
  and g28093 (n17054, n_10963, n_10962);
  and g28094 (n17055, \asqrt[12] , n17054);
  not g28095 (n_11390, n17055);
  and g28096 (n17056, n_10961, n_11390);
  not g28097 (n_11391, n17053);
  not g28098 (n_11392, n17056);
  and g28099 (n17057, n_11391, n_11392);
  and g28100 (n17058, n_162, n_11387);
  and g28101 (n17059, n_11388, n17058);
  not g28102 (n_11393, n17057);
  not g28103 (n_11394, n17059);
  and g28104 (n17060, n_11393, n_11394);
  not g28105 (n_11395, n17050);
  not g28106 (n_11396, n17060);
  and g28107 (n17061, n_11395, n_11396);
  not g28108 (n_11397, n17061);
  and g28109 (n17062, \asqrt[61] , n_11397);
  and g28113 (n17066, n_10971, n_10970);
  and g28114 (n17067, \asqrt[12] , n17066);
  not g28115 (n_11398, n17067);
  and g28116 (n17068, n_10969, n_11398);
  not g28117 (n_11399, n17065);
  not g28118 (n_11400, n17068);
  and g28119 (n17069, n_11399, n_11400);
  and g28120 (n17070, n_115, n_11395);
  and g28121 (n17071, n_11396, n17070);
  not g28122 (n_11401, n17069);
  not g28123 (n_11402, n17071);
  and g28124 (n17072, n_11401, n_11402);
  not g28125 (n_11403, n17062);
  not g28126 (n_11404, n17072);
  and g28127 (n17073, n_11403, n_11404);
  not g28128 (n_11405, n17073);
  and g28129 (n17074, \asqrt[62] , n_11405);
  and g28133 (n17078, n_10979, n_10978);
  and g28134 (n17079, \asqrt[12] , n17078);
  not g28135 (n_11406, n17079);
  and g28136 (n17080, n_10977, n_11406);
  not g28137 (n_11407, n17077);
  not g28138 (n_11408, n17080);
  and g28139 (n17081, n_11407, n_11408);
  and g28140 (n17082, n_76, n_11403);
  and g28141 (n17083, n_11404, n17082);
  not g28142 (n_11409, n17081);
  not g28143 (n_11410, n17083);
  and g28144 (n17084, n_11409, n_11410);
  not g28145 (n_11411, n17074);
  not g28146 (n_11412, n17084);
  and g28147 (n17085, n_11411, n_11412);
  and g28151 (n17089, n_10987, n_10986);
  and g28152 (n17090, \asqrt[12] , n17089);
  not g28153 (n_11413, n17090);
  and g28154 (n17091, n_10985, n_11413);
  not g28155 (n_11414, n17088);
  not g28156 (n_11415, n17091);
  and g28157 (n17092, n_11414, n_11415);
  and g28158 (n17093, n_10994, n_10993);
  and g28159 (n17094, \asqrt[12] , n17093);
  not g28162 (n_11417, n17092);
  not g28164 (n_11418, n17085);
  not g28166 (n_11419, n17097);
  and g28167 (n17098, n_21, n_11419);
  and g28168 (n17099, n_11411, n17092);
  and g28169 (n17100, n_11412, n17099);
  and g28170 (n17101, n_10993, \asqrt[12] );
  not g28171 (n_11420, n17101);
  and g28172 (n17102, n16453, n_11420);
  not g28173 (n_11421, n17093);
  and g28174 (n17103, \asqrt[63] , n_11421);
  not g28175 (n_11422, n17102);
  and g28176 (n17104, n_11422, n17103);
  not g28182 (n_11423, n17104);
  not g28183 (n_11424, n17109);
  not g28185 (n_11425, n17100);
  and g28189 (n17113, \a[22] , \asqrt[11] );
  not g28190 (n_11430, \a[20] );
  not g28191 (n_11431, \a[21] );
  and g28192 (n17114, n_11430, n_11431);
  and g28193 (n17115, n_11006, n17114);
  not g28194 (n_11432, n17113);
  not g28195 (n_11433, n17115);
  and g28196 (n17116, n_11432, n_11433);
  not g28197 (n_11434, n17116);
  and g28198 (n17117, \asqrt[12] , n_11434);
  and g28204 (n17123, n_11006, \asqrt[11] );
  not g28205 (n_11435, n17123);
  and g28206 (n17124, \a[23] , n_11435);
  and g28207 (n17125, n16482, \asqrt[11] );
  not g28208 (n_11436, n17124);
  not g28209 (n_11437, n17125);
  and g28210 (n17126, n_11436, n_11437);
  not g28211 (n_11438, n17122);
  and g28212 (n17127, n_11438, n17126);
  not g28213 (n_11439, n17117);
  not g28214 (n_11440, n17127);
  and g28215 (n17128, n_11439, n_11440);
  not g28216 (n_11441, n17128);
  and g28217 (n17129, \asqrt[13] , n_11441);
  not g28218 (n_11442, \asqrt[13] );
  and g28219 (n17130, n_11442, n_11439);
  and g28220 (n17131, n_11440, n17130);
  not g28224 (n_11443, n17098);
  not g28226 (n_11444, n17135);
  and g28227 (n17136, n_11437, n_11444);
  not g28228 (n_11445, n17136);
  and g28229 (n17137, \a[24] , n_11445);
  and g28230 (n17138, n_10590, n_11444);
  and g28231 (n17139, n_11437, n17138);
  not g28232 (n_11446, n17137);
  not g28233 (n_11447, n17139);
  and g28234 (n17140, n_11446, n_11447);
  not g28235 (n_11448, n17131);
  not g28236 (n_11449, n17140);
  and g28237 (n17141, n_11448, n_11449);
  not g28238 (n_11450, n17129);
  not g28239 (n_11451, n17141);
  and g28240 (n17142, n_11450, n_11451);
  not g28241 (n_11452, n17142);
  and g28242 (n17143, \asqrt[14] , n_11452);
  and g28243 (n17144, n_11015, n_11014);
  not g28244 (n_11453, n16494);
  and g28245 (n17145, n_11453, n17144);
  and g28246 (n17146, \asqrt[11] , n17145);
  and g28247 (n17147, \asqrt[11] , n17144);
  not g28248 (n_11454, n17147);
  and g28249 (n17148, n16494, n_11454);
  not g28250 (n_11455, n17146);
  not g28251 (n_11456, n17148);
  and g28252 (n17149, n_11455, n_11456);
  and g28253 (n17150, n_11018, n_11450);
  and g28254 (n17151, n_11451, n17150);
  not g28255 (n_11457, n17149);
  not g28256 (n_11458, n17151);
  and g28257 (n17152, n_11457, n_11458);
  not g28258 (n_11459, n17143);
  not g28259 (n_11460, n17152);
  and g28260 (n17153, n_11459, n_11460);
  not g28261 (n_11461, n17153);
  and g28262 (n17154, \asqrt[15] , n_11461);
  and g28266 (n17158, n_11026, n_11024);
  and g28267 (n17159, \asqrt[11] , n17158);
  not g28268 (n_11462, n17159);
  and g28269 (n17160, n_11025, n_11462);
  not g28270 (n_11463, n17157);
  not g28271 (n_11464, n17160);
  and g28272 (n17161, n_11463, n_11464);
  and g28273 (n17162, n_10602, n_11459);
  and g28274 (n17163, n_11460, n17162);
  not g28275 (n_11465, n17161);
  not g28276 (n_11466, n17163);
  and g28277 (n17164, n_11465, n_11466);
  not g28278 (n_11467, n17154);
  not g28279 (n_11468, n17164);
  and g28280 (n17165, n_11467, n_11468);
  not g28281 (n_11469, n17165);
  and g28282 (n17166, \asqrt[16] , n_11469);
  and g28286 (n17170, n_11035, n_11034);
  and g28287 (n17171, \asqrt[11] , n17170);
  not g28288 (n_11470, n17171);
  and g28289 (n17172, n_11033, n_11470);
  not g28290 (n_11471, n17169);
  not g28291 (n_11472, n17172);
  and g28292 (n17173, n_11471, n_11472);
  and g28293 (n17174, n_10194, n_11467);
  and g28294 (n17175, n_11468, n17174);
  not g28295 (n_11473, n17173);
  not g28296 (n_11474, n17175);
  and g28297 (n17176, n_11473, n_11474);
  not g28298 (n_11475, n17166);
  not g28299 (n_11476, n17176);
  and g28300 (n17177, n_11475, n_11476);
  not g28301 (n_11477, n17177);
  and g28302 (n17178, \asqrt[17] , n_11477);
  and g28306 (n17182, n_11043, n_11042);
  and g28307 (n17183, \asqrt[11] , n17182);
  not g28308 (n_11478, n17183);
  and g28309 (n17184, n_11041, n_11478);
  not g28310 (n_11479, n17181);
  not g28311 (n_11480, n17184);
  and g28312 (n17185, n_11479, n_11480);
  and g28313 (n17186, n_9794, n_11475);
  and g28314 (n17187, n_11476, n17186);
  not g28315 (n_11481, n17185);
  not g28316 (n_11482, n17187);
  and g28317 (n17188, n_11481, n_11482);
  not g28318 (n_11483, n17178);
  not g28319 (n_11484, n17188);
  and g28320 (n17189, n_11483, n_11484);
  not g28321 (n_11485, n17189);
  and g28322 (n17190, \asqrt[18] , n_11485);
  and g28326 (n17194, n_11051, n_11050);
  and g28327 (n17195, \asqrt[11] , n17194);
  not g28328 (n_11486, n17195);
  and g28329 (n17196, n_11049, n_11486);
  not g28330 (n_11487, n17193);
  not g28331 (n_11488, n17196);
  and g28332 (n17197, n_11487, n_11488);
  and g28333 (n17198, n_9402, n_11483);
  and g28334 (n17199, n_11484, n17198);
  not g28335 (n_11489, n17197);
  not g28336 (n_11490, n17199);
  and g28337 (n17200, n_11489, n_11490);
  not g28338 (n_11491, n17190);
  not g28339 (n_11492, n17200);
  and g28340 (n17201, n_11491, n_11492);
  not g28341 (n_11493, n17201);
  and g28342 (n17202, \asqrt[19] , n_11493);
  and g28346 (n17206, n_11059, n_11058);
  and g28347 (n17207, \asqrt[11] , n17206);
  not g28348 (n_11494, n17207);
  and g28349 (n17208, n_11057, n_11494);
  not g28350 (n_11495, n17205);
  not g28351 (n_11496, n17208);
  and g28352 (n17209, n_11495, n_11496);
  and g28353 (n17210, n_9018, n_11491);
  and g28354 (n17211, n_11492, n17210);
  not g28355 (n_11497, n17209);
  not g28356 (n_11498, n17211);
  and g28357 (n17212, n_11497, n_11498);
  not g28358 (n_11499, n17202);
  not g28359 (n_11500, n17212);
  and g28360 (n17213, n_11499, n_11500);
  not g28361 (n_11501, n17213);
  and g28362 (n17214, \asqrt[20] , n_11501);
  and g28366 (n17218, n_11067, n_11066);
  and g28367 (n17219, \asqrt[11] , n17218);
  not g28368 (n_11502, n17219);
  and g28369 (n17220, n_11065, n_11502);
  not g28370 (n_11503, n17217);
  not g28371 (n_11504, n17220);
  and g28372 (n17221, n_11503, n_11504);
  and g28373 (n17222, n_8642, n_11499);
  and g28374 (n17223, n_11500, n17222);
  not g28375 (n_11505, n17221);
  not g28376 (n_11506, n17223);
  and g28377 (n17224, n_11505, n_11506);
  not g28378 (n_11507, n17214);
  not g28379 (n_11508, n17224);
  and g28380 (n17225, n_11507, n_11508);
  not g28381 (n_11509, n17225);
  and g28382 (n17226, \asqrt[21] , n_11509);
  and g28386 (n17230, n_11075, n_11074);
  and g28387 (n17231, \asqrt[11] , n17230);
  not g28388 (n_11510, n17231);
  and g28389 (n17232, n_11073, n_11510);
  not g28390 (n_11511, n17229);
  not g28391 (n_11512, n17232);
  and g28392 (n17233, n_11511, n_11512);
  and g28393 (n17234, n_8274, n_11507);
  and g28394 (n17235, n_11508, n17234);
  not g28395 (n_11513, n17233);
  not g28396 (n_11514, n17235);
  and g28397 (n17236, n_11513, n_11514);
  not g28398 (n_11515, n17226);
  not g28399 (n_11516, n17236);
  and g28400 (n17237, n_11515, n_11516);
  not g28401 (n_11517, n17237);
  and g28402 (n17238, \asqrt[22] , n_11517);
  and g28406 (n17242, n_11083, n_11082);
  and g28407 (n17243, \asqrt[11] , n17242);
  not g28408 (n_11518, n17243);
  and g28409 (n17244, n_11081, n_11518);
  not g28410 (n_11519, n17241);
  not g28411 (n_11520, n17244);
  and g28412 (n17245, n_11519, n_11520);
  and g28413 (n17246, n_7914, n_11515);
  and g28414 (n17247, n_11516, n17246);
  not g28415 (n_11521, n17245);
  not g28416 (n_11522, n17247);
  and g28417 (n17248, n_11521, n_11522);
  not g28418 (n_11523, n17238);
  not g28419 (n_11524, n17248);
  and g28420 (n17249, n_11523, n_11524);
  not g28421 (n_11525, n17249);
  and g28422 (n17250, \asqrt[23] , n_11525);
  and g28426 (n17254, n_11091, n_11090);
  and g28427 (n17255, \asqrt[11] , n17254);
  not g28428 (n_11526, n17255);
  and g28429 (n17256, n_11089, n_11526);
  not g28430 (n_11527, n17253);
  not g28431 (n_11528, n17256);
  and g28432 (n17257, n_11527, n_11528);
  and g28433 (n17258, n_7562, n_11523);
  and g28434 (n17259, n_11524, n17258);
  not g28435 (n_11529, n17257);
  not g28436 (n_11530, n17259);
  and g28437 (n17260, n_11529, n_11530);
  not g28438 (n_11531, n17250);
  not g28439 (n_11532, n17260);
  and g28440 (n17261, n_11531, n_11532);
  not g28441 (n_11533, n17261);
  and g28442 (n17262, \asqrt[24] , n_11533);
  and g28446 (n17266, n_11099, n_11098);
  and g28447 (n17267, \asqrt[11] , n17266);
  not g28448 (n_11534, n17267);
  and g28449 (n17268, n_11097, n_11534);
  not g28450 (n_11535, n17265);
  not g28451 (n_11536, n17268);
  and g28452 (n17269, n_11535, n_11536);
  and g28453 (n17270, n_7218, n_11531);
  and g28454 (n17271, n_11532, n17270);
  not g28455 (n_11537, n17269);
  not g28456 (n_11538, n17271);
  and g28457 (n17272, n_11537, n_11538);
  not g28458 (n_11539, n17262);
  not g28459 (n_11540, n17272);
  and g28460 (n17273, n_11539, n_11540);
  not g28461 (n_11541, n17273);
  and g28462 (n17274, \asqrt[25] , n_11541);
  and g28466 (n17278, n_11107, n_11106);
  and g28467 (n17279, \asqrt[11] , n17278);
  not g28468 (n_11542, n17279);
  and g28469 (n17280, n_11105, n_11542);
  not g28470 (n_11543, n17277);
  not g28471 (n_11544, n17280);
  and g28472 (n17281, n_11543, n_11544);
  and g28473 (n17282, n_6882, n_11539);
  and g28474 (n17283, n_11540, n17282);
  not g28475 (n_11545, n17281);
  not g28476 (n_11546, n17283);
  and g28477 (n17284, n_11545, n_11546);
  not g28478 (n_11547, n17274);
  not g28479 (n_11548, n17284);
  and g28480 (n17285, n_11547, n_11548);
  not g28481 (n_11549, n17285);
  and g28482 (n17286, \asqrt[26] , n_11549);
  and g28486 (n17290, n_11115, n_11114);
  and g28487 (n17291, \asqrt[11] , n17290);
  not g28488 (n_11550, n17291);
  and g28489 (n17292, n_11113, n_11550);
  not g28490 (n_11551, n17289);
  not g28491 (n_11552, n17292);
  and g28492 (n17293, n_11551, n_11552);
  and g28493 (n17294, n_6554, n_11547);
  and g28494 (n17295, n_11548, n17294);
  not g28495 (n_11553, n17293);
  not g28496 (n_11554, n17295);
  and g28497 (n17296, n_11553, n_11554);
  not g28498 (n_11555, n17286);
  not g28499 (n_11556, n17296);
  and g28500 (n17297, n_11555, n_11556);
  not g28501 (n_11557, n17297);
  and g28502 (n17298, \asqrt[27] , n_11557);
  and g28506 (n17302, n_11123, n_11122);
  and g28507 (n17303, \asqrt[11] , n17302);
  not g28508 (n_11558, n17303);
  and g28509 (n17304, n_11121, n_11558);
  not g28510 (n_11559, n17301);
  not g28511 (n_11560, n17304);
  and g28512 (n17305, n_11559, n_11560);
  and g28513 (n17306, n_6234, n_11555);
  and g28514 (n17307, n_11556, n17306);
  not g28515 (n_11561, n17305);
  not g28516 (n_11562, n17307);
  and g28517 (n17308, n_11561, n_11562);
  not g28518 (n_11563, n17298);
  not g28519 (n_11564, n17308);
  and g28520 (n17309, n_11563, n_11564);
  not g28521 (n_11565, n17309);
  and g28522 (n17310, \asqrt[28] , n_11565);
  and g28526 (n17314, n_11131, n_11130);
  and g28527 (n17315, \asqrt[11] , n17314);
  not g28528 (n_11566, n17315);
  and g28529 (n17316, n_11129, n_11566);
  not g28530 (n_11567, n17313);
  not g28531 (n_11568, n17316);
  and g28532 (n17317, n_11567, n_11568);
  and g28533 (n17318, n_5922, n_11563);
  and g28534 (n17319, n_11564, n17318);
  not g28535 (n_11569, n17317);
  not g28536 (n_11570, n17319);
  and g28537 (n17320, n_11569, n_11570);
  not g28538 (n_11571, n17310);
  not g28539 (n_11572, n17320);
  and g28540 (n17321, n_11571, n_11572);
  not g28541 (n_11573, n17321);
  and g28542 (n17322, \asqrt[29] , n_11573);
  and g28546 (n17326, n_11139, n_11138);
  and g28547 (n17327, \asqrt[11] , n17326);
  not g28548 (n_11574, n17327);
  and g28549 (n17328, n_11137, n_11574);
  not g28550 (n_11575, n17325);
  not g28551 (n_11576, n17328);
  and g28552 (n17329, n_11575, n_11576);
  and g28553 (n17330, n_5618, n_11571);
  and g28554 (n17331, n_11572, n17330);
  not g28555 (n_11577, n17329);
  not g28556 (n_11578, n17331);
  and g28557 (n17332, n_11577, n_11578);
  not g28558 (n_11579, n17322);
  not g28559 (n_11580, n17332);
  and g28560 (n17333, n_11579, n_11580);
  not g28561 (n_11581, n17333);
  and g28562 (n17334, \asqrt[30] , n_11581);
  and g28566 (n17338, n_11147, n_11146);
  and g28567 (n17339, \asqrt[11] , n17338);
  not g28568 (n_11582, n17339);
  and g28569 (n17340, n_11145, n_11582);
  not g28570 (n_11583, n17337);
  not g28571 (n_11584, n17340);
  and g28572 (n17341, n_11583, n_11584);
  and g28573 (n17342, n_5322, n_11579);
  and g28574 (n17343, n_11580, n17342);
  not g28575 (n_11585, n17341);
  not g28576 (n_11586, n17343);
  and g28577 (n17344, n_11585, n_11586);
  not g28578 (n_11587, n17334);
  not g28579 (n_11588, n17344);
  and g28580 (n17345, n_11587, n_11588);
  not g28581 (n_11589, n17345);
  and g28582 (n17346, \asqrt[31] , n_11589);
  and g28586 (n17350, n_11155, n_11154);
  and g28587 (n17351, \asqrt[11] , n17350);
  not g28588 (n_11590, n17351);
  and g28589 (n17352, n_11153, n_11590);
  not g28590 (n_11591, n17349);
  not g28591 (n_11592, n17352);
  and g28592 (n17353, n_11591, n_11592);
  and g28593 (n17354, n_5034, n_11587);
  and g28594 (n17355, n_11588, n17354);
  not g28595 (n_11593, n17353);
  not g28596 (n_11594, n17355);
  and g28597 (n17356, n_11593, n_11594);
  not g28598 (n_11595, n17346);
  not g28599 (n_11596, n17356);
  and g28600 (n17357, n_11595, n_11596);
  not g28601 (n_11597, n17357);
  and g28602 (n17358, \asqrt[32] , n_11597);
  and g28606 (n17362, n_11163, n_11162);
  and g28607 (n17363, \asqrt[11] , n17362);
  not g28608 (n_11598, n17363);
  and g28609 (n17364, n_11161, n_11598);
  not g28610 (n_11599, n17361);
  not g28611 (n_11600, n17364);
  and g28612 (n17365, n_11599, n_11600);
  and g28613 (n17366, n_4754, n_11595);
  and g28614 (n17367, n_11596, n17366);
  not g28615 (n_11601, n17365);
  not g28616 (n_11602, n17367);
  and g28617 (n17368, n_11601, n_11602);
  not g28618 (n_11603, n17358);
  not g28619 (n_11604, n17368);
  and g28620 (n17369, n_11603, n_11604);
  not g28621 (n_11605, n17369);
  and g28622 (n17370, \asqrt[33] , n_11605);
  and g28626 (n17374, n_11171, n_11170);
  and g28627 (n17375, \asqrt[11] , n17374);
  not g28628 (n_11606, n17375);
  and g28629 (n17376, n_11169, n_11606);
  not g28630 (n_11607, n17373);
  not g28631 (n_11608, n17376);
  and g28632 (n17377, n_11607, n_11608);
  and g28633 (n17378, n_4482, n_11603);
  and g28634 (n17379, n_11604, n17378);
  not g28635 (n_11609, n17377);
  not g28636 (n_11610, n17379);
  and g28637 (n17380, n_11609, n_11610);
  not g28638 (n_11611, n17370);
  not g28639 (n_11612, n17380);
  and g28640 (n17381, n_11611, n_11612);
  not g28641 (n_11613, n17381);
  and g28642 (n17382, \asqrt[34] , n_11613);
  and g28646 (n17386, n_11179, n_11178);
  and g28647 (n17387, \asqrt[11] , n17386);
  not g28648 (n_11614, n17387);
  and g28649 (n17388, n_11177, n_11614);
  not g28650 (n_11615, n17385);
  not g28651 (n_11616, n17388);
  and g28652 (n17389, n_11615, n_11616);
  and g28653 (n17390, n_4218, n_11611);
  and g28654 (n17391, n_11612, n17390);
  not g28655 (n_11617, n17389);
  not g28656 (n_11618, n17391);
  and g28657 (n17392, n_11617, n_11618);
  not g28658 (n_11619, n17382);
  not g28659 (n_11620, n17392);
  and g28660 (n17393, n_11619, n_11620);
  not g28661 (n_11621, n17393);
  and g28662 (n17394, \asqrt[35] , n_11621);
  and g28666 (n17398, n_11187, n_11186);
  and g28667 (n17399, \asqrt[11] , n17398);
  not g28668 (n_11622, n17399);
  and g28669 (n17400, n_11185, n_11622);
  not g28670 (n_11623, n17397);
  not g28671 (n_11624, n17400);
  and g28672 (n17401, n_11623, n_11624);
  and g28673 (n17402, n_3962, n_11619);
  and g28674 (n17403, n_11620, n17402);
  not g28675 (n_11625, n17401);
  not g28676 (n_11626, n17403);
  and g28677 (n17404, n_11625, n_11626);
  not g28678 (n_11627, n17394);
  not g28679 (n_11628, n17404);
  and g28680 (n17405, n_11627, n_11628);
  not g28681 (n_11629, n17405);
  and g28682 (n17406, \asqrt[36] , n_11629);
  and g28686 (n17410, n_11195, n_11194);
  and g28687 (n17411, \asqrt[11] , n17410);
  not g28688 (n_11630, n17411);
  and g28689 (n17412, n_11193, n_11630);
  not g28690 (n_11631, n17409);
  not g28691 (n_11632, n17412);
  and g28692 (n17413, n_11631, n_11632);
  and g28693 (n17414, n_3714, n_11627);
  and g28694 (n17415, n_11628, n17414);
  not g28695 (n_11633, n17413);
  not g28696 (n_11634, n17415);
  and g28697 (n17416, n_11633, n_11634);
  not g28698 (n_11635, n17406);
  not g28699 (n_11636, n17416);
  and g28700 (n17417, n_11635, n_11636);
  not g28701 (n_11637, n17417);
  and g28702 (n17418, \asqrt[37] , n_11637);
  and g28706 (n17422, n_11203, n_11202);
  and g28707 (n17423, \asqrt[11] , n17422);
  not g28708 (n_11638, n17423);
  and g28709 (n17424, n_11201, n_11638);
  not g28710 (n_11639, n17421);
  not g28711 (n_11640, n17424);
  and g28712 (n17425, n_11639, n_11640);
  and g28713 (n17426, n_3474, n_11635);
  and g28714 (n17427, n_11636, n17426);
  not g28715 (n_11641, n17425);
  not g28716 (n_11642, n17427);
  and g28717 (n17428, n_11641, n_11642);
  not g28718 (n_11643, n17418);
  not g28719 (n_11644, n17428);
  and g28720 (n17429, n_11643, n_11644);
  not g28721 (n_11645, n17429);
  and g28722 (n17430, \asqrt[38] , n_11645);
  and g28726 (n17434, n_11211, n_11210);
  and g28727 (n17435, \asqrt[11] , n17434);
  not g28728 (n_11646, n17435);
  and g28729 (n17436, n_11209, n_11646);
  not g28730 (n_11647, n17433);
  not g28731 (n_11648, n17436);
  and g28732 (n17437, n_11647, n_11648);
  and g28733 (n17438, n_3242, n_11643);
  and g28734 (n17439, n_11644, n17438);
  not g28735 (n_11649, n17437);
  not g28736 (n_11650, n17439);
  and g28737 (n17440, n_11649, n_11650);
  not g28738 (n_11651, n17430);
  not g28739 (n_11652, n17440);
  and g28740 (n17441, n_11651, n_11652);
  not g28741 (n_11653, n17441);
  and g28742 (n17442, \asqrt[39] , n_11653);
  and g28746 (n17446, n_11219, n_11218);
  and g28747 (n17447, \asqrt[11] , n17446);
  not g28748 (n_11654, n17447);
  and g28749 (n17448, n_11217, n_11654);
  not g28750 (n_11655, n17445);
  not g28751 (n_11656, n17448);
  and g28752 (n17449, n_11655, n_11656);
  and g28753 (n17450, n_3018, n_11651);
  and g28754 (n17451, n_11652, n17450);
  not g28755 (n_11657, n17449);
  not g28756 (n_11658, n17451);
  and g28757 (n17452, n_11657, n_11658);
  not g28758 (n_11659, n17442);
  not g28759 (n_11660, n17452);
  and g28760 (n17453, n_11659, n_11660);
  not g28761 (n_11661, n17453);
  and g28762 (n17454, \asqrt[40] , n_11661);
  and g28766 (n17458, n_11227, n_11226);
  and g28767 (n17459, \asqrt[11] , n17458);
  not g28768 (n_11662, n17459);
  and g28769 (n17460, n_11225, n_11662);
  not g28770 (n_11663, n17457);
  not g28771 (n_11664, n17460);
  and g28772 (n17461, n_11663, n_11664);
  and g28773 (n17462, n_2802, n_11659);
  and g28774 (n17463, n_11660, n17462);
  not g28775 (n_11665, n17461);
  not g28776 (n_11666, n17463);
  and g28777 (n17464, n_11665, n_11666);
  not g28778 (n_11667, n17454);
  not g28779 (n_11668, n17464);
  and g28780 (n17465, n_11667, n_11668);
  not g28781 (n_11669, n17465);
  and g28782 (n17466, \asqrt[41] , n_11669);
  and g28786 (n17470, n_11235, n_11234);
  and g28787 (n17471, \asqrt[11] , n17470);
  not g28788 (n_11670, n17471);
  and g28789 (n17472, n_11233, n_11670);
  not g28790 (n_11671, n17469);
  not g28791 (n_11672, n17472);
  and g28792 (n17473, n_11671, n_11672);
  and g28793 (n17474, n_2594, n_11667);
  and g28794 (n17475, n_11668, n17474);
  not g28795 (n_11673, n17473);
  not g28796 (n_11674, n17475);
  and g28797 (n17476, n_11673, n_11674);
  not g28798 (n_11675, n17466);
  not g28799 (n_11676, n17476);
  and g28800 (n17477, n_11675, n_11676);
  not g28801 (n_11677, n17477);
  and g28802 (n17478, \asqrt[42] , n_11677);
  and g28806 (n17482, n_11243, n_11242);
  and g28807 (n17483, \asqrt[11] , n17482);
  not g28808 (n_11678, n17483);
  and g28809 (n17484, n_11241, n_11678);
  not g28810 (n_11679, n17481);
  not g28811 (n_11680, n17484);
  and g28812 (n17485, n_11679, n_11680);
  and g28813 (n17486, n_2394, n_11675);
  and g28814 (n17487, n_11676, n17486);
  not g28815 (n_11681, n17485);
  not g28816 (n_11682, n17487);
  and g28817 (n17488, n_11681, n_11682);
  not g28818 (n_11683, n17478);
  not g28819 (n_11684, n17488);
  and g28820 (n17489, n_11683, n_11684);
  not g28821 (n_11685, n17489);
  and g28822 (n17490, \asqrt[43] , n_11685);
  and g28826 (n17494, n_11251, n_11250);
  and g28827 (n17495, \asqrt[11] , n17494);
  not g28828 (n_11686, n17495);
  and g28829 (n17496, n_11249, n_11686);
  not g28830 (n_11687, n17493);
  not g28831 (n_11688, n17496);
  and g28832 (n17497, n_11687, n_11688);
  and g28833 (n17498, n_2202, n_11683);
  and g28834 (n17499, n_11684, n17498);
  not g28835 (n_11689, n17497);
  not g28836 (n_11690, n17499);
  and g28837 (n17500, n_11689, n_11690);
  not g28838 (n_11691, n17490);
  not g28839 (n_11692, n17500);
  and g28840 (n17501, n_11691, n_11692);
  not g28841 (n_11693, n17501);
  and g28842 (n17502, \asqrt[44] , n_11693);
  and g28846 (n17506, n_11259, n_11258);
  and g28847 (n17507, \asqrt[11] , n17506);
  not g28848 (n_11694, n17507);
  and g28849 (n17508, n_11257, n_11694);
  not g28850 (n_11695, n17505);
  not g28851 (n_11696, n17508);
  and g28852 (n17509, n_11695, n_11696);
  and g28853 (n17510, n_2018, n_11691);
  and g28854 (n17511, n_11692, n17510);
  not g28855 (n_11697, n17509);
  not g28856 (n_11698, n17511);
  and g28857 (n17512, n_11697, n_11698);
  not g28858 (n_11699, n17502);
  not g28859 (n_11700, n17512);
  and g28860 (n17513, n_11699, n_11700);
  not g28861 (n_11701, n17513);
  and g28862 (n17514, \asqrt[45] , n_11701);
  and g28866 (n17518, n_11267, n_11266);
  and g28867 (n17519, \asqrt[11] , n17518);
  not g28868 (n_11702, n17519);
  and g28869 (n17520, n_11265, n_11702);
  not g28870 (n_11703, n17517);
  not g28871 (n_11704, n17520);
  and g28872 (n17521, n_11703, n_11704);
  and g28873 (n17522, n_1842, n_11699);
  and g28874 (n17523, n_11700, n17522);
  not g28875 (n_11705, n17521);
  not g28876 (n_11706, n17523);
  and g28877 (n17524, n_11705, n_11706);
  not g28878 (n_11707, n17514);
  not g28879 (n_11708, n17524);
  and g28880 (n17525, n_11707, n_11708);
  not g28881 (n_11709, n17525);
  and g28882 (n17526, \asqrt[46] , n_11709);
  and g28886 (n17530, n_11275, n_11274);
  and g28887 (n17531, \asqrt[11] , n17530);
  not g28888 (n_11710, n17531);
  and g28889 (n17532, n_11273, n_11710);
  not g28890 (n_11711, n17529);
  not g28891 (n_11712, n17532);
  and g28892 (n17533, n_11711, n_11712);
  and g28893 (n17534, n_1674, n_11707);
  and g28894 (n17535, n_11708, n17534);
  not g28895 (n_11713, n17533);
  not g28896 (n_11714, n17535);
  and g28897 (n17536, n_11713, n_11714);
  not g28898 (n_11715, n17526);
  not g28899 (n_11716, n17536);
  and g28900 (n17537, n_11715, n_11716);
  not g28901 (n_11717, n17537);
  and g28902 (n17538, \asqrt[47] , n_11717);
  and g28906 (n17542, n_11283, n_11282);
  and g28907 (n17543, \asqrt[11] , n17542);
  not g28908 (n_11718, n17543);
  and g28909 (n17544, n_11281, n_11718);
  not g28910 (n_11719, n17541);
  not g28911 (n_11720, n17544);
  and g28912 (n17545, n_11719, n_11720);
  and g28913 (n17546, n_1514, n_11715);
  and g28914 (n17547, n_11716, n17546);
  not g28915 (n_11721, n17545);
  not g28916 (n_11722, n17547);
  and g28917 (n17548, n_11721, n_11722);
  not g28918 (n_11723, n17538);
  not g28919 (n_11724, n17548);
  and g28920 (n17549, n_11723, n_11724);
  not g28921 (n_11725, n17549);
  and g28922 (n17550, \asqrt[48] , n_11725);
  and g28926 (n17554, n_11291, n_11290);
  and g28927 (n17555, \asqrt[11] , n17554);
  not g28928 (n_11726, n17555);
  and g28929 (n17556, n_11289, n_11726);
  not g28930 (n_11727, n17553);
  not g28931 (n_11728, n17556);
  and g28932 (n17557, n_11727, n_11728);
  and g28933 (n17558, n_1362, n_11723);
  and g28934 (n17559, n_11724, n17558);
  not g28935 (n_11729, n17557);
  not g28936 (n_11730, n17559);
  and g28937 (n17560, n_11729, n_11730);
  not g28938 (n_11731, n17550);
  not g28939 (n_11732, n17560);
  and g28940 (n17561, n_11731, n_11732);
  not g28941 (n_11733, n17561);
  and g28942 (n17562, \asqrt[49] , n_11733);
  and g28946 (n17566, n_11299, n_11298);
  and g28947 (n17567, \asqrt[11] , n17566);
  not g28948 (n_11734, n17567);
  and g28949 (n17568, n_11297, n_11734);
  not g28950 (n_11735, n17565);
  not g28951 (n_11736, n17568);
  and g28952 (n17569, n_11735, n_11736);
  and g28953 (n17570, n_1218, n_11731);
  and g28954 (n17571, n_11732, n17570);
  not g28955 (n_11737, n17569);
  not g28956 (n_11738, n17571);
  and g28957 (n17572, n_11737, n_11738);
  not g28958 (n_11739, n17562);
  not g28959 (n_11740, n17572);
  and g28960 (n17573, n_11739, n_11740);
  not g28961 (n_11741, n17573);
  and g28962 (n17574, \asqrt[50] , n_11741);
  and g28966 (n17578, n_11307, n_11306);
  and g28967 (n17579, \asqrt[11] , n17578);
  not g28968 (n_11742, n17579);
  and g28969 (n17580, n_11305, n_11742);
  not g28970 (n_11743, n17577);
  not g28971 (n_11744, n17580);
  and g28972 (n17581, n_11743, n_11744);
  and g28973 (n17582, n_1082, n_11739);
  and g28974 (n17583, n_11740, n17582);
  not g28975 (n_11745, n17581);
  not g28976 (n_11746, n17583);
  and g28977 (n17584, n_11745, n_11746);
  not g28978 (n_11747, n17574);
  not g28979 (n_11748, n17584);
  and g28980 (n17585, n_11747, n_11748);
  not g28981 (n_11749, n17585);
  and g28982 (n17586, \asqrt[51] , n_11749);
  and g28986 (n17590, n_11315, n_11314);
  and g28987 (n17591, \asqrt[11] , n17590);
  not g28988 (n_11750, n17591);
  and g28989 (n17592, n_11313, n_11750);
  not g28990 (n_11751, n17589);
  not g28991 (n_11752, n17592);
  and g28992 (n17593, n_11751, n_11752);
  and g28993 (n17594, n_954, n_11747);
  and g28994 (n17595, n_11748, n17594);
  not g28995 (n_11753, n17593);
  not g28996 (n_11754, n17595);
  and g28997 (n17596, n_11753, n_11754);
  not g28998 (n_11755, n17586);
  not g28999 (n_11756, n17596);
  and g29000 (n17597, n_11755, n_11756);
  not g29001 (n_11757, n17597);
  and g29002 (n17598, \asqrt[52] , n_11757);
  and g29006 (n17602, n_11323, n_11322);
  and g29007 (n17603, \asqrt[11] , n17602);
  not g29008 (n_11758, n17603);
  and g29009 (n17604, n_11321, n_11758);
  not g29010 (n_11759, n17601);
  not g29011 (n_11760, n17604);
  and g29012 (n17605, n_11759, n_11760);
  and g29013 (n17606, n_834, n_11755);
  and g29014 (n17607, n_11756, n17606);
  not g29015 (n_11761, n17605);
  not g29016 (n_11762, n17607);
  and g29017 (n17608, n_11761, n_11762);
  not g29018 (n_11763, n17598);
  not g29019 (n_11764, n17608);
  and g29020 (n17609, n_11763, n_11764);
  not g29021 (n_11765, n17609);
  and g29022 (n17610, \asqrt[53] , n_11765);
  and g29026 (n17614, n_11331, n_11330);
  and g29027 (n17615, \asqrt[11] , n17614);
  not g29028 (n_11766, n17615);
  and g29029 (n17616, n_11329, n_11766);
  not g29030 (n_11767, n17613);
  not g29031 (n_11768, n17616);
  and g29032 (n17617, n_11767, n_11768);
  and g29033 (n17618, n_722, n_11763);
  and g29034 (n17619, n_11764, n17618);
  not g29035 (n_11769, n17617);
  not g29036 (n_11770, n17619);
  and g29037 (n17620, n_11769, n_11770);
  not g29038 (n_11771, n17610);
  not g29039 (n_11772, n17620);
  and g29040 (n17621, n_11771, n_11772);
  not g29041 (n_11773, n17621);
  and g29042 (n17622, \asqrt[54] , n_11773);
  and g29043 (n17623, n_618, n_11771);
  and g29044 (n17624, n_11772, n17623);
  and g29048 (n17628, n_11339, n_11337);
  and g29049 (n17629, \asqrt[11] , n17628);
  not g29050 (n_11774, n17629);
  and g29051 (n17630, n_11338, n_11774);
  not g29052 (n_11775, n17627);
  not g29053 (n_11776, n17630);
  and g29054 (n17631, n_11775, n_11776);
  not g29055 (n_11777, n17624);
  not g29056 (n_11778, n17631);
  and g29057 (n17632, n_11777, n_11778);
  not g29058 (n_11779, n17622);
  not g29059 (n_11780, n17632);
  and g29060 (n17633, n_11779, n_11780);
  not g29061 (n_11781, n17633);
  and g29062 (n17634, \asqrt[55] , n_11781);
  and g29066 (n17638, n_11347, n_11346);
  and g29067 (n17639, \asqrt[11] , n17638);
  not g29068 (n_11782, n17639);
  and g29069 (n17640, n_11345, n_11782);
  not g29070 (n_11783, n17637);
  not g29071 (n_11784, n17640);
  and g29072 (n17641, n_11783, n_11784);
  and g29073 (n17642, n_522, n_11779);
  and g29074 (n17643, n_11780, n17642);
  not g29075 (n_11785, n17641);
  not g29076 (n_11786, n17643);
  and g29077 (n17644, n_11785, n_11786);
  not g29078 (n_11787, n17634);
  not g29079 (n_11788, n17644);
  and g29080 (n17645, n_11787, n_11788);
  not g29081 (n_11789, n17645);
  and g29082 (n17646, \asqrt[56] , n_11789);
  and g29086 (n17650, n_11355, n_11354);
  and g29087 (n17651, \asqrt[11] , n17650);
  not g29088 (n_11790, n17651);
  and g29089 (n17652, n_11353, n_11790);
  not g29090 (n_11791, n17649);
  not g29091 (n_11792, n17652);
  and g29092 (n17653, n_11791, n_11792);
  and g29093 (n17654, n_434, n_11787);
  and g29094 (n17655, n_11788, n17654);
  not g29095 (n_11793, n17653);
  not g29096 (n_11794, n17655);
  and g29097 (n17656, n_11793, n_11794);
  not g29098 (n_11795, n17646);
  not g29099 (n_11796, n17656);
  and g29100 (n17657, n_11795, n_11796);
  not g29101 (n_11797, n17657);
  and g29102 (n17658, \asqrt[57] , n_11797);
  and g29106 (n17662, n_11363, n_11362);
  and g29107 (n17663, \asqrt[11] , n17662);
  not g29108 (n_11798, n17663);
  and g29109 (n17664, n_11361, n_11798);
  not g29110 (n_11799, n17661);
  not g29111 (n_11800, n17664);
  and g29112 (n17665, n_11799, n_11800);
  and g29113 (n17666, n_354, n_11795);
  and g29114 (n17667, n_11796, n17666);
  not g29115 (n_11801, n17665);
  not g29116 (n_11802, n17667);
  and g29117 (n17668, n_11801, n_11802);
  not g29118 (n_11803, n17658);
  not g29119 (n_11804, n17668);
  and g29120 (n17669, n_11803, n_11804);
  not g29121 (n_11805, n17669);
  and g29122 (n17670, \asqrt[58] , n_11805);
  and g29126 (n17674, n_11371, n_11370);
  and g29127 (n17675, \asqrt[11] , n17674);
  not g29128 (n_11806, n17675);
  and g29129 (n17676, n_11369, n_11806);
  not g29130 (n_11807, n17673);
  not g29131 (n_11808, n17676);
  and g29132 (n17677, n_11807, n_11808);
  and g29133 (n17678, n_282, n_11803);
  and g29134 (n17679, n_11804, n17678);
  not g29135 (n_11809, n17677);
  not g29136 (n_11810, n17679);
  and g29137 (n17680, n_11809, n_11810);
  not g29138 (n_11811, n17670);
  not g29139 (n_11812, n17680);
  and g29140 (n17681, n_11811, n_11812);
  not g29141 (n_11813, n17681);
  and g29142 (n17682, \asqrt[59] , n_11813);
  and g29146 (n17686, n_11379, n_11378);
  and g29147 (n17687, \asqrt[11] , n17686);
  not g29148 (n_11814, n17687);
  and g29149 (n17688, n_11377, n_11814);
  not g29150 (n_11815, n17685);
  not g29151 (n_11816, n17688);
  and g29152 (n17689, n_11815, n_11816);
  and g29153 (n17690, n_218, n_11811);
  and g29154 (n17691, n_11812, n17690);
  not g29155 (n_11817, n17689);
  not g29156 (n_11818, n17691);
  and g29157 (n17692, n_11817, n_11818);
  not g29158 (n_11819, n17682);
  not g29159 (n_11820, n17692);
  and g29160 (n17693, n_11819, n_11820);
  not g29161 (n_11821, n17693);
  and g29162 (n17694, \asqrt[60] , n_11821);
  and g29166 (n17698, n_11387, n_11386);
  and g29167 (n17699, \asqrt[11] , n17698);
  not g29168 (n_11822, n17699);
  and g29169 (n17700, n_11385, n_11822);
  not g29170 (n_11823, n17697);
  not g29171 (n_11824, n17700);
  and g29172 (n17701, n_11823, n_11824);
  and g29173 (n17702, n_162, n_11819);
  and g29174 (n17703, n_11820, n17702);
  not g29175 (n_11825, n17701);
  not g29176 (n_11826, n17703);
  and g29177 (n17704, n_11825, n_11826);
  not g29178 (n_11827, n17694);
  not g29179 (n_11828, n17704);
  and g29180 (n17705, n_11827, n_11828);
  not g29181 (n_11829, n17705);
  and g29182 (n17706, \asqrt[61] , n_11829);
  and g29186 (n17710, n_11395, n_11394);
  and g29187 (n17711, \asqrt[11] , n17710);
  not g29188 (n_11830, n17711);
  and g29189 (n17712, n_11393, n_11830);
  not g29190 (n_11831, n17709);
  not g29191 (n_11832, n17712);
  and g29192 (n17713, n_11831, n_11832);
  and g29193 (n17714, n_115, n_11827);
  and g29194 (n17715, n_11828, n17714);
  not g29195 (n_11833, n17713);
  not g29196 (n_11834, n17715);
  and g29197 (n17716, n_11833, n_11834);
  not g29198 (n_11835, n17706);
  not g29199 (n_11836, n17716);
  and g29200 (n17717, n_11835, n_11836);
  not g29201 (n_11837, n17717);
  and g29202 (n17718, \asqrt[62] , n_11837);
  and g29206 (n17722, n_11403, n_11402);
  and g29207 (n17723, \asqrt[11] , n17722);
  not g29208 (n_11838, n17723);
  and g29209 (n17724, n_11401, n_11838);
  not g29210 (n_11839, n17721);
  not g29211 (n_11840, n17724);
  and g29212 (n17725, n_11839, n_11840);
  and g29213 (n17726, n_76, n_11835);
  and g29214 (n17727, n_11836, n17726);
  not g29215 (n_11841, n17725);
  not g29216 (n_11842, n17727);
  and g29217 (n17728, n_11841, n_11842);
  not g29218 (n_11843, n17718);
  not g29219 (n_11844, n17728);
  and g29220 (n17729, n_11843, n_11844);
  and g29224 (n17733, n_11411, n_11410);
  and g29225 (n17734, \asqrt[11] , n17733);
  not g29226 (n_11845, n17734);
  and g29227 (n17735, n_11409, n_11845);
  not g29228 (n_11846, n17732);
  not g29229 (n_11847, n17735);
  and g29230 (n17736, n_11846, n_11847);
  and g29231 (n17737, n_11418, n_11417);
  and g29232 (n17738, \asqrt[11] , n17737);
  not g29235 (n_11849, n17736);
  not g29237 (n_11850, n17729);
  not g29239 (n_11851, n17741);
  and g29240 (n17742, n_21, n_11851);
  and g29241 (n17743, n_11843, n17736);
  and g29242 (n17744, n_11844, n17743);
  and g29243 (n17745, n_11417, \asqrt[11] );
  not g29244 (n_11852, n17745);
  and g29245 (n17746, n17085, n_11852);
  not g29246 (n_11853, n17737);
  and g29247 (n17747, \asqrt[63] , n_11853);
  not g29248 (n_11854, n17746);
  and g29249 (n17748, n_11854, n17747);
  not g29255 (n_11855, n17748);
  not g29256 (n_11856, n17753);
  not g29258 (n_11857, n17744);
  and g29262 (n17757, \a[20] , \asqrt[10] );
  not g29263 (n_11862, \a[18] );
  not g29264 (n_11863, \a[19] );
  and g29265 (n17758, n_11862, n_11863);
  and g29266 (n17759, n_11430, n17758);
  not g29267 (n_11864, n17757);
  not g29268 (n_11865, n17759);
  and g29269 (n17760, n_11864, n_11865);
  not g29270 (n_11866, n17760);
  and g29271 (n17761, \asqrt[11] , n_11866);
  and g29277 (n17767, n_11430, \asqrt[10] );
  not g29278 (n_11867, n17767);
  and g29279 (n17768, \a[21] , n_11867);
  and g29280 (n17769, n17114, \asqrt[10] );
  not g29281 (n_11868, n17768);
  not g29282 (n_11869, n17769);
  and g29283 (n17770, n_11868, n_11869);
  not g29284 (n_11870, n17766);
  and g29285 (n17771, n_11870, n17770);
  not g29286 (n_11871, n17761);
  not g29287 (n_11872, n17771);
  and g29288 (n17772, n_11871, n_11872);
  not g29289 (n_11873, n17772);
  and g29290 (n17773, \asqrt[12] , n_11873);
  not g29291 (n_11874, \asqrt[12] );
  and g29292 (n17774, n_11874, n_11871);
  and g29293 (n17775, n_11872, n17774);
  not g29297 (n_11875, n17742);
  not g29299 (n_11876, n17779);
  and g29300 (n17780, n_11869, n_11876);
  not g29301 (n_11877, n17780);
  and g29302 (n17781, \a[22] , n_11877);
  and g29303 (n17782, n_11006, n_11876);
  and g29304 (n17783, n_11869, n17782);
  not g29305 (n_11878, n17781);
  not g29306 (n_11879, n17783);
  and g29307 (n17784, n_11878, n_11879);
  not g29308 (n_11880, n17775);
  not g29309 (n_11881, n17784);
  and g29310 (n17785, n_11880, n_11881);
  not g29311 (n_11882, n17773);
  not g29312 (n_11883, n17785);
  and g29313 (n17786, n_11882, n_11883);
  not g29314 (n_11884, n17786);
  and g29315 (n17787, \asqrt[13] , n_11884);
  and g29316 (n17788, n_11439, n_11438);
  not g29317 (n_11885, n17126);
  and g29318 (n17789, n_11885, n17788);
  and g29319 (n17790, \asqrt[10] , n17789);
  and g29320 (n17791, \asqrt[10] , n17788);
  not g29321 (n_11886, n17791);
  and g29322 (n17792, n17126, n_11886);
  not g29323 (n_11887, n17790);
  not g29324 (n_11888, n17792);
  and g29325 (n17793, n_11887, n_11888);
  and g29326 (n17794, n_11442, n_11882);
  and g29327 (n17795, n_11883, n17794);
  not g29328 (n_11889, n17793);
  not g29329 (n_11890, n17795);
  and g29330 (n17796, n_11889, n_11890);
  not g29331 (n_11891, n17787);
  not g29332 (n_11892, n17796);
  and g29333 (n17797, n_11891, n_11892);
  not g29334 (n_11893, n17797);
  and g29335 (n17798, \asqrt[14] , n_11893);
  and g29339 (n17802, n_11450, n_11448);
  and g29340 (n17803, \asqrt[10] , n17802);
  not g29341 (n_11894, n17803);
  and g29342 (n17804, n_11449, n_11894);
  not g29343 (n_11895, n17801);
  not g29344 (n_11896, n17804);
  and g29345 (n17805, n_11895, n_11896);
  and g29346 (n17806, n_11018, n_11891);
  and g29347 (n17807, n_11892, n17806);
  not g29348 (n_11897, n17805);
  not g29349 (n_11898, n17807);
  and g29350 (n17808, n_11897, n_11898);
  not g29351 (n_11899, n17798);
  not g29352 (n_11900, n17808);
  and g29353 (n17809, n_11899, n_11900);
  not g29354 (n_11901, n17809);
  and g29355 (n17810, \asqrt[15] , n_11901);
  and g29359 (n17814, n_11459, n_11458);
  and g29360 (n17815, \asqrt[10] , n17814);
  not g29361 (n_11902, n17815);
  and g29362 (n17816, n_11457, n_11902);
  not g29363 (n_11903, n17813);
  not g29364 (n_11904, n17816);
  and g29365 (n17817, n_11903, n_11904);
  and g29366 (n17818, n_10602, n_11899);
  and g29367 (n17819, n_11900, n17818);
  not g29368 (n_11905, n17817);
  not g29369 (n_11906, n17819);
  and g29370 (n17820, n_11905, n_11906);
  not g29371 (n_11907, n17810);
  not g29372 (n_11908, n17820);
  and g29373 (n17821, n_11907, n_11908);
  not g29374 (n_11909, n17821);
  and g29375 (n17822, \asqrt[16] , n_11909);
  and g29379 (n17826, n_11467, n_11466);
  and g29380 (n17827, \asqrt[10] , n17826);
  not g29381 (n_11910, n17827);
  and g29382 (n17828, n_11465, n_11910);
  not g29383 (n_11911, n17825);
  not g29384 (n_11912, n17828);
  and g29385 (n17829, n_11911, n_11912);
  and g29386 (n17830, n_10194, n_11907);
  and g29387 (n17831, n_11908, n17830);
  not g29388 (n_11913, n17829);
  not g29389 (n_11914, n17831);
  and g29390 (n17832, n_11913, n_11914);
  not g29391 (n_11915, n17822);
  not g29392 (n_11916, n17832);
  and g29393 (n17833, n_11915, n_11916);
  not g29394 (n_11917, n17833);
  and g29395 (n17834, \asqrt[17] , n_11917);
  and g29399 (n17838, n_11475, n_11474);
  and g29400 (n17839, \asqrt[10] , n17838);
  not g29401 (n_11918, n17839);
  and g29402 (n17840, n_11473, n_11918);
  not g29403 (n_11919, n17837);
  not g29404 (n_11920, n17840);
  and g29405 (n17841, n_11919, n_11920);
  and g29406 (n17842, n_9794, n_11915);
  and g29407 (n17843, n_11916, n17842);
  not g29408 (n_11921, n17841);
  not g29409 (n_11922, n17843);
  and g29410 (n17844, n_11921, n_11922);
  not g29411 (n_11923, n17834);
  not g29412 (n_11924, n17844);
  and g29413 (n17845, n_11923, n_11924);
  not g29414 (n_11925, n17845);
  and g29415 (n17846, \asqrt[18] , n_11925);
  and g29419 (n17850, n_11483, n_11482);
  and g29420 (n17851, \asqrt[10] , n17850);
  not g29421 (n_11926, n17851);
  and g29422 (n17852, n_11481, n_11926);
  not g29423 (n_11927, n17849);
  not g29424 (n_11928, n17852);
  and g29425 (n17853, n_11927, n_11928);
  and g29426 (n17854, n_9402, n_11923);
  and g29427 (n17855, n_11924, n17854);
  not g29428 (n_11929, n17853);
  not g29429 (n_11930, n17855);
  and g29430 (n17856, n_11929, n_11930);
  not g29431 (n_11931, n17846);
  not g29432 (n_11932, n17856);
  and g29433 (n17857, n_11931, n_11932);
  not g29434 (n_11933, n17857);
  and g29435 (n17858, \asqrt[19] , n_11933);
  and g29439 (n17862, n_11491, n_11490);
  and g29440 (n17863, \asqrt[10] , n17862);
  not g29441 (n_11934, n17863);
  and g29442 (n17864, n_11489, n_11934);
  not g29443 (n_11935, n17861);
  not g29444 (n_11936, n17864);
  and g29445 (n17865, n_11935, n_11936);
  and g29446 (n17866, n_9018, n_11931);
  and g29447 (n17867, n_11932, n17866);
  not g29448 (n_11937, n17865);
  not g29449 (n_11938, n17867);
  and g29450 (n17868, n_11937, n_11938);
  not g29451 (n_11939, n17858);
  not g29452 (n_11940, n17868);
  and g29453 (n17869, n_11939, n_11940);
  not g29454 (n_11941, n17869);
  and g29455 (n17870, \asqrt[20] , n_11941);
  and g29459 (n17874, n_11499, n_11498);
  and g29460 (n17875, \asqrt[10] , n17874);
  not g29461 (n_11942, n17875);
  and g29462 (n17876, n_11497, n_11942);
  not g29463 (n_11943, n17873);
  not g29464 (n_11944, n17876);
  and g29465 (n17877, n_11943, n_11944);
  and g29466 (n17878, n_8642, n_11939);
  and g29467 (n17879, n_11940, n17878);
  not g29468 (n_11945, n17877);
  not g29469 (n_11946, n17879);
  and g29470 (n17880, n_11945, n_11946);
  not g29471 (n_11947, n17870);
  not g29472 (n_11948, n17880);
  and g29473 (n17881, n_11947, n_11948);
  not g29474 (n_11949, n17881);
  and g29475 (n17882, \asqrt[21] , n_11949);
  and g29479 (n17886, n_11507, n_11506);
  and g29480 (n17887, \asqrt[10] , n17886);
  not g29481 (n_11950, n17887);
  and g29482 (n17888, n_11505, n_11950);
  not g29483 (n_11951, n17885);
  not g29484 (n_11952, n17888);
  and g29485 (n17889, n_11951, n_11952);
  and g29486 (n17890, n_8274, n_11947);
  and g29487 (n17891, n_11948, n17890);
  not g29488 (n_11953, n17889);
  not g29489 (n_11954, n17891);
  and g29490 (n17892, n_11953, n_11954);
  not g29491 (n_11955, n17882);
  not g29492 (n_11956, n17892);
  and g29493 (n17893, n_11955, n_11956);
  not g29494 (n_11957, n17893);
  and g29495 (n17894, \asqrt[22] , n_11957);
  and g29499 (n17898, n_11515, n_11514);
  and g29500 (n17899, \asqrt[10] , n17898);
  not g29501 (n_11958, n17899);
  and g29502 (n17900, n_11513, n_11958);
  not g29503 (n_11959, n17897);
  not g29504 (n_11960, n17900);
  and g29505 (n17901, n_11959, n_11960);
  and g29506 (n17902, n_7914, n_11955);
  and g29507 (n17903, n_11956, n17902);
  not g29508 (n_11961, n17901);
  not g29509 (n_11962, n17903);
  and g29510 (n17904, n_11961, n_11962);
  not g29511 (n_11963, n17894);
  not g29512 (n_11964, n17904);
  and g29513 (n17905, n_11963, n_11964);
  not g29514 (n_11965, n17905);
  and g29515 (n17906, \asqrt[23] , n_11965);
  and g29519 (n17910, n_11523, n_11522);
  and g29520 (n17911, \asqrt[10] , n17910);
  not g29521 (n_11966, n17911);
  and g29522 (n17912, n_11521, n_11966);
  not g29523 (n_11967, n17909);
  not g29524 (n_11968, n17912);
  and g29525 (n17913, n_11967, n_11968);
  and g29526 (n17914, n_7562, n_11963);
  and g29527 (n17915, n_11964, n17914);
  not g29528 (n_11969, n17913);
  not g29529 (n_11970, n17915);
  and g29530 (n17916, n_11969, n_11970);
  not g29531 (n_11971, n17906);
  not g29532 (n_11972, n17916);
  and g29533 (n17917, n_11971, n_11972);
  not g29534 (n_11973, n17917);
  and g29535 (n17918, \asqrt[24] , n_11973);
  and g29539 (n17922, n_11531, n_11530);
  and g29540 (n17923, \asqrt[10] , n17922);
  not g29541 (n_11974, n17923);
  and g29542 (n17924, n_11529, n_11974);
  not g29543 (n_11975, n17921);
  not g29544 (n_11976, n17924);
  and g29545 (n17925, n_11975, n_11976);
  and g29546 (n17926, n_7218, n_11971);
  and g29547 (n17927, n_11972, n17926);
  not g29548 (n_11977, n17925);
  not g29549 (n_11978, n17927);
  and g29550 (n17928, n_11977, n_11978);
  not g29551 (n_11979, n17918);
  not g29552 (n_11980, n17928);
  and g29553 (n17929, n_11979, n_11980);
  not g29554 (n_11981, n17929);
  and g29555 (n17930, \asqrt[25] , n_11981);
  and g29559 (n17934, n_11539, n_11538);
  and g29560 (n17935, \asqrt[10] , n17934);
  not g29561 (n_11982, n17935);
  and g29562 (n17936, n_11537, n_11982);
  not g29563 (n_11983, n17933);
  not g29564 (n_11984, n17936);
  and g29565 (n17937, n_11983, n_11984);
  and g29566 (n17938, n_6882, n_11979);
  and g29567 (n17939, n_11980, n17938);
  not g29568 (n_11985, n17937);
  not g29569 (n_11986, n17939);
  and g29570 (n17940, n_11985, n_11986);
  not g29571 (n_11987, n17930);
  not g29572 (n_11988, n17940);
  and g29573 (n17941, n_11987, n_11988);
  not g29574 (n_11989, n17941);
  and g29575 (n17942, \asqrt[26] , n_11989);
  and g29579 (n17946, n_11547, n_11546);
  and g29580 (n17947, \asqrt[10] , n17946);
  not g29581 (n_11990, n17947);
  and g29582 (n17948, n_11545, n_11990);
  not g29583 (n_11991, n17945);
  not g29584 (n_11992, n17948);
  and g29585 (n17949, n_11991, n_11992);
  and g29586 (n17950, n_6554, n_11987);
  and g29587 (n17951, n_11988, n17950);
  not g29588 (n_11993, n17949);
  not g29589 (n_11994, n17951);
  and g29590 (n17952, n_11993, n_11994);
  not g29591 (n_11995, n17942);
  not g29592 (n_11996, n17952);
  and g29593 (n17953, n_11995, n_11996);
  not g29594 (n_11997, n17953);
  and g29595 (n17954, \asqrt[27] , n_11997);
  and g29599 (n17958, n_11555, n_11554);
  and g29600 (n17959, \asqrt[10] , n17958);
  not g29601 (n_11998, n17959);
  and g29602 (n17960, n_11553, n_11998);
  not g29603 (n_11999, n17957);
  not g29604 (n_12000, n17960);
  and g29605 (n17961, n_11999, n_12000);
  and g29606 (n17962, n_6234, n_11995);
  and g29607 (n17963, n_11996, n17962);
  not g29608 (n_12001, n17961);
  not g29609 (n_12002, n17963);
  and g29610 (n17964, n_12001, n_12002);
  not g29611 (n_12003, n17954);
  not g29612 (n_12004, n17964);
  and g29613 (n17965, n_12003, n_12004);
  not g29614 (n_12005, n17965);
  and g29615 (n17966, \asqrt[28] , n_12005);
  and g29619 (n17970, n_11563, n_11562);
  and g29620 (n17971, \asqrt[10] , n17970);
  not g29621 (n_12006, n17971);
  and g29622 (n17972, n_11561, n_12006);
  not g29623 (n_12007, n17969);
  not g29624 (n_12008, n17972);
  and g29625 (n17973, n_12007, n_12008);
  and g29626 (n17974, n_5922, n_12003);
  and g29627 (n17975, n_12004, n17974);
  not g29628 (n_12009, n17973);
  not g29629 (n_12010, n17975);
  and g29630 (n17976, n_12009, n_12010);
  not g29631 (n_12011, n17966);
  not g29632 (n_12012, n17976);
  and g29633 (n17977, n_12011, n_12012);
  not g29634 (n_12013, n17977);
  and g29635 (n17978, \asqrt[29] , n_12013);
  and g29639 (n17982, n_11571, n_11570);
  and g29640 (n17983, \asqrt[10] , n17982);
  not g29641 (n_12014, n17983);
  and g29642 (n17984, n_11569, n_12014);
  not g29643 (n_12015, n17981);
  not g29644 (n_12016, n17984);
  and g29645 (n17985, n_12015, n_12016);
  and g29646 (n17986, n_5618, n_12011);
  and g29647 (n17987, n_12012, n17986);
  not g29648 (n_12017, n17985);
  not g29649 (n_12018, n17987);
  and g29650 (n17988, n_12017, n_12018);
  not g29651 (n_12019, n17978);
  not g29652 (n_12020, n17988);
  and g29653 (n17989, n_12019, n_12020);
  not g29654 (n_12021, n17989);
  and g29655 (n17990, \asqrt[30] , n_12021);
  and g29659 (n17994, n_11579, n_11578);
  and g29660 (n17995, \asqrt[10] , n17994);
  not g29661 (n_12022, n17995);
  and g29662 (n17996, n_11577, n_12022);
  not g29663 (n_12023, n17993);
  not g29664 (n_12024, n17996);
  and g29665 (n17997, n_12023, n_12024);
  and g29666 (n17998, n_5322, n_12019);
  and g29667 (n17999, n_12020, n17998);
  not g29668 (n_12025, n17997);
  not g29669 (n_12026, n17999);
  and g29670 (n18000, n_12025, n_12026);
  not g29671 (n_12027, n17990);
  not g29672 (n_12028, n18000);
  and g29673 (n18001, n_12027, n_12028);
  not g29674 (n_12029, n18001);
  and g29675 (n18002, \asqrt[31] , n_12029);
  and g29679 (n18006, n_11587, n_11586);
  and g29680 (n18007, \asqrt[10] , n18006);
  not g29681 (n_12030, n18007);
  and g29682 (n18008, n_11585, n_12030);
  not g29683 (n_12031, n18005);
  not g29684 (n_12032, n18008);
  and g29685 (n18009, n_12031, n_12032);
  and g29686 (n18010, n_5034, n_12027);
  and g29687 (n18011, n_12028, n18010);
  not g29688 (n_12033, n18009);
  not g29689 (n_12034, n18011);
  and g29690 (n18012, n_12033, n_12034);
  not g29691 (n_12035, n18002);
  not g29692 (n_12036, n18012);
  and g29693 (n18013, n_12035, n_12036);
  not g29694 (n_12037, n18013);
  and g29695 (n18014, \asqrt[32] , n_12037);
  and g29699 (n18018, n_11595, n_11594);
  and g29700 (n18019, \asqrt[10] , n18018);
  not g29701 (n_12038, n18019);
  and g29702 (n18020, n_11593, n_12038);
  not g29703 (n_12039, n18017);
  not g29704 (n_12040, n18020);
  and g29705 (n18021, n_12039, n_12040);
  and g29706 (n18022, n_4754, n_12035);
  and g29707 (n18023, n_12036, n18022);
  not g29708 (n_12041, n18021);
  not g29709 (n_12042, n18023);
  and g29710 (n18024, n_12041, n_12042);
  not g29711 (n_12043, n18014);
  not g29712 (n_12044, n18024);
  and g29713 (n18025, n_12043, n_12044);
  not g29714 (n_12045, n18025);
  and g29715 (n18026, \asqrt[33] , n_12045);
  and g29719 (n18030, n_11603, n_11602);
  and g29720 (n18031, \asqrt[10] , n18030);
  not g29721 (n_12046, n18031);
  and g29722 (n18032, n_11601, n_12046);
  not g29723 (n_12047, n18029);
  not g29724 (n_12048, n18032);
  and g29725 (n18033, n_12047, n_12048);
  and g29726 (n18034, n_4482, n_12043);
  and g29727 (n18035, n_12044, n18034);
  not g29728 (n_12049, n18033);
  not g29729 (n_12050, n18035);
  and g29730 (n18036, n_12049, n_12050);
  not g29731 (n_12051, n18026);
  not g29732 (n_12052, n18036);
  and g29733 (n18037, n_12051, n_12052);
  not g29734 (n_12053, n18037);
  and g29735 (n18038, \asqrt[34] , n_12053);
  and g29739 (n18042, n_11611, n_11610);
  and g29740 (n18043, \asqrt[10] , n18042);
  not g29741 (n_12054, n18043);
  and g29742 (n18044, n_11609, n_12054);
  not g29743 (n_12055, n18041);
  not g29744 (n_12056, n18044);
  and g29745 (n18045, n_12055, n_12056);
  and g29746 (n18046, n_4218, n_12051);
  and g29747 (n18047, n_12052, n18046);
  not g29748 (n_12057, n18045);
  not g29749 (n_12058, n18047);
  and g29750 (n18048, n_12057, n_12058);
  not g29751 (n_12059, n18038);
  not g29752 (n_12060, n18048);
  and g29753 (n18049, n_12059, n_12060);
  not g29754 (n_12061, n18049);
  and g29755 (n18050, \asqrt[35] , n_12061);
  and g29759 (n18054, n_11619, n_11618);
  and g29760 (n18055, \asqrt[10] , n18054);
  not g29761 (n_12062, n18055);
  and g29762 (n18056, n_11617, n_12062);
  not g29763 (n_12063, n18053);
  not g29764 (n_12064, n18056);
  and g29765 (n18057, n_12063, n_12064);
  and g29766 (n18058, n_3962, n_12059);
  and g29767 (n18059, n_12060, n18058);
  not g29768 (n_12065, n18057);
  not g29769 (n_12066, n18059);
  and g29770 (n18060, n_12065, n_12066);
  not g29771 (n_12067, n18050);
  not g29772 (n_12068, n18060);
  and g29773 (n18061, n_12067, n_12068);
  not g29774 (n_12069, n18061);
  and g29775 (n18062, \asqrt[36] , n_12069);
  and g29779 (n18066, n_11627, n_11626);
  and g29780 (n18067, \asqrt[10] , n18066);
  not g29781 (n_12070, n18067);
  and g29782 (n18068, n_11625, n_12070);
  not g29783 (n_12071, n18065);
  not g29784 (n_12072, n18068);
  and g29785 (n18069, n_12071, n_12072);
  and g29786 (n18070, n_3714, n_12067);
  and g29787 (n18071, n_12068, n18070);
  not g29788 (n_12073, n18069);
  not g29789 (n_12074, n18071);
  and g29790 (n18072, n_12073, n_12074);
  not g29791 (n_12075, n18062);
  not g29792 (n_12076, n18072);
  and g29793 (n18073, n_12075, n_12076);
  not g29794 (n_12077, n18073);
  and g29795 (n18074, \asqrt[37] , n_12077);
  and g29799 (n18078, n_11635, n_11634);
  and g29800 (n18079, \asqrt[10] , n18078);
  not g29801 (n_12078, n18079);
  and g29802 (n18080, n_11633, n_12078);
  not g29803 (n_12079, n18077);
  not g29804 (n_12080, n18080);
  and g29805 (n18081, n_12079, n_12080);
  and g29806 (n18082, n_3474, n_12075);
  and g29807 (n18083, n_12076, n18082);
  not g29808 (n_12081, n18081);
  not g29809 (n_12082, n18083);
  and g29810 (n18084, n_12081, n_12082);
  not g29811 (n_12083, n18074);
  not g29812 (n_12084, n18084);
  and g29813 (n18085, n_12083, n_12084);
  not g29814 (n_12085, n18085);
  and g29815 (n18086, \asqrt[38] , n_12085);
  and g29819 (n18090, n_11643, n_11642);
  and g29820 (n18091, \asqrt[10] , n18090);
  not g29821 (n_12086, n18091);
  and g29822 (n18092, n_11641, n_12086);
  not g29823 (n_12087, n18089);
  not g29824 (n_12088, n18092);
  and g29825 (n18093, n_12087, n_12088);
  and g29826 (n18094, n_3242, n_12083);
  and g29827 (n18095, n_12084, n18094);
  not g29828 (n_12089, n18093);
  not g29829 (n_12090, n18095);
  and g29830 (n18096, n_12089, n_12090);
  not g29831 (n_12091, n18086);
  not g29832 (n_12092, n18096);
  and g29833 (n18097, n_12091, n_12092);
  not g29834 (n_12093, n18097);
  and g29835 (n18098, \asqrt[39] , n_12093);
  and g29839 (n18102, n_11651, n_11650);
  and g29840 (n18103, \asqrt[10] , n18102);
  not g29841 (n_12094, n18103);
  and g29842 (n18104, n_11649, n_12094);
  not g29843 (n_12095, n18101);
  not g29844 (n_12096, n18104);
  and g29845 (n18105, n_12095, n_12096);
  and g29846 (n18106, n_3018, n_12091);
  and g29847 (n18107, n_12092, n18106);
  not g29848 (n_12097, n18105);
  not g29849 (n_12098, n18107);
  and g29850 (n18108, n_12097, n_12098);
  not g29851 (n_12099, n18098);
  not g29852 (n_12100, n18108);
  and g29853 (n18109, n_12099, n_12100);
  not g29854 (n_12101, n18109);
  and g29855 (n18110, \asqrt[40] , n_12101);
  and g29859 (n18114, n_11659, n_11658);
  and g29860 (n18115, \asqrt[10] , n18114);
  not g29861 (n_12102, n18115);
  and g29862 (n18116, n_11657, n_12102);
  not g29863 (n_12103, n18113);
  not g29864 (n_12104, n18116);
  and g29865 (n18117, n_12103, n_12104);
  and g29866 (n18118, n_2802, n_12099);
  and g29867 (n18119, n_12100, n18118);
  not g29868 (n_12105, n18117);
  not g29869 (n_12106, n18119);
  and g29870 (n18120, n_12105, n_12106);
  not g29871 (n_12107, n18110);
  not g29872 (n_12108, n18120);
  and g29873 (n18121, n_12107, n_12108);
  not g29874 (n_12109, n18121);
  and g29875 (n18122, \asqrt[41] , n_12109);
  and g29879 (n18126, n_11667, n_11666);
  and g29880 (n18127, \asqrt[10] , n18126);
  not g29881 (n_12110, n18127);
  and g29882 (n18128, n_11665, n_12110);
  not g29883 (n_12111, n18125);
  not g29884 (n_12112, n18128);
  and g29885 (n18129, n_12111, n_12112);
  and g29886 (n18130, n_2594, n_12107);
  and g29887 (n18131, n_12108, n18130);
  not g29888 (n_12113, n18129);
  not g29889 (n_12114, n18131);
  and g29890 (n18132, n_12113, n_12114);
  not g29891 (n_12115, n18122);
  not g29892 (n_12116, n18132);
  and g29893 (n18133, n_12115, n_12116);
  not g29894 (n_12117, n18133);
  and g29895 (n18134, \asqrt[42] , n_12117);
  and g29899 (n18138, n_11675, n_11674);
  and g29900 (n18139, \asqrt[10] , n18138);
  not g29901 (n_12118, n18139);
  and g29902 (n18140, n_11673, n_12118);
  not g29903 (n_12119, n18137);
  not g29904 (n_12120, n18140);
  and g29905 (n18141, n_12119, n_12120);
  and g29906 (n18142, n_2394, n_12115);
  and g29907 (n18143, n_12116, n18142);
  not g29908 (n_12121, n18141);
  not g29909 (n_12122, n18143);
  and g29910 (n18144, n_12121, n_12122);
  not g29911 (n_12123, n18134);
  not g29912 (n_12124, n18144);
  and g29913 (n18145, n_12123, n_12124);
  not g29914 (n_12125, n18145);
  and g29915 (n18146, \asqrt[43] , n_12125);
  and g29919 (n18150, n_11683, n_11682);
  and g29920 (n18151, \asqrt[10] , n18150);
  not g29921 (n_12126, n18151);
  and g29922 (n18152, n_11681, n_12126);
  not g29923 (n_12127, n18149);
  not g29924 (n_12128, n18152);
  and g29925 (n18153, n_12127, n_12128);
  and g29926 (n18154, n_2202, n_12123);
  and g29927 (n18155, n_12124, n18154);
  not g29928 (n_12129, n18153);
  not g29929 (n_12130, n18155);
  and g29930 (n18156, n_12129, n_12130);
  not g29931 (n_12131, n18146);
  not g29932 (n_12132, n18156);
  and g29933 (n18157, n_12131, n_12132);
  not g29934 (n_12133, n18157);
  and g29935 (n18158, \asqrt[44] , n_12133);
  and g29939 (n18162, n_11691, n_11690);
  and g29940 (n18163, \asqrt[10] , n18162);
  not g29941 (n_12134, n18163);
  and g29942 (n18164, n_11689, n_12134);
  not g29943 (n_12135, n18161);
  not g29944 (n_12136, n18164);
  and g29945 (n18165, n_12135, n_12136);
  and g29946 (n18166, n_2018, n_12131);
  and g29947 (n18167, n_12132, n18166);
  not g29948 (n_12137, n18165);
  not g29949 (n_12138, n18167);
  and g29950 (n18168, n_12137, n_12138);
  not g29951 (n_12139, n18158);
  not g29952 (n_12140, n18168);
  and g29953 (n18169, n_12139, n_12140);
  not g29954 (n_12141, n18169);
  and g29955 (n18170, \asqrt[45] , n_12141);
  and g29959 (n18174, n_11699, n_11698);
  and g29960 (n18175, \asqrt[10] , n18174);
  not g29961 (n_12142, n18175);
  and g29962 (n18176, n_11697, n_12142);
  not g29963 (n_12143, n18173);
  not g29964 (n_12144, n18176);
  and g29965 (n18177, n_12143, n_12144);
  and g29966 (n18178, n_1842, n_12139);
  and g29967 (n18179, n_12140, n18178);
  not g29968 (n_12145, n18177);
  not g29969 (n_12146, n18179);
  and g29970 (n18180, n_12145, n_12146);
  not g29971 (n_12147, n18170);
  not g29972 (n_12148, n18180);
  and g29973 (n18181, n_12147, n_12148);
  not g29974 (n_12149, n18181);
  and g29975 (n18182, \asqrt[46] , n_12149);
  and g29979 (n18186, n_11707, n_11706);
  and g29980 (n18187, \asqrt[10] , n18186);
  not g29981 (n_12150, n18187);
  and g29982 (n18188, n_11705, n_12150);
  not g29983 (n_12151, n18185);
  not g29984 (n_12152, n18188);
  and g29985 (n18189, n_12151, n_12152);
  and g29986 (n18190, n_1674, n_12147);
  and g29987 (n18191, n_12148, n18190);
  not g29988 (n_12153, n18189);
  not g29989 (n_12154, n18191);
  and g29990 (n18192, n_12153, n_12154);
  not g29991 (n_12155, n18182);
  not g29992 (n_12156, n18192);
  and g29993 (n18193, n_12155, n_12156);
  not g29994 (n_12157, n18193);
  and g29995 (n18194, \asqrt[47] , n_12157);
  and g29999 (n18198, n_11715, n_11714);
  and g30000 (n18199, \asqrt[10] , n18198);
  not g30001 (n_12158, n18199);
  and g30002 (n18200, n_11713, n_12158);
  not g30003 (n_12159, n18197);
  not g30004 (n_12160, n18200);
  and g30005 (n18201, n_12159, n_12160);
  and g30006 (n18202, n_1514, n_12155);
  and g30007 (n18203, n_12156, n18202);
  not g30008 (n_12161, n18201);
  not g30009 (n_12162, n18203);
  and g30010 (n18204, n_12161, n_12162);
  not g30011 (n_12163, n18194);
  not g30012 (n_12164, n18204);
  and g30013 (n18205, n_12163, n_12164);
  not g30014 (n_12165, n18205);
  and g30015 (n18206, \asqrt[48] , n_12165);
  and g30019 (n18210, n_11723, n_11722);
  and g30020 (n18211, \asqrt[10] , n18210);
  not g30021 (n_12166, n18211);
  and g30022 (n18212, n_11721, n_12166);
  not g30023 (n_12167, n18209);
  not g30024 (n_12168, n18212);
  and g30025 (n18213, n_12167, n_12168);
  and g30026 (n18214, n_1362, n_12163);
  and g30027 (n18215, n_12164, n18214);
  not g30028 (n_12169, n18213);
  not g30029 (n_12170, n18215);
  and g30030 (n18216, n_12169, n_12170);
  not g30031 (n_12171, n18206);
  not g30032 (n_12172, n18216);
  and g30033 (n18217, n_12171, n_12172);
  not g30034 (n_12173, n18217);
  and g30035 (n18218, \asqrt[49] , n_12173);
  and g30039 (n18222, n_11731, n_11730);
  and g30040 (n18223, \asqrt[10] , n18222);
  not g30041 (n_12174, n18223);
  and g30042 (n18224, n_11729, n_12174);
  not g30043 (n_12175, n18221);
  not g30044 (n_12176, n18224);
  and g30045 (n18225, n_12175, n_12176);
  and g30046 (n18226, n_1218, n_12171);
  and g30047 (n18227, n_12172, n18226);
  not g30048 (n_12177, n18225);
  not g30049 (n_12178, n18227);
  and g30050 (n18228, n_12177, n_12178);
  not g30051 (n_12179, n18218);
  not g30052 (n_12180, n18228);
  and g30053 (n18229, n_12179, n_12180);
  not g30054 (n_12181, n18229);
  and g30055 (n18230, \asqrt[50] , n_12181);
  and g30059 (n18234, n_11739, n_11738);
  and g30060 (n18235, \asqrt[10] , n18234);
  not g30061 (n_12182, n18235);
  and g30062 (n18236, n_11737, n_12182);
  not g30063 (n_12183, n18233);
  not g30064 (n_12184, n18236);
  and g30065 (n18237, n_12183, n_12184);
  and g30066 (n18238, n_1082, n_12179);
  and g30067 (n18239, n_12180, n18238);
  not g30068 (n_12185, n18237);
  not g30069 (n_12186, n18239);
  and g30070 (n18240, n_12185, n_12186);
  not g30071 (n_12187, n18230);
  not g30072 (n_12188, n18240);
  and g30073 (n18241, n_12187, n_12188);
  not g30074 (n_12189, n18241);
  and g30075 (n18242, \asqrt[51] , n_12189);
  and g30079 (n18246, n_11747, n_11746);
  and g30080 (n18247, \asqrt[10] , n18246);
  not g30081 (n_12190, n18247);
  and g30082 (n18248, n_11745, n_12190);
  not g30083 (n_12191, n18245);
  not g30084 (n_12192, n18248);
  and g30085 (n18249, n_12191, n_12192);
  and g30086 (n18250, n_954, n_12187);
  and g30087 (n18251, n_12188, n18250);
  not g30088 (n_12193, n18249);
  not g30089 (n_12194, n18251);
  and g30090 (n18252, n_12193, n_12194);
  not g30091 (n_12195, n18242);
  not g30092 (n_12196, n18252);
  and g30093 (n18253, n_12195, n_12196);
  not g30094 (n_12197, n18253);
  and g30095 (n18254, \asqrt[52] , n_12197);
  and g30099 (n18258, n_11755, n_11754);
  and g30100 (n18259, \asqrt[10] , n18258);
  not g30101 (n_12198, n18259);
  and g30102 (n18260, n_11753, n_12198);
  not g30103 (n_12199, n18257);
  not g30104 (n_12200, n18260);
  and g30105 (n18261, n_12199, n_12200);
  and g30106 (n18262, n_834, n_12195);
  and g30107 (n18263, n_12196, n18262);
  not g30108 (n_12201, n18261);
  not g30109 (n_12202, n18263);
  and g30110 (n18264, n_12201, n_12202);
  not g30111 (n_12203, n18254);
  not g30112 (n_12204, n18264);
  and g30113 (n18265, n_12203, n_12204);
  not g30114 (n_12205, n18265);
  and g30115 (n18266, \asqrt[53] , n_12205);
  and g30119 (n18270, n_11763, n_11762);
  and g30120 (n18271, \asqrt[10] , n18270);
  not g30121 (n_12206, n18271);
  and g30122 (n18272, n_11761, n_12206);
  not g30123 (n_12207, n18269);
  not g30124 (n_12208, n18272);
  and g30125 (n18273, n_12207, n_12208);
  and g30126 (n18274, n_722, n_12203);
  and g30127 (n18275, n_12204, n18274);
  not g30128 (n_12209, n18273);
  not g30129 (n_12210, n18275);
  and g30130 (n18276, n_12209, n_12210);
  not g30131 (n_12211, n18266);
  not g30132 (n_12212, n18276);
  and g30133 (n18277, n_12211, n_12212);
  not g30134 (n_12213, n18277);
  and g30135 (n18278, \asqrt[54] , n_12213);
  and g30139 (n18282, n_11771, n_11770);
  and g30140 (n18283, \asqrt[10] , n18282);
  not g30141 (n_12214, n18283);
  and g30142 (n18284, n_11769, n_12214);
  not g30143 (n_12215, n18281);
  not g30144 (n_12216, n18284);
  and g30145 (n18285, n_12215, n_12216);
  and g30146 (n18286, n_618, n_12211);
  and g30147 (n18287, n_12212, n18286);
  not g30148 (n_12217, n18285);
  not g30149 (n_12218, n18287);
  and g30150 (n18288, n_12217, n_12218);
  not g30151 (n_12219, n18278);
  not g30152 (n_12220, n18288);
  and g30153 (n18289, n_12219, n_12220);
  not g30154 (n_12221, n18289);
  and g30155 (n18290, \asqrt[55] , n_12221);
  and g30156 (n18291, n_522, n_12219);
  and g30157 (n18292, n_12220, n18291);
  and g30161 (n18296, n_11779, n_11777);
  and g30162 (n18297, \asqrt[10] , n18296);
  not g30163 (n_12222, n18297);
  and g30164 (n18298, n_11778, n_12222);
  not g30165 (n_12223, n18295);
  not g30166 (n_12224, n18298);
  and g30167 (n18299, n_12223, n_12224);
  not g30168 (n_12225, n18292);
  not g30169 (n_12226, n18299);
  and g30170 (n18300, n_12225, n_12226);
  not g30171 (n_12227, n18290);
  not g30172 (n_12228, n18300);
  and g30173 (n18301, n_12227, n_12228);
  not g30174 (n_12229, n18301);
  and g30175 (n18302, \asqrt[56] , n_12229);
  and g30179 (n18306, n_11787, n_11786);
  and g30180 (n18307, \asqrt[10] , n18306);
  not g30181 (n_12230, n18307);
  and g30182 (n18308, n_11785, n_12230);
  not g30183 (n_12231, n18305);
  not g30184 (n_12232, n18308);
  and g30185 (n18309, n_12231, n_12232);
  and g30186 (n18310, n_434, n_12227);
  and g30187 (n18311, n_12228, n18310);
  not g30188 (n_12233, n18309);
  not g30189 (n_12234, n18311);
  and g30190 (n18312, n_12233, n_12234);
  not g30191 (n_12235, n18302);
  not g30192 (n_12236, n18312);
  and g30193 (n18313, n_12235, n_12236);
  not g30194 (n_12237, n18313);
  and g30195 (n18314, \asqrt[57] , n_12237);
  and g30199 (n18318, n_11795, n_11794);
  and g30200 (n18319, \asqrt[10] , n18318);
  not g30201 (n_12238, n18319);
  and g30202 (n18320, n_11793, n_12238);
  not g30203 (n_12239, n18317);
  not g30204 (n_12240, n18320);
  and g30205 (n18321, n_12239, n_12240);
  and g30206 (n18322, n_354, n_12235);
  and g30207 (n18323, n_12236, n18322);
  not g30208 (n_12241, n18321);
  not g30209 (n_12242, n18323);
  and g30210 (n18324, n_12241, n_12242);
  not g30211 (n_12243, n18314);
  not g30212 (n_12244, n18324);
  and g30213 (n18325, n_12243, n_12244);
  not g30214 (n_12245, n18325);
  and g30215 (n18326, \asqrt[58] , n_12245);
  and g30219 (n18330, n_11803, n_11802);
  and g30220 (n18331, \asqrt[10] , n18330);
  not g30221 (n_12246, n18331);
  and g30222 (n18332, n_11801, n_12246);
  not g30223 (n_12247, n18329);
  not g30224 (n_12248, n18332);
  and g30225 (n18333, n_12247, n_12248);
  and g30226 (n18334, n_282, n_12243);
  and g30227 (n18335, n_12244, n18334);
  not g30228 (n_12249, n18333);
  not g30229 (n_12250, n18335);
  and g30230 (n18336, n_12249, n_12250);
  not g30231 (n_12251, n18326);
  not g30232 (n_12252, n18336);
  and g30233 (n18337, n_12251, n_12252);
  not g30234 (n_12253, n18337);
  and g30235 (n18338, \asqrt[59] , n_12253);
  and g30239 (n18342, n_11811, n_11810);
  and g30240 (n18343, \asqrt[10] , n18342);
  not g30241 (n_12254, n18343);
  and g30242 (n18344, n_11809, n_12254);
  not g30243 (n_12255, n18341);
  not g30244 (n_12256, n18344);
  and g30245 (n18345, n_12255, n_12256);
  and g30246 (n18346, n_218, n_12251);
  and g30247 (n18347, n_12252, n18346);
  not g30248 (n_12257, n18345);
  not g30249 (n_12258, n18347);
  and g30250 (n18348, n_12257, n_12258);
  not g30251 (n_12259, n18338);
  not g30252 (n_12260, n18348);
  and g30253 (n18349, n_12259, n_12260);
  not g30254 (n_12261, n18349);
  and g30255 (n18350, \asqrt[60] , n_12261);
  and g30259 (n18354, n_11819, n_11818);
  and g30260 (n18355, \asqrt[10] , n18354);
  not g30261 (n_12262, n18355);
  and g30262 (n18356, n_11817, n_12262);
  not g30263 (n_12263, n18353);
  not g30264 (n_12264, n18356);
  and g30265 (n18357, n_12263, n_12264);
  and g30266 (n18358, n_162, n_12259);
  and g30267 (n18359, n_12260, n18358);
  not g30268 (n_12265, n18357);
  not g30269 (n_12266, n18359);
  and g30270 (n18360, n_12265, n_12266);
  not g30271 (n_12267, n18350);
  not g30272 (n_12268, n18360);
  and g30273 (n18361, n_12267, n_12268);
  not g30274 (n_12269, n18361);
  and g30275 (n18362, \asqrt[61] , n_12269);
  and g30279 (n18366, n_11827, n_11826);
  and g30280 (n18367, \asqrt[10] , n18366);
  not g30281 (n_12270, n18367);
  and g30282 (n18368, n_11825, n_12270);
  not g30283 (n_12271, n18365);
  not g30284 (n_12272, n18368);
  and g30285 (n18369, n_12271, n_12272);
  and g30286 (n18370, n_115, n_12267);
  and g30287 (n18371, n_12268, n18370);
  not g30288 (n_12273, n18369);
  not g30289 (n_12274, n18371);
  and g30290 (n18372, n_12273, n_12274);
  not g30291 (n_12275, n18362);
  not g30292 (n_12276, n18372);
  and g30293 (n18373, n_12275, n_12276);
  not g30294 (n_12277, n18373);
  and g30295 (n18374, \asqrt[62] , n_12277);
  and g30299 (n18378, n_11835, n_11834);
  and g30300 (n18379, \asqrt[10] , n18378);
  not g30301 (n_12278, n18379);
  and g30302 (n18380, n_11833, n_12278);
  not g30303 (n_12279, n18377);
  not g30304 (n_12280, n18380);
  and g30305 (n18381, n_12279, n_12280);
  and g30306 (n18382, n_76, n_12275);
  and g30307 (n18383, n_12276, n18382);
  not g30308 (n_12281, n18381);
  not g30309 (n_12282, n18383);
  and g30310 (n18384, n_12281, n_12282);
  not g30311 (n_12283, n18374);
  not g30312 (n_12284, n18384);
  and g30313 (n18385, n_12283, n_12284);
  and g30317 (n18389, n_11843, n_11842);
  and g30318 (n18390, \asqrt[10] , n18389);
  not g30319 (n_12285, n18390);
  and g30320 (n18391, n_11841, n_12285);
  not g30321 (n_12286, n18388);
  not g30322 (n_12287, n18391);
  and g30323 (n18392, n_12286, n_12287);
  and g30324 (n18393, n_11850, n_11849);
  and g30325 (n18394, \asqrt[10] , n18393);
  not g30328 (n_12289, n18392);
  not g30330 (n_12290, n18385);
  not g30332 (n_12291, n18397);
  and g30333 (n18398, n_21, n_12291);
  and g30334 (n18399, n_12283, n18392);
  and g30335 (n18400, n_12284, n18399);
  and g30336 (n18401, n_11849, \asqrt[10] );
  not g30337 (n_12292, n18401);
  and g30338 (n18402, n17729, n_12292);
  not g30339 (n_12293, n18393);
  and g30340 (n18403, \asqrt[63] , n_12293);
  not g30341 (n_12294, n18402);
  and g30342 (n18404, n_12294, n18403);
  not g30348 (n_12295, n18404);
  not g30349 (n_12296, n18409);
  not g30351 (n_12297, n18400);
  and g30355 (n18413, \a[18] , \asqrt[9] );
  not g30356 (n_12302, \a[16] );
  not g30357 (n_12303, \a[17] );
  and g30358 (n18414, n_12302, n_12303);
  and g30359 (n18415, n_11862, n18414);
  not g30360 (n_12304, n18413);
  not g30361 (n_12305, n18415);
  and g30362 (n18416, n_12304, n_12305);
  not g30363 (n_12306, n18416);
  and g30364 (n18417, \asqrt[10] , n_12306);
  and g30370 (n18423, n_11862, \asqrt[9] );
  not g30371 (n_12307, n18423);
  and g30372 (n18424, \a[19] , n_12307);
  and g30373 (n18425, n17758, \asqrt[9] );
  not g30374 (n_12308, n18424);
  not g30375 (n_12309, n18425);
  and g30376 (n18426, n_12308, n_12309);
  not g30377 (n_12310, n18422);
  and g30378 (n18427, n_12310, n18426);
  not g30379 (n_12311, n18417);
  not g30380 (n_12312, n18427);
  and g30381 (n18428, n_12311, n_12312);
  not g30382 (n_12313, n18428);
  and g30383 (n18429, \asqrt[11] , n_12313);
  not g30384 (n_12314, \asqrt[11] );
  and g30385 (n18430, n_12314, n_12311);
  and g30386 (n18431, n_12312, n18430);
  not g30390 (n_12315, n18398);
  not g30392 (n_12316, n18435);
  and g30393 (n18436, n_12309, n_12316);
  not g30394 (n_12317, n18436);
  and g30395 (n18437, \a[20] , n_12317);
  and g30396 (n18438, n_11430, n_12316);
  and g30397 (n18439, n_12309, n18438);
  not g30398 (n_12318, n18437);
  not g30399 (n_12319, n18439);
  and g30400 (n18440, n_12318, n_12319);
  not g30401 (n_12320, n18431);
  not g30402 (n_12321, n18440);
  and g30403 (n18441, n_12320, n_12321);
  not g30404 (n_12322, n18429);
  not g30405 (n_12323, n18441);
  and g30406 (n18442, n_12322, n_12323);
  not g30407 (n_12324, n18442);
  and g30408 (n18443, \asqrt[12] , n_12324);
  and g30409 (n18444, n_11871, n_11870);
  not g30410 (n_12325, n17770);
  and g30411 (n18445, n_12325, n18444);
  and g30412 (n18446, \asqrt[9] , n18445);
  and g30413 (n18447, \asqrt[9] , n18444);
  not g30414 (n_12326, n18447);
  and g30415 (n18448, n17770, n_12326);
  not g30416 (n_12327, n18446);
  not g30417 (n_12328, n18448);
  and g30418 (n18449, n_12327, n_12328);
  and g30419 (n18450, n_11874, n_12322);
  and g30420 (n18451, n_12323, n18450);
  not g30421 (n_12329, n18449);
  not g30422 (n_12330, n18451);
  and g30423 (n18452, n_12329, n_12330);
  not g30424 (n_12331, n18443);
  not g30425 (n_12332, n18452);
  and g30426 (n18453, n_12331, n_12332);
  not g30427 (n_12333, n18453);
  and g30428 (n18454, \asqrt[13] , n_12333);
  and g30432 (n18458, n_11882, n_11880);
  and g30433 (n18459, \asqrt[9] , n18458);
  not g30434 (n_12334, n18459);
  and g30435 (n18460, n_11881, n_12334);
  not g30436 (n_12335, n18457);
  not g30437 (n_12336, n18460);
  and g30438 (n18461, n_12335, n_12336);
  and g30439 (n18462, n_11442, n_12331);
  and g30440 (n18463, n_12332, n18462);
  not g30441 (n_12337, n18461);
  not g30442 (n_12338, n18463);
  and g30443 (n18464, n_12337, n_12338);
  not g30444 (n_12339, n18454);
  not g30445 (n_12340, n18464);
  and g30446 (n18465, n_12339, n_12340);
  not g30447 (n_12341, n18465);
  and g30448 (n18466, \asqrt[14] , n_12341);
  and g30452 (n18470, n_11891, n_11890);
  and g30453 (n18471, \asqrt[9] , n18470);
  not g30454 (n_12342, n18471);
  and g30455 (n18472, n_11889, n_12342);
  not g30456 (n_12343, n18469);
  not g30457 (n_12344, n18472);
  and g30458 (n18473, n_12343, n_12344);
  and g30459 (n18474, n_11018, n_12339);
  and g30460 (n18475, n_12340, n18474);
  not g30461 (n_12345, n18473);
  not g30462 (n_12346, n18475);
  and g30463 (n18476, n_12345, n_12346);
  not g30464 (n_12347, n18466);
  not g30465 (n_12348, n18476);
  and g30466 (n18477, n_12347, n_12348);
  not g30467 (n_12349, n18477);
  and g30468 (n18478, \asqrt[15] , n_12349);
  and g30472 (n18482, n_11899, n_11898);
  and g30473 (n18483, \asqrt[9] , n18482);
  not g30474 (n_12350, n18483);
  and g30475 (n18484, n_11897, n_12350);
  not g30476 (n_12351, n18481);
  not g30477 (n_12352, n18484);
  and g30478 (n18485, n_12351, n_12352);
  and g30479 (n18486, n_10602, n_12347);
  and g30480 (n18487, n_12348, n18486);
  not g30481 (n_12353, n18485);
  not g30482 (n_12354, n18487);
  and g30483 (n18488, n_12353, n_12354);
  not g30484 (n_12355, n18478);
  not g30485 (n_12356, n18488);
  and g30486 (n18489, n_12355, n_12356);
  not g30487 (n_12357, n18489);
  and g30488 (n18490, \asqrt[16] , n_12357);
  and g30492 (n18494, n_11907, n_11906);
  and g30493 (n18495, \asqrt[9] , n18494);
  not g30494 (n_12358, n18495);
  and g30495 (n18496, n_11905, n_12358);
  not g30496 (n_12359, n18493);
  not g30497 (n_12360, n18496);
  and g30498 (n18497, n_12359, n_12360);
  and g30499 (n18498, n_10194, n_12355);
  and g30500 (n18499, n_12356, n18498);
  not g30501 (n_12361, n18497);
  not g30502 (n_12362, n18499);
  and g30503 (n18500, n_12361, n_12362);
  not g30504 (n_12363, n18490);
  not g30505 (n_12364, n18500);
  and g30506 (n18501, n_12363, n_12364);
  not g30507 (n_12365, n18501);
  and g30508 (n18502, \asqrt[17] , n_12365);
  and g30512 (n18506, n_11915, n_11914);
  and g30513 (n18507, \asqrt[9] , n18506);
  not g30514 (n_12366, n18507);
  and g30515 (n18508, n_11913, n_12366);
  not g30516 (n_12367, n18505);
  not g30517 (n_12368, n18508);
  and g30518 (n18509, n_12367, n_12368);
  and g30519 (n18510, n_9794, n_12363);
  and g30520 (n18511, n_12364, n18510);
  not g30521 (n_12369, n18509);
  not g30522 (n_12370, n18511);
  and g30523 (n18512, n_12369, n_12370);
  not g30524 (n_12371, n18502);
  not g30525 (n_12372, n18512);
  and g30526 (n18513, n_12371, n_12372);
  not g30527 (n_12373, n18513);
  and g30528 (n18514, \asqrt[18] , n_12373);
  and g30532 (n18518, n_11923, n_11922);
  and g30533 (n18519, \asqrt[9] , n18518);
  not g30534 (n_12374, n18519);
  and g30535 (n18520, n_11921, n_12374);
  not g30536 (n_12375, n18517);
  not g30537 (n_12376, n18520);
  and g30538 (n18521, n_12375, n_12376);
  and g30539 (n18522, n_9402, n_12371);
  and g30540 (n18523, n_12372, n18522);
  not g30541 (n_12377, n18521);
  not g30542 (n_12378, n18523);
  and g30543 (n18524, n_12377, n_12378);
  not g30544 (n_12379, n18514);
  not g30545 (n_12380, n18524);
  and g30546 (n18525, n_12379, n_12380);
  not g30547 (n_12381, n18525);
  and g30548 (n18526, \asqrt[19] , n_12381);
  and g30552 (n18530, n_11931, n_11930);
  and g30553 (n18531, \asqrt[9] , n18530);
  not g30554 (n_12382, n18531);
  and g30555 (n18532, n_11929, n_12382);
  not g30556 (n_12383, n18529);
  not g30557 (n_12384, n18532);
  and g30558 (n18533, n_12383, n_12384);
  and g30559 (n18534, n_9018, n_12379);
  and g30560 (n18535, n_12380, n18534);
  not g30561 (n_12385, n18533);
  not g30562 (n_12386, n18535);
  and g30563 (n18536, n_12385, n_12386);
  not g30564 (n_12387, n18526);
  not g30565 (n_12388, n18536);
  and g30566 (n18537, n_12387, n_12388);
  not g30567 (n_12389, n18537);
  and g30568 (n18538, \asqrt[20] , n_12389);
  and g30572 (n18542, n_11939, n_11938);
  and g30573 (n18543, \asqrt[9] , n18542);
  not g30574 (n_12390, n18543);
  and g30575 (n18544, n_11937, n_12390);
  not g30576 (n_12391, n18541);
  not g30577 (n_12392, n18544);
  and g30578 (n18545, n_12391, n_12392);
  and g30579 (n18546, n_8642, n_12387);
  and g30580 (n18547, n_12388, n18546);
  not g30581 (n_12393, n18545);
  not g30582 (n_12394, n18547);
  and g30583 (n18548, n_12393, n_12394);
  not g30584 (n_12395, n18538);
  not g30585 (n_12396, n18548);
  and g30586 (n18549, n_12395, n_12396);
  not g30587 (n_12397, n18549);
  and g30588 (n18550, \asqrt[21] , n_12397);
  and g30592 (n18554, n_11947, n_11946);
  and g30593 (n18555, \asqrt[9] , n18554);
  not g30594 (n_12398, n18555);
  and g30595 (n18556, n_11945, n_12398);
  not g30596 (n_12399, n18553);
  not g30597 (n_12400, n18556);
  and g30598 (n18557, n_12399, n_12400);
  and g30599 (n18558, n_8274, n_12395);
  and g30600 (n18559, n_12396, n18558);
  not g30601 (n_12401, n18557);
  not g30602 (n_12402, n18559);
  and g30603 (n18560, n_12401, n_12402);
  not g30604 (n_12403, n18550);
  not g30605 (n_12404, n18560);
  and g30606 (n18561, n_12403, n_12404);
  not g30607 (n_12405, n18561);
  and g30608 (n18562, \asqrt[22] , n_12405);
  and g30612 (n18566, n_11955, n_11954);
  and g30613 (n18567, \asqrt[9] , n18566);
  not g30614 (n_12406, n18567);
  and g30615 (n18568, n_11953, n_12406);
  not g30616 (n_12407, n18565);
  not g30617 (n_12408, n18568);
  and g30618 (n18569, n_12407, n_12408);
  and g30619 (n18570, n_7914, n_12403);
  and g30620 (n18571, n_12404, n18570);
  not g30621 (n_12409, n18569);
  not g30622 (n_12410, n18571);
  and g30623 (n18572, n_12409, n_12410);
  not g30624 (n_12411, n18562);
  not g30625 (n_12412, n18572);
  and g30626 (n18573, n_12411, n_12412);
  not g30627 (n_12413, n18573);
  and g30628 (n18574, \asqrt[23] , n_12413);
  and g30632 (n18578, n_11963, n_11962);
  and g30633 (n18579, \asqrt[9] , n18578);
  not g30634 (n_12414, n18579);
  and g30635 (n18580, n_11961, n_12414);
  not g30636 (n_12415, n18577);
  not g30637 (n_12416, n18580);
  and g30638 (n18581, n_12415, n_12416);
  and g30639 (n18582, n_7562, n_12411);
  and g30640 (n18583, n_12412, n18582);
  not g30641 (n_12417, n18581);
  not g30642 (n_12418, n18583);
  and g30643 (n18584, n_12417, n_12418);
  not g30644 (n_12419, n18574);
  not g30645 (n_12420, n18584);
  and g30646 (n18585, n_12419, n_12420);
  not g30647 (n_12421, n18585);
  and g30648 (n18586, \asqrt[24] , n_12421);
  and g30652 (n18590, n_11971, n_11970);
  and g30653 (n18591, \asqrt[9] , n18590);
  not g30654 (n_12422, n18591);
  and g30655 (n18592, n_11969, n_12422);
  not g30656 (n_12423, n18589);
  not g30657 (n_12424, n18592);
  and g30658 (n18593, n_12423, n_12424);
  and g30659 (n18594, n_7218, n_12419);
  and g30660 (n18595, n_12420, n18594);
  not g30661 (n_12425, n18593);
  not g30662 (n_12426, n18595);
  and g30663 (n18596, n_12425, n_12426);
  not g30664 (n_12427, n18586);
  not g30665 (n_12428, n18596);
  and g30666 (n18597, n_12427, n_12428);
  not g30667 (n_12429, n18597);
  and g30668 (n18598, \asqrt[25] , n_12429);
  and g30672 (n18602, n_11979, n_11978);
  and g30673 (n18603, \asqrt[9] , n18602);
  not g30674 (n_12430, n18603);
  and g30675 (n18604, n_11977, n_12430);
  not g30676 (n_12431, n18601);
  not g30677 (n_12432, n18604);
  and g30678 (n18605, n_12431, n_12432);
  and g30679 (n18606, n_6882, n_12427);
  and g30680 (n18607, n_12428, n18606);
  not g30681 (n_12433, n18605);
  not g30682 (n_12434, n18607);
  and g30683 (n18608, n_12433, n_12434);
  not g30684 (n_12435, n18598);
  not g30685 (n_12436, n18608);
  and g30686 (n18609, n_12435, n_12436);
  not g30687 (n_12437, n18609);
  and g30688 (n18610, \asqrt[26] , n_12437);
  and g30692 (n18614, n_11987, n_11986);
  and g30693 (n18615, \asqrt[9] , n18614);
  not g30694 (n_12438, n18615);
  and g30695 (n18616, n_11985, n_12438);
  not g30696 (n_12439, n18613);
  not g30697 (n_12440, n18616);
  and g30698 (n18617, n_12439, n_12440);
  and g30699 (n18618, n_6554, n_12435);
  and g30700 (n18619, n_12436, n18618);
  not g30701 (n_12441, n18617);
  not g30702 (n_12442, n18619);
  and g30703 (n18620, n_12441, n_12442);
  not g30704 (n_12443, n18610);
  not g30705 (n_12444, n18620);
  and g30706 (n18621, n_12443, n_12444);
  not g30707 (n_12445, n18621);
  and g30708 (n18622, \asqrt[27] , n_12445);
  and g30712 (n18626, n_11995, n_11994);
  and g30713 (n18627, \asqrt[9] , n18626);
  not g30714 (n_12446, n18627);
  and g30715 (n18628, n_11993, n_12446);
  not g30716 (n_12447, n18625);
  not g30717 (n_12448, n18628);
  and g30718 (n18629, n_12447, n_12448);
  and g30719 (n18630, n_6234, n_12443);
  and g30720 (n18631, n_12444, n18630);
  not g30721 (n_12449, n18629);
  not g30722 (n_12450, n18631);
  and g30723 (n18632, n_12449, n_12450);
  not g30724 (n_12451, n18622);
  not g30725 (n_12452, n18632);
  and g30726 (n18633, n_12451, n_12452);
  not g30727 (n_12453, n18633);
  and g30728 (n18634, \asqrt[28] , n_12453);
  and g30732 (n18638, n_12003, n_12002);
  and g30733 (n18639, \asqrt[9] , n18638);
  not g30734 (n_12454, n18639);
  and g30735 (n18640, n_12001, n_12454);
  not g30736 (n_12455, n18637);
  not g30737 (n_12456, n18640);
  and g30738 (n18641, n_12455, n_12456);
  and g30739 (n18642, n_5922, n_12451);
  and g30740 (n18643, n_12452, n18642);
  not g30741 (n_12457, n18641);
  not g30742 (n_12458, n18643);
  and g30743 (n18644, n_12457, n_12458);
  not g30744 (n_12459, n18634);
  not g30745 (n_12460, n18644);
  and g30746 (n18645, n_12459, n_12460);
  not g30747 (n_12461, n18645);
  and g30748 (n18646, \asqrt[29] , n_12461);
  and g30752 (n18650, n_12011, n_12010);
  and g30753 (n18651, \asqrt[9] , n18650);
  not g30754 (n_12462, n18651);
  and g30755 (n18652, n_12009, n_12462);
  not g30756 (n_12463, n18649);
  not g30757 (n_12464, n18652);
  and g30758 (n18653, n_12463, n_12464);
  and g30759 (n18654, n_5618, n_12459);
  and g30760 (n18655, n_12460, n18654);
  not g30761 (n_12465, n18653);
  not g30762 (n_12466, n18655);
  and g30763 (n18656, n_12465, n_12466);
  not g30764 (n_12467, n18646);
  not g30765 (n_12468, n18656);
  and g30766 (n18657, n_12467, n_12468);
  not g30767 (n_12469, n18657);
  and g30768 (n18658, \asqrt[30] , n_12469);
  and g30772 (n18662, n_12019, n_12018);
  and g30773 (n18663, \asqrt[9] , n18662);
  not g30774 (n_12470, n18663);
  and g30775 (n18664, n_12017, n_12470);
  not g30776 (n_12471, n18661);
  not g30777 (n_12472, n18664);
  and g30778 (n18665, n_12471, n_12472);
  and g30779 (n18666, n_5322, n_12467);
  and g30780 (n18667, n_12468, n18666);
  not g30781 (n_12473, n18665);
  not g30782 (n_12474, n18667);
  and g30783 (n18668, n_12473, n_12474);
  not g30784 (n_12475, n18658);
  not g30785 (n_12476, n18668);
  and g30786 (n18669, n_12475, n_12476);
  not g30787 (n_12477, n18669);
  and g30788 (n18670, \asqrt[31] , n_12477);
  and g30792 (n18674, n_12027, n_12026);
  and g30793 (n18675, \asqrt[9] , n18674);
  not g30794 (n_12478, n18675);
  and g30795 (n18676, n_12025, n_12478);
  not g30796 (n_12479, n18673);
  not g30797 (n_12480, n18676);
  and g30798 (n18677, n_12479, n_12480);
  and g30799 (n18678, n_5034, n_12475);
  and g30800 (n18679, n_12476, n18678);
  not g30801 (n_12481, n18677);
  not g30802 (n_12482, n18679);
  and g30803 (n18680, n_12481, n_12482);
  not g30804 (n_12483, n18670);
  not g30805 (n_12484, n18680);
  and g30806 (n18681, n_12483, n_12484);
  not g30807 (n_12485, n18681);
  and g30808 (n18682, \asqrt[32] , n_12485);
  and g30812 (n18686, n_12035, n_12034);
  and g30813 (n18687, \asqrt[9] , n18686);
  not g30814 (n_12486, n18687);
  and g30815 (n18688, n_12033, n_12486);
  not g30816 (n_12487, n18685);
  not g30817 (n_12488, n18688);
  and g30818 (n18689, n_12487, n_12488);
  and g30819 (n18690, n_4754, n_12483);
  and g30820 (n18691, n_12484, n18690);
  not g30821 (n_12489, n18689);
  not g30822 (n_12490, n18691);
  and g30823 (n18692, n_12489, n_12490);
  not g30824 (n_12491, n18682);
  not g30825 (n_12492, n18692);
  and g30826 (n18693, n_12491, n_12492);
  not g30827 (n_12493, n18693);
  and g30828 (n18694, \asqrt[33] , n_12493);
  and g30832 (n18698, n_12043, n_12042);
  and g30833 (n18699, \asqrt[9] , n18698);
  not g30834 (n_12494, n18699);
  and g30835 (n18700, n_12041, n_12494);
  not g30836 (n_12495, n18697);
  not g30837 (n_12496, n18700);
  and g30838 (n18701, n_12495, n_12496);
  and g30839 (n18702, n_4482, n_12491);
  and g30840 (n18703, n_12492, n18702);
  not g30841 (n_12497, n18701);
  not g30842 (n_12498, n18703);
  and g30843 (n18704, n_12497, n_12498);
  not g30844 (n_12499, n18694);
  not g30845 (n_12500, n18704);
  and g30846 (n18705, n_12499, n_12500);
  not g30847 (n_12501, n18705);
  and g30848 (n18706, \asqrt[34] , n_12501);
  and g30852 (n18710, n_12051, n_12050);
  and g30853 (n18711, \asqrt[9] , n18710);
  not g30854 (n_12502, n18711);
  and g30855 (n18712, n_12049, n_12502);
  not g30856 (n_12503, n18709);
  not g30857 (n_12504, n18712);
  and g30858 (n18713, n_12503, n_12504);
  and g30859 (n18714, n_4218, n_12499);
  and g30860 (n18715, n_12500, n18714);
  not g30861 (n_12505, n18713);
  not g30862 (n_12506, n18715);
  and g30863 (n18716, n_12505, n_12506);
  not g30864 (n_12507, n18706);
  not g30865 (n_12508, n18716);
  and g30866 (n18717, n_12507, n_12508);
  not g30867 (n_12509, n18717);
  and g30868 (n18718, \asqrt[35] , n_12509);
  and g30872 (n18722, n_12059, n_12058);
  and g30873 (n18723, \asqrt[9] , n18722);
  not g30874 (n_12510, n18723);
  and g30875 (n18724, n_12057, n_12510);
  not g30876 (n_12511, n18721);
  not g30877 (n_12512, n18724);
  and g30878 (n18725, n_12511, n_12512);
  and g30879 (n18726, n_3962, n_12507);
  and g30880 (n18727, n_12508, n18726);
  not g30881 (n_12513, n18725);
  not g30882 (n_12514, n18727);
  and g30883 (n18728, n_12513, n_12514);
  not g30884 (n_12515, n18718);
  not g30885 (n_12516, n18728);
  and g30886 (n18729, n_12515, n_12516);
  not g30887 (n_12517, n18729);
  and g30888 (n18730, \asqrt[36] , n_12517);
  and g30892 (n18734, n_12067, n_12066);
  and g30893 (n18735, \asqrt[9] , n18734);
  not g30894 (n_12518, n18735);
  and g30895 (n18736, n_12065, n_12518);
  not g30896 (n_12519, n18733);
  not g30897 (n_12520, n18736);
  and g30898 (n18737, n_12519, n_12520);
  and g30899 (n18738, n_3714, n_12515);
  and g30900 (n18739, n_12516, n18738);
  not g30901 (n_12521, n18737);
  not g30902 (n_12522, n18739);
  and g30903 (n18740, n_12521, n_12522);
  not g30904 (n_12523, n18730);
  not g30905 (n_12524, n18740);
  and g30906 (n18741, n_12523, n_12524);
  not g30907 (n_12525, n18741);
  and g30908 (n18742, \asqrt[37] , n_12525);
  and g30912 (n18746, n_12075, n_12074);
  and g30913 (n18747, \asqrt[9] , n18746);
  not g30914 (n_12526, n18747);
  and g30915 (n18748, n_12073, n_12526);
  not g30916 (n_12527, n18745);
  not g30917 (n_12528, n18748);
  and g30918 (n18749, n_12527, n_12528);
  and g30919 (n18750, n_3474, n_12523);
  and g30920 (n18751, n_12524, n18750);
  not g30921 (n_12529, n18749);
  not g30922 (n_12530, n18751);
  and g30923 (n18752, n_12529, n_12530);
  not g30924 (n_12531, n18742);
  not g30925 (n_12532, n18752);
  and g30926 (n18753, n_12531, n_12532);
  not g30927 (n_12533, n18753);
  and g30928 (n18754, \asqrt[38] , n_12533);
  and g30932 (n18758, n_12083, n_12082);
  and g30933 (n18759, \asqrt[9] , n18758);
  not g30934 (n_12534, n18759);
  and g30935 (n18760, n_12081, n_12534);
  not g30936 (n_12535, n18757);
  not g30937 (n_12536, n18760);
  and g30938 (n18761, n_12535, n_12536);
  and g30939 (n18762, n_3242, n_12531);
  and g30940 (n18763, n_12532, n18762);
  not g30941 (n_12537, n18761);
  not g30942 (n_12538, n18763);
  and g30943 (n18764, n_12537, n_12538);
  not g30944 (n_12539, n18754);
  not g30945 (n_12540, n18764);
  and g30946 (n18765, n_12539, n_12540);
  not g30947 (n_12541, n18765);
  and g30948 (n18766, \asqrt[39] , n_12541);
  and g30952 (n18770, n_12091, n_12090);
  and g30953 (n18771, \asqrt[9] , n18770);
  not g30954 (n_12542, n18771);
  and g30955 (n18772, n_12089, n_12542);
  not g30956 (n_12543, n18769);
  not g30957 (n_12544, n18772);
  and g30958 (n18773, n_12543, n_12544);
  and g30959 (n18774, n_3018, n_12539);
  and g30960 (n18775, n_12540, n18774);
  not g30961 (n_12545, n18773);
  not g30962 (n_12546, n18775);
  and g30963 (n18776, n_12545, n_12546);
  not g30964 (n_12547, n18766);
  not g30965 (n_12548, n18776);
  and g30966 (n18777, n_12547, n_12548);
  not g30967 (n_12549, n18777);
  and g30968 (n18778, \asqrt[40] , n_12549);
  and g30972 (n18782, n_12099, n_12098);
  and g30973 (n18783, \asqrt[9] , n18782);
  not g30974 (n_12550, n18783);
  and g30975 (n18784, n_12097, n_12550);
  not g30976 (n_12551, n18781);
  not g30977 (n_12552, n18784);
  and g30978 (n18785, n_12551, n_12552);
  and g30979 (n18786, n_2802, n_12547);
  and g30980 (n18787, n_12548, n18786);
  not g30981 (n_12553, n18785);
  not g30982 (n_12554, n18787);
  and g30983 (n18788, n_12553, n_12554);
  not g30984 (n_12555, n18778);
  not g30985 (n_12556, n18788);
  and g30986 (n18789, n_12555, n_12556);
  not g30987 (n_12557, n18789);
  and g30988 (n18790, \asqrt[41] , n_12557);
  and g30992 (n18794, n_12107, n_12106);
  and g30993 (n18795, \asqrt[9] , n18794);
  not g30994 (n_12558, n18795);
  and g30995 (n18796, n_12105, n_12558);
  not g30996 (n_12559, n18793);
  not g30997 (n_12560, n18796);
  and g30998 (n18797, n_12559, n_12560);
  and g30999 (n18798, n_2594, n_12555);
  and g31000 (n18799, n_12556, n18798);
  not g31001 (n_12561, n18797);
  not g31002 (n_12562, n18799);
  and g31003 (n18800, n_12561, n_12562);
  not g31004 (n_12563, n18790);
  not g31005 (n_12564, n18800);
  and g31006 (n18801, n_12563, n_12564);
  not g31007 (n_12565, n18801);
  and g31008 (n18802, \asqrt[42] , n_12565);
  and g31012 (n18806, n_12115, n_12114);
  and g31013 (n18807, \asqrt[9] , n18806);
  not g31014 (n_12566, n18807);
  and g31015 (n18808, n_12113, n_12566);
  not g31016 (n_12567, n18805);
  not g31017 (n_12568, n18808);
  and g31018 (n18809, n_12567, n_12568);
  and g31019 (n18810, n_2394, n_12563);
  and g31020 (n18811, n_12564, n18810);
  not g31021 (n_12569, n18809);
  not g31022 (n_12570, n18811);
  and g31023 (n18812, n_12569, n_12570);
  not g31024 (n_12571, n18802);
  not g31025 (n_12572, n18812);
  and g31026 (n18813, n_12571, n_12572);
  not g31027 (n_12573, n18813);
  and g31028 (n18814, \asqrt[43] , n_12573);
  and g31032 (n18818, n_12123, n_12122);
  and g31033 (n18819, \asqrt[9] , n18818);
  not g31034 (n_12574, n18819);
  and g31035 (n18820, n_12121, n_12574);
  not g31036 (n_12575, n18817);
  not g31037 (n_12576, n18820);
  and g31038 (n18821, n_12575, n_12576);
  and g31039 (n18822, n_2202, n_12571);
  and g31040 (n18823, n_12572, n18822);
  not g31041 (n_12577, n18821);
  not g31042 (n_12578, n18823);
  and g31043 (n18824, n_12577, n_12578);
  not g31044 (n_12579, n18814);
  not g31045 (n_12580, n18824);
  and g31046 (n18825, n_12579, n_12580);
  not g31047 (n_12581, n18825);
  and g31048 (n18826, \asqrt[44] , n_12581);
  and g31052 (n18830, n_12131, n_12130);
  and g31053 (n18831, \asqrt[9] , n18830);
  not g31054 (n_12582, n18831);
  and g31055 (n18832, n_12129, n_12582);
  not g31056 (n_12583, n18829);
  not g31057 (n_12584, n18832);
  and g31058 (n18833, n_12583, n_12584);
  and g31059 (n18834, n_2018, n_12579);
  and g31060 (n18835, n_12580, n18834);
  not g31061 (n_12585, n18833);
  not g31062 (n_12586, n18835);
  and g31063 (n18836, n_12585, n_12586);
  not g31064 (n_12587, n18826);
  not g31065 (n_12588, n18836);
  and g31066 (n18837, n_12587, n_12588);
  not g31067 (n_12589, n18837);
  and g31068 (n18838, \asqrt[45] , n_12589);
  and g31072 (n18842, n_12139, n_12138);
  and g31073 (n18843, \asqrt[9] , n18842);
  not g31074 (n_12590, n18843);
  and g31075 (n18844, n_12137, n_12590);
  not g31076 (n_12591, n18841);
  not g31077 (n_12592, n18844);
  and g31078 (n18845, n_12591, n_12592);
  and g31079 (n18846, n_1842, n_12587);
  and g31080 (n18847, n_12588, n18846);
  not g31081 (n_12593, n18845);
  not g31082 (n_12594, n18847);
  and g31083 (n18848, n_12593, n_12594);
  not g31084 (n_12595, n18838);
  not g31085 (n_12596, n18848);
  and g31086 (n18849, n_12595, n_12596);
  not g31087 (n_12597, n18849);
  and g31088 (n18850, \asqrt[46] , n_12597);
  and g31092 (n18854, n_12147, n_12146);
  and g31093 (n18855, \asqrt[9] , n18854);
  not g31094 (n_12598, n18855);
  and g31095 (n18856, n_12145, n_12598);
  not g31096 (n_12599, n18853);
  not g31097 (n_12600, n18856);
  and g31098 (n18857, n_12599, n_12600);
  and g31099 (n18858, n_1674, n_12595);
  and g31100 (n18859, n_12596, n18858);
  not g31101 (n_12601, n18857);
  not g31102 (n_12602, n18859);
  and g31103 (n18860, n_12601, n_12602);
  not g31104 (n_12603, n18850);
  not g31105 (n_12604, n18860);
  and g31106 (n18861, n_12603, n_12604);
  not g31107 (n_12605, n18861);
  and g31108 (n18862, \asqrt[47] , n_12605);
  and g31112 (n18866, n_12155, n_12154);
  and g31113 (n18867, \asqrt[9] , n18866);
  not g31114 (n_12606, n18867);
  and g31115 (n18868, n_12153, n_12606);
  not g31116 (n_12607, n18865);
  not g31117 (n_12608, n18868);
  and g31118 (n18869, n_12607, n_12608);
  and g31119 (n18870, n_1514, n_12603);
  and g31120 (n18871, n_12604, n18870);
  not g31121 (n_12609, n18869);
  not g31122 (n_12610, n18871);
  and g31123 (n18872, n_12609, n_12610);
  not g31124 (n_12611, n18862);
  not g31125 (n_12612, n18872);
  and g31126 (n18873, n_12611, n_12612);
  not g31127 (n_12613, n18873);
  and g31128 (n18874, \asqrt[48] , n_12613);
  and g31132 (n18878, n_12163, n_12162);
  and g31133 (n18879, \asqrt[9] , n18878);
  not g31134 (n_12614, n18879);
  and g31135 (n18880, n_12161, n_12614);
  not g31136 (n_12615, n18877);
  not g31137 (n_12616, n18880);
  and g31138 (n18881, n_12615, n_12616);
  and g31139 (n18882, n_1362, n_12611);
  and g31140 (n18883, n_12612, n18882);
  not g31141 (n_12617, n18881);
  not g31142 (n_12618, n18883);
  and g31143 (n18884, n_12617, n_12618);
  not g31144 (n_12619, n18874);
  not g31145 (n_12620, n18884);
  and g31146 (n18885, n_12619, n_12620);
  not g31147 (n_12621, n18885);
  and g31148 (n18886, \asqrt[49] , n_12621);
  and g31152 (n18890, n_12171, n_12170);
  and g31153 (n18891, \asqrt[9] , n18890);
  not g31154 (n_12622, n18891);
  and g31155 (n18892, n_12169, n_12622);
  not g31156 (n_12623, n18889);
  not g31157 (n_12624, n18892);
  and g31158 (n18893, n_12623, n_12624);
  and g31159 (n18894, n_1218, n_12619);
  and g31160 (n18895, n_12620, n18894);
  not g31161 (n_12625, n18893);
  not g31162 (n_12626, n18895);
  and g31163 (n18896, n_12625, n_12626);
  not g31164 (n_12627, n18886);
  not g31165 (n_12628, n18896);
  and g31166 (n18897, n_12627, n_12628);
  not g31167 (n_12629, n18897);
  and g31168 (n18898, \asqrt[50] , n_12629);
  and g31172 (n18902, n_12179, n_12178);
  and g31173 (n18903, \asqrt[9] , n18902);
  not g31174 (n_12630, n18903);
  and g31175 (n18904, n_12177, n_12630);
  not g31176 (n_12631, n18901);
  not g31177 (n_12632, n18904);
  and g31178 (n18905, n_12631, n_12632);
  and g31179 (n18906, n_1082, n_12627);
  and g31180 (n18907, n_12628, n18906);
  not g31181 (n_12633, n18905);
  not g31182 (n_12634, n18907);
  and g31183 (n18908, n_12633, n_12634);
  not g31184 (n_12635, n18898);
  not g31185 (n_12636, n18908);
  and g31186 (n18909, n_12635, n_12636);
  not g31187 (n_12637, n18909);
  and g31188 (n18910, \asqrt[51] , n_12637);
  and g31192 (n18914, n_12187, n_12186);
  and g31193 (n18915, \asqrt[9] , n18914);
  not g31194 (n_12638, n18915);
  and g31195 (n18916, n_12185, n_12638);
  not g31196 (n_12639, n18913);
  not g31197 (n_12640, n18916);
  and g31198 (n18917, n_12639, n_12640);
  and g31199 (n18918, n_954, n_12635);
  and g31200 (n18919, n_12636, n18918);
  not g31201 (n_12641, n18917);
  not g31202 (n_12642, n18919);
  and g31203 (n18920, n_12641, n_12642);
  not g31204 (n_12643, n18910);
  not g31205 (n_12644, n18920);
  and g31206 (n18921, n_12643, n_12644);
  not g31207 (n_12645, n18921);
  and g31208 (n18922, \asqrt[52] , n_12645);
  and g31212 (n18926, n_12195, n_12194);
  and g31213 (n18927, \asqrt[9] , n18926);
  not g31214 (n_12646, n18927);
  and g31215 (n18928, n_12193, n_12646);
  not g31216 (n_12647, n18925);
  not g31217 (n_12648, n18928);
  and g31218 (n18929, n_12647, n_12648);
  and g31219 (n18930, n_834, n_12643);
  and g31220 (n18931, n_12644, n18930);
  not g31221 (n_12649, n18929);
  not g31222 (n_12650, n18931);
  and g31223 (n18932, n_12649, n_12650);
  not g31224 (n_12651, n18922);
  not g31225 (n_12652, n18932);
  and g31226 (n18933, n_12651, n_12652);
  not g31227 (n_12653, n18933);
  and g31228 (n18934, \asqrt[53] , n_12653);
  and g31232 (n18938, n_12203, n_12202);
  and g31233 (n18939, \asqrt[9] , n18938);
  not g31234 (n_12654, n18939);
  and g31235 (n18940, n_12201, n_12654);
  not g31236 (n_12655, n18937);
  not g31237 (n_12656, n18940);
  and g31238 (n18941, n_12655, n_12656);
  and g31239 (n18942, n_722, n_12651);
  and g31240 (n18943, n_12652, n18942);
  not g31241 (n_12657, n18941);
  not g31242 (n_12658, n18943);
  and g31243 (n18944, n_12657, n_12658);
  not g31244 (n_12659, n18934);
  not g31245 (n_12660, n18944);
  and g31246 (n18945, n_12659, n_12660);
  not g31247 (n_12661, n18945);
  and g31248 (n18946, \asqrt[54] , n_12661);
  and g31252 (n18950, n_12211, n_12210);
  and g31253 (n18951, \asqrt[9] , n18950);
  not g31254 (n_12662, n18951);
  and g31255 (n18952, n_12209, n_12662);
  not g31256 (n_12663, n18949);
  not g31257 (n_12664, n18952);
  and g31258 (n18953, n_12663, n_12664);
  and g31259 (n18954, n_618, n_12659);
  and g31260 (n18955, n_12660, n18954);
  not g31261 (n_12665, n18953);
  not g31262 (n_12666, n18955);
  and g31263 (n18956, n_12665, n_12666);
  not g31264 (n_12667, n18946);
  not g31265 (n_12668, n18956);
  and g31266 (n18957, n_12667, n_12668);
  not g31267 (n_12669, n18957);
  and g31268 (n18958, \asqrt[55] , n_12669);
  and g31272 (n18962, n_12219, n_12218);
  and g31273 (n18963, \asqrt[9] , n18962);
  not g31274 (n_12670, n18963);
  and g31275 (n18964, n_12217, n_12670);
  not g31276 (n_12671, n18961);
  not g31277 (n_12672, n18964);
  and g31278 (n18965, n_12671, n_12672);
  and g31279 (n18966, n_522, n_12667);
  and g31280 (n18967, n_12668, n18966);
  not g31281 (n_12673, n18965);
  not g31282 (n_12674, n18967);
  and g31283 (n18968, n_12673, n_12674);
  not g31284 (n_12675, n18958);
  not g31285 (n_12676, n18968);
  and g31286 (n18969, n_12675, n_12676);
  not g31287 (n_12677, n18969);
  and g31288 (n18970, \asqrt[56] , n_12677);
  and g31289 (n18971, n_434, n_12675);
  and g31290 (n18972, n_12676, n18971);
  and g31294 (n18976, n_12227, n_12225);
  and g31295 (n18977, \asqrt[9] , n18976);
  not g31296 (n_12678, n18977);
  and g31297 (n18978, n_12226, n_12678);
  not g31298 (n_12679, n18975);
  not g31299 (n_12680, n18978);
  and g31300 (n18979, n_12679, n_12680);
  not g31301 (n_12681, n18972);
  not g31302 (n_12682, n18979);
  and g31303 (n18980, n_12681, n_12682);
  not g31304 (n_12683, n18970);
  not g31305 (n_12684, n18980);
  and g31306 (n18981, n_12683, n_12684);
  not g31307 (n_12685, n18981);
  and g31308 (n18982, \asqrt[57] , n_12685);
  and g31312 (n18986, n_12235, n_12234);
  and g31313 (n18987, \asqrt[9] , n18986);
  not g31314 (n_12686, n18987);
  and g31315 (n18988, n_12233, n_12686);
  not g31316 (n_12687, n18985);
  not g31317 (n_12688, n18988);
  and g31318 (n18989, n_12687, n_12688);
  and g31319 (n18990, n_354, n_12683);
  and g31320 (n18991, n_12684, n18990);
  not g31321 (n_12689, n18989);
  not g31322 (n_12690, n18991);
  and g31323 (n18992, n_12689, n_12690);
  not g31324 (n_12691, n18982);
  not g31325 (n_12692, n18992);
  and g31326 (n18993, n_12691, n_12692);
  not g31327 (n_12693, n18993);
  and g31328 (n18994, \asqrt[58] , n_12693);
  and g31332 (n18998, n_12243, n_12242);
  and g31333 (n18999, \asqrt[9] , n18998);
  not g31334 (n_12694, n18999);
  and g31335 (n19000, n_12241, n_12694);
  not g31336 (n_12695, n18997);
  not g31337 (n_12696, n19000);
  and g31338 (n19001, n_12695, n_12696);
  and g31339 (n19002, n_282, n_12691);
  and g31340 (n19003, n_12692, n19002);
  not g31341 (n_12697, n19001);
  not g31342 (n_12698, n19003);
  and g31343 (n19004, n_12697, n_12698);
  not g31344 (n_12699, n18994);
  not g31345 (n_12700, n19004);
  and g31346 (n19005, n_12699, n_12700);
  not g31347 (n_12701, n19005);
  and g31348 (n19006, \asqrt[59] , n_12701);
  and g31352 (n19010, n_12251, n_12250);
  and g31353 (n19011, \asqrt[9] , n19010);
  not g31354 (n_12702, n19011);
  and g31355 (n19012, n_12249, n_12702);
  not g31356 (n_12703, n19009);
  not g31357 (n_12704, n19012);
  and g31358 (n19013, n_12703, n_12704);
  and g31359 (n19014, n_218, n_12699);
  and g31360 (n19015, n_12700, n19014);
  not g31361 (n_12705, n19013);
  not g31362 (n_12706, n19015);
  and g31363 (n19016, n_12705, n_12706);
  not g31364 (n_12707, n19006);
  not g31365 (n_12708, n19016);
  and g31366 (n19017, n_12707, n_12708);
  not g31367 (n_12709, n19017);
  and g31368 (n19018, \asqrt[60] , n_12709);
  and g31372 (n19022, n_12259, n_12258);
  and g31373 (n19023, \asqrt[9] , n19022);
  not g31374 (n_12710, n19023);
  and g31375 (n19024, n_12257, n_12710);
  not g31376 (n_12711, n19021);
  not g31377 (n_12712, n19024);
  and g31378 (n19025, n_12711, n_12712);
  and g31379 (n19026, n_162, n_12707);
  and g31380 (n19027, n_12708, n19026);
  not g31381 (n_12713, n19025);
  not g31382 (n_12714, n19027);
  and g31383 (n19028, n_12713, n_12714);
  not g31384 (n_12715, n19018);
  not g31385 (n_12716, n19028);
  and g31386 (n19029, n_12715, n_12716);
  not g31387 (n_12717, n19029);
  and g31388 (n19030, \asqrt[61] , n_12717);
  and g31392 (n19034, n_12267, n_12266);
  and g31393 (n19035, \asqrt[9] , n19034);
  not g31394 (n_12718, n19035);
  and g31395 (n19036, n_12265, n_12718);
  not g31396 (n_12719, n19033);
  not g31397 (n_12720, n19036);
  and g31398 (n19037, n_12719, n_12720);
  and g31399 (n19038, n_115, n_12715);
  and g31400 (n19039, n_12716, n19038);
  not g31401 (n_12721, n19037);
  not g31402 (n_12722, n19039);
  and g31403 (n19040, n_12721, n_12722);
  not g31404 (n_12723, n19030);
  not g31405 (n_12724, n19040);
  and g31406 (n19041, n_12723, n_12724);
  not g31407 (n_12725, n19041);
  and g31408 (n19042, \asqrt[62] , n_12725);
  and g31412 (n19046, n_12275, n_12274);
  and g31413 (n19047, \asqrt[9] , n19046);
  not g31414 (n_12726, n19047);
  and g31415 (n19048, n_12273, n_12726);
  not g31416 (n_12727, n19045);
  not g31417 (n_12728, n19048);
  and g31418 (n19049, n_12727, n_12728);
  and g31419 (n19050, n_76, n_12723);
  and g31420 (n19051, n_12724, n19050);
  not g31421 (n_12729, n19049);
  not g31422 (n_12730, n19051);
  and g31423 (n19052, n_12729, n_12730);
  not g31424 (n_12731, n19042);
  not g31425 (n_12732, n19052);
  and g31426 (n19053, n_12731, n_12732);
  and g31430 (n19057, n_12283, n_12282);
  and g31431 (n19058, \asqrt[9] , n19057);
  not g31432 (n_12733, n19058);
  and g31433 (n19059, n_12281, n_12733);
  not g31434 (n_12734, n19056);
  not g31435 (n_12735, n19059);
  and g31436 (n19060, n_12734, n_12735);
  and g31437 (n19061, n_12290, n_12289);
  and g31438 (n19062, \asqrt[9] , n19061);
  not g31441 (n_12737, n19060);
  not g31443 (n_12738, n19053);
  not g31445 (n_12739, n19065);
  and g31446 (n19066, n_21, n_12739);
  and g31447 (n19067, n_12731, n19060);
  and g31448 (n19068, n_12732, n19067);
  and g31449 (n19069, n_12289, \asqrt[9] );
  not g31450 (n_12740, n19069);
  and g31451 (n19070, n18385, n_12740);
  not g31452 (n_12741, n19061);
  and g31453 (n19071, \asqrt[63] , n_12741);
  not g31454 (n_12742, n19070);
  and g31455 (n19072, n_12742, n19071);
  not g31461 (n_12743, n19072);
  not g31462 (n_12744, n19077);
  not g31464 (n_12745, n19068);
  and g31468 (n19081, \a[16] , \asqrt[8] );
  not g31469 (n_12750, \a[14] );
  not g31470 (n_12751, \a[15] );
  and g31471 (n19082, n_12750, n_12751);
  and g31472 (n19083, n_12302, n19082);
  not g31473 (n_12752, n19081);
  not g31474 (n_12753, n19083);
  and g31475 (n19084, n_12752, n_12753);
  not g31476 (n_12754, n19084);
  and g31477 (n19085, \asqrt[9] , n_12754);
  and g31483 (n19091, n_12302, \asqrt[8] );
  not g31484 (n_12755, n19091);
  and g31485 (n19092, \a[17] , n_12755);
  and g31486 (n19093, n18414, \asqrt[8] );
  not g31487 (n_12756, n19092);
  not g31488 (n_12757, n19093);
  and g31489 (n19094, n_12756, n_12757);
  not g31490 (n_12758, n19090);
  and g31491 (n19095, n_12758, n19094);
  not g31492 (n_12759, n19085);
  not g31493 (n_12760, n19095);
  and g31494 (n19096, n_12759, n_12760);
  not g31495 (n_12761, n19096);
  and g31496 (n19097, \asqrt[10] , n_12761);
  not g31497 (n_12762, \asqrt[10] );
  and g31498 (n19098, n_12762, n_12759);
  and g31499 (n19099, n_12760, n19098);
  not g31503 (n_12763, n19066);
  not g31505 (n_12764, n19103);
  and g31506 (n19104, n_12757, n_12764);
  not g31507 (n_12765, n19104);
  and g31508 (n19105, \a[18] , n_12765);
  and g31509 (n19106, n_11862, n_12764);
  and g31510 (n19107, n_12757, n19106);
  not g31511 (n_12766, n19105);
  not g31512 (n_12767, n19107);
  and g31513 (n19108, n_12766, n_12767);
  not g31514 (n_12768, n19099);
  not g31515 (n_12769, n19108);
  and g31516 (n19109, n_12768, n_12769);
  not g31517 (n_12770, n19097);
  not g31518 (n_12771, n19109);
  and g31519 (n19110, n_12770, n_12771);
  not g31520 (n_12772, n19110);
  and g31521 (n19111, \asqrt[11] , n_12772);
  and g31522 (n19112, n_12311, n_12310);
  not g31523 (n_12773, n18426);
  and g31524 (n19113, n_12773, n19112);
  and g31525 (n19114, \asqrt[8] , n19113);
  and g31526 (n19115, \asqrt[8] , n19112);
  not g31527 (n_12774, n19115);
  and g31528 (n19116, n18426, n_12774);
  not g31529 (n_12775, n19114);
  not g31530 (n_12776, n19116);
  and g31531 (n19117, n_12775, n_12776);
  and g31532 (n19118, n_12314, n_12770);
  and g31533 (n19119, n_12771, n19118);
  not g31534 (n_12777, n19117);
  not g31535 (n_12778, n19119);
  and g31536 (n19120, n_12777, n_12778);
  not g31537 (n_12779, n19111);
  not g31538 (n_12780, n19120);
  and g31539 (n19121, n_12779, n_12780);
  not g31540 (n_12781, n19121);
  and g31541 (n19122, \asqrt[12] , n_12781);
  and g31545 (n19126, n_12322, n_12320);
  and g31546 (n19127, \asqrt[8] , n19126);
  not g31547 (n_12782, n19127);
  and g31548 (n19128, n_12321, n_12782);
  not g31549 (n_12783, n19125);
  not g31550 (n_12784, n19128);
  and g31551 (n19129, n_12783, n_12784);
  and g31552 (n19130, n_11874, n_12779);
  and g31553 (n19131, n_12780, n19130);
  not g31554 (n_12785, n19129);
  not g31555 (n_12786, n19131);
  and g31556 (n19132, n_12785, n_12786);
  not g31557 (n_12787, n19122);
  not g31558 (n_12788, n19132);
  and g31559 (n19133, n_12787, n_12788);
  not g31560 (n_12789, n19133);
  and g31561 (n19134, \asqrt[13] , n_12789);
  and g31565 (n19138, n_12331, n_12330);
  and g31566 (n19139, \asqrt[8] , n19138);
  not g31567 (n_12790, n19139);
  and g31568 (n19140, n_12329, n_12790);
  not g31569 (n_12791, n19137);
  not g31570 (n_12792, n19140);
  and g31571 (n19141, n_12791, n_12792);
  and g31572 (n19142, n_11442, n_12787);
  and g31573 (n19143, n_12788, n19142);
  not g31574 (n_12793, n19141);
  not g31575 (n_12794, n19143);
  and g31576 (n19144, n_12793, n_12794);
  not g31577 (n_12795, n19134);
  not g31578 (n_12796, n19144);
  and g31579 (n19145, n_12795, n_12796);
  not g31580 (n_12797, n19145);
  and g31581 (n19146, \asqrt[14] , n_12797);
  and g31585 (n19150, n_12339, n_12338);
  and g31586 (n19151, \asqrt[8] , n19150);
  not g31587 (n_12798, n19151);
  and g31588 (n19152, n_12337, n_12798);
  not g31589 (n_12799, n19149);
  not g31590 (n_12800, n19152);
  and g31591 (n19153, n_12799, n_12800);
  and g31592 (n19154, n_11018, n_12795);
  and g31593 (n19155, n_12796, n19154);
  not g31594 (n_12801, n19153);
  not g31595 (n_12802, n19155);
  and g31596 (n19156, n_12801, n_12802);
  not g31597 (n_12803, n19146);
  not g31598 (n_12804, n19156);
  and g31599 (n19157, n_12803, n_12804);
  not g31600 (n_12805, n19157);
  and g31601 (n19158, \asqrt[15] , n_12805);
  and g31605 (n19162, n_12347, n_12346);
  and g31606 (n19163, \asqrt[8] , n19162);
  not g31607 (n_12806, n19163);
  and g31608 (n19164, n_12345, n_12806);
  not g31609 (n_12807, n19161);
  not g31610 (n_12808, n19164);
  and g31611 (n19165, n_12807, n_12808);
  and g31612 (n19166, n_10602, n_12803);
  and g31613 (n19167, n_12804, n19166);
  not g31614 (n_12809, n19165);
  not g31615 (n_12810, n19167);
  and g31616 (n19168, n_12809, n_12810);
  not g31617 (n_12811, n19158);
  not g31618 (n_12812, n19168);
  and g31619 (n19169, n_12811, n_12812);
  not g31620 (n_12813, n19169);
  and g31621 (n19170, \asqrt[16] , n_12813);
  and g31625 (n19174, n_12355, n_12354);
  and g31626 (n19175, \asqrt[8] , n19174);
  not g31627 (n_12814, n19175);
  and g31628 (n19176, n_12353, n_12814);
  not g31629 (n_12815, n19173);
  not g31630 (n_12816, n19176);
  and g31631 (n19177, n_12815, n_12816);
  and g31632 (n19178, n_10194, n_12811);
  and g31633 (n19179, n_12812, n19178);
  not g31634 (n_12817, n19177);
  not g31635 (n_12818, n19179);
  and g31636 (n19180, n_12817, n_12818);
  not g31637 (n_12819, n19170);
  not g31638 (n_12820, n19180);
  and g31639 (n19181, n_12819, n_12820);
  not g31640 (n_12821, n19181);
  and g31641 (n19182, \asqrt[17] , n_12821);
  and g31645 (n19186, n_12363, n_12362);
  and g31646 (n19187, \asqrt[8] , n19186);
  not g31647 (n_12822, n19187);
  and g31648 (n19188, n_12361, n_12822);
  not g31649 (n_12823, n19185);
  not g31650 (n_12824, n19188);
  and g31651 (n19189, n_12823, n_12824);
  and g31652 (n19190, n_9794, n_12819);
  and g31653 (n19191, n_12820, n19190);
  not g31654 (n_12825, n19189);
  not g31655 (n_12826, n19191);
  and g31656 (n19192, n_12825, n_12826);
  not g31657 (n_12827, n19182);
  not g31658 (n_12828, n19192);
  and g31659 (n19193, n_12827, n_12828);
  not g31660 (n_12829, n19193);
  and g31661 (n19194, \asqrt[18] , n_12829);
  and g31665 (n19198, n_12371, n_12370);
  and g31666 (n19199, \asqrt[8] , n19198);
  not g31667 (n_12830, n19199);
  and g31668 (n19200, n_12369, n_12830);
  not g31669 (n_12831, n19197);
  not g31670 (n_12832, n19200);
  and g31671 (n19201, n_12831, n_12832);
  and g31672 (n19202, n_9402, n_12827);
  and g31673 (n19203, n_12828, n19202);
  not g31674 (n_12833, n19201);
  not g31675 (n_12834, n19203);
  and g31676 (n19204, n_12833, n_12834);
  not g31677 (n_12835, n19194);
  not g31678 (n_12836, n19204);
  and g31679 (n19205, n_12835, n_12836);
  not g31680 (n_12837, n19205);
  and g31681 (n19206, \asqrt[19] , n_12837);
  and g31685 (n19210, n_12379, n_12378);
  and g31686 (n19211, \asqrt[8] , n19210);
  not g31687 (n_12838, n19211);
  and g31688 (n19212, n_12377, n_12838);
  not g31689 (n_12839, n19209);
  not g31690 (n_12840, n19212);
  and g31691 (n19213, n_12839, n_12840);
  and g31692 (n19214, n_9018, n_12835);
  and g31693 (n19215, n_12836, n19214);
  not g31694 (n_12841, n19213);
  not g31695 (n_12842, n19215);
  and g31696 (n19216, n_12841, n_12842);
  not g31697 (n_12843, n19206);
  not g31698 (n_12844, n19216);
  and g31699 (n19217, n_12843, n_12844);
  not g31700 (n_12845, n19217);
  and g31701 (n19218, \asqrt[20] , n_12845);
  and g31705 (n19222, n_12387, n_12386);
  and g31706 (n19223, \asqrt[8] , n19222);
  not g31707 (n_12846, n19223);
  and g31708 (n19224, n_12385, n_12846);
  not g31709 (n_12847, n19221);
  not g31710 (n_12848, n19224);
  and g31711 (n19225, n_12847, n_12848);
  and g31712 (n19226, n_8642, n_12843);
  and g31713 (n19227, n_12844, n19226);
  not g31714 (n_12849, n19225);
  not g31715 (n_12850, n19227);
  and g31716 (n19228, n_12849, n_12850);
  not g31717 (n_12851, n19218);
  not g31718 (n_12852, n19228);
  and g31719 (n19229, n_12851, n_12852);
  not g31720 (n_12853, n19229);
  and g31721 (n19230, \asqrt[21] , n_12853);
  and g31725 (n19234, n_12395, n_12394);
  and g31726 (n19235, \asqrt[8] , n19234);
  not g31727 (n_12854, n19235);
  and g31728 (n19236, n_12393, n_12854);
  not g31729 (n_12855, n19233);
  not g31730 (n_12856, n19236);
  and g31731 (n19237, n_12855, n_12856);
  and g31732 (n19238, n_8274, n_12851);
  and g31733 (n19239, n_12852, n19238);
  not g31734 (n_12857, n19237);
  not g31735 (n_12858, n19239);
  and g31736 (n19240, n_12857, n_12858);
  not g31737 (n_12859, n19230);
  not g31738 (n_12860, n19240);
  and g31739 (n19241, n_12859, n_12860);
  not g31740 (n_12861, n19241);
  and g31741 (n19242, \asqrt[22] , n_12861);
  and g31745 (n19246, n_12403, n_12402);
  and g31746 (n19247, \asqrt[8] , n19246);
  not g31747 (n_12862, n19247);
  and g31748 (n19248, n_12401, n_12862);
  not g31749 (n_12863, n19245);
  not g31750 (n_12864, n19248);
  and g31751 (n19249, n_12863, n_12864);
  and g31752 (n19250, n_7914, n_12859);
  and g31753 (n19251, n_12860, n19250);
  not g31754 (n_12865, n19249);
  not g31755 (n_12866, n19251);
  and g31756 (n19252, n_12865, n_12866);
  not g31757 (n_12867, n19242);
  not g31758 (n_12868, n19252);
  and g31759 (n19253, n_12867, n_12868);
  not g31760 (n_12869, n19253);
  and g31761 (n19254, \asqrt[23] , n_12869);
  and g31765 (n19258, n_12411, n_12410);
  and g31766 (n19259, \asqrt[8] , n19258);
  not g31767 (n_12870, n19259);
  and g31768 (n19260, n_12409, n_12870);
  not g31769 (n_12871, n19257);
  not g31770 (n_12872, n19260);
  and g31771 (n19261, n_12871, n_12872);
  and g31772 (n19262, n_7562, n_12867);
  and g31773 (n19263, n_12868, n19262);
  not g31774 (n_12873, n19261);
  not g31775 (n_12874, n19263);
  and g31776 (n19264, n_12873, n_12874);
  not g31777 (n_12875, n19254);
  not g31778 (n_12876, n19264);
  and g31779 (n19265, n_12875, n_12876);
  not g31780 (n_12877, n19265);
  and g31781 (n19266, \asqrt[24] , n_12877);
  and g31785 (n19270, n_12419, n_12418);
  and g31786 (n19271, \asqrt[8] , n19270);
  not g31787 (n_12878, n19271);
  and g31788 (n19272, n_12417, n_12878);
  not g31789 (n_12879, n19269);
  not g31790 (n_12880, n19272);
  and g31791 (n19273, n_12879, n_12880);
  and g31792 (n19274, n_7218, n_12875);
  and g31793 (n19275, n_12876, n19274);
  not g31794 (n_12881, n19273);
  not g31795 (n_12882, n19275);
  and g31796 (n19276, n_12881, n_12882);
  not g31797 (n_12883, n19266);
  not g31798 (n_12884, n19276);
  and g31799 (n19277, n_12883, n_12884);
  not g31800 (n_12885, n19277);
  and g31801 (n19278, \asqrt[25] , n_12885);
  and g31805 (n19282, n_12427, n_12426);
  and g31806 (n19283, \asqrt[8] , n19282);
  not g31807 (n_12886, n19283);
  and g31808 (n19284, n_12425, n_12886);
  not g31809 (n_12887, n19281);
  not g31810 (n_12888, n19284);
  and g31811 (n19285, n_12887, n_12888);
  and g31812 (n19286, n_6882, n_12883);
  and g31813 (n19287, n_12884, n19286);
  not g31814 (n_12889, n19285);
  not g31815 (n_12890, n19287);
  and g31816 (n19288, n_12889, n_12890);
  not g31817 (n_12891, n19278);
  not g31818 (n_12892, n19288);
  and g31819 (n19289, n_12891, n_12892);
  not g31820 (n_12893, n19289);
  and g31821 (n19290, \asqrt[26] , n_12893);
  and g31825 (n19294, n_12435, n_12434);
  and g31826 (n19295, \asqrt[8] , n19294);
  not g31827 (n_12894, n19295);
  and g31828 (n19296, n_12433, n_12894);
  not g31829 (n_12895, n19293);
  not g31830 (n_12896, n19296);
  and g31831 (n19297, n_12895, n_12896);
  and g31832 (n19298, n_6554, n_12891);
  and g31833 (n19299, n_12892, n19298);
  not g31834 (n_12897, n19297);
  not g31835 (n_12898, n19299);
  and g31836 (n19300, n_12897, n_12898);
  not g31837 (n_12899, n19290);
  not g31838 (n_12900, n19300);
  and g31839 (n19301, n_12899, n_12900);
  not g31840 (n_12901, n19301);
  and g31841 (n19302, \asqrt[27] , n_12901);
  and g31845 (n19306, n_12443, n_12442);
  and g31846 (n19307, \asqrt[8] , n19306);
  not g31847 (n_12902, n19307);
  and g31848 (n19308, n_12441, n_12902);
  not g31849 (n_12903, n19305);
  not g31850 (n_12904, n19308);
  and g31851 (n19309, n_12903, n_12904);
  and g31852 (n19310, n_6234, n_12899);
  and g31853 (n19311, n_12900, n19310);
  not g31854 (n_12905, n19309);
  not g31855 (n_12906, n19311);
  and g31856 (n19312, n_12905, n_12906);
  not g31857 (n_12907, n19302);
  not g31858 (n_12908, n19312);
  and g31859 (n19313, n_12907, n_12908);
  not g31860 (n_12909, n19313);
  and g31861 (n19314, \asqrt[28] , n_12909);
  and g31865 (n19318, n_12451, n_12450);
  and g31866 (n19319, \asqrt[8] , n19318);
  not g31867 (n_12910, n19319);
  and g31868 (n19320, n_12449, n_12910);
  not g31869 (n_12911, n19317);
  not g31870 (n_12912, n19320);
  and g31871 (n19321, n_12911, n_12912);
  and g31872 (n19322, n_5922, n_12907);
  and g31873 (n19323, n_12908, n19322);
  not g31874 (n_12913, n19321);
  not g31875 (n_12914, n19323);
  and g31876 (n19324, n_12913, n_12914);
  not g31877 (n_12915, n19314);
  not g31878 (n_12916, n19324);
  and g31879 (n19325, n_12915, n_12916);
  not g31880 (n_12917, n19325);
  and g31881 (n19326, \asqrt[29] , n_12917);
  and g31885 (n19330, n_12459, n_12458);
  and g31886 (n19331, \asqrt[8] , n19330);
  not g31887 (n_12918, n19331);
  and g31888 (n19332, n_12457, n_12918);
  not g31889 (n_12919, n19329);
  not g31890 (n_12920, n19332);
  and g31891 (n19333, n_12919, n_12920);
  and g31892 (n19334, n_5618, n_12915);
  and g31893 (n19335, n_12916, n19334);
  not g31894 (n_12921, n19333);
  not g31895 (n_12922, n19335);
  and g31896 (n19336, n_12921, n_12922);
  not g31897 (n_12923, n19326);
  not g31898 (n_12924, n19336);
  and g31899 (n19337, n_12923, n_12924);
  not g31900 (n_12925, n19337);
  and g31901 (n19338, \asqrt[30] , n_12925);
  and g31905 (n19342, n_12467, n_12466);
  and g31906 (n19343, \asqrt[8] , n19342);
  not g31907 (n_12926, n19343);
  and g31908 (n19344, n_12465, n_12926);
  not g31909 (n_12927, n19341);
  not g31910 (n_12928, n19344);
  and g31911 (n19345, n_12927, n_12928);
  and g31912 (n19346, n_5322, n_12923);
  and g31913 (n19347, n_12924, n19346);
  not g31914 (n_12929, n19345);
  not g31915 (n_12930, n19347);
  and g31916 (n19348, n_12929, n_12930);
  not g31917 (n_12931, n19338);
  not g31918 (n_12932, n19348);
  and g31919 (n19349, n_12931, n_12932);
  not g31920 (n_12933, n19349);
  and g31921 (n19350, \asqrt[31] , n_12933);
  and g31925 (n19354, n_12475, n_12474);
  and g31926 (n19355, \asqrt[8] , n19354);
  not g31927 (n_12934, n19355);
  and g31928 (n19356, n_12473, n_12934);
  not g31929 (n_12935, n19353);
  not g31930 (n_12936, n19356);
  and g31931 (n19357, n_12935, n_12936);
  and g31932 (n19358, n_5034, n_12931);
  and g31933 (n19359, n_12932, n19358);
  not g31934 (n_12937, n19357);
  not g31935 (n_12938, n19359);
  and g31936 (n19360, n_12937, n_12938);
  not g31937 (n_12939, n19350);
  not g31938 (n_12940, n19360);
  and g31939 (n19361, n_12939, n_12940);
  not g31940 (n_12941, n19361);
  and g31941 (n19362, \asqrt[32] , n_12941);
  and g31945 (n19366, n_12483, n_12482);
  and g31946 (n19367, \asqrt[8] , n19366);
  not g31947 (n_12942, n19367);
  and g31948 (n19368, n_12481, n_12942);
  not g31949 (n_12943, n19365);
  not g31950 (n_12944, n19368);
  and g31951 (n19369, n_12943, n_12944);
  and g31952 (n19370, n_4754, n_12939);
  and g31953 (n19371, n_12940, n19370);
  not g31954 (n_12945, n19369);
  not g31955 (n_12946, n19371);
  and g31956 (n19372, n_12945, n_12946);
  not g31957 (n_12947, n19362);
  not g31958 (n_12948, n19372);
  and g31959 (n19373, n_12947, n_12948);
  not g31960 (n_12949, n19373);
  and g31961 (n19374, \asqrt[33] , n_12949);
  and g31965 (n19378, n_12491, n_12490);
  and g31966 (n19379, \asqrt[8] , n19378);
  not g31967 (n_12950, n19379);
  and g31968 (n19380, n_12489, n_12950);
  not g31969 (n_12951, n19377);
  not g31970 (n_12952, n19380);
  and g31971 (n19381, n_12951, n_12952);
  and g31972 (n19382, n_4482, n_12947);
  and g31973 (n19383, n_12948, n19382);
  not g31974 (n_12953, n19381);
  not g31975 (n_12954, n19383);
  and g31976 (n19384, n_12953, n_12954);
  not g31977 (n_12955, n19374);
  not g31978 (n_12956, n19384);
  and g31979 (n19385, n_12955, n_12956);
  not g31980 (n_12957, n19385);
  and g31981 (n19386, \asqrt[34] , n_12957);
  and g31985 (n19390, n_12499, n_12498);
  and g31986 (n19391, \asqrt[8] , n19390);
  not g31987 (n_12958, n19391);
  and g31988 (n19392, n_12497, n_12958);
  not g31989 (n_12959, n19389);
  not g31990 (n_12960, n19392);
  and g31991 (n19393, n_12959, n_12960);
  and g31992 (n19394, n_4218, n_12955);
  and g31993 (n19395, n_12956, n19394);
  not g31994 (n_12961, n19393);
  not g31995 (n_12962, n19395);
  and g31996 (n19396, n_12961, n_12962);
  not g31997 (n_12963, n19386);
  not g31998 (n_12964, n19396);
  and g31999 (n19397, n_12963, n_12964);
  not g32000 (n_12965, n19397);
  and g32001 (n19398, \asqrt[35] , n_12965);
  and g32005 (n19402, n_12507, n_12506);
  and g32006 (n19403, \asqrt[8] , n19402);
  not g32007 (n_12966, n19403);
  and g32008 (n19404, n_12505, n_12966);
  not g32009 (n_12967, n19401);
  not g32010 (n_12968, n19404);
  and g32011 (n19405, n_12967, n_12968);
  and g32012 (n19406, n_3962, n_12963);
  and g32013 (n19407, n_12964, n19406);
  not g32014 (n_12969, n19405);
  not g32015 (n_12970, n19407);
  and g32016 (n19408, n_12969, n_12970);
  not g32017 (n_12971, n19398);
  not g32018 (n_12972, n19408);
  and g32019 (n19409, n_12971, n_12972);
  not g32020 (n_12973, n19409);
  and g32021 (n19410, \asqrt[36] , n_12973);
  and g32025 (n19414, n_12515, n_12514);
  and g32026 (n19415, \asqrt[8] , n19414);
  not g32027 (n_12974, n19415);
  and g32028 (n19416, n_12513, n_12974);
  not g32029 (n_12975, n19413);
  not g32030 (n_12976, n19416);
  and g32031 (n19417, n_12975, n_12976);
  and g32032 (n19418, n_3714, n_12971);
  and g32033 (n19419, n_12972, n19418);
  not g32034 (n_12977, n19417);
  not g32035 (n_12978, n19419);
  and g32036 (n19420, n_12977, n_12978);
  not g32037 (n_12979, n19410);
  not g32038 (n_12980, n19420);
  and g32039 (n19421, n_12979, n_12980);
  not g32040 (n_12981, n19421);
  and g32041 (n19422, \asqrt[37] , n_12981);
  and g32045 (n19426, n_12523, n_12522);
  and g32046 (n19427, \asqrt[8] , n19426);
  not g32047 (n_12982, n19427);
  and g32048 (n19428, n_12521, n_12982);
  not g32049 (n_12983, n19425);
  not g32050 (n_12984, n19428);
  and g32051 (n19429, n_12983, n_12984);
  and g32052 (n19430, n_3474, n_12979);
  and g32053 (n19431, n_12980, n19430);
  not g32054 (n_12985, n19429);
  not g32055 (n_12986, n19431);
  and g32056 (n19432, n_12985, n_12986);
  not g32057 (n_12987, n19422);
  not g32058 (n_12988, n19432);
  and g32059 (n19433, n_12987, n_12988);
  not g32060 (n_12989, n19433);
  and g32061 (n19434, \asqrt[38] , n_12989);
  and g32065 (n19438, n_12531, n_12530);
  and g32066 (n19439, \asqrt[8] , n19438);
  not g32067 (n_12990, n19439);
  and g32068 (n19440, n_12529, n_12990);
  not g32069 (n_12991, n19437);
  not g32070 (n_12992, n19440);
  and g32071 (n19441, n_12991, n_12992);
  and g32072 (n19442, n_3242, n_12987);
  and g32073 (n19443, n_12988, n19442);
  not g32074 (n_12993, n19441);
  not g32075 (n_12994, n19443);
  and g32076 (n19444, n_12993, n_12994);
  not g32077 (n_12995, n19434);
  not g32078 (n_12996, n19444);
  and g32079 (n19445, n_12995, n_12996);
  not g32080 (n_12997, n19445);
  and g32081 (n19446, \asqrt[39] , n_12997);
  and g32085 (n19450, n_12539, n_12538);
  and g32086 (n19451, \asqrt[8] , n19450);
  not g32087 (n_12998, n19451);
  and g32088 (n19452, n_12537, n_12998);
  not g32089 (n_12999, n19449);
  not g32090 (n_13000, n19452);
  and g32091 (n19453, n_12999, n_13000);
  and g32092 (n19454, n_3018, n_12995);
  and g32093 (n19455, n_12996, n19454);
  not g32094 (n_13001, n19453);
  not g32095 (n_13002, n19455);
  and g32096 (n19456, n_13001, n_13002);
  not g32097 (n_13003, n19446);
  not g32098 (n_13004, n19456);
  and g32099 (n19457, n_13003, n_13004);
  not g32100 (n_13005, n19457);
  and g32101 (n19458, \asqrt[40] , n_13005);
  and g32105 (n19462, n_12547, n_12546);
  and g32106 (n19463, \asqrt[8] , n19462);
  not g32107 (n_13006, n19463);
  and g32108 (n19464, n_12545, n_13006);
  not g32109 (n_13007, n19461);
  not g32110 (n_13008, n19464);
  and g32111 (n19465, n_13007, n_13008);
  and g32112 (n19466, n_2802, n_13003);
  and g32113 (n19467, n_13004, n19466);
  not g32114 (n_13009, n19465);
  not g32115 (n_13010, n19467);
  and g32116 (n19468, n_13009, n_13010);
  not g32117 (n_13011, n19458);
  not g32118 (n_13012, n19468);
  and g32119 (n19469, n_13011, n_13012);
  not g32120 (n_13013, n19469);
  and g32121 (n19470, \asqrt[41] , n_13013);
  and g32125 (n19474, n_12555, n_12554);
  and g32126 (n19475, \asqrt[8] , n19474);
  not g32127 (n_13014, n19475);
  and g32128 (n19476, n_12553, n_13014);
  not g32129 (n_13015, n19473);
  not g32130 (n_13016, n19476);
  and g32131 (n19477, n_13015, n_13016);
  and g32132 (n19478, n_2594, n_13011);
  and g32133 (n19479, n_13012, n19478);
  not g32134 (n_13017, n19477);
  not g32135 (n_13018, n19479);
  and g32136 (n19480, n_13017, n_13018);
  not g32137 (n_13019, n19470);
  not g32138 (n_13020, n19480);
  and g32139 (n19481, n_13019, n_13020);
  not g32140 (n_13021, n19481);
  and g32141 (n19482, \asqrt[42] , n_13021);
  and g32145 (n19486, n_12563, n_12562);
  and g32146 (n19487, \asqrt[8] , n19486);
  not g32147 (n_13022, n19487);
  and g32148 (n19488, n_12561, n_13022);
  not g32149 (n_13023, n19485);
  not g32150 (n_13024, n19488);
  and g32151 (n19489, n_13023, n_13024);
  and g32152 (n19490, n_2394, n_13019);
  and g32153 (n19491, n_13020, n19490);
  not g32154 (n_13025, n19489);
  not g32155 (n_13026, n19491);
  and g32156 (n19492, n_13025, n_13026);
  not g32157 (n_13027, n19482);
  not g32158 (n_13028, n19492);
  and g32159 (n19493, n_13027, n_13028);
  not g32160 (n_13029, n19493);
  and g32161 (n19494, \asqrt[43] , n_13029);
  and g32165 (n19498, n_12571, n_12570);
  and g32166 (n19499, \asqrt[8] , n19498);
  not g32167 (n_13030, n19499);
  and g32168 (n19500, n_12569, n_13030);
  not g32169 (n_13031, n19497);
  not g32170 (n_13032, n19500);
  and g32171 (n19501, n_13031, n_13032);
  and g32172 (n19502, n_2202, n_13027);
  and g32173 (n19503, n_13028, n19502);
  not g32174 (n_13033, n19501);
  not g32175 (n_13034, n19503);
  and g32176 (n19504, n_13033, n_13034);
  not g32177 (n_13035, n19494);
  not g32178 (n_13036, n19504);
  and g32179 (n19505, n_13035, n_13036);
  not g32180 (n_13037, n19505);
  and g32181 (n19506, \asqrt[44] , n_13037);
  and g32185 (n19510, n_12579, n_12578);
  and g32186 (n19511, \asqrt[8] , n19510);
  not g32187 (n_13038, n19511);
  and g32188 (n19512, n_12577, n_13038);
  not g32189 (n_13039, n19509);
  not g32190 (n_13040, n19512);
  and g32191 (n19513, n_13039, n_13040);
  and g32192 (n19514, n_2018, n_13035);
  and g32193 (n19515, n_13036, n19514);
  not g32194 (n_13041, n19513);
  not g32195 (n_13042, n19515);
  and g32196 (n19516, n_13041, n_13042);
  not g32197 (n_13043, n19506);
  not g32198 (n_13044, n19516);
  and g32199 (n19517, n_13043, n_13044);
  not g32200 (n_13045, n19517);
  and g32201 (n19518, \asqrt[45] , n_13045);
  and g32205 (n19522, n_12587, n_12586);
  and g32206 (n19523, \asqrt[8] , n19522);
  not g32207 (n_13046, n19523);
  and g32208 (n19524, n_12585, n_13046);
  not g32209 (n_13047, n19521);
  not g32210 (n_13048, n19524);
  and g32211 (n19525, n_13047, n_13048);
  and g32212 (n19526, n_1842, n_13043);
  and g32213 (n19527, n_13044, n19526);
  not g32214 (n_13049, n19525);
  not g32215 (n_13050, n19527);
  and g32216 (n19528, n_13049, n_13050);
  not g32217 (n_13051, n19518);
  not g32218 (n_13052, n19528);
  and g32219 (n19529, n_13051, n_13052);
  not g32220 (n_13053, n19529);
  and g32221 (n19530, \asqrt[46] , n_13053);
  and g32225 (n19534, n_12595, n_12594);
  and g32226 (n19535, \asqrt[8] , n19534);
  not g32227 (n_13054, n19535);
  and g32228 (n19536, n_12593, n_13054);
  not g32229 (n_13055, n19533);
  not g32230 (n_13056, n19536);
  and g32231 (n19537, n_13055, n_13056);
  and g32232 (n19538, n_1674, n_13051);
  and g32233 (n19539, n_13052, n19538);
  not g32234 (n_13057, n19537);
  not g32235 (n_13058, n19539);
  and g32236 (n19540, n_13057, n_13058);
  not g32237 (n_13059, n19530);
  not g32238 (n_13060, n19540);
  and g32239 (n19541, n_13059, n_13060);
  not g32240 (n_13061, n19541);
  and g32241 (n19542, \asqrt[47] , n_13061);
  and g32245 (n19546, n_12603, n_12602);
  and g32246 (n19547, \asqrt[8] , n19546);
  not g32247 (n_13062, n19547);
  and g32248 (n19548, n_12601, n_13062);
  not g32249 (n_13063, n19545);
  not g32250 (n_13064, n19548);
  and g32251 (n19549, n_13063, n_13064);
  and g32252 (n19550, n_1514, n_13059);
  and g32253 (n19551, n_13060, n19550);
  not g32254 (n_13065, n19549);
  not g32255 (n_13066, n19551);
  and g32256 (n19552, n_13065, n_13066);
  not g32257 (n_13067, n19542);
  not g32258 (n_13068, n19552);
  and g32259 (n19553, n_13067, n_13068);
  not g32260 (n_13069, n19553);
  and g32261 (n19554, \asqrt[48] , n_13069);
  and g32265 (n19558, n_12611, n_12610);
  and g32266 (n19559, \asqrt[8] , n19558);
  not g32267 (n_13070, n19559);
  and g32268 (n19560, n_12609, n_13070);
  not g32269 (n_13071, n19557);
  not g32270 (n_13072, n19560);
  and g32271 (n19561, n_13071, n_13072);
  and g32272 (n19562, n_1362, n_13067);
  and g32273 (n19563, n_13068, n19562);
  not g32274 (n_13073, n19561);
  not g32275 (n_13074, n19563);
  and g32276 (n19564, n_13073, n_13074);
  not g32277 (n_13075, n19554);
  not g32278 (n_13076, n19564);
  and g32279 (n19565, n_13075, n_13076);
  not g32280 (n_13077, n19565);
  and g32281 (n19566, \asqrt[49] , n_13077);
  and g32285 (n19570, n_12619, n_12618);
  and g32286 (n19571, \asqrt[8] , n19570);
  not g32287 (n_13078, n19571);
  and g32288 (n19572, n_12617, n_13078);
  not g32289 (n_13079, n19569);
  not g32290 (n_13080, n19572);
  and g32291 (n19573, n_13079, n_13080);
  and g32292 (n19574, n_1218, n_13075);
  and g32293 (n19575, n_13076, n19574);
  not g32294 (n_13081, n19573);
  not g32295 (n_13082, n19575);
  and g32296 (n19576, n_13081, n_13082);
  not g32297 (n_13083, n19566);
  not g32298 (n_13084, n19576);
  and g32299 (n19577, n_13083, n_13084);
  not g32300 (n_13085, n19577);
  and g32301 (n19578, \asqrt[50] , n_13085);
  and g32305 (n19582, n_12627, n_12626);
  and g32306 (n19583, \asqrt[8] , n19582);
  not g32307 (n_13086, n19583);
  and g32308 (n19584, n_12625, n_13086);
  not g32309 (n_13087, n19581);
  not g32310 (n_13088, n19584);
  and g32311 (n19585, n_13087, n_13088);
  and g32312 (n19586, n_1082, n_13083);
  and g32313 (n19587, n_13084, n19586);
  not g32314 (n_13089, n19585);
  not g32315 (n_13090, n19587);
  and g32316 (n19588, n_13089, n_13090);
  not g32317 (n_13091, n19578);
  not g32318 (n_13092, n19588);
  and g32319 (n19589, n_13091, n_13092);
  not g32320 (n_13093, n19589);
  and g32321 (n19590, \asqrt[51] , n_13093);
  and g32325 (n19594, n_12635, n_12634);
  and g32326 (n19595, \asqrt[8] , n19594);
  not g32327 (n_13094, n19595);
  and g32328 (n19596, n_12633, n_13094);
  not g32329 (n_13095, n19593);
  not g32330 (n_13096, n19596);
  and g32331 (n19597, n_13095, n_13096);
  and g32332 (n19598, n_954, n_13091);
  and g32333 (n19599, n_13092, n19598);
  not g32334 (n_13097, n19597);
  not g32335 (n_13098, n19599);
  and g32336 (n19600, n_13097, n_13098);
  not g32337 (n_13099, n19590);
  not g32338 (n_13100, n19600);
  and g32339 (n19601, n_13099, n_13100);
  not g32340 (n_13101, n19601);
  and g32341 (n19602, \asqrt[52] , n_13101);
  and g32345 (n19606, n_12643, n_12642);
  and g32346 (n19607, \asqrt[8] , n19606);
  not g32347 (n_13102, n19607);
  and g32348 (n19608, n_12641, n_13102);
  not g32349 (n_13103, n19605);
  not g32350 (n_13104, n19608);
  and g32351 (n19609, n_13103, n_13104);
  and g32352 (n19610, n_834, n_13099);
  and g32353 (n19611, n_13100, n19610);
  not g32354 (n_13105, n19609);
  not g32355 (n_13106, n19611);
  and g32356 (n19612, n_13105, n_13106);
  not g32357 (n_13107, n19602);
  not g32358 (n_13108, n19612);
  and g32359 (n19613, n_13107, n_13108);
  not g32360 (n_13109, n19613);
  and g32361 (n19614, \asqrt[53] , n_13109);
  and g32365 (n19618, n_12651, n_12650);
  and g32366 (n19619, \asqrt[8] , n19618);
  not g32367 (n_13110, n19619);
  and g32368 (n19620, n_12649, n_13110);
  not g32369 (n_13111, n19617);
  not g32370 (n_13112, n19620);
  and g32371 (n19621, n_13111, n_13112);
  and g32372 (n19622, n_722, n_13107);
  and g32373 (n19623, n_13108, n19622);
  not g32374 (n_13113, n19621);
  not g32375 (n_13114, n19623);
  and g32376 (n19624, n_13113, n_13114);
  not g32377 (n_13115, n19614);
  not g32378 (n_13116, n19624);
  and g32379 (n19625, n_13115, n_13116);
  not g32380 (n_13117, n19625);
  and g32381 (n19626, \asqrt[54] , n_13117);
  and g32385 (n19630, n_12659, n_12658);
  and g32386 (n19631, \asqrt[8] , n19630);
  not g32387 (n_13118, n19631);
  and g32388 (n19632, n_12657, n_13118);
  not g32389 (n_13119, n19629);
  not g32390 (n_13120, n19632);
  and g32391 (n19633, n_13119, n_13120);
  and g32392 (n19634, n_618, n_13115);
  and g32393 (n19635, n_13116, n19634);
  not g32394 (n_13121, n19633);
  not g32395 (n_13122, n19635);
  and g32396 (n19636, n_13121, n_13122);
  not g32397 (n_13123, n19626);
  not g32398 (n_13124, n19636);
  and g32399 (n19637, n_13123, n_13124);
  not g32400 (n_13125, n19637);
  and g32401 (n19638, \asqrt[55] , n_13125);
  and g32405 (n19642, n_12667, n_12666);
  and g32406 (n19643, \asqrt[8] , n19642);
  not g32407 (n_13126, n19643);
  and g32408 (n19644, n_12665, n_13126);
  not g32409 (n_13127, n19641);
  not g32410 (n_13128, n19644);
  and g32411 (n19645, n_13127, n_13128);
  and g32412 (n19646, n_522, n_13123);
  and g32413 (n19647, n_13124, n19646);
  not g32414 (n_13129, n19645);
  not g32415 (n_13130, n19647);
  and g32416 (n19648, n_13129, n_13130);
  not g32417 (n_13131, n19638);
  not g32418 (n_13132, n19648);
  and g32419 (n19649, n_13131, n_13132);
  not g32420 (n_13133, n19649);
  and g32421 (n19650, \asqrt[56] , n_13133);
  and g32425 (n19654, n_12675, n_12674);
  and g32426 (n19655, \asqrt[8] , n19654);
  not g32427 (n_13134, n19655);
  and g32428 (n19656, n_12673, n_13134);
  not g32429 (n_13135, n19653);
  not g32430 (n_13136, n19656);
  and g32431 (n19657, n_13135, n_13136);
  and g32432 (n19658, n_434, n_13131);
  and g32433 (n19659, n_13132, n19658);
  not g32434 (n_13137, n19657);
  not g32435 (n_13138, n19659);
  and g32436 (n19660, n_13137, n_13138);
  not g32437 (n_13139, n19650);
  not g32438 (n_13140, n19660);
  and g32439 (n19661, n_13139, n_13140);
  not g32440 (n_13141, n19661);
  and g32441 (n19662, \asqrt[57] , n_13141);
  and g32442 (n19663, n_354, n_13139);
  and g32443 (n19664, n_13140, n19663);
  and g32447 (n19668, n_12683, n_12681);
  and g32448 (n19669, \asqrt[8] , n19668);
  not g32449 (n_13142, n19669);
  and g32450 (n19670, n_12682, n_13142);
  not g32451 (n_13143, n19667);
  not g32452 (n_13144, n19670);
  and g32453 (n19671, n_13143, n_13144);
  not g32454 (n_13145, n19664);
  not g32455 (n_13146, n19671);
  and g32456 (n19672, n_13145, n_13146);
  not g32457 (n_13147, n19662);
  not g32458 (n_13148, n19672);
  and g32459 (n19673, n_13147, n_13148);
  not g32460 (n_13149, n19673);
  and g32461 (n19674, \asqrt[58] , n_13149);
  and g32465 (n19678, n_12691, n_12690);
  and g32466 (n19679, \asqrt[8] , n19678);
  not g32467 (n_13150, n19679);
  and g32468 (n19680, n_12689, n_13150);
  not g32469 (n_13151, n19677);
  not g32470 (n_13152, n19680);
  and g32471 (n19681, n_13151, n_13152);
  and g32472 (n19682, n_282, n_13147);
  and g32473 (n19683, n_13148, n19682);
  not g32474 (n_13153, n19681);
  not g32475 (n_13154, n19683);
  and g32476 (n19684, n_13153, n_13154);
  not g32477 (n_13155, n19674);
  not g32478 (n_13156, n19684);
  and g32479 (n19685, n_13155, n_13156);
  not g32480 (n_13157, n19685);
  and g32481 (n19686, \asqrt[59] , n_13157);
  and g32485 (n19690, n_12699, n_12698);
  and g32486 (n19691, \asqrt[8] , n19690);
  not g32487 (n_13158, n19691);
  and g32488 (n19692, n_12697, n_13158);
  not g32489 (n_13159, n19689);
  not g32490 (n_13160, n19692);
  and g32491 (n19693, n_13159, n_13160);
  and g32492 (n19694, n_218, n_13155);
  and g32493 (n19695, n_13156, n19694);
  not g32494 (n_13161, n19693);
  not g32495 (n_13162, n19695);
  and g32496 (n19696, n_13161, n_13162);
  not g32497 (n_13163, n19686);
  not g32498 (n_13164, n19696);
  and g32499 (n19697, n_13163, n_13164);
  not g32500 (n_13165, n19697);
  and g32501 (n19698, \asqrt[60] , n_13165);
  and g32505 (n19702, n_12707, n_12706);
  and g32506 (n19703, \asqrt[8] , n19702);
  not g32507 (n_13166, n19703);
  and g32508 (n19704, n_12705, n_13166);
  not g32509 (n_13167, n19701);
  not g32510 (n_13168, n19704);
  and g32511 (n19705, n_13167, n_13168);
  and g32512 (n19706, n_162, n_13163);
  and g32513 (n19707, n_13164, n19706);
  not g32514 (n_13169, n19705);
  not g32515 (n_13170, n19707);
  and g32516 (n19708, n_13169, n_13170);
  not g32517 (n_13171, n19698);
  not g32518 (n_13172, n19708);
  and g32519 (n19709, n_13171, n_13172);
  not g32520 (n_13173, n19709);
  and g32521 (n19710, \asqrt[61] , n_13173);
  and g32525 (n19714, n_12715, n_12714);
  and g32526 (n19715, \asqrt[8] , n19714);
  not g32527 (n_13174, n19715);
  and g32528 (n19716, n_12713, n_13174);
  not g32529 (n_13175, n19713);
  not g32530 (n_13176, n19716);
  and g32531 (n19717, n_13175, n_13176);
  and g32532 (n19718, n_115, n_13171);
  and g32533 (n19719, n_13172, n19718);
  not g32534 (n_13177, n19717);
  not g32535 (n_13178, n19719);
  and g32536 (n19720, n_13177, n_13178);
  not g32537 (n_13179, n19710);
  not g32538 (n_13180, n19720);
  and g32539 (n19721, n_13179, n_13180);
  not g32540 (n_13181, n19721);
  and g32541 (n19722, \asqrt[62] , n_13181);
  and g32545 (n19726, n_12723, n_12722);
  and g32546 (n19727, \asqrt[8] , n19726);
  not g32547 (n_13182, n19727);
  and g32548 (n19728, n_12721, n_13182);
  not g32549 (n_13183, n19725);
  not g32550 (n_13184, n19728);
  and g32551 (n19729, n_13183, n_13184);
  and g32552 (n19730, n_76, n_13179);
  and g32553 (n19731, n_13180, n19730);
  not g32554 (n_13185, n19729);
  not g32555 (n_13186, n19731);
  and g32556 (n19732, n_13185, n_13186);
  not g32557 (n_13187, n19722);
  not g32558 (n_13188, n19732);
  and g32559 (n19733, n_13187, n_13188);
  and g32563 (n19737, n_12731, n_12730);
  and g32564 (n19738, \asqrt[8] , n19737);
  not g32565 (n_13189, n19738);
  and g32566 (n19739, n_12729, n_13189);
  not g32567 (n_13190, n19736);
  not g32568 (n_13191, n19739);
  and g32569 (n19740, n_13190, n_13191);
  and g32570 (n19741, n_12738, n_12737);
  and g32571 (n19742, \asqrt[8] , n19741);
  not g32574 (n_13193, n19740);
  not g32576 (n_13194, n19733);
  not g32578 (n_13195, n19745);
  and g32579 (n19746, n_21, n_13195);
  and g32580 (n19747, n_13187, n19740);
  and g32581 (n19748, n_13188, n19747);
  and g32582 (n19749, n_12737, \asqrt[8] );
  not g32583 (n_13196, n19749);
  and g32584 (n19750, n19053, n_13196);
  not g32585 (n_13197, n19741);
  and g32586 (n19751, \asqrt[63] , n_13197);
  not g32587 (n_13198, n19750);
  and g32588 (n19752, n_13198, n19751);
  not g32594 (n_13199, n19752);
  not g32595 (n_13200, n19757);
  not g32597 (n_13201, n19748);
  and g32601 (n19761, \a[14] , \asqrt[7] );
  not g32602 (n_13206, \a[12] );
  not g32603 (n_13207, \a[13] );
  and g32604 (n19762, n_13206, n_13207);
  and g32605 (n19763, n_12750, n19762);
  not g32606 (n_13208, n19761);
  not g32607 (n_13209, n19763);
  and g32608 (n19764, n_13208, n_13209);
  not g32609 (n_13210, n19764);
  and g32610 (n19765, \asqrt[8] , n_13210);
  and g32616 (n19771, n_12750, \asqrt[7] );
  not g32617 (n_13211, n19771);
  and g32618 (n19772, \a[15] , n_13211);
  and g32619 (n19773, n19082, \asqrt[7] );
  not g32620 (n_13212, n19772);
  not g32621 (n_13213, n19773);
  and g32622 (n19774, n_13212, n_13213);
  not g32623 (n_13214, n19770);
  and g32624 (n19775, n_13214, n19774);
  not g32625 (n_13215, n19765);
  not g32626 (n_13216, n19775);
  and g32627 (n19776, n_13215, n_13216);
  not g32628 (n_13217, n19776);
  and g32629 (n19777, \asqrt[9] , n_13217);
  not g32630 (n_13218, \asqrt[9] );
  and g32631 (n19778, n_13218, n_13215);
  and g32632 (n19779, n_13216, n19778);
  not g32636 (n_13219, n19746);
  not g32638 (n_13220, n19783);
  and g32639 (n19784, n_13213, n_13220);
  not g32640 (n_13221, n19784);
  and g32641 (n19785, \a[16] , n_13221);
  and g32642 (n19786, n_12302, n_13220);
  and g32643 (n19787, n_13213, n19786);
  not g32644 (n_13222, n19785);
  not g32645 (n_13223, n19787);
  and g32646 (n19788, n_13222, n_13223);
  not g32647 (n_13224, n19779);
  not g32648 (n_13225, n19788);
  and g32649 (n19789, n_13224, n_13225);
  not g32650 (n_13226, n19777);
  not g32651 (n_13227, n19789);
  and g32652 (n19790, n_13226, n_13227);
  not g32653 (n_13228, n19790);
  and g32654 (n19791, \asqrt[10] , n_13228);
  and g32655 (n19792, n_12759, n_12758);
  not g32656 (n_13229, n19094);
  and g32657 (n19793, n_13229, n19792);
  and g32658 (n19794, \asqrt[7] , n19793);
  and g32659 (n19795, \asqrt[7] , n19792);
  not g32660 (n_13230, n19795);
  and g32661 (n19796, n19094, n_13230);
  not g32662 (n_13231, n19794);
  not g32663 (n_13232, n19796);
  and g32664 (n19797, n_13231, n_13232);
  and g32665 (n19798, n_12762, n_13226);
  and g32666 (n19799, n_13227, n19798);
  not g32667 (n_13233, n19797);
  not g32668 (n_13234, n19799);
  and g32669 (n19800, n_13233, n_13234);
  not g32670 (n_13235, n19791);
  not g32671 (n_13236, n19800);
  and g32672 (n19801, n_13235, n_13236);
  not g32673 (n_13237, n19801);
  and g32674 (n19802, \asqrt[11] , n_13237);
  and g32678 (n19806, n_12770, n_12768);
  and g32679 (n19807, \asqrt[7] , n19806);
  not g32680 (n_13238, n19807);
  and g32681 (n19808, n_12769, n_13238);
  not g32682 (n_13239, n19805);
  not g32683 (n_13240, n19808);
  and g32684 (n19809, n_13239, n_13240);
  and g32685 (n19810, n_12314, n_13235);
  and g32686 (n19811, n_13236, n19810);
  not g32687 (n_13241, n19809);
  not g32688 (n_13242, n19811);
  and g32689 (n19812, n_13241, n_13242);
  not g32690 (n_13243, n19802);
  not g32691 (n_13244, n19812);
  and g32692 (n19813, n_13243, n_13244);
  not g32693 (n_13245, n19813);
  and g32694 (n19814, \asqrt[12] , n_13245);
  and g32698 (n19818, n_12779, n_12778);
  and g32699 (n19819, \asqrt[7] , n19818);
  not g32700 (n_13246, n19819);
  and g32701 (n19820, n_12777, n_13246);
  not g32702 (n_13247, n19817);
  not g32703 (n_13248, n19820);
  and g32704 (n19821, n_13247, n_13248);
  and g32705 (n19822, n_11874, n_13243);
  and g32706 (n19823, n_13244, n19822);
  not g32707 (n_13249, n19821);
  not g32708 (n_13250, n19823);
  and g32709 (n19824, n_13249, n_13250);
  not g32710 (n_13251, n19814);
  not g32711 (n_13252, n19824);
  and g32712 (n19825, n_13251, n_13252);
  not g32713 (n_13253, n19825);
  and g32714 (n19826, \asqrt[13] , n_13253);
  and g32718 (n19830, n_12787, n_12786);
  and g32719 (n19831, \asqrt[7] , n19830);
  not g32720 (n_13254, n19831);
  and g32721 (n19832, n_12785, n_13254);
  not g32722 (n_13255, n19829);
  not g32723 (n_13256, n19832);
  and g32724 (n19833, n_13255, n_13256);
  and g32725 (n19834, n_11442, n_13251);
  and g32726 (n19835, n_13252, n19834);
  not g32727 (n_13257, n19833);
  not g32728 (n_13258, n19835);
  and g32729 (n19836, n_13257, n_13258);
  not g32730 (n_13259, n19826);
  not g32731 (n_13260, n19836);
  and g32732 (n19837, n_13259, n_13260);
  not g32733 (n_13261, n19837);
  and g32734 (n19838, \asqrt[14] , n_13261);
  and g32738 (n19842, n_12795, n_12794);
  and g32739 (n19843, \asqrt[7] , n19842);
  not g32740 (n_13262, n19843);
  and g32741 (n19844, n_12793, n_13262);
  not g32742 (n_13263, n19841);
  not g32743 (n_13264, n19844);
  and g32744 (n19845, n_13263, n_13264);
  and g32745 (n19846, n_11018, n_13259);
  and g32746 (n19847, n_13260, n19846);
  not g32747 (n_13265, n19845);
  not g32748 (n_13266, n19847);
  and g32749 (n19848, n_13265, n_13266);
  not g32750 (n_13267, n19838);
  not g32751 (n_13268, n19848);
  and g32752 (n19849, n_13267, n_13268);
  not g32753 (n_13269, n19849);
  and g32754 (n19850, \asqrt[15] , n_13269);
  and g32758 (n19854, n_12803, n_12802);
  and g32759 (n19855, \asqrt[7] , n19854);
  not g32760 (n_13270, n19855);
  and g32761 (n19856, n_12801, n_13270);
  not g32762 (n_13271, n19853);
  not g32763 (n_13272, n19856);
  and g32764 (n19857, n_13271, n_13272);
  and g32765 (n19858, n_10602, n_13267);
  and g32766 (n19859, n_13268, n19858);
  not g32767 (n_13273, n19857);
  not g32768 (n_13274, n19859);
  and g32769 (n19860, n_13273, n_13274);
  not g32770 (n_13275, n19850);
  not g32771 (n_13276, n19860);
  and g32772 (n19861, n_13275, n_13276);
  not g32773 (n_13277, n19861);
  and g32774 (n19862, \asqrt[16] , n_13277);
  and g32778 (n19866, n_12811, n_12810);
  and g32779 (n19867, \asqrt[7] , n19866);
  not g32780 (n_13278, n19867);
  and g32781 (n19868, n_12809, n_13278);
  not g32782 (n_13279, n19865);
  not g32783 (n_13280, n19868);
  and g32784 (n19869, n_13279, n_13280);
  and g32785 (n19870, n_10194, n_13275);
  and g32786 (n19871, n_13276, n19870);
  not g32787 (n_13281, n19869);
  not g32788 (n_13282, n19871);
  and g32789 (n19872, n_13281, n_13282);
  not g32790 (n_13283, n19862);
  not g32791 (n_13284, n19872);
  and g32792 (n19873, n_13283, n_13284);
  not g32793 (n_13285, n19873);
  and g32794 (n19874, \asqrt[17] , n_13285);
  and g32798 (n19878, n_12819, n_12818);
  and g32799 (n19879, \asqrt[7] , n19878);
  not g32800 (n_13286, n19879);
  and g32801 (n19880, n_12817, n_13286);
  not g32802 (n_13287, n19877);
  not g32803 (n_13288, n19880);
  and g32804 (n19881, n_13287, n_13288);
  and g32805 (n19882, n_9794, n_13283);
  and g32806 (n19883, n_13284, n19882);
  not g32807 (n_13289, n19881);
  not g32808 (n_13290, n19883);
  and g32809 (n19884, n_13289, n_13290);
  not g32810 (n_13291, n19874);
  not g32811 (n_13292, n19884);
  and g32812 (n19885, n_13291, n_13292);
  not g32813 (n_13293, n19885);
  and g32814 (n19886, \asqrt[18] , n_13293);
  and g32818 (n19890, n_12827, n_12826);
  and g32819 (n19891, \asqrt[7] , n19890);
  not g32820 (n_13294, n19891);
  and g32821 (n19892, n_12825, n_13294);
  not g32822 (n_13295, n19889);
  not g32823 (n_13296, n19892);
  and g32824 (n19893, n_13295, n_13296);
  and g32825 (n19894, n_9402, n_13291);
  and g32826 (n19895, n_13292, n19894);
  not g32827 (n_13297, n19893);
  not g32828 (n_13298, n19895);
  and g32829 (n19896, n_13297, n_13298);
  not g32830 (n_13299, n19886);
  not g32831 (n_13300, n19896);
  and g32832 (n19897, n_13299, n_13300);
  not g32833 (n_13301, n19897);
  and g32834 (n19898, \asqrt[19] , n_13301);
  and g32838 (n19902, n_12835, n_12834);
  and g32839 (n19903, \asqrt[7] , n19902);
  not g32840 (n_13302, n19903);
  and g32841 (n19904, n_12833, n_13302);
  not g32842 (n_13303, n19901);
  not g32843 (n_13304, n19904);
  and g32844 (n19905, n_13303, n_13304);
  and g32845 (n19906, n_9018, n_13299);
  and g32846 (n19907, n_13300, n19906);
  not g32847 (n_13305, n19905);
  not g32848 (n_13306, n19907);
  and g32849 (n19908, n_13305, n_13306);
  not g32850 (n_13307, n19898);
  not g32851 (n_13308, n19908);
  and g32852 (n19909, n_13307, n_13308);
  not g32853 (n_13309, n19909);
  and g32854 (n19910, \asqrt[20] , n_13309);
  and g32858 (n19914, n_12843, n_12842);
  and g32859 (n19915, \asqrt[7] , n19914);
  not g32860 (n_13310, n19915);
  and g32861 (n19916, n_12841, n_13310);
  not g32862 (n_13311, n19913);
  not g32863 (n_13312, n19916);
  and g32864 (n19917, n_13311, n_13312);
  and g32865 (n19918, n_8642, n_13307);
  and g32866 (n19919, n_13308, n19918);
  not g32867 (n_13313, n19917);
  not g32868 (n_13314, n19919);
  and g32869 (n19920, n_13313, n_13314);
  not g32870 (n_13315, n19910);
  not g32871 (n_13316, n19920);
  and g32872 (n19921, n_13315, n_13316);
  not g32873 (n_13317, n19921);
  and g32874 (n19922, \asqrt[21] , n_13317);
  and g32878 (n19926, n_12851, n_12850);
  and g32879 (n19927, \asqrt[7] , n19926);
  not g32880 (n_13318, n19927);
  and g32881 (n19928, n_12849, n_13318);
  not g32882 (n_13319, n19925);
  not g32883 (n_13320, n19928);
  and g32884 (n19929, n_13319, n_13320);
  and g32885 (n19930, n_8274, n_13315);
  and g32886 (n19931, n_13316, n19930);
  not g32887 (n_13321, n19929);
  not g32888 (n_13322, n19931);
  and g32889 (n19932, n_13321, n_13322);
  not g32890 (n_13323, n19922);
  not g32891 (n_13324, n19932);
  and g32892 (n19933, n_13323, n_13324);
  not g32893 (n_13325, n19933);
  and g32894 (n19934, \asqrt[22] , n_13325);
  and g32898 (n19938, n_12859, n_12858);
  and g32899 (n19939, \asqrt[7] , n19938);
  not g32900 (n_13326, n19939);
  and g32901 (n19940, n_12857, n_13326);
  not g32902 (n_13327, n19937);
  not g32903 (n_13328, n19940);
  and g32904 (n19941, n_13327, n_13328);
  and g32905 (n19942, n_7914, n_13323);
  and g32906 (n19943, n_13324, n19942);
  not g32907 (n_13329, n19941);
  not g32908 (n_13330, n19943);
  and g32909 (n19944, n_13329, n_13330);
  not g32910 (n_13331, n19934);
  not g32911 (n_13332, n19944);
  and g32912 (n19945, n_13331, n_13332);
  not g32913 (n_13333, n19945);
  and g32914 (n19946, \asqrt[23] , n_13333);
  and g32918 (n19950, n_12867, n_12866);
  and g32919 (n19951, \asqrt[7] , n19950);
  not g32920 (n_13334, n19951);
  and g32921 (n19952, n_12865, n_13334);
  not g32922 (n_13335, n19949);
  not g32923 (n_13336, n19952);
  and g32924 (n19953, n_13335, n_13336);
  and g32925 (n19954, n_7562, n_13331);
  and g32926 (n19955, n_13332, n19954);
  not g32927 (n_13337, n19953);
  not g32928 (n_13338, n19955);
  and g32929 (n19956, n_13337, n_13338);
  not g32930 (n_13339, n19946);
  not g32931 (n_13340, n19956);
  and g32932 (n19957, n_13339, n_13340);
  not g32933 (n_13341, n19957);
  and g32934 (n19958, \asqrt[24] , n_13341);
  and g32938 (n19962, n_12875, n_12874);
  and g32939 (n19963, \asqrt[7] , n19962);
  not g32940 (n_13342, n19963);
  and g32941 (n19964, n_12873, n_13342);
  not g32942 (n_13343, n19961);
  not g32943 (n_13344, n19964);
  and g32944 (n19965, n_13343, n_13344);
  and g32945 (n19966, n_7218, n_13339);
  and g32946 (n19967, n_13340, n19966);
  not g32947 (n_13345, n19965);
  not g32948 (n_13346, n19967);
  and g32949 (n19968, n_13345, n_13346);
  not g32950 (n_13347, n19958);
  not g32951 (n_13348, n19968);
  and g32952 (n19969, n_13347, n_13348);
  not g32953 (n_13349, n19969);
  and g32954 (n19970, \asqrt[25] , n_13349);
  and g32958 (n19974, n_12883, n_12882);
  and g32959 (n19975, \asqrt[7] , n19974);
  not g32960 (n_13350, n19975);
  and g32961 (n19976, n_12881, n_13350);
  not g32962 (n_13351, n19973);
  not g32963 (n_13352, n19976);
  and g32964 (n19977, n_13351, n_13352);
  and g32965 (n19978, n_6882, n_13347);
  and g32966 (n19979, n_13348, n19978);
  not g32967 (n_13353, n19977);
  not g32968 (n_13354, n19979);
  and g32969 (n19980, n_13353, n_13354);
  not g32970 (n_13355, n19970);
  not g32971 (n_13356, n19980);
  and g32972 (n19981, n_13355, n_13356);
  not g32973 (n_13357, n19981);
  and g32974 (n19982, \asqrt[26] , n_13357);
  and g32978 (n19986, n_12891, n_12890);
  and g32979 (n19987, \asqrt[7] , n19986);
  not g32980 (n_13358, n19987);
  and g32981 (n19988, n_12889, n_13358);
  not g32982 (n_13359, n19985);
  not g32983 (n_13360, n19988);
  and g32984 (n19989, n_13359, n_13360);
  and g32985 (n19990, n_6554, n_13355);
  and g32986 (n19991, n_13356, n19990);
  not g32987 (n_13361, n19989);
  not g32988 (n_13362, n19991);
  and g32989 (n19992, n_13361, n_13362);
  not g32990 (n_13363, n19982);
  not g32991 (n_13364, n19992);
  and g32992 (n19993, n_13363, n_13364);
  not g32993 (n_13365, n19993);
  and g32994 (n19994, \asqrt[27] , n_13365);
  and g32998 (n19998, n_12899, n_12898);
  and g32999 (n19999, \asqrt[7] , n19998);
  not g33000 (n_13366, n19999);
  and g33001 (n20000, n_12897, n_13366);
  not g33002 (n_13367, n19997);
  not g33003 (n_13368, n20000);
  and g33004 (n20001, n_13367, n_13368);
  and g33005 (n20002, n_6234, n_13363);
  and g33006 (n20003, n_13364, n20002);
  not g33007 (n_13369, n20001);
  not g33008 (n_13370, n20003);
  and g33009 (n20004, n_13369, n_13370);
  not g33010 (n_13371, n19994);
  not g33011 (n_13372, n20004);
  and g33012 (n20005, n_13371, n_13372);
  not g33013 (n_13373, n20005);
  and g33014 (n20006, \asqrt[28] , n_13373);
  and g33018 (n20010, n_12907, n_12906);
  and g33019 (n20011, \asqrt[7] , n20010);
  not g33020 (n_13374, n20011);
  and g33021 (n20012, n_12905, n_13374);
  not g33022 (n_13375, n20009);
  not g33023 (n_13376, n20012);
  and g33024 (n20013, n_13375, n_13376);
  and g33025 (n20014, n_5922, n_13371);
  and g33026 (n20015, n_13372, n20014);
  not g33027 (n_13377, n20013);
  not g33028 (n_13378, n20015);
  and g33029 (n20016, n_13377, n_13378);
  not g33030 (n_13379, n20006);
  not g33031 (n_13380, n20016);
  and g33032 (n20017, n_13379, n_13380);
  not g33033 (n_13381, n20017);
  and g33034 (n20018, \asqrt[29] , n_13381);
  and g33038 (n20022, n_12915, n_12914);
  and g33039 (n20023, \asqrt[7] , n20022);
  not g33040 (n_13382, n20023);
  and g33041 (n20024, n_12913, n_13382);
  not g33042 (n_13383, n20021);
  not g33043 (n_13384, n20024);
  and g33044 (n20025, n_13383, n_13384);
  and g33045 (n20026, n_5618, n_13379);
  and g33046 (n20027, n_13380, n20026);
  not g33047 (n_13385, n20025);
  not g33048 (n_13386, n20027);
  and g33049 (n20028, n_13385, n_13386);
  not g33050 (n_13387, n20018);
  not g33051 (n_13388, n20028);
  and g33052 (n20029, n_13387, n_13388);
  not g33053 (n_13389, n20029);
  and g33054 (n20030, \asqrt[30] , n_13389);
  and g33058 (n20034, n_12923, n_12922);
  and g33059 (n20035, \asqrt[7] , n20034);
  not g33060 (n_13390, n20035);
  and g33061 (n20036, n_12921, n_13390);
  not g33062 (n_13391, n20033);
  not g33063 (n_13392, n20036);
  and g33064 (n20037, n_13391, n_13392);
  and g33065 (n20038, n_5322, n_13387);
  and g33066 (n20039, n_13388, n20038);
  not g33067 (n_13393, n20037);
  not g33068 (n_13394, n20039);
  and g33069 (n20040, n_13393, n_13394);
  not g33070 (n_13395, n20030);
  not g33071 (n_13396, n20040);
  and g33072 (n20041, n_13395, n_13396);
  not g33073 (n_13397, n20041);
  and g33074 (n20042, \asqrt[31] , n_13397);
  and g33078 (n20046, n_12931, n_12930);
  and g33079 (n20047, \asqrt[7] , n20046);
  not g33080 (n_13398, n20047);
  and g33081 (n20048, n_12929, n_13398);
  not g33082 (n_13399, n20045);
  not g33083 (n_13400, n20048);
  and g33084 (n20049, n_13399, n_13400);
  and g33085 (n20050, n_5034, n_13395);
  and g33086 (n20051, n_13396, n20050);
  not g33087 (n_13401, n20049);
  not g33088 (n_13402, n20051);
  and g33089 (n20052, n_13401, n_13402);
  not g33090 (n_13403, n20042);
  not g33091 (n_13404, n20052);
  and g33092 (n20053, n_13403, n_13404);
  not g33093 (n_13405, n20053);
  and g33094 (n20054, \asqrt[32] , n_13405);
  and g33098 (n20058, n_12939, n_12938);
  and g33099 (n20059, \asqrt[7] , n20058);
  not g33100 (n_13406, n20059);
  and g33101 (n20060, n_12937, n_13406);
  not g33102 (n_13407, n20057);
  not g33103 (n_13408, n20060);
  and g33104 (n20061, n_13407, n_13408);
  and g33105 (n20062, n_4754, n_13403);
  and g33106 (n20063, n_13404, n20062);
  not g33107 (n_13409, n20061);
  not g33108 (n_13410, n20063);
  and g33109 (n20064, n_13409, n_13410);
  not g33110 (n_13411, n20054);
  not g33111 (n_13412, n20064);
  and g33112 (n20065, n_13411, n_13412);
  not g33113 (n_13413, n20065);
  and g33114 (n20066, \asqrt[33] , n_13413);
  and g33118 (n20070, n_12947, n_12946);
  and g33119 (n20071, \asqrt[7] , n20070);
  not g33120 (n_13414, n20071);
  and g33121 (n20072, n_12945, n_13414);
  not g33122 (n_13415, n20069);
  not g33123 (n_13416, n20072);
  and g33124 (n20073, n_13415, n_13416);
  and g33125 (n20074, n_4482, n_13411);
  and g33126 (n20075, n_13412, n20074);
  not g33127 (n_13417, n20073);
  not g33128 (n_13418, n20075);
  and g33129 (n20076, n_13417, n_13418);
  not g33130 (n_13419, n20066);
  not g33131 (n_13420, n20076);
  and g33132 (n20077, n_13419, n_13420);
  not g33133 (n_13421, n20077);
  and g33134 (n20078, \asqrt[34] , n_13421);
  and g33138 (n20082, n_12955, n_12954);
  and g33139 (n20083, \asqrt[7] , n20082);
  not g33140 (n_13422, n20083);
  and g33141 (n20084, n_12953, n_13422);
  not g33142 (n_13423, n20081);
  not g33143 (n_13424, n20084);
  and g33144 (n20085, n_13423, n_13424);
  and g33145 (n20086, n_4218, n_13419);
  and g33146 (n20087, n_13420, n20086);
  not g33147 (n_13425, n20085);
  not g33148 (n_13426, n20087);
  and g33149 (n20088, n_13425, n_13426);
  not g33150 (n_13427, n20078);
  not g33151 (n_13428, n20088);
  and g33152 (n20089, n_13427, n_13428);
  not g33153 (n_13429, n20089);
  and g33154 (n20090, \asqrt[35] , n_13429);
  and g33158 (n20094, n_12963, n_12962);
  and g33159 (n20095, \asqrt[7] , n20094);
  not g33160 (n_13430, n20095);
  and g33161 (n20096, n_12961, n_13430);
  not g33162 (n_13431, n20093);
  not g33163 (n_13432, n20096);
  and g33164 (n20097, n_13431, n_13432);
  and g33165 (n20098, n_3962, n_13427);
  and g33166 (n20099, n_13428, n20098);
  not g33167 (n_13433, n20097);
  not g33168 (n_13434, n20099);
  and g33169 (n20100, n_13433, n_13434);
  not g33170 (n_13435, n20090);
  not g33171 (n_13436, n20100);
  and g33172 (n20101, n_13435, n_13436);
  not g33173 (n_13437, n20101);
  and g33174 (n20102, \asqrt[36] , n_13437);
  and g33178 (n20106, n_12971, n_12970);
  and g33179 (n20107, \asqrt[7] , n20106);
  not g33180 (n_13438, n20107);
  and g33181 (n20108, n_12969, n_13438);
  not g33182 (n_13439, n20105);
  not g33183 (n_13440, n20108);
  and g33184 (n20109, n_13439, n_13440);
  and g33185 (n20110, n_3714, n_13435);
  and g33186 (n20111, n_13436, n20110);
  not g33187 (n_13441, n20109);
  not g33188 (n_13442, n20111);
  and g33189 (n20112, n_13441, n_13442);
  not g33190 (n_13443, n20102);
  not g33191 (n_13444, n20112);
  and g33192 (n20113, n_13443, n_13444);
  not g33193 (n_13445, n20113);
  and g33194 (n20114, \asqrt[37] , n_13445);
  and g33198 (n20118, n_12979, n_12978);
  and g33199 (n20119, \asqrt[7] , n20118);
  not g33200 (n_13446, n20119);
  and g33201 (n20120, n_12977, n_13446);
  not g33202 (n_13447, n20117);
  not g33203 (n_13448, n20120);
  and g33204 (n20121, n_13447, n_13448);
  and g33205 (n20122, n_3474, n_13443);
  and g33206 (n20123, n_13444, n20122);
  not g33207 (n_13449, n20121);
  not g33208 (n_13450, n20123);
  and g33209 (n20124, n_13449, n_13450);
  not g33210 (n_13451, n20114);
  not g33211 (n_13452, n20124);
  and g33212 (n20125, n_13451, n_13452);
  not g33213 (n_13453, n20125);
  and g33214 (n20126, \asqrt[38] , n_13453);
  and g33218 (n20130, n_12987, n_12986);
  and g33219 (n20131, \asqrt[7] , n20130);
  not g33220 (n_13454, n20131);
  and g33221 (n20132, n_12985, n_13454);
  not g33222 (n_13455, n20129);
  not g33223 (n_13456, n20132);
  and g33224 (n20133, n_13455, n_13456);
  and g33225 (n20134, n_3242, n_13451);
  and g33226 (n20135, n_13452, n20134);
  not g33227 (n_13457, n20133);
  not g33228 (n_13458, n20135);
  and g33229 (n20136, n_13457, n_13458);
  not g33230 (n_13459, n20126);
  not g33231 (n_13460, n20136);
  and g33232 (n20137, n_13459, n_13460);
  not g33233 (n_13461, n20137);
  and g33234 (n20138, \asqrt[39] , n_13461);
  and g33238 (n20142, n_12995, n_12994);
  and g33239 (n20143, \asqrt[7] , n20142);
  not g33240 (n_13462, n20143);
  and g33241 (n20144, n_12993, n_13462);
  not g33242 (n_13463, n20141);
  not g33243 (n_13464, n20144);
  and g33244 (n20145, n_13463, n_13464);
  and g33245 (n20146, n_3018, n_13459);
  and g33246 (n20147, n_13460, n20146);
  not g33247 (n_13465, n20145);
  not g33248 (n_13466, n20147);
  and g33249 (n20148, n_13465, n_13466);
  not g33250 (n_13467, n20138);
  not g33251 (n_13468, n20148);
  and g33252 (n20149, n_13467, n_13468);
  not g33253 (n_13469, n20149);
  and g33254 (n20150, \asqrt[40] , n_13469);
  and g33258 (n20154, n_13003, n_13002);
  and g33259 (n20155, \asqrt[7] , n20154);
  not g33260 (n_13470, n20155);
  and g33261 (n20156, n_13001, n_13470);
  not g33262 (n_13471, n20153);
  not g33263 (n_13472, n20156);
  and g33264 (n20157, n_13471, n_13472);
  and g33265 (n20158, n_2802, n_13467);
  and g33266 (n20159, n_13468, n20158);
  not g33267 (n_13473, n20157);
  not g33268 (n_13474, n20159);
  and g33269 (n20160, n_13473, n_13474);
  not g33270 (n_13475, n20150);
  not g33271 (n_13476, n20160);
  and g33272 (n20161, n_13475, n_13476);
  not g33273 (n_13477, n20161);
  and g33274 (n20162, \asqrt[41] , n_13477);
  and g33278 (n20166, n_13011, n_13010);
  and g33279 (n20167, \asqrt[7] , n20166);
  not g33280 (n_13478, n20167);
  and g33281 (n20168, n_13009, n_13478);
  not g33282 (n_13479, n20165);
  not g33283 (n_13480, n20168);
  and g33284 (n20169, n_13479, n_13480);
  and g33285 (n20170, n_2594, n_13475);
  and g33286 (n20171, n_13476, n20170);
  not g33287 (n_13481, n20169);
  not g33288 (n_13482, n20171);
  and g33289 (n20172, n_13481, n_13482);
  not g33290 (n_13483, n20162);
  not g33291 (n_13484, n20172);
  and g33292 (n20173, n_13483, n_13484);
  not g33293 (n_13485, n20173);
  and g33294 (n20174, \asqrt[42] , n_13485);
  and g33298 (n20178, n_13019, n_13018);
  and g33299 (n20179, \asqrt[7] , n20178);
  not g33300 (n_13486, n20179);
  and g33301 (n20180, n_13017, n_13486);
  not g33302 (n_13487, n20177);
  not g33303 (n_13488, n20180);
  and g33304 (n20181, n_13487, n_13488);
  and g33305 (n20182, n_2394, n_13483);
  and g33306 (n20183, n_13484, n20182);
  not g33307 (n_13489, n20181);
  not g33308 (n_13490, n20183);
  and g33309 (n20184, n_13489, n_13490);
  not g33310 (n_13491, n20174);
  not g33311 (n_13492, n20184);
  and g33312 (n20185, n_13491, n_13492);
  not g33313 (n_13493, n20185);
  and g33314 (n20186, \asqrt[43] , n_13493);
  and g33318 (n20190, n_13027, n_13026);
  and g33319 (n20191, \asqrt[7] , n20190);
  not g33320 (n_13494, n20191);
  and g33321 (n20192, n_13025, n_13494);
  not g33322 (n_13495, n20189);
  not g33323 (n_13496, n20192);
  and g33324 (n20193, n_13495, n_13496);
  and g33325 (n20194, n_2202, n_13491);
  and g33326 (n20195, n_13492, n20194);
  not g33327 (n_13497, n20193);
  not g33328 (n_13498, n20195);
  and g33329 (n20196, n_13497, n_13498);
  not g33330 (n_13499, n20186);
  not g33331 (n_13500, n20196);
  and g33332 (n20197, n_13499, n_13500);
  not g33333 (n_13501, n20197);
  and g33334 (n20198, \asqrt[44] , n_13501);
  and g33338 (n20202, n_13035, n_13034);
  and g33339 (n20203, \asqrt[7] , n20202);
  not g33340 (n_13502, n20203);
  and g33341 (n20204, n_13033, n_13502);
  not g33342 (n_13503, n20201);
  not g33343 (n_13504, n20204);
  and g33344 (n20205, n_13503, n_13504);
  and g33345 (n20206, n_2018, n_13499);
  and g33346 (n20207, n_13500, n20206);
  not g33347 (n_13505, n20205);
  not g33348 (n_13506, n20207);
  and g33349 (n20208, n_13505, n_13506);
  not g33350 (n_13507, n20198);
  not g33351 (n_13508, n20208);
  and g33352 (n20209, n_13507, n_13508);
  not g33353 (n_13509, n20209);
  and g33354 (n20210, \asqrt[45] , n_13509);
  and g33358 (n20214, n_13043, n_13042);
  and g33359 (n20215, \asqrt[7] , n20214);
  not g33360 (n_13510, n20215);
  and g33361 (n20216, n_13041, n_13510);
  not g33362 (n_13511, n20213);
  not g33363 (n_13512, n20216);
  and g33364 (n20217, n_13511, n_13512);
  and g33365 (n20218, n_1842, n_13507);
  and g33366 (n20219, n_13508, n20218);
  not g33367 (n_13513, n20217);
  not g33368 (n_13514, n20219);
  and g33369 (n20220, n_13513, n_13514);
  not g33370 (n_13515, n20210);
  not g33371 (n_13516, n20220);
  and g33372 (n20221, n_13515, n_13516);
  not g33373 (n_13517, n20221);
  and g33374 (n20222, \asqrt[46] , n_13517);
  and g33378 (n20226, n_13051, n_13050);
  and g33379 (n20227, \asqrt[7] , n20226);
  not g33380 (n_13518, n20227);
  and g33381 (n20228, n_13049, n_13518);
  not g33382 (n_13519, n20225);
  not g33383 (n_13520, n20228);
  and g33384 (n20229, n_13519, n_13520);
  and g33385 (n20230, n_1674, n_13515);
  and g33386 (n20231, n_13516, n20230);
  not g33387 (n_13521, n20229);
  not g33388 (n_13522, n20231);
  and g33389 (n20232, n_13521, n_13522);
  not g33390 (n_13523, n20222);
  not g33391 (n_13524, n20232);
  and g33392 (n20233, n_13523, n_13524);
  not g33393 (n_13525, n20233);
  and g33394 (n20234, \asqrt[47] , n_13525);
  and g33398 (n20238, n_13059, n_13058);
  and g33399 (n20239, \asqrt[7] , n20238);
  not g33400 (n_13526, n20239);
  and g33401 (n20240, n_13057, n_13526);
  not g33402 (n_13527, n20237);
  not g33403 (n_13528, n20240);
  and g33404 (n20241, n_13527, n_13528);
  and g33405 (n20242, n_1514, n_13523);
  and g33406 (n20243, n_13524, n20242);
  not g33407 (n_13529, n20241);
  not g33408 (n_13530, n20243);
  and g33409 (n20244, n_13529, n_13530);
  not g33410 (n_13531, n20234);
  not g33411 (n_13532, n20244);
  and g33412 (n20245, n_13531, n_13532);
  not g33413 (n_13533, n20245);
  and g33414 (n20246, \asqrt[48] , n_13533);
  and g33418 (n20250, n_13067, n_13066);
  and g33419 (n20251, \asqrt[7] , n20250);
  not g33420 (n_13534, n20251);
  and g33421 (n20252, n_13065, n_13534);
  not g33422 (n_13535, n20249);
  not g33423 (n_13536, n20252);
  and g33424 (n20253, n_13535, n_13536);
  and g33425 (n20254, n_1362, n_13531);
  and g33426 (n20255, n_13532, n20254);
  not g33427 (n_13537, n20253);
  not g33428 (n_13538, n20255);
  and g33429 (n20256, n_13537, n_13538);
  not g33430 (n_13539, n20246);
  not g33431 (n_13540, n20256);
  and g33432 (n20257, n_13539, n_13540);
  not g33433 (n_13541, n20257);
  and g33434 (n20258, \asqrt[49] , n_13541);
  and g33438 (n20262, n_13075, n_13074);
  and g33439 (n20263, \asqrt[7] , n20262);
  not g33440 (n_13542, n20263);
  and g33441 (n20264, n_13073, n_13542);
  not g33442 (n_13543, n20261);
  not g33443 (n_13544, n20264);
  and g33444 (n20265, n_13543, n_13544);
  and g33445 (n20266, n_1218, n_13539);
  and g33446 (n20267, n_13540, n20266);
  not g33447 (n_13545, n20265);
  not g33448 (n_13546, n20267);
  and g33449 (n20268, n_13545, n_13546);
  not g33450 (n_13547, n20258);
  not g33451 (n_13548, n20268);
  and g33452 (n20269, n_13547, n_13548);
  not g33453 (n_13549, n20269);
  and g33454 (n20270, \asqrt[50] , n_13549);
  and g33458 (n20274, n_13083, n_13082);
  and g33459 (n20275, \asqrt[7] , n20274);
  not g33460 (n_13550, n20275);
  and g33461 (n20276, n_13081, n_13550);
  not g33462 (n_13551, n20273);
  not g33463 (n_13552, n20276);
  and g33464 (n20277, n_13551, n_13552);
  and g33465 (n20278, n_1082, n_13547);
  and g33466 (n20279, n_13548, n20278);
  not g33467 (n_13553, n20277);
  not g33468 (n_13554, n20279);
  and g33469 (n20280, n_13553, n_13554);
  not g33470 (n_13555, n20270);
  not g33471 (n_13556, n20280);
  and g33472 (n20281, n_13555, n_13556);
  not g33473 (n_13557, n20281);
  and g33474 (n20282, \asqrt[51] , n_13557);
  and g33478 (n20286, n_13091, n_13090);
  and g33479 (n20287, \asqrt[7] , n20286);
  not g33480 (n_13558, n20287);
  and g33481 (n20288, n_13089, n_13558);
  not g33482 (n_13559, n20285);
  not g33483 (n_13560, n20288);
  and g33484 (n20289, n_13559, n_13560);
  and g33485 (n20290, n_954, n_13555);
  and g33486 (n20291, n_13556, n20290);
  not g33487 (n_13561, n20289);
  not g33488 (n_13562, n20291);
  and g33489 (n20292, n_13561, n_13562);
  not g33490 (n_13563, n20282);
  not g33491 (n_13564, n20292);
  and g33492 (n20293, n_13563, n_13564);
  not g33493 (n_13565, n20293);
  and g33494 (n20294, \asqrt[52] , n_13565);
  and g33498 (n20298, n_13099, n_13098);
  and g33499 (n20299, \asqrt[7] , n20298);
  not g33500 (n_13566, n20299);
  and g33501 (n20300, n_13097, n_13566);
  not g33502 (n_13567, n20297);
  not g33503 (n_13568, n20300);
  and g33504 (n20301, n_13567, n_13568);
  and g33505 (n20302, n_834, n_13563);
  and g33506 (n20303, n_13564, n20302);
  not g33507 (n_13569, n20301);
  not g33508 (n_13570, n20303);
  and g33509 (n20304, n_13569, n_13570);
  not g33510 (n_13571, n20294);
  not g33511 (n_13572, n20304);
  and g33512 (n20305, n_13571, n_13572);
  not g33513 (n_13573, n20305);
  and g33514 (n20306, \asqrt[53] , n_13573);
  and g33518 (n20310, n_13107, n_13106);
  and g33519 (n20311, \asqrt[7] , n20310);
  not g33520 (n_13574, n20311);
  and g33521 (n20312, n_13105, n_13574);
  not g33522 (n_13575, n20309);
  not g33523 (n_13576, n20312);
  and g33524 (n20313, n_13575, n_13576);
  and g33525 (n20314, n_722, n_13571);
  and g33526 (n20315, n_13572, n20314);
  not g33527 (n_13577, n20313);
  not g33528 (n_13578, n20315);
  and g33529 (n20316, n_13577, n_13578);
  not g33530 (n_13579, n20306);
  not g33531 (n_13580, n20316);
  and g33532 (n20317, n_13579, n_13580);
  not g33533 (n_13581, n20317);
  and g33534 (n20318, \asqrt[54] , n_13581);
  and g33538 (n20322, n_13115, n_13114);
  and g33539 (n20323, \asqrt[7] , n20322);
  not g33540 (n_13582, n20323);
  and g33541 (n20324, n_13113, n_13582);
  not g33542 (n_13583, n20321);
  not g33543 (n_13584, n20324);
  and g33544 (n20325, n_13583, n_13584);
  and g33545 (n20326, n_618, n_13579);
  and g33546 (n20327, n_13580, n20326);
  not g33547 (n_13585, n20325);
  not g33548 (n_13586, n20327);
  and g33549 (n20328, n_13585, n_13586);
  not g33550 (n_13587, n20318);
  not g33551 (n_13588, n20328);
  and g33552 (n20329, n_13587, n_13588);
  not g33553 (n_13589, n20329);
  and g33554 (n20330, \asqrt[55] , n_13589);
  and g33558 (n20334, n_13123, n_13122);
  and g33559 (n20335, \asqrt[7] , n20334);
  not g33560 (n_13590, n20335);
  and g33561 (n20336, n_13121, n_13590);
  not g33562 (n_13591, n20333);
  not g33563 (n_13592, n20336);
  and g33564 (n20337, n_13591, n_13592);
  and g33565 (n20338, n_522, n_13587);
  and g33566 (n20339, n_13588, n20338);
  not g33567 (n_13593, n20337);
  not g33568 (n_13594, n20339);
  and g33569 (n20340, n_13593, n_13594);
  not g33570 (n_13595, n20330);
  not g33571 (n_13596, n20340);
  and g33572 (n20341, n_13595, n_13596);
  not g33573 (n_13597, n20341);
  and g33574 (n20342, \asqrt[56] , n_13597);
  and g33578 (n20346, n_13131, n_13130);
  and g33579 (n20347, \asqrt[7] , n20346);
  not g33580 (n_13598, n20347);
  and g33581 (n20348, n_13129, n_13598);
  not g33582 (n_13599, n20345);
  not g33583 (n_13600, n20348);
  and g33584 (n20349, n_13599, n_13600);
  and g33585 (n20350, n_434, n_13595);
  and g33586 (n20351, n_13596, n20350);
  not g33587 (n_13601, n20349);
  not g33588 (n_13602, n20351);
  and g33589 (n20352, n_13601, n_13602);
  not g33590 (n_13603, n20342);
  not g33591 (n_13604, n20352);
  and g33592 (n20353, n_13603, n_13604);
  not g33593 (n_13605, n20353);
  and g33594 (n20354, \asqrt[57] , n_13605);
  and g33598 (n20358, n_13139, n_13138);
  and g33599 (n20359, \asqrt[7] , n20358);
  not g33600 (n_13606, n20359);
  and g33601 (n20360, n_13137, n_13606);
  not g33602 (n_13607, n20357);
  not g33603 (n_13608, n20360);
  and g33604 (n20361, n_13607, n_13608);
  and g33605 (n20362, n_354, n_13603);
  and g33606 (n20363, n_13604, n20362);
  not g33607 (n_13609, n20361);
  not g33608 (n_13610, n20363);
  and g33609 (n20364, n_13609, n_13610);
  not g33610 (n_13611, n20354);
  not g33611 (n_13612, n20364);
  and g33612 (n20365, n_13611, n_13612);
  not g33613 (n_13613, n20365);
  and g33614 (n20366, \asqrt[58] , n_13613);
  and g33615 (n20367, n_282, n_13611);
  and g33616 (n20368, n_13612, n20367);
  and g33620 (n20372, n_13147, n_13145);
  and g33621 (n20373, \asqrt[7] , n20372);
  not g33622 (n_13614, n20373);
  and g33623 (n20374, n_13146, n_13614);
  not g33624 (n_13615, n20371);
  not g33625 (n_13616, n20374);
  and g33626 (n20375, n_13615, n_13616);
  not g33627 (n_13617, n20368);
  not g33628 (n_13618, n20375);
  and g33629 (n20376, n_13617, n_13618);
  not g33630 (n_13619, n20366);
  not g33631 (n_13620, n20376);
  and g33632 (n20377, n_13619, n_13620);
  not g33633 (n_13621, n20377);
  and g33634 (n20378, \asqrt[59] , n_13621);
  and g33638 (n20382, n_13155, n_13154);
  and g33639 (n20383, \asqrt[7] , n20382);
  not g33640 (n_13622, n20383);
  and g33641 (n20384, n_13153, n_13622);
  not g33642 (n_13623, n20381);
  not g33643 (n_13624, n20384);
  and g33644 (n20385, n_13623, n_13624);
  and g33645 (n20386, n_218, n_13619);
  and g33646 (n20387, n_13620, n20386);
  not g33647 (n_13625, n20385);
  not g33648 (n_13626, n20387);
  and g33649 (n20388, n_13625, n_13626);
  not g33650 (n_13627, n20378);
  not g33651 (n_13628, n20388);
  and g33652 (n20389, n_13627, n_13628);
  not g33653 (n_13629, n20389);
  and g33654 (n20390, \asqrt[60] , n_13629);
  and g33658 (n20394, n_13163, n_13162);
  and g33659 (n20395, \asqrt[7] , n20394);
  not g33660 (n_13630, n20395);
  and g33661 (n20396, n_13161, n_13630);
  not g33662 (n_13631, n20393);
  not g33663 (n_13632, n20396);
  and g33664 (n20397, n_13631, n_13632);
  and g33665 (n20398, n_162, n_13627);
  and g33666 (n20399, n_13628, n20398);
  not g33667 (n_13633, n20397);
  not g33668 (n_13634, n20399);
  and g33669 (n20400, n_13633, n_13634);
  not g33670 (n_13635, n20390);
  not g33671 (n_13636, n20400);
  and g33672 (n20401, n_13635, n_13636);
  not g33673 (n_13637, n20401);
  and g33674 (n20402, \asqrt[61] , n_13637);
  and g33678 (n20406, n_13171, n_13170);
  and g33679 (n20407, \asqrt[7] , n20406);
  not g33680 (n_13638, n20407);
  and g33681 (n20408, n_13169, n_13638);
  not g33682 (n_13639, n20405);
  not g33683 (n_13640, n20408);
  and g33684 (n20409, n_13639, n_13640);
  and g33685 (n20410, n_115, n_13635);
  and g33686 (n20411, n_13636, n20410);
  not g33687 (n_13641, n20409);
  not g33688 (n_13642, n20411);
  and g33689 (n20412, n_13641, n_13642);
  not g33690 (n_13643, n20402);
  not g33691 (n_13644, n20412);
  and g33692 (n20413, n_13643, n_13644);
  not g33693 (n_13645, n20413);
  and g33694 (n20414, \asqrt[62] , n_13645);
  and g33698 (n20418, n_13179, n_13178);
  and g33699 (n20419, \asqrt[7] , n20418);
  not g33700 (n_13646, n20419);
  and g33701 (n20420, n_13177, n_13646);
  not g33702 (n_13647, n20417);
  not g33703 (n_13648, n20420);
  and g33704 (n20421, n_13647, n_13648);
  and g33705 (n20422, n_76, n_13643);
  and g33706 (n20423, n_13644, n20422);
  not g33707 (n_13649, n20421);
  not g33708 (n_13650, n20423);
  and g33709 (n20424, n_13649, n_13650);
  not g33710 (n_13651, n20414);
  not g33711 (n_13652, n20424);
  and g33712 (n20425, n_13651, n_13652);
  and g33716 (n20429, n_13187, n_13186);
  and g33717 (n20430, \asqrt[7] , n20429);
  not g33718 (n_13653, n20430);
  and g33719 (n20431, n_13185, n_13653);
  not g33720 (n_13654, n20428);
  not g33721 (n_13655, n20431);
  and g33722 (n20432, n_13654, n_13655);
  and g33723 (n20433, n_13194, n_13193);
  and g33724 (n20434, \asqrt[7] , n20433);
  not g33727 (n_13657, n20432);
  not g33729 (n_13658, n20425);
  not g33731 (n_13659, n20437);
  and g33732 (n20438, n_21, n_13659);
  and g33733 (n20439, n_13651, n20432);
  and g33734 (n20440, n_13652, n20439);
  and g33735 (n20441, n_13193, \asqrt[7] );
  not g33736 (n_13660, n20441);
  and g33737 (n20442, n19733, n_13660);
  not g33738 (n_13661, n20433);
  and g33739 (n20443, \asqrt[63] , n_13661);
  not g33740 (n_13662, n20442);
  and g33741 (n20444, n_13662, n20443);
  not g33747 (n_13663, n20444);
  not g33748 (n_13664, n20449);
  not g33750 (n_13665, n20440);
  and g33754 (n20453, \a[12] , \asqrt[6] );
  not g33755 (n_13670, \a[10] );
  not g33756 (n_13671, \a[11] );
  and g33757 (n20454, n_13670, n_13671);
  and g33758 (n20455, n_13206, n20454);
  not g33759 (n_13672, n20453);
  not g33760 (n_13673, n20455);
  and g33761 (n20456, n_13672, n_13673);
  not g33762 (n_13674, n20456);
  and g33763 (n20457, \asqrt[7] , n_13674);
  and g33769 (n20463, n_13206, \asqrt[6] );
  not g33770 (n_13675, n20463);
  and g33771 (n20464, \a[13] , n_13675);
  and g33772 (n20465, n19762, \asqrt[6] );
  not g33773 (n_13676, n20464);
  not g33774 (n_13677, n20465);
  and g33775 (n20466, n_13676, n_13677);
  not g33776 (n_13678, n20462);
  and g33777 (n20467, n_13678, n20466);
  not g33778 (n_13679, n20457);
  not g33779 (n_13680, n20467);
  and g33780 (n20468, n_13679, n_13680);
  not g33781 (n_13681, n20468);
  and g33782 (n20469, \asqrt[8] , n_13681);
  not g33783 (n_13682, \asqrt[8] );
  and g33784 (n20470, n_13682, n_13679);
  and g33785 (n20471, n_13680, n20470);
  not g33789 (n_13683, n20438);
  not g33791 (n_13684, n20475);
  and g33792 (n20476, n_13677, n_13684);
  not g33793 (n_13685, n20476);
  and g33794 (n20477, \a[14] , n_13685);
  and g33795 (n20478, n_12750, n_13684);
  and g33796 (n20479, n_13677, n20478);
  not g33797 (n_13686, n20477);
  not g33798 (n_13687, n20479);
  and g33799 (n20480, n_13686, n_13687);
  not g33800 (n_13688, n20471);
  not g33801 (n_13689, n20480);
  and g33802 (n20481, n_13688, n_13689);
  not g33803 (n_13690, n20469);
  not g33804 (n_13691, n20481);
  and g33805 (n20482, n_13690, n_13691);
  not g33806 (n_13692, n20482);
  and g33807 (n20483, \asqrt[9] , n_13692);
  and g33808 (n20484, n_13215, n_13214);
  not g33809 (n_13693, n19774);
  and g33810 (n20485, n_13693, n20484);
  and g33811 (n20486, \asqrt[6] , n20485);
  and g33812 (n20487, \asqrt[6] , n20484);
  not g33813 (n_13694, n20487);
  and g33814 (n20488, n19774, n_13694);
  not g33815 (n_13695, n20486);
  not g33816 (n_13696, n20488);
  and g33817 (n20489, n_13695, n_13696);
  and g33818 (n20490, n_13218, n_13690);
  and g33819 (n20491, n_13691, n20490);
  not g33820 (n_13697, n20489);
  not g33821 (n_13698, n20491);
  and g33822 (n20492, n_13697, n_13698);
  not g33823 (n_13699, n20483);
  not g33824 (n_13700, n20492);
  and g33825 (n20493, n_13699, n_13700);
  not g33826 (n_13701, n20493);
  and g33827 (n20494, \asqrt[10] , n_13701);
  and g33831 (n20498, n_13226, n_13224);
  and g33832 (n20499, \asqrt[6] , n20498);
  not g33833 (n_13702, n20499);
  and g33834 (n20500, n_13225, n_13702);
  not g33835 (n_13703, n20497);
  not g33836 (n_13704, n20500);
  and g33837 (n20501, n_13703, n_13704);
  and g33838 (n20502, n_12762, n_13699);
  and g33839 (n20503, n_13700, n20502);
  not g33840 (n_13705, n20501);
  not g33841 (n_13706, n20503);
  and g33842 (n20504, n_13705, n_13706);
  not g33843 (n_13707, n20494);
  not g33844 (n_13708, n20504);
  and g33845 (n20505, n_13707, n_13708);
  not g33846 (n_13709, n20505);
  and g33847 (n20506, \asqrt[11] , n_13709);
  and g33851 (n20510, n_13235, n_13234);
  and g33852 (n20511, \asqrt[6] , n20510);
  not g33853 (n_13710, n20511);
  and g33854 (n20512, n_13233, n_13710);
  not g33855 (n_13711, n20509);
  not g33856 (n_13712, n20512);
  and g33857 (n20513, n_13711, n_13712);
  and g33858 (n20514, n_12314, n_13707);
  and g33859 (n20515, n_13708, n20514);
  not g33860 (n_13713, n20513);
  not g33861 (n_13714, n20515);
  and g33862 (n20516, n_13713, n_13714);
  not g33863 (n_13715, n20506);
  not g33864 (n_13716, n20516);
  and g33865 (n20517, n_13715, n_13716);
  not g33866 (n_13717, n20517);
  and g33867 (n20518, \asqrt[12] , n_13717);
  and g33871 (n20522, n_13243, n_13242);
  and g33872 (n20523, \asqrt[6] , n20522);
  not g33873 (n_13718, n20523);
  and g33874 (n20524, n_13241, n_13718);
  not g33875 (n_13719, n20521);
  not g33876 (n_13720, n20524);
  and g33877 (n20525, n_13719, n_13720);
  and g33878 (n20526, n_11874, n_13715);
  and g33879 (n20527, n_13716, n20526);
  not g33880 (n_13721, n20525);
  not g33881 (n_13722, n20527);
  and g33882 (n20528, n_13721, n_13722);
  not g33883 (n_13723, n20518);
  not g33884 (n_13724, n20528);
  and g33885 (n20529, n_13723, n_13724);
  not g33886 (n_13725, n20529);
  and g33887 (n20530, \asqrt[13] , n_13725);
  and g33891 (n20534, n_13251, n_13250);
  and g33892 (n20535, \asqrt[6] , n20534);
  not g33893 (n_13726, n20535);
  and g33894 (n20536, n_13249, n_13726);
  not g33895 (n_13727, n20533);
  not g33896 (n_13728, n20536);
  and g33897 (n20537, n_13727, n_13728);
  and g33898 (n20538, n_11442, n_13723);
  and g33899 (n20539, n_13724, n20538);
  not g33900 (n_13729, n20537);
  not g33901 (n_13730, n20539);
  and g33902 (n20540, n_13729, n_13730);
  not g33903 (n_13731, n20530);
  not g33904 (n_13732, n20540);
  and g33905 (n20541, n_13731, n_13732);
  not g33906 (n_13733, n20541);
  and g33907 (n20542, \asqrt[14] , n_13733);
  and g33911 (n20546, n_13259, n_13258);
  and g33912 (n20547, \asqrt[6] , n20546);
  not g33913 (n_13734, n20547);
  and g33914 (n20548, n_13257, n_13734);
  not g33915 (n_13735, n20545);
  not g33916 (n_13736, n20548);
  and g33917 (n20549, n_13735, n_13736);
  and g33918 (n20550, n_11018, n_13731);
  and g33919 (n20551, n_13732, n20550);
  not g33920 (n_13737, n20549);
  not g33921 (n_13738, n20551);
  and g33922 (n20552, n_13737, n_13738);
  not g33923 (n_13739, n20542);
  not g33924 (n_13740, n20552);
  and g33925 (n20553, n_13739, n_13740);
  not g33926 (n_13741, n20553);
  and g33927 (n20554, \asqrt[15] , n_13741);
  and g33931 (n20558, n_13267, n_13266);
  and g33932 (n20559, \asqrt[6] , n20558);
  not g33933 (n_13742, n20559);
  and g33934 (n20560, n_13265, n_13742);
  not g33935 (n_13743, n20557);
  not g33936 (n_13744, n20560);
  and g33937 (n20561, n_13743, n_13744);
  and g33938 (n20562, n_10602, n_13739);
  and g33939 (n20563, n_13740, n20562);
  not g33940 (n_13745, n20561);
  not g33941 (n_13746, n20563);
  and g33942 (n20564, n_13745, n_13746);
  not g33943 (n_13747, n20554);
  not g33944 (n_13748, n20564);
  and g33945 (n20565, n_13747, n_13748);
  not g33946 (n_13749, n20565);
  and g33947 (n20566, \asqrt[16] , n_13749);
  and g33951 (n20570, n_13275, n_13274);
  and g33952 (n20571, \asqrt[6] , n20570);
  not g33953 (n_13750, n20571);
  and g33954 (n20572, n_13273, n_13750);
  not g33955 (n_13751, n20569);
  not g33956 (n_13752, n20572);
  and g33957 (n20573, n_13751, n_13752);
  and g33958 (n20574, n_10194, n_13747);
  and g33959 (n20575, n_13748, n20574);
  not g33960 (n_13753, n20573);
  not g33961 (n_13754, n20575);
  and g33962 (n20576, n_13753, n_13754);
  not g33963 (n_13755, n20566);
  not g33964 (n_13756, n20576);
  and g33965 (n20577, n_13755, n_13756);
  not g33966 (n_13757, n20577);
  and g33967 (n20578, \asqrt[17] , n_13757);
  and g33971 (n20582, n_13283, n_13282);
  and g33972 (n20583, \asqrt[6] , n20582);
  not g33973 (n_13758, n20583);
  and g33974 (n20584, n_13281, n_13758);
  not g33975 (n_13759, n20581);
  not g33976 (n_13760, n20584);
  and g33977 (n20585, n_13759, n_13760);
  and g33978 (n20586, n_9794, n_13755);
  and g33979 (n20587, n_13756, n20586);
  not g33980 (n_13761, n20585);
  not g33981 (n_13762, n20587);
  and g33982 (n20588, n_13761, n_13762);
  not g33983 (n_13763, n20578);
  not g33984 (n_13764, n20588);
  and g33985 (n20589, n_13763, n_13764);
  not g33986 (n_13765, n20589);
  and g33987 (n20590, \asqrt[18] , n_13765);
  and g33991 (n20594, n_13291, n_13290);
  and g33992 (n20595, \asqrt[6] , n20594);
  not g33993 (n_13766, n20595);
  and g33994 (n20596, n_13289, n_13766);
  not g33995 (n_13767, n20593);
  not g33996 (n_13768, n20596);
  and g33997 (n20597, n_13767, n_13768);
  and g33998 (n20598, n_9402, n_13763);
  and g33999 (n20599, n_13764, n20598);
  not g34000 (n_13769, n20597);
  not g34001 (n_13770, n20599);
  and g34002 (n20600, n_13769, n_13770);
  not g34003 (n_13771, n20590);
  not g34004 (n_13772, n20600);
  and g34005 (n20601, n_13771, n_13772);
  not g34006 (n_13773, n20601);
  and g34007 (n20602, \asqrt[19] , n_13773);
  and g34011 (n20606, n_13299, n_13298);
  and g34012 (n20607, \asqrt[6] , n20606);
  not g34013 (n_13774, n20607);
  and g34014 (n20608, n_13297, n_13774);
  not g34015 (n_13775, n20605);
  not g34016 (n_13776, n20608);
  and g34017 (n20609, n_13775, n_13776);
  and g34018 (n20610, n_9018, n_13771);
  and g34019 (n20611, n_13772, n20610);
  not g34020 (n_13777, n20609);
  not g34021 (n_13778, n20611);
  and g34022 (n20612, n_13777, n_13778);
  not g34023 (n_13779, n20602);
  not g34024 (n_13780, n20612);
  and g34025 (n20613, n_13779, n_13780);
  not g34026 (n_13781, n20613);
  and g34027 (n20614, \asqrt[20] , n_13781);
  and g34031 (n20618, n_13307, n_13306);
  and g34032 (n20619, \asqrt[6] , n20618);
  not g34033 (n_13782, n20619);
  and g34034 (n20620, n_13305, n_13782);
  not g34035 (n_13783, n20617);
  not g34036 (n_13784, n20620);
  and g34037 (n20621, n_13783, n_13784);
  and g34038 (n20622, n_8642, n_13779);
  and g34039 (n20623, n_13780, n20622);
  not g34040 (n_13785, n20621);
  not g34041 (n_13786, n20623);
  and g34042 (n20624, n_13785, n_13786);
  not g34043 (n_13787, n20614);
  not g34044 (n_13788, n20624);
  and g34045 (n20625, n_13787, n_13788);
  not g34046 (n_13789, n20625);
  and g34047 (n20626, \asqrt[21] , n_13789);
  and g34051 (n20630, n_13315, n_13314);
  and g34052 (n20631, \asqrt[6] , n20630);
  not g34053 (n_13790, n20631);
  and g34054 (n20632, n_13313, n_13790);
  not g34055 (n_13791, n20629);
  not g34056 (n_13792, n20632);
  and g34057 (n20633, n_13791, n_13792);
  and g34058 (n20634, n_8274, n_13787);
  and g34059 (n20635, n_13788, n20634);
  not g34060 (n_13793, n20633);
  not g34061 (n_13794, n20635);
  and g34062 (n20636, n_13793, n_13794);
  not g34063 (n_13795, n20626);
  not g34064 (n_13796, n20636);
  and g34065 (n20637, n_13795, n_13796);
  not g34066 (n_13797, n20637);
  and g34067 (n20638, \asqrt[22] , n_13797);
  and g34071 (n20642, n_13323, n_13322);
  and g34072 (n20643, \asqrt[6] , n20642);
  not g34073 (n_13798, n20643);
  and g34074 (n20644, n_13321, n_13798);
  not g34075 (n_13799, n20641);
  not g34076 (n_13800, n20644);
  and g34077 (n20645, n_13799, n_13800);
  and g34078 (n20646, n_7914, n_13795);
  and g34079 (n20647, n_13796, n20646);
  not g34080 (n_13801, n20645);
  not g34081 (n_13802, n20647);
  and g34082 (n20648, n_13801, n_13802);
  not g34083 (n_13803, n20638);
  not g34084 (n_13804, n20648);
  and g34085 (n20649, n_13803, n_13804);
  not g34086 (n_13805, n20649);
  and g34087 (n20650, \asqrt[23] , n_13805);
  and g34091 (n20654, n_13331, n_13330);
  and g34092 (n20655, \asqrt[6] , n20654);
  not g34093 (n_13806, n20655);
  and g34094 (n20656, n_13329, n_13806);
  not g34095 (n_13807, n20653);
  not g34096 (n_13808, n20656);
  and g34097 (n20657, n_13807, n_13808);
  and g34098 (n20658, n_7562, n_13803);
  and g34099 (n20659, n_13804, n20658);
  not g34100 (n_13809, n20657);
  not g34101 (n_13810, n20659);
  and g34102 (n20660, n_13809, n_13810);
  not g34103 (n_13811, n20650);
  not g34104 (n_13812, n20660);
  and g34105 (n20661, n_13811, n_13812);
  not g34106 (n_13813, n20661);
  and g34107 (n20662, \asqrt[24] , n_13813);
  and g34111 (n20666, n_13339, n_13338);
  and g34112 (n20667, \asqrt[6] , n20666);
  not g34113 (n_13814, n20667);
  and g34114 (n20668, n_13337, n_13814);
  not g34115 (n_13815, n20665);
  not g34116 (n_13816, n20668);
  and g34117 (n20669, n_13815, n_13816);
  and g34118 (n20670, n_7218, n_13811);
  and g34119 (n20671, n_13812, n20670);
  not g34120 (n_13817, n20669);
  not g34121 (n_13818, n20671);
  and g34122 (n20672, n_13817, n_13818);
  not g34123 (n_13819, n20662);
  not g34124 (n_13820, n20672);
  and g34125 (n20673, n_13819, n_13820);
  not g34126 (n_13821, n20673);
  and g34127 (n20674, \asqrt[25] , n_13821);
  and g34131 (n20678, n_13347, n_13346);
  and g34132 (n20679, \asqrt[6] , n20678);
  not g34133 (n_13822, n20679);
  and g34134 (n20680, n_13345, n_13822);
  not g34135 (n_13823, n20677);
  not g34136 (n_13824, n20680);
  and g34137 (n20681, n_13823, n_13824);
  and g34138 (n20682, n_6882, n_13819);
  and g34139 (n20683, n_13820, n20682);
  not g34140 (n_13825, n20681);
  not g34141 (n_13826, n20683);
  and g34142 (n20684, n_13825, n_13826);
  not g34143 (n_13827, n20674);
  not g34144 (n_13828, n20684);
  and g34145 (n20685, n_13827, n_13828);
  not g34146 (n_13829, n20685);
  and g34147 (n20686, \asqrt[26] , n_13829);
  and g34151 (n20690, n_13355, n_13354);
  and g34152 (n20691, \asqrt[6] , n20690);
  not g34153 (n_13830, n20691);
  and g34154 (n20692, n_13353, n_13830);
  not g34155 (n_13831, n20689);
  not g34156 (n_13832, n20692);
  and g34157 (n20693, n_13831, n_13832);
  and g34158 (n20694, n_6554, n_13827);
  and g34159 (n20695, n_13828, n20694);
  not g34160 (n_13833, n20693);
  not g34161 (n_13834, n20695);
  and g34162 (n20696, n_13833, n_13834);
  not g34163 (n_13835, n20686);
  not g34164 (n_13836, n20696);
  and g34165 (n20697, n_13835, n_13836);
  not g34166 (n_13837, n20697);
  and g34167 (n20698, \asqrt[27] , n_13837);
  and g34171 (n20702, n_13363, n_13362);
  and g34172 (n20703, \asqrt[6] , n20702);
  not g34173 (n_13838, n20703);
  and g34174 (n20704, n_13361, n_13838);
  not g34175 (n_13839, n20701);
  not g34176 (n_13840, n20704);
  and g34177 (n20705, n_13839, n_13840);
  and g34178 (n20706, n_6234, n_13835);
  and g34179 (n20707, n_13836, n20706);
  not g34180 (n_13841, n20705);
  not g34181 (n_13842, n20707);
  and g34182 (n20708, n_13841, n_13842);
  not g34183 (n_13843, n20698);
  not g34184 (n_13844, n20708);
  and g34185 (n20709, n_13843, n_13844);
  not g34186 (n_13845, n20709);
  and g34187 (n20710, \asqrt[28] , n_13845);
  and g34191 (n20714, n_13371, n_13370);
  and g34192 (n20715, \asqrt[6] , n20714);
  not g34193 (n_13846, n20715);
  and g34194 (n20716, n_13369, n_13846);
  not g34195 (n_13847, n20713);
  not g34196 (n_13848, n20716);
  and g34197 (n20717, n_13847, n_13848);
  and g34198 (n20718, n_5922, n_13843);
  and g34199 (n20719, n_13844, n20718);
  not g34200 (n_13849, n20717);
  not g34201 (n_13850, n20719);
  and g34202 (n20720, n_13849, n_13850);
  not g34203 (n_13851, n20710);
  not g34204 (n_13852, n20720);
  and g34205 (n20721, n_13851, n_13852);
  not g34206 (n_13853, n20721);
  and g34207 (n20722, \asqrt[29] , n_13853);
  and g34211 (n20726, n_13379, n_13378);
  and g34212 (n20727, \asqrt[6] , n20726);
  not g34213 (n_13854, n20727);
  and g34214 (n20728, n_13377, n_13854);
  not g34215 (n_13855, n20725);
  not g34216 (n_13856, n20728);
  and g34217 (n20729, n_13855, n_13856);
  and g34218 (n20730, n_5618, n_13851);
  and g34219 (n20731, n_13852, n20730);
  not g34220 (n_13857, n20729);
  not g34221 (n_13858, n20731);
  and g34222 (n20732, n_13857, n_13858);
  not g34223 (n_13859, n20722);
  not g34224 (n_13860, n20732);
  and g34225 (n20733, n_13859, n_13860);
  not g34226 (n_13861, n20733);
  and g34227 (n20734, \asqrt[30] , n_13861);
  and g34231 (n20738, n_13387, n_13386);
  and g34232 (n20739, \asqrt[6] , n20738);
  not g34233 (n_13862, n20739);
  and g34234 (n20740, n_13385, n_13862);
  not g34235 (n_13863, n20737);
  not g34236 (n_13864, n20740);
  and g34237 (n20741, n_13863, n_13864);
  and g34238 (n20742, n_5322, n_13859);
  and g34239 (n20743, n_13860, n20742);
  not g34240 (n_13865, n20741);
  not g34241 (n_13866, n20743);
  and g34242 (n20744, n_13865, n_13866);
  not g34243 (n_13867, n20734);
  not g34244 (n_13868, n20744);
  and g34245 (n20745, n_13867, n_13868);
  not g34246 (n_13869, n20745);
  and g34247 (n20746, \asqrt[31] , n_13869);
  and g34251 (n20750, n_13395, n_13394);
  and g34252 (n20751, \asqrt[6] , n20750);
  not g34253 (n_13870, n20751);
  and g34254 (n20752, n_13393, n_13870);
  not g34255 (n_13871, n20749);
  not g34256 (n_13872, n20752);
  and g34257 (n20753, n_13871, n_13872);
  and g34258 (n20754, n_5034, n_13867);
  and g34259 (n20755, n_13868, n20754);
  not g34260 (n_13873, n20753);
  not g34261 (n_13874, n20755);
  and g34262 (n20756, n_13873, n_13874);
  not g34263 (n_13875, n20746);
  not g34264 (n_13876, n20756);
  and g34265 (n20757, n_13875, n_13876);
  not g34266 (n_13877, n20757);
  and g34267 (n20758, \asqrt[32] , n_13877);
  and g34271 (n20762, n_13403, n_13402);
  and g34272 (n20763, \asqrt[6] , n20762);
  not g34273 (n_13878, n20763);
  and g34274 (n20764, n_13401, n_13878);
  not g34275 (n_13879, n20761);
  not g34276 (n_13880, n20764);
  and g34277 (n20765, n_13879, n_13880);
  and g34278 (n20766, n_4754, n_13875);
  and g34279 (n20767, n_13876, n20766);
  not g34280 (n_13881, n20765);
  not g34281 (n_13882, n20767);
  and g34282 (n20768, n_13881, n_13882);
  not g34283 (n_13883, n20758);
  not g34284 (n_13884, n20768);
  and g34285 (n20769, n_13883, n_13884);
  not g34286 (n_13885, n20769);
  and g34287 (n20770, \asqrt[33] , n_13885);
  and g34291 (n20774, n_13411, n_13410);
  and g34292 (n20775, \asqrt[6] , n20774);
  not g34293 (n_13886, n20775);
  and g34294 (n20776, n_13409, n_13886);
  not g34295 (n_13887, n20773);
  not g34296 (n_13888, n20776);
  and g34297 (n20777, n_13887, n_13888);
  and g34298 (n20778, n_4482, n_13883);
  and g34299 (n20779, n_13884, n20778);
  not g34300 (n_13889, n20777);
  not g34301 (n_13890, n20779);
  and g34302 (n20780, n_13889, n_13890);
  not g34303 (n_13891, n20770);
  not g34304 (n_13892, n20780);
  and g34305 (n20781, n_13891, n_13892);
  not g34306 (n_13893, n20781);
  and g34307 (n20782, \asqrt[34] , n_13893);
  and g34311 (n20786, n_13419, n_13418);
  and g34312 (n20787, \asqrt[6] , n20786);
  not g34313 (n_13894, n20787);
  and g34314 (n20788, n_13417, n_13894);
  not g34315 (n_13895, n20785);
  not g34316 (n_13896, n20788);
  and g34317 (n20789, n_13895, n_13896);
  and g34318 (n20790, n_4218, n_13891);
  and g34319 (n20791, n_13892, n20790);
  not g34320 (n_13897, n20789);
  not g34321 (n_13898, n20791);
  and g34322 (n20792, n_13897, n_13898);
  not g34323 (n_13899, n20782);
  not g34324 (n_13900, n20792);
  and g34325 (n20793, n_13899, n_13900);
  not g34326 (n_13901, n20793);
  and g34327 (n20794, \asqrt[35] , n_13901);
  and g34331 (n20798, n_13427, n_13426);
  and g34332 (n20799, \asqrt[6] , n20798);
  not g34333 (n_13902, n20799);
  and g34334 (n20800, n_13425, n_13902);
  not g34335 (n_13903, n20797);
  not g34336 (n_13904, n20800);
  and g34337 (n20801, n_13903, n_13904);
  and g34338 (n20802, n_3962, n_13899);
  and g34339 (n20803, n_13900, n20802);
  not g34340 (n_13905, n20801);
  not g34341 (n_13906, n20803);
  and g34342 (n20804, n_13905, n_13906);
  not g34343 (n_13907, n20794);
  not g34344 (n_13908, n20804);
  and g34345 (n20805, n_13907, n_13908);
  not g34346 (n_13909, n20805);
  and g34347 (n20806, \asqrt[36] , n_13909);
  and g34351 (n20810, n_13435, n_13434);
  and g34352 (n20811, \asqrt[6] , n20810);
  not g34353 (n_13910, n20811);
  and g34354 (n20812, n_13433, n_13910);
  not g34355 (n_13911, n20809);
  not g34356 (n_13912, n20812);
  and g34357 (n20813, n_13911, n_13912);
  and g34358 (n20814, n_3714, n_13907);
  and g34359 (n20815, n_13908, n20814);
  not g34360 (n_13913, n20813);
  not g34361 (n_13914, n20815);
  and g34362 (n20816, n_13913, n_13914);
  not g34363 (n_13915, n20806);
  not g34364 (n_13916, n20816);
  and g34365 (n20817, n_13915, n_13916);
  not g34366 (n_13917, n20817);
  and g34367 (n20818, \asqrt[37] , n_13917);
  and g34371 (n20822, n_13443, n_13442);
  and g34372 (n20823, \asqrt[6] , n20822);
  not g34373 (n_13918, n20823);
  and g34374 (n20824, n_13441, n_13918);
  not g34375 (n_13919, n20821);
  not g34376 (n_13920, n20824);
  and g34377 (n20825, n_13919, n_13920);
  and g34378 (n20826, n_3474, n_13915);
  and g34379 (n20827, n_13916, n20826);
  not g34380 (n_13921, n20825);
  not g34381 (n_13922, n20827);
  and g34382 (n20828, n_13921, n_13922);
  not g34383 (n_13923, n20818);
  not g34384 (n_13924, n20828);
  and g34385 (n20829, n_13923, n_13924);
  not g34386 (n_13925, n20829);
  and g34387 (n20830, \asqrt[38] , n_13925);
  and g34391 (n20834, n_13451, n_13450);
  and g34392 (n20835, \asqrt[6] , n20834);
  not g34393 (n_13926, n20835);
  and g34394 (n20836, n_13449, n_13926);
  not g34395 (n_13927, n20833);
  not g34396 (n_13928, n20836);
  and g34397 (n20837, n_13927, n_13928);
  and g34398 (n20838, n_3242, n_13923);
  and g34399 (n20839, n_13924, n20838);
  not g34400 (n_13929, n20837);
  not g34401 (n_13930, n20839);
  and g34402 (n20840, n_13929, n_13930);
  not g34403 (n_13931, n20830);
  not g34404 (n_13932, n20840);
  and g34405 (n20841, n_13931, n_13932);
  not g34406 (n_13933, n20841);
  and g34407 (n20842, \asqrt[39] , n_13933);
  and g34411 (n20846, n_13459, n_13458);
  and g34412 (n20847, \asqrt[6] , n20846);
  not g34413 (n_13934, n20847);
  and g34414 (n20848, n_13457, n_13934);
  not g34415 (n_13935, n20845);
  not g34416 (n_13936, n20848);
  and g34417 (n20849, n_13935, n_13936);
  and g34418 (n20850, n_3018, n_13931);
  and g34419 (n20851, n_13932, n20850);
  not g34420 (n_13937, n20849);
  not g34421 (n_13938, n20851);
  and g34422 (n20852, n_13937, n_13938);
  not g34423 (n_13939, n20842);
  not g34424 (n_13940, n20852);
  and g34425 (n20853, n_13939, n_13940);
  not g34426 (n_13941, n20853);
  and g34427 (n20854, \asqrt[40] , n_13941);
  and g34431 (n20858, n_13467, n_13466);
  and g34432 (n20859, \asqrt[6] , n20858);
  not g34433 (n_13942, n20859);
  and g34434 (n20860, n_13465, n_13942);
  not g34435 (n_13943, n20857);
  not g34436 (n_13944, n20860);
  and g34437 (n20861, n_13943, n_13944);
  and g34438 (n20862, n_2802, n_13939);
  and g34439 (n20863, n_13940, n20862);
  not g34440 (n_13945, n20861);
  not g34441 (n_13946, n20863);
  and g34442 (n20864, n_13945, n_13946);
  not g34443 (n_13947, n20854);
  not g34444 (n_13948, n20864);
  and g34445 (n20865, n_13947, n_13948);
  not g34446 (n_13949, n20865);
  and g34447 (n20866, \asqrt[41] , n_13949);
  and g34451 (n20870, n_13475, n_13474);
  and g34452 (n20871, \asqrt[6] , n20870);
  not g34453 (n_13950, n20871);
  and g34454 (n20872, n_13473, n_13950);
  not g34455 (n_13951, n20869);
  not g34456 (n_13952, n20872);
  and g34457 (n20873, n_13951, n_13952);
  and g34458 (n20874, n_2594, n_13947);
  and g34459 (n20875, n_13948, n20874);
  not g34460 (n_13953, n20873);
  not g34461 (n_13954, n20875);
  and g34462 (n20876, n_13953, n_13954);
  not g34463 (n_13955, n20866);
  not g34464 (n_13956, n20876);
  and g34465 (n20877, n_13955, n_13956);
  not g34466 (n_13957, n20877);
  and g34467 (n20878, \asqrt[42] , n_13957);
  and g34471 (n20882, n_13483, n_13482);
  and g34472 (n20883, \asqrt[6] , n20882);
  not g34473 (n_13958, n20883);
  and g34474 (n20884, n_13481, n_13958);
  not g34475 (n_13959, n20881);
  not g34476 (n_13960, n20884);
  and g34477 (n20885, n_13959, n_13960);
  and g34478 (n20886, n_2394, n_13955);
  and g34479 (n20887, n_13956, n20886);
  not g34480 (n_13961, n20885);
  not g34481 (n_13962, n20887);
  and g34482 (n20888, n_13961, n_13962);
  not g34483 (n_13963, n20878);
  not g34484 (n_13964, n20888);
  and g34485 (n20889, n_13963, n_13964);
  not g34486 (n_13965, n20889);
  and g34487 (n20890, \asqrt[43] , n_13965);
  and g34491 (n20894, n_13491, n_13490);
  and g34492 (n20895, \asqrt[6] , n20894);
  not g34493 (n_13966, n20895);
  and g34494 (n20896, n_13489, n_13966);
  not g34495 (n_13967, n20893);
  not g34496 (n_13968, n20896);
  and g34497 (n20897, n_13967, n_13968);
  and g34498 (n20898, n_2202, n_13963);
  and g34499 (n20899, n_13964, n20898);
  not g34500 (n_13969, n20897);
  not g34501 (n_13970, n20899);
  and g34502 (n20900, n_13969, n_13970);
  not g34503 (n_13971, n20890);
  not g34504 (n_13972, n20900);
  and g34505 (n20901, n_13971, n_13972);
  not g34506 (n_13973, n20901);
  and g34507 (n20902, \asqrt[44] , n_13973);
  and g34511 (n20906, n_13499, n_13498);
  and g34512 (n20907, \asqrt[6] , n20906);
  not g34513 (n_13974, n20907);
  and g34514 (n20908, n_13497, n_13974);
  not g34515 (n_13975, n20905);
  not g34516 (n_13976, n20908);
  and g34517 (n20909, n_13975, n_13976);
  and g34518 (n20910, n_2018, n_13971);
  and g34519 (n20911, n_13972, n20910);
  not g34520 (n_13977, n20909);
  not g34521 (n_13978, n20911);
  and g34522 (n20912, n_13977, n_13978);
  not g34523 (n_13979, n20902);
  not g34524 (n_13980, n20912);
  and g34525 (n20913, n_13979, n_13980);
  not g34526 (n_13981, n20913);
  and g34527 (n20914, \asqrt[45] , n_13981);
  and g34531 (n20918, n_13507, n_13506);
  and g34532 (n20919, \asqrt[6] , n20918);
  not g34533 (n_13982, n20919);
  and g34534 (n20920, n_13505, n_13982);
  not g34535 (n_13983, n20917);
  not g34536 (n_13984, n20920);
  and g34537 (n20921, n_13983, n_13984);
  and g34538 (n20922, n_1842, n_13979);
  and g34539 (n20923, n_13980, n20922);
  not g34540 (n_13985, n20921);
  not g34541 (n_13986, n20923);
  and g34542 (n20924, n_13985, n_13986);
  not g34543 (n_13987, n20914);
  not g34544 (n_13988, n20924);
  and g34545 (n20925, n_13987, n_13988);
  not g34546 (n_13989, n20925);
  and g34547 (n20926, \asqrt[46] , n_13989);
  and g34551 (n20930, n_13515, n_13514);
  and g34552 (n20931, \asqrt[6] , n20930);
  not g34553 (n_13990, n20931);
  and g34554 (n20932, n_13513, n_13990);
  not g34555 (n_13991, n20929);
  not g34556 (n_13992, n20932);
  and g34557 (n20933, n_13991, n_13992);
  and g34558 (n20934, n_1674, n_13987);
  and g34559 (n20935, n_13988, n20934);
  not g34560 (n_13993, n20933);
  not g34561 (n_13994, n20935);
  and g34562 (n20936, n_13993, n_13994);
  not g34563 (n_13995, n20926);
  not g34564 (n_13996, n20936);
  and g34565 (n20937, n_13995, n_13996);
  not g34566 (n_13997, n20937);
  and g34567 (n20938, \asqrt[47] , n_13997);
  and g34571 (n20942, n_13523, n_13522);
  and g34572 (n20943, \asqrt[6] , n20942);
  not g34573 (n_13998, n20943);
  and g34574 (n20944, n_13521, n_13998);
  not g34575 (n_13999, n20941);
  not g34576 (n_14000, n20944);
  and g34577 (n20945, n_13999, n_14000);
  and g34578 (n20946, n_1514, n_13995);
  and g34579 (n20947, n_13996, n20946);
  not g34580 (n_14001, n20945);
  not g34581 (n_14002, n20947);
  and g34582 (n20948, n_14001, n_14002);
  not g34583 (n_14003, n20938);
  not g34584 (n_14004, n20948);
  and g34585 (n20949, n_14003, n_14004);
  not g34586 (n_14005, n20949);
  and g34587 (n20950, \asqrt[48] , n_14005);
  and g34591 (n20954, n_13531, n_13530);
  and g34592 (n20955, \asqrt[6] , n20954);
  not g34593 (n_14006, n20955);
  and g34594 (n20956, n_13529, n_14006);
  not g34595 (n_14007, n20953);
  not g34596 (n_14008, n20956);
  and g34597 (n20957, n_14007, n_14008);
  and g34598 (n20958, n_1362, n_14003);
  and g34599 (n20959, n_14004, n20958);
  not g34600 (n_14009, n20957);
  not g34601 (n_14010, n20959);
  and g34602 (n20960, n_14009, n_14010);
  not g34603 (n_14011, n20950);
  not g34604 (n_14012, n20960);
  and g34605 (n20961, n_14011, n_14012);
  not g34606 (n_14013, n20961);
  and g34607 (n20962, \asqrt[49] , n_14013);
  and g34611 (n20966, n_13539, n_13538);
  and g34612 (n20967, \asqrt[6] , n20966);
  not g34613 (n_14014, n20967);
  and g34614 (n20968, n_13537, n_14014);
  not g34615 (n_14015, n20965);
  not g34616 (n_14016, n20968);
  and g34617 (n20969, n_14015, n_14016);
  and g34618 (n20970, n_1218, n_14011);
  and g34619 (n20971, n_14012, n20970);
  not g34620 (n_14017, n20969);
  not g34621 (n_14018, n20971);
  and g34622 (n20972, n_14017, n_14018);
  not g34623 (n_14019, n20962);
  not g34624 (n_14020, n20972);
  and g34625 (n20973, n_14019, n_14020);
  not g34626 (n_14021, n20973);
  and g34627 (n20974, \asqrt[50] , n_14021);
  and g34631 (n20978, n_13547, n_13546);
  and g34632 (n20979, \asqrt[6] , n20978);
  not g34633 (n_14022, n20979);
  and g34634 (n20980, n_13545, n_14022);
  not g34635 (n_14023, n20977);
  not g34636 (n_14024, n20980);
  and g34637 (n20981, n_14023, n_14024);
  and g34638 (n20982, n_1082, n_14019);
  and g34639 (n20983, n_14020, n20982);
  not g34640 (n_14025, n20981);
  not g34641 (n_14026, n20983);
  and g34642 (n20984, n_14025, n_14026);
  not g34643 (n_14027, n20974);
  not g34644 (n_14028, n20984);
  and g34645 (n20985, n_14027, n_14028);
  not g34646 (n_14029, n20985);
  and g34647 (n20986, \asqrt[51] , n_14029);
  and g34651 (n20990, n_13555, n_13554);
  and g34652 (n20991, \asqrt[6] , n20990);
  not g34653 (n_14030, n20991);
  and g34654 (n20992, n_13553, n_14030);
  not g34655 (n_14031, n20989);
  not g34656 (n_14032, n20992);
  and g34657 (n20993, n_14031, n_14032);
  and g34658 (n20994, n_954, n_14027);
  and g34659 (n20995, n_14028, n20994);
  not g34660 (n_14033, n20993);
  not g34661 (n_14034, n20995);
  and g34662 (n20996, n_14033, n_14034);
  not g34663 (n_14035, n20986);
  not g34664 (n_14036, n20996);
  and g34665 (n20997, n_14035, n_14036);
  not g34666 (n_14037, n20997);
  and g34667 (n20998, \asqrt[52] , n_14037);
  and g34671 (n21002, n_13563, n_13562);
  and g34672 (n21003, \asqrt[6] , n21002);
  not g34673 (n_14038, n21003);
  and g34674 (n21004, n_13561, n_14038);
  not g34675 (n_14039, n21001);
  not g34676 (n_14040, n21004);
  and g34677 (n21005, n_14039, n_14040);
  and g34678 (n21006, n_834, n_14035);
  and g34679 (n21007, n_14036, n21006);
  not g34680 (n_14041, n21005);
  not g34681 (n_14042, n21007);
  and g34682 (n21008, n_14041, n_14042);
  not g34683 (n_14043, n20998);
  not g34684 (n_14044, n21008);
  and g34685 (n21009, n_14043, n_14044);
  not g34686 (n_14045, n21009);
  and g34687 (n21010, \asqrt[53] , n_14045);
  and g34691 (n21014, n_13571, n_13570);
  and g34692 (n21015, \asqrt[6] , n21014);
  not g34693 (n_14046, n21015);
  and g34694 (n21016, n_13569, n_14046);
  not g34695 (n_14047, n21013);
  not g34696 (n_14048, n21016);
  and g34697 (n21017, n_14047, n_14048);
  and g34698 (n21018, n_722, n_14043);
  and g34699 (n21019, n_14044, n21018);
  not g34700 (n_14049, n21017);
  not g34701 (n_14050, n21019);
  and g34702 (n21020, n_14049, n_14050);
  not g34703 (n_14051, n21010);
  not g34704 (n_14052, n21020);
  and g34705 (n21021, n_14051, n_14052);
  not g34706 (n_14053, n21021);
  and g34707 (n21022, \asqrt[54] , n_14053);
  and g34711 (n21026, n_13579, n_13578);
  and g34712 (n21027, \asqrt[6] , n21026);
  not g34713 (n_14054, n21027);
  and g34714 (n21028, n_13577, n_14054);
  not g34715 (n_14055, n21025);
  not g34716 (n_14056, n21028);
  and g34717 (n21029, n_14055, n_14056);
  and g34718 (n21030, n_618, n_14051);
  and g34719 (n21031, n_14052, n21030);
  not g34720 (n_14057, n21029);
  not g34721 (n_14058, n21031);
  and g34722 (n21032, n_14057, n_14058);
  not g34723 (n_14059, n21022);
  not g34724 (n_14060, n21032);
  and g34725 (n21033, n_14059, n_14060);
  not g34726 (n_14061, n21033);
  and g34727 (n21034, \asqrt[55] , n_14061);
  and g34731 (n21038, n_13587, n_13586);
  and g34732 (n21039, \asqrt[6] , n21038);
  not g34733 (n_14062, n21039);
  and g34734 (n21040, n_13585, n_14062);
  not g34735 (n_14063, n21037);
  not g34736 (n_14064, n21040);
  and g34737 (n21041, n_14063, n_14064);
  and g34738 (n21042, n_522, n_14059);
  and g34739 (n21043, n_14060, n21042);
  not g34740 (n_14065, n21041);
  not g34741 (n_14066, n21043);
  and g34742 (n21044, n_14065, n_14066);
  not g34743 (n_14067, n21034);
  not g34744 (n_14068, n21044);
  and g34745 (n21045, n_14067, n_14068);
  not g34746 (n_14069, n21045);
  and g34747 (n21046, \asqrt[56] , n_14069);
  and g34751 (n21050, n_13595, n_13594);
  and g34752 (n21051, \asqrt[6] , n21050);
  not g34753 (n_14070, n21051);
  and g34754 (n21052, n_13593, n_14070);
  not g34755 (n_14071, n21049);
  not g34756 (n_14072, n21052);
  and g34757 (n21053, n_14071, n_14072);
  and g34758 (n21054, n_434, n_14067);
  and g34759 (n21055, n_14068, n21054);
  not g34760 (n_14073, n21053);
  not g34761 (n_14074, n21055);
  and g34762 (n21056, n_14073, n_14074);
  not g34763 (n_14075, n21046);
  not g34764 (n_14076, n21056);
  and g34765 (n21057, n_14075, n_14076);
  not g34766 (n_14077, n21057);
  and g34767 (n21058, \asqrt[57] , n_14077);
  and g34771 (n21062, n_13603, n_13602);
  and g34772 (n21063, \asqrt[6] , n21062);
  not g34773 (n_14078, n21063);
  and g34774 (n21064, n_13601, n_14078);
  not g34775 (n_14079, n21061);
  not g34776 (n_14080, n21064);
  and g34777 (n21065, n_14079, n_14080);
  and g34778 (n21066, n_354, n_14075);
  and g34779 (n21067, n_14076, n21066);
  not g34780 (n_14081, n21065);
  not g34781 (n_14082, n21067);
  and g34782 (n21068, n_14081, n_14082);
  not g34783 (n_14083, n21058);
  not g34784 (n_14084, n21068);
  and g34785 (n21069, n_14083, n_14084);
  not g34786 (n_14085, n21069);
  and g34787 (n21070, \asqrt[58] , n_14085);
  and g34791 (n21074, n_13611, n_13610);
  and g34792 (n21075, \asqrt[6] , n21074);
  not g34793 (n_14086, n21075);
  and g34794 (n21076, n_13609, n_14086);
  not g34795 (n_14087, n21073);
  not g34796 (n_14088, n21076);
  and g34797 (n21077, n_14087, n_14088);
  and g34798 (n21078, n_282, n_14083);
  and g34799 (n21079, n_14084, n21078);
  not g34800 (n_14089, n21077);
  not g34801 (n_14090, n21079);
  and g34802 (n21080, n_14089, n_14090);
  not g34803 (n_14091, n21070);
  not g34804 (n_14092, n21080);
  and g34805 (n21081, n_14091, n_14092);
  not g34806 (n_14093, n21081);
  and g34807 (n21082, \asqrt[59] , n_14093);
  and g34808 (n21083, n_218, n_14091);
  and g34809 (n21084, n_14092, n21083);
  and g34813 (n21088, n_13619, n_13617);
  and g34814 (n21089, \asqrt[6] , n21088);
  not g34815 (n_14094, n21089);
  and g34816 (n21090, n_13618, n_14094);
  not g34817 (n_14095, n21087);
  not g34818 (n_14096, n21090);
  and g34819 (n21091, n_14095, n_14096);
  not g34820 (n_14097, n21084);
  not g34821 (n_14098, n21091);
  and g34822 (n21092, n_14097, n_14098);
  not g34823 (n_14099, n21082);
  not g34824 (n_14100, n21092);
  and g34825 (n21093, n_14099, n_14100);
  not g34826 (n_14101, n21093);
  and g34827 (n21094, \asqrt[60] , n_14101);
  and g34831 (n21098, n_13627, n_13626);
  and g34832 (n21099, \asqrt[6] , n21098);
  not g34833 (n_14102, n21099);
  and g34834 (n21100, n_13625, n_14102);
  not g34835 (n_14103, n21097);
  not g34836 (n_14104, n21100);
  and g34837 (n21101, n_14103, n_14104);
  and g34838 (n21102, n_162, n_14099);
  and g34839 (n21103, n_14100, n21102);
  not g34840 (n_14105, n21101);
  not g34841 (n_14106, n21103);
  and g34842 (n21104, n_14105, n_14106);
  not g34843 (n_14107, n21094);
  not g34844 (n_14108, n21104);
  and g34845 (n21105, n_14107, n_14108);
  not g34846 (n_14109, n21105);
  and g34847 (n21106, \asqrt[61] , n_14109);
  and g34851 (n21110, n_13635, n_13634);
  and g34852 (n21111, \asqrt[6] , n21110);
  not g34853 (n_14110, n21111);
  and g34854 (n21112, n_13633, n_14110);
  not g34855 (n_14111, n21109);
  not g34856 (n_14112, n21112);
  and g34857 (n21113, n_14111, n_14112);
  and g34858 (n21114, n_115, n_14107);
  and g34859 (n21115, n_14108, n21114);
  not g34860 (n_14113, n21113);
  not g34861 (n_14114, n21115);
  and g34862 (n21116, n_14113, n_14114);
  not g34863 (n_14115, n21106);
  not g34864 (n_14116, n21116);
  and g34865 (n21117, n_14115, n_14116);
  not g34866 (n_14117, n21117);
  and g34867 (n21118, \asqrt[62] , n_14117);
  and g34871 (n21122, n_13643, n_13642);
  and g34872 (n21123, \asqrt[6] , n21122);
  not g34873 (n_14118, n21123);
  and g34874 (n21124, n_13641, n_14118);
  not g34875 (n_14119, n21121);
  not g34876 (n_14120, n21124);
  and g34877 (n21125, n_14119, n_14120);
  and g34878 (n21126, n_76, n_14115);
  and g34879 (n21127, n_14116, n21126);
  not g34880 (n_14121, n21125);
  not g34881 (n_14122, n21127);
  and g34882 (n21128, n_14121, n_14122);
  not g34883 (n_14123, n21118);
  not g34884 (n_14124, n21128);
  and g34885 (n21129, n_14123, n_14124);
  and g34889 (n21133, n_13651, n_13650);
  and g34890 (n21134, \asqrt[6] , n21133);
  not g34891 (n_14125, n21134);
  and g34892 (n21135, n_13649, n_14125);
  not g34893 (n_14126, n21132);
  not g34894 (n_14127, n21135);
  and g34895 (n21136, n_14126, n_14127);
  and g34896 (n21137, n_13658, n_13657);
  and g34897 (n21138, \asqrt[6] , n21137);
  not g34900 (n_14129, n21136);
  not g34902 (n_14130, n21129);
  not g34904 (n_14131, n21141);
  and g34905 (n21142, n_21, n_14131);
  and g34906 (n21143, n_14123, n21136);
  and g34907 (n21144, n_14124, n21143);
  and g34908 (n21145, n_13657, \asqrt[6] );
  not g34909 (n_14132, n21145);
  and g34910 (n21146, n20425, n_14132);
  not g34911 (n_14133, n21137);
  and g34912 (n21147, \asqrt[63] , n_14133);
  not g34913 (n_14134, n21146);
  and g34914 (n21148, n_14134, n21147);
  not g34915 (n_14135, n21144);
  not g34916 (n_14136, n21148);
  and g34917 (n21149, n_14135, n_14136);
  not g34918 (n_14137, n21149);
  or g34919 (\asqrt[5] , n21142, n_14137);
  and g34920 (n21151, \a[10] , \asqrt[5] );
  not g34921 (n_14141, \a[8] );
  not g34922 (n_14142, \a[9] );
  and g34923 (n21152, n_14141, n_14142);
  and g34924 (n21153, n_13670, n21152);
  not g34925 (n_14143, n21151);
  not g34926 (n_14144, n21153);
  and g34927 (n21154, n_14143, n_14144);
  not g34928 (n_14145, n21154);
  and g34929 (n21155, \asqrt[6] , n_14145);
  and g34935 (n21161, n_13670, \asqrt[5] );
  not g34936 (n_14146, n21161);
  and g34937 (n21162, \a[11] , n_14146);
  and g34938 (n21163, n20454, \asqrt[5] );
  not g34939 (n_14147, n21162);
  not g34940 (n_14148, n21163);
  and g34941 (n21164, n_14147, n_14148);
  not g34942 (n_14149, n21160);
  and g34943 (n21165, n_14149, n21164);
  not g34944 (n_14150, n21155);
  not g34945 (n_14151, n21165);
  and g34946 (n21166, n_14150, n_14151);
  not g34947 (n_14152, n21166);
  and g34948 (n21167, \asqrt[7] , n_14152);
  not g34949 (n_14153, \asqrt[7] );
  and g34950 (n21168, n_14153, n_14150);
  and g34951 (n21169, n_14151, n21168);
  not g34954 (n_14154, n21142);
  not g34956 (n_14155, n21172);
  and g34957 (n21173, n_14148, n_14155);
  not g34958 (n_14156, n21173);
  and g34959 (n21174, \a[12] , n_14156);
  and g34960 (n21175, n_13206, n_14155);
  and g34961 (n21176, n_14148, n21175);
  not g34962 (n_14157, n21174);
  not g34963 (n_14158, n21176);
  and g34964 (n21177, n_14157, n_14158);
  not g34965 (n_14159, n21169);
  not g34966 (n_14160, n21177);
  and g34967 (n21178, n_14159, n_14160);
  not g34968 (n_14161, n21167);
  not g34969 (n_14162, n21178);
  and g34970 (n21179, n_14161, n_14162);
  not g34971 (n_14163, n21179);
  and g34972 (n21180, \asqrt[8] , n_14163);
  and g34973 (n21181, n_13679, n_13678);
  not g34974 (n_14164, n20466);
  and g34975 (n21182, n_14164, n21181);
  and g34976 (n21183, \asqrt[5] , n21182);
  and g34977 (n21184, \asqrt[5] , n21181);
  not g34978 (n_14165, n21184);
  and g34979 (n21185, n20466, n_14165);
  not g34980 (n_14166, n21183);
  not g34981 (n_14167, n21185);
  and g34982 (n21186, n_14166, n_14167);
  and g34983 (n21187, n_13682, n_14161);
  and g34984 (n21188, n_14162, n21187);
  not g34985 (n_14168, n21186);
  not g34986 (n_14169, n21188);
  and g34987 (n21189, n_14168, n_14169);
  not g34988 (n_14170, n21180);
  not g34989 (n_14171, n21189);
  and g34990 (n21190, n_14170, n_14171);
  not g34991 (n_14172, n21190);
  and g34992 (n21191, \asqrt[9] , n_14172);
  and g34996 (n21195, n_13690, n_13688);
  and g34997 (n21196, \asqrt[5] , n21195);
  not g34998 (n_14173, n21196);
  and g34999 (n21197, n_13689, n_14173);
  not g35000 (n_14174, n21194);
  not g35001 (n_14175, n21197);
  and g35002 (n21198, n_14174, n_14175);
  and g35003 (n21199, n_13218, n_14170);
  and g35004 (n21200, n_14171, n21199);
  not g35005 (n_14176, n21198);
  not g35006 (n_14177, n21200);
  and g35007 (n21201, n_14176, n_14177);
  not g35008 (n_14178, n21191);
  not g35009 (n_14179, n21201);
  and g35010 (n21202, n_14178, n_14179);
  not g35011 (n_14180, n21202);
  and g35012 (n21203, \asqrt[10] , n_14180);
  and g35016 (n21207, n_13699, n_13698);
  and g35017 (n21208, \asqrt[5] , n21207);
  not g35018 (n_14181, n21208);
  and g35019 (n21209, n_13697, n_14181);
  not g35020 (n_14182, n21206);
  not g35021 (n_14183, n21209);
  and g35022 (n21210, n_14182, n_14183);
  and g35023 (n21211, n_12762, n_14178);
  and g35024 (n21212, n_14179, n21211);
  not g35025 (n_14184, n21210);
  not g35026 (n_14185, n21212);
  and g35027 (n21213, n_14184, n_14185);
  not g35028 (n_14186, n21203);
  not g35029 (n_14187, n21213);
  and g35030 (n21214, n_14186, n_14187);
  not g35031 (n_14188, n21214);
  and g35032 (n21215, \asqrt[11] , n_14188);
  and g35036 (n21219, n_13707, n_13706);
  and g35037 (n21220, \asqrt[5] , n21219);
  not g35038 (n_14189, n21220);
  and g35039 (n21221, n_13705, n_14189);
  not g35040 (n_14190, n21218);
  not g35041 (n_14191, n21221);
  and g35042 (n21222, n_14190, n_14191);
  and g35043 (n21223, n_12314, n_14186);
  and g35044 (n21224, n_14187, n21223);
  not g35045 (n_14192, n21222);
  not g35046 (n_14193, n21224);
  and g35047 (n21225, n_14192, n_14193);
  not g35048 (n_14194, n21215);
  not g35049 (n_14195, n21225);
  and g35050 (n21226, n_14194, n_14195);
  not g35051 (n_14196, n21226);
  and g35052 (n21227, \asqrt[12] , n_14196);
  and g35056 (n21231, n_13715, n_13714);
  and g35057 (n21232, \asqrt[5] , n21231);
  not g35058 (n_14197, n21232);
  and g35059 (n21233, n_13713, n_14197);
  not g35060 (n_14198, n21230);
  not g35061 (n_14199, n21233);
  and g35062 (n21234, n_14198, n_14199);
  and g35063 (n21235, n_11874, n_14194);
  and g35064 (n21236, n_14195, n21235);
  not g35065 (n_14200, n21234);
  not g35066 (n_14201, n21236);
  and g35067 (n21237, n_14200, n_14201);
  not g35068 (n_14202, n21227);
  not g35069 (n_14203, n21237);
  and g35070 (n21238, n_14202, n_14203);
  not g35071 (n_14204, n21238);
  and g35072 (n21239, \asqrt[13] , n_14204);
  and g35076 (n21243, n_13723, n_13722);
  and g35077 (n21244, \asqrt[5] , n21243);
  not g35078 (n_14205, n21244);
  and g35079 (n21245, n_13721, n_14205);
  not g35080 (n_14206, n21242);
  not g35081 (n_14207, n21245);
  and g35082 (n21246, n_14206, n_14207);
  and g35083 (n21247, n_11442, n_14202);
  and g35084 (n21248, n_14203, n21247);
  not g35085 (n_14208, n21246);
  not g35086 (n_14209, n21248);
  and g35087 (n21249, n_14208, n_14209);
  not g35088 (n_14210, n21239);
  not g35089 (n_14211, n21249);
  and g35090 (n21250, n_14210, n_14211);
  not g35091 (n_14212, n21250);
  and g35092 (n21251, \asqrt[14] , n_14212);
  and g35096 (n21255, n_13731, n_13730);
  and g35097 (n21256, \asqrt[5] , n21255);
  not g35098 (n_14213, n21256);
  and g35099 (n21257, n_13729, n_14213);
  not g35100 (n_14214, n21254);
  not g35101 (n_14215, n21257);
  and g35102 (n21258, n_14214, n_14215);
  and g35103 (n21259, n_11018, n_14210);
  and g35104 (n21260, n_14211, n21259);
  not g35105 (n_14216, n21258);
  not g35106 (n_14217, n21260);
  and g35107 (n21261, n_14216, n_14217);
  not g35108 (n_14218, n21251);
  not g35109 (n_14219, n21261);
  and g35110 (n21262, n_14218, n_14219);
  not g35111 (n_14220, n21262);
  and g35112 (n21263, \asqrt[15] , n_14220);
  and g35116 (n21267, n_13739, n_13738);
  and g35117 (n21268, \asqrt[5] , n21267);
  not g35118 (n_14221, n21268);
  and g35119 (n21269, n_13737, n_14221);
  not g35120 (n_14222, n21266);
  not g35121 (n_14223, n21269);
  and g35122 (n21270, n_14222, n_14223);
  and g35123 (n21271, n_10602, n_14218);
  and g35124 (n21272, n_14219, n21271);
  not g35125 (n_14224, n21270);
  not g35126 (n_14225, n21272);
  and g35127 (n21273, n_14224, n_14225);
  not g35128 (n_14226, n21263);
  not g35129 (n_14227, n21273);
  and g35130 (n21274, n_14226, n_14227);
  not g35131 (n_14228, n21274);
  and g35132 (n21275, \asqrt[16] , n_14228);
  and g35136 (n21279, n_13747, n_13746);
  and g35137 (n21280, \asqrt[5] , n21279);
  not g35138 (n_14229, n21280);
  and g35139 (n21281, n_13745, n_14229);
  not g35140 (n_14230, n21278);
  not g35141 (n_14231, n21281);
  and g35142 (n21282, n_14230, n_14231);
  and g35143 (n21283, n_10194, n_14226);
  and g35144 (n21284, n_14227, n21283);
  not g35145 (n_14232, n21282);
  not g35146 (n_14233, n21284);
  and g35147 (n21285, n_14232, n_14233);
  not g35148 (n_14234, n21275);
  not g35149 (n_14235, n21285);
  and g35150 (n21286, n_14234, n_14235);
  not g35151 (n_14236, n21286);
  and g35152 (n21287, \asqrt[17] , n_14236);
  and g35156 (n21291, n_13755, n_13754);
  and g35157 (n21292, \asqrt[5] , n21291);
  not g35158 (n_14237, n21292);
  and g35159 (n21293, n_13753, n_14237);
  not g35160 (n_14238, n21290);
  not g35161 (n_14239, n21293);
  and g35162 (n21294, n_14238, n_14239);
  and g35163 (n21295, n_9794, n_14234);
  and g35164 (n21296, n_14235, n21295);
  not g35165 (n_14240, n21294);
  not g35166 (n_14241, n21296);
  and g35167 (n21297, n_14240, n_14241);
  not g35168 (n_14242, n21287);
  not g35169 (n_14243, n21297);
  and g35170 (n21298, n_14242, n_14243);
  not g35171 (n_14244, n21298);
  and g35172 (n21299, \asqrt[18] , n_14244);
  and g35176 (n21303, n_13763, n_13762);
  and g35177 (n21304, \asqrt[5] , n21303);
  not g35178 (n_14245, n21304);
  and g35179 (n21305, n_13761, n_14245);
  not g35180 (n_14246, n21302);
  not g35181 (n_14247, n21305);
  and g35182 (n21306, n_14246, n_14247);
  and g35183 (n21307, n_9402, n_14242);
  and g35184 (n21308, n_14243, n21307);
  not g35185 (n_14248, n21306);
  not g35186 (n_14249, n21308);
  and g35187 (n21309, n_14248, n_14249);
  not g35188 (n_14250, n21299);
  not g35189 (n_14251, n21309);
  and g35190 (n21310, n_14250, n_14251);
  not g35191 (n_14252, n21310);
  and g35192 (n21311, \asqrt[19] , n_14252);
  and g35196 (n21315, n_13771, n_13770);
  and g35197 (n21316, \asqrt[5] , n21315);
  not g35198 (n_14253, n21316);
  and g35199 (n21317, n_13769, n_14253);
  not g35200 (n_14254, n21314);
  not g35201 (n_14255, n21317);
  and g35202 (n21318, n_14254, n_14255);
  and g35203 (n21319, n_9018, n_14250);
  and g35204 (n21320, n_14251, n21319);
  not g35205 (n_14256, n21318);
  not g35206 (n_14257, n21320);
  and g35207 (n21321, n_14256, n_14257);
  not g35208 (n_14258, n21311);
  not g35209 (n_14259, n21321);
  and g35210 (n21322, n_14258, n_14259);
  not g35211 (n_14260, n21322);
  and g35212 (n21323, \asqrt[20] , n_14260);
  and g35216 (n21327, n_13779, n_13778);
  and g35217 (n21328, \asqrt[5] , n21327);
  not g35218 (n_14261, n21328);
  and g35219 (n21329, n_13777, n_14261);
  not g35220 (n_14262, n21326);
  not g35221 (n_14263, n21329);
  and g35222 (n21330, n_14262, n_14263);
  and g35223 (n21331, n_8642, n_14258);
  and g35224 (n21332, n_14259, n21331);
  not g35225 (n_14264, n21330);
  not g35226 (n_14265, n21332);
  and g35227 (n21333, n_14264, n_14265);
  not g35228 (n_14266, n21323);
  not g35229 (n_14267, n21333);
  and g35230 (n21334, n_14266, n_14267);
  not g35231 (n_14268, n21334);
  and g35232 (n21335, \asqrt[21] , n_14268);
  and g35236 (n21339, n_13787, n_13786);
  and g35237 (n21340, \asqrt[5] , n21339);
  not g35238 (n_14269, n21340);
  and g35239 (n21341, n_13785, n_14269);
  not g35240 (n_14270, n21338);
  not g35241 (n_14271, n21341);
  and g35242 (n21342, n_14270, n_14271);
  and g35243 (n21343, n_8274, n_14266);
  and g35244 (n21344, n_14267, n21343);
  not g35245 (n_14272, n21342);
  not g35246 (n_14273, n21344);
  and g35247 (n21345, n_14272, n_14273);
  not g35248 (n_14274, n21335);
  not g35249 (n_14275, n21345);
  and g35250 (n21346, n_14274, n_14275);
  not g35251 (n_14276, n21346);
  and g35252 (n21347, \asqrt[22] , n_14276);
  and g35256 (n21351, n_13795, n_13794);
  and g35257 (n21352, \asqrt[5] , n21351);
  not g35258 (n_14277, n21352);
  and g35259 (n21353, n_13793, n_14277);
  not g35260 (n_14278, n21350);
  not g35261 (n_14279, n21353);
  and g35262 (n21354, n_14278, n_14279);
  and g35263 (n21355, n_7914, n_14274);
  and g35264 (n21356, n_14275, n21355);
  not g35265 (n_14280, n21354);
  not g35266 (n_14281, n21356);
  and g35267 (n21357, n_14280, n_14281);
  not g35268 (n_14282, n21347);
  not g35269 (n_14283, n21357);
  and g35270 (n21358, n_14282, n_14283);
  not g35271 (n_14284, n21358);
  and g35272 (n21359, \asqrt[23] , n_14284);
  and g35276 (n21363, n_13803, n_13802);
  and g35277 (n21364, \asqrt[5] , n21363);
  not g35278 (n_14285, n21364);
  and g35279 (n21365, n_13801, n_14285);
  not g35280 (n_14286, n21362);
  not g35281 (n_14287, n21365);
  and g35282 (n21366, n_14286, n_14287);
  and g35283 (n21367, n_7562, n_14282);
  and g35284 (n21368, n_14283, n21367);
  not g35285 (n_14288, n21366);
  not g35286 (n_14289, n21368);
  and g35287 (n21369, n_14288, n_14289);
  not g35288 (n_14290, n21359);
  not g35289 (n_14291, n21369);
  and g35290 (n21370, n_14290, n_14291);
  not g35291 (n_14292, n21370);
  and g35292 (n21371, \asqrt[24] , n_14292);
  and g35296 (n21375, n_13811, n_13810);
  and g35297 (n21376, \asqrt[5] , n21375);
  not g35298 (n_14293, n21376);
  and g35299 (n21377, n_13809, n_14293);
  not g35300 (n_14294, n21374);
  not g35301 (n_14295, n21377);
  and g35302 (n21378, n_14294, n_14295);
  and g35303 (n21379, n_7218, n_14290);
  and g35304 (n21380, n_14291, n21379);
  not g35305 (n_14296, n21378);
  not g35306 (n_14297, n21380);
  and g35307 (n21381, n_14296, n_14297);
  not g35308 (n_14298, n21371);
  not g35309 (n_14299, n21381);
  and g35310 (n21382, n_14298, n_14299);
  not g35311 (n_14300, n21382);
  and g35312 (n21383, \asqrt[25] , n_14300);
  and g35316 (n21387, n_13819, n_13818);
  and g35317 (n21388, \asqrt[5] , n21387);
  not g35318 (n_14301, n21388);
  and g35319 (n21389, n_13817, n_14301);
  not g35320 (n_14302, n21386);
  not g35321 (n_14303, n21389);
  and g35322 (n21390, n_14302, n_14303);
  and g35323 (n21391, n_6882, n_14298);
  and g35324 (n21392, n_14299, n21391);
  not g35325 (n_14304, n21390);
  not g35326 (n_14305, n21392);
  and g35327 (n21393, n_14304, n_14305);
  not g35328 (n_14306, n21383);
  not g35329 (n_14307, n21393);
  and g35330 (n21394, n_14306, n_14307);
  not g35331 (n_14308, n21394);
  and g35332 (n21395, \asqrt[26] , n_14308);
  and g35336 (n21399, n_13827, n_13826);
  and g35337 (n21400, \asqrt[5] , n21399);
  not g35338 (n_14309, n21400);
  and g35339 (n21401, n_13825, n_14309);
  not g35340 (n_14310, n21398);
  not g35341 (n_14311, n21401);
  and g35342 (n21402, n_14310, n_14311);
  and g35343 (n21403, n_6554, n_14306);
  and g35344 (n21404, n_14307, n21403);
  not g35345 (n_14312, n21402);
  not g35346 (n_14313, n21404);
  and g35347 (n21405, n_14312, n_14313);
  not g35348 (n_14314, n21395);
  not g35349 (n_14315, n21405);
  and g35350 (n21406, n_14314, n_14315);
  not g35351 (n_14316, n21406);
  and g35352 (n21407, \asqrt[27] , n_14316);
  and g35356 (n21411, n_13835, n_13834);
  and g35357 (n21412, \asqrt[5] , n21411);
  not g35358 (n_14317, n21412);
  and g35359 (n21413, n_13833, n_14317);
  not g35360 (n_14318, n21410);
  not g35361 (n_14319, n21413);
  and g35362 (n21414, n_14318, n_14319);
  and g35363 (n21415, n_6234, n_14314);
  and g35364 (n21416, n_14315, n21415);
  not g35365 (n_14320, n21414);
  not g35366 (n_14321, n21416);
  and g35367 (n21417, n_14320, n_14321);
  not g35368 (n_14322, n21407);
  not g35369 (n_14323, n21417);
  and g35370 (n21418, n_14322, n_14323);
  not g35371 (n_14324, n21418);
  and g35372 (n21419, \asqrt[28] , n_14324);
  and g35376 (n21423, n_13843, n_13842);
  and g35377 (n21424, \asqrt[5] , n21423);
  not g35378 (n_14325, n21424);
  and g35379 (n21425, n_13841, n_14325);
  not g35380 (n_14326, n21422);
  not g35381 (n_14327, n21425);
  and g35382 (n21426, n_14326, n_14327);
  and g35383 (n21427, n_5922, n_14322);
  and g35384 (n21428, n_14323, n21427);
  not g35385 (n_14328, n21426);
  not g35386 (n_14329, n21428);
  and g35387 (n21429, n_14328, n_14329);
  not g35388 (n_14330, n21419);
  not g35389 (n_14331, n21429);
  and g35390 (n21430, n_14330, n_14331);
  not g35391 (n_14332, n21430);
  and g35392 (n21431, \asqrt[29] , n_14332);
  and g35396 (n21435, n_13851, n_13850);
  and g35397 (n21436, \asqrt[5] , n21435);
  not g35398 (n_14333, n21436);
  and g35399 (n21437, n_13849, n_14333);
  not g35400 (n_14334, n21434);
  not g35401 (n_14335, n21437);
  and g35402 (n21438, n_14334, n_14335);
  and g35403 (n21439, n_5618, n_14330);
  and g35404 (n21440, n_14331, n21439);
  not g35405 (n_14336, n21438);
  not g35406 (n_14337, n21440);
  and g35407 (n21441, n_14336, n_14337);
  not g35408 (n_14338, n21431);
  not g35409 (n_14339, n21441);
  and g35410 (n21442, n_14338, n_14339);
  not g35411 (n_14340, n21442);
  and g35412 (n21443, \asqrt[30] , n_14340);
  and g35416 (n21447, n_13859, n_13858);
  and g35417 (n21448, \asqrt[5] , n21447);
  not g35418 (n_14341, n21448);
  and g35419 (n21449, n_13857, n_14341);
  not g35420 (n_14342, n21446);
  not g35421 (n_14343, n21449);
  and g35422 (n21450, n_14342, n_14343);
  and g35423 (n21451, n_5322, n_14338);
  and g35424 (n21452, n_14339, n21451);
  not g35425 (n_14344, n21450);
  not g35426 (n_14345, n21452);
  and g35427 (n21453, n_14344, n_14345);
  not g35428 (n_14346, n21443);
  not g35429 (n_14347, n21453);
  and g35430 (n21454, n_14346, n_14347);
  not g35431 (n_14348, n21454);
  and g35432 (n21455, \asqrt[31] , n_14348);
  and g35436 (n21459, n_13867, n_13866);
  and g35437 (n21460, \asqrt[5] , n21459);
  not g35438 (n_14349, n21460);
  and g35439 (n21461, n_13865, n_14349);
  not g35440 (n_14350, n21458);
  not g35441 (n_14351, n21461);
  and g35442 (n21462, n_14350, n_14351);
  and g35443 (n21463, n_5034, n_14346);
  and g35444 (n21464, n_14347, n21463);
  not g35445 (n_14352, n21462);
  not g35446 (n_14353, n21464);
  and g35447 (n21465, n_14352, n_14353);
  not g35448 (n_14354, n21455);
  not g35449 (n_14355, n21465);
  and g35450 (n21466, n_14354, n_14355);
  not g35451 (n_14356, n21466);
  and g35452 (n21467, \asqrt[32] , n_14356);
  and g35456 (n21471, n_13875, n_13874);
  and g35457 (n21472, \asqrt[5] , n21471);
  not g35458 (n_14357, n21472);
  and g35459 (n21473, n_13873, n_14357);
  not g35460 (n_14358, n21470);
  not g35461 (n_14359, n21473);
  and g35462 (n21474, n_14358, n_14359);
  and g35463 (n21475, n_4754, n_14354);
  and g35464 (n21476, n_14355, n21475);
  not g35465 (n_14360, n21474);
  not g35466 (n_14361, n21476);
  and g35467 (n21477, n_14360, n_14361);
  not g35468 (n_14362, n21467);
  not g35469 (n_14363, n21477);
  and g35470 (n21478, n_14362, n_14363);
  not g35471 (n_14364, n21478);
  and g35472 (n21479, \asqrt[33] , n_14364);
  and g35476 (n21483, n_13883, n_13882);
  and g35477 (n21484, \asqrt[5] , n21483);
  not g35478 (n_14365, n21484);
  and g35479 (n21485, n_13881, n_14365);
  not g35480 (n_14366, n21482);
  not g35481 (n_14367, n21485);
  and g35482 (n21486, n_14366, n_14367);
  and g35483 (n21487, n_4482, n_14362);
  and g35484 (n21488, n_14363, n21487);
  not g35485 (n_14368, n21486);
  not g35486 (n_14369, n21488);
  and g35487 (n21489, n_14368, n_14369);
  not g35488 (n_14370, n21479);
  not g35489 (n_14371, n21489);
  and g35490 (n21490, n_14370, n_14371);
  not g35491 (n_14372, n21490);
  and g35492 (n21491, \asqrt[34] , n_14372);
  and g35496 (n21495, n_13891, n_13890);
  and g35497 (n21496, \asqrt[5] , n21495);
  not g35498 (n_14373, n21496);
  and g35499 (n21497, n_13889, n_14373);
  not g35500 (n_14374, n21494);
  not g35501 (n_14375, n21497);
  and g35502 (n21498, n_14374, n_14375);
  and g35503 (n21499, n_4218, n_14370);
  and g35504 (n21500, n_14371, n21499);
  not g35505 (n_14376, n21498);
  not g35506 (n_14377, n21500);
  and g35507 (n21501, n_14376, n_14377);
  not g35508 (n_14378, n21491);
  not g35509 (n_14379, n21501);
  and g35510 (n21502, n_14378, n_14379);
  not g35511 (n_14380, n21502);
  and g35512 (n21503, \asqrt[35] , n_14380);
  and g35516 (n21507, n_13899, n_13898);
  and g35517 (n21508, \asqrt[5] , n21507);
  not g35518 (n_14381, n21508);
  and g35519 (n21509, n_13897, n_14381);
  not g35520 (n_14382, n21506);
  not g35521 (n_14383, n21509);
  and g35522 (n21510, n_14382, n_14383);
  and g35523 (n21511, n_3962, n_14378);
  and g35524 (n21512, n_14379, n21511);
  not g35525 (n_14384, n21510);
  not g35526 (n_14385, n21512);
  and g35527 (n21513, n_14384, n_14385);
  not g35528 (n_14386, n21503);
  not g35529 (n_14387, n21513);
  and g35530 (n21514, n_14386, n_14387);
  not g35531 (n_14388, n21514);
  and g35532 (n21515, \asqrt[36] , n_14388);
  and g35536 (n21519, n_13907, n_13906);
  and g35537 (n21520, \asqrt[5] , n21519);
  not g35538 (n_14389, n21520);
  and g35539 (n21521, n_13905, n_14389);
  not g35540 (n_14390, n21518);
  not g35541 (n_14391, n21521);
  and g35542 (n21522, n_14390, n_14391);
  and g35543 (n21523, n_3714, n_14386);
  and g35544 (n21524, n_14387, n21523);
  not g35545 (n_14392, n21522);
  not g35546 (n_14393, n21524);
  and g35547 (n21525, n_14392, n_14393);
  not g35548 (n_14394, n21515);
  not g35549 (n_14395, n21525);
  and g35550 (n21526, n_14394, n_14395);
  not g35551 (n_14396, n21526);
  and g35552 (n21527, \asqrt[37] , n_14396);
  and g35556 (n21531, n_13915, n_13914);
  and g35557 (n21532, \asqrt[5] , n21531);
  not g35558 (n_14397, n21532);
  and g35559 (n21533, n_13913, n_14397);
  not g35560 (n_14398, n21530);
  not g35561 (n_14399, n21533);
  and g35562 (n21534, n_14398, n_14399);
  and g35563 (n21535, n_3474, n_14394);
  and g35564 (n21536, n_14395, n21535);
  not g35565 (n_14400, n21534);
  not g35566 (n_14401, n21536);
  and g35567 (n21537, n_14400, n_14401);
  not g35568 (n_14402, n21527);
  not g35569 (n_14403, n21537);
  and g35570 (n21538, n_14402, n_14403);
  not g35571 (n_14404, n21538);
  and g35572 (n21539, \asqrt[38] , n_14404);
  and g35576 (n21543, n_13923, n_13922);
  and g35577 (n21544, \asqrt[5] , n21543);
  not g35578 (n_14405, n21544);
  and g35579 (n21545, n_13921, n_14405);
  not g35580 (n_14406, n21542);
  not g35581 (n_14407, n21545);
  and g35582 (n21546, n_14406, n_14407);
  and g35583 (n21547, n_3242, n_14402);
  and g35584 (n21548, n_14403, n21547);
  not g35585 (n_14408, n21546);
  not g35586 (n_14409, n21548);
  and g35587 (n21549, n_14408, n_14409);
  not g35588 (n_14410, n21539);
  not g35589 (n_14411, n21549);
  and g35590 (n21550, n_14410, n_14411);
  not g35591 (n_14412, n21550);
  and g35592 (n21551, \asqrt[39] , n_14412);
  and g35596 (n21555, n_13931, n_13930);
  and g35597 (n21556, \asqrt[5] , n21555);
  not g35598 (n_14413, n21556);
  and g35599 (n21557, n_13929, n_14413);
  not g35600 (n_14414, n21554);
  not g35601 (n_14415, n21557);
  and g35602 (n21558, n_14414, n_14415);
  and g35603 (n21559, n_3018, n_14410);
  and g35604 (n21560, n_14411, n21559);
  not g35605 (n_14416, n21558);
  not g35606 (n_14417, n21560);
  and g35607 (n21561, n_14416, n_14417);
  not g35608 (n_14418, n21551);
  not g35609 (n_14419, n21561);
  and g35610 (n21562, n_14418, n_14419);
  not g35611 (n_14420, n21562);
  and g35612 (n21563, \asqrt[40] , n_14420);
  and g35616 (n21567, n_13939, n_13938);
  and g35617 (n21568, \asqrt[5] , n21567);
  not g35618 (n_14421, n21568);
  and g35619 (n21569, n_13937, n_14421);
  not g35620 (n_14422, n21566);
  not g35621 (n_14423, n21569);
  and g35622 (n21570, n_14422, n_14423);
  and g35623 (n21571, n_2802, n_14418);
  and g35624 (n21572, n_14419, n21571);
  not g35625 (n_14424, n21570);
  not g35626 (n_14425, n21572);
  and g35627 (n21573, n_14424, n_14425);
  not g35628 (n_14426, n21563);
  not g35629 (n_14427, n21573);
  and g35630 (n21574, n_14426, n_14427);
  not g35631 (n_14428, n21574);
  and g35632 (n21575, \asqrt[41] , n_14428);
  and g35636 (n21579, n_13947, n_13946);
  and g35637 (n21580, \asqrt[5] , n21579);
  not g35638 (n_14429, n21580);
  and g35639 (n21581, n_13945, n_14429);
  not g35640 (n_14430, n21578);
  not g35641 (n_14431, n21581);
  and g35642 (n21582, n_14430, n_14431);
  and g35643 (n21583, n_2594, n_14426);
  and g35644 (n21584, n_14427, n21583);
  not g35645 (n_14432, n21582);
  not g35646 (n_14433, n21584);
  and g35647 (n21585, n_14432, n_14433);
  not g35648 (n_14434, n21575);
  not g35649 (n_14435, n21585);
  and g35650 (n21586, n_14434, n_14435);
  not g35651 (n_14436, n21586);
  and g35652 (n21587, \asqrt[42] , n_14436);
  and g35656 (n21591, n_13955, n_13954);
  and g35657 (n21592, \asqrt[5] , n21591);
  not g35658 (n_14437, n21592);
  and g35659 (n21593, n_13953, n_14437);
  not g35660 (n_14438, n21590);
  not g35661 (n_14439, n21593);
  and g35662 (n21594, n_14438, n_14439);
  and g35663 (n21595, n_2394, n_14434);
  and g35664 (n21596, n_14435, n21595);
  not g35665 (n_14440, n21594);
  not g35666 (n_14441, n21596);
  and g35667 (n21597, n_14440, n_14441);
  not g35668 (n_14442, n21587);
  not g35669 (n_14443, n21597);
  and g35670 (n21598, n_14442, n_14443);
  not g35671 (n_14444, n21598);
  and g35672 (n21599, \asqrt[43] , n_14444);
  and g35676 (n21603, n_13963, n_13962);
  and g35677 (n21604, \asqrt[5] , n21603);
  not g35678 (n_14445, n21604);
  and g35679 (n21605, n_13961, n_14445);
  not g35680 (n_14446, n21602);
  not g35681 (n_14447, n21605);
  and g35682 (n21606, n_14446, n_14447);
  and g35683 (n21607, n_2202, n_14442);
  and g35684 (n21608, n_14443, n21607);
  not g35685 (n_14448, n21606);
  not g35686 (n_14449, n21608);
  and g35687 (n21609, n_14448, n_14449);
  not g35688 (n_14450, n21599);
  not g35689 (n_14451, n21609);
  and g35690 (n21610, n_14450, n_14451);
  not g35691 (n_14452, n21610);
  and g35692 (n21611, \asqrt[44] , n_14452);
  and g35696 (n21615, n_13971, n_13970);
  and g35697 (n21616, \asqrt[5] , n21615);
  not g35698 (n_14453, n21616);
  and g35699 (n21617, n_13969, n_14453);
  not g35700 (n_14454, n21614);
  not g35701 (n_14455, n21617);
  and g35702 (n21618, n_14454, n_14455);
  and g35703 (n21619, n_2018, n_14450);
  and g35704 (n21620, n_14451, n21619);
  not g35705 (n_14456, n21618);
  not g35706 (n_14457, n21620);
  and g35707 (n21621, n_14456, n_14457);
  not g35708 (n_14458, n21611);
  not g35709 (n_14459, n21621);
  and g35710 (n21622, n_14458, n_14459);
  not g35711 (n_14460, n21622);
  and g35712 (n21623, \asqrt[45] , n_14460);
  and g35716 (n21627, n_13979, n_13978);
  and g35717 (n21628, \asqrt[5] , n21627);
  not g35718 (n_14461, n21628);
  and g35719 (n21629, n_13977, n_14461);
  not g35720 (n_14462, n21626);
  not g35721 (n_14463, n21629);
  and g35722 (n21630, n_14462, n_14463);
  and g35723 (n21631, n_1842, n_14458);
  and g35724 (n21632, n_14459, n21631);
  not g35725 (n_14464, n21630);
  not g35726 (n_14465, n21632);
  and g35727 (n21633, n_14464, n_14465);
  not g35728 (n_14466, n21623);
  not g35729 (n_14467, n21633);
  and g35730 (n21634, n_14466, n_14467);
  not g35731 (n_14468, n21634);
  and g35732 (n21635, \asqrt[46] , n_14468);
  and g35736 (n21639, n_13987, n_13986);
  and g35737 (n21640, \asqrt[5] , n21639);
  not g35738 (n_14469, n21640);
  and g35739 (n21641, n_13985, n_14469);
  not g35740 (n_14470, n21638);
  not g35741 (n_14471, n21641);
  and g35742 (n21642, n_14470, n_14471);
  and g35743 (n21643, n_1674, n_14466);
  and g35744 (n21644, n_14467, n21643);
  not g35745 (n_14472, n21642);
  not g35746 (n_14473, n21644);
  and g35747 (n21645, n_14472, n_14473);
  not g35748 (n_14474, n21635);
  not g35749 (n_14475, n21645);
  and g35750 (n21646, n_14474, n_14475);
  not g35751 (n_14476, n21646);
  and g35752 (n21647, \asqrt[47] , n_14476);
  and g35756 (n21651, n_13995, n_13994);
  and g35757 (n21652, \asqrt[5] , n21651);
  not g35758 (n_14477, n21652);
  and g35759 (n21653, n_13993, n_14477);
  not g35760 (n_14478, n21650);
  not g35761 (n_14479, n21653);
  and g35762 (n21654, n_14478, n_14479);
  and g35763 (n21655, n_1514, n_14474);
  and g35764 (n21656, n_14475, n21655);
  not g35765 (n_14480, n21654);
  not g35766 (n_14481, n21656);
  and g35767 (n21657, n_14480, n_14481);
  not g35768 (n_14482, n21647);
  not g35769 (n_14483, n21657);
  and g35770 (n21658, n_14482, n_14483);
  not g35771 (n_14484, n21658);
  and g35772 (n21659, \asqrt[48] , n_14484);
  and g35776 (n21663, n_14003, n_14002);
  and g35777 (n21664, \asqrt[5] , n21663);
  not g35778 (n_14485, n21664);
  and g35779 (n21665, n_14001, n_14485);
  not g35780 (n_14486, n21662);
  not g35781 (n_14487, n21665);
  and g35782 (n21666, n_14486, n_14487);
  and g35783 (n21667, n_1362, n_14482);
  and g35784 (n21668, n_14483, n21667);
  not g35785 (n_14488, n21666);
  not g35786 (n_14489, n21668);
  and g35787 (n21669, n_14488, n_14489);
  not g35788 (n_14490, n21659);
  not g35789 (n_14491, n21669);
  and g35790 (n21670, n_14490, n_14491);
  not g35791 (n_14492, n21670);
  and g35792 (n21671, \asqrt[49] , n_14492);
  and g35796 (n21675, n_14011, n_14010);
  and g35797 (n21676, \asqrt[5] , n21675);
  not g35798 (n_14493, n21676);
  and g35799 (n21677, n_14009, n_14493);
  not g35800 (n_14494, n21674);
  not g35801 (n_14495, n21677);
  and g35802 (n21678, n_14494, n_14495);
  and g35803 (n21679, n_1218, n_14490);
  and g35804 (n21680, n_14491, n21679);
  not g35805 (n_14496, n21678);
  not g35806 (n_14497, n21680);
  and g35807 (n21681, n_14496, n_14497);
  not g35808 (n_14498, n21671);
  not g35809 (n_14499, n21681);
  and g35810 (n21682, n_14498, n_14499);
  not g35811 (n_14500, n21682);
  and g35812 (n21683, \asqrt[50] , n_14500);
  and g35816 (n21687, n_14019, n_14018);
  and g35817 (n21688, \asqrt[5] , n21687);
  not g35818 (n_14501, n21688);
  and g35819 (n21689, n_14017, n_14501);
  not g35820 (n_14502, n21686);
  not g35821 (n_14503, n21689);
  and g35822 (n21690, n_14502, n_14503);
  and g35823 (n21691, n_1082, n_14498);
  and g35824 (n21692, n_14499, n21691);
  not g35825 (n_14504, n21690);
  not g35826 (n_14505, n21692);
  and g35827 (n21693, n_14504, n_14505);
  not g35828 (n_14506, n21683);
  not g35829 (n_14507, n21693);
  and g35830 (n21694, n_14506, n_14507);
  not g35831 (n_14508, n21694);
  and g35832 (n21695, \asqrt[51] , n_14508);
  and g35836 (n21699, n_14027, n_14026);
  and g35837 (n21700, \asqrt[5] , n21699);
  not g35838 (n_14509, n21700);
  and g35839 (n21701, n_14025, n_14509);
  not g35840 (n_14510, n21698);
  not g35841 (n_14511, n21701);
  and g35842 (n21702, n_14510, n_14511);
  and g35843 (n21703, n_954, n_14506);
  and g35844 (n21704, n_14507, n21703);
  not g35845 (n_14512, n21702);
  not g35846 (n_14513, n21704);
  and g35847 (n21705, n_14512, n_14513);
  not g35848 (n_14514, n21695);
  not g35849 (n_14515, n21705);
  and g35850 (n21706, n_14514, n_14515);
  not g35851 (n_14516, n21706);
  and g35852 (n21707, \asqrt[52] , n_14516);
  and g35856 (n21711, n_14035, n_14034);
  and g35857 (n21712, \asqrt[5] , n21711);
  not g35858 (n_14517, n21712);
  and g35859 (n21713, n_14033, n_14517);
  not g35860 (n_14518, n21710);
  not g35861 (n_14519, n21713);
  and g35862 (n21714, n_14518, n_14519);
  and g35863 (n21715, n_834, n_14514);
  and g35864 (n21716, n_14515, n21715);
  not g35865 (n_14520, n21714);
  not g35866 (n_14521, n21716);
  and g35867 (n21717, n_14520, n_14521);
  not g35868 (n_14522, n21707);
  not g35869 (n_14523, n21717);
  and g35870 (n21718, n_14522, n_14523);
  not g35871 (n_14524, n21718);
  and g35872 (n21719, \asqrt[53] , n_14524);
  and g35876 (n21723, n_14043, n_14042);
  and g35877 (n21724, \asqrt[5] , n21723);
  not g35878 (n_14525, n21724);
  and g35879 (n21725, n_14041, n_14525);
  not g35880 (n_14526, n21722);
  not g35881 (n_14527, n21725);
  and g35882 (n21726, n_14526, n_14527);
  and g35883 (n21727, n_722, n_14522);
  and g35884 (n21728, n_14523, n21727);
  not g35885 (n_14528, n21726);
  not g35886 (n_14529, n21728);
  and g35887 (n21729, n_14528, n_14529);
  not g35888 (n_14530, n21719);
  not g35889 (n_14531, n21729);
  and g35890 (n21730, n_14530, n_14531);
  not g35891 (n_14532, n21730);
  and g35892 (n21731, \asqrt[54] , n_14532);
  and g35896 (n21735, n_14051, n_14050);
  and g35897 (n21736, \asqrt[5] , n21735);
  not g35898 (n_14533, n21736);
  and g35899 (n21737, n_14049, n_14533);
  not g35900 (n_14534, n21734);
  not g35901 (n_14535, n21737);
  and g35902 (n21738, n_14534, n_14535);
  and g35903 (n21739, n_618, n_14530);
  and g35904 (n21740, n_14531, n21739);
  not g35905 (n_14536, n21738);
  not g35906 (n_14537, n21740);
  and g35907 (n21741, n_14536, n_14537);
  not g35908 (n_14538, n21731);
  not g35909 (n_14539, n21741);
  and g35910 (n21742, n_14538, n_14539);
  not g35911 (n_14540, n21742);
  and g35912 (n21743, \asqrt[55] , n_14540);
  and g35916 (n21747, n_14059, n_14058);
  and g35917 (n21748, \asqrt[5] , n21747);
  not g35918 (n_14541, n21748);
  and g35919 (n21749, n_14057, n_14541);
  not g35920 (n_14542, n21746);
  not g35921 (n_14543, n21749);
  and g35922 (n21750, n_14542, n_14543);
  and g35923 (n21751, n_522, n_14538);
  and g35924 (n21752, n_14539, n21751);
  not g35925 (n_14544, n21750);
  not g35926 (n_14545, n21752);
  and g35927 (n21753, n_14544, n_14545);
  not g35928 (n_14546, n21743);
  not g35929 (n_14547, n21753);
  and g35930 (n21754, n_14546, n_14547);
  not g35931 (n_14548, n21754);
  and g35932 (n21755, \asqrt[56] , n_14548);
  and g35936 (n21759, n_14067, n_14066);
  and g35937 (n21760, \asqrt[5] , n21759);
  not g35938 (n_14549, n21760);
  and g35939 (n21761, n_14065, n_14549);
  not g35940 (n_14550, n21758);
  not g35941 (n_14551, n21761);
  and g35942 (n21762, n_14550, n_14551);
  and g35943 (n21763, n_434, n_14546);
  and g35944 (n21764, n_14547, n21763);
  not g35945 (n_14552, n21762);
  not g35946 (n_14553, n21764);
  and g35947 (n21765, n_14552, n_14553);
  not g35948 (n_14554, n21755);
  not g35949 (n_14555, n21765);
  and g35950 (n21766, n_14554, n_14555);
  not g35951 (n_14556, n21766);
  and g35952 (n21767, \asqrt[57] , n_14556);
  and g35956 (n21771, n_14075, n_14074);
  and g35957 (n21772, \asqrt[5] , n21771);
  not g35958 (n_14557, n21772);
  and g35959 (n21773, n_14073, n_14557);
  not g35960 (n_14558, n21770);
  not g35961 (n_14559, n21773);
  and g35962 (n21774, n_14558, n_14559);
  and g35963 (n21775, n_354, n_14554);
  and g35964 (n21776, n_14555, n21775);
  not g35965 (n_14560, n21774);
  not g35966 (n_14561, n21776);
  and g35967 (n21777, n_14560, n_14561);
  not g35968 (n_14562, n21767);
  not g35969 (n_14563, n21777);
  and g35970 (n21778, n_14562, n_14563);
  not g35971 (n_14564, n21778);
  and g35972 (n21779, \asqrt[58] , n_14564);
  and g35976 (n21783, n_14083, n_14082);
  and g35977 (n21784, \asqrt[5] , n21783);
  not g35978 (n_14565, n21784);
  and g35979 (n21785, n_14081, n_14565);
  not g35980 (n_14566, n21782);
  not g35981 (n_14567, n21785);
  and g35982 (n21786, n_14566, n_14567);
  and g35983 (n21787, n_282, n_14562);
  and g35984 (n21788, n_14563, n21787);
  not g35985 (n_14568, n21786);
  not g35986 (n_14569, n21788);
  and g35987 (n21789, n_14568, n_14569);
  not g35988 (n_14570, n21779);
  not g35989 (n_14571, n21789);
  and g35990 (n21790, n_14570, n_14571);
  not g35991 (n_14572, n21790);
  and g35992 (n21791, \asqrt[59] , n_14572);
  and g35996 (n21795, n_14091, n_14090);
  and g35997 (n21796, \asqrt[5] , n21795);
  not g35998 (n_14573, n21796);
  and g35999 (n21797, n_14089, n_14573);
  not g36000 (n_14574, n21794);
  not g36001 (n_14575, n21797);
  and g36002 (n21798, n_14574, n_14575);
  and g36003 (n21799, n_218, n_14570);
  and g36004 (n21800, n_14571, n21799);
  not g36005 (n_14576, n21798);
  not g36006 (n_14577, n21800);
  and g36007 (n21801, n_14576, n_14577);
  not g36008 (n_14578, n21791);
  not g36009 (n_14579, n21801);
  and g36010 (n21802, n_14578, n_14579);
  not g36011 (n_14580, n21802);
  and g36012 (n21803, \asqrt[60] , n_14580);
  and g36013 (n21804, n_162, n_14578);
  and g36014 (n21805, n_14579, n21804);
  and g36018 (n21809, n_14099, n_14097);
  and g36019 (n21810, \asqrt[5] , n21809);
  not g36020 (n_14581, n21810);
  and g36021 (n21811, n_14098, n_14581);
  not g36022 (n_14582, n21808);
  not g36023 (n_14583, n21811);
  and g36024 (n21812, n_14582, n_14583);
  not g36025 (n_14584, n21805);
  not g36026 (n_14585, n21812);
  and g36027 (n21813, n_14584, n_14585);
  not g36028 (n_14586, n21803);
  not g36029 (n_14587, n21813);
  and g36030 (n21814, n_14586, n_14587);
  not g36031 (n_14588, n21814);
  and g36032 (n21815, \asqrt[61] , n_14588);
  and g36036 (n21819, n_14107, n_14106);
  and g36037 (n21820, \asqrt[5] , n21819);
  not g36038 (n_14589, n21820);
  and g36039 (n21821, n_14105, n_14589);
  not g36040 (n_14590, n21818);
  not g36041 (n_14591, n21821);
  and g36042 (n21822, n_14590, n_14591);
  and g36043 (n21823, n_115, n_14586);
  and g36044 (n21824, n_14587, n21823);
  not g36045 (n_14592, n21822);
  not g36046 (n_14593, n21824);
  and g36047 (n21825, n_14592, n_14593);
  not g36048 (n_14594, n21815);
  not g36049 (n_14595, n21825);
  and g36050 (n21826, n_14594, n_14595);
  not g36051 (n_14596, n21826);
  and g36052 (n21827, \asqrt[62] , n_14596);
  and g36056 (n21831, n_14115, n_14114);
  and g36057 (n21832, \asqrt[5] , n21831);
  not g36058 (n_14597, n21832);
  and g36059 (n21833, n_14113, n_14597);
  not g36060 (n_14598, n21830);
  not g36061 (n_14599, n21833);
  and g36062 (n21834, n_14598, n_14599);
  and g36063 (n21835, n_76, n_14594);
  and g36064 (n21836, n_14595, n21835);
  not g36065 (n_14600, n21834);
  not g36066 (n_14601, n21836);
  and g36067 (n21837, n_14600, n_14601);
  not g36068 (n_14602, n21827);
  not g36069 (n_14603, n21837);
  and g36070 (n21838, n_14602, n_14603);
  and g36074 (n21842, n_14123, n_14122);
  and g36075 (n21843, \asqrt[5] , n21842);
  not g36076 (n_14604, n21843);
  and g36077 (n21844, n_14121, n_14604);
  not g36078 (n_14605, n21841);
  not g36079 (n_14606, n21844);
  and g36080 (n21845, n_14605, n_14606);
  and g36081 (n21846, n_14130, n_14129);
  and g36082 (n21847, \asqrt[5] , n21846);
  not g36085 (n_14608, n21845);
  not g36087 (n_14609, n21838);
  not g36089 (n_14610, n21850);
  and g36090 (n21851, n_21, n_14610);
  and g36091 (n21852, n_14602, n21845);
  and g36092 (n21853, n_14603, n21852);
  and g36093 (n21854, n_14129, \asqrt[5] );
  not g36094 (n_14611, n21854);
  and g36095 (n21855, n21129, n_14611);
  not g36096 (n_14612, n21846);
  and g36097 (n21856, \asqrt[63] , n_14612);
  not g36098 (n_14613, n21855);
  and g36099 (n21857, n_14613, n21856);
  not g36100 (n_14614, n21853);
  not g36101 (n_14615, n21857);
  and g36102 (n21858, n_14614, n_14615);
  not g36103 (n_14616, n21858);
  or g36104 (\asqrt[4] , n21851, n_14616);
  and g36105 (n21860, \a[8] , \asqrt[4] );
  not g36106 (n_14620, \a[6] );
  not g36107 (n_14621, \a[7] );
  and g36108 (n21861, n_14620, n_14621);
  and g36109 (n21862, n_14141, n21861);
  not g36110 (n_14622, n21860);
  not g36111 (n_14623, n21862);
  and g36112 (n21863, n_14622, n_14623);
  not g36113 (n_14624, n21863);
  and g36114 (n21864, \asqrt[5] , n_14624);
  and g36119 (n21869, n_14141, \asqrt[4] );
  not g36120 (n_14625, n21869);
  and g36121 (n21870, \a[9] , n_14625);
  and g36122 (n21871, n21152, \asqrt[4] );
  not g36123 (n_14626, n21870);
  not g36124 (n_14627, n21871);
  and g36125 (n21872, n_14626, n_14627);
  not g36126 (n_14628, n21868);
  and g36127 (n21873, n_14628, n21872);
  not g36128 (n_14629, n21864);
  not g36129 (n_14630, n21873);
  and g36130 (n21874, n_14629, n_14630);
  not g36131 (n_14631, n21874);
  and g36132 (n21875, \asqrt[6] , n_14631);
  not g36133 (n_14632, \asqrt[6] );
  and g36134 (n21876, n_14632, n_14629);
  and g36135 (n21877, n_14630, n21876);
  not g36138 (n_14633, n21851);
  not g36140 (n_14634, n21880);
  and g36141 (n21881, n_14627, n_14634);
  not g36142 (n_14635, n21881);
  and g36143 (n21882, \a[10] , n_14635);
  and g36144 (n21883, n_13670, n_14634);
  and g36145 (n21884, n_14627, n21883);
  not g36146 (n_14636, n21882);
  not g36147 (n_14637, n21884);
  and g36148 (n21885, n_14636, n_14637);
  not g36149 (n_14638, n21877);
  not g36150 (n_14639, n21885);
  and g36151 (n21886, n_14638, n_14639);
  not g36152 (n_14640, n21875);
  not g36153 (n_14641, n21886);
  and g36154 (n21887, n_14640, n_14641);
  not g36155 (n_14642, n21887);
  and g36156 (n21888, \asqrt[7] , n_14642);
  and g36157 (n21889, n_14150, n_14149);
  not g36158 (n_14643, n21164);
  and g36159 (n21890, n_14643, n21889);
  and g36160 (n21891, \asqrt[4] , n21890);
  and g36161 (n21892, \asqrt[4] , n21889);
  not g36162 (n_14644, n21892);
  and g36163 (n21893, n21164, n_14644);
  not g36164 (n_14645, n21891);
  not g36165 (n_14646, n21893);
  and g36166 (n21894, n_14645, n_14646);
  and g36167 (n21895, n_14153, n_14640);
  and g36168 (n21896, n_14641, n21895);
  not g36169 (n_14647, n21894);
  not g36170 (n_14648, n21896);
  and g36171 (n21897, n_14647, n_14648);
  not g36172 (n_14649, n21888);
  not g36173 (n_14650, n21897);
  and g36174 (n21898, n_14649, n_14650);
  not g36175 (n_14651, n21898);
  and g36176 (n21899, \asqrt[8] , n_14651);
  and g36180 (n21903, n_14161, n_14159);
  and g36181 (n21904, \asqrt[4] , n21903);
  not g36182 (n_14652, n21904);
  and g36183 (n21905, n_14160, n_14652);
  not g36184 (n_14653, n21902);
  not g36185 (n_14654, n21905);
  and g36186 (n21906, n_14653, n_14654);
  and g36187 (n21907, n_13682, n_14649);
  and g36188 (n21908, n_14650, n21907);
  not g36189 (n_14655, n21906);
  not g36190 (n_14656, n21908);
  and g36191 (n21909, n_14655, n_14656);
  not g36192 (n_14657, n21899);
  not g36193 (n_14658, n21909);
  and g36194 (n21910, n_14657, n_14658);
  not g36195 (n_14659, n21910);
  and g36196 (n21911, \asqrt[9] , n_14659);
  and g36200 (n21915, n_14170, n_14169);
  and g36201 (n21916, \asqrt[4] , n21915);
  not g36202 (n_14660, n21916);
  and g36203 (n21917, n_14168, n_14660);
  not g36204 (n_14661, n21914);
  not g36205 (n_14662, n21917);
  and g36206 (n21918, n_14661, n_14662);
  and g36207 (n21919, n_13218, n_14657);
  and g36208 (n21920, n_14658, n21919);
  not g36209 (n_14663, n21918);
  not g36210 (n_14664, n21920);
  and g36211 (n21921, n_14663, n_14664);
  not g36212 (n_14665, n21911);
  not g36213 (n_14666, n21921);
  and g36214 (n21922, n_14665, n_14666);
  not g36215 (n_14667, n21922);
  and g36216 (n21923, \asqrt[10] , n_14667);
  and g36220 (n21927, n_14178, n_14177);
  and g36221 (n21928, \asqrt[4] , n21927);
  not g36222 (n_14668, n21928);
  and g36223 (n21929, n_14176, n_14668);
  not g36224 (n_14669, n21926);
  not g36225 (n_14670, n21929);
  and g36226 (n21930, n_14669, n_14670);
  and g36227 (n21931, n_12762, n_14665);
  and g36228 (n21932, n_14666, n21931);
  not g36229 (n_14671, n21930);
  not g36230 (n_14672, n21932);
  and g36231 (n21933, n_14671, n_14672);
  not g36232 (n_14673, n21923);
  not g36233 (n_14674, n21933);
  and g36234 (n21934, n_14673, n_14674);
  not g36235 (n_14675, n21934);
  and g36236 (n21935, \asqrt[11] , n_14675);
  and g36240 (n21939, n_14186, n_14185);
  and g36241 (n21940, \asqrt[4] , n21939);
  not g36242 (n_14676, n21940);
  and g36243 (n21941, n_14184, n_14676);
  not g36244 (n_14677, n21938);
  not g36245 (n_14678, n21941);
  and g36246 (n21942, n_14677, n_14678);
  and g36247 (n21943, n_12314, n_14673);
  and g36248 (n21944, n_14674, n21943);
  not g36249 (n_14679, n21942);
  not g36250 (n_14680, n21944);
  and g36251 (n21945, n_14679, n_14680);
  not g36252 (n_14681, n21935);
  not g36253 (n_14682, n21945);
  and g36254 (n21946, n_14681, n_14682);
  not g36255 (n_14683, n21946);
  and g36256 (n21947, \asqrt[12] , n_14683);
  and g36260 (n21951, n_14194, n_14193);
  and g36261 (n21952, \asqrt[4] , n21951);
  not g36262 (n_14684, n21952);
  and g36263 (n21953, n_14192, n_14684);
  not g36264 (n_14685, n21950);
  not g36265 (n_14686, n21953);
  and g36266 (n21954, n_14685, n_14686);
  and g36267 (n21955, n_11874, n_14681);
  and g36268 (n21956, n_14682, n21955);
  not g36269 (n_14687, n21954);
  not g36270 (n_14688, n21956);
  and g36271 (n21957, n_14687, n_14688);
  not g36272 (n_14689, n21947);
  not g36273 (n_14690, n21957);
  and g36274 (n21958, n_14689, n_14690);
  not g36275 (n_14691, n21958);
  and g36276 (n21959, \asqrt[13] , n_14691);
  and g36280 (n21963, n_14202, n_14201);
  and g36281 (n21964, \asqrt[4] , n21963);
  not g36282 (n_14692, n21964);
  and g36283 (n21965, n_14200, n_14692);
  not g36284 (n_14693, n21962);
  not g36285 (n_14694, n21965);
  and g36286 (n21966, n_14693, n_14694);
  and g36287 (n21967, n_11442, n_14689);
  and g36288 (n21968, n_14690, n21967);
  not g36289 (n_14695, n21966);
  not g36290 (n_14696, n21968);
  and g36291 (n21969, n_14695, n_14696);
  not g36292 (n_14697, n21959);
  not g36293 (n_14698, n21969);
  and g36294 (n21970, n_14697, n_14698);
  not g36295 (n_14699, n21970);
  and g36296 (n21971, \asqrt[14] , n_14699);
  and g36300 (n21975, n_14210, n_14209);
  and g36301 (n21976, \asqrt[4] , n21975);
  not g36302 (n_14700, n21976);
  and g36303 (n21977, n_14208, n_14700);
  not g36304 (n_14701, n21974);
  not g36305 (n_14702, n21977);
  and g36306 (n21978, n_14701, n_14702);
  and g36307 (n21979, n_11018, n_14697);
  and g36308 (n21980, n_14698, n21979);
  not g36309 (n_14703, n21978);
  not g36310 (n_14704, n21980);
  and g36311 (n21981, n_14703, n_14704);
  not g36312 (n_14705, n21971);
  not g36313 (n_14706, n21981);
  and g36314 (n21982, n_14705, n_14706);
  not g36315 (n_14707, n21982);
  and g36316 (n21983, \asqrt[15] , n_14707);
  and g36320 (n21987, n_14218, n_14217);
  and g36321 (n21988, \asqrt[4] , n21987);
  not g36322 (n_14708, n21988);
  and g36323 (n21989, n_14216, n_14708);
  not g36324 (n_14709, n21986);
  not g36325 (n_14710, n21989);
  and g36326 (n21990, n_14709, n_14710);
  and g36327 (n21991, n_10602, n_14705);
  and g36328 (n21992, n_14706, n21991);
  not g36329 (n_14711, n21990);
  not g36330 (n_14712, n21992);
  and g36331 (n21993, n_14711, n_14712);
  not g36332 (n_14713, n21983);
  not g36333 (n_14714, n21993);
  and g36334 (n21994, n_14713, n_14714);
  not g36335 (n_14715, n21994);
  and g36336 (n21995, \asqrt[16] , n_14715);
  and g36340 (n21999, n_14226, n_14225);
  and g36341 (n22000, \asqrt[4] , n21999);
  not g36342 (n_14716, n22000);
  and g36343 (n22001, n_14224, n_14716);
  not g36344 (n_14717, n21998);
  not g36345 (n_14718, n22001);
  and g36346 (n22002, n_14717, n_14718);
  and g36347 (n22003, n_10194, n_14713);
  and g36348 (n22004, n_14714, n22003);
  not g36349 (n_14719, n22002);
  not g36350 (n_14720, n22004);
  and g36351 (n22005, n_14719, n_14720);
  not g36352 (n_14721, n21995);
  not g36353 (n_14722, n22005);
  and g36354 (n22006, n_14721, n_14722);
  not g36355 (n_14723, n22006);
  and g36356 (n22007, \asqrt[17] , n_14723);
  and g36360 (n22011, n_14234, n_14233);
  and g36361 (n22012, \asqrt[4] , n22011);
  not g36362 (n_14724, n22012);
  and g36363 (n22013, n_14232, n_14724);
  not g36364 (n_14725, n22010);
  not g36365 (n_14726, n22013);
  and g36366 (n22014, n_14725, n_14726);
  and g36367 (n22015, n_9794, n_14721);
  and g36368 (n22016, n_14722, n22015);
  not g36369 (n_14727, n22014);
  not g36370 (n_14728, n22016);
  and g36371 (n22017, n_14727, n_14728);
  not g36372 (n_14729, n22007);
  not g36373 (n_14730, n22017);
  and g36374 (n22018, n_14729, n_14730);
  not g36375 (n_14731, n22018);
  and g36376 (n22019, \asqrt[18] , n_14731);
  and g36380 (n22023, n_14242, n_14241);
  and g36381 (n22024, \asqrt[4] , n22023);
  not g36382 (n_14732, n22024);
  and g36383 (n22025, n_14240, n_14732);
  not g36384 (n_14733, n22022);
  not g36385 (n_14734, n22025);
  and g36386 (n22026, n_14733, n_14734);
  and g36387 (n22027, n_9402, n_14729);
  and g36388 (n22028, n_14730, n22027);
  not g36389 (n_14735, n22026);
  not g36390 (n_14736, n22028);
  and g36391 (n22029, n_14735, n_14736);
  not g36392 (n_14737, n22019);
  not g36393 (n_14738, n22029);
  and g36394 (n22030, n_14737, n_14738);
  not g36395 (n_14739, n22030);
  and g36396 (n22031, \asqrt[19] , n_14739);
  and g36400 (n22035, n_14250, n_14249);
  and g36401 (n22036, \asqrt[4] , n22035);
  not g36402 (n_14740, n22036);
  and g36403 (n22037, n_14248, n_14740);
  not g36404 (n_14741, n22034);
  not g36405 (n_14742, n22037);
  and g36406 (n22038, n_14741, n_14742);
  and g36407 (n22039, n_9018, n_14737);
  and g36408 (n22040, n_14738, n22039);
  not g36409 (n_14743, n22038);
  not g36410 (n_14744, n22040);
  and g36411 (n22041, n_14743, n_14744);
  not g36412 (n_14745, n22031);
  not g36413 (n_14746, n22041);
  and g36414 (n22042, n_14745, n_14746);
  not g36415 (n_14747, n22042);
  and g36416 (n22043, \asqrt[20] , n_14747);
  and g36420 (n22047, n_14258, n_14257);
  and g36421 (n22048, \asqrt[4] , n22047);
  not g36422 (n_14748, n22048);
  and g36423 (n22049, n_14256, n_14748);
  not g36424 (n_14749, n22046);
  not g36425 (n_14750, n22049);
  and g36426 (n22050, n_14749, n_14750);
  and g36427 (n22051, n_8642, n_14745);
  and g36428 (n22052, n_14746, n22051);
  not g36429 (n_14751, n22050);
  not g36430 (n_14752, n22052);
  and g36431 (n22053, n_14751, n_14752);
  not g36432 (n_14753, n22043);
  not g36433 (n_14754, n22053);
  and g36434 (n22054, n_14753, n_14754);
  not g36435 (n_14755, n22054);
  and g36436 (n22055, \asqrt[21] , n_14755);
  and g36440 (n22059, n_14266, n_14265);
  and g36441 (n22060, \asqrt[4] , n22059);
  not g36442 (n_14756, n22060);
  and g36443 (n22061, n_14264, n_14756);
  not g36444 (n_14757, n22058);
  not g36445 (n_14758, n22061);
  and g36446 (n22062, n_14757, n_14758);
  and g36447 (n22063, n_8274, n_14753);
  and g36448 (n22064, n_14754, n22063);
  not g36449 (n_14759, n22062);
  not g36450 (n_14760, n22064);
  and g36451 (n22065, n_14759, n_14760);
  not g36452 (n_14761, n22055);
  not g36453 (n_14762, n22065);
  and g36454 (n22066, n_14761, n_14762);
  not g36455 (n_14763, n22066);
  and g36456 (n22067, \asqrt[22] , n_14763);
  and g36460 (n22071, n_14274, n_14273);
  and g36461 (n22072, \asqrt[4] , n22071);
  not g36462 (n_14764, n22072);
  and g36463 (n22073, n_14272, n_14764);
  not g36464 (n_14765, n22070);
  not g36465 (n_14766, n22073);
  and g36466 (n22074, n_14765, n_14766);
  and g36467 (n22075, n_7914, n_14761);
  and g36468 (n22076, n_14762, n22075);
  not g36469 (n_14767, n22074);
  not g36470 (n_14768, n22076);
  and g36471 (n22077, n_14767, n_14768);
  not g36472 (n_14769, n22067);
  not g36473 (n_14770, n22077);
  and g36474 (n22078, n_14769, n_14770);
  not g36475 (n_14771, n22078);
  and g36476 (n22079, \asqrt[23] , n_14771);
  and g36480 (n22083, n_14282, n_14281);
  and g36481 (n22084, \asqrt[4] , n22083);
  not g36482 (n_14772, n22084);
  and g36483 (n22085, n_14280, n_14772);
  not g36484 (n_14773, n22082);
  not g36485 (n_14774, n22085);
  and g36486 (n22086, n_14773, n_14774);
  and g36487 (n22087, n_7562, n_14769);
  and g36488 (n22088, n_14770, n22087);
  not g36489 (n_14775, n22086);
  not g36490 (n_14776, n22088);
  and g36491 (n22089, n_14775, n_14776);
  not g36492 (n_14777, n22079);
  not g36493 (n_14778, n22089);
  and g36494 (n22090, n_14777, n_14778);
  not g36495 (n_14779, n22090);
  and g36496 (n22091, \asqrt[24] , n_14779);
  and g36500 (n22095, n_14290, n_14289);
  and g36501 (n22096, \asqrt[4] , n22095);
  not g36502 (n_14780, n22096);
  and g36503 (n22097, n_14288, n_14780);
  not g36504 (n_14781, n22094);
  not g36505 (n_14782, n22097);
  and g36506 (n22098, n_14781, n_14782);
  and g36507 (n22099, n_7218, n_14777);
  and g36508 (n22100, n_14778, n22099);
  not g36509 (n_14783, n22098);
  not g36510 (n_14784, n22100);
  and g36511 (n22101, n_14783, n_14784);
  not g36512 (n_14785, n22091);
  not g36513 (n_14786, n22101);
  and g36514 (n22102, n_14785, n_14786);
  not g36515 (n_14787, n22102);
  and g36516 (n22103, \asqrt[25] , n_14787);
  and g36520 (n22107, n_14298, n_14297);
  and g36521 (n22108, \asqrt[4] , n22107);
  not g36522 (n_14788, n22108);
  and g36523 (n22109, n_14296, n_14788);
  not g36524 (n_14789, n22106);
  not g36525 (n_14790, n22109);
  and g36526 (n22110, n_14789, n_14790);
  and g36527 (n22111, n_6882, n_14785);
  and g36528 (n22112, n_14786, n22111);
  not g36529 (n_14791, n22110);
  not g36530 (n_14792, n22112);
  and g36531 (n22113, n_14791, n_14792);
  not g36532 (n_14793, n22103);
  not g36533 (n_14794, n22113);
  and g36534 (n22114, n_14793, n_14794);
  not g36535 (n_14795, n22114);
  and g36536 (n22115, \asqrt[26] , n_14795);
  and g36540 (n22119, n_14306, n_14305);
  and g36541 (n22120, \asqrt[4] , n22119);
  not g36542 (n_14796, n22120);
  and g36543 (n22121, n_14304, n_14796);
  not g36544 (n_14797, n22118);
  not g36545 (n_14798, n22121);
  and g36546 (n22122, n_14797, n_14798);
  and g36547 (n22123, n_6554, n_14793);
  and g36548 (n22124, n_14794, n22123);
  not g36549 (n_14799, n22122);
  not g36550 (n_14800, n22124);
  and g36551 (n22125, n_14799, n_14800);
  not g36552 (n_14801, n22115);
  not g36553 (n_14802, n22125);
  and g36554 (n22126, n_14801, n_14802);
  not g36555 (n_14803, n22126);
  and g36556 (n22127, \asqrt[27] , n_14803);
  and g36560 (n22131, n_14314, n_14313);
  and g36561 (n22132, \asqrt[4] , n22131);
  not g36562 (n_14804, n22132);
  and g36563 (n22133, n_14312, n_14804);
  not g36564 (n_14805, n22130);
  not g36565 (n_14806, n22133);
  and g36566 (n22134, n_14805, n_14806);
  and g36567 (n22135, n_6234, n_14801);
  and g36568 (n22136, n_14802, n22135);
  not g36569 (n_14807, n22134);
  not g36570 (n_14808, n22136);
  and g36571 (n22137, n_14807, n_14808);
  not g36572 (n_14809, n22127);
  not g36573 (n_14810, n22137);
  and g36574 (n22138, n_14809, n_14810);
  not g36575 (n_14811, n22138);
  and g36576 (n22139, \asqrt[28] , n_14811);
  and g36580 (n22143, n_14322, n_14321);
  and g36581 (n22144, \asqrt[4] , n22143);
  not g36582 (n_14812, n22144);
  and g36583 (n22145, n_14320, n_14812);
  not g36584 (n_14813, n22142);
  not g36585 (n_14814, n22145);
  and g36586 (n22146, n_14813, n_14814);
  and g36587 (n22147, n_5922, n_14809);
  and g36588 (n22148, n_14810, n22147);
  not g36589 (n_14815, n22146);
  not g36590 (n_14816, n22148);
  and g36591 (n22149, n_14815, n_14816);
  not g36592 (n_14817, n22139);
  not g36593 (n_14818, n22149);
  and g36594 (n22150, n_14817, n_14818);
  not g36595 (n_14819, n22150);
  and g36596 (n22151, \asqrt[29] , n_14819);
  and g36600 (n22155, n_14330, n_14329);
  and g36601 (n22156, \asqrt[4] , n22155);
  not g36602 (n_14820, n22156);
  and g36603 (n22157, n_14328, n_14820);
  not g36604 (n_14821, n22154);
  not g36605 (n_14822, n22157);
  and g36606 (n22158, n_14821, n_14822);
  and g36607 (n22159, n_5618, n_14817);
  and g36608 (n22160, n_14818, n22159);
  not g36609 (n_14823, n22158);
  not g36610 (n_14824, n22160);
  and g36611 (n22161, n_14823, n_14824);
  not g36612 (n_14825, n22151);
  not g36613 (n_14826, n22161);
  and g36614 (n22162, n_14825, n_14826);
  not g36615 (n_14827, n22162);
  and g36616 (n22163, \asqrt[30] , n_14827);
  and g36620 (n22167, n_14338, n_14337);
  and g36621 (n22168, \asqrt[4] , n22167);
  not g36622 (n_14828, n22168);
  and g36623 (n22169, n_14336, n_14828);
  not g36624 (n_14829, n22166);
  not g36625 (n_14830, n22169);
  and g36626 (n22170, n_14829, n_14830);
  and g36627 (n22171, n_5322, n_14825);
  and g36628 (n22172, n_14826, n22171);
  not g36629 (n_14831, n22170);
  not g36630 (n_14832, n22172);
  and g36631 (n22173, n_14831, n_14832);
  not g36632 (n_14833, n22163);
  not g36633 (n_14834, n22173);
  and g36634 (n22174, n_14833, n_14834);
  not g36635 (n_14835, n22174);
  and g36636 (n22175, \asqrt[31] , n_14835);
  and g36640 (n22179, n_14346, n_14345);
  and g36641 (n22180, \asqrt[4] , n22179);
  not g36642 (n_14836, n22180);
  and g36643 (n22181, n_14344, n_14836);
  not g36644 (n_14837, n22178);
  not g36645 (n_14838, n22181);
  and g36646 (n22182, n_14837, n_14838);
  and g36647 (n22183, n_5034, n_14833);
  and g36648 (n22184, n_14834, n22183);
  not g36649 (n_14839, n22182);
  not g36650 (n_14840, n22184);
  and g36651 (n22185, n_14839, n_14840);
  not g36652 (n_14841, n22175);
  not g36653 (n_14842, n22185);
  and g36654 (n22186, n_14841, n_14842);
  not g36655 (n_14843, n22186);
  and g36656 (n22187, \asqrt[32] , n_14843);
  and g36660 (n22191, n_14354, n_14353);
  and g36661 (n22192, \asqrt[4] , n22191);
  not g36662 (n_14844, n22192);
  and g36663 (n22193, n_14352, n_14844);
  not g36664 (n_14845, n22190);
  not g36665 (n_14846, n22193);
  and g36666 (n22194, n_14845, n_14846);
  and g36667 (n22195, n_4754, n_14841);
  and g36668 (n22196, n_14842, n22195);
  not g36669 (n_14847, n22194);
  not g36670 (n_14848, n22196);
  and g36671 (n22197, n_14847, n_14848);
  not g36672 (n_14849, n22187);
  not g36673 (n_14850, n22197);
  and g36674 (n22198, n_14849, n_14850);
  not g36675 (n_14851, n22198);
  and g36676 (n22199, \asqrt[33] , n_14851);
  and g36680 (n22203, n_14362, n_14361);
  and g36681 (n22204, \asqrt[4] , n22203);
  not g36682 (n_14852, n22204);
  and g36683 (n22205, n_14360, n_14852);
  not g36684 (n_14853, n22202);
  not g36685 (n_14854, n22205);
  and g36686 (n22206, n_14853, n_14854);
  and g36687 (n22207, n_4482, n_14849);
  and g36688 (n22208, n_14850, n22207);
  not g36689 (n_14855, n22206);
  not g36690 (n_14856, n22208);
  and g36691 (n22209, n_14855, n_14856);
  not g36692 (n_14857, n22199);
  not g36693 (n_14858, n22209);
  and g36694 (n22210, n_14857, n_14858);
  not g36695 (n_14859, n22210);
  and g36696 (n22211, \asqrt[34] , n_14859);
  and g36700 (n22215, n_14370, n_14369);
  and g36701 (n22216, \asqrt[4] , n22215);
  not g36702 (n_14860, n22216);
  and g36703 (n22217, n_14368, n_14860);
  not g36704 (n_14861, n22214);
  not g36705 (n_14862, n22217);
  and g36706 (n22218, n_14861, n_14862);
  and g36707 (n22219, n_4218, n_14857);
  and g36708 (n22220, n_14858, n22219);
  not g36709 (n_14863, n22218);
  not g36710 (n_14864, n22220);
  and g36711 (n22221, n_14863, n_14864);
  not g36712 (n_14865, n22211);
  not g36713 (n_14866, n22221);
  and g36714 (n22222, n_14865, n_14866);
  not g36715 (n_14867, n22222);
  and g36716 (n22223, \asqrt[35] , n_14867);
  and g36720 (n22227, n_14378, n_14377);
  and g36721 (n22228, \asqrt[4] , n22227);
  not g36722 (n_14868, n22228);
  and g36723 (n22229, n_14376, n_14868);
  not g36724 (n_14869, n22226);
  not g36725 (n_14870, n22229);
  and g36726 (n22230, n_14869, n_14870);
  and g36727 (n22231, n_3962, n_14865);
  and g36728 (n22232, n_14866, n22231);
  not g36729 (n_14871, n22230);
  not g36730 (n_14872, n22232);
  and g36731 (n22233, n_14871, n_14872);
  not g36732 (n_14873, n22223);
  not g36733 (n_14874, n22233);
  and g36734 (n22234, n_14873, n_14874);
  not g36735 (n_14875, n22234);
  and g36736 (n22235, \asqrt[36] , n_14875);
  and g36740 (n22239, n_14386, n_14385);
  and g36741 (n22240, \asqrt[4] , n22239);
  not g36742 (n_14876, n22240);
  and g36743 (n22241, n_14384, n_14876);
  not g36744 (n_14877, n22238);
  not g36745 (n_14878, n22241);
  and g36746 (n22242, n_14877, n_14878);
  and g36747 (n22243, n_3714, n_14873);
  and g36748 (n22244, n_14874, n22243);
  not g36749 (n_14879, n22242);
  not g36750 (n_14880, n22244);
  and g36751 (n22245, n_14879, n_14880);
  not g36752 (n_14881, n22235);
  not g36753 (n_14882, n22245);
  and g36754 (n22246, n_14881, n_14882);
  not g36755 (n_14883, n22246);
  and g36756 (n22247, \asqrt[37] , n_14883);
  and g36760 (n22251, n_14394, n_14393);
  and g36761 (n22252, \asqrt[4] , n22251);
  not g36762 (n_14884, n22252);
  and g36763 (n22253, n_14392, n_14884);
  not g36764 (n_14885, n22250);
  not g36765 (n_14886, n22253);
  and g36766 (n22254, n_14885, n_14886);
  and g36767 (n22255, n_3474, n_14881);
  and g36768 (n22256, n_14882, n22255);
  not g36769 (n_14887, n22254);
  not g36770 (n_14888, n22256);
  and g36771 (n22257, n_14887, n_14888);
  not g36772 (n_14889, n22247);
  not g36773 (n_14890, n22257);
  and g36774 (n22258, n_14889, n_14890);
  not g36775 (n_14891, n22258);
  and g36776 (n22259, \asqrt[38] , n_14891);
  and g36780 (n22263, n_14402, n_14401);
  and g36781 (n22264, \asqrt[4] , n22263);
  not g36782 (n_14892, n22264);
  and g36783 (n22265, n_14400, n_14892);
  not g36784 (n_14893, n22262);
  not g36785 (n_14894, n22265);
  and g36786 (n22266, n_14893, n_14894);
  and g36787 (n22267, n_3242, n_14889);
  and g36788 (n22268, n_14890, n22267);
  not g36789 (n_14895, n22266);
  not g36790 (n_14896, n22268);
  and g36791 (n22269, n_14895, n_14896);
  not g36792 (n_14897, n22259);
  not g36793 (n_14898, n22269);
  and g36794 (n22270, n_14897, n_14898);
  not g36795 (n_14899, n22270);
  and g36796 (n22271, \asqrt[39] , n_14899);
  and g36800 (n22275, n_14410, n_14409);
  and g36801 (n22276, \asqrt[4] , n22275);
  not g36802 (n_14900, n22276);
  and g36803 (n22277, n_14408, n_14900);
  not g36804 (n_14901, n22274);
  not g36805 (n_14902, n22277);
  and g36806 (n22278, n_14901, n_14902);
  and g36807 (n22279, n_3018, n_14897);
  and g36808 (n22280, n_14898, n22279);
  not g36809 (n_14903, n22278);
  not g36810 (n_14904, n22280);
  and g36811 (n22281, n_14903, n_14904);
  not g36812 (n_14905, n22271);
  not g36813 (n_14906, n22281);
  and g36814 (n22282, n_14905, n_14906);
  not g36815 (n_14907, n22282);
  and g36816 (n22283, \asqrt[40] , n_14907);
  and g36820 (n22287, n_14418, n_14417);
  and g36821 (n22288, \asqrt[4] , n22287);
  not g36822 (n_14908, n22288);
  and g36823 (n22289, n_14416, n_14908);
  not g36824 (n_14909, n22286);
  not g36825 (n_14910, n22289);
  and g36826 (n22290, n_14909, n_14910);
  and g36827 (n22291, n_2802, n_14905);
  and g36828 (n22292, n_14906, n22291);
  not g36829 (n_14911, n22290);
  not g36830 (n_14912, n22292);
  and g36831 (n22293, n_14911, n_14912);
  not g36832 (n_14913, n22283);
  not g36833 (n_14914, n22293);
  and g36834 (n22294, n_14913, n_14914);
  not g36835 (n_14915, n22294);
  and g36836 (n22295, \asqrt[41] , n_14915);
  and g36840 (n22299, n_14426, n_14425);
  and g36841 (n22300, \asqrt[4] , n22299);
  not g36842 (n_14916, n22300);
  and g36843 (n22301, n_14424, n_14916);
  not g36844 (n_14917, n22298);
  not g36845 (n_14918, n22301);
  and g36846 (n22302, n_14917, n_14918);
  and g36847 (n22303, n_2594, n_14913);
  and g36848 (n22304, n_14914, n22303);
  not g36849 (n_14919, n22302);
  not g36850 (n_14920, n22304);
  and g36851 (n22305, n_14919, n_14920);
  not g36852 (n_14921, n22295);
  not g36853 (n_14922, n22305);
  and g36854 (n22306, n_14921, n_14922);
  not g36855 (n_14923, n22306);
  and g36856 (n22307, \asqrt[42] , n_14923);
  and g36860 (n22311, n_14434, n_14433);
  and g36861 (n22312, \asqrt[4] , n22311);
  not g36862 (n_14924, n22312);
  and g36863 (n22313, n_14432, n_14924);
  not g36864 (n_14925, n22310);
  not g36865 (n_14926, n22313);
  and g36866 (n22314, n_14925, n_14926);
  and g36867 (n22315, n_2394, n_14921);
  and g36868 (n22316, n_14922, n22315);
  not g36869 (n_14927, n22314);
  not g36870 (n_14928, n22316);
  and g36871 (n22317, n_14927, n_14928);
  not g36872 (n_14929, n22307);
  not g36873 (n_14930, n22317);
  and g36874 (n22318, n_14929, n_14930);
  not g36875 (n_14931, n22318);
  and g36876 (n22319, \asqrt[43] , n_14931);
  and g36880 (n22323, n_14442, n_14441);
  and g36881 (n22324, \asqrt[4] , n22323);
  not g36882 (n_14932, n22324);
  and g36883 (n22325, n_14440, n_14932);
  not g36884 (n_14933, n22322);
  not g36885 (n_14934, n22325);
  and g36886 (n22326, n_14933, n_14934);
  and g36887 (n22327, n_2202, n_14929);
  and g36888 (n22328, n_14930, n22327);
  not g36889 (n_14935, n22326);
  not g36890 (n_14936, n22328);
  and g36891 (n22329, n_14935, n_14936);
  not g36892 (n_14937, n22319);
  not g36893 (n_14938, n22329);
  and g36894 (n22330, n_14937, n_14938);
  not g36895 (n_14939, n22330);
  and g36896 (n22331, \asqrt[44] , n_14939);
  and g36900 (n22335, n_14450, n_14449);
  and g36901 (n22336, \asqrt[4] , n22335);
  not g36902 (n_14940, n22336);
  and g36903 (n22337, n_14448, n_14940);
  not g36904 (n_14941, n22334);
  not g36905 (n_14942, n22337);
  and g36906 (n22338, n_14941, n_14942);
  and g36907 (n22339, n_2018, n_14937);
  and g36908 (n22340, n_14938, n22339);
  not g36909 (n_14943, n22338);
  not g36910 (n_14944, n22340);
  and g36911 (n22341, n_14943, n_14944);
  not g36912 (n_14945, n22331);
  not g36913 (n_14946, n22341);
  and g36914 (n22342, n_14945, n_14946);
  not g36915 (n_14947, n22342);
  and g36916 (n22343, \asqrt[45] , n_14947);
  and g36920 (n22347, n_14458, n_14457);
  and g36921 (n22348, \asqrt[4] , n22347);
  not g36922 (n_14948, n22348);
  and g36923 (n22349, n_14456, n_14948);
  not g36924 (n_14949, n22346);
  not g36925 (n_14950, n22349);
  and g36926 (n22350, n_14949, n_14950);
  and g36927 (n22351, n_1842, n_14945);
  and g36928 (n22352, n_14946, n22351);
  not g36929 (n_14951, n22350);
  not g36930 (n_14952, n22352);
  and g36931 (n22353, n_14951, n_14952);
  not g36932 (n_14953, n22343);
  not g36933 (n_14954, n22353);
  and g36934 (n22354, n_14953, n_14954);
  not g36935 (n_14955, n22354);
  and g36936 (n22355, \asqrt[46] , n_14955);
  and g36940 (n22359, n_14466, n_14465);
  and g36941 (n22360, \asqrt[4] , n22359);
  not g36942 (n_14956, n22360);
  and g36943 (n22361, n_14464, n_14956);
  not g36944 (n_14957, n22358);
  not g36945 (n_14958, n22361);
  and g36946 (n22362, n_14957, n_14958);
  and g36947 (n22363, n_1674, n_14953);
  and g36948 (n22364, n_14954, n22363);
  not g36949 (n_14959, n22362);
  not g36950 (n_14960, n22364);
  and g36951 (n22365, n_14959, n_14960);
  not g36952 (n_14961, n22355);
  not g36953 (n_14962, n22365);
  and g36954 (n22366, n_14961, n_14962);
  not g36955 (n_14963, n22366);
  and g36956 (n22367, \asqrt[47] , n_14963);
  and g36960 (n22371, n_14474, n_14473);
  and g36961 (n22372, \asqrt[4] , n22371);
  not g36962 (n_14964, n22372);
  and g36963 (n22373, n_14472, n_14964);
  not g36964 (n_14965, n22370);
  not g36965 (n_14966, n22373);
  and g36966 (n22374, n_14965, n_14966);
  and g36967 (n22375, n_1514, n_14961);
  and g36968 (n22376, n_14962, n22375);
  not g36969 (n_14967, n22374);
  not g36970 (n_14968, n22376);
  and g36971 (n22377, n_14967, n_14968);
  not g36972 (n_14969, n22367);
  not g36973 (n_14970, n22377);
  and g36974 (n22378, n_14969, n_14970);
  not g36975 (n_14971, n22378);
  and g36976 (n22379, \asqrt[48] , n_14971);
  and g36980 (n22383, n_14482, n_14481);
  and g36981 (n22384, \asqrt[4] , n22383);
  not g36982 (n_14972, n22384);
  and g36983 (n22385, n_14480, n_14972);
  not g36984 (n_14973, n22382);
  not g36985 (n_14974, n22385);
  and g36986 (n22386, n_14973, n_14974);
  and g36987 (n22387, n_1362, n_14969);
  and g36988 (n22388, n_14970, n22387);
  not g36989 (n_14975, n22386);
  not g36990 (n_14976, n22388);
  and g36991 (n22389, n_14975, n_14976);
  not g36992 (n_14977, n22379);
  not g36993 (n_14978, n22389);
  and g36994 (n22390, n_14977, n_14978);
  not g36995 (n_14979, n22390);
  and g36996 (n22391, \asqrt[49] , n_14979);
  and g37000 (n22395, n_14490, n_14489);
  and g37001 (n22396, \asqrt[4] , n22395);
  not g37002 (n_14980, n22396);
  and g37003 (n22397, n_14488, n_14980);
  not g37004 (n_14981, n22394);
  not g37005 (n_14982, n22397);
  and g37006 (n22398, n_14981, n_14982);
  and g37007 (n22399, n_1218, n_14977);
  and g37008 (n22400, n_14978, n22399);
  not g37009 (n_14983, n22398);
  not g37010 (n_14984, n22400);
  and g37011 (n22401, n_14983, n_14984);
  not g37012 (n_14985, n22391);
  not g37013 (n_14986, n22401);
  and g37014 (n22402, n_14985, n_14986);
  not g37015 (n_14987, n22402);
  and g37016 (n22403, \asqrt[50] , n_14987);
  and g37020 (n22407, n_14498, n_14497);
  and g37021 (n22408, \asqrt[4] , n22407);
  not g37022 (n_14988, n22408);
  and g37023 (n22409, n_14496, n_14988);
  not g37024 (n_14989, n22406);
  not g37025 (n_14990, n22409);
  and g37026 (n22410, n_14989, n_14990);
  and g37027 (n22411, n_1082, n_14985);
  and g37028 (n22412, n_14986, n22411);
  not g37029 (n_14991, n22410);
  not g37030 (n_14992, n22412);
  and g37031 (n22413, n_14991, n_14992);
  not g37032 (n_14993, n22403);
  not g37033 (n_14994, n22413);
  and g37034 (n22414, n_14993, n_14994);
  not g37035 (n_14995, n22414);
  and g37036 (n22415, \asqrt[51] , n_14995);
  and g37040 (n22419, n_14506, n_14505);
  and g37041 (n22420, \asqrt[4] , n22419);
  not g37042 (n_14996, n22420);
  and g37043 (n22421, n_14504, n_14996);
  not g37044 (n_14997, n22418);
  not g37045 (n_14998, n22421);
  and g37046 (n22422, n_14997, n_14998);
  and g37047 (n22423, n_954, n_14993);
  and g37048 (n22424, n_14994, n22423);
  not g37049 (n_14999, n22422);
  not g37050 (n_15000, n22424);
  and g37051 (n22425, n_14999, n_15000);
  not g37052 (n_15001, n22415);
  not g37053 (n_15002, n22425);
  and g37054 (n22426, n_15001, n_15002);
  not g37055 (n_15003, n22426);
  and g37056 (n22427, \asqrt[52] , n_15003);
  and g37060 (n22431, n_14514, n_14513);
  and g37061 (n22432, \asqrt[4] , n22431);
  not g37062 (n_15004, n22432);
  and g37063 (n22433, n_14512, n_15004);
  not g37064 (n_15005, n22430);
  not g37065 (n_15006, n22433);
  and g37066 (n22434, n_15005, n_15006);
  and g37067 (n22435, n_834, n_15001);
  and g37068 (n22436, n_15002, n22435);
  not g37069 (n_15007, n22434);
  not g37070 (n_15008, n22436);
  and g37071 (n22437, n_15007, n_15008);
  not g37072 (n_15009, n22427);
  not g37073 (n_15010, n22437);
  and g37074 (n22438, n_15009, n_15010);
  not g37075 (n_15011, n22438);
  and g37076 (n22439, \asqrt[53] , n_15011);
  and g37080 (n22443, n_14522, n_14521);
  and g37081 (n22444, \asqrt[4] , n22443);
  not g37082 (n_15012, n22444);
  and g37083 (n22445, n_14520, n_15012);
  not g37084 (n_15013, n22442);
  not g37085 (n_15014, n22445);
  and g37086 (n22446, n_15013, n_15014);
  and g37087 (n22447, n_722, n_15009);
  and g37088 (n22448, n_15010, n22447);
  not g37089 (n_15015, n22446);
  not g37090 (n_15016, n22448);
  and g37091 (n22449, n_15015, n_15016);
  not g37092 (n_15017, n22439);
  not g37093 (n_15018, n22449);
  and g37094 (n22450, n_15017, n_15018);
  not g37095 (n_15019, n22450);
  and g37096 (n22451, \asqrt[54] , n_15019);
  and g37100 (n22455, n_14530, n_14529);
  and g37101 (n22456, \asqrt[4] , n22455);
  not g37102 (n_15020, n22456);
  and g37103 (n22457, n_14528, n_15020);
  not g37104 (n_15021, n22454);
  not g37105 (n_15022, n22457);
  and g37106 (n22458, n_15021, n_15022);
  and g37107 (n22459, n_618, n_15017);
  and g37108 (n22460, n_15018, n22459);
  not g37109 (n_15023, n22458);
  not g37110 (n_15024, n22460);
  and g37111 (n22461, n_15023, n_15024);
  not g37112 (n_15025, n22451);
  not g37113 (n_15026, n22461);
  and g37114 (n22462, n_15025, n_15026);
  not g37115 (n_15027, n22462);
  and g37116 (n22463, \asqrt[55] , n_15027);
  and g37120 (n22467, n_14538, n_14537);
  and g37121 (n22468, \asqrt[4] , n22467);
  not g37122 (n_15028, n22468);
  and g37123 (n22469, n_14536, n_15028);
  not g37124 (n_15029, n22466);
  not g37125 (n_15030, n22469);
  and g37126 (n22470, n_15029, n_15030);
  and g37127 (n22471, n_522, n_15025);
  and g37128 (n22472, n_15026, n22471);
  not g37129 (n_15031, n22470);
  not g37130 (n_15032, n22472);
  and g37131 (n22473, n_15031, n_15032);
  not g37132 (n_15033, n22463);
  not g37133 (n_15034, n22473);
  and g37134 (n22474, n_15033, n_15034);
  not g37135 (n_15035, n22474);
  and g37136 (n22475, \asqrt[56] , n_15035);
  and g37140 (n22479, n_14546, n_14545);
  and g37141 (n22480, \asqrt[4] , n22479);
  not g37142 (n_15036, n22480);
  and g37143 (n22481, n_14544, n_15036);
  not g37144 (n_15037, n22478);
  not g37145 (n_15038, n22481);
  and g37146 (n22482, n_15037, n_15038);
  and g37147 (n22483, n_434, n_15033);
  and g37148 (n22484, n_15034, n22483);
  not g37149 (n_15039, n22482);
  not g37150 (n_15040, n22484);
  and g37151 (n22485, n_15039, n_15040);
  not g37152 (n_15041, n22475);
  not g37153 (n_15042, n22485);
  and g37154 (n22486, n_15041, n_15042);
  not g37155 (n_15043, n22486);
  and g37156 (n22487, \asqrt[57] , n_15043);
  and g37160 (n22491, n_14554, n_14553);
  and g37161 (n22492, \asqrt[4] , n22491);
  not g37162 (n_15044, n22492);
  and g37163 (n22493, n_14552, n_15044);
  not g37164 (n_15045, n22490);
  not g37165 (n_15046, n22493);
  and g37166 (n22494, n_15045, n_15046);
  and g37167 (n22495, n_354, n_15041);
  and g37168 (n22496, n_15042, n22495);
  not g37169 (n_15047, n22494);
  not g37170 (n_15048, n22496);
  and g37171 (n22497, n_15047, n_15048);
  not g37172 (n_15049, n22487);
  not g37173 (n_15050, n22497);
  and g37174 (n22498, n_15049, n_15050);
  not g37175 (n_15051, n22498);
  and g37176 (n22499, \asqrt[58] , n_15051);
  and g37180 (n22503, n_14562, n_14561);
  and g37181 (n22504, \asqrt[4] , n22503);
  not g37182 (n_15052, n22504);
  and g37183 (n22505, n_14560, n_15052);
  not g37184 (n_15053, n22502);
  not g37185 (n_15054, n22505);
  and g37186 (n22506, n_15053, n_15054);
  and g37187 (n22507, n_282, n_15049);
  and g37188 (n22508, n_15050, n22507);
  not g37189 (n_15055, n22506);
  not g37190 (n_15056, n22508);
  and g37191 (n22509, n_15055, n_15056);
  not g37192 (n_15057, n22499);
  not g37193 (n_15058, n22509);
  and g37194 (n22510, n_15057, n_15058);
  not g37195 (n_15059, n22510);
  and g37196 (n22511, \asqrt[59] , n_15059);
  and g37200 (n22515, n_14570, n_14569);
  and g37201 (n22516, \asqrt[4] , n22515);
  not g37202 (n_15060, n22516);
  and g37203 (n22517, n_14568, n_15060);
  not g37204 (n_15061, n22514);
  not g37205 (n_15062, n22517);
  and g37206 (n22518, n_15061, n_15062);
  and g37207 (n22519, n_218, n_15057);
  and g37208 (n22520, n_15058, n22519);
  not g37209 (n_15063, n22518);
  not g37210 (n_15064, n22520);
  and g37211 (n22521, n_15063, n_15064);
  not g37212 (n_15065, n22511);
  not g37213 (n_15066, n22521);
  and g37214 (n22522, n_15065, n_15066);
  not g37215 (n_15067, n22522);
  and g37216 (n22523, \asqrt[60] , n_15067);
  and g37220 (n22527, n_14578, n_14577);
  and g37221 (n22528, \asqrt[4] , n22527);
  not g37222 (n_15068, n22528);
  and g37223 (n22529, n_14576, n_15068);
  not g37224 (n_15069, n22526);
  not g37225 (n_15070, n22529);
  and g37226 (n22530, n_15069, n_15070);
  and g37227 (n22531, n_162, n_15065);
  and g37228 (n22532, n_15066, n22531);
  not g37229 (n_15071, n22530);
  not g37230 (n_15072, n22532);
  and g37231 (n22533, n_15071, n_15072);
  not g37232 (n_15073, n22523);
  not g37233 (n_15074, n22533);
  and g37234 (n22534, n_15073, n_15074);
  not g37235 (n_15075, n22534);
  and g37236 (n22535, \asqrt[61] , n_15075);
  and g37237 (n22536, n_115, n_15073);
  and g37238 (n22537, n_15074, n22536);
  and g37242 (n22541, n_14586, n_14584);
  and g37243 (n22542, \asqrt[4] , n22541);
  not g37244 (n_15076, n22542);
  and g37245 (n22543, n_14585, n_15076);
  not g37246 (n_15077, n22540);
  not g37247 (n_15078, n22543);
  and g37248 (n22544, n_15077, n_15078);
  not g37249 (n_15079, n22537);
  not g37250 (n_15080, n22544);
  and g37251 (n22545, n_15079, n_15080);
  not g37252 (n_15081, n22535);
  not g37253 (n_15082, n22545);
  and g37254 (n22546, n_15081, n_15082);
  not g37255 (n_15083, n22546);
  and g37256 (n22547, \asqrt[62] , n_15083);
  and g37260 (n22551, n_14594, n_14593);
  and g37261 (n22552, \asqrt[4] , n22551);
  not g37262 (n_15084, n22552);
  and g37263 (n22553, n_14592, n_15084);
  not g37264 (n_15085, n22550);
  not g37265 (n_15086, n22553);
  and g37266 (n22554, n_15085, n_15086);
  and g37267 (n22555, n_76, n_15081);
  and g37268 (n22556, n_15082, n22555);
  not g37269 (n_15087, n22554);
  not g37270 (n_15088, n22556);
  and g37271 (n22557, n_15087, n_15088);
  not g37272 (n_15089, n22547);
  not g37273 (n_15090, n22557);
  and g37274 (n22558, n_15089, n_15090);
  and g37278 (n22562, n_14602, n_14601);
  and g37279 (n22563, \asqrt[4] , n22562);
  not g37280 (n_15091, n22563);
  and g37281 (n22564, n_14600, n_15091);
  not g37282 (n_15092, n22561);
  not g37283 (n_15093, n22564);
  and g37284 (n22565, n_15092, n_15093);
  and g37285 (n22566, n_14609, n_14608);
  and g37286 (n22567, \asqrt[4] , n22566);
  not g37289 (n_15095, n22565);
  not g37291 (n_15096, n22558);
  not g37293 (n_15097, n22570);
  and g37294 (n22571, n_21, n_15097);
  and g37295 (n22572, n_15089, n22565);
  and g37296 (n22573, n_15090, n22572);
  and g37297 (n22574, n_14608, \asqrt[4] );
  not g37298 (n_15098, n22574);
  and g37299 (n22575, n21838, n_15098);
  not g37300 (n_15099, n22566);
  and g37301 (n22576, \asqrt[63] , n_15099);
  not g37302 (n_15100, n22575);
  and g37303 (n22577, n_15100, n22576);
  not g37304 (n_15101, n22573);
  not g37305 (n_15102, n22577);
  and g37306 (n22578, n_15101, n_15102);
  not g37307 (n_15103, n22578);
  or g37308 (\asqrt[3] , n22571, n_15103);
  and g37309 (n22580, \a[6] , \asqrt[3] );
  not g37310 (n_15107, \a[4] );
  not g37311 (n_15108, \a[5] );
  and g37312 (n22581, n_15107, n_15108);
  and g37313 (n22582, n_14620, n22581);
  not g37314 (n_15109, n22580);
  not g37315 (n_15110, n22582);
  and g37316 (n22583, n_15109, n_15110);
  not g37317 (n_15111, n22583);
  and g37318 (n22584, \asqrt[4] , n_15111);
  and g37323 (n22589, n_14620, \asqrt[3] );
  not g37324 (n_15112, n22589);
  and g37325 (n22590, \a[7] , n_15112);
  and g37326 (n22591, n21861, \asqrt[3] );
  not g37327 (n_15113, n22590);
  not g37328 (n_15114, n22591);
  and g37329 (n22592, n_15113, n_15114);
  not g37330 (n_15115, n22588);
  and g37331 (n22593, n_15115, n22592);
  not g37332 (n_15116, n22584);
  not g37333 (n_15117, n22593);
  and g37334 (n22594, n_15116, n_15117);
  not g37335 (n_15118, n22594);
  and g37336 (n22595, \asqrt[5] , n_15118);
  not g37337 (n_15119, \asqrt[5] );
  and g37338 (n22596, n_15119, n_15116);
  and g37339 (n22597, n_15117, n22596);
  not g37342 (n_15120, n22571);
  not g37344 (n_15121, n22600);
  and g37345 (n22601, n_15114, n_15121);
  not g37346 (n_15122, n22601);
  and g37347 (n22602, \a[8] , n_15122);
  and g37348 (n22603, n_14141, n_15121);
  and g37349 (n22604, n_15114, n22603);
  not g37350 (n_15123, n22602);
  not g37351 (n_15124, n22604);
  and g37352 (n22605, n_15123, n_15124);
  not g37353 (n_15125, n22597);
  not g37354 (n_15126, n22605);
  and g37355 (n22606, n_15125, n_15126);
  not g37356 (n_15127, n22595);
  not g37357 (n_15128, n22606);
  and g37358 (n22607, n_15127, n_15128);
  not g37359 (n_15129, n22607);
  and g37360 (n22608, \asqrt[6] , n_15129);
  and g37361 (n22609, n_14629, n_14628);
  not g37362 (n_15130, n21872);
  and g37363 (n22610, n_15130, n22609);
  and g37364 (n22611, \asqrt[3] , n22610);
  and g37365 (n22612, \asqrt[3] , n22609);
  not g37366 (n_15131, n22612);
  and g37367 (n22613, n21872, n_15131);
  not g37368 (n_15132, n22611);
  not g37369 (n_15133, n22613);
  and g37370 (n22614, n_15132, n_15133);
  and g37371 (n22615, n_14632, n_15127);
  and g37372 (n22616, n_15128, n22615);
  not g37373 (n_15134, n22614);
  not g37374 (n_15135, n22616);
  and g37375 (n22617, n_15134, n_15135);
  not g37376 (n_15136, n22608);
  not g37377 (n_15137, n22617);
  and g37378 (n22618, n_15136, n_15137);
  not g37379 (n_15138, n22618);
  and g37380 (n22619, \asqrt[7] , n_15138);
  and g37384 (n22623, n_14640, n_14638);
  and g37385 (n22624, \asqrt[3] , n22623);
  not g37386 (n_15139, n22624);
  and g37387 (n22625, n_14639, n_15139);
  not g37388 (n_15140, n22622);
  not g37389 (n_15141, n22625);
  and g37390 (n22626, n_15140, n_15141);
  and g37391 (n22627, n_14153, n_15136);
  and g37392 (n22628, n_15137, n22627);
  not g37393 (n_15142, n22626);
  not g37394 (n_15143, n22628);
  and g37395 (n22629, n_15142, n_15143);
  not g37396 (n_15144, n22619);
  not g37397 (n_15145, n22629);
  and g37398 (n22630, n_15144, n_15145);
  not g37399 (n_15146, n22630);
  and g37400 (n22631, \asqrt[8] , n_15146);
  and g37404 (n22635, n_14649, n_14648);
  and g37405 (n22636, \asqrt[3] , n22635);
  not g37406 (n_15147, n22636);
  and g37407 (n22637, n_14647, n_15147);
  not g37408 (n_15148, n22634);
  not g37409 (n_15149, n22637);
  and g37410 (n22638, n_15148, n_15149);
  and g37411 (n22639, n_13682, n_15144);
  and g37412 (n22640, n_15145, n22639);
  not g37413 (n_15150, n22638);
  not g37414 (n_15151, n22640);
  and g37415 (n22641, n_15150, n_15151);
  not g37416 (n_15152, n22631);
  not g37417 (n_15153, n22641);
  and g37418 (n22642, n_15152, n_15153);
  not g37419 (n_15154, n22642);
  and g37420 (n22643, \asqrt[9] , n_15154);
  and g37424 (n22647, n_14657, n_14656);
  and g37425 (n22648, \asqrt[3] , n22647);
  not g37426 (n_15155, n22648);
  and g37427 (n22649, n_14655, n_15155);
  not g37428 (n_15156, n22646);
  not g37429 (n_15157, n22649);
  and g37430 (n22650, n_15156, n_15157);
  and g37431 (n22651, n_13218, n_15152);
  and g37432 (n22652, n_15153, n22651);
  not g37433 (n_15158, n22650);
  not g37434 (n_15159, n22652);
  and g37435 (n22653, n_15158, n_15159);
  not g37436 (n_15160, n22643);
  not g37437 (n_15161, n22653);
  and g37438 (n22654, n_15160, n_15161);
  not g37439 (n_15162, n22654);
  and g37440 (n22655, \asqrt[10] , n_15162);
  and g37444 (n22659, n_14665, n_14664);
  and g37445 (n22660, \asqrt[3] , n22659);
  not g37446 (n_15163, n22660);
  and g37447 (n22661, n_14663, n_15163);
  not g37448 (n_15164, n22658);
  not g37449 (n_15165, n22661);
  and g37450 (n22662, n_15164, n_15165);
  and g37451 (n22663, n_12762, n_15160);
  and g37452 (n22664, n_15161, n22663);
  not g37453 (n_15166, n22662);
  not g37454 (n_15167, n22664);
  and g37455 (n22665, n_15166, n_15167);
  not g37456 (n_15168, n22655);
  not g37457 (n_15169, n22665);
  and g37458 (n22666, n_15168, n_15169);
  not g37459 (n_15170, n22666);
  and g37460 (n22667, \asqrt[11] , n_15170);
  and g37464 (n22671, n_14673, n_14672);
  and g37465 (n22672, \asqrt[3] , n22671);
  not g37466 (n_15171, n22672);
  and g37467 (n22673, n_14671, n_15171);
  not g37468 (n_15172, n22670);
  not g37469 (n_15173, n22673);
  and g37470 (n22674, n_15172, n_15173);
  and g37471 (n22675, n_12314, n_15168);
  and g37472 (n22676, n_15169, n22675);
  not g37473 (n_15174, n22674);
  not g37474 (n_15175, n22676);
  and g37475 (n22677, n_15174, n_15175);
  not g37476 (n_15176, n22667);
  not g37477 (n_15177, n22677);
  and g37478 (n22678, n_15176, n_15177);
  not g37479 (n_15178, n22678);
  and g37480 (n22679, \asqrt[12] , n_15178);
  and g37484 (n22683, n_14681, n_14680);
  and g37485 (n22684, \asqrt[3] , n22683);
  not g37486 (n_15179, n22684);
  and g37487 (n22685, n_14679, n_15179);
  not g37488 (n_15180, n22682);
  not g37489 (n_15181, n22685);
  and g37490 (n22686, n_15180, n_15181);
  and g37491 (n22687, n_11874, n_15176);
  and g37492 (n22688, n_15177, n22687);
  not g37493 (n_15182, n22686);
  not g37494 (n_15183, n22688);
  and g37495 (n22689, n_15182, n_15183);
  not g37496 (n_15184, n22679);
  not g37497 (n_15185, n22689);
  and g37498 (n22690, n_15184, n_15185);
  not g37499 (n_15186, n22690);
  and g37500 (n22691, \asqrt[13] , n_15186);
  and g37504 (n22695, n_14689, n_14688);
  and g37505 (n22696, \asqrt[3] , n22695);
  not g37506 (n_15187, n22696);
  and g37507 (n22697, n_14687, n_15187);
  not g37508 (n_15188, n22694);
  not g37509 (n_15189, n22697);
  and g37510 (n22698, n_15188, n_15189);
  and g37511 (n22699, n_11442, n_15184);
  and g37512 (n22700, n_15185, n22699);
  not g37513 (n_15190, n22698);
  not g37514 (n_15191, n22700);
  and g37515 (n22701, n_15190, n_15191);
  not g37516 (n_15192, n22691);
  not g37517 (n_15193, n22701);
  and g37518 (n22702, n_15192, n_15193);
  not g37519 (n_15194, n22702);
  and g37520 (n22703, \asqrt[14] , n_15194);
  and g37524 (n22707, n_14697, n_14696);
  and g37525 (n22708, \asqrt[3] , n22707);
  not g37526 (n_15195, n22708);
  and g37527 (n22709, n_14695, n_15195);
  not g37528 (n_15196, n22706);
  not g37529 (n_15197, n22709);
  and g37530 (n22710, n_15196, n_15197);
  and g37531 (n22711, n_11018, n_15192);
  and g37532 (n22712, n_15193, n22711);
  not g37533 (n_15198, n22710);
  not g37534 (n_15199, n22712);
  and g37535 (n22713, n_15198, n_15199);
  not g37536 (n_15200, n22703);
  not g37537 (n_15201, n22713);
  and g37538 (n22714, n_15200, n_15201);
  not g37539 (n_15202, n22714);
  and g37540 (n22715, \asqrt[15] , n_15202);
  and g37544 (n22719, n_14705, n_14704);
  and g37545 (n22720, \asqrt[3] , n22719);
  not g37546 (n_15203, n22720);
  and g37547 (n22721, n_14703, n_15203);
  not g37548 (n_15204, n22718);
  not g37549 (n_15205, n22721);
  and g37550 (n22722, n_15204, n_15205);
  and g37551 (n22723, n_10602, n_15200);
  and g37552 (n22724, n_15201, n22723);
  not g37553 (n_15206, n22722);
  not g37554 (n_15207, n22724);
  and g37555 (n22725, n_15206, n_15207);
  not g37556 (n_15208, n22715);
  not g37557 (n_15209, n22725);
  and g37558 (n22726, n_15208, n_15209);
  not g37559 (n_15210, n22726);
  and g37560 (n22727, \asqrt[16] , n_15210);
  and g37564 (n22731, n_14713, n_14712);
  and g37565 (n22732, \asqrt[3] , n22731);
  not g37566 (n_15211, n22732);
  and g37567 (n22733, n_14711, n_15211);
  not g37568 (n_15212, n22730);
  not g37569 (n_15213, n22733);
  and g37570 (n22734, n_15212, n_15213);
  and g37571 (n22735, n_10194, n_15208);
  and g37572 (n22736, n_15209, n22735);
  not g37573 (n_15214, n22734);
  not g37574 (n_15215, n22736);
  and g37575 (n22737, n_15214, n_15215);
  not g37576 (n_15216, n22727);
  not g37577 (n_15217, n22737);
  and g37578 (n22738, n_15216, n_15217);
  not g37579 (n_15218, n22738);
  and g37580 (n22739, \asqrt[17] , n_15218);
  and g37584 (n22743, n_14721, n_14720);
  and g37585 (n22744, \asqrt[3] , n22743);
  not g37586 (n_15219, n22744);
  and g37587 (n22745, n_14719, n_15219);
  not g37588 (n_15220, n22742);
  not g37589 (n_15221, n22745);
  and g37590 (n22746, n_15220, n_15221);
  and g37591 (n22747, n_9794, n_15216);
  and g37592 (n22748, n_15217, n22747);
  not g37593 (n_15222, n22746);
  not g37594 (n_15223, n22748);
  and g37595 (n22749, n_15222, n_15223);
  not g37596 (n_15224, n22739);
  not g37597 (n_15225, n22749);
  and g37598 (n22750, n_15224, n_15225);
  not g37599 (n_15226, n22750);
  and g37600 (n22751, \asqrt[18] , n_15226);
  and g37604 (n22755, n_14729, n_14728);
  and g37605 (n22756, \asqrt[3] , n22755);
  not g37606 (n_15227, n22756);
  and g37607 (n22757, n_14727, n_15227);
  not g37608 (n_15228, n22754);
  not g37609 (n_15229, n22757);
  and g37610 (n22758, n_15228, n_15229);
  and g37611 (n22759, n_9402, n_15224);
  and g37612 (n22760, n_15225, n22759);
  not g37613 (n_15230, n22758);
  not g37614 (n_15231, n22760);
  and g37615 (n22761, n_15230, n_15231);
  not g37616 (n_15232, n22751);
  not g37617 (n_15233, n22761);
  and g37618 (n22762, n_15232, n_15233);
  not g37619 (n_15234, n22762);
  and g37620 (n22763, \asqrt[19] , n_15234);
  and g37624 (n22767, n_14737, n_14736);
  and g37625 (n22768, \asqrt[3] , n22767);
  not g37626 (n_15235, n22768);
  and g37627 (n22769, n_14735, n_15235);
  not g37628 (n_15236, n22766);
  not g37629 (n_15237, n22769);
  and g37630 (n22770, n_15236, n_15237);
  and g37631 (n22771, n_9018, n_15232);
  and g37632 (n22772, n_15233, n22771);
  not g37633 (n_15238, n22770);
  not g37634 (n_15239, n22772);
  and g37635 (n22773, n_15238, n_15239);
  not g37636 (n_15240, n22763);
  not g37637 (n_15241, n22773);
  and g37638 (n22774, n_15240, n_15241);
  not g37639 (n_15242, n22774);
  and g37640 (n22775, \asqrt[20] , n_15242);
  and g37644 (n22779, n_14745, n_14744);
  and g37645 (n22780, \asqrt[3] , n22779);
  not g37646 (n_15243, n22780);
  and g37647 (n22781, n_14743, n_15243);
  not g37648 (n_15244, n22778);
  not g37649 (n_15245, n22781);
  and g37650 (n22782, n_15244, n_15245);
  and g37651 (n22783, n_8642, n_15240);
  and g37652 (n22784, n_15241, n22783);
  not g37653 (n_15246, n22782);
  not g37654 (n_15247, n22784);
  and g37655 (n22785, n_15246, n_15247);
  not g37656 (n_15248, n22775);
  not g37657 (n_15249, n22785);
  and g37658 (n22786, n_15248, n_15249);
  not g37659 (n_15250, n22786);
  and g37660 (n22787, \asqrt[21] , n_15250);
  and g37664 (n22791, n_14753, n_14752);
  and g37665 (n22792, \asqrt[3] , n22791);
  not g37666 (n_15251, n22792);
  and g37667 (n22793, n_14751, n_15251);
  not g37668 (n_15252, n22790);
  not g37669 (n_15253, n22793);
  and g37670 (n22794, n_15252, n_15253);
  and g37671 (n22795, n_8274, n_15248);
  and g37672 (n22796, n_15249, n22795);
  not g37673 (n_15254, n22794);
  not g37674 (n_15255, n22796);
  and g37675 (n22797, n_15254, n_15255);
  not g37676 (n_15256, n22787);
  not g37677 (n_15257, n22797);
  and g37678 (n22798, n_15256, n_15257);
  not g37679 (n_15258, n22798);
  and g37680 (n22799, \asqrt[22] , n_15258);
  and g37684 (n22803, n_14761, n_14760);
  and g37685 (n22804, \asqrt[3] , n22803);
  not g37686 (n_15259, n22804);
  and g37687 (n22805, n_14759, n_15259);
  not g37688 (n_15260, n22802);
  not g37689 (n_15261, n22805);
  and g37690 (n22806, n_15260, n_15261);
  and g37691 (n22807, n_7914, n_15256);
  and g37692 (n22808, n_15257, n22807);
  not g37693 (n_15262, n22806);
  not g37694 (n_15263, n22808);
  and g37695 (n22809, n_15262, n_15263);
  not g37696 (n_15264, n22799);
  not g37697 (n_15265, n22809);
  and g37698 (n22810, n_15264, n_15265);
  not g37699 (n_15266, n22810);
  and g37700 (n22811, \asqrt[23] , n_15266);
  and g37704 (n22815, n_14769, n_14768);
  and g37705 (n22816, \asqrt[3] , n22815);
  not g37706 (n_15267, n22816);
  and g37707 (n22817, n_14767, n_15267);
  not g37708 (n_15268, n22814);
  not g37709 (n_15269, n22817);
  and g37710 (n22818, n_15268, n_15269);
  and g37711 (n22819, n_7562, n_15264);
  and g37712 (n22820, n_15265, n22819);
  not g37713 (n_15270, n22818);
  not g37714 (n_15271, n22820);
  and g37715 (n22821, n_15270, n_15271);
  not g37716 (n_15272, n22811);
  not g37717 (n_15273, n22821);
  and g37718 (n22822, n_15272, n_15273);
  not g37719 (n_15274, n22822);
  and g37720 (n22823, \asqrt[24] , n_15274);
  and g37724 (n22827, n_14777, n_14776);
  and g37725 (n22828, \asqrt[3] , n22827);
  not g37726 (n_15275, n22828);
  and g37727 (n22829, n_14775, n_15275);
  not g37728 (n_15276, n22826);
  not g37729 (n_15277, n22829);
  and g37730 (n22830, n_15276, n_15277);
  and g37731 (n22831, n_7218, n_15272);
  and g37732 (n22832, n_15273, n22831);
  not g37733 (n_15278, n22830);
  not g37734 (n_15279, n22832);
  and g37735 (n22833, n_15278, n_15279);
  not g37736 (n_15280, n22823);
  not g37737 (n_15281, n22833);
  and g37738 (n22834, n_15280, n_15281);
  not g37739 (n_15282, n22834);
  and g37740 (n22835, \asqrt[25] , n_15282);
  and g37744 (n22839, n_14785, n_14784);
  and g37745 (n22840, \asqrt[3] , n22839);
  not g37746 (n_15283, n22840);
  and g37747 (n22841, n_14783, n_15283);
  not g37748 (n_15284, n22838);
  not g37749 (n_15285, n22841);
  and g37750 (n22842, n_15284, n_15285);
  and g37751 (n22843, n_6882, n_15280);
  and g37752 (n22844, n_15281, n22843);
  not g37753 (n_15286, n22842);
  not g37754 (n_15287, n22844);
  and g37755 (n22845, n_15286, n_15287);
  not g37756 (n_15288, n22835);
  not g37757 (n_15289, n22845);
  and g37758 (n22846, n_15288, n_15289);
  not g37759 (n_15290, n22846);
  and g37760 (n22847, \asqrt[26] , n_15290);
  and g37764 (n22851, n_14793, n_14792);
  and g37765 (n22852, \asqrt[3] , n22851);
  not g37766 (n_15291, n22852);
  and g37767 (n22853, n_14791, n_15291);
  not g37768 (n_15292, n22850);
  not g37769 (n_15293, n22853);
  and g37770 (n22854, n_15292, n_15293);
  and g37771 (n22855, n_6554, n_15288);
  and g37772 (n22856, n_15289, n22855);
  not g37773 (n_15294, n22854);
  not g37774 (n_15295, n22856);
  and g37775 (n22857, n_15294, n_15295);
  not g37776 (n_15296, n22847);
  not g37777 (n_15297, n22857);
  and g37778 (n22858, n_15296, n_15297);
  not g37779 (n_15298, n22858);
  and g37780 (n22859, \asqrt[27] , n_15298);
  and g37784 (n22863, n_14801, n_14800);
  and g37785 (n22864, \asqrt[3] , n22863);
  not g37786 (n_15299, n22864);
  and g37787 (n22865, n_14799, n_15299);
  not g37788 (n_15300, n22862);
  not g37789 (n_15301, n22865);
  and g37790 (n22866, n_15300, n_15301);
  and g37791 (n22867, n_6234, n_15296);
  and g37792 (n22868, n_15297, n22867);
  not g37793 (n_15302, n22866);
  not g37794 (n_15303, n22868);
  and g37795 (n22869, n_15302, n_15303);
  not g37796 (n_15304, n22859);
  not g37797 (n_15305, n22869);
  and g37798 (n22870, n_15304, n_15305);
  not g37799 (n_15306, n22870);
  and g37800 (n22871, \asqrt[28] , n_15306);
  and g37804 (n22875, n_14809, n_14808);
  and g37805 (n22876, \asqrt[3] , n22875);
  not g37806 (n_15307, n22876);
  and g37807 (n22877, n_14807, n_15307);
  not g37808 (n_15308, n22874);
  not g37809 (n_15309, n22877);
  and g37810 (n22878, n_15308, n_15309);
  and g37811 (n22879, n_5922, n_15304);
  and g37812 (n22880, n_15305, n22879);
  not g37813 (n_15310, n22878);
  not g37814 (n_15311, n22880);
  and g37815 (n22881, n_15310, n_15311);
  not g37816 (n_15312, n22871);
  not g37817 (n_15313, n22881);
  and g37818 (n22882, n_15312, n_15313);
  not g37819 (n_15314, n22882);
  and g37820 (n22883, \asqrt[29] , n_15314);
  and g37824 (n22887, n_14817, n_14816);
  and g37825 (n22888, \asqrt[3] , n22887);
  not g37826 (n_15315, n22888);
  and g37827 (n22889, n_14815, n_15315);
  not g37828 (n_15316, n22886);
  not g37829 (n_15317, n22889);
  and g37830 (n22890, n_15316, n_15317);
  and g37831 (n22891, n_5618, n_15312);
  and g37832 (n22892, n_15313, n22891);
  not g37833 (n_15318, n22890);
  not g37834 (n_15319, n22892);
  and g37835 (n22893, n_15318, n_15319);
  not g37836 (n_15320, n22883);
  not g37837 (n_15321, n22893);
  and g37838 (n22894, n_15320, n_15321);
  not g37839 (n_15322, n22894);
  and g37840 (n22895, \asqrt[30] , n_15322);
  and g37844 (n22899, n_14825, n_14824);
  and g37845 (n22900, \asqrt[3] , n22899);
  not g37846 (n_15323, n22900);
  and g37847 (n22901, n_14823, n_15323);
  not g37848 (n_15324, n22898);
  not g37849 (n_15325, n22901);
  and g37850 (n22902, n_15324, n_15325);
  and g37851 (n22903, n_5322, n_15320);
  and g37852 (n22904, n_15321, n22903);
  not g37853 (n_15326, n22902);
  not g37854 (n_15327, n22904);
  and g37855 (n22905, n_15326, n_15327);
  not g37856 (n_15328, n22895);
  not g37857 (n_15329, n22905);
  and g37858 (n22906, n_15328, n_15329);
  not g37859 (n_15330, n22906);
  and g37860 (n22907, \asqrt[31] , n_15330);
  and g37864 (n22911, n_14833, n_14832);
  and g37865 (n22912, \asqrt[3] , n22911);
  not g37866 (n_15331, n22912);
  and g37867 (n22913, n_14831, n_15331);
  not g37868 (n_15332, n22910);
  not g37869 (n_15333, n22913);
  and g37870 (n22914, n_15332, n_15333);
  and g37871 (n22915, n_5034, n_15328);
  and g37872 (n22916, n_15329, n22915);
  not g37873 (n_15334, n22914);
  not g37874 (n_15335, n22916);
  and g37875 (n22917, n_15334, n_15335);
  not g37876 (n_15336, n22907);
  not g37877 (n_15337, n22917);
  and g37878 (n22918, n_15336, n_15337);
  not g37879 (n_15338, n22918);
  and g37880 (n22919, \asqrt[32] , n_15338);
  and g37884 (n22923, n_14841, n_14840);
  and g37885 (n22924, \asqrt[3] , n22923);
  not g37886 (n_15339, n22924);
  and g37887 (n22925, n_14839, n_15339);
  not g37888 (n_15340, n22922);
  not g37889 (n_15341, n22925);
  and g37890 (n22926, n_15340, n_15341);
  and g37891 (n22927, n_4754, n_15336);
  and g37892 (n22928, n_15337, n22927);
  not g37893 (n_15342, n22926);
  not g37894 (n_15343, n22928);
  and g37895 (n22929, n_15342, n_15343);
  not g37896 (n_15344, n22919);
  not g37897 (n_15345, n22929);
  and g37898 (n22930, n_15344, n_15345);
  not g37899 (n_15346, n22930);
  and g37900 (n22931, \asqrt[33] , n_15346);
  and g37904 (n22935, n_14849, n_14848);
  and g37905 (n22936, \asqrt[3] , n22935);
  not g37906 (n_15347, n22936);
  and g37907 (n22937, n_14847, n_15347);
  not g37908 (n_15348, n22934);
  not g37909 (n_15349, n22937);
  and g37910 (n22938, n_15348, n_15349);
  and g37911 (n22939, n_4482, n_15344);
  and g37912 (n22940, n_15345, n22939);
  not g37913 (n_15350, n22938);
  not g37914 (n_15351, n22940);
  and g37915 (n22941, n_15350, n_15351);
  not g37916 (n_15352, n22931);
  not g37917 (n_15353, n22941);
  and g37918 (n22942, n_15352, n_15353);
  not g37919 (n_15354, n22942);
  and g37920 (n22943, \asqrt[34] , n_15354);
  and g37924 (n22947, n_14857, n_14856);
  and g37925 (n22948, \asqrt[3] , n22947);
  not g37926 (n_15355, n22948);
  and g37927 (n22949, n_14855, n_15355);
  not g37928 (n_15356, n22946);
  not g37929 (n_15357, n22949);
  and g37930 (n22950, n_15356, n_15357);
  and g37931 (n22951, n_4218, n_15352);
  and g37932 (n22952, n_15353, n22951);
  not g37933 (n_15358, n22950);
  not g37934 (n_15359, n22952);
  and g37935 (n22953, n_15358, n_15359);
  not g37936 (n_15360, n22943);
  not g37937 (n_15361, n22953);
  and g37938 (n22954, n_15360, n_15361);
  not g37939 (n_15362, n22954);
  and g37940 (n22955, \asqrt[35] , n_15362);
  and g37944 (n22959, n_14865, n_14864);
  and g37945 (n22960, \asqrt[3] , n22959);
  not g37946 (n_15363, n22960);
  and g37947 (n22961, n_14863, n_15363);
  not g37948 (n_15364, n22958);
  not g37949 (n_15365, n22961);
  and g37950 (n22962, n_15364, n_15365);
  and g37951 (n22963, n_3962, n_15360);
  and g37952 (n22964, n_15361, n22963);
  not g37953 (n_15366, n22962);
  not g37954 (n_15367, n22964);
  and g37955 (n22965, n_15366, n_15367);
  not g37956 (n_15368, n22955);
  not g37957 (n_15369, n22965);
  and g37958 (n22966, n_15368, n_15369);
  not g37959 (n_15370, n22966);
  and g37960 (n22967, \asqrt[36] , n_15370);
  and g37964 (n22971, n_14873, n_14872);
  and g37965 (n22972, \asqrt[3] , n22971);
  not g37966 (n_15371, n22972);
  and g37967 (n22973, n_14871, n_15371);
  not g37968 (n_15372, n22970);
  not g37969 (n_15373, n22973);
  and g37970 (n22974, n_15372, n_15373);
  and g37971 (n22975, n_3714, n_15368);
  and g37972 (n22976, n_15369, n22975);
  not g37973 (n_15374, n22974);
  not g37974 (n_15375, n22976);
  and g37975 (n22977, n_15374, n_15375);
  not g37976 (n_15376, n22967);
  not g37977 (n_15377, n22977);
  and g37978 (n22978, n_15376, n_15377);
  not g37979 (n_15378, n22978);
  and g37980 (n22979, \asqrt[37] , n_15378);
  and g37984 (n22983, n_14881, n_14880);
  and g37985 (n22984, \asqrt[3] , n22983);
  not g37986 (n_15379, n22984);
  and g37987 (n22985, n_14879, n_15379);
  not g37988 (n_15380, n22982);
  not g37989 (n_15381, n22985);
  and g37990 (n22986, n_15380, n_15381);
  and g37991 (n22987, n_3474, n_15376);
  and g37992 (n22988, n_15377, n22987);
  not g37993 (n_15382, n22986);
  not g37994 (n_15383, n22988);
  and g37995 (n22989, n_15382, n_15383);
  not g37996 (n_15384, n22979);
  not g37997 (n_15385, n22989);
  and g37998 (n22990, n_15384, n_15385);
  not g37999 (n_15386, n22990);
  and g38000 (n22991, \asqrt[38] , n_15386);
  and g38004 (n22995, n_14889, n_14888);
  and g38005 (n22996, \asqrt[3] , n22995);
  not g38006 (n_15387, n22996);
  and g38007 (n22997, n_14887, n_15387);
  not g38008 (n_15388, n22994);
  not g38009 (n_15389, n22997);
  and g38010 (n22998, n_15388, n_15389);
  and g38011 (n22999, n_3242, n_15384);
  and g38012 (n23000, n_15385, n22999);
  not g38013 (n_15390, n22998);
  not g38014 (n_15391, n23000);
  and g38015 (n23001, n_15390, n_15391);
  not g38016 (n_15392, n22991);
  not g38017 (n_15393, n23001);
  and g38018 (n23002, n_15392, n_15393);
  not g38019 (n_15394, n23002);
  and g38020 (n23003, \asqrt[39] , n_15394);
  and g38024 (n23007, n_14897, n_14896);
  and g38025 (n23008, \asqrt[3] , n23007);
  not g38026 (n_15395, n23008);
  and g38027 (n23009, n_14895, n_15395);
  not g38028 (n_15396, n23006);
  not g38029 (n_15397, n23009);
  and g38030 (n23010, n_15396, n_15397);
  and g38031 (n23011, n_3018, n_15392);
  and g38032 (n23012, n_15393, n23011);
  not g38033 (n_15398, n23010);
  not g38034 (n_15399, n23012);
  and g38035 (n23013, n_15398, n_15399);
  not g38036 (n_15400, n23003);
  not g38037 (n_15401, n23013);
  and g38038 (n23014, n_15400, n_15401);
  not g38039 (n_15402, n23014);
  and g38040 (n23015, \asqrt[40] , n_15402);
  and g38044 (n23019, n_14905, n_14904);
  and g38045 (n23020, \asqrt[3] , n23019);
  not g38046 (n_15403, n23020);
  and g38047 (n23021, n_14903, n_15403);
  not g38048 (n_15404, n23018);
  not g38049 (n_15405, n23021);
  and g38050 (n23022, n_15404, n_15405);
  and g38051 (n23023, n_2802, n_15400);
  and g38052 (n23024, n_15401, n23023);
  not g38053 (n_15406, n23022);
  not g38054 (n_15407, n23024);
  and g38055 (n23025, n_15406, n_15407);
  not g38056 (n_15408, n23015);
  not g38057 (n_15409, n23025);
  and g38058 (n23026, n_15408, n_15409);
  not g38059 (n_15410, n23026);
  and g38060 (n23027, \asqrt[41] , n_15410);
  and g38064 (n23031, n_14913, n_14912);
  and g38065 (n23032, \asqrt[3] , n23031);
  not g38066 (n_15411, n23032);
  and g38067 (n23033, n_14911, n_15411);
  not g38068 (n_15412, n23030);
  not g38069 (n_15413, n23033);
  and g38070 (n23034, n_15412, n_15413);
  and g38071 (n23035, n_2594, n_15408);
  and g38072 (n23036, n_15409, n23035);
  not g38073 (n_15414, n23034);
  not g38074 (n_15415, n23036);
  and g38075 (n23037, n_15414, n_15415);
  not g38076 (n_15416, n23027);
  not g38077 (n_15417, n23037);
  and g38078 (n23038, n_15416, n_15417);
  not g38079 (n_15418, n23038);
  and g38080 (n23039, \asqrt[42] , n_15418);
  and g38084 (n23043, n_14921, n_14920);
  and g38085 (n23044, \asqrt[3] , n23043);
  not g38086 (n_15419, n23044);
  and g38087 (n23045, n_14919, n_15419);
  not g38088 (n_15420, n23042);
  not g38089 (n_15421, n23045);
  and g38090 (n23046, n_15420, n_15421);
  and g38091 (n23047, n_2394, n_15416);
  and g38092 (n23048, n_15417, n23047);
  not g38093 (n_15422, n23046);
  not g38094 (n_15423, n23048);
  and g38095 (n23049, n_15422, n_15423);
  not g38096 (n_15424, n23039);
  not g38097 (n_15425, n23049);
  and g38098 (n23050, n_15424, n_15425);
  not g38099 (n_15426, n23050);
  and g38100 (n23051, \asqrt[43] , n_15426);
  and g38104 (n23055, n_14929, n_14928);
  and g38105 (n23056, \asqrt[3] , n23055);
  not g38106 (n_15427, n23056);
  and g38107 (n23057, n_14927, n_15427);
  not g38108 (n_15428, n23054);
  not g38109 (n_15429, n23057);
  and g38110 (n23058, n_15428, n_15429);
  and g38111 (n23059, n_2202, n_15424);
  and g38112 (n23060, n_15425, n23059);
  not g38113 (n_15430, n23058);
  not g38114 (n_15431, n23060);
  and g38115 (n23061, n_15430, n_15431);
  not g38116 (n_15432, n23051);
  not g38117 (n_15433, n23061);
  and g38118 (n23062, n_15432, n_15433);
  not g38119 (n_15434, n23062);
  and g38120 (n23063, \asqrt[44] , n_15434);
  and g38124 (n23067, n_14937, n_14936);
  and g38125 (n23068, \asqrt[3] , n23067);
  not g38126 (n_15435, n23068);
  and g38127 (n23069, n_14935, n_15435);
  not g38128 (n_15436, n23066);
  not g38129 (n_15437, n23069);
  and g38130 (n23070, n_15436, n_15437);
  and g38131 (n23071, n_2018, n_15432);
  and g38132 (n23072, n_15433, n23071);
  not g38133 (n_15438, n23070);
  not g38134 (n_15439, n23072);
  and g38135 (n23073, n_15438, n_15439);
  not g38136 (n_15440, n23063);
  not g38137 (n_15441, n23073);
  and g38138 (n23074, n_15440, n_15441);
  not g38139 (n_15442, n23074);
  and g38140 (n23075, \asqrt[45] , n_15442);
  and g38144 (n23079, n_14945, n_14944);
  and g38145 (n23080, \asqrt[3] , n23079);
  not g38146 (n_15443, n23080);
  and g38147 (n23081, n_14943, n_15443);
  not g38148 (n_15444, n23078);
  not g38149 (n_15445, n23081);
  and g38150 (n23082, n_15444, n_15445);
  and g38151 (n23083, n_1842, n_15440);
  and g38152 (n23084, n_15441, n23083);
  not g38153 (n_15446, n23082);
  not g38154 (n_15447, n23084);
  and g38155 (n23085, n_15446, n_15447);
  not g38156 (n_15448, n23075);
  not g38157 (n_15449, n23085);
  and g38158 (n23086, n_15448, n_15449);
  not g38159 (n_15450, n23086);
  and g38160 (n23087, \asqrt[46] , n_15450);
  and g38164 (n23091, n_14953, n_14952);
  and g38165 (n23092, \asqrt[3] , n23091);
  not g38166 (n_15451, n23092);
  and g38167 (n23093, n_14951, n_15451);
  not g38168 (n_15452, n23090);
  not g38169 (n_15453, n23093);
  and g38170 (n23094, n_15452, n_15453);
  and g38171 (n23095, n_1674, n_15448);
  and g38172 (n23096, n_15449, n23095);
  not g38173 (n_15454, n23094);
  not g38174 (n_15455, n23096);
  and g38175 (n23097, n_15454, n_15455);
  not g38176 (n_15456, n23087);
  not g38177 (n_15457, n23097);
  and g38178 (n23098, n_15456, n_15457);
  not g38179 (n_15458, n23098);
  and g38180 (n23099, \asqrt[47] , n_15458);
  and g38184 (n23103, n_14961, n_14960);
  and g38185 (n23104, \asqrt[3] , n23103);
  not g38186 (n_15459, n23104);
  and g38187 (n23105, n_14959, n_15459);
  not g38188 (n_15460, n23102);
  not g38189 (n_15461, n23105);
  and g38190 (n23106, n_15460, n_15461);
  and g38191 (n23107, n_1514, n_15456);
  and g38192 (n23108, n_15457, n23107);
  not g38193 (n_15462, n23106);
  not g38194 (n_15463, n23108);
  and g38195 (n23109, n_15462, n_15463);
  not g38196 (n_15464, n23099);
  not g38197 (n_15465, n23109);
  and g38198 (n23110, n_15464, n_15465);
  not g38199 (n_15466, n23110);
  and g38200 (n23111, \asqrt[48] , n_15466);
  and g38204 (n23115, n_14969, n_14968);
  and g38205 (n23116, \asqrt[3] , n23115);
  not g38206 (n_15467, n23116);
  and g38207 (n23117, n_14967, n_15467);
  not g38208 (n_15468, n23114);
  not g38209 (n_15469, n23117);
  and g38210 (n23118, n_15468, n_15469);
  and g38211 (n23119, n_1362, n_15464);
  and g38212 (n23120, n_15465, n23119);
  not g38213 (n_15470, n23118);
  not g38214 (n_15471, n23120);
  and g38215 (n23121, n_15470, n_15471);
  not g38216 (n_15472, n23111);
  not g38217 (n_15473, n23121);
  and g38218 (n23122, n_15472, n_15473);
  not g38219 (n_15474, n23122);
  and g38220 (n23123, \asqrt[49] , n_15474);
  and g38224 (n23127, n_14977, n_14976);
  and g38225 (n23128, \asqrt[3] , n23127);
  not g38226 (n_15475, n23128);
  and g38227 (n23129, n_14975, n_15475);
  not g38228 (n_15476, n23126);
  not g38229 (n_15477, n23129);
  and g38230 (n23130, n_15476, n_15477);
  and g38231 (n23131, n_1218, n_15472);
  and g38232 (n23132, n_15473, n23131);
  not g38233 (n_15478, n23130);
  not g38234 (n_15479, n23132);
  and g38235 (n23133, n_15478, n_15479);
  not g38236 (n_15480, n23123);
  not g38237 (n_15481, n23133);
  and g38238 (n23134, n_15480, n_15481);
  not g38239 (n_15482, n23134);
  and g38240 (n23135, \asqrt[50] , n_15482);
  and g38244 (n23139, n_14985, n_14984);
  and g38245 (n23140, \asqrt[3] , n23139);
  not g38246 (n_15483, n23140);
  and g38247 (n23141, n_14983, n_15483);
  not g38248 (n_15484, n23138);
  not g38249 (n_15485, n23141);
  and g38250 (n23142, n_15484, n_15485);
  and g38251 (n23143, n_1082, n_15480);
  and g38252 (n23144, n_15481, n23143);
  not g38253 (n_15486, n23142);
  not g38254 (n_15487, n23144);
  and g38255 (n23145, n_15486, n_15487);
  not g38256 (n_15488, n23135);
  not g38257 (n_15489, n23145);
  and g38258 (n23146, n_15488, n_15489);
  not g38259 (n_15490, n23146);
  and g38260 (n23147, \asqrt[51] , n_15490);
  and g38264 (n23151, n_14993, n_14992);
  and g38265 (n23152, \asqrt[3] , n23151);
  not g38266 (n_15491, n23152);
  and g38267 (n23153, n_14991, n_15491);
  not g38268 (n_15492, n23150);
  not g38269 (n_15493, n23153);
  and g38270 (n23154, n_15492, n_15493);
  and g38271 (n23155, n_954, n_15488);
  and g38272 (n23156, n_15489, n23155);
  not g38273 (n_15494, n23154);
  not g38274 (n_15495, n23156);
  and g38275 (n23157, n_15494, n_15495);
  not g38276 (n_15496, n23147);
  not g38277 (n_15497, n23157);
  and g38278 (n23158, n_15496, n_15497);
  not g38279 (n_15498, n23158);
  and g38280 (n23159, \asqrt[52] , n_15498);
  and g38284 (n23163, n_15001, n_15000);
  and g38285 (n23164, \asqrt[3] , n23163);
  not g38286 (n_15499, n23164);
  and g38287 (n23165, n_14999, n_15499);
  not g38288 (n_15500, n23162);
  not g38289 (n_15501, n23165);
  and g38290 (n23166, n_15500, n_15501);
  and g38291 (n23167, n_834, n_15496);
  and g38292 (n23168, n_15497, n23167);
  not g38293 (n_15502, n23166);
  not g38294 (n_15503, n23168);
  and g38295 (n23169, n_15502, n_15503);
  not g38296 (n_15504, n23159);
  not g38297 (n_15505, n23169);
  and g38298 (n23170, n_15504, n_15505);
  not g38299 (n_15506, n23170);
  and g38300 (n23171, \asqrt[53] , n_15506);
  and g38304 (n23175, n_15009, n_15008);
  and g38305 (n23176, \asqrt[3] , n23175);
  not g38306 (n_15507, n23176);
  and g38307 (n23177, n_15007, n_15507);
  not g38308 (n_15508, n23174);
  not g38309 (n_15509, n23177);
  and g38310 (n23178, n_15508, n_15509);
  and g38311 (n23179, n_722, n_15504);
  and g38312 (n23180, n_15505, n23179);
  not g38313 (n_15510, n23178);
  not g38314 (n_15511, n23180);
  and g38315 (n23181, n_15510, n_15511);
  not g38316 (n_15512, n23171);
  not g38317 (n_15513, n23181);
  and g38318 (n23182, n_15512, n_15513);
  not g38319 (n_15514, n23182);
  and g38320 (n23183, \asqrt[54] , n_15514);
  and g38324 (n23187, n_15017, n_15016);
  and g38325 (n23188, \asqrt[3] , n23187);
  not g38326 (n_15515, n23188);
  and g38327 (n23189, n_15015, n_15515);
  not g38328 (n_15516, n23186);
  not g38329 (n_15517, n23189);
  and g38330 (n23190, n_15516, n_15517);
  and g38331 (n23191, n_618, n_15512);
  and g38332 (n23192, n_15513, n23191);
  not g38333 (n_15518, n23190);
  not g38334 (n_15519, n23192);
  and g38335 (n23193, n_15518, n_15519);
  not g38336 (n_15520, n23183);
  not g38337 (n_15521, n23193);
  and g38338 (n23194, n_15520, n_15521);
  not g38339 (n_15522, n23194);
  and g38340 (n23195, \asqrt[55] , n_15522);
  and g38344 (n23199, n_15025, n_15024);
  and g38345 (n23200, \asqrt[3] , n23199);
  not g38346 (n_15523, n23200);
  and g38347 (n23201, n_15023, n_15523);
  not g38348 (n_15524, n23198);
  not g38349 (n_15525, n23201);
  and g38350 (n23202, n_15524, n_15525);
  and g38351 (n23203, n_522, n_15520);
  and g38352 (n23204, n_15521, n23203);
  not g38353 (n_15526, n23202);
  not g38354 (n_15527, n23204);
  and g38355 (n23205, n_15526, n_15527);
  not g38356 (n_15528, n23195);
  not g38357 (n_15529, n23205);
  and g38358 (n23206, n_15528, n_15529);
  not g38359 (n_15530, n23206);
  and g38360 (n23207, \asqrt[56] , n_15530);
  and g38364 (n23211, n_15033, n_15032);
  and g38365 (n23212, \asqrt[3] , n23211);
  not g38366 (n_15531, n23212);
  and g38367 (n23213, n_15031, n_15531);
  not g38368 (n_15532, n23210);
  not g38369 (n_15533, n23213);
  and g38370 (n23214, n_15532, n_15533);
  and g38371 (n23215, n_434, n_15528);
  and g38372 (n23216, n_15529, n23215);
  not g38373 (n_15534, n23214);
  not g38374 (n_15535, n23216);
  and g38375 (n23217, n_15534, n_15535);
  not g38376 (n_15536, n23207);
  not g38377 (n_15537, n23217);
  and g38378 (n23218, n_15536, n_15537);
  not g38379 (n_15538, n23218);
  and g38380 (n23219, \asqrt[57] , n_15538);
  and g38384 (n23223, n_15041, n_15040);
  and g38385 (n23224, \asqrt[3] , n23223);
  not g38386 (n_15539, n23224);
  and g38387 (n23225, n_15039, n_15539);
  not g38388 (n_15540, n23222);
  not g38389 (n_15541, n23225);
  and g38390 (n23226, n_15540, n_15541);
  and g38391 (n23227, n_354, n_15536);
  and g38392 (n23228, n_15537, n23227);
  not g38393 (n_15542, n23226);
  not g38394 (n_15543, n23228);
  and g38395 (n23229, n_15542, n_15543);
  not g38396 (n_15544, n23219);
  not g38397 (n_15545, n23229);
  and g38398 (n23230, n_15544, n_15545);
  not g38399 (n_15546, n23230);
  and g38400 (n23231, \asqrt[58] , n_15546);
  and g38404 (n23235, n_15049, n_15048);
  and g38405 (n23236, \asqrt[3] , n23235);
  not g38406 (n_15547, n23236);
  and g38407 (n23237, n_15047, n_15547);
  not g38408 (n_15548, n23234);
  not g38409 (n_15549, n23237);
  and g38410 (n23238, n_15548, n_15549);
  and g38411 (n23239, n_282, n_15544);
  and g38412 (n23240, n_15545, n23239);
  not g38413 (n_15550, n23238);
  not g38414 (n_15551, n23240);
  and g38415 (n23241, n_15550, n_15551);
  not g38416 (n_15552, n23231);
  not g38417 (n_15553, n23241);
  and g38418 (n23242, n_15552, n_15553);
  not g38419 (n_15554, n23242);
  and g38420 (n23243, \asqrt[59] , n_15554);
  and g38424 (n23247, n_15057, n_15056);
  and g38425 (n23248, \asqrt[3] , n23247);
  not g38426 (n_15555, n23248);
  and g38427 (n23249, n_15055, n_15555);
  not g38428 (n_15556, n23246);
  not g38429 (n_15557, n23249);
  and g38430 (n23250, n_15556, n_15557);
  and g38431 (n23251, n_218, n_15552);
  and g38432 (n23252, n_15553, n23251);
  not g38433 (n_15558, n23250);
  not g38434 (n_15559, n23252);
  and g38435 (n23253, n_15558, n_15559);
  not g38436 (n_15560, n23243);
  not g38437 (n_15561, n23253);
  and g38438 (n23254, n_15560, n_15561);
  not g38439 (n_15562, n23254);
  and g38440 (n23255, \asqrt[60] , n_15562);
  and g38444 (n23259, n_15065, n_15064);
  and g38445 (n23260, \asqrt[3] , n23259);
  not g38446 (n_15563, n23260);
  and g38447 (n23261, n_15063, n_15563);
  not g38448 (n_15564, n23258);
  not g38449 (n_15565, n23261);
  and g38450 (n23262, n_15564, n_15565);
  and g38451 (n23263, n_162, n_15560);
  and g38452 (n23264, n_15561, n23263);
  not g38453 (n_15566, n23262);
  not g38454 (n_15567, n23264);
  and g38455 (n23265, n_15566, n_15567);
  not g38456 (n_15568, n23255);
  not g38457 (n_15569, n23265);
  and g38458 (n23266, n_15568, n_15569);
  not g38459 (n_15570, n23266);
  and g38460 (n23267, \asqrt[61] , n_15570);
  and g38464 (n23271, n_15073, n_15072);
  and g38465 (n23272, \asqrt[3] , n23271);
  not g38466 (n_15571, n23272);
  and g38467 (n23273, n_15071, n_15571);
  not g38468 (n_15572, n23270);
  not g38469 (n_15573, n23273);
  and g38470 (n23274, n_15572, n_15573);
  and g38471 (n23275, n_115, n_15568);
  and g38472 (n23276, n_15569, n23275);
  not g38473 (n_15574, n23274);
  not g38474 (n_15575, n23276);
  and g38475 (n23277, n_15574, n_15575);
  not g38476 (n_15576, n23267);
  not g38477 (n_15577, n23277);
  and g38478 (n23278, n_15576, n_15577);
  not g38479 (n_15578, n23278);
  and g38480 (n23279, \asqrt[62] , n_15578);
  and g38481 (n23280, n_76, n_15576);
  and g38482 (n23281, n_15577, n23280);
  and g38486 (n23285, n_15081, n_15079);
  and g38487 (n23286, \asqrt[3] , n23285);
  not g38488 (n_15579, n23286);
  and g38489 (n23287, n_15080, n_15579);
  not g38490 (n_15580, n23284);
  not g38491 (n_15581, n23287);
  and g38492 (n23288, n_15580, n_15581);
  not g38493 (n_15582, n23281);
  not g38494 (n_15583, n23288);
  and g38495 (n23289, n_15582, n_15583);
  not g38496 (n_15584, n23279);
  not g38497 (n_15585, n23289);
  and g38498 (n23290, n_15584, n_15585);
  and g38502 (n23294, n_15089, n_15088);
  and g38503 (n23295, \asqrt[3] , n23294);
  not g38504 (n_15586, n23295);
  and g38505 (n23296, n_15087, n_15586);
  not g38506 (n_15587, n23293);
  not g38507 (n_15588, n23296);
  and g38508 (n23297, n_15587, n_15588);
  and g38509 (n23298, n_15096, n_15095);
  and g38510 (n23299, \asqrt[3] , n23298);
  not g38513 (n_15590, n23297);
  not g38515 (n_15591, n23290);
  not g38517 (n_15592, n23302);
  and g38518 (n23303, n_21, n_15592);
  and g38519 (n23304, n_15584, n23297);
  and g38520 (n23305, n_15585, n23304);
  and g38521 (n23306, n_15095, \asqrt[3] );
  not g38522 (n_15593, n23306);
  and g38523 (n23307, n22558, n_15593);
  not g38524 (n_15594, n23298);
  and g38525 (n23308, \asqrt[63] , n_15594);
  not g38526 (n_15595, n23307);
  and g38527 (n23309, n_15595, n23308);
  not g38528 (n_15596, n23305);
  not g38529 (n_15597, n23309);
  and g38530 (n23310, n_15596, n_15597);
  not g38531 (n_15598, n23310);
  or g38532 (\asqrt[2] , n23303, n_15598);
  and g38536 (n23315, n_15568, n_15567);
  and g38537 (n23316, \asqrt[2] , n23315);
  not g38538 (n_15600, n23316);
  and g38539 (n23317, n_15566, n_15600);
  not g38540 (n_15601, n23314);
  not g38541 (n_15602, n23317);
  and g38542 (n23318, n_15601, n_15602);
  and g38543 (n23319, \a[4] , \asqrt[2] );
  not g38544 (n_15605, \a[2] );
  not g38545 (n_15606, \a[3] );
  and g38546 (n23320, n_15605, n_15606);
  and g38547 (n23321, n_15107, n23320);
  not g38548 (n_15607, n23319);
  not g38549 (n_15608, n23321);
  and g38550 (n23322, n_15607, n_15608);
  not g38551 (n_15609, n23322);
  and g38552 (n23323, \asqrt[3] , n_15609);
  and g38557 (n23328, n_15107, \asqrt[2] );
  not g38558 (n_15610, n23328);
  and g38559 (n23329, \a[5] , n_15610);
  and g38560 (n23330, n22581, \asqrt[2] );
  not g38561 (n_15611, n23329);
  not g38562 (n_15612, n23330);
  and g38563 (n23331, n_15611, n_15612);
  not g38564 (n_15613, n23327);
  and g38565 (n23332, n_15613, n23331);
  not g38566 (n_15614, n23323);
  not g38567 (n_15615, n23332);
  and g38568 (n23333, n_15614, n_15615);
  not g38569 (n_15616, n23333);
  and g38570 (n23334, \asqrt[4] , n_15616);
  not g38571 (n_15617, \asqrt[4] );
  and g38572 (n23335, n_15617, n_15614);
  and g38573 (n23336, n_15615, n23335);
  not g38578 (n_15619, n23339);
  and g38579 (n23340, n_15612, n_15619);
  not g38580 (n_15620, n23340);
  and g38581 (n23341, \a[6] , n_15620);
  and g38582 (n23342, n_14620, n_15619);
  and g38583 (n23343, n_15612, n23342);
  not g38584 (n_15621, n23341);
  not g38585 (n_15622, n23343);
  and g38586 (n23344, n_15621, n_15622);
  not g38587 (n_15623, n23336);
  not g38588 (n_15624, n23344);
  and g38589 (n23345, n_15623, n_15624);
  not g38590 (n_15625, n23334);
  not g38591 (n_15626, n23345);
  and g38592 (n23346, n_15625, n_15626);
  not g38593 (n_15627, n23346);
  and g38594 (n23347, \asqrt[5] , n_15627);
  and g38595 (n23348, n_15116, n_15115);
  not g38596 (n_15628, n22592);
  and g38597 (n23349, n_15628, n23348);
  and g38598 (n23350, \asqrt[2] , n23349);
  and g38599 (n23351, \asqrt[2] , n23348);
  not g38600 (n_15629, n23351);
  and g38601 (n23352, n22592, n_15629);
  not g38602 (n_15630, n23350);
  not g38603 (n_15631, n23352);
  and g38604 (n23353, n_15630, n_15631);
  and g38605 (n23354, n_15119, n_15625);
  and g38606 (n23355, n_15626, n23354);
  not g38607 (n_15632, n23353);
  not g38608 (n_15633, n23355);
  and g38609 (n23356, n_15632, n_15633);
  not g38610 (n_15634, n23347);
  not g38611 (n_15635, n23356);
  and g38612 (n23357, n_15634, n_15635);
  not g38613 (n_15636, n23357);
  and g38614 (n23358, \asqrt[6] , n_15636);
  and g38618 (n23362, n_15127, n_15125);
  and g38619 (n23363, \asqrt[2] , n23362);
  not g38620 (n_15637, n23363);
  and g38621 (n23364, n_15126, n_15637);
  not g38622 (n_15638, n23361);
  not g38623 (n_15639, n23364);
  and g38624 (n23365, n_15638, n_15639);
  and g38625 (n23366, n_14632, n_15634);
  and g38626 (n23367, n_15635, n23366);
  not g38627 (n_15640, n23365);
  not g38628 (n_15641, n23367);
  and g38629 (n23368, n_15640, n_15641);
  not g38630 (n_15642, n23358);
  not g38631 (n_15643, n23368);
  and g38632 (n23369, n_15642, n_15643);
  not g38633 (n_15644, n23369);
  and g38634 (n23370, \asqrt[7] , n_15644);
  and g38638 (n23374, n_15136, n_15135);
  and g38639 (n23375, \asqrt[2] , n23374);
  not g38640 (n_15645, n23375);
  and g38641 (n23376, n_15134, n_15645);
  not g38642 (n_15646, n23373);
  not g38643 (n_15647, n23376);
  and g38644 (n23377, n_15646, n_15647);
  and g38645 (n23378, n_14153, n_15642);
  and g38646 (n23379, n_15643, n23378);
  not g38647 (n_15648, n23377);
  not g38648 (n_15649, n23379);
  and g38649 (n23380, n_15648, n_15649);
  not g38650 (n_15650, n23370);
  not g38651 (n_15651, n23380);
  and g38652 (n23381, n_15650, n_15651);
  not g38653 (n_15652, n23381);
  and g38654 (n23382, \asqrt[8] , n_15652);
  and g38658 (n23386, n_15144, n_15143);
  and g38659 (n23387, \asqrt[2] , n23386);
  not g38660 (n_15653, n23387);
  and g38661 (n23388, n_15142, n_15653);
  not g38662 (n_15654, n23385);
  not g38663 (n_15655, n23388);
  and g38664 (n23389, n_15654, n_15655);
  and g38665 (n23390, n_13682, n_15650);
  and g38666 (n23391, n_15651, n23390);
  not g38667 (n_15656, n23389);
  not g38668 (n_15657, n23391);
  and g38669 (n23392, n_15656, n_15657);
  not g38670 (n_15658, n23382);
  not g38671 (n_15659, n23392);
  and g38672 (n23393, n_15658, n_15659);
  not g38673 (n_15660, n23393);
  and g38674 (n23394, \asqrt[9] , n_15660);
  and g38678 (n23398, n_15152, n_15151);
  and g38679 (n23399, \asqrt[2] , n23398);
  not g38680 (n_15661, n23399);
  and g38681 (n23400, n_15150, n_15661);
  not g38682 (n_15662, n23397);
  not g38683 (n_15663, n23400);
  and g38684 (n23401, n_15662, n_15663);
  and g38685 (n23402, n_13218, n_15658);
  and g38686 (n23403, n_15659, n23402);
  not g38687 (n_15664, n23401);
  not g38688 (n_15665, n23403);
  and g38689 (n23404, n_15664, n_15665);
  not g38690 (n_15666, n23394);
  not g38691 (n_15667, n23404);
  and g38692 (n23405, n_15666, n_15667);
  not g38693 (n_15668, n23405);
  and g38694 (n23406, \asqrt[10] , n_15668);
  and g38698 (n23410, n_15160, n_15159);
  and g38699 (n23411, \asqrt[2] , n23410);
  not g38700 (n_15669, n23411);
  and g38701 (n23412, n_15158, n_15669);
  not g38702 (n_15670, n23409);
  not g38703 (n_15671, n23412);
  and g38704 (n23413, n_15670, n_15671);
  and g38705 (n23414, n_12762, n_15666);
  and g38706 (n23415, n_15667, n23414);
  not g38707 (n_15672, n23413);
  not g38708 (n_15673, n23415);
  and g38709 (n23416, n_15672, n_15673);
  not g38710 (n_15674, n23406);
  not g38711 (n_15675, n23416);
  and g38712 (n23417, n_15674, n_15675);
  not g38713 (n_15676, n23417);
  and g38714 (n23418, \asqrt[11] , n_15676);
  and g38718 (n23422, n_15168, n_15167);
  and g38719 (n23423, \asqrt[2] , n23422);
  not g38720 (n_15677, n23423);
  and g38721 (n23424, n_15166, n_15677);
  not g38722 (n_15678, n23421);
  not g38723 (n_15679, n23424);
  and g38724 (n23425, n_15678, n_15679);
  and g38725 (n23426, n_12314, n_15674);
  and g38726 (n23427, n_15675, n23426);
  not g38727 (n_15680, n23425);
  not g38728 (n_15681, n23427);
  and g38729 (n23428, n_15680, n_15681);
  not g38730 (n_15682, n23418);
  not g38731 (n_15683, n23428);
  and g38732 (n23429, n_15682, n_15683);
  not g38733 (n_15684, n23429);
  and g38734 (n23430, \asqrt[12] , n_15684);
  and g38738 (n23434, n_15176, n_15175);
  and g38739 (n23435, \asqrt[2] , n23434);
  not g38740 (n_15685, n23435);
  and g38741 (n23436, n_15174, n_15685);
  not g38742 (n_15686, n23433);
  not g38743 (n_15687, n23436);
  and g38744 (n23437, n_15686, n_15687);
  and g38745 (n23438, n_11874, n_15682);
  and g38746 (n23439, n_15683, n23438);
  not g38747 (n_15688, n23437);
  not g38748 (n_15689, n23439);
  and g38749 (n23440, n_15688, n_15689);
  not g38750 (n_15690, n23430);
  not g38751 (n_15691, n23440);
  and g38752 (n23441, n_15690, n_15691);
  not g38753 (n_15692, n23441);
  and g38754 (n23442, \asqrt[13] , n_15692);
  and g38758 (n23446, n_15184, n_15183);
  and g38759 (n23447, \asqrt[2] , n23446);
  not g38760 (n_15693, n23447);
  and g38761 (n23448, n_15182, n_15693);
  not g38762 (n_15694, n23445);
  not g38763 (n_15695, n23448);
  and g38764 (n23449, n_15694, n_15695);
  and g38765 (n23450, n_11442, n_15690);
  and g38766 (n23451, n_15691, n23450);
  not g38767 (n_15696, n23449);
  not g38768 (n_15697, n23451);
  and g38769 (n23452, n_15696, n_15697);
  not g38770 (n_15698, n23442);
  not g38771 (n_15699, n23452);
  and g38772 (n23453, n_15698, n_15699);
  not g38773 (n_15700, n23453);
  and g38774 (n23454, \asqrt[14] , n_15700);
  and g38778 (n23458, n_15192, n_15191);
  and g38779 (n23459, \asqrt[2] , n23458);
  not g38780 (n_15701, n23459);
  and g38781 (n23460, n_15190, n_15701);
  not g38782 (n_15702, n23457);
  not g38783 (n_15703, n23460);
  and g38784 (n23461, n_15702, n_15703);
  and g38785 (n23462, n_11018, n_15698);
  and g38786 (n23463, n_15699, n23462);
  not g38787 (n_15704, n23461);
  not g38788 (n_15705, n23463);
  and g38789 (n23464, n_15704, n_15705);
  not g38790 (n_15706, n23454);
  not g38791 (n_15707, n23464);
  and g38792 (n23465, n_15706, n_15707);
  not g38793 (n_15708, n23465);
  and g38794 (n23466, \asqrt[15] , n_15708);
  and g38798 (n23470, n_15200, n_15199);
  and g38799 (n23471, \asqrt[2] , n23470);
  not g38800 (n_15709, n23471);
  and g38801 (n23472, n_15198, n_15709);
  not g38802 (n_15710, n23469);
  not g38803 (n_15711, n23472);
  and g38804 (n23473, n_15710, n_15711);
  and g38805 (n23474, n_10602, n_15706);
  and g38806 (n23475, n_15707, n23474);
  not g38807 (n_15712, n23473);
  not g38808 (n_15713, n23475);
  and g38809 (n23476, n_15712, n_15713);
  not g38810 (n_15714, n23466);
  not g38811 (n_15715, n23476);
  and g38812 (n23477, n_15714, n_15715);
  not g38813 (n_15716, n23477);
  and g38814 (n23478, \asqrt[16] , n_15716);
  and g38818 (n23482, n_15208, n_15207);
  and g38819 (n23483, \asqrt[2] , n23482);
  not g38820 (n_15717, n23483);
  and g38821 (n23484, n_15206, n_15717);
  not g38822 (n_15718, n23481);
  not g38823 (n_15719, n23484);
  and g38824 (n23485, n_15718, n_15719);
  and g38825 (n23486, n_10194, n_15714);
  and g38826 (n23487, n_15715, n23486);
  not g38827 (n_15720, n23485);
  not g38828 (n_15721, n23487);
  and g38829 (n23488, n_15720, n_15721);
  not g38830 (n_15722, n23478);
  not g38831 (n_15723, n23488);
  and g38832 (n23489, n_15722, n_15723);
  not g38833 (n_15724, n23489);
  and g38834 (n23490, \asqrt[17] , n_15724);
  and g38838 (n23494, n_15216, n_15215);
  and g38839 (n23495, \asqrt[2] , n23494);
  not g38840 (n_15725, n23495);
  and g38841 (n23496, n_15214, n_15725);
  not g38842 (n_15726, n23493);
  not g38843 (n_15727, n23496);
  and g38844 (n23497, n_15726, n_15727);
  and g38845 (n23498, n_9794, n_15722);
  and g38846 (n23499, n_15723, n23498);
  not g38847 (n_15728, n23497);
  not g38848 (n_15729, n23499);
  and g38849 (n23500, n_15728, n_15729);
  not g38850 (n_15730, n23490);
  not g38851 (n_15731, n23500);
  and g38852 (n23501, n_15730, n_15731);
  not g38853 (n_15732, n23501);
  and g38854 (n23502, \asqrt[18] , n_15732);
  and g38858 (n23506, n_15224, n_15223);
  and g38859 (n23507, \asqrt[2] , n23506);
  not g38860 (n_15733, n23507);
  and g38861 (n23508, n_15222, n_15733);
  not g38862 (n_15734, n23505);
  not g38863 (n_15735, n23508);
  and g38864 (n23509, n_15734, n_15735);
  and g38865 (n23510, n_9402, n_15730);
  and g38866 (n23511, n_15731, n23510);
  not g38867 (n_15736, n23509);
  not g38868 (n_15737, n23511);
  and g38869 (n23512, n_15736, n_15737);
  not g38870 (n_15738, n23502);
  not g38871 (n_15739, n23512);
  and g38872 (n23513, n_15738, n_15739);
  not g38873 (n_15740, n23513);
  and g38874 (n23514, \asqrt[19] , n_15740);
  and g38878 (n23518, n_15232, n_15231);
  and g38879 (n23519, \asqrt[2] , n23518);
  not g38880 (n_15741, n23519);
  and g38881 (n23520, n_15230, n_15741);
  not g38882 (n_15742, n23517);
  not g38883 (n_15743, n23520);
  and g38884 (n23521, n_15742, n_15743);
  and g38885 (n23522, n_9018, n_15738);
  and g38886 (n23523, n_15739, n23522);
  not g38887 (n_15744, n23521);
  not g38888 (n_15745, n23523);
  and g38889 (n23524, n_15744, n_15745);
  not g38890 (n_15746, n23514);
  not g38891 (n_15747, n23524);
  and g38892 (n23525, n_15746, n_15747);
  not g38893 (n_15748, n23525);
  and g38894 (n23526, \asqrt[20] , n_15748);
  and g38898 (n23530, n_15240, n_15239);
  and g38899 (n23531, \asqrt[2] , n23530);
  not g38900 (n_15749, n23531);
  and g38901 (n23532, n_15238, n_15749);
  not g38902 (n_15750, n23529);
  not g38903 (n_15751, n23532);
  and g38904 (n23533, n_15750, n_15751);
  and g38905 (n23534, n_8642, n_15746);
  and g38906 (n23535, n_15747, n23534);
  not g38907 (n_15752, n23533);
  not g38908 (n_15753, n23535);
  and g38909 (n23536, n_15752, n_15753);
  not g38910 (n_15754, n23526);
  not g38911 (n_15755, n23536);
  and g38912 (n23537, n_15754, n_15755);
  not g38913 (n_15756, n23537);
  and g38914 (n23538, \asqrt[21] , n_15756);
  and g38918 (n23542, n_15248, n_15247);
  and g38919 (n23543, \asqrt[2] , n23542);
  not g38920 (n_15757, n23543);
  and g38921 (n23544, n_15246, n_15757);
  not g38922 (n_15758, n23541);
  not g38923 (n_15759, n23544);
  and g38924 (n23545, n_15758, n_15759);
  and g38925 (n23546, n_8274, n_15754);
  and g38926 (n23547, n_15755, n23546);
  not g38927 (n_15760, n23545);
  not g38928 (n_15761, n23547);
  and g38929 (n23548, n_15760, n_15761);
  not g38930 (n_15762, n23538);
  not g38931 (n_15763, n23548);
  and g38932 (n23549, n_15762, n_15763);
  not g38933 (n_15764, n23549);
  and g38934 (n23550, \asqrt[22] , n_15764);
  and g38938 (n23554, n_15256, n_15255);
  and g38939 (n23555, \asqrt[2] , n23554);
  not g38940 (n_15765, n23555);
  and g38941 (n23556, n_15254, n_15765);
  not g38942 (n_15766, n23553);
  not g38943 (n_15767, n23556);
  and g38944 (n23557, n_15766, n_15767);
  and g38945 (n23558, n_7914, n_15762);
  and g38946 (n23559, n_15763, n23558);
  not g38947 (n_15768, n23557);
  not g38948 (n_15769, n23559);
  and g38949 (n23560, n_15768, n_15769);
  not g38950 (n_15770, n23550);
  not g38951 (n_15771, n23560);
  and g38952 (n23561, n_15770, n_15771);
  not g38953 (n_15772, n23561);
  and g38954 (n23562, \asqrt[23] , n_15772);
  and g38958 (n23566, n_15264, n_15263);
  and g38959 (n23567, \asqrt[2] , n23566);
  not g38960 (n_15773, n23567);
  and g38961 (n23568, n_15262, n_15773);
  not g38962 (n_15774, n23565);
  not g38963 (n_15775, n23568);
  and g38964 (n23569, n_15774, n_15775);
  and g38965 (n23570, n_7562, n_15770);
  and g38966 (n23571, n_15771, n23570);
  not g38967 (n_15776, n23569);
  not g38968 (n_15777, n23571);
  and g38969 (n23572, n_15776, n_15777);
  not g38970 (n_15778, n23562);
  not g38971 (n_15779, n23572);
  and g38972 (n23573, n_15778, n_15779);
  not g38973 (n_15780, n23573);
  and g38974 (n23574, \asqrt[24] , n_15780);
  and g38978 (n23578, n_15272, n_15271);
  and g38979 (n23579, \asqrt[2] , n23578);
  not g38980 (n_15781, n23579);
  and g38981 (n23580, n_15270, n_15781);
  not g38982 (n_15782, n23577);
  not g38983 (n_15783, n23580);
  and g38984 (n23581, n_15782, n_15783);
  and g38985 (n23582, n_7218, n_15778);
  and g38986 (n23583, n_15779, n23582);
  not g38987 (n_15784, n23581);
  not g38988 (n_15785, n23583);
  and g38989 (n23584, n_15784, n_15785);
  not g38990 (n_15786, n23574);
  not g38991 (n_15787, n23584);
  and g38992 (n23585, n_15786, n_15787);
  not g38993 (n_15788, n23585);
  and g38994 (n23586, \asqrt[25] , n_15788);
  and g38998 (n23590, n_15280, n_15279);
  and g38999 (n23591, \asqrt[2] , n23590);
  not g39000 (n_15789, n23591);
  and g39001 (n23592, n_15278, n_15789);
  not g39002 (n_15790, n23589);
  not g39003 (n_15791, n23592);
  and g39004 (n23593, n_15790, n_15791);
  and g39005 (n23594, n_6882, n_15786);
  and g39006 (n23595, n_15787, n23594);
  not g39007 (n_15792, n23593);
  not g39008 (n_15793, n23595);
  and g39009 (n23596, n_15792, n_15793);
  not g39010 (n_15794, n23586);
  not g39011 (n_15795, n23596);
  and g39012 (n23597, n_15794, n_15795);
  not g39013 (n_15796, n23597);
  and g39014 (n23598, \asqrt[26] , n_15796);
  and g39018 (n23602, n_15288, n_15287);
  and g39019 (n23603, \asqrt[2] , n23602);
  not g39020 (n_15797, n23603);
  and g39021 (n23604, n_15286, n_15797);
  not g39022 (n_15798, n23601);
  not g39023 (n_15799, n23604);
  and g39024 (n23605, n_15798, n_15799);
  and g39025 (n23606, n_6554, n_15794);
  and g39026 (n23607, n_15795, n23606);
  not g39027 (n_15800, n23605);
  not g39028 (n_15801, n23607);
  and g39029 (n23608, n_15800, n_15801);
  not g39030 (n_15802, n23598);
  not g39031 (n_15803, n23608);
  and g39032 (n23609, n_15802, n_15803);
  not g39033 (n_15804, n23609);
  and g39034 (n23610, \asqrt[27] , n_15804);
  and g39038 (n23614, n_15296, n_15295);
  and g39039 (n23615, \asqrt[2] , n23614);
  not g39040 (n_15805, n23615);
  and g39041 (n23616, n_15294, n_15805);
  not g39042 (n_15806, n23613);
  not g39043 (n_15807, n23616);
  and g39044 (n23617, n_15806, n_15807);
  and g39045 (n23618, n_6234, n_15802);
  and g39046 (n23619, n_15803, n23618);
  not g39047 (n_15808, n23617);
  not g39048 (n_15809, n23619);
  and g39049 (n23620, n_15808, n_15809);
  not g39050 (n_15810, n23610);
  not g39051 (n_15811, n23620);
  and g39052 (n23621, n_15810, n_15811);
  not g39053 (n_15812, n23621);
  and g39054 (n23622, \asqrt[28] , n_15812);
  and g39058 (n23626, n_15304, n_15303);
  and g39059 (n23627, \asqrt[2] , n23626);
  not g39060 (n_15813, n23627);
  and g39061 (n23628, n_15302, n_15813);
  not g39062 (n_15814, n23625);
  not g39063 (n_15815, n23628);
  and g39064 (n23629, n_15814, n_15815);
  and g39065 (n23630, n_5922, n_15810);
  and g39066 (n23631, n_15811, n23630);
  not g39067 (n_15816, n23629);
  not g39068 (n_15817, n23631);
  and g39069 (n23632, n_15816, n_15817);
  not g39070 (n_15818, n23622);
  not g39071 (n_15819, n23632);
  and g39072 (n23633, n_15818, n_15819);
  not g39073 (n_15820, n23633);
  and g39074 (n23634, \asqrt[29] , n_15820);
  and g39078 (n23638, n_15312, n_15311);
  and g39079 (n23639, \asqrt[2] , n23638);
  not g39080 (n_15821, n23639);
  and g39081 (n23640, n_15310, n_15821);
  not g39082 (n_15822, n23637);
  not g39083 (n_15823, n23640);
  and g39084 (n23641, n_15822, n_15823);
  and g39085 (n23642, n_5618, n_15818);
  and g39086 (n23643, n_15819, n23642);
  not g39087 (n_15824, n23641);
  not g39088 (n_15825, n23643);
  and g39089 (n23644, n_15824, n_15825);
  not g39090 (n_15826, n23634);
  not g39091 (n_15827, n23644);
  and g39092 (n23645, n_15826, n_15827);
  not g39093 (n_15828, n23645);
  and g39094 (n23646, \asqrt[30] , n_15828);
  and g39098 (n23650, n_15320, n_15319);
  and g39099 (n23651, \asqrt[2] , n23650);
  not g39100 (n_15829, n23651);
  and g39101 (n23652, n_15318, n_15829);
  not g39102 (n_15830, n23649);
  not g39103 (n_15831, n23652);
  and g39104 (n23653, n_15830, n_15831);
  and g39105 (n23654, n_5322, n_15826);
  and g39106 (n23655, n_15827, n23654);
  not g39107 (n_15832, n23653);
  not g39108 (n_15833, n23655);
  and g39109 (n23656, n_15832, n_15833);
  not g39110 (n_15834, n23646);
  not g39111 (n_15835, n23656);
  and g39112 (n23657, n_15834, n_15835);
  not g39113 (n_15836, n23657);
  and g39114 (n23658, \asqrt[31] , n_15836);
  and g39118 (n23662, n_15328, n_15327);
  and g39119 (n23663, \asqrt[2] , n23662);
  not g39120 (n_15837, n23663);
  and g39121 (n23664, n_15326, n_15837);
  not g39122 (n_15838, n23661);
  not g39123 (n_15839, n23664);
  and g39124 (n23665, n_15838, n_15839);
  and g39125 (n23666, n_5034, n_15834);
  and g39126 (n23667, n_15835, n23666);
  not g39127 (n_15840, n23665);
  not g39128 (n_15841, n23667);
  and g39129 (n23668, n_15840, n_15841);
  not g39130 (n_15842, n23658);
  not g39131 (n_15843, n23668);
  and g39132 (n23669, n_15842, n_15843);
  not g39133 (n_15844, n23669);
  and g39134 (n23670, \asqrt[32] , n_15844);
  and g39138 (n23674, n_15336, n_15335);
  and g39139 (n23675, \asqrt[2] , n23674);
  not g39140 (n_15845, n23675);
  and g39141 (n23676, n_15334, n_15845);
  not g39142 (n_15846, n23673);
  not g39143 (n_15847, n23676);
  and g39144 (n23677, n_15846, n_15847);
  and g39145 (n23678, n_4754, n_15842);
  and g39146 (n23679, n_15843, n23678);
  not g39147 (n_15848, n23677);
  not g39148 (n_15849, n23679);
  and g39149 (n23680, n_15848, n_15849);
  not g39150 (n_15850, n23670);
  not g39151 (n_15851, n23680);
  and g39152 (n23681, n_15850, n_15851);
  not g39153 (n_15852, n23681);
  and g39154 (n23682, \asqrt[33] , n_15852);
  and g39158 (n23686, n_15344, n_15343);
  and g39159 (n23687, \asqrt[2] , n23686);
  not g39160 (n_15853, n23687);
  and g39161 (n23688, n_15342, n_15853);
  not g39162 (n_15854, n23685);
  not g39163 (n_15855, n23688);
  and g39164 (n23689, n_15854, n_15855);
  and g39165 (n23690, n_4482, n_15850);
  and g39166 (n23691, n_15851, n23690);
  not g39167 (n_15856, n23689);
  not g39168 (n_15857, n23691);
  and g39169 (n23692, n_15856, n_15857);
  not g39170 (n_15858, n23682);
  not g39171 (n_15859, n23692);
  and g39172 (n23693, n_15858, n_15859);
  not g39173 (n_15860, n23693);
  and g39174 (n23694, \asqrt[34] , n_15860);
  and g39178 (n23698, n_15352, n_15351);
  and g39179 (n23699, \asqrt[2] , n23698);
  not g39180 (n_15861, n23699);
  and g39181 (n23700, n_15350, n_15861);
  not g39182 (n_15862, n23697);
  not g39183 (n_15863, n23700);
  and g39184 (n23701, n_15862, n_15863);
  and g39185 (n23702, n_4218, n_15858);
  and g39186 (n23703, n_15859, n23702);
  not g39187 (n_15864, n23701);
  not g39188 (n_15865, n23703);
  and g39189 (n23704, n_15864, n_15865);
  not g39190 (n_15866, n23694);
  not g39191 (n_15867, n23704);
  and g39192 (n23705, n_15866, n_15867);
  not g39193 (n_15868, n23705);
  and g39194 (n23706, \asqrt[35] , n_15868);
  and g39198 (n23710, n_15360, n_15359);
  and g39199 (n23711, \asqrt[2] , n23710);
  not g39200 (n_15869, n23711);
  and g39201 (n23712, n_15358, n_15869);
  not g39202 (n_15870, n23709);
  not g39203 (n_15871, n23712);
  and g39204 (n23713, n_15870, n_15871);
  and g39205 (n23714, n_3962, n_15866);
  and g39206 (n23715, n_15867, n23714);
  not g39207 (n_15872, n23713);
  not g39208 (n_15873, n23715);
  and g39209 (n23716, n_15872, n_15873);
  not g39210 (n_15874, n23706);
  not g39211 (n_15875, n23716);
  and g39212 (n23717, n_15874, n_15875);
  not g39213 (n_15876, n23717);
  and g39214 (n23718, \asqrt[36] , n_15876);
  and g39218 (n23722, n_15368, n_15367);
  and g39219 (n23723, \asqrt[2] , n23722);
  not g39220 (n_15877, n23723);
  and g39221 (n23724, n_15366, n_15877);
  not g39222 (n_15878, n23721);
  not g39223 (n_15879, n23724);
  and g39224 (n23725, n_15878, n_15879);
  and g39225 (n23726, n_3714, n_15874);
  and g39226 (n23727, n_15875, n23726);
  not g39227 (n_15880, n23725);
  not g39228 (n_15881, n23727);
  and g39229 (n23728, n_15880, n_15881);
  not g39230 (n_15882, n23718);
  not g39231 (n_15883, n23728);
  and g39232 (n23729, n_15882, n_15883);
  not g39233 (n_15884, n23729);
  and g39234 (n23730, \asqrt[37] , n_15884);
  and g39238 (n23734, n_15376, n_15375);
  and g39239 (n23735, \asqrt[2] , n23734);
  not g39240 (n_15885, n23735);
  and g39241 (n23736, n_15374, n_15885);
  not g39242 (n_15886, n23733);
  not g39243 (n_15887, n23736);
  and g39244 (n23737, n_15886, n_15887);
  and g39245 (n23738, n_3474, n_15882);
  and g39246 (n23739, n_15883, n23738);
  not g39247 (n_15888, n23737);
  not g39248 (n_15889, n23739);
  and g39249 (n23740, n_15888, n_15889);
  not g39250 (n_15890, n23730);
  not g39251 (n_15891, n23740);
  and g39252 (n23741, n_15890, n_15891);
  not g39253 (n_15892, n23741);
  and g39254 (n23742, \asqrt[38] , n_15892);
  and g39258 (n23746, n_15384, n_15383);
  and g39259 (n23747, \asqrt[2] , n23746);
  not g39260 (n_15893, n23747);
  and g39261 (n23748, n_15382, n_15893);
  not g39262 (n_15894, n23745);
  not g39263 (n_15895, n23748);
  and g39264 (n23749, n_15894, n_15895);
  and g39265 (n23750, n_3242, n_15890);
  and g39266 (n23751, n_15891, n23750);
  not g39267 (n_15896, n23749);
  not g39268 (n_15897, n23751);
  and g39269 (n23752, n_15896, n_15897);
  not g39270 (n_15898, n23742);
  not g39271 (n_15899, n23752);
  and g39272 (n23753, n_15898, n_15899);
  not g39273 (n_15900, n23753);
  and g39274 (n23754, \asqrt[39] , n_15900);
  and g39278 (n23758, n_15392, n_15391);
  and g39279 (n23759, \asqrt[2] , n23758);
  not g39280 (n_15901, n23759);
  and g39281 (n23760, n_15390, n_15901);
  not g39282 (n_15902, n23757);
  not g39283 (n_15903, n23760);
  and g39284 (n23761, n_15902, n_15903);
  and g39285 (n23762, n_3018, n_15898);
  and g39286 (n23763, n_15899, n23762);
  not g39287 (n_15904, n23761);
  not g39288 (n_15905, n23763);
  and g39289 (n23764, n_15904, n_15905);
  not g39290 (n_15906, n23754);
  not g39291 (n_15907, n23764);
  and g39292 (n23765, n_15906, n_15907);
  not g39293 (n_15908, n23765);
  and g39294 (n23766, \asqrt[40] , n_15908);
  and g39298 (n23770, n_15400, n_15399);
  and g39299 (n23771, \asqrt[2] , n23770);
  not g39300 (n_15909, n23771);
  and g39301 (n23772, n_15398, n_15909);
  not g39302 (n_15910, n23769);
  not g39303 (n_15911, n23772);
  and g39304 (n23773, n_15910, n_15911);
  and g39305 (n23774, n_2802, n_15906);
  and g39306 (n23775, n_15907, n23774);
  not g39307 (n_15912, n23773);
  not g39308 (n_15913, n23775);
  and g39309 (n23776, n_15912, n_15913);
  not g39310 (n_15914, n23766);
  not g39311 (n_15915, n23776);
  and g39312 (n23777, n_15914, n_15915);
  not g39313 (n_15916, n23777);
  and g39314 (n23778, \asqrt[41] , n_15916);
  and g39318 (n23782, n_15408, n_15407);
  and g39319 (n23783, \asqrt[2] , n23782);
  not g39320 (n_15917, n23783);
  and g39321 (n23784, n_15406, n_15917);
  not g39322 (n_15918, n23781);
  not g39323 (n_15919, n23784);
  and g39324 (n23785, n_15918, n_15919);
  and g39325 (n23786, n_2594, n_15914);
  and g39326 (n23787, n_15915, n23786);
  not g39327 (n_15920, n23785);
  not g39328 (n_15921, n23787);
  and g39329 (n23788, n_15920, n_15921);
  not g39330 (n_15922, n23778);
  not g39331 (n_15923, n23788);
  and g39332 (n23789, n_15922, n_15923);
  not g39333 (n_15924, n23789);
  and g39334 (n23790, \asqrt[42] , n_15924);
  and g39338 (n23794, n_15416, n_15415);
  and g39339 (n23795, \asqrt[2] , n23794);
  not g39340 (n_15925, n23795);
  and g39341 (n23796, n_15414, n_15925);
  not g39342 (n_15926, n23793);
  not g39343 (n_15927, n23796);
  and g39344 (n23797, n_15926, n_15927);
  and g39345 (n23798, n_2394, n_15922);
  and g39346 (n23799, n_15923, n23798);
  not g39347 (n_15928, n23797);
  not g39348 (n_15929, n23799);
  and g39349 (n23800, n_15928, n_15929);
  not g39350 (n_15930, n23790);
  not g39351 (n_15931, n23800);
  and g39352 (n23801, n_15930, n_15931);
  not g39353 (n_15932, n23801);
  and g39354 (n23802, \asqrt[43] , n_15932);
  and g39358 (n23806, n_15424, n_15423);
  and g39359 (n23807, \asqrt[2] , n23806);
  not g39360 (n_15933, n23807);
  and g39361 (n23808, n_15422, n_15933);
  not g39362 (n_15934, n23805);
  not g39363 (n_15935, n23808);
  and g39364 (n23809, n_15934, n_15935);
  and g39365 (n23810, n_2202, n_15930);
  and g39366 (n23811, n_15931, n23810);
  not g39367 (n_15936, n23809);
  not g39368 (n_15937, n23811);
  and g39369 (n23812, n_15936, n_15937);
  not g39370 (n_15938, n23802);
  not g39371 (n_15939, n23812);
  and g39372 (n23813, n_15938, n_15939);
  not g39373 (n_15940, n23813);
  and g39374 (n23814, \asqrt[44] , n_15940);
  and g39378 (n23818, n_15432, n_15431);
  and g39379 (n23819, \asqrt[2] , n23818);
  not g39380 (n_15941, n23819);
  and g39381 (n23820, n_15430, n_15941);
  not g39382 (n_15942, n23817);
  not g39383 (n_15943, n23820);
  and g39384 (n23821, n_15942, n_15943);
  and g39385 (n23822, n_2018, n_15938);
  and g39386 (n23823, n_15939, n23822);
  not g39387 (n_15944, n23821);
  not g39388 (n_15945, n23823);
  and g39389 (n23824, n_15944, n_15945);
  not g39390 (n_15946, n23814);
  not g39391 (n_15947, n23824);
  and g39392 (n23825, n_15946, n_15947);
  not g39393 (n_15948, n23825);
  and g39394 (n23826, \asqrt[45] , n_15948);
  and g39398 (n23830, n_15440, n_15439);
  and g39399 (n23831, \asqrt[2] , n23830);
  not g39400 (n_15949, n23831);
  and g39401 (n23832, n_15438, n_15949);
  not g39402 (n_15950, n23829);
  not g39403 (n_15951, n23832);
  and g39404 (n23833, n_15950, n_15951);
  and g39405 (n23834, n_1842, n_15946);
  and g39406 (n23835, n_15947, n23834);
  not g39407 (n_15952, n23833);
  not g39408 (n_15953, n23835);
  and g39409 (n23836, n_15952, n_15953);
  not g39410 (n_15954, n23826);
  not g39411 (n_15955, n23836);
  and g39412 (n23837, n_15954, n_15955);
  not g39413 (n_15956, n23837);
  and g39414 (n23838, \asqrt[46] , n_15956);
  and g39418 (n23842, n_15448, n_15447);
  and g39419 (n23843, \asqrt[2] , n23842);
  not g39420 (n_15957, n23843);
  and g39421 (n23844, n_15446, n_15957);
  not g39422 (n_15958, n23841);
  not g39423 (n_15959, n23844);
  and g39424 (n23845, n_15958, n_15959);
  and g39425 (n23846, n_1674, n_15954);
  and g39426 (n23847, n_15955, n23846);
  not g39427 (n_15960, n23845);
  not g39428 (n_15961, n23847);
  and g39429 (n23848, n_15960, n_15961);
  not g39430 (n_15962, n23838);
  not g39431 (n_15963, n23848);
  and g39432 (n23849, n_15962, n_15963);
  not g39433 (n_15964, n23849);
  and g39434 (n23850, \asqrt[47] , n_15964);
  and g39438 (n23854, n_15456, n_15455);
  and g39439 (n23855, \asqrt[2] , n23854);
  not g39440 (n_15965, n23855);
  and g39441 (n23856, n_15454, n_15965);
  not g39442 (n_15966, n23853);
  not g39443 (n_15967, n23856);
  and g39444 (n23857, n_15966, n_15967);
  and g39445 (n23858, n_1514, n_15962);
  and g39446 (n23859, n_15963, n23858);
  not g39447 (n_15968, n23857);
  not g39448 (n_15969, n23859);
  and g39449 (n23860, n_15968, n_15969);
  not g39450 (n_15970, n23850);
  not g39451 (n_15971, n23860);
  and g39452 (n23861, n_15970, n_15971);
  not g39453 (n_15972, n23861);
  and g39454 (n23862, \asqrt[48] , n_15972);
  and g39458 (n23866, n_15464, n_15463);
  and g39459 (n23867, \asqrt[2] , n23866);
  not g39460 (n_15973, n23867);
  and g39461 (n23868, n_15462, n_15973);
  not g39462 (n_15974, n23865);
  not g39463 (n_15975, n23868);
  and g39464 (n23869, n_15974, n_15975);
  and g39465 (n23870, n_1362, n_15970);
  and g39466 (n23871, n_15971, n23870);
  not g39467 (n_15976, n23869);
  not g39468 (n_15977, n23871);
  and g39469 (n23872, n_15976, n_15977);
  not g39470 (n_15978, n23862);
  not g39471 (n_15979, n23872);
  and g39472 (n23873, n_15978, n_15979);
  not g39473 (n_15980, n23873);
  and g39474 (n23874, \asqrt[49] , n_15980);
  and g39478 (n23878, n_15472, n_15471);
  and g39479 (n23879, \asqrt[2] , n23878);
  not g39480 (n_15981, n23879);
  and g39481 (n23880, n_15470, n_15981);
  not g39482 (n_15982, n23877);
  not g39483 (n_15983, n23880);
  and g39484 (n23881, n_15982, n_15983);
  and g39485 (n23882, n_1218, n_15978);
  and g39486 (n23883, n_15979, n23882);
  not g39487 (n_15984, n23881);
  not g39488 (n_15985, n23883);
  and g39489 (n23884, n_15984, n_15985);
  not g39490 (n_15986, n23874);
  not g39491 (n_15987, n23884);
  and g39492 (n23885, n_15986, n_15987);
  not g39493 (n_15988, n23885);
  and g39494 (n23886, \asqrt[50] , n_15988);
  and g39498 (n23890, n_15480, n_15479);
  and g39499 (n23891, \asqrt[2] , n23890);
  not g39500 (n_15989, n23891);
  and g39501 (n23892, n_15478, n_15989);
  not g39502 (n_15990, n23889);
  not g39503 (n_15991, n23892);
  and g39504 (n23893, n_15990, n_15991);
  and g39505 (n23894, n_1082, n_15986);
  and g39506 (n23895, n_15987, n23894);
  not g39507 (n_15992, n23893);
  not g39508 (n_15993, n23895);
  and g39509 (n23896, n_15992, n_15993);
  not g39510 (n_15994, n23886);
  not g39511 (n_15995, n23896);
  and g39512 (n23897, n_15994, n_15995);
  not g39513 (n_15996, n23897);
  and g39514 (n23898, \asqrt[51] , n_15996);
  and g39518 (n23902, n_15488, n_15487);
  and g39519 (n23903, \asqrt[2] , n23902);
  not g39520 (n_15997, n23903);
  and g39521 (n23904, n_15486, n_15997);
  not g39522 (n_15998, n23901);
  not g39523 (n_15999, n23904);
  and g39524 (n23905, n_15998, n_15999);
  and g39525 (n23906, n_954, n_15994);
  and g39526 (n23907, n_15995, n23906);
  not g39527 (n_16000, n23905);
  not g39528 (n_16001, n23907);
  and g39529 (n23908, n_16000, n_16001);
  not g39530 (n_16002, n23898);
  not g39531 (n_16003, n23908);
  and g39532 (n23909, n_16002, n_16003);
  not g39533 (n_16004, n23909);
  and g39534 (n23910, \asqrt[52] , n_16004);
  and g39538 (n23914, n_15496, n_15495);
  and g39539 (n23915, \asqrt[2] , n23914);
  not g39540 (n_16005, n23915);
  and g39541 (n23916, n_15494, n_16005);
  not g39542 (n_16006, n23913);
  not g39543 (n_16007, n23916);
  and g39544 (n23917, n_16006, n_16007);
  and g39545 (n23918, n_834, n_16002);
  and g39546 (n23919, n_16003, n23918);
  not g39547 (n_16008, n23917);
  not g39548 (n_16009, n23919);
  and g39549 (n23920, n_16008, n_16009);
  not g39550 (n_16010, n23910);
  not g39551 (n_16011, n23920);
  and g39552 (n23921, n_16010, n_16011);
  not g39553 (n_16012, n23921);
  and g39554 (n23922, \asqrt[53] , n_16012);
  and g39558 (n23926, n_15504, n_15503);
  and g39559 (n23927, \asqrt[2] , n23926);
  not g39560 (n_16013, n23927);
  and g39561 (n23928, n_15502, n_16013);
  not g39562 (n_16014, n23925);
  not g39563 (n_16015, n23928);
  and g39564 (n23929, n_16014, n_16015);
  and g39565 (n23930, n_722, n_16010);
  and g39566 (n23931, n_16011, n23930);
  not g39567 (n_16016, n23929);
  not g39568 (n_16017, n23931);
  and g39569 (n23932, n_16016, n_16017);
  not g39570 (n_16018, n23922);
  not g39571 (n_16019, n23932);
  and g39572 (n23933, n_16018, n_16019);
  not g39573 (n_16020, n23933);
  and g39574 (n23934, \asqrt[54] , n_16020);
  and g39578 (n23938, n_15512, n_15511);
  and g39579 (n23939, \asqrt[2] , n23938);
  not g39580 (n_16021, n23939);
  and g39581 (n23940, n_15510, n_16021);
  not g39582 (n_16022, n23937);
  not g39583 (n_16023, n23940);
  and g39584 (n23941, n_16022, n_16023);
  and g39585 (n23942, n_618, n_16018);
  and g39586 (n23943, n_16019, n23942);
  not g39587 (n_16024, n23941);
  not g39588 (n_16025, n23943);
  and g39589 (n23944, n_16024, n_16025);
  not g39590 (n_16026, n23934);
  not g39591 (n_16027, n23944);
  and g39592 (n23945, n_16026, n_16027);
  not g39593 (n_16028, n23945);
  and g39594 (n23946, \asqrt[55] , n_16028);
  and g39598 (n23950, n_15520, n_15519);
  and g39599 (n23951, \asqrt[2] , n23950);
  not g39600 (n_16029, n23951);
  and g39601 (n23952, n_15518, n_16029);
  not g39602 (n_16030, n23949);
  not g39603 (n_16031, n23952);
  and g39604 (n23953, n_16030, n_16031);
  and g39605 (n23954, n_522, n_16026);
  and g39606 (n23955, n_16027, n23954);
  not g39607 (n_16032, n23953);
  not g39608 (n_16033, n23955);
  and g39609 (n23956, n_16032, n_16033);
  not g39610 (n_16034, n23946);
  not g39611 (n_16035, n23956);
  and g39612 (n23957, n_16034, n_16035);
  not g39613 (n_16036, n23957);
  and g39614 (n23958, \asqrt[56] , n_16036);
  and g39618 (n23962, n_15528, n_15527);
  and g39619 (n23963, \asqrt[2] , n23962);
  not g39620 (n_16037, n23963);
  and g39621 (n23964, n_15526, n_16037);
  not g39622 (n_16038, n23961);
  not g39623 (n_16039, n23964);
  and g39624 (n23965, n_16038, n_16039);
  and g39625 (n23966, n_434, n_16034);
  and g39626 (n23967, n_16035, n23966);
  not g39627 (n_16040, n23965);
  not g39628 (n_16041, n23967);
  and g39629 (n23968, n_16040, n_16041);
  not g39630 (n_16042, n23958);
  not g39631 (n_16043, n23968);
  and g39632 (n23969, n_16042, n_16043);
  not g39633 (n_16044, n23969);
  and g39634 (n23970, \asqrt[57] , n_16044);
  and g39638 (n23974, n_15536, n_15535);
  and g39639 (n23975, \asqrt[2] , n23974);
  not g39640 (n_16045, n23975);
  and g39641 (n23976, n_15534, n_16045);
  not g39642 (n_16046, n23973);
  not g39643 (n_16047, n23976);
  and g39644 (n23977, n_16046, n_16047);
  and g39645 (n23978, n_354, n_16042);
  and g39646 (n23979, n_16043, n23978);
  not g39647 (n_16048, n23977);
  not g39648 (n_16049, n23979);
  and g39649 (n23980, n_16048, n_16049);
  not g39650 (n_16050, n23970);
  not g39651 (n_16051, n23980);
  and g39652 (n23981, n_16050, n_16051);
  not g39653 (n_16052, n23981);
  and g39654 (n23982, \asqrt[58] , n_16052);
  and g39658 (n23986, n_15544, n_15543);
  and g39659 (n23987, \asqrt[2] , n23986);
  not g39660 (n_16053, n23987);
  and g39661 (n23988, n_15542, n_16053);
  not g39662 (n_16054, n23985);
  not g39663 (n_16055, n23988);
  and g39664 (n23989, n_16054, n_16055);
  and g39665 (n23990, n_282, n_16050);
  and g39666 (n23991, n_16051, n23990);
  not g39667 (n_16056, n23989);
  not g39668 (n_16057, n23991);
  and g39669 (n23992, n_16056, n_16057);
  not g39670 (n_16058, n23982);
  not g39671 (n_16059, n23992);
  and g39672 (n23993, n_16058, n_16059);
  not g39673 (n_16060, n23993);
  and g39674 (n23994, \asqrt[59] , n_16060);
  and g39678 (n23998, n_15552, n_15551);
  and g39679 (n23999, \asqrt[2] , n23998);
  not g39680 (n_16061, n23999);
  and g39681 (n24000, n_15550, n_16061);
  not g39682 (n_16062, n23997);
  not g39683 (n_16063, n24000);
  and g39684 (n24001, n_16062, n_16063);
  and g39685 (n24002, n_218, n_16058);
  and g39686 (n24003, n_16059, n24002);
  not g39687 (n_16064, n24001);
  not g39688 (n_16065, n24003);
  and g39689 (n24004, n_16064, n_16065);
  not g39690 (n_16066, n23994);
  not g39691 (n_16067, n24004);
  and g39692 (n24005, n_16066, n_16067);
  not g39693 (n_16068, n24005);
  and g39694 (n24006, \asqrt[60] , n_16068);
  and g39698 (n24010, n_15560, n_15559);
  and g39699 (n24011, \asqrt[2] , n24010);
  not g39700 (n_16069, n24011);
  and g39701 (n24012, n_15558, n_16069);
  not g39702 (n_16070, n24009);
  not g39703 (n_16071, n24012);
  and g39704 (n24013, n_16070, n_16071);
  and g39705 (n24014, n_162, n_16066);
  and g39706 (n24015, n_16067, n24014);
  not g39707 (n_16072, n24013);
  not g39708 (n_16073, n24015);
  and g39709 (n24016, n_16072, n_16073);
  not g39710 (n_16074, n24006);
  not g39711 (n_16075, n24016);
  and g39712 (n24017, n_16074, n_16075);
  not g39713 (n_16076, n24017);
  and g39714 (n24018, \asqrt[61] , n_16076);
  and g39715 (n24019, n_115, n_16074);
  and g39716 (n24020, n_16075, n24019);
  not g39717 (n_16077, n23318);
  not g39718 (n_16078, n24020);
  and g39719 (n24021, n_16077, n_16078);
  not g39720 (n_16079, n24018);
  not g39721 (n_16080, n24021);
  and g39722 (n24022, n_16079, n_16080);
  not g39723 (n_16081, n24022);
  and g39724 (n24023, \asqrt[62] , n_16081);
  and g39728 (n24027, n_15576, n_15575);
  and g39729 (n24028, \asqrt[2] , n24027);
  not g39730 (n_16082, n24028);
  and g39731 (n24029, n_15574, n_16082);
  not g39732 (n_16083, n24026);
  not g39733 (n_16084, n24029);
  and g39734 (n24030, n_16083, n_16084);
  and g39735 (n24031, n_76, n_16079);
  and g39736 (n24032, n_16080, n24031);
  not g39737 (n_16085, n24030);
  not g39738 (n_16086, n24032);
  and g39739 (n24033, n_16085, n_16086);
  not g39740 (n_16087, n24023);
  not g39741 (n_16088, n24033);
  and g39742 (n24034, n_16087, n_16088);
  and g39746 (n24038, n_15584, n_15582);
  and g39747 (n24039, \asqrt[2] , n24038);
  not g39748 (n_16089, n24039);
  and g39749 (n24040, n_15583, n_16089);
  not g39750 (n_16090, n24037);
  not g39751 (n_16091, n24040);
  and g39752 (n24041, n_16090, n_16091);
  and g39753 (n24042, n_15591, n_15590);
  and g39754 (n24043, \asqrt[2] , n24042);
  not g39757 (n_16093, n24041);
  not g39759 (n_16094, n24034);
  not g39761 (n_16095, n24046);
  and g39762 (n24047, n_21, n_16095);
  and g39763 (n24048, n_16087, n24041);
  and g39764 (n24049, n_16088, n24048);
  and g39765 (n24050, n_15590, \asqrt[2] );
  not g39766 (n_16096, n24050);
  and g39767 (n24051, n23290, n_16096);
  not g39768 (n_16097, n24042);
  and g39769 (n24052, \asqrt[63] , n_16097);
  not g39770 (n_16098, n24051);
  and g39771 (n24053, n_16098, n24052);
  not g39772 (n_16099, n24049);
  not g39773 (n_16100, n24053);
  and g39774 (n24054, n_16099, n_16100);
  not g39775 (n_16101, n24054);
  or g39776 (\asqrt[1] , n24047, n_16101);
  and g39777 (n24056, n_16079, n_16078);
  and g39778 (n24057, \asqrt[1] , n24056);
  not g39779 (n_16103, n24057);
  and g39780 (n24058, n_16077, n_16103);
  not g39784 (n_16104, n24058);
  not g39785 (n_16105, n24061);
  and g39786 (n24062, n_16104, n_16105);
  and g39787 (n24063, n_16066, n_16065);
  and g39788 (n24064, \asqrt[1] , n24063);
  not g39789 (n_16106, n24064);
  and g39790 (n24065, n_16064, n_16106);
  not g39794 (n_16107, n24065);
  not g39795 (n_16108, n24068);
  and g39796 (n24069, n_16107, n_16108);
  and g39797 (n24070, n_16050, n_16049);
  and g39798 (n24071, \asqrt[1] , n24070);
  not g39799 (n_16109, n24071);
  and g39800 (n24072, n_16048, n_16109);
  not g39804 (n_16110, n24072);
  not g39805 (n_16111, n24075);
  and g39806 (n24076, n_16110, n_16111);
  and g39807 (n24077, n_16034, n_16033);
  and g39808 (n24078, \asqrt[1] , n24077);
  not g39809 (n_16112, n24078);
  and g39810 (n24079, n_16032, n_16112);
  not g39814 (n_16113, n24079);
  not g39815 (n_16114, n24082);
  and g39816 (n24083, n_16113, n_16114);
  and g39817 (n24084, n_16018, n_16017);
  and g39818 (n24085, \asqrt[1] , n24084);
  not g39819 (n_16115, n24085);
  and g39820 (n24086, n_16016, n_16115);
  not g39824 (n_16116, n24086);
  not g39825 (n_16117, n24089);
  and g39826 (n24090, n_16116, n_16117);
  and g39827 (n24091, n_16002, n_16001);
  and g39828 (n24092, \asqrt[1] , n24091);
  not g39829 (n_16118, n24092);
  and g39830 (n24093, n_16000, n_16118);
  not g39834 (n_16119, n24093);
  not g39835 (n_16120, n24096);
  and g39836 (n24097, n_16119, n_16120);
  and g39837 (n24098, n_15986, n_15985);
  and g39838 (n24099, \asqrt[1] , n24098);
  not g39839 (n_16121, n24099);
  and g39840 (n24100, n_15984, n_16121);
  not g39844 (n_16122, n24100);
  not g39845 (n_16123, n24103);
  and g39846 (n24104, n_16122, n_16123);
  and g39847 (n24105, n_15970, n_15969);
  and g39848 (n24106, \asqrt[1] , n24105);
  not g39849 (n_16124, n24106);
  and g39850 (n24107, n_15968, n_16124);
  not g39854 (n_16125, n24107);
  not g39855 (n_16126, n24110);
  and g39856 (n24111, n_16125, n_16126);
  and g39857 (n24112, n_15954, n_15953);
  and g39858 (n24113, \asqrt[1] , n24112);
  not g39859 (n_16127, n24113);
  and g39860 (n24114, n_15952, n_16127);
  not g39864 (n_16128, n24114);
  not g39865 (n_16129, n24117);
  and g39866 (n24118, n_16128, n_16129);
  and g39867 (n24119, n_15938, n_15937);
  and g39868 (n24120, \asqrt[1] , n24119);
  not g39869 (n_16130, n24120);
  and g39870 (n24121, n_15936, n_16130);
  not g39874 (n_16131, n24121);
  not g39875 (n_16132, n24124);
  and g39876 (n24125, n_16131, n_16132);
  and g39877 (n24126, n_15922, n_15921);
  and g39878 (n24127, \asqrt[1] , n24126);
  not g39879 (n_16133, n24127);
  and g39880 (n24128, n_15920, n_16133);
  not g39884 (n_16134, n24128);
  not g39885 (n_16135, n24131);
  and g39886 (n24132, n_16134, n_16135);
  and g39887 (n24133, n_15906, n_15905);
  and g39888 (n24134, \asqrt[1] , n24133);
  not g39889 (n_16136, n24134);
  and g39890 (n24135, n_15904, n_16136);
  not g39894 (n_16137, n24135);
  not g39895 (n_16138, n24138);
  and g39896 (n24139, n_16137, n_16138);
  and g39897 (n24140, n_15890, n_15889);
  and g39898 (n24141, \asqrt[1] , n24140);
  not g39899 (n_16139, n24141);
  and g39900 (n24142, n_15888, n_16139);
  not g39904 (n_16140, n24142);
  not g39905 (n_16141, n24145);
  and g39906 (n24146, n_16140, n_16141);
  and g39907 (n24147, n_15874, n_15873);
  and g39908 (n24148, \asqrt[1] , n24147);
  not g39909 (n_16142, n24148);
  and g39910 (n24149, n_15872, n_16142);
  not g39914 (n_16143, n24149);
  not g39915 (n_16144, n24152);
  and g39916 (n24153, n_16143, n_16144);
  and g39917 (n24154, n_15858, n_15857);
  and g39918 (n24155, \asqrt[1] , n24154);
  not g39919 (n_16145, n24155);
  and g39920 (n24156, n_15856, n_16145);
  not g39924 (n_16146, n24156);
  not g39925 (n_16147, n24159);
  and g39926 (n24160, n_16146, n_16147);
  and g39927 (n24161, n_15842, n_15841);
  and g39928 (n24162, \asqrt[1] , n24161);
  not g39929 (n_16148, n24162);
  and g39930 (n24163, n_15840, n_16148);
  not g39934 (n_16149, n24163);
  not g39935 (n_16150, n24166);
  and g39936 (n24167, n_16149, n_16150);
  and g39937 (n24168, n_15826, n_15825);
  and g39938 (n24169, \asqrt[1] , n24168);
  not g39939 (n_16151, n24169);
  and g39940 (n24170, n_15824, n_16151);
  not g39944 (n_16152, n24170);
  not g39945 (n_16153, n24173);
  and g39946 (n24174, n_16152, n_16153);
  and g39947 (n24175, n_15810, n_15809);
  and g39948 (n24176, \asqrt[1] , n24175);
  not g39949 (n_16154, n24176);
  and g39950 (n24177, n_15808, n_16154);
  not g39954 (n_16155, n24177);
  not g39955 (n_16156, n24180);
  and g39956 (n24181, n_16155, n_16156);
  and g39957 (n24182, n_15794, n_15793);
  and g39958 (n24183, \asqrt[1] , n24182);
  not g39959 (n_16157, n24183);
  and g39960 (n24184, n_15792, n_16157);
  not g39964 (n_16158, n24184);
  not g39965 (n_16159, n24187);
  and g39966 (n24188, n_16158, n_16159);
  and g39967 (n24189, n_15778, n_15777);
  and g39968 (n24190, \asqrt[1] , n24189);
  not g39969 (n_16160, n24190);
  and g39970 (n24191, n_15776, n_16160);
  not g39974 (n_16161, n24191);
  not g39975 (n_16162, n24194);
  and g39976 (n24195, n_16161, n_16162);
  and g39977 (n24196, n_15762, n_15761);
  and g39978 (n24197, \asqrt[1] , n24196);
  not g39979 (n_16163, n24197);
  and g39980 (n24198, n_15760, n_16163);
  not g39984 (n_16164, n24198);
  not g39985 (n_16165, n24201);
  and g39986 (n24202, n_16164, n_16165);
  and g39987 (n24203, n_15746, n_15745);
  and g39988 (n24204, \asqrt[1] , n24203);
  not g39989 (n_16166, n24204);
  and g39990 (n24205, n_15744, n_16166);
  not g39994 (n_16167, n24205);
  not g39995 (n_16168, n24208);
  and g39996 (n24209, n_16167, n_16168);
  and g39997 (n24210, n_15730, n_15729);
  and g39998 (n24211, \asqrt[1] , n24210);
  not g39999 (n_16169, n24211);
  and g40000 (n24212, n_15728, n_16169);
  not g40004 (n_16170, n24212);
  not g40005 (n_16171, n24215);
  and g40006 (n24216, n_16170, n_16171);
  and g40007 (n24217, n_15714, n_15713);
  and g40008 (n24218, \asqrt[1] , n24217);
  not g40009 (n_16172, n24218);
  and g40010 (n24219, n_15712, n_16172);
  not g40014 (n_16173, n24219);
  not g40015 (n_16174, n24222);
  and g40016 (n24223, n_16173, n_16174);
  and g40017 (n24224, n_15698, n_15697);
  and g40018 (n24225, \asqrt[1] , n24224);
  not g40019 (n_16175, n24225);
  and g40020 (n24226, n_15696, n_16175);
  not g40024 (n_16176, n24226);
  not g40025 (n_16177, n24229);
  and g40026 (n24230, n_16176, n_16177);
  and g40027 (n24231, n_15682, n_15681);
  and g40028 (n24232, \asqrt[1] , n24231);
  not g40029 (n_16178, n24232);
  and g40030 (n24233, n_15680, n_16178);
  not g40034 (n_16179, n24233);
  not g40035 (n_16180, n24236);
  and g40036 (n24237, n_16179, n_16180);
  and g40037 (n24238, n_15666, n_15665);
  and g40038 (n24239, \asqrt[1] , n24238);
  not g40039 (n_16181, n24239);
  and g40040 (n24240, n_15664, n_16181);
  not g40044 (n_16182, n24240);
  not g40045 (n_16183, n24243);
  and g40046 (n24244, n_16182, n_16183);
  and g40047 (n24245, n_15650, n_15649);
  and g40048 (n24246, \asqrt[1] , n24245);
  not g40049 (n_16184, n24246);
  and g40050 (n24247, n_15648, n_16184);
  not g40054 (n_16185, n24247);
  not g40055 (n_16186, n24250);
  and g40056 (n24251, n_16185, n_16186);
  and g40060 (n24255, n_15634, n_15633);
  and g40061 (n24256, \asqrt[1] , n24255);
  not g40062 (n_16187, n24256);
  and g40063 (n24257, n_15632, n_16187);
  not g40064 (n_16188, n24254);
  not g40065 (n_16189, n24257);
  and g40066 (n24258, n_16188, n_16189);
  and g40067 (n24259, n_15614, n_15613);
  not g40068 (n_16190, n23331);
  and g40069 (n24260, n_16190, n24259);
  and g40070 (n24261, \asqrt[1] , n24260);
  and g40071 (n24262, \asqrt[1] , n24259);
  not g40072 (n_16191, n24262);
  and g40073 (n24263, n23331, n_16191);
  not g40074 (n_16192, n24261);
  not g40075 (n_16193, n24263);
  and g40076 (n24264, n_16192, n_16193);
  and g40077 (n24265, n23320, \asqrt[1] );
  not g40080 (n_16194, n24047);
  not g40082 (n_16195, n24265);
  not g40083 (n_16196, n24268);
  and g40084 (n24269, n_16195, n_16196);
  not g40085 (n_16197, n24269);
  and g40086 (n24270, \a[4] , n_16197);
  and g40087 (n24271, n_15107, n_16196);
  and g40088 (n24272, n_16195, n24271);
  not g40089 (n_16198, n24270);
  not g40090 (n_16199, n24272);
  and g40091 (n24273, n_16198, n_16199);
  and g40092 (n24274, n_15605, \asqrt[1] );
  not g40093 (n_16200, n24274);
  and g40094 (n24275, \a[3] , n_16200);
  not g40095 (n_16203, \a[0] );
  not g40096 (n_16204, \a[1] );
  and g40097 (n24276, n_16203, n_16204);
  not g40098 (n_16205, n24276);
  and g40099 (n24277, n_15605, n_16205);
  not g40103 (n_16206, n24277);
  not g40104 (n_16207, n24280);
  and g40105 (n24281, n_16206, n_16207);
  and g40106 (n24282, n_16195, n24281);
  not g40107 (n_16208, n24275);
  and g40108 (n24283, n_16208, n24282);
  not g40109 (n_16209, \asqrt[2] );
  not g40110 (n_16210, n24283);
  and g40111 (n24284, n_16209, n_16210);
  and g40112 (n24285, n_16195, n_16208);
  not g40113 (n_16211, n24281);
  not g40114 (n_16212, n24285);
  and g40115 (n24286, n_16211, n_16212);
  not g40116 (n_16213, n24284);
  not g40117 (n_16214, n24286);
  and g40118 (n24287, n_16213, n_16214);
  not g40119 (n_16215, n24273);
  and g40120 (n24288, n_16215, n24287);
  not g40121 (n_16216, \asqrt[3] );
  not g40122 (n_16217, n24288);
  and g40123 (n24289, n_16216, n_16217);
  not g40124 (n_16218, n24287);
  and g40125 (n24290, n24273, n_16218);
  not g40126 (n_16219, n24289);
  not g40127 (n_16220, n24290);
  and g40128 (n24291, n_16219, n_16220);
  not g40129 (n_16221, n24291);
  and g40130 (n24292, n24264, n_16221);
  not g40131 (n_16222, n24264);
  and g40132 (n24293, n_16222, n_16220);
  and g40133 (n24294, n_16219, n24293);
  not g40134 (n_16223, n24294);
  and g40135 (n24295, n_15617, n_16223);
  and g40136 (n24296, n_15625, n_15623);
  and g40137 (n24297, \asqrt[1] , n24296);
  not g40138 (n_16224, n24297);
  and g40139 (n24298, n_15624, n_16224);
  not g40143 (n_16225, n24298);
  not g40144 (n_16226, n24301);
  and g40145 (n24302, n_16225, n_16226);
  not g40146 (n_16227, n24295);
  not g40147 (n_16228, n24302);
  and g40148 (n24303, n_16227, n_16228);
  not g40149 (n_16229, n24292);
  and g40150 (n24304, n_16229, n24303);
  not g40151 (n_16230, n24304);
  and g40152 (n24305, n_15119, n_16230);
  and g40153 (n24306, n_16229, n_16227);
  not g40154 (n_16231, n24306);
  and g40155 (n24307, n24302, n_16231);
  not g40156 (n_16232, n24305);
  not g40157 (n_16233, n24307);
  and g40158 (n24308, n_16232, n_16233);
  not g40159 (n_16234, n24308);
  and g40160 (n24309, n24258, n_16234);
  not g40161 (n_16235, n24258);
  and g40162 (n24310, n_16235, n_16233);
  and g40163 (n24311, n_16232, n24310);
  not g40164 (n_16236, n24311);
  and g40165 (n24312, n_14632, n_16236);
  and g40166 (n24313, n_15642, n_15641);
  and g40167 (n24314, \asqrt[1] , n24313);
  not g40168 (n_16237, n24314);
  and g40169 (n24315, n_15640, n_16237);
  not g40173 (n_16238, n24315);
  not g40174 (n_16239, n24318);
  and g40175 (n24319, n_16238, n_16239);
  not g40176 (n_16240, n24312);
  not g40177 (n_16241, n24319);
  and g40178 (n24320, n_16240, n_16241);
  not g40179 (n_16242, n24309);
  and g40180 (n24321, n_16242, n24320);
  not g40181 (n_16243, n24321);
  and g40182 (n24322, n_14153, n_16243);
  and g40183 (n24323, n_16242, n_16240);
  not g40184 (n_16244, n24323);
  and g40185 (n24324, n24319, n_16244);
  not g40186 (n_16245, n24322);
  not g40187 (n_16246, n24324);
  and g40188 (n24325, n_16245, n_16246);
  not g40189 (n_16247, n24325);
  and g40190 (n24326, n24251, n_16247);
  not g40191 (n_16248, n24251);
  and g40192 (n24327, n_16248, n_16246);
  and g40193 (n24328, n_16245, n24327);
  not g40194 (n_16249, n24328);
  and g40195 (n24329, n_13682, n_16249);
  and g40196 (n24330, n_15658, n_15657);
  and g40197 (n24331, \asqrt[1] , n24330);
  not g40198 (n_16250, n24331);
  and g40199 (n24332, n_15656, n_16250);
  not g40203 (n_16251, n24332);
  not g40204 (n_16252, n24335);
  and g40205 (n24336, n_16251, n_16252);
  not g40206 (n_16253, n24329);
  not g40207 (n_16254, n24336);
  and g40208 (n24337, n_16253, n_16254);
  not g40209 (n_16255, n24326);
  and g40210 (n24338, n_16255, n24337);
  not g40211 (n_16256, n24338);
  and g40212 (n24339, n_13218, n_16256);
  and g40213 (n24340, n_16255, n_16253);
  not g40214 (n_16257, n24340);
  and g40215 (n24341, n24336, n_16257);
  not g40216 (n_16258, n24339);
  not g40217 (n_16259, n24341);
  and g40218 (n24342, n_16258, n_16259);
  not g40219 (n_16260, n24342);
  and g40220 (n24343, n24244, n_16260);
  not g40221 (n_16261, n24244);
  and g40222 (n24344, n_16261, n_16259);
  and g40223 (n24345, n_16258, n24344);
  not g40224 (n_16262, n24345);
  and g40225 (n24346, n_12762, n_16262);
  and g40226 (n24347, n_15674, n_15673);
  and g40227 (n24348, \asqrt[1] , n24347);
  not g40228 (n_16263, n24348);
  and g40229 (n24349, n_15672, n_16263);
  not g40233 (n_16264, n24349);
  not g40234 (n_16265, n24352);
  and g40235 (n24353, n_16264, n_16265);
  not g40236 (n_16266, n24346);
  not g40237 (n_16267, n24353);
  and g40238 (n24354, n_16266, n_16267);
  not g40239 (n_16268, n24343);
  and g40240 (n24355, n_16268, n24354);
  not g40241 (n_16269, n24355);
  and g40242 (n24356, n_12314, n_16269);
  and g40243 (n24357, n_16268, n_16266);
  not g40244 (n_16270, n24357);
  and g40245 (n24358, n24353, n_16270);
  not g40246 (n_16271, n24356);
  not g40247 (n_16272, n24358);
  and g40248 (n24359, n_16271, n_16272);
  not g40249 (n_16273, n24359);
  and g40250 (n24360, n24237, n_16273);
  not g40251 (n_16274, n24237);
  and g40252 (n24361, n_16274, n_16272);
  and g40253 (n24362, n_16271, n24361);
  not g40254 (n_16275, n24362);
  and g40255 (n24363, n_11874, n_16275);
  and g40256 (n24364, n_15690, n_15689);
  and g40257 (n24365, \asqrt[1] , n24364);
  not g40258 (n_16276, n24365);
  and g40259 (n24366, n_15688, n_16276);
  not g40263 (n_16277, n24366);
  not g40264 (n_16278, n24369);
  and g40265 (n24370, n_16277, n_16278);
  not g40266 (n_16279, n24363);
  not g40267 (n_16280, n24370);
  and g40268 (n24371, n_16279, n_16280);
  not g40269 (n_16281, n24360);
  and g40270 (n24372, n_16281, n24371);
  not g40271 (n_16282, n24372);
  and g40272 (n24373, n_11442, n_16282);
  and g40273 (n24374, n_16281, n_16279);
  not g40274 (n_16283, n24374);
  and g40275 (n24375, n24370, n_16283);
  not g40276 (n_16284, n24373);
  not g40277 (n_16285, n24375);
  and g40278 (n24376, n_16284, n_16285);
  not g40279 (n_16286, n24376);
  and g40280 (n24377, n24230, n_16286);
  not g40281 (n_16287, n24230);
  and g40282 (n24378, n_16287, n_16285);
  and g40283 (n24379, n_16284, n24378);
  not g40284 (n_16288, n24379);
  and g40285 (n24380, n_11018, n_16288);
  and g40286 (n24381, n_15706, n_15705);
  and g40287 (n24382, \asqrt[1] , n24381);
  not g40288 (n_16289, n24382);
  and g40289 (n24383, n_15704, n_16289);
  not g40293 (n_16290, n24383);
  not g40294 (n_16291, n24386);
  and g40295 (n24387, n_16290, n_16291);
  not g40296 (n_16292, n24380);
  not g40297 (n_16293, n24387);
  and g40298 (n24388, n_16292, n_16293);
  not g40299 (n_16294, n24377);
  and g40300 (n24389, n_16294, n24388);
  not g40301 (n_16295, n24389);
  and g40302 (n24390, n_10602, n_16295);
  and g40303 (n24391, n_16294, n_16292);
  not g40304 (n_16296, n24391);
  and g40305 (n24392, n24387, n_16296);
  not g40306 (n_16297, n24390);
  not g40307 (n_16298, n24392);
  and g40308 (n24393, n_16297, n_16298);
  not g40309 (n_16299, n24393);
  and g40310 (n24394, n24223, n_16299);
  not g40311 (n_16300, n24223);
  and g40312 (n24395, n_16300, n_16298);
  and g40313 (n24396, n_16297, n24395);
  not g40314 (n_16301, n24396);
  and g40315 (n24397, n_10194, n_16301);
  and g40316 (n24398, n_15722, n_15721);
  and g40317 (n24399, \asqrt[1] , n24398);
  not g40318 (n_16302, n24399);
  and g40319 (n24400, n_15720, n_16302);
  not g40323 (n_16303, n24400);
  not g40324 (n_16304, n24403);
  and g40325 (n24404, n_16303, n_16304);
  not g40326 (n_16305, n24397);
  not g40327 (n_16306, n24404);
  and g40328 (n24405, n_16305, n_16306);
  not g40329 (n_16307, n24394);
  and g40330 (n24406, n_16307, n24405);
  not g40331 (n_16308, n24406);
  and g40332 (n24407, n_9794, n_16308);
  and g40333 (n24408, n_16307, n_16305);
  not g40334 (n_16309, n24408);
  and g40335 (n24409, n24404, n_16309);
  not g40336 (n_16310, n24407);
  not g40337 (n_16311, n24409);
  and g40338 (n24410, n_16310, n_16311);
  not g40339 (n_16312, n24410);
  and g40340 (n24411, n24216, n_16312);
  not g40341 (n_16313, n24216);
  and g40342 (n24412, n_16313, n_16311);
  and g40343 (n24413, n_16310, n24412);
  not g40344 (n_16314, n24413);
  and g40345 (n24414, n_9402, n_16314);
  and g40346 (n24415, n_15738, n_15737);
  and g40347 (n24416, \asqrt[1] , n24415);
  not g40348 (n_16315, n24416);
  and g40349 (n24417, n_15736, n_16315);
  not g40353 (n_16316, n24417);
  not g40354 (n_16317, n24420);
  and g40355 (n24421, n_16316, n_16317);
  not g40356 (n_16318, n24414);
  not g40357 (n_16319, n24421);
  and g40358 (n24422, n_16318, n_16319);
  not g40359 (n_16320, n24411);
  and g40360 (n24423, n_16320, n24422);
  not g40361 (n_16321, n24423);
  and g40362 (n24424, n_9018, n_16321);
  and g40363 (n24425, n_16320, n_16318);
  not g40364 (n_16322, n24425);
  and g40365 (n24426, n24421, n_16322);
  not g40366 (n_16323, n24424);
  not g40367 (n_16324, n24426);
  and g40368 (n24427, n_16323, n_16324);
  not g40369 (n_16325, n24427);
  and g40370 (n24428, n24209, n_16325);
  not g40371 (n_16326, n24209);
  and g40372 (n24429, n_16326, n_16324);
  and g40373 (n24430, n_16323, n24429);
  not g40374 (n_16327, n24430);
  and g40375 (n24431, n_8642, n_16327);
  and g40376 (n24432, n_15754, n_15753);
  and g40377 (n24433, \asqrt[1] , n24432);
  not g40378 (n_16328, n24433);
  and g40379 (n24434, n_15752, n_16328);
  not g40383 (n_16329, n24434);
  not g40384 (n_16330, n24437);
  and g40385 (n24438, n_16329, n_16330);
  not g40386 (n_16331, n24431);
  not g40387 (n_16332, n24438);
  and g40388 (n24439, n_16331, n_16332);
  not g40389 (n_16333, n24428);
  and g40390 (n24440, n_16333, n24439);
  not g40391 (n_16334, n24440);
  and g40392 (n24441, n_8274, n_16334);
  and g40393 (n24442, n_16333, n_16331);
  not g40394 (n_16335, n24442);
  and g40395 (n24443, n24438, n_16335);
  not g40396 (n_16336, n24441);
  not g40397 (n_16337, n24443);
  and g40398 (n24444, n_16336, n_16337);
  not g40399 (n_16338, n24444);
  and g40400 (n24445, n24202, n_16338);
  not g40401 (n_16339, n24202);
  and g40402 (n24446, n_16339, n_16337);
  and g40403 (n24447, n_16336, n24446);
  not g40404 (n_16340, n24447);
  and g40405 (n24448, n_7914, n_16340);
  and g40406 (n24449, n_15770, n_15769);
  and g40407 (n24450, \asqrt[1] , n24449);
  not g40408 (n_16341, n24450);
  and g40409 (n24451, n_15768, n_16341);
  not g40413 (n_16342, n24451);
  not g40414 (n_16343, n24454);
  and g40415 (n24455, n_16342, n_16343);
  not g40416 (n_16344, n24448);
  not g40417 (n_16345, n24455);
  and g40418 (n24456, n_16344, n_16345);
  not g40419 (n_16346, n24445);
  and g40420 (n24457, n_16346, n24456);
  not g40421 (n_16347, n24457);
  and g40422 (n24458, n_7562, n_16347);
  and g40423 (n24459, n_16346, n_16344);
  not g40424 (n_16348, n24459);
  and g40425 (n24460, n24455, n_16348);
  not g40426 (n_16349, n24458);
  not g40427 (n_16350, n24460);
  and g40428 (n24461, n_16349, n_16350);
  not g40429 (n_16351, n24461);
  and g40430 (n24462, n24195, n_16351);
  not g40431 (n_16352, n24195);
  and g40432 (n24463, n_16352, n_16350);
  and g40433 (n24464, n_16349, n24463);
  not g40434 (n_16353, n24464);
  and g40435 (n24465, n_7218, n_16353);
  and g40436 (n24466, n_15786, n_15785);
  and g40437 (n24467, \asqrt[1] , n24466);
  not g40438 (n_16354, n24467);
  and g40439 (n24468, n_15784, n_16354);
  not g40443 (n_16355, n24468);
  not g40444 (n_16356, n24471);
  and g40445 (n24472, n_16355, n_16356);
  not g40446 (n_16357, n24465);
  not g40447 (n_16358, n24472);
  and g40448 (n24473, n_16357, n_16358);
  not g40449 (n_16359, n24462);
  and g40450 (n24474, n_16359, n24473);
  not g40451 (n_16360, n24474);
  and g40452 (n24475, n_6882, n_16360);
  and g40453 (n24476, n_16359, n_16357);
  not g40454 (n_16361, n24476);
  and g40455 (n24477, n24472, n_16361);
  not g40456 (n_16362, n24475);
  not g40457 (n_16363, n24477);
  and g40458 (n24478, n_16362, n_16363);
  not g40459 (n_16364, n24478);
  and g40460 (n24479, n24188, n_16364);
  not g40461 (n_16365, n24188);
  and g40462 (n24480, n_16365, n_16363);
  and g40463 (n24481, n_16362, n24480);
  not g40464 (n_16366, n24481);
  and g40465 (n24482, n_6554, n_16366);
  and g40466 (n24483, n_15802, n_15801);
  and g40467 (n24484, \asqrt[1] , n24483);
  not g40468 (n_16367, n24484);
  and g40469 (n24485, n_15800, n_16367);
  not g40473 (n_16368, n24485);
  not g40474 (n_16369, n24488);
  and g40475 (n24489, n_16368, n_16369);
  not g40476 (n_16370, n24482);
  not g40477 (n_16371, n24489);
  and g40478 (n24490, n_16370, n_16371);
  not g40479 (n_16372, n24479);
  and g40480 (n24491, n_16372, n24490);
  not g40481 (n_16373, n24491);
  and g40482 (n24492, n_6234, n_16373);
  and g40483 (n24493, n_16372, n_16370);
  not g40484 (n_16374, n24493);
  and g40485 (n24494, n24489, n_16374);
  not g40486 (n_16375, n24492);
  not g40487 (n_16376, n24494);
  and g40488 (n24495, n_16375, n_16376);
  not g40489 (n_16377, n24495);
  and g40490 (n24496, n24181, n_16377);
  not g40491 (n_16378, n24181);
  and g40492 (n24497, n_16378, n_16376);
  and g40493 (n24498, n_16375, n24497);
  not g40494 (n_16379, n24498);
  and g40495 (n24499, n_5922, n_16379);
  and g40496 (n24500, n_15818, n_15817);
  and g40497 (n24501, \asqrt[1] , n24500);
  not g40498 (n_16380, n24501);
  and g40499 (n24502, n_15816, n_16380);
  not g40503 (n_16381, n24502);
  not g40504 (n_16382, n24505);
  and g40505 (n24506, n_16381, n_16382);
  not g40506 (n_16383, n24499);
  not g40507 (n_16384, n24506);
  and g40508 (n24507, n_16383, n_16384);
  not g40509 (n_16385, n24496);
  and g40510 (n24508, n_16385, n24507);
  not g40511 (n_16386, n24508);
  and g40512 (n24509, n_5618, n_16386);
  and g40513 (n24510, n_16385, n_16383);
  not g40514 (n_16387, n24510);
  and g40515 (n24511, n24506, n_16387);
  not g40516 (n_16388, n24509);
  not g40517 (n_16389, n24511);
  and g40518 (n24512, n_16388, n_16389);
  not g40519 (n_16390, n24512);
  and g40520 (n24513, n24174, n_16390);
  not g40521 (n_16391, n24174);
  and g40522 (n24514, n_16391, n_16389);
  and g40523 (n24515, n_16388, n24514);
  not g40524 (n_16392, n24515);
  and g40525 (n24516, n_5322, n_16392);
  and g40526 (n24517, n_15834, n_15833);
  and g40527 (n24518, \asqrt[1] , n24517);
  not g40528 (n_16393, n24518);
  and g40529 (n24519, n_15832, n_16393);
  not g40533 (n_16394, n24519);
  not g40534 (n_16395, n24522);
  and g40535 (n24523, n_16394, n_16395);
  not g40536 (n_16396, n24516);
  not g40537 (n_16397, n24523);
  and g40538 (n24524, n_16396, n_16397);
  not g40539 (n_16398, n24513);
  and g40540 (n24525, n_16398, n24524);
  not g40541 (n_16399, n24525);
  and g40542 (n24526, n_5034, n_16399);
  and g40543 (n24527, n_16398, n_16396);
  not g40544 (n_16400, n24527);
  and g40545 (n24528, n24523, n_16400);
  not g40546 (n_16401, n24526);
  not g40547 (n_16402, n24528);
  and g40548 (n24529, n_16401, n_16402);
  not g40549 (n_16403, n24529);
  and g40550 (n24530, n24167, n_16403);
  not g40551 (n_16404, n24167);
  and g40552 (n24531, n_16404, n_16402);
  and g40553 (n24532, n_16401, n24531);
  not g40554 (n_16405, n24532);
  and g40555 (n24533, n_4754, n_16405);
  and g40556 (n24534, n_15850, n_15849);
  and g40557 (n24535, \asqrt[1] , n24534);
  not g40558 (n_16406, n24535);
  and g40559 (n24536, n_15848, n_16406);
  not g40563 (n_16407, n24536);
  not g40564 (n_16408, n24539);
  and g40565 (n24540, n_16407, n_16408);
  not g40566 (n_16409, n24533);
  not g40567 (n_16410, n24540);
  and g40568 (n24541, n_16409, n_16410);
  not g40569 (n_16411, n24530);
  and g40570 (n24542, n_16411, n24541);
  not g40571 (n_16412, n24542);
  and g40572 (n24543, n_4482, n_16412);
  and g40573 (n24544, n_16411, n_16409);
  not g40574 (n_16413, n24544);
  and g40575 (n24545, n24540, n_16413);
  not g40576 (n_16414, n24543);
  not g40577 (n_16415, n24545);
  and g40578 (n24546, n_16414, n_16415);
  not g40579 (n_16416, n24546);
  and g40580 (n24547, n24160, n_16416);
  not g40581 (n_16417, n24160);
  and g40582 (n24548, n_16417, n_16415);
  and g40583 (n24549, n_16414, n24548);
  not g40584 (n_16418, n24549);
  and g40585 (n24550, n_4218, n_16418);
  and g40586 (n24551, n_15866, n_15865);
  and g40587 (n24552, \asqrt[1] , n24551);
  not g40588 (n_16419, n24552);
  and g40589 (n24553, n_15864, n_16419);
  not g40593 (n_16420, n24553);
  not g40594 (n_16421, n24556);
  and g40595 (n24557, n_16420, n_16421);
  not g40596 (n_16422, n24550);
  not g40597 (n_16423, n24557);
  and g40598 (n24558, n_16422, n_16423);
  not g40599 (n_16424, n24547);
  and g40600 (n24559, n_16424, n24558);
  not g40601 (n_16425, n24559);
  and g40602 (n24560, n_3962, n_16425);
  and g40603 (n24561, n_16424, n_16422);
  not g40604 (n_16426, n24561);
  and g40605 (n24562, n24557, n_16426);
  not g40606 (n_16427, n24560);
  not g40607 (n_16428, n24562);
  and g40608 (n24563, n_16427, n_16428);
  not g40609 (n_16429, n24563);
  and g40610 (n24564, n24153, n_16429);
  not g40611 (n_16430, n24153);
  and g40612 (n24565, n_16430, n_16428);
  and g40613 (n24566, n_16427, n24565);
  not g40614 (n_16431, n24566);
  and g40615 (n24567, n_3714, n_16431);
  and g40616 (n24568, n_15882, n_15881);
  and g40617 (n24569, \asqrt[1] , n24568);
  not g40618 (n_16432, n24569);
  and g40619 (n24570, n_15880, n_16432);
  not g40623 (n_16433, n24570);
  not g40624 (n_16434, n24573);
  and g40625 (n24574, n_16433, n_16434);
  not g40626 (n_16435, n24567);
  not g40627 (n_16436, n24574);
  and g40628 (n24575, n_16435, n_16436);
  not g40629 (n_16437, n24564);
  and g40630 (n24576, n_16437, n24575);
  not g40631 (n_16438, n24576);
  and g40632 (n24577, n_3474, n_16438);
  and g40633 (n24578, n_16437, n_16435);
  not g40634 (n_16439, n24578);
  and g40635 (n24579, n24574, n_16439);
  not g40636 (n_16440, n24577);
  not g40637 (n_16441, n24579);
  and g40638 (n24580, n_16440, n_16441);
  not g40639 (n_16442, n24580);
  and g40640 (n24581, n24146, n_16442);
  not g40641 (n_16443, n24146);
  and g40642 (n24582, n_16443, n_16441);
  and g40643 (n24583, n_16440, n24582);
  not g40644 (n_16444, n24583);
  and g40645 (n24584, n_3242, n_16444);
  and g40646 (n24585, n_15898, n_15897);
  and g40647 (n24586, \asqrt[1] , n24585);
  not g40648 (n_16445, n24586);
  and g40649 (n24587, n_15896, n_16445);
  not g40653 (n_16446, n24587);
  not g40654 (n_16447, n24590);
  and g40655 (n24591, n_16446, n_16447);
  not g40656 (n_16448, n24584);
  not g40657 (n_16449, n24591);
  and g40658 (n24592, n_16448, n_16449);
  not g40659 (n_16450, n24581);
  and g40660 (n24593, n_16450, n24592);
  not g40661 (n_16451, n24593);
  and g40662 (n24594, n_3018, n_16451);
  and g40663 (n24595, n_16450, n_16448);
  not g40664 (n_16452, n24595);
  and g40665 (n24596, n24591, n_16452);
  not g40666 (n_16453, n24594);
  not g40667 (n_16454, n24596);
  and g40668 (n24597, n_16453, n_16454);
  not g40669 (n_16455, n24597);
  and g40670 (n24598, n24139, n_16455);
  not g40671 (n_16456, n24139);
  and g40672 (n24599, n_16456, n_16454);
  and g40673 (n24600, n_16453, n24599);
  not g40674 (n_16457, n24600);
  and g40675 (n24601, n_2802, n_16457);
  and g40676 (n24602, n_15914, n_15913);
  and g40677 (n24603, \asqrt[1] , n24602);
  not g40678 (n_16458, n24603);
  and g40679 (n24604, n_15912, n_16458);
  not g40683 (n_16459, n24604);
  not g40684 (n_16460, n24607);
  and g40685 (n24608, n_16459, n_16460);
  not g40686 (n_16461, n24601);
  not g40687 (n_16462, n24608);
  and g40688 (n24609, n_16461, n_16462);
  not g40689 (n_16463, n24598);
  and g40690 (n24610, n_16463, n24609);
  not g40691 (n_16464, n24610);
  and g40692 (n24611, n_2594, n_16464);
  and g40693 (n24612, n_16463, n_16461);
  not g40694 (n_16465, n24612);
  and g40695 (n24613, n24608, n_16465);
  not g40696 (n_16466, n24611);
  not g40697 (n_16467, n24613);
  and g40698 (n24614, n_16466, n_16467);
  not g40699 (n_16468, n24614);
  and g40700 (n24615, n24132, n_16468);
  not g40701 (n_16469, n24132);
  and g40702 (n24616, n_16469, n_16467);
  and g40703 (n24617, n_16466, n24616);
  not g40704 (n_16470, n24617);
  and g40705 (n24618, n_2394, n_16470);
  and g40706 (n24619, n_15930, n_15929);
  and g40707 (n24620, \asqrt[1] , n24619);
  not g40708 (n_16471, n24620);
  and g40709 (n24621, n_15928, n_16471);
  not g40713 (n_16472, n24621);
  not g40714 (n_16473, n24624);
  and g40715 (n24625, n_16472, n_16473);
  not g40716 (n_16474, n24618);
  not g40717 (n_16475, n24625);
  and g40718 (n24626, n_16474, n_16475);
  not g40719 (n_16476, n24615);
  and g40720 (n24627, n_16476, n24626);
  not g40721 (n_16477, n24627);
  and g40722 (n24628, n_2202, n_16477);
  and g40723 (n24629, n_16476, n_16474);
  not g40724 (n_16478, n24629);
  and g40725 (n24630, n24625, n_16478);
  not g40726 (n_16479, n24628);
  not g40727 (n_16480, n24630);
  and g40728 (n24631, n_16479, n_16480);
  not g40729 (n_16481, n24631);
  and g40730 (n24632, n24125, n_16481);
  not g40731 (n_16482, n24125);
  and g40732 (n24633, n_16482, n_16480);
  and g40733 (n24634, n_16479, n24633);
  not g40734 (n_16483, n24634);
  and g40735 (n24635, n_2018, n_16483);
  and g40736 (n24636, n_15946, n_15945);
  and g40737 (n24637, \asqrt[1] , n24636);
  not g40738 (n_16484, n24637);
  and g40739 (n24638, n_15944, n_16484);
  not g40743 (n_16485, n24638);
  not g40744 (n_16486, n24641);
  and g40745 (n24642, n_16485, n_16486);
  not g40746 (n_16487, n24635);
  not g40747 (n_16488, n24642);
  and g40748 (n24643, n_16487, n_16488);
  not g40749 (n_16489, n24632);
  and g40750 (n24644, n_16489, n24643);
  not g40751 (n_16490, n24644);
  and g40752 (n24645, n_1842, n_16490);
  and g40753 (n24646, n_16489, n_16487);
  not g40754 (n_16491, n24646);
  and g40755 (n24647, n24642, n_16491);
  not g40756 (n_16492, n24645);
  not g40757 (n_16493, n24647);
  and g40758 (n24648, n_16492, n_16493);
  not g40759 (n_16494, n24648);
  and g40760 (n24649, n24118, n_16494);
  not g40761 (n_16495, n24118);
  and g40762 (n24650, n_16495, n_16493);
  and g40763 (n24651, n_16492, n24650);
  not g40764 (n_16496, n24651);
  and g40765 (n24652, n_1674, n_16496);
  and g40766 (n24653, n_15962, n_15961);
  and g40767 (n24654, \asqrt[1] , n24653);
  not g40768 (n_16497, n24654);
  and g40769 (n24655, n_15960, n_16497);
  not g40773 (n_16498, n24655);
  not g40774 (n_16499, n24658);
  and g40775 (n24659, n_16498, n_16499);
  not g40776 (n_16500, n24652);
  not g40777 (n_16501, n24659);
  and g40778 (n24660, n_16500, n_16501);
  not g40779 (n_16502, n24649);
  and g40780 (n24661, n_16502, n24660);
  not g40781 (n_16503, n24661);
  and g40782 (n24662, n_1514, n_16503);
  and g40783 (n24663, n_16502, n_16500);
  not g40784 (n_16504, n24663);
  and g40785 (n24664, n24659, n_16504);
  not g40786 (n_16505, n24662);
  not g40787 (n_16506, n24664);
  and g40788 (n24665, n_16505, n_16506);
  not g40789 (n_16507, n24665);
  and g40790 (n24666, n24111, n_16507);
  not g40791 (n_16508, n24111);
  and g40792 (n24667, n_16508, n_16506);
  and g40793 (n24668, n_16505, n24667);
  not g40794 (n_16509, n24668);
  and g40795 (n24669, n_1362, n_16509);
  and g40796 (n24670, n_15978, n_15977);
  and g40797 (n24671, \asqrt[1] , n24670);
  not g40798 (n_16510, n24671);
  and g40799 (n24672, n_15976, n_16510);
  not g40803 (n_16511, n24672);
  not g40804 (n_16512, n24675);
  and g40805 (n24676, n_16511, n_16512);
  not g40806 (n_16513, n24669);
  not g40807 (n_16514, n24676);
  and g40808 (n24677, n_16513, n_16514);
  not g40809 (n_16515, n24666);
  and g40810 (n24678, n_16515, n24677);
  not g40811 (n_16516, n24678);
  and g40812 (n24679, n_1218, n_16516);
  and g40813 (n24680, n_16515, n_16513);
  not g40814 (n_16517, n24680);
  and g40815 (n24681, n24676, n_16517);
  not g40816 (n_16518, n24679);
  not g40817 (n_16519, n24681);
  and g40818 (n24682, n_16518, n_16519);
  not g40819 (n_16520, n24682);
  and g40820 (n24683, n24104, n_16520);
  not g40821 (n_16521, n24104);
  and g40822 (n24684, n_16521, n_16519);
  and g40823 (n24685, n_16518, n24684);
  not g40824 (n_16522, n24685);
  and g40825 (n24686, n_1082, n_16522);
  and g40826 (n24687, n_15994, n_15993);
  and g40827 (n24688, \asqrt[1] , n24687);
  not g40828 (n_16523, n24688);
  and g40829 (n24689, n_15992, n_16523);
  not g40833 (n_16524, n24689);
  not g40834 (n_16525, n24692);
  and g40835 (n24693, n_16524, n_16525);
  not g40836 (n_16526, n24686);
  not g40837 (n_16527, n24693);
  and g40838 (n24694, n_16526, n_16527);
  not g40839 (n_16528, n24683);
  and g40840 (n24695, n_16528, n24694);
  not g40841 (n_16529, n24695);
  and g40842 (n24696, n_954, n_16529);
  and g40843 (n24697, n_16528, n_16526);
  not g40844 (n_16530, n24697);
  and g40845 (n24698, n24693, n_16530);
  not g40846 (n_16531, n24696);
  not g40847 (n_16532, n24698);
  and g40848 (n24699, n_16531, n_16532);
  not g40849 (n_16533, n24699);
  and g40850 (n24700, n24097, n_16533);
  not g40851 (n_16534, n24097);
  and g40852 (n24701, n_16534, n_16532);
  and g40853 (n24702, n_16531, n24701);
  not g40854 (n_16535, n24702);
  and g40855 (n24703, n_834, n_16535);
  and g40856 (n24704, n_16010, n_16009);
  and g40857 (n24705, \asqrt[1] , n24704);
  not g40858 (n_16536, n24705);
  and g40859 (n24706, n_16008, n_16536);
  not g40863 (n_16537, n24706);
  not g40864 (n_16538, n24709);
  and g40865 (n24710, n_16537, n_16538);
  not g40866 (n_16539, n24703);
  not g40867 (n_16540, n24710);
  and g40868 (n24711, n_16539, n_16540);
  not g40869 (n_16541, n24700);
  and g40870 (n24712, n_16541, n24711);
  not g40871 (n_16542, n24712);
  and g40872 (n24713, n_722, n_16542);
  and g40873 (n24714, n_16541, n_16539);
  not g40874 (n_16543, n24714);
  and g40875 (n24715, n24710, n_16543);
  not g40876 (n_16544, n24713);
  not g40877 (n_16545, n24715);
  and g40878 (n24716, n_16544, n_16545);
  not g40879 (n_16546, n24716);
  and g40880 (n24717, n24090, n_16546);
  not g40881 (n_16547, n24090);
  and g40882 (n24718, n_16547, n_16545);
  and g40883 (n24719, n_16544, n24718);
  not g40884 (n_16548, n24719);
  and g40885 (n24720, n_618, n_16548);
  and g40886 (n24721, n_16026, n_16025);
  and g40887 (n24722, \asqrt[1] , n24721);
  not g40888 (n_16549, n24722);
  and g40889 (n24723, n_16024, n_16549);
  not g40893 (n_16550, n24723);
  not g40894 (n_16551, n24726);
  and g40895 (n24727, n_16550, n_16551);
  not g40896 (n_16552, n24720);
  not g40897 (n_16553, n24727);
  and g40898 (n24728, n_16552, n_16553);
  not g40899 (n_16554, n24717);
  and g40900 (n24729, n_16554, n24728);
  not g40901 (n_16555, n24729);
  and g40902 (n24730, n_522, n_16555);
  and g40903 (n24731, n_16554, n_16552);
  not g40904 (n_16556, n24731);
  and g40905 (n24732, n24727, n_16556);
  not g40906 (n_16557, n24730);
  not g40907 (n_16558, n24732);
  and g40908 (n24733, n_16557, n_16558);
  not g40909 (n_16559, n24733);
  and g40910 (n24734, n24083, n_16559);
  not g40911 (n_16560, n24083);
  and g40912 (n24735, n_16560, n_16558);
  and g40913 (n24736, n_16557, n24735);
  not g40914 (n_16561, n24736);
  and g40915 (n24737, n_434, n_16561);
  and g40916 (n24738, n_16042, n_16041);
  and g40917 (n24739, \asqrt[1] , n24738);
  not g40918 (n_16562, n24739);
  and g40919 (n24740, n_16040, n_16562);
  not g40923 (n_16563, n24740);
  not g40924 (n_16564, n24743);
  and g40925 (n24744, n_16563, n_16564);
  not g40926 (n_16565, n24737);
  not g40927 (n_16566, n24744);
  and g40928 (n24745, n_16565, n_16566);
  not g40929 (n_16567, n24734);
  and g40930 (n24746, n_16567, n24745);
  not g40931 (n_16568, n24746);
  and g40932 (n24747, n_354, n_16568);
  and g40933 (n24748, n_16567, n_16565);
  not g40934 (n_16569, n24748);
  and g40935 (n24749, n24744, n_16569);
  not g40936 (n_16570, n24747);
  not g40937 (n_16571, n24749);
  and g40938 (n24750, n_16570, n_16571);
  not g40939 (n_16572, n24750);
  and g40940 (n24751, n24076, n_16572);
  not g40941 (n_16573, n24076);
  and g40942 (n24752, n_16573, n_16571);
  and g40943 (n24753, n_16570, n24752);
  not g40944 (n_16574, n24753);
  and g40945 (n24754, n_282, n_16574);
  and g40946 (n24755, n_16058, n_16057);
  and g40947 (n24756, \asqrt[1] , n24755);
  not g40948 (n_16575, n24756);
  and g40949 (n24757, n_16056, n_16575);
  not g40953 (n_16576, n24757);
  not g40954 (n_16577, n24760);
  and g40955 (n24761, n_16576, n_16577);
  not g40956 (n_16578, n24754);
  not g40957 (n_16579, n24761);
  and g40958 (n24762, n_16578, n_16579);
  not g40959 (n_16580, n24751);
  and g40960 (n24763, n_16580, n24762);
  not g40961 (n_16581, n24763);
  and g40962 (n24764, n_218, n_16581);
  and g40963 (n24765, n_16580, n_16578);
  not g40964 (n_16582, n24765);
  and g40965 (n24766, n24761, n_16582);
  not g40966 (n_16583, n24764);
  not g40967 (n_16584, n24766);
  and g40968 (n24767, n_16583, n_16584);
  not g40969 (n_16585, n24767);
  and g40970 (n24768, n24069, n_16585);
  not g40971 (n_16586, n24069);
  and g40972 (n24769, n_16586, n_16584);
  and g40973 (n24770, n_16583, n24769);
  not g40974 (n_16587, n24770);
  and g40975 (n24771, n_162, n_16587);
  and g40976 (n24772, n_16074, n_16073);
  and g40977 (n24773, \asqrt[1] , n24772);
  not g40978 (n_16588, n24773);
  and g40979 (n24774, n_16072, n_16588);
  not g40983 (n_16589, n24774);
  not g40984 (n_16590, n24777);
  and g40985 (n24778, n_16589, n_16590);
  not g40986 (n_16591, n24771);
  not g40987 (n_16592, n24778);
  and g40988 (n24779, n_16591, n_16592);
  not g40989 (n_16593, n24768);
  and g40990 (n24780, n_16593, n24779);
  not g40991 (n_16594, n24780);
  and g40992 (n24781, n_115, n_16594);
  and g40993 (n24782, n_16593, n_16591);
  not g40994 (n_16595, n24782);
  and g40995 (n24783, n24778, n_16595);
  not g40996 (n_16596, n24781);
  not g40997 (n_16597, n24783);
  and g40998 (n24784, n_16596, n_16597);
  not g40999 (n_16598, n24784);
  and g41000 (n24785, n24062, n_16598);
  not g41001 (n_16599, n24062);
  and g41002 (n24786, n_16599, n_16597);
  and g41003 (n24787, n_16596, n24786);
  not g41004 (n_16600, n24787);
  and g41005 (n24788, n_76, n_16600);
  and g41006 (n24789, n_16087, n_16086);
  and g41007 (n24790, \asqrt[1] , n24789);
  not g41008 (n_16601, n24790);
  and g41009 (n24791, n_16085, n_16601);
  not g41013 (n_16602, n24791);
  not g41014 (n_16603, n24794);
  and g41015 (n24795, n_16602, n_16603);
  and g41016 (n24796, n_16094, n_16093);
  and g41017 (n24797, \asqrt[1] , n24796);
  not g41022 (n_16606, n24788);
  not g41024 (n_16607, n24785);
  not g41026 (n_16608, n24801);
  and g41027 (n24802, n_21, n_16608);
  and g41028 (n24803, n_16607, n_16606);
  not g41029 (n_16609, n24803);
  and g41030 (n24804, n24795, n_16609);
  and g41031 (n24805, n_16093, \asqrt[1] );
  not g41032 (n_16610, n24805);
  and g41033 (n24806, n24034, n_16610);
  not g41034 (n_16611, n24796);
  and g41035 (n24807, \asqrt[63] , n_16611);
  not g41036 (n_16612, n24806);
  and g41037 (n24808, n_16612, n24807);
  not g41038 (n_16613, n24804);
  not g41039 (n_16614, n24808);
  and g41040 (n24809, n_16613, n_16614);
  not g41041 (n_16615, n24809);
  or g41042 (\asqrt[0] , n24802, n_16615);
  nor g41043 (n_16617, n24795, n24797);
  and g41044 (n24801, n_16607, n_16606, n_16099, n_16617);
  and g41045 (n24794, \asqrt[1] , n_16087, n24030, n_16086);
  and g41046 (n24026, \asqrt[2] , n_15576, n23274, n_15575);
  and g41047 (n24037, \asqrt[2] , n_15582, n_15584, n23288);
  and g41048 (n24061, \asqrt[1] , n_16078, n23318, n_16079);
  and g41049 (n24046, n_16618, n_16094, n_16093, n_15596);
  not g41050 (n_16618, n24043);
  and g41051 (n23270, \asqrt[3] , n_15073, n22530, n_15072);
  and g41052 (n23284, \asqrt[3] , n_15079, n_15081, n22544);
  and g41053 (n23314, \asqrt[2] , n_15567, n_15568, n23262);
  and g41054 (n23302, n_16619, n_15591, n_15590, n_15101);
  not g41055 (n_16619, n23299);
  and g41056 (n24777, \asqrt[1] , n_16074, n24013, n_16073);
  and g41057 (n22526, \asqrt[4] , n_14578, n21798, n_14577);
  and g41058 (n22540, \asqrt[4] , n_14584, n_14586, n21812);
  and g41059 (n23258, \asqrt[3] , n_15064, n_15065, n22518);
  and g41060 (n23293, \asqrt[3] , n_15089, n22554, n_15088);
  and g41061 (n22570, n_16620, n_15096, n_15095, n_14614);
  not g41062 (n_16620, n22567);
  or g41063 (\asqrt[60] , n243, n247, n250, n242);
  and g41067 (n24009, \asqrt[2] , n_15560, n23250, n_15559);
  and g41068 (n21794, \asqrt[5] , n_14091, n21077, n_14090);
  and g41069 (n21808, \asqrt[5] , n_14097, n_14099, n21091);
  and g41070 (n22514, \asqrt[4] , n_14569, n_14570, n21786);
  and g41071 (n24068, \asqrt[1] , n_16065, n_16066, n24001);
  and g41072 (n22550, \asqrt[4] , n_14594, n21822, n_14593);
  and g41073 (n22561, \asqrt[4] , n_14601, n_14602, n21834);
  and g41074 (n241, n_16624, n_53, n_52, n_27);
  not g41075 (n_16624, n238);
  and g41076 (n250, n_46, n_27, n_23, n_28);
  and g41077 (n21850, n_16625, n_14609, n_14608, n_14135);
  not g41078 (n_16625, n21847);
  or g41079 (\asqrt[59] , n296, n300, n305, n294);
  and g41083 (n23246, \asqrt[3] , n_15057, n22506, n_15056);
  and g41084 (n21073, \asqrt[6] , n_13611, n20361, n_13610);
  and g41085 (n21087, \asqrt[6] , n_13617, n_13619, n20375);
  and g41086 (n21782, \asqrt[5] , n_14082, n_14083, n21065);
  and g41087 (n23997, \asqrt[2] , n_15551, n_15552, n23238);
  and g41088 (n21818, \asqrt[5] , n_14107, n21101, n_14106);
  and g41089 (n21830, \asqrt[5] , n_14114, n_14115, n21113);
  and g41090 (n21841, \asqrt[5] , n_14123, n21125, n_14122);
  and g41091 (n293, n_16629, n_92, n_91, n_59);
  not g41092 (n_16629, n290);
  and g41094 (n_16631, n_57, n_49);
  and g41095 (n305, n_50, n_58, n_16630, n_16631);
  and g41096 (n21141, n_16632, n_14130, n_14129, n_13665);
  not g41097 (n_16632, n21138);
  or g41098 (\asqrt[58] , n365, n369, n374, n363);
  or g41102 (\asqrt[6] , n20440, n20444, n20449, n20438);
  and g41106 (n24760, \asqrt[1] , n_16058, n23989, n_16057);
  and g41107 (n22502, \asqrt[4] , n_14562, n21774, n_14561);
  and g41108 (n20357, \asqrt[7] , n_13139, n19657, n_13138);
  and g41109 (n20371, \asqrt[7] , n_13145, n_13147, n19671);
  and g41110 (n21061, \asqrt[6] , n_13602, n_13603, n20349);
  and g41111 (n23234, \asqrt[3] , n_15048, n_15049, n22494);
  and g41112 (n21097, \asqrt[6] , n_13627, n20385, n_13626);
  and g41113 (n21109, \asqrt[6] , n_13634, n_13635, n20397);
  and g41114 (n21121, \asqrt[6] , n_13643, n20409, n_13642);
  and g41115 (n223, n_16639, n_16640, n_35, n_36);
  not g41116 (n_16639, n197);
  not g41117 (n_16640, n194);
  and g41118 (n21132, \asqrt[6] , n_13650, n_13651, n20421);
  and g41119 (n362, n_16641, n_139, n_138, n_98);
  not g41120 (n_16641, n359);
  and g41122 (n_16643, n_96, n_89);
  and g41123 (n374, n_88, n_97, n_16642, n_16643);
  and g41124 (n20437, n_16644, n_13658, n_13657, n_13201);
  not g41125 (n_16644, n20434);
  and g41127 (n_16646, n_13199, n_13191);
  and g41128 (n20449, n_13190, n_13200, n_16645, n_16646);
  or g41129 (\asqrt[57] , n445, n449, n454, n443);
  or g41133 (\asqrt[7] , n19748, n19752, n19757, n19746);
  and g41137 (n23985, \asqrt[2] , n_15544, n23226, n_15543);
  and g41138 (n21770, \asqrt[5] , n_14075, n21053, n_14074);
  and g41139 (n232, n_46, n_27, \asqrt[62] , n_28);
  and g41140 (n19653, \asqrt[8] , n_12675, n18965, n_12674);
  and g41141 (n19667, \asqrt[8] , n_12681, n_12683, n18979);
  and g41142 (n20345, \asqrt[7] , n_13130, n_13131, n19645);
  and g41143 (n22490, \asqrt[4] , n_14553, n_14554, n21762);
  and g41144 (n24075, \asqrt[1] , n_16049, n_16050, n23977);
  and g41145 (n20381, \asqrt[7] , n_13155, n19681, n_13154);
  and g41146 (n20393, \asqrt[7] , n_13162, n_13163, n19693);
  and g41147 (n20405, \asqrt[7] , n_13171, n19705, n_13170);
  and g41148 (n20417, \asqrt[7] , n_13178, n_13179, n19717);
  and g41149 (n20428, \asqrt[7] , n_13187, n19729, n_13186);
  and g41150 (n19736, \asqrt[8] , n_12730, n_12731, n19049);
  and g41152 (n_16654, n_12743, n_12735);
  and g41153 (n19757, n_12734, n_12744, n_16653, n_16654);
  and g41154 (n442, n_16655, n_194, n_193, n_145);
  not g41155 (n_16655, n439);
  and g41157 (n_16657, n_143, n_136);
  and g41158 (n454, n_135, n_144, n_16656, n_16657);
  and g41159 (n19745, n_16658, n_13194, n_13193, n_12745);
  not g41160 (n_16658, n19742);
  or g41161 (\asqrt[56] , n537, n541, n546, n535);
  or g41165 (\asqrt[8] , n19068, n19072, n19077, n19066);
  and g41169 (n23222, \asqrt[3] , n_15041, n22482, n_15040);
  and g41170 (n21049, \asqrt[6] , n_13595, n20337, n_13594);
  and g41171 (n353, \asqrt[59] , n_84, n_82, n280);
  and g41172 (n18961, \asqrt[9] , n_12219, n18285, n_12218);
  and g41173 (n18975, \asqrt[9] , n_12225, n_12227, n18299);
  and g41174 (n19641, \asqrt[8] , n_12666, n_12667, n18953);
  and g41175 (n21758, \asqrt[5] , n_14066, n_14067, n21041);
  and g41176 (n23973, \asqrt[2] , n_15535, n_15536, n23214);
  and g41177 (n19677, \asqrt[8] , n_12691, n18989, n_12690);
  and g41178 (n19689, \asqrt[8] , n_12698, n_12699, n19001);
  and g41179 (n19701, \asqrt[8] , n_12707, n19013, n_12706);
  and g41180 (n19713, \asqrt[8] , n_12714, n_12715, n19025);
  and g41181 (n19725, \asqrt[8] , n_12723, n19037, n_12722);
  and g41182 (n19045, \asqrt[9] , n_12274, n_12275, n18369);
  and g41183 (n19056, \asqrt[9] , n_12283, n18381, n_12282);
  and g41185 (n_16666, n_12295, n_12287);
  and g41186 (n19077, n_12286, n_12296, n_16665, n_16666);
  and g41187 (n534, n_16667, n_258, n_257, n_201);
  not g41188 (n_16667, n531);
  and g41190 (n_16669, n_199, n_191);
  and g41191 (n546, n_190, n_200, n_16668, n_16669);
  and g41192 (n19065, n_16670, n_12738, n_12737, n_12297);
  not g41193 (n_16670, n19062);
  or g41194 (\asqrt[55] , n641, n645, n650, n639);
  or g41198 (\asqrt[9] , n18400, n18404, n18409, n18398);
  and g41202 (n24743, \asqrt[1] , n_16042, n23965, n_16041);
  and g41203 (n22478, \asqrt[4] , n_14546, n21750, n_14545);
  and g41204 (n20333, \asqrt[7] , n_13123, n19633, n_13122);
  and g41205 (n_16630, n_77, n_59);
  and g41206 (n275, n_57, \asqrt[61] , n_58, n_16630);
  and g41207 (n_16678, n_66, n_46);
  and g41208 (n266, n_27, n_28, n_67, n_16678);
  and g41209 (n344, n_16679, \asqrt[59] , n_73, n_72);
  not g41210 (n_16679, n262);
  and g41211 (n433, \asqrt[58] , n_130, n_132, n348);
  and g41212 (n18281, \asqrt[10] , n_11771, n17617, n_11770);
  and g41213 (n18295, \asqrt[10] , n_11777, n_11779, n17631);
  and g41214 (n18949, \asqrt[9] , n_12210, n_12211, n18273);
  and g41215 (n21037, \asqrt[6] , n_13586, n_13587, n20325);
  and g41216 (n23210, \asqrt[3] , n_15032, n_15033, n22470);
  and g41217 (n18985, \asqrt[9] , n_12235, n18309, n_12234);
  and g41218 (n18997, \asqrt[9] , n_12242, n_12243, n18321);
  and g41219 (n19009, \asqrt[9] , n_12251, n18333, n_12250);
  and g41220 (n19021, \asqrt[9] , n_12258, n_12259, n18345);
  and g41221 (n19033, \asqrt[9] , n_12267, n18357, n_12266);
  and g41222 (n18365, \asqrt[10] , n_11826, n_11827, n17701);
  and g41223 (n18377, \asqrt[10] , n_11835, n17713, n_11834);
  and g41224 (n18388, \asqrt[10] , n_11842, n_11843, n17725);
  and g41226 (n_16681, n_11855, n_11847);
  and g41227 (n18409, n_11846, n_11856, n_16680, n_16681);
  and g41228 (n638, n_16682, n_330, n_329, n_265);
  not g41229 (n_16682, n635);
  and g41231 (n_16684, n_263, n_255);
  and g41232 (n650, n_254, n_264, n_16683, n_16684);
  and g41233 (n18397, n_16685, n_12290, n_12289, n_11857);
  not g41234 (n_16685, n18394);
  or g41235 (\asqrt[54] , n758, n762, n767, n756);
  or g41239 (\asqrt[10] , n17744, n17748, n17753, n17742);
  and g41243 (n23961, \asqrt[2] , n_15528, n23202, n_15527);
  and g41244 (n21746, \asqrt[5] , n_14059, n21029, n_14058);
  and g41245 (n19629, \asqrt[8] , n_12659, n18941, n_12658);
  and g41246 (n422, \asqrt[58] , n_123, n_121, n336);
  and g41247 (n525, \asqrt[57] , n_187, n426, n_186);
  and g41248 (n17613, \asqrt[11] , n_11331, n16961, n_11330);
  and g41249 (n17627, \asqrt[11] , n_11337, n_11339, n16975);
  and g41250 (n18269, \asqrt[10] , n_11762, n_11763, n17605);
  and g41251 (n20321, \asqrt[7] , n_13114, n_13115, n19621);
  and g41252 (n22466, \asqrt[4] , n_14537, n_14538, n21738);
  and g41253 (n24082, \asqrt[1] , n_16033, n_16034, n23953);
  and g41254 (n18305, \asqrt[10] , n_11787, n17641, n_11786);
  and g41255 (n18317, \asqrt[10] , n_11794, n_11795, n17653);
  and g41256 (n18329, \asqrt[10] , n_11803, n17665, n_11802);
  and g41257 (n18341, \asqrt[10] , n_11810, n_11811, n17677);
  and g41258 (n18353, \asqrt[10] , n_11819, n17689, n_11818);
  and g41259 (n17697, \asqrt[11] , n_11386, n_11387, n17045);
  and g41260 (n17709, \asqrt[11] , n_11395, n17057, n_11394);
  and g41261 (n17721, \asqrt[11] , n_11402, n_11403, n17069);
  and g41262 (n17732, \asqrt[11] , n_11411, n17081, n_11410);
  and g41264 (n_16693, n_11423, n_11415);
  and g41265 (n17753, n_11414, n_11424, n_16692, n_16693);
  and g41266 (n755, n_16694, n_410, n_409, n_337);
  not g41267 (n_16694, n752);
  and g41269 (n_16696, n_335, n_327);
  and g41270 (n767, n_326, n_336, n_16695, n_16696);
  and g41271 (n17741, n_16697, n_11850, n_11849, n_11425);
  not g41272 (n_16697, n17738);
  or g41273 (\asqrt[53] , n886, n890, n895, n884);
  or g41277 (\asqrt[11] , n17100, n17104, n17109, n17098);
  and g41281 (n23198, \asqrt[3] , n_15025, n22458, n_15024);
  and g41282 (n21025, \asqrt[6] , n_13579, n20313, n_13578);
  and g41283 (n18937, \asqrt[9] , n_12203, n18261, n_12202);
  and g41284 (n514, \asqrt[57] , n_178, n_179, n414);
  and g41285 (n629, \asqrt[56] , n_250, n_251, n518);
  and g41286 (n16957, \asqrt[12] , n_10899, n16317, n_10898);
  and g41287 (n16971, \asqrt[12] , n_10905, n_10907, n16331);
  and g41288 (n17601, \asqrt[11] , n_11322, n_11323, n16949);
  and g41289 (n19617, \asqrt[8] , n_12650, n_12651, n18929);
  and g41290 (n21734, \asqrt[5] , n_14050, n_14051, n21017);
  and g41291 (n23949, \asqrt[2] , n_15519, n_15520, n23190);
  and g41292 (n17637, \asqrt[11] , n_11347, n16985, n_11346);
  and g41293 (n17649, \asqrt[11] , n_11354, n_11355, n16997);
  and g41294 (n17661, \asqrt[11] , n_11363, n17009, n_11362);
  and g41295 (n17673, \asqrt[11] , n_11370, n_11371, n17021);
  and g41296 (n17685, \asqrt[11] , n_11379, n17033, n_11378);
  and g41297 (n_16704, n_105, n_77);
  and g41298 (n_16705, n_59, n_57);
  and g41299 (n318, n_58, n_106, n_16704, n_16705);
  and g41300 (n_16642, n_116, n_98);
  and g41301 (n331, n_96, \asqrt[60] , n_97, n_16642);
  and g41302 (n17041, \asqrt[12] , n_10954, n_10955, n16401);
  and g41303 (n17053, \asqrt[12] , n_10963, n16413, n_10962);
  and g41304 (n17065, \asqrt[12] , n_10970, n_10971, n16425);
  and g41305 (n17077, \asqrt[12] , n_10979, n16437, n_10978);
  and g41306 (n17088, \asqrt[12] , n_10986, n_10987, n16449);
  and g41308 (n_16708, n_10999, n_10991);
  and g41309 (n17109, n_10990, n_11000, n_16707, n_16708);
  and g41310 (n883, n_16709, n_498, n_497, n_417);
  not g41311 (n_16709, n880);
  and g41313 (n_16711, n_415, n_407);
  and g41314 (n895, n_406, n_416, n_16710, n_16711);
  and g41315 (n17097, n_16712, n_11418, n_11417, n_11001);
  not g41316 (n_16712, n17094);
  or g41317 (\asqrt[52] , n1026, n1030, n1035, n1024);
  or g41321 (\asqrt[12] , n16468, n16472, n16477, n16466);
  and g41325 (n24726, \asqrt[1] , n_16026, n23941, n_16025);
  and g41326 (n22454, \asqrt[4] , n_14530, n21726, n_14529);
  and g41327 (n20309, \asqrt[7] , n_13107, n19609, n_13106);
  and g41328 (n18257, \asqrt[10] , n_11755, n17593, n_11754);
  and g41329 (n618, \asqrt[56] , n_243, n506, n_242);
  and g41330 (n746, \asqrt[55] , n_323, n622, n_322);
  and g41331 (n16313, \asqrt[13] , n_10475, n15685, n_10474);
  and g41332 (n16327, \asqrt[13] , n_10481, n_10483, n15699);
  and g41333 (n16945, \asqrt[12] , n_10890, n_10891, n16305);
  and g41334 (n18925, \asqrt[9] , n_12194, n_12195, n18249);
  and g41335 (n21013, \asqrt[6] , n_13570, n_13571, n20301);
  and g41336 (n23186, \asqrt[3] , n_15016, n_15017, n22446);
  and g41337 (n16981, \asqrt[12] , n_10915, n16341, n_10914);
  and g41338 (n16993, \asqrt[12] , n_10922, n_10923, n16353);
  and g41339 (n17005, \asqrt[12] , n_10931, n16365, n_10930);
  and g41340 (n17017, \asqrt[12] , n_10938, n_10939, n16377);
  and g41341 (n17029, \asqrt[12] , n_10947, n16389, n_10946);
  and g41342 (n16397, \asqrt[13] , n_10530, n_10531, n15769);
  and g41343 (n16409, \asqrt[13] , n_10539, n15781, n_10538);
  and g41344 (n16421, \asqrt[13] , n_10546, n_10547, n15793);
  and g41345 (n16433, \asqrt[13] , n_10555, n15805, n_10554);
  and g41346 (n16445, \asqrt[13] , n_10562, n_10563, n15817);
  and g41347 (n16456, \asqrt[13] , n_10571, n15829, n_10570);
  and g41349 (n_16720, n_10583, n_10575);
  and g41350 (n16477, n_10574, n_10584, n_16719, n_16720);
  and g41351 (n502, \asqrt[57] , n_170, n_168, n405);
  and g41352 (n1023, n_16721, n_594, n_593, n_505);
  not g41353 (n_16721, n1020);
  and g41355 (n_16723, n_503, n_495);
  and g41356 (n1035, n_494, n_504, n_16722, n_16723);
  and g41357 (n16465, n_16724, n_10994, n_10993, n_10585);
  not g41358 (n_16724, n16462);
  or g41359 (\asqrt[51] , n1178, n1182, n1187, n1176);
  or g41363 (\asqrt[13] , n15848, n15852, n15857, n15846);
  and g41367 (n23937, \asqrt[2] , n_15512, n23178, n_15511);
  and g41368 (n21722, \asqrt[5] , n_14043, n21005, n_14042);
  and g41369 (n19605, \asqrt[8] , n_12643, n18917, n_12642);
  and g41370 (n17589, \asqrt[11] , n_11315, n16937, n_11314);
  and g41371 (n735, \asqrt[55] , n_314, n_315, n610);
  and g41372 (n874, \asqrt[54] , n_402, n_403, n739);
  and g41373 (n15681, \asqrt[14] , n_10059, n15065, n_10058);
  and g41374 (n15695, \asqrt[14] , n_10065, n_10067, n15079);
  and g41375 (n16301, \asqrt[13] , n_10466, n_10467, n15673);
  and g41376 (n18245, \asqrt[10] , n_11746, n_11747, n17581);
  and g41377 (n20297, \asqrt[7] , n_13098, n_13099, n19597);
  and g41378 (n22442, \asqrt[4] , n_14521, n_14522, n21714);
  and g41379 (n24089, \asqrt[1] , n_16017, n_16018, n23929);
  and g41380 (n16337, \asqrt[13] , n_10491, n15709, n_10490);
  and g41381 (n16349, \asqrt[13] , n_10498, n_10499, n15721);
  and g41382 (n16361, \asqrt[13] , n_10507, n15733, n_10506);
  and g41383 (n16373, \asqrt[13] , n_10514, n_10515, n15745);
  and g41384 (n16385, \asqrt[13] , n_10523, n15757, n_10522);
  and g41385 (n15765, \asqrt[14] , n_10114, n_10115, n15149);
  and g41386 (n15777, \asqrt[14] , n_10123, n15161, n_10122);
  and g41387 (n15789, \asqrt[14] , n_10130, n_10131, n15173);
  and g41388 (n15801, \asqrt[14] , n_10139, n15185, n_10138);
  and g41389 (n15813, \asqrt[14] , n_10146, n_10147, n15197);
  and g41390 (n15825, \asqrt[14] , n_10155, n15209, n_10154);
  and g41391 (n15836, \asqrt[14] , n_10162, n_10163, n15221);
  and g41393 (n_16732, n_10175, n_10167);
  and g41394 (n15857, n_10166, n_10176, n_16731, n_16732);
  and g41395 (n606, \asqrt[56] , n_234, n_235, n494);
  and g41396 (n1175, n_16733, n_698, n_697, n_601);
  not g41397 (n_16733, n1172);
  and g41399 (n_16735, n_599, n_591);
  and g41400 (n1187, n_590, n_600, n_16734, n_16735);
  and g41401 (n15845, n_16736, n_10578, n_10577, n_10177);
  not g41402 (n_16736, n15842);
  or g41403 (\asqrt[50] , n1342, n1346, n1351, n1340);
  or g41407 (\asqrt[14] , n15240, n15244, n15249, n15238);
  and g41411 (n23174, \asqrt[3] , n_15009, n22434, n_15008);
  and g41412 (n21001, \asqrt[6] , n_13563, n20289, n_13562);
  and g41413 (n18913, \asqrt[9] , n_12187, n18237, n_12186);
  and g41414 (n16933, \asqrt[12] , n_10883, n16293, n_10882);
  and g41415 (n_16743, n_152, n_116);
  and g41416 (n_16744, n_98, n_96);
  and g41417 (n387, n_97, n_153, n_16743, n_16744);
  and g41418 (n_16656, n_163, n_145);
  and g41419 (n400, n_143, \asqrt[59] , n_144, n_16656);
  and g41420 (n863, \asqrt[54] , n_395, n727, n_394);
  and g41421 (n1014, \asqrt[53] , n_491, n867, n_490);
  and g41422 (n15061, \asqrt[15] , n_9651, n14457, n_9650);
  and g41423 (n15075, \asqrt[15] , n_9657, n_9659, n14471);
  and g41424 (n15669, \asqrt[14] , n_10050, n_10051, n15053);
  and g41425 (n17577, \asqrt[11] , n_11306, n_11307, n16925);
  and g41426 (n19593, \asqrt[8] , n_12634, n_12635, n18905);
  and g41427 (n21710, \asqrt[5] , n_14034, n_14035, n20993);
  and g41428 (n23925, \asqrt[2] , n_15503, n_15504, n23166);
  and g41429 (n15705, \asqrt[14] , n_10075, n15089, n_10074);
  and g41430 (n15717, \asqrt[14] , n_10082, n_10083, n15101);
  and g41431 (n15729, \asqrt[14] , n_10091, n15113, n_10090);
  and g41432 (n15741, \asqrt[14] , n_10098, n_10099, n15125);
  and g41433 (n15753, \asqrt[14] , n_10107, n15137, n_10106);
  and g41434 (n15145, \asqrt[15] , n_9706, n_9707, n14541);
  and g41435 (n15157, \asqrt[15] , n_9715, n14553, n_9714);
  and g41436 (n15169, \asqrt[15] , n_9722, n_9723, n14565);
  and g41437 (n15181, \asqrt[15] , n_9731, n14577, n_9730);
  and g41438 (n15193, \asqrt[15] , n_9738, n_9739, n14589);
  and g41439 (n15205, \asqrt[15] , n_9747, n14601, n_9746);
  and g41440 (n15217, \asqrt[15] , n_9754, n_9755, n14613);
  and g41441 (n15228, \asqrt[15] , n_9763, n14625, n_9762);
  and g41443 (n_16747, n_9775, n_9767);
  and g41444 (n15249, n_9766, n_9776, n_16746, n_16747);
  and g41445 (n723, \asqrt[55] , n_307, n598, n_306);
  and g41446 (n1339, n_16748, n_810, n_809, n_705);
  not g41447 (n_16748, n1336);
  and g41449 (n_16750, n_703, n_695);
  and g41450 (n1351, n_694, n_704, n_16749, n_16750);
  and g41451 (n15237, n_16751, n_10170, n_10169, n_9777);
  not g41452 (n_16751, n15234);
  or g41453 (\asqrt[49] , n1518, n1522, n1527, n1516);
  or g41457 (\asqrt[15] , n14644, n14648, n14653, n14642);
  and g41461 (n24709, \asqrt[1] , n_16010, n23917, n_16009);
  and g41462 (n22430, \asqrt[4] , n_14514, n21702, n_14513);
  and g41463 (n20285, \asqrt[7] , n_13091, n19585, n_13090);
  and g41464 (n18233, \asqrt[10] , n_11739, n17569, n_11738);
  and g41465 (n16289, \asqrt[13] , n_10459, n15661, n_10458);
  and g41466 (n594, \asqrt[56] , n_226, n_224, n485);
  and g41467 (n1003, \asqrt[53] , n_482, n_483, n855);
  and g41468 (n1166, \asqrt[52] , n_586, n_587, n1007);
  and g41469 (n14453, \asqrt[16] , n_9251, n13861, n_9250);
  and g41470 (n14467, \asqrt[16] , n_9257, n_9259, n13875);
  and g41471 (n15049, \asqrt[15] , n_9642, n_9643, n14445);
  and g41472 (n16921, \asqrt[12] , n_10874, n_10875, n16281);
  and g41473 (n18901, \asqrt[9] , n_12178, n_12179, n18225);
  and g41474 (n20989, \asqrt[6] , n_13554, n_13555, n20277);
  and g41475 (n23162, \asqrt[3] , n_15000, n_15001, n22422);
  and g41476 (n15085, \asqrt[15] , n_9667, n14481, n_9666);
  and g41477 (n15097, \asqrt[15] , n_9674, n_9675, n14493);
  and g41478 (n15109, \asqrt[15] , n_9683, n14505, n_9682);
  and g41479 (n15121, \asqrt[15] , n_9690, n_9691, n14517);
  and g41480 (n15133, \asqrt[15] , n_9699, n14529, n_9698);
  and g41481 (n14537, \asqrt[16] , n_9306, n_9307, n13945);
  and g41482 (n14549, \asqrt[16] , n_9315, n13957, n_9314);
  and g41483 (n14561, \asqrt[16] , n_9322, n_9323, n13969);
  and g41484 (n14573, \asqrt[16] , n_9331, n13981, n_9330);
  and g41485 (n14585, \asqrt[16] , n_9338, n_9339, n13993);
  and g41486 (n14597, \asqrt[16] , n_9347, n14005, n_9346);
  and g41487 (n14609, \asqrt[16] , n_9354, n_9355, n14017);
  and g41488 (n14621, \asqrt[16] , n_9363, n14029, n_9362);
  and g41489 (n14632, \asqrt[16] , n_9370, n_9371, n14041);
  and g41491 (n_16759, n_9383, n_9375);
  and g41492 (n14653, n_9374, n_9384, n_16758, n_16759);
  and g41493 (n851, \asqrt[54] , n_386, n_387, n715);
  and g41494 (n1515, n_16760, n_930, n_929, n_817);
  not g41495 (n_16760, n1512);
  and g41497 (n_16762, n_815, n_807);
  and g41498 (n1527, n_806, n_816, n_16761, n_16762);
  and g41499 (n14641, n_16763, n_9770, n_9769, n_9385);
  not g41500 (n_16763, n14638);
  or g41501 (\asqrt[48] , n1706, n1710, n1715, n1704);
  or g41505 (\asqrt[16] , n14060, n14064, n14069, n14058);
  and g41509 (n23913, \asqrt[2] , n_15496, n23154, n_15495);
  and g41510 (n21698, \asqrt[5] , n_14027, n20981, n_14026);
  and g41511 (n19581, \asqrt[8] , n_12627, n18893, n_12626);
  and g41512 (n17565, \asqrt[11] , n_11299, n16913, n_11298);
  and g41513 (n15657, \asqrt[14] , n_10043, n15041, n_10042);
  and g41514 (n711, \asqrt[55] , n_298, n_299, n586);
  and g41515 (n1155, \asqrt[52] , n_579, n995, n_578);
  and g41516 (n1330, \asqrt[51] , n_691, n1159, n_690);
  and g41517 (n13857, \asqrt[17] , n_8859, n13277, n_8858);
  and g41518 (n13871, \asqrt[17] , n_8865, n_8867, n13291);
  and g41519 (n14441, \asqrt[16] , n_9242, n_9243, n13849);
  and g41520 (n16277, \asqrt[13] , n_10450, n_10451, n15649);
  and g41521 (n18221, \asqrt[10] , n_11730, n_11731, n17557);
  and g41522 (n20273, \asqrt[7] , n_13082, n_13083, n19573);
  and g41523 (n22418, \asqrt[4] , n_14505, n_14506, n21690);
  and g41524 (n24096, \asqrt[1] , n_16001, n_16002, n23905);
  and g41525 (n14477, \asqrt[16] , n_9267, n13885, n_9266);
  and g41526 (n14489, \asqrt[16] , n_9274, n_9275, n13897);
  and g41527 (n14501, \asqrt[16] , n_9283, n13909, n_9282);
  and g41528 (n14513, \asqrt[16] , n_9290, n_9291, n13921);
  and g41529 (n14525, \asqrt[16] , n_9299, n13933, n_9298);
  and g41530 (n13941, \asqrt[17] , n_8914, n_8915, n13361);
  and g41531 (n13953, \asqrt[17] , n_8923, n13373, n_8922);
  and g41532 (n13965, \asqrt[17] , n_8930, n_8931, n13385);
  and g41533 (n13977, \asqrt[17] , n_8939, n13397, n_8938);
  and g41534 (n13989, \asqrt[17] , n_8946, n_8947, n13409);
  and g41535 (n14001, \asqrt[17] , n_8955, n13421, n_8954);
  and g41536 (n14013, \asqrt[17] , n_8962, n_8963, n13433);
  and g41537 (n14025, \asqrt[17] , n_8971, n13445, n_8970);
  and g41538 (n14037, \asqrt[17] , n_8978, n_8979, n13457);
  and g41539 (n14048, \asqrt[17] , n_8987, n13469, n_8986);
  and g41541 (n_16771, n_8999, n_8991);
  and g41542 (n14069, n_8990, n_9000, n_16770, n_16771);
  and g41543 (n_16772, n_208, n_163);
  and g41544 (n_16773, n_145, n_143);
  and g41545 (n467, n_144, n_209, n_16772, n_16773);
  and g41546 (n_16668, n_219, n_201);
  and g41547 (n480, n_199, \asqrt[58] , n_200, n_16668);
  and g41548 (n991, \asqrt[53] , n_475, n843, n_474);
  and g41549 (n1703, n_16775, n_1058, n_1057, n_937);
  not g41550 (n_16775, n1700);
  and g41552 (n_16777, n_935, n_927);
  and g41553 (n1715, n_926, n_936, n_16776, n_16777);
  and g41554 (n14057, n_16778, n_9378, n_9377, n_9001);
  not g41555 (n_16778, n14054);
  or g41556 (\asqrt[47] , n1906, n1910, n1915, n1904);
  or g41560 (\asqrt[17] , n13488, n13492, n13497, n13486);
  and g41564 (n23150, \asqrt[3] , n_14993, n22410, n_14992);
  and g41565 (n20977, \asqrt[6] , n_13547, n20265, n_13546);
  and g41566 (n18889, \asqrt[9] , n_12171, n18213, n_12170);
  and g41567 (n16909, \asqrt[12] , n_10867, n16269, n_10866);
  and g41568 (n15037, \asqrt[15] , n_9635, n14433, n_9634);
  and g41569 (n839, \asqrt[54] , n_379, n703, n_378);
  and g41570 (n1321, \asqrt[51] , n_681, n_683, n1149);
  and g41571 (n1506, \asqrt[50] , n_801, n_803, n1325);
  and g41572 (n13273, \asqrt[18] , n_8475, n12705, n_8474);
  and g41573 (n13287, \asqrt[18] , n_8481, n_8483, n12719);
  and g41574 (n13845, \asqrt[17] , n_8850, n_8851, n13265);
  and g41575 (n15645, \asqrt[14] , n_10034, n_10035, n15029);
  and g41576 (n17553, \asqrt[11] , n_11290, n_11291, n16901);
  and g41577 (n19569, \asqrt[8] , n_12618, n_12619, n18881);
  and g41578 (n21686, \asqrt[5] , n_14018, n_14019, n20969);
  and g41579 (n23901, \asqrt[2] , n_15487, n_15488, n23142);
  and g41580 (n13881, \asqrt[17] , n_8875, n13301, n_8874);
  and g41581 (n13893, \asqrt[17] , n_8882, n_8883, n13313);
  and g41582 (n13905, \asqrt[17] , n_8891, n13325, n_8890);
  and g41583 (n13917, \asqrt[17] , n_8898, n_8899, n13337);
  and g41584 (n13929, \asqrt[17] , n_8907, n13349, n_8906);
  and g41585 (n13357, \asqrt[18] , n_8530, n_8531, n12789);
  and g41586 (n13369, \asqrt[18] , n_8539, n12801, n_8538);
  and g41587 (n13381, \asqrt[18] , n_8546, n_8547, n12813);
  and g41588 (n13393, \asqrt[18] , n_8555, n12825, n_8554);
  and g41589 (n13405, \asqrt[18] , n_8562, n_8563, n12837);
  and g41590 (n13417, \asqrt[18] , n_8571, n12849, n_8570);
  and g41591 (n13429, \asqrt[18] , n_8578, n_8579, n12861);
  and g41592 (n13441, \asqrt[18] , n_8587, n12873, n_8586);
  and g41593 (n13453, \asqrt[18] , n_8594, n_8595, n12885);
  and g41594 (n13465, \asqrt[18] , n_8603, n12897, n_8602);
  and g41595 (n13476, \asqrt[18] , n_8610, n_8611, n12909);
  and g41597 (n_16786, n_8623, n_8615);
  and g41598 (n13497, n_8614, n_8624, n_16785, n_16786);
  and g41599 (n699, \asqrt[55] , n_290, n_288, n577);
  and g41600 (n1145, \asqrt[52] , n_569, n_571, n985);
  and g41601 (n1903, n_16787, n_1194, n_1193, n_1065);
  not g41602 (n_16787, n1900);
  and g41604 (n_16789, n_1063, n_1055);
  and g41605 (n1915, n_1054, n_1064, n_16788, n_16789);
  and g41606 (n13485, n_16790, n_8994, n_8993, n_8625);
  not g41607 (n_16790, n13482);
  or g41608 (\asqrt[46] , n2119, n2123, n2128, n2117);
  or g41612 (\asqrt[18] , n12928, n12932, n12937, n12926);
  and g41616 (n24692, \asqrt[1] , n_15994, n23893, n_15993);
  and g41617 (n22406, \asqrt[4] , n_14498, n21678, n_14497);
  and g41618 (n20261, \asqrt[7] , n_13075, n19561, n_13074);
  and g41619 (n18209, \asqrt[10] , n_11723, n17545, n_11722);
  and g41620 (n16265, \asqrt[13] , n_10443, n15637, n_10442);
  and g41621 (n14429, \asqrt[16] , n_9235, n13837, n_9234);
  and g41622 (n981, \asqrt[53] , n_465, n_467, n833);
  and g41623 (n1495, \asqrt[50] , n_795, n1311, n_794);
  and g41624 (n1694, \asqrt[49] , n_923, n1499, n_922);
  and g41625 (n12701, \asqrt[19] , n_8099, n12145, n_8098);
  and g41626 (n12715, \asqrt[19] , n_8105, n_8107, n12159);
  and g41627 (n13261, \asqrt[18] , n_8466, n_8467, n12693);
  and g41628 (n15025, \asqrt[15] , n_9626, n_9627, n14421);
  and g41629 (n16897, \asqrt[12] , n_10858, n_10859, n16257);
  and g41630 (n18877, \asqrt[9] , n_12162, n_12163, n18201);
  and g41631 (n20965, \asqrt[6] , n_13538, n_13539, n20253);
  and g41632 (n23138, \asqrt[3] , n_14984, n_14985, n22398);
  and g41633 (n13297, \asqrt[18] , n_8491, n12729, n_8490);
  and g41634 (n13309, \asqrt[18] , n_8498, n_8499, n12741);
  and g41635 (n13321, \asqrt[18] , n_8507, n12753, n_8506);
  and g41636 (n13333, \asqrt[18] , n_8514, n_8515, n12765);
  and g41637 (n13345, \asqrt[18] , n_8523, n12777, n_8522);
  and g41638 (n12785, \asqrt[19] , n_8154, n_8155, n12229);
  and g41639 (n12797, \asqrt[19] , n_8163, n12241, n_8162);
  and g41640 (n12809, \asqrt[19] , n_8170, n_8171, n12253);
  and g41641 (n12821, \asqrt[19] , n_8179, n12265, n_8178);
  and g41642 (n12833, \asqrt[19] , n_8186, n_8187, n12277);
  and g41643 (n12845, \asqrt[19] , n_8195, n12289, n_8194);
  and g41644 (n12857, \asqrt[19] , n_8202, n_8203, n12301);
  and g41645 (n12869, \asqrt[19] , n_8211, n12313, n_8210);
  and g41646 (n12881, \asqrt[19] , n_8218, n_8219, n12325);
  and g41647 (n12893, \asqrt[19] , n_8227, n12337, n_8226);
  and g41648 (n12905, \asqrt[19] , n_8234, n_8235, n12349);
  and g41649 (n12916, \asqrt[19] , n_8243, n12361, n_8242);
  and g41651 (n_16798, n_8255, n_8247);
  and g41652 (n12937, n_8246, n_8256, n_16797, n_16798);
  and g41653 (n829, \asqrt[54] , n_369, n_371, n693);
  and g41654 (n1307, \asqrt[51] , n_675, n1135, n_674);
  and g41655 (n2116, n_16799, n_1338, n_1337, n_1201);
  not g41656 (n_16799, n2113);
  and g41658 (n_16801, n_1199, n_1191);
  and g41659 (n2128, n_1190, n_1200, n_16800, n_16801);
  and g41660 (n12925, n_16802, n_8618, n_8617, n_8257);
  not g41661 (n_16802, n12922);
  or g41662 (\asqrt[45] , n2343, n2347, n2352, n2341);
  or g41666 (\asqrt[19] , n12380, n12384, n12389, n12378);
  and g41670 (n23889, \asqrt[2] , n_15480, n23130, n_15479);
  and g41671 (n21674, \asqrt[5] , n_14011, n20957, n_14010);
  and g41672 (n19557, \asqrt[8] , n_12611, n18869, n_12610);
  and g41673 (n17541, \asqrt[11] , n_11283, n16889, n_11282);
  and g41674 (n15633, \asqrt[14] , n_10027, n15017, n_10026);
  and g41675 (n13833, \asqrt[17] , n_8843, n13253, n_8842);
  and g41676 (n_16809, n_272, n_219);
  and g41677 (n_16810, n_201, n_199);
  and g41678 (n563, n_200, n_273, n_16809, n_16810);
  and g41679 (n_16683, n_283, n_265);
  and g41680 (n572, n_263, \asqrt[57] , n_264, n_16683);
  and g41681 (n689, n_16812, \asqrt[55] , n_279, n_278);
  not g41682 (n_16812, n558);
  and g41683 (n1131, \asqrt[52] , n_563, n971, n_562);
  and g41684 (n1683, \asqrt[49] , n_914, n_915, n1487);
  and g41685 (n1894, \asqrt[48] , n_1050, n_1051, n1687);
  and g41686 (n12141, \asqrt[20] , n_7731, n11597, n_7730);
  and g41687 (n12155, \asqrt[20] , n_7737, n_7739, n11611);
  and g41688 (n12689, \asqrt[19] , n_8090, n_8091, n12133);
  and g41689 (n14417, \asqrt[16] , n_9226, n_9227, n13825);
  and g41690 (n16253, \asqrt[13] , n_10434, n_10435, n15625);
  and g41691 (n18197, \asqrt[10] , n_11714, n_11715, n17533);
  and g41692 (n20249, \asqrt[7] , n_13066, n_13067, n19549);
  and g41693 (n22394, \asqrt[4] , n_14489, n_14490, n21666);
  and g41694 (n24103, \asqrt[1] , n_15985, n_15986, n23881);
  and g41695 (n12725, \asqrt[19] , n_8115, n12169, n_8114);
  and g41696 (n12737, \asqrt[19] , n_8122, n_8123, n12181);
  and g41697 (n12749, \asqrt[19] , n_8131, n12193, n_8130);
  and g41698 (n12761, \asqrt[19] , n_8138, n_8139, n12205);
  and g41699 (n12773, \asqrt[19] , n_8147, n12217, n_8146);
  and g41700 (n12225, \asqrt[20] , n_7786, n_7787, n11681);
  and g41701 (n12237, \asqrt[20] , n_7795, n11693, n_7794);
  and g41702 (n12249, \asqrt[20] , n_7802, n_7803, n11705);
  and g41703 (n12261, \asqrt[20] , n_7811, n11717, n_7810);
  and g41704 (n12273, \asqrt[20] , n_7818, n_7819, n11729);
  and g41705 (n12285, \asqrt[20] , n_7827, n11741, n_7826);
  and g41706 (n12297, \asqrt[20] , n_7834, n_7835, n11753);
  and g41707 (n12309, \asqrt[20] , n_7843, n11765, n_7842);
  and g41708 (n12321, \asqrt[20] , n_7850, n_7851, n11777);
  and g41709 (n12333, \asqrt[20] , n_7859, n11789, n_7858);
  and g41710 (n12345, \asqrt[20] , n_7866, n_7867, n11801);
  and g41711 (n12357, \asqrt[20] , n_7875, n11813, n_7874);
  and g41712 (n12368, \asqrt[20] , n_7882, n_7883, n11825);
  and g41714 (n_16814, n_7895, n_7887);
  and g41715 (n12389, n_7886, n_7896, n_16813, n_16814);
  and g41716 (n967, \asqrt[53] , n_459, n819, n_458);
  and g41717 (n1483, \asqrt[50] , n_786, n_787, n1299);
  and g41718 (n2340, n_16815, n_1490, n_1489, n_1345);
  not g41719 (n_16815, n2337);
  and g41721 (n_16817, n_1343, n_1335);
  and g41722 (n2352, n_1334, n_1344, n_16816, n_16817);
  and g41723 (n12377, n_16818, n_8250, n_8249, n_7897);
  not g41724 (n_16818, n12374);
  or g41725 (\asqrt[44] , n2579, n2583, n2588, n2577);
  or g41729 (\asqrt[20] , n11844, n11848, n11853, n11842);
  and g41733 (n23126, \asqrt[3] , n_14977, n22386, n_14976);
  and g41734 (n20953, \asqrt[6] , n_13531, n20241, n_13530);
  and g41735 (n18865, \asqrt[9] , n_12155, n18189, n_12154);
  and g41736 (n16885, \asqrt[12] , n_10851, n16245, n_10850);
  and g41737 (n15013, \asqrt[15] , n_9619, n14409, n_9618);
  and g41738 (n13249, \asqrt[18] , n_8459, n12681, n_8458);
  and g41739 (n815, \asqrt[54] , n_362, n_360, n681);
  and g41740 (n1295, \asqrt[51] , n_666, n_667, n1123);
  and g41741 (n1883, \asqrt[48] , n_1043, n1675, n_1042);
  and g41742 (n2107, \asqrt[47] , n_1187, n1887, n_1186);
  and g41743 (n11593, \asqrt[21] , n_7371, n11061, n_7370);
  and g41744 (n11607, \asqrt[21] , n_7377, n_7379, n11075);
  and g41745 (n12129, \asqrt[20] , n_7722, n_7723, n11585);
  and g41746 (n13821, \asqrt[17] , n_8834, n_8835, n13241);
  and g41747 (n15621, \asqrt[14] , n_10018, n_10019, n15005);
  and g41748 (n17529, \asqrt[11] , n_11274, n_11275, n16877);
  and g41749 (n19545, \asqrt[8] , n_12602, n_12603, n18857);
  and g41750 (n21662, \asqrt[5] , n_14002, n_14003, n20945);
  and g41751 (n23877, \asqrt[2] , n_15471, n_15472, n23118);
  and g41752 (n12165, \asqrt[20] , n_7747, n11621, n_7746);
  and g41753 (n12177, \asqrt[20] , n_7754, n_7755, n11633);
  and g41754 (n12189, \asqrt[20] , n_7763, n11645, n_7762);
  and g41755 (n12201, \asqrt[20] , n_7770, n_7771, n11657);
  and g41756 (n12213, \asqrt[20] , n_7779, n11669, n_7778);
  and g41757 (n11677, \asqrt[21] , n_7426, n_7427, n11145);
  and g41758 (n11689, \asqrt[21] , n_7435, n11157, n_7434);
  and g41759 (n11701, \asqrt[21] , n_7442, n_7443, n11169);
  and g41760 (n11713, \asqrt[21] , n_7451, n11181, n_7450);
  and g41761 (n11725, \asqrt[21] , n_7458, n_7459, n11193);
  and g41762 (n11737, \asqrt[21] , n_7467, n11205, n_7466);
  and g41763 (n11749, \asqrt[21] , n_7474, n_7475, n11217);
  and g41764 (n11761, \asqrt[21] , n_7483, n11229, n_7482);
  and g41765 (n11773, \asqrt[21] , n_7490, n_7491, n11241);
  and g41766 (n11785, \asqrt[21] , n_7499, n11253, n_7498);
  and g41767 (n11797, \asqrt[21] , n_7506, n_7507, n11265);
  and g41768 (n11809, \asqrt[21] , n_7515, n11277, n_7514);
  and g41769 (n11821, \asqrt[21] , n_7522, n_7523, n11289);
  and g41770 (n11832, \asqrt[21] , n_7531, n11301, n_7530);
  and g41772 (n_16826, n_7543, n_7535);
  and g41773 (n11853, n_7534, n_7544, n_16825, n_16826);
  and g41774 (n1119, \asqrt[52] , n_554, n_555, n959);
  and g41775 (n1671, \asqrt[49] , n_907, n1475, n_906);
  and g41776 (n2576, n_16827, n_1650, n_1649, n_1497);
  not g41777 (n_16827, n2573);
  and g41779 (n_16829, n_1495, n_1487);
  and g41780 (n2588, n_1486, n_1496, n_16828, n_16829);
  and g41781 (n11841, n_16830, n_7890, n_7889, n_7545);
  not g41782 (n_16830, n11838);
  or g41783 (\asqrt[43] , n2827, n2831, n2836, n2825);
  or g41787 (\asqrt[21] , n11320, n11324, n11329, n11318);
  and g41791 (n24675, \asqrt[1] , n_15978, n23869, n_15977);
  and g41792 (n22382, \asqrt[4] , n_14482, n21654, n_14481);
  and g41793 (n20237, \asqrt[7] , n_13059, n19537, n_13058);
  and g41794 (n18185, \asqrt[10] , n_11707, n17521, n_11706);
  and g41795 (n16241, \asqrt[13] , n_10427, n15613, n_10426);
  and g41796 (n14405, \asqrt[16] , n_9219, n13813, n_9218);
  and g41797 (n12677, \asqrt[19] , n_8083, n12121, n_8082);
  and g41798 (n955, \asqrt[53] , n_450, n_451, n807);
  and g41799 (n1471, \asqrt[50] , n_779, n1287, n_778);
  and g41800 (n2096, \asqrt[47] , n_1178, n_1179, n1875);
  and g41801 (n2331, \asqrt[46] , n_1330, n_1331, n2100);
  and g41802 (n11057, \asqrt[22] , n_7019, n10537, n_7018);
  and g41803 (n11071, \asqrt[22] , n_7025, n_7027, n10551);
  and g41804 (n11581, \asqrt[21] , n_7362, n_7363, n11049);
  and g41805 (n13237, \asqrt[18] , n_8450, n_8451, n12669);
  and g41806 (n15001, \asqrt[15] , n_9610, n_9611, n14397);
  and g41807 (n16873, \asqrt[12] , n_10842, n_10843, n16233);
  and g41808 (n18853, \asqrt[9] , n_12146, n_12147, n18177);
  and g41809 (n20941, \asqrt[6] , n_13522, n_13523, n20229);
  and g41810 (n23114, \asqrt[3] , n_14968, n_14969, n22374);
  and g41811 (n11617, \asqrt[21] , n_7387, n11085, n_7386);
  and g41812 (n11629, \asqrt[21] , n_7394, n_7395, n11097);
  and g41813 (n11641, \asqrt[21] , n_7403, n11109, n_7402);
  and g41814 (n11653, \asqrt[21] , n_7410, n_7411, n11121);
  and g41815 (n11665, \asqrt[21] , n_7419, n11133, n_7418);
  and g41816 (n11141, \asqrt[22] , n_7074, n_7075, n10621);
  and g41817 (n11153, \asqrt[22] , n_7083, n10633, n_7082);
  and g41818 (n11165, \asqrt[22] , n_7090, n_7091, n10645);
  and g41819 (n11177, \asqrt[22] , n_7099, n10657, n_7098);
  and g41820 (n11189, \asqrt[22] , n_7106, n_7107, n10669);
  and g41821 (n11201, \asqrt[22] , n_7115, n10681, n_7114);
  and g41822 (n11213, \asqrt[22] , n_7122, n_7123, n10693);
  and g41823 (n11225, \asqrt[22] , n_7131, n10705, n_7130);
  and g41824 (n11237, \asqrt[22] , n_7138, n_7139, n10717);
  and g41825 (n11249, \asqrt[22] , n_7147, n10729, n_7146);
  and g41826 (n11261, \asqrt[22] , n_7154, n_7155, n10741);
  and g41827 (n11273, \asqrt[22] , n_7163, n10753, n_7162);
  and g41828 (n11285, \asqrt[22] , n_7170, n_7171, n10765);
  and g41829 (n11297, \asqrt[22] , n_7179, n10777, n_7178);
  and g41830 (n11308, \asqrt[22] , n_7186, n_7187, n10789);
  and g41832 (n_16838, n_7199, n_7191);
  and g41833 (n11329, n_7190, n_7200, n_16837, n_16838);
  and g41834 (n_16839, n_344, n_283);
  and g41835 (n_16840, n_265, n_263);
  and g41836 (n663, n_264, n_345, n_16839, n_16840);
  and g41837 (n_16695, n_355, n_337);
  and g41838 (n676, n_335, \asqrt[56] , n_336, n_16695);
  and g41839 (n1283, \asqrt[51] , n_659, n1111, n_658);
  and g41840 (n1871, \asqrt[48] , n_1034, n_1035, n1663);
  and g41841 (n2824, n_16842, n_1818, n_1817, n_1657);
  not g41842 (n_16842, n2821);
  and g41844 (n_16844, n_1655, n_1647);
  and g41845 (n2836, n_1646, n_1656, n_16843, n_16844);
  and g41846 (n11317, n_16845, n_7538, n_7537, n_7201);
  not g41847 (n_16845, n11314);
  or g41848 (\asqrt[42] , n3087, n3091, n3096, n3085);
  or g41852 (\asqrt[22] , n10808, n10812, n10817, n10806);
  and g41856 (n23865, \asqrt[2] , n_15464, n23106, n_15463);
  and g41857 (n21650, \asqrt[5] , n_13995, n20933, n_13994);
  and g41858 (n19533, \asqrt[8] , n_12595, n18845, n_12594);
  and g41859 (n17517, \asqrt[11] , n_11267, n16865, n_11266);
  and g41860 (n15609, \asqrt[14] , n_10011, n14993, n_10010);
  and g41861 (n13809, \asqrt[17] , n_8827, n13229, n_8826);
  and g41862 (n12117, \asqrt[20] , n_7715, n11573, n_7714);
  and g41863 (n1107, \asqrt[52] , n_547, n947, n_546);
  and g41864 (n1659, \asqrt[49] , n_898, n_899, n1463);
  and g41865 (n2320, \asqrt[46] , n_1323, n2088, n_1322);
  and g41866 (n2567, \asqrt[45] , n_1483, n2324, n_1482);
  and g41867 (n10533, \asqrt[23] , n_6675, n10025, n_6674);
  and g41868 (n10547, \asqrt[23] , n_6681, n_6683, n10039);
  and g41869 (n11045, \asqrt[22] , n_7010, n_7011, n10525);
  and g41870 (n12665, \asqrt[19] , n_8074, n_8075, n12109);
  and g41871 (n14393, \asqrt[16] , n_9210, n_9211, n13801);
  and g41872 (n16229, \asqrt[13] , n_10418, n_10419, n15601);
  and g41873 (n18173, \asqrt[10] , n_11698, n_11699, n17509);
  and g41874 (n20225, \asqrt[7] , n_13050, n_13051, n19525);
  and g41875 (n22370, \asqrt[4] , n_14473, n_14474, n21642);
  and g41876 (n24110, \asqrt[1] , n_15969, n_15970, n23857);
  and g41877 (n11081, \asqrt[22] , n_7035, n10561, n_7034);
  and g41878 (n11093, \asqrt[22] , n_7042, n_7043, n10573);
  and g41879 (n11105, \asqrt[22] , n_7051, n10585, n_7050);
  and g41880 (n11117, \asqrt[22] , n_7058, n_7059, n10597);
  and g41881 (n11129, \asqrt[22] , n_7067, n10609, n_7066);
  and g41882 (n10617, \asqrt[23] , n_6730, n_6731, n10109);
  and g41883 (n10629, \asqrt[23] , n_6739, n10121, n_6738);
  and g41884 (n10641, \asqrt[23] , n_6746, n_6747, n10133);
  and g41885 (n10653, \asqrt[23] , n_6755, n10145, n_6754);
  and g41886 (n10665, \asqrt[23] , n_6762, n_6763, n10157);
  and g41887 (n10677, \asqrt[23] , n_6771, n10169, n_6770);
  and g41888 (n10689, \asqrt[23] , n_6778, n_6779, n10181);
  and g41889 (n10701, \asqrt[23] , n_6787, n10193, n_6786);
  and g41890 (n10713, \asqrt[23] , n_6794, n_6795, n10205);
  and g41891 (n10725, \asqrt[23] , n_6803, n10217, n_6802);
  and g41892 (n10737, \asqrt[23] , n_6810, n_6811, n10229);
  and g41893 (n10749, \asqrt[23] , n_6819, n10241, n_6818);
  and g41894 (n10761, \asqrt[23] , n_6826, n_6827, n10253);
  and g41895 (n10773, \asqrt[23] , n_6835, n10265, n_6834);
  and g41896 (n10785, \asqrt[23] , n_6842, n_6843, n10277);
  and g41897 (n10796, \asqrt[23] , n_6851, n10289, n_6850);
  and g41899 (n_16853, n_6863, n_6855);
  and g41900 (n10817, n_6854, n_6864, n_16852, n_16853);
  and g41901 (n943, \asqrt[53] , n_442, n_440, n798);
  and g41902 (n1459, \asqrt[50] , n_770, n_771, n1275);
  and g41903 (n2084, \asqrt[47] , n_1171, n1863, n_1170);
  and g41904 (n3084, n_16854, n_1994, n_1993, n_1825);
  not g41905 (n_16854, n3081);
  and g41907 (n_16856, n_1823, n_1815);
  and g41908 (n3096, n_1814, n_1824, n_16855, n_16856);
  and g41909 (n10805, n_16857, n_7194, n_7193, n_6865);
  not g41910 (n_16857, n10802);
  or g41911 (\asqrt[41] , n3359, n3363, n3368, n3357);
  or g41915 (\asqrt[23] , n10308, n10312, n10317, n10306);
  and g41919 (n23102, \asqrt[3] , n_14961, n22362, n_14960);
  and g41920 (n20929, \asqrt[6] , n_13515, n20217, n_13514);
  and g41921 (n18841, \asqrt[9] , n_12139, n18165, n_12138);
  and g41922 (n16861, \asqrt[12] , n_10835, n16221, n_10834);
  and g41923 (n14989, \asqrt[15] , n_9603, n14385, n_9602);
  and g41924 (n13225, \asqrt[18] , n_8443, n12657, n_8442);
  and g41925 (n11569, \asqrt[21] , n_7355, n11037, n_7354);
  and g41926 (n1271, \asqrt[51] , n_650, n_651, n1099);
  and g41927 (n1859, \asqrt[48] , n_1027, n1651, n_1026);
  and g41928 (n2556, \asqrt[45] , n_1474, n_1475, n2312);
  and g41929 (n2815, \asqrt[44] , n_1642, n_1643, n2560);
  and g41930 (n10021, \asqrt[24] , n_6339, n9525, n_6338);
  and g41931 (n10035, \asqrt[24] , n_6345, n_6347, n9539);
  and g41932 (n10521, \asqrt[23] , n_6666, n_6667, n10013);
  and g41933 (n12105, \asqrt[20] , n_7706, n_7707, n11561);
  and g41934 (n13797, \asqrt[17] , n_8818, n_8819, n13217);
  and g41935 (n15597, \asqrt[14] , n_10002, n_10003, n14981);
  and g41936 (n17505, \asqrt[11] , n_11258, n_11259, n16853);
  and g41937 (n19521, \asqrt[8] , n_12586, n_12587, n18833);
  and g41938 (n21638, \asqrt[5] , n_13986, n_13987, n20921);
  and g41939 (n23853, \asqrt[2] , n_15455, n_15456, n23094);
  and g41940 (n10557, \asqrt[23] , n_6691, n10049, n_6690);
  and g41941 (n10569, \asqrt[23] , n_6698, n_6699, n10061);
  and g41942 (n10581, \asqrt[23] , n_6707, n10073, n_6706);
  and g41943 (n10593, \asqrt[23] , n_6714, n_6715, n10085);
  and g41944 (n10605, \asqrt[23] , n_6723, n10097, n_6722);
  and g41945 (n10105, \asqrt[24] , n_6394, n_6395, n9609);
  and g41946 (n10117, \asqrt[24] , n_6403, n9621, n_6402);
  and g41947 (n10129, \asqrt[24] , n_6410, n_6411, n9633);
  and g41948 (n10141, \asqrt[24] , n_6419, n9645, n_6418);
  and g41949 (n10153, \asqrt[24] , n_6426, n_6427, n9657);
  and g41950 (n10165, \asqrt[24] , n_6435, n9669, n_6434);
  and g41951 (n10177, \asqrt[24] , n_6442, n_6443, n9681);
  and g41952 (n10189, \asqrt[24] , n_6451, n9693, n_6450);
  and g41953 (n10201, \asqrt[24] , n_6458, n_6459, n9705);
  and g41954 (n10213, \asqrt[24] , n_6467, n9717, n_6466);
  and g41955 (n10225, \asqrt[24] , n_6474, n_6475, n9729);
  and g41956 (n10237, \asqrt[24] , n_6483, n9741, n_6482);
  and g41957 (n10249, \asqrt[24] , n_6490, n_6491, n9753);
  and g41958 (n10261, \asqrt[24] , n_6499, n9765, n_6498);
  and g41959 (n10273, \asqrt[24] , n_6506, n_6507, n9777);
  and g41960 (n10285, \asqrt[24] , n_6515, n9789, n_6514);
  and g41961 (n10296, \asqrt[24] , n_6522, n_6523, n9801);
  and g41963 (n_16865, n_6535, n_6527);
  and g41964 (n10317, n_6526, n_6536, n_16864, n_16865);
  and g41965 (n1095, \asqrt[52] , n_538, n_539, n935);
  and g41966 (n1647, \asqrt[49] , n_891, n1451, n_890);
  and g41967 (n2308, \asqrt[46] , n_1314, n_1315, n2076);
  and g41968 (n3356, n_16866, n_2178, n_2177, n_2001);
  not g41969 (n_16866, n3353);
  and g41971 (n_16868, n_1999, n_1991);
  and g41972 (n3368, n_1990, n_2000, n_16867, n_16868);
  and g41973 (n10305, n_16869, n_6858, n_6857, n_6537);
  not g41974 (n_16869, n10302);
  or g41975 (\asqrt[40] , n3643, n3647, n3652, n3641);
  or g41979 (\asqrt[24] , n9820, n9824, n9829, n9818);
  and g41983 (n24658, \asqrt[1] , n_15962, n23845, n_15961);
  and g41984 (n22358, \asqrt[4] , n_14466, n21630, n_14465);
  and g41985 (n20213, \asqrt[7] , n_13043, n19513, n_13042);
  and g41986 (n18161, \asqrt[10] , n_11691, n17497, n_11690);
  and g41987 (n16217, \asqrt[13] , n_10411, n15589, n_10410);
  and g41988 (n14381, \asqrt[16] , n_9203, n13789, n_9202);
  and g41989 (n12653, \asqrt[19] , n_8067, n12097, n_8066);
  and g41990 (n11033, \asqrt[22] , n_7003, n10513, n_7002);
  and g41991 (n_16876, n_424, n_355);
  and g41992 (n_16877, n_337, n_335);
  and g41993 (n780, n_336, n_425, n_16876, n_16877);
  and g41994 (n_16710, n_435, n_417);
  and g41995 (n793, n_415, \asqrt[55] , n_416, n_16710);
  and g41996 (n1447, \asqrt[50] , n_763, n1263, n_762);
  and g41997 (n2072, \asqrt[47] , n_1162, n_1163, n1851);
  and g41998 (n2804, \asqrt[44] , n_1635, n2548, n_1634);
  and g41999 (n3075, \asqrt[43] , n_1811, n2808, n_1810);
  and g42000 (n9521, \asqrt[25] , n_6011, n9037, n_6010);
  and g42001 (n9535, \asqrt[25] , n_6017, n_6019, n9051);
  and g42002 (n10009, \asqrt[24] , n_6330, n_6331, n9513);
  and g42003 (n11557, \asqrt[21] , n_7346, n_7347, n11025);
  and g42004 (n13213, \asqrt[18] , n_8434, n_8435, n12645);
  and g42005 (n14977, \asqrt[15] , n_9594, n_9595, n14373);
  and g42006 (n16849, \asqrt[12] , n_10826, n_10827, n16209);
  and g42007 (n18829, \asqrt[9] , n_12130, n_12131, n18153);
  and g42008 (n20917, \asqrt[6] , n_13506, n_13507, n20205);
  and g42009 (n23090, \asqrt[3] , n_14952, n_14953, n22350);
  and g42010 (n10045, \asqrt[24] , n_6355, n9549, n_6354);
  and g42011 (n10057, \asqrt[24] , n_6362, n_6363, n9561);
  and g42012 (n10069, \asqrt[24] , n_6371, n9573, n_6370);
  and g42013 (n10081, \asqrt[24] , n_6378, n_6379, n9585);
  and g42014 (n10093, \asqrt[24] , n_6387, n9597, n_6386);
  and g42015 (n9605, \asqrt[25] , n_6066, n_6067, n9121);
  and g42016 (n9617, \asqrt[25] , n_6075, n9133, n_6074);
  and g42017 (n9629, \asqrt[25] , n_6082, n_6083, n9145);
  and g42018 (n9641, \asqrt[25] , n_6091, n9157, n_6090);
  and g42019 (n9653, \asqrt[25] , n_6098, n_6099, n9169);
  and g42020 (n9665, \asqrt[25] , n_6107, n9181, n_6106);
  and g42021 (n9677, \asqrt[25] , n_6114, n_6115, n9193);
  and g42022 (n9689, \asqrt[25] , n_6123, n9205, n_6122);
  and g42023 (n9701, \asqrt[25] , n_6130, n_6131, n9217);
  and g42024 (n9713, \asqrt[25] , n_6139, n9229, n_6138);
  and g42025 (n9725, \asqrt[25] , n_6146, n_6147, n9241);
  and g42026 (n9737, \asqrt[25] , n_6155, n9253, n_6154);
  and g42027 (n9749, \asqrt[25] , n_6162, n_6163, n9265);
  and g42028 (n9761, \asqrt[25] , n_6171, n9277, n_6170);
  and g42029 (n9773, \asqrt[25] , n_6178, n_6179, n9289);
  and g42030 (n9785, \asqrt[25] , n_6187, n9301, n_6186);
  and g42031 (n9797, \asqrt[25] , n_6194, n_6195, n9313);
  and g42032 (n9808, \asqrt[25] , n_6203, n9325, n_6202);
  and g42034 (n_16880, n_6215, n_6207);
  and g42035 (n9829, n_6206, n_6216, n_16879, n_16880);
  and g42036 (n1259, \asqrt[51] , n_643, n1087, n_642);
  and g42037 (n1847, \asqrt[48] , n_1018, n_1019, n1639);
  and g42038 (n2544, \asqrt[45] , n_1467, n2300, n_1466);
  and g42039 (n3640, n_16881, n_2370, n_2369, n_2185);
  not g42040 (n_16881, n3637);
  and g42042 (n_16883, n_2183, n_2175);
  and g42043 (n3652, n_2174, n_2184, n_16882, n_16883);
  and g42044 (n9817, n_16884, n_6530, n_6529, n_6217);
  not g42045 (n_16884, n9814);
  or g42046 (\asqrt[39] , n3939, n3943, n3948, n3937);
  or g42050 (\asqrt[25] , n9344, n9348, n9353, n9342);
  and g42054 (n23841, \asqrt[2] , n_15448, n23082, n_15447);
  and g42055 (n21626, \asqrt[5] , n_13979, n20909, n_13978);
  and g42056 (n19509, \asqrt[8] , n_12579, n18821, n_12578);
  and g42057 (n17493, \asqrt[11] , n_11251, n16841, n_11250);
  and g42058 (n15585, \asqrt[14] , n_9995, n14969, n_9994);
  and g42059 (n13785, \asqrt[17] , n_8811, n13205, n_8810);
  and g42060 (n12093, \asqrt[20] , n_7699, n11549, n_7698);
  and g42061 (n10509, \asqrt[23] , n_6659, n10001, n_6658);
  and g42062 (n1083, \asqrt[52] , n_530, n_528, n926);
  and g42063 (n1635, \asqrt[49] , n_882, n_883, n1439);
  and g42064 (n2296, \asqrt[46] , n_1307, n2064, n_1306);
  and g42065 (n3064, \asqrt[43] , n_1802, n_1803, n2796);
  and g42066 (n3347, \asqrt[42] , n_1986, n_1987, n3068);
  and g42067 (n9033, \asqrt[26] , n_5691, n8561, n_5690);
  and g42068 (n9047, \asqrt[26] , n_5697, n_5699, n8575);
  and g42069 (n9509, \asqrt[25] , n_6002, n_6003, n9025);
  and g42070 (n11021, \asqrt[22] , n_6994, n_6995, n10501);
  and g42071 (n12641, \asqrt[19] , n_8058, n_8059, n12085);
  and g42072 (n14369, \asqrt[16] , n_9194, n_9195, n13777);
  and g42073 (n16205, \asqrt[13] , n_10402, n_10403, n15577);
  and g42074 (n18149, \asqrt[10] , n_11682, n_11683, n17485);
  and g42075 (n20201, \asqrt[7] , n_13034, n_13035, n19501);
  and g42076 (n22346, \asqrt[4] , n_14457, n_14458, n21618);
  and g42077 (n24117, \asqrt[1] , n_15953, n_15954, n23833);
  and g42078 (n9545, \asqrt[25] , n_6027, n9061, n_6026);
  and g42079 (n9557, \asqrt[25] , n_6034, n_6035, n9073);
  and g42080 (n9569, \asqrt[25] , n_6043, n9085, n_6042);
  and g42081 (n9581, \asqrt[25] , n_6050, n_6051, n9097);
  and g42082 (n9593, \asqrt[25] , n_6059, n9109, n_6058);
  and g42083 (n9117, \asqrt[26] , n_5746, n_5747, n8645);
  and g42084 (n9129, \asqrt[26] , n_5755, n8657, n_5754);
  and g42085 (n9141, \asqrt[26] , n_5762, n_5763, n8669);
  and g42086 (n9153, \asqrt[26] , n_5771, n8681, n_5770);
  and g42087 (n9165, \asqrt[26] , n_5778, n_5779, n8693);
  and g42088 (n9177, \asqrt[26] , n_5787, n8705, n_5786);
  and g42089 (n9189, \asqrt[26] , n_5794, n_5795, n8717);
  and g42090 (n9201, \asqrt[26] , n_5803, n8729, n_5802);
  and g42091 (n9213, \asqrt[26] , n_5810, n_5811, n8741);
  and g42092 (n9225, \asqrt[26] , n_5819, n8753, n_5818);
  and g42093 (n9237, \asqrt[26] , n_5826, n_5827, n8765);
  and g42094 (n9249, \asqrt[26] , n_5835, n8777, n_5834);
  and g42095 (n9261, \asqrt[26] , n_5842, n_5843, n8789);
  and g42096 (n9273, \asqrt[26] , n_5851, n8801, n_5850);
  and g42097 (n9285, \asqrt[26] , n_5858, n_5859, n8813);
  and g42098 (n9297, \asqrt[26] , n_5867, n8825, n_5866);
  and g42099 (n9309, \asqrt[26] , n_5874, n_5875, n8837);
  and g42100 (n9321, \asqrt[26] , n_5883, n8849, n_5882);
  and g42101 (n9332, \asqrt[26] , n_5890, n_5891, n8861);
  and g42103 (n_16892, n_5903, n_5895);
  and g42104 (n9353, n_5894, n_5904, n_16891, n_16892);
  and g42105 (n1435, \asqrt[50] , n_754, n_755, n1251);
  and g42106 (n2060, \asqrt[47] , n_1155, n1839, n_1154);
  and g42107 (n2792, \asqrt[44] , n_1626, n_1627, n2536);
  and g42108 (n3936, n_16893, n_2570, n_2569, n_2377);
  not g42109 (n_16893, n3933);
  and g42111 (n_16895, n_2375, n_2367);
  and g42112 (n3948, n_2366, n_2376, n_16894, n_16895);
  and g42113 (n9341, n_16896, n_6210, n_6209, n_5905);
  not g42114 (n_16896, n9338);
  or g42115 (\asqrt[38] , n4247, n4251, n4256, n4245);
  or g42119 (\asqrt[26] , n8880, n8884, n8889, n8878);
  and g42123 (n23078, \asqrt[3] , n_14945, n22338, n_14944);
  and g42124 (n20905, \asqrt[6] , n_13499, n20193, n_13498);
  and g42125 (n18817, \asqrt[9] , n_12123, n18141, n_12122);
  and g42126 (n16837, \asqrt[12] , n_10819, n16197, n_10818);
  and g42127 (n14965, \asqrt[15] , n_9587, n14361, n_9586);
  and g42128 (n13201, \asqrt[18] , n_8427, n12633, n_8426);
  and g42129 (n11545, \asqrt[21] , n_7339, n11013, n_7338);
  and g42130 (n9997, \asqrt[24] , n_6323, n9501, n_6322);
  and g42131 (n1247, \asqrt[51] , n_634, n_635, n1075);
  and g42132 (n1835, \asqrt[48] , n_1011, n1627, n_1010);
  and g42133 (n2532, \asqrt[45] , n_1458, n_1459, n2288);
  and g42134 (n3336, \asqrt[42] , n_1979, n3056, n_1978);
  and g42135 (n3631, \asqrt[41] , n_2171, n3340, n_2170);
  and g42136 (n8557, \asqrt[27] , n_5379, n8097, n_5378);
  and g42137 (n8571, \asqrt[27] , n_5385, n_5387, n8111);
  and g42138 (n9021, \asqrt[26] , n_5682, n_5683, n8549);
  and g42139 (n10497, \asqrt[23] , n_6650, n_6651, n9989);
  and g42140 (n12081, \asqrt[20] , n_7690, n_7691, n11537);
  and g42141 (n13773, \asqrt[17] , n_8802, n_8803, n13193);
  and g42142 (n15573, \asqrt[14] , n_9986, n_9987, n14957);
  and g42143 (n17481, \asqrt[11] , n_11242, n_11243, n16829);
  and g42144 (n19497, \asqrt[8] , n_12570, n_12571, n18809);
  and g42145 (n21614, \asqrt[5] , n_13970, n_13971, n20897);
  and g42146 (n23829, \asqrt[2] , n_15439, n_15440, n23070);
  and g42147 (n9057, \asqrt[26] , n_5707, n8585, n_5706);
  and g42148 (n9069, \asqrt[26] , n_5714, n_5715, n8597);
  and g42149 (n9081, \asqrt[26] , n_5723, n8609, n_5722);
  and g42150 (n9093, \asqrt[26] , n_5730, n_5731, n8621);
  and g42151 (n9105, \asqrt[26] , n_5739, n8633, n_5738);
  and g42152 (n8641, \asqrt[27] , n_5434, n_5435, n8181);
  and g42153 (n8653, \asqrt[27] , n_5443, n8193, n_5442);
  and g42154 (n8665, \asqrt[27] , n_5450, n_5451, n8205);
  and g42155 (n8677, \asqrt[27] , n_5459, n8217, n_5458);
  and g42156 (n8689, \asqrt[27] , n_5466, n_5467, n8229);
  and g42157 (n8701, \asqrt[27] , n_5475, n8241, n_5474);
  and g42158 (n8713, \asqrt[27] , n_5482, n_5483, n8253);
  and g42159 (n8725, \asqrt[27] , n_5491, n8265, n_5490);
  and g42160 (n8737, \asqrt[27] , n_5498, n_5499, n8277);
  and g42161 (n8749, \asqrt[27] , n_5507, n8289, n_5506);
  and g42162 (n8761, \asqrt[27] , n_5514, n_5515, n8301);
  and g42163 (n8773, \asqrt[27] , n_5523, n8313, n_5522);
  and g42164 (n8785, \asqrt[27] , n_5530, n_5531, n8325);
  and g42165 (n8797, \asqrt[27] , n_5539, n8337, n_5538);
  and g42166 (n8809, \asqrt[27] , n_5546, n_5547, n8349);
  and g42167 (n8821, \asqrt[27] , n_5555, n8361, n_5554);
  and g42168 (n8833, \asqrt[27] , n_5562, n_5563, n8373);
  and g42169 (n8845, \asqrt[27] , n_5571, n8385, n_5570);
  and g42170 (n8857, \asqrt[27] , n_5578, n_5579, n8397);
  and g42171 (n8868, \asqrt[27] , n_5587, n8409, n_5586);
  and g42173 (n_16904, n_5599, n_5591);
  and g42174 (n8889, n_5590, n_5600, n_16903, n_16904);
  and g42175 (n_16905, n_512, n_435);
  and g42176 (n_16906, n_417, n_415);
  and g42177 (n908, n_416, n_513, n_16905, n_16906);
  and g42178 (n_16722, n_523, n_505);
  and g42179 (n921, n_503, \asqrt[54] , n_504, n_16722);
  and g42180 (n1623, \asqrt[49] , n_875, n1427, n_874);
  and g42181 (n2284, \asqrt[46] , n_1298, n_1299, n2052);
  and g42182 (n3052, \asqrt[43] , n_1795, n2784, n_1794);
  and g42183 (n4244, n_16908, n_2778, n_2777, n_2577);
  not g42184 (n_16908, n4241);
  and g42186 (n_16910, n_2575, n_2567);
  and g42187 (n4256, n_2566, n_2576, n_16909, n_16910);
  and g42188 (n8877, n_16911, n_5898, n_5897, n_5601);
  not g42189 (n_16911, n8874);
  or g42190 (\asqrt[37] , n4567, n4571, n4576, n4565);
  or g42194 (\asqrt[27] , n8428, n8432, n8437, n8426);
  and g42198 (n24641, \asqrt[1] , n_15946, n23821, n_15945);
  and g42199 (n22334, \asqrt[4] , n_14450, n21606, n_14449);
  and g42200 (n20189, \asqrt[7] , n_13027, n19489, n_13026);
  and g42201 (n18137, \asqrt[10] , n_11675, n17473, n_11674);
  and g42202 (n16193, \asqrt[13] , n_10395, n15565, n_10394);
  and g42203 (n14357, \asqrt[16] , n_9187, n13765, n_9186);
  and g42204 (n12629, \asqrt[19] , n_8051, n12073, n_8050);
  and g42205 (n11009, \asqrt[22] , n_6987, n10489, n_6986);
  and g42206 (n9497, \asqrt[25] , n_5995, n9013, n_5994);
  and g42207 (n1423, \asqrt[50] , n_747, n1239, n_746);
  and g42208 (n2048, \asqrt[47] , n_1146, n_1147, n1827);
  and g42209 (n2780, \asqrt[44] , n_1619, n2524, n_1618);
  and g42210 (n3620, \asqrt[41] , n_2162, n_2163, n3328);
  and g42211 (n3927, \asqrt[40] , n_2362, n_2363, n3624);
  and g42212 (n8093, \asqrt[28] , n_5075, n7645, n_5074);
  and g42213 (n8107, \asqrt[28] , n_5081, n_5083, n7659);
  and g42214 (n8545, \asqrt[27] , n_5370, n_5371, n8085);
  and g42215 (n9985, \asqrt[24] , n_6314, n_6315, n9489);
  and g42216 (n11533, \asqrt[21] , n_7330, n_7331, n11001);
  and g42217 (n13189, \asqrt[18] , n_8418, n_8419, n12621);
  and g42218 (n14953, \asqrt[15] , n_9578, n_9579, n14349);
  and g42219 (n16825, \asqrt[12] , n_10810, n_10811, n16185);
  and g42220 (n18805, \asqrt[9] , n_12114, n_12115, n18129);
  and g42221 (n20893, \asqrt[6] , n_13490, n_13491, n20181);
  and g42222 (n23066, \asqrt[3] , n_14936, n_14937, n22326);
  and g42223 (n8581, \asqrt[27] , n_5395, n8121, n_5394);
  and g42224 (n8593, \asqrt[27] , n_5402, n_5403, n8133);
  and g42225 (n8605, \asqrt[27] , n_5411, n8145, n_5410);
  and g42226 (n8617, \asqrt[27] , n_5418, n_5419, n8157);
  and g42227 (n8629, \asqrt[27] , n_5427, n8169, n_5426);
  and g42228 (n8177, \asqrt[28] , n_5130, n_5131, n7729);
  and g42229 (n8189, \asqrt[28] , n_5139, n7741, n_5138);
  and g42230 (n8201, \asqrt[28] , n_5146, n_5147, n7753);
  and g42231 (n8213, \asqrt[28] , n_5155, n7765, n_5154);
  and g42232 (n8225, \asqrt[28] , n_5162, n_5163, n7777);
  and g42233 (n8237, \asqrt[28] , n_5171, n7789, n_5170);
  and g42234 (n8249, \asqrt[28] , n_5178, n_5179, n7801);
  and g42235 (n8261, \asqrt[28] , n_5187, n7813, n_5186);
  and g42236 (n8273, \asqrt[28] , n_5194, n_5195, n7825);
  and g42237 (n8285, \asqrt[28] , n_5203, n7837, n_5202);
  and g42238 (n8297, \asqrt[28] , n_5210, n_5211, n7849);
  and g42239 (n8309, \asqrt[28] , n_5219, n7861, n_5218);
  and g42240 (n8321, \asqrt[28] , n_5226, n_5227, n7873);
  and g42241 (n8333, \asqrt[28] , n_5235, n7885, n_5234);
  and g42242 (n8345, \asqrt[28] , n_5242, n_5243, n7897);
  and g42243 (n8357, \asqrt[28] , n_5251, n7909, n_5250);
  and g42244 (n8369, \asqrt[28] , n_5258, n_5259, n7921);
  and g42245 (n8381, \asqrt[28] , n_5267, n7933, n_5266);
  and g42246 (n8393, \asqrt[28] , n_5274, n_5275, n7945);
  and g42247 (n8405, \asqrt[28] , n_5283, n7957, n_5282);
  and g42248 (n8416, \asqrt[28] , n_5290, n_5291, n7969);
  and g42250 (n_16919, n_5303, n_5295);
  and g42251 (n8437, n_5294, n_5304, n_16918, n_16919);
  and g42252 (n1235, \asqrt[51] , n_626, n_624, n1066);
  and g42253 (n1823, \asqrt[48] , n_1002, n_1003, n1615);
  and g42254 (n2520, \asqrt[45] , n_1451, n2276, n_1450);
  and g42255 (n3324, \asqrt[42] , n_1970, n_1971, n3044);
  and g42256 (n4564, n_16920, n_2994, n_2993, n_2785);
  not g42257 (n_16920, n4561);
  and g42259 (n_16922, n_2783, n_2775);
  and g42260 (n4576, n_2774, n_2784, n_16921, n_16922);
  and g42261 (n8425, n_16923, n_5594, n_5593, n_5305);
  not g42262 (n_16923, n8422);
  or g42263 (\asqrt[36] , n4899, n4903, n4908, n4897);
  or g42267 (\asqrt[28] , n7988, n7992, n7997, n7986);
  and g42271 (n23817, \asqrt[2] , n_15432, n23058, n_15431);
  and g42272 (n21602, \asqrt[5] , n_13963, n20885, n_13962);
  and g42273 (n19485, \asqrt[8] , n_12563, n18797, n_12562);
  and g42274 (n17469, \asqrt[11] , n_11235, n16817, n_11234);
  and g42275 (n15561, \asqrt[14] , n_9979, n14945, n_9978);
  and g42276 (n13761, \asqrt[17] , n_8795, n13181, n_8794);
  and g42277 (n12069, \asqrt[20] , n_7683, n11525, n_7682);
  and g42278 (n10485, \asqrt[23] , n_6643, n9977, n_6642);
  and g42279 (n9009, \asqrt[26] , n_5675, n8537, n_5674);
  and g42280 (n1611, \asqrt[49] , n_866, n_867, n1415);
  and g42281 (n2272, \asqrt[46] , n_1291, n2040, n_1290);
  and g42282 (n3040, \asqrt[43] , n_1786, n_1787, n2772);
  and g42283 (n3916, \asqrt[40] , n_2355, n3612, n_2354);
  and g42284 (n4235, \asqrt[39] , n_2563, n3920, n_2562);
  and g42285 (n7641, \asqrt[29] , n_4779, n7205, n_4778);
  and g42286 (n7655, \asqrt[29] , n_4785, n_4787, n7219);
  and g42287 (n8081, \asqrt[28] , n_5066, n_5067, n7633);
  and g42288 (n9485, \asqrt[25] , n_5986, n_5987, n9001);
  and g42289 (n10997, \asqrt[22] , n_6978, n_6979, n10477);
  and g42290 (n12617, \asqrt[19] , n_8042, n_8043, n12061);
  and g42291 (n14345, \asqrt[16] , n_9178, n_9179, n13753);
  and g42292 (n16181, \asqrt[13] , n_10386, n_10387, n15553);
  and g42293 (n18125, \asqrt[10] , n_11666, n_11667, n17461);
  and g42294 (n20177, \asqrt[7] , n_13018, n_13019, n19477);
  and g42295 (n22322, \asqrt[4] , n_14441, n_14442, n21594);
  and g42296 (n24124, \asqrt[1] , n_15937, n_15938, n23809);
  and g42297 (n8117, \asqrt[28] , n_5091, n7669, n_5090);
  and g42298 (n8129, \asqrt[28] , n_5098, n_5099, n7681);
  and g42299 (n8141, \asqrt[28] , n_5107, n7693, n_5106);
  and g42300 (n8153, \asqrt[28] , n_5114, n_5115, n7705);
  and g42301 (n8165, \asqrt[28] , n_5123, n7717, n_5122);
  and g42302 (n7725, \asqrt[29] , n_4834, n_4835, n7289);
  and g42303 (n7737, \asqrt[29] , n_4843, n7301, n_4842);
  and g42304 (n7749, \asqrt[29] , n_4850, n_4851, n7313);
  and g42305 (n7761, \asqrt[29] , n_4859, n7325, n_4858);
  and g42306 (n7773, \asqrt[29] , n_4866, n_4867, n7337);
  and g42307 (n7785, \asqrt[29] , n_4875, n7349, n_4874);
  and g42308 (n7797, \asqrt[29] , n_4882, n_4883, n7361);
  and g42309 (n7809, \asqrt[29] , n_4891, n7373, n_4890);
  and g42310 (n7821, \asqrt[29] , n_4898, n_4899, n7385);
  and g42311 (n7833, \asqrt[29] , n_4907, n7397, n_4906);
  and g42312 (n7845, \asqrt[29] , n_4914, n_4915, n7409);
  and g42313 (n7857, \asqrt[29] , n_4923, n7421, n_4922);
  and g42314 (n7869, \asqrt[29] , n_4930, n_4931, n7433);
  and g42315 (n7881, \asqrt[29] , n_4939, n7445, n_4938);
  and g42316 (n7893, \asqrt[29] , n_4946, n_4947, n7457);
  and g42317 (n7905, \asqrt[29] , n_4955, n7469, n_4954);
  and g42318 (n7917, \asqrt[29] , n_4962, n_4963, n7481);
  and g42319 (n7929, \asqrt[29] , n_4971, n7493, n_4970);
  and g42320 (n7941, \asqrt[29] , n_4978, n_4979, n7505);
  and g42321 (n7953, \asqrt[29] , n_4987, n7517, n_4986);
  and g42322 (n7965, \asqrt[29] , n_4994, n_4995, n7529);
  and g42323 (n7976, \asqrt[29] , n_5003, n7541, n_5002);
  and g42325 (n_16931, n_5015, n_5007);
  and g42326 (n7997, n_5006, n_5016, n_16930, n_16931);
  and g42327 (n1411, \asqrt[50] , n_738, n_739, n1227);
  and g42328 (n2036, \asqrt[47] , n_1139, n1815, n_1138);
  and g42329 (n2768, \asqrt[44] , n_1610, n_1611, n2512);
  and g42330 (n3608, \asqrt[41] , n_2155, n3316, n_2154);
  and g42331 (n4896, n_16932, n_3218, n_3217, n_3001);
  not g42332 (n_16932, n4893);
  and g42334 (n_16934, n_2999, n_2991);
  and g42335 (n4908, n_2990, n_3000, n_16933, n_16934);
  and g42336 (n7985, n_16935, n_5298, n_5297, n_5017);
  not g42337 (n_16935, n7982);
  or g42338 (\asqrt[35] , n5243, n5247, n5252, n5241);
  or g42342 (\asqrt[29] , n7560, n7564, n7569, n7558);
  and g42346 (n23054, \asqrt[3] , n_14929, n22314, n_14928);
  and g42347 (n20881, \asqrt[6] , n_13483, n20169, n_13482);
  and g42348 (n18793, \asqrt[9] , n_12107, n18117, n_12106);
  and g42349 (n16813, \asqrt[12] , n_10803, n16173, n_10802);
  and g42350 (n14941, \asqrt[15] , n_9571, n14337, n_9570);
  and g42351 (n13177, \asqrt[18] , n_8411, n12609, n_8410);
  and g42352 (n11521, \asqrt[21] , n_7323, n10989, n_7322);
  and g42353 (n9973, \asqrt[24] , n_6307, n9477, n_6306);
  and g42354 (n8533, \asqrt[27] , n_5363, n8073, n_5362);
  and g42355 (n_16942, n_608, n_523);
  and g42356 (n_16943, n_505, n_503);
  and g42357 (n1048, n_504, n_609, n_16942, n_16943);
  and g42358 (n_16734, n_619, n_601);
  and g42359 (n1061, n_599, \asqrt[53] , n_600, n_16734);
  and g42360 (n1811, \asqrt[48] , n_995, n1603, n_994);
  and g42361 (n2508, \asqrt[45] , n_1442, n_1443, n2264);
  and g42362 (n3312, \asqrt[42] , n_1963, n3032, n_1962);
  and g42363 (n4224, \asqrt[39] , n_2554, n_2555, n3908);
  and g42364 (n4555, \asqrt[38] , n_2770, n_2771, n4228);
  and g42365 (n7201, \asqrt[30] , n_4490, n_4488, n6779);
  and g42366 (n7215, \asqrt[30] , n_4497, n_4499, n6791);
  and g42367 (n7629, \asqrt[29] , n_4770, n_4771, n7193);
  and g42368 (n8997, \asqrt[26] , n_5666, n_5667, n8525);
  and g42369 (n10473, \asqrt[23] , n_6634, n_6635, n9965);
  and g42370 (n12057, \asqrt[20] , n_7674, n_7675, n11513);
  and g42371 (n13749, \asqrt[17] , n_8786, n_8787, n13169);
  and g42372 (n15549, \asqrt[14] , n_9970, n_9971, n14933);
  and g42373 (n17457, \asqrt[11] , n_11226, n_11227, n16805);
  and g42374 (n19473, \asqrt[8] , n_12554, n_12555, n18785);
  and g42375 (n21590, \asqrt[5] , n_13954, n_13955, n20873);
  and g42376 (n23805, \asqrt[2] , n_15423, n_15424, n23046);
  and g42377 (n7665, \asqrt[29] , n_4795, n7229, n_4794);
  and g42378 (n7677, \asqrt[29] , n_4802, n_4803, n7241);
  and g42379 (n7689, \asqrt[29] , n_4811, n7253, n_4810);
  and g42380 (n7701, \asqrt[29] , n_4818, n_4819, n7265);
  and g42381 (n7713, \asqrt[29] , n_4827, n7277, n_4826);
  and g42382 (n7285, \asqrt[30] , n_4546, n_4547, n6861);
  and g42383 (n7297, \asqrt[30] , n_4555, n6873, n_4554);
  and g42384 (n7309, \asqrt[30] , n_4562, n_4563, n6885);
  and g42385 (n7321, \asqrt[30] , n_4571, n6897, n_4570);
  and g42386 (n7333, \asqrt[30] , n_4578, n_4579, n6909);
  and g42387 (n7345, \asqrt[30] , n_4587, n6921, n_4586);
  and g42388 (n7357, \asqrt[30] , n_4594, n_4595, n6933);
  and g42389 (n7369, \asqrt[30] , n_4603, n6945, n_4602);
  and g42390 (n7381, \asqrt[30] , n_4610, n_4611, n6957);
  and g42391 (n7393, \asqrt[30] , n_4619, n6969, n_4618);
  and g42392 (n7405, \asqrt[30] , n_4626, n_4627, n6981);
  and g42393 (n7417, \asqrt[30] , n_4635, n6993, n_4634);
  and g42394 (n7429, \asqrt[30] , n_4642, n_4643, n7005);
  and g42395 (n7441, \asqrt[30] , n_4651, n7017, n_4650);
  and g42396 (n7453, \asqrt[30] , n_4658, n_4659, n7029);
  and g42397 (n7465, \asqrt[30] , n_4667, n7041, n_4666);
  and g42398 (n7477, \asqrt[30] , n_4674, n_4675, n7053);
  and g42399 (n7489, \asqrt[30] , n_4683, n7065, n_4682);
  and g42400 (n7501, \asqrt[30] , n_4690, n_4691, n7077);
  and g42401 (n7513, \asqrt[30] , n_4699, n7089, n_4698);
  and g42402 (n7525, \asqrt[30] , n_4706, n_4707, n7101);
  and g42403 (n7537, \asqrt[30] , n_4715, n7113, n_4714);
  and g42404 (n7548, \asqrt[30] , n_4722, n_4723, n7125);
  and g42406 (n_16946, n_4735, n_4727);
  and g42407 (n7569, n_4726, n_4736, n_16945, n_16946);
  and g42408 (n1599, \asqrt[49] , n_859, n1403, n_858);
  and g42409 (n2260, \asqrt[46] , n_1282, n_1283, n2028);
  and g42410 (n3028, \asqrt[43] , n_1779, n2760, n_1778);
  and g42411 (n3904, \asqrt[40] , n_2346, n_2347, n3600);
  and g42412 (n5240, n_16947, n_3450, n_3449, n_3225);
  not g42413 (n_16947, n5237);
  and g42415 (n_16949, n_3223, n_3215);
  and g42416 (n5252, n_3214, n_3224, n_16948, n_16949);
  and g42417 (n7557, n_16950, n_5010, n_5009, n_4737);
  not g42418 (n_16950, n7554);
  or g42419 (\asqrt[34] , n5599, n5603, n5608, n5597);
  or g42423 (\asqrt[30] , n7144, n7148, n7153, n7142);
  and g42427 (n24624, \asqrt[1] , n_15930, n23797, n_15929);
  and g42428 (n22310, \asqrt[4] , n_14434, n21582, n_14433);
  and g42429 (n20165, \asqrt[7] , n_13011, n19465, n_13010);
  and g42430 (n18113, \asqrt[10] , n_11659, n17449, n_11658);
  and g42431 (n16169, \asqrt[13] , n_10379, n15541, n_10378);
  and g42432 (n14333, \asqrt[16] , n_9171, n13741, n_9170);
  and g42433 (n12605, \asqrt[19] , n_8035, n12049, n_8034);
  and g42434 (n10985, \asqrt[22] , n_6971, n10465, n_6970);
  and g42435 (n9473, \asqrt[25] , n_5979, n8989, n_5978);
  and g42436 (n8069, \asqrt[28] , n_5059, n7621, n_5058);
  and g42437 (n1399, \asqrt[50] , n_730, n_728, n1218);
  and g42438 (n2024, \asqrt[47] , n_1130, n_1131, n1803);
  and g42439 (n2756, \asqrt[44] , n_1603, n2500, n_1602);
  and g42440 (n3596, \asqrt[41] , n_2146, n_2147, n3304);
  and g42441 (n4544, \asqrt[38] , n_2763, n4216, n_2762);
  and g42442 (n4887, \asqrt[37] , n_2987, n4548, n_2986);
  and g42443 (n6787, n_16957, \asqrt[31] , n_4215, n_4214);
  not g42444 (n_16957, n6368);
  and g42445 (n8521, \asqrt[27] , n_5354, n_5355, n8061);
  and g42446 (n9961, \asqrt[24] , n_6298, n_6299, n9465);
  and g42447 (n11509, \asqrt[21] , n_7314, n_7315, n10977);
  and g42448 (n13165, \asqrt[18] , n_8402, n_8403, n12597);
  and g42449 (n14929, \asqrt[15] , n_9562, n_9563, n14325);
  and g42450 (n16801, \asqrt[12] , n_10794, n_10795, n16161);
  and g42451 (n18781, \asqrt[9] , n_12098, n_12099, n18105);
  and g42452 (n20869, \asqrt[6] , n_13474, n_13475, n20157);
  and g42453 (n23042, \asqrt[3] , n_14920, n_14921, n22302);
  and g42454 (n7225, \asqrt[30] , n_4507, n6801, n_4506);
  and g42455 (n7237, \asqrt[30] , n_4514, n_4515, n6813);
  and g42456 (n7249, \asqrt[30] , n_4523, n6825, n_4522);
  and g42457 (n7261, \asqrt[30] , n_4530, n_4531, n6837);
  and g42458 (n7273, \asqrt[30] , n_4539, n6849, n_4538);
  and g42459 (n6857, \asqrt[31] , n_4266, n_4267, n6444);
  and g42460 (n6869, \asqrt[31] , n_4275, n6456, n_4274);
  and g42461 (n6881, \asqrt[31] , n_4282, n_4283, n6468);
  and g42462 (n6893, \asqrt[31] , n_4291, n6480, n_4290);
  and g42463 (n6905, \asqrt[31] , n_4298, n_4299, n6492);
  and g42464 (n6917, \asqrt[31] , n_4307, n6504, n_4306);
  and g42465 (n6929, \asqrt[31] , n_4314, n_4315, n6516);
  and g42466 (n6941, \asqrt[31] , n_4323, n6528, n_4322);
  and g42467 (n6953, \asqrt[31] , n_4330, n_4331, n6540);
  and g42468 (n6965, \asqrt[31] , n_4339, n6552, n_4338);
  and g42469 (n6977, \asqrt[31] , n_4346, n_4347, n6564);
  and g42470 (n6989, \asqrt[31] , n_4355, n6576, n_4354);
  and g42471 (n7001, \asqrt[31] , n_4362, n_4363, n6588);
  and g42472 (n7013, \asqrt[31] , n_4371, n6600, n_4370);
  and g42473 (n7025, \asqrt[31] , n_4378, n_4379, n6612);
  and g42474 (n7037, \asqrt[31] , n_4387, n6624, n_4386);
  and g42475 (n7049, \asqrt[31] , n_4394, n_4395, n6636);
  and g42476 (n7061, \asqrt[31] , n_4403, n6648, n_4402);
  and g42477 (n7073, \asqrt[31] , n_4410, n_4411, n6660);
  and g42478 (n7085, \asqrt[31] , n_4419, n6672, n_4418);
  and g42479 (n7097, \asqrt[31] , n_4426, n_4427, n6684);
  and g42480 (n7109, \asqrt[31] , n_4435, n6696, n_4434);
  and g42481 (n7121, \asqrt[31] , n_4442, n_4443, n6708);
  and g42482 (n7132, \asqrt[31] , n_4451, n6720, n_4450);
  and g42484 (n_16959, n_4463, n_4455);
  and g42485 (n7153, n_4454, n_4464, n_16958, n_16959);
  and g42486 (n1799, \asqrt[48] , n_986, n_987, n1591);
  and g42487 (n2496, \asqrt[45] , n_1435, n2252, n_1434);
  and g42488 (n3300, \asqrt[42] , n_1954, n_1955, n3020);
  and g42489 (n4212, \asqrt[39] , n_2547, n3896, n_2546);
  and g42490 (n5596, n_16960, n_3690, n_3689, n_3457);
  not g42491 (n_16960, n5593);
  and g42493 (n_16962, n_3455, n_3447);
  and g42494 (n5608, n_3446, n_3456, n_16961, n_16962);
  and g42495 (n7141, n_16963, n_4730, n_4729, n_4465);
  not g42496 (n_16963, n7138);
  or g42497 (\asqrt[33] , n5967, n5971, n5976, n5965);
  or g42501 (\asqrt[31] , n6739, n6743, n6748, n6737);
  and g42505 (n23793, \asqrt[2] , n_15416, n23034, n_15415);
  and g42506 (n21578, \asqrt[5] , n_13947, n20861, n_13946);
  and g42507 (n19461, \asqrt[8] , n_12547, n18773, n_12546);
  and g42508 (n17445, \asqrt[11] , n_11219, n16793, n_11218);
  and g42509 (n15537, \asqrt[14] , n_9963, n14921, n_9962);
  and g42510 (n13737, \asqrt[17] , n_8779, n13157, n_8778);
  and g42511 (n12045, \asqrt[20] , n_7667, n11501, n_7666);
  and g42512 (n10461, \asqrt[23] , n_6627, n9953, n_6626);
  and g42513 (n8985, \asqrt[26] , n_5659, n8513, n_5658);
  and g42514 (n7617, \asqrt[29] , n_4762, n_4760, n7184);
  and g42515 (n1587, \asqrt[49] , n_850, n_851, n1391);
  and g42516 (n2248, \asqrt[46] , n_1275, n2016, n_1274);
  and g42517 (n3016, \asqrt[43] , n_1770, n_1771, n2748);
  and g42518 (n3892, \asqrt[40] , n_2339, n3588, n_2338);
  and g42519 (n4876, \asqrt[37] , n_2978, n_2979, n4536);
  and g42520 (n5231, \asqrt[36] , n_3210, n_3211, n4880);
  and g42521 (n_16958, n_4483, n_4465);
  and g42522 (n6774, n_4463, \asqrt[32] , n_4464, n_16958);
  and g42523 (n_16971, n_4208, n_3963);
  and g42524 (n_16972, n_3945, n_3943);
  and g42525 (n6373, n_3944, n_4209, n_16971, n_16972);
  and g42526 (n8057, \asqrt[28] , n_5050, n_5051, n7609);
  and g42527 (n9461, \asqrt[25] , n_5970, n_5971, n8977);
  and g42528 (n10973, \asqrt[22] , n_6962, n_6963, n10453);
  and g42529 (n12593, \asqrt[19] , n_8026, n_8027, n12037);
  and g42530 (n14321, \asqrt[16] , n_9162, n_9163, n13729);
  and g42531 (n16157, \asqrt[13] , n_10370, n_10371, n15529);
  and g42532 (n18101, \asqrt[10] , n_11650, n_11651, n17437);
  and g42533 (n20153, \asqrt[7] , n_13002, n_13003, n19453);
  and g42534 (n22298, \asqrt[4] , n_14425, n_14426, n21570);
  and g42535 (n24131, \asqrt[1] , n_15921, n_15922, n23785);
  and g42536 (n6797, \asqrt[31] , n_4226, n_4224, n6387);
  and g42537 (n6809, \asqrt[31] , n_4234, n_4235, n6396);
  and g42538 (n6821, \asqrt[31] , n_4243, n6408, n_4242);
  and g42539 (n6833, \asqrt[31] , n_4250, n_4251, n6420);
  and g42540 (n6845, \asqrt[31] , n_4259, n6432, n_4258);
  and g42541 (n6440, \asqrt[32] , n_3994, n_3995, n6040);
  and g42542 (n6452, \asqrt[32] , n_4003, n6052, n_4002);
  and g42543 (n6464, \asqrt[32] , n_4010, n_4011, n6064);
  and g42544 (n6476, \asqrt[32] , n_4019, n6076, n_4018);
  and g42545 (n6488, \asqrt[32] , n_4026, n_4027, n6088);
  and g42546 (n6500, \asqrt[32] , n_4035, n6100, n_4034);
  and g42547 (n6512, \asqrt[32] , n_4042, n_4043, n6112);
  and g42548 (n6524, \asqrt[32] , n_4051, n6124, n_4050);
  and g42549 (n6536, \asqrt[32] , n_4058, n_4059, n6136);
  and g42550 (n6548, \asqrt[32] , n_4067, n6148, n_4066);
  and g42551 (n6560, \asqrt[32] , n_4074, n_4075, n6160);
  and g42552 (n6572, \asqrt[32] , n_4083, n6172, n_4082);
  and g42553 (n6584, \asqrt[32] , n_4090, n_4091, n6184);
  and g42554 (n6596, \asqrt[32] , n_4099, n6196, n_4098);
  and g42555 (n6608, \asqrt[32] , n_4106, n_4107, n6208);
  and g42556 (n6620, \asqrt[32] , n_4115, n6220, n_4114);
  and g42557 (n6632, \asqrt[32] , n_4122, n_4123, n6232);
  and g42558 (n6644, \asqrt[32] , n_4131, n6244, n_4130);
  and g42559 (n6656, \asqrt[32] , n_4138, n_4139, n6256);
  and g42560 (n6668, \asqrt[32] , n_4147, n6268, n_4146);
  and g42561 (n6680, \asqrt[32] , n_4154, n_4155, n6280);
  and g42562 (n6692, \asqrt[32] , n_4163, n6292, n_4162);
  and g42563 (n6704, \asqrt[32] , n_4170, n_4171, n6304);
  and g42564 (n6716, \asqrt[32] , n_4179, n6316, n_4178);
  and g42565 (n6727, \asqrt[32] , n_4186, n_4187, n6328);
  and g42567 (n_16974, n_4199, n_4191);
  and g42568 (n6748, n_4190, n_4200, n_16973, n_16974);
  and g42569 (n_16975, n_712, n_619);
  and g42570 (n_16976, n_601, n_599);
  and g42571 (n1200, n_600, n_713, n_16975, n_16976);
  and g42572 (n_16749, n_723, n_705);
  and g42573 (n1213, n_703, \asqrt[52] , n_704, n_16749);
  and g42574 (n2012, \asqrt[47] , n_1123, n1791, n_1122);
  and g42575 (n2744, \asqrt[44] , n_1594, n_1595, n2488);
  and g42576 (n3584, \asqrt[41] , n_2139, n3292, n_2138);
  and g42577 (n4532, \asqrt[38] , n_2754, n_2755, n4204);
  and g42578 (n5964, n_16978, n_3938, n_3937, n_3697);
  not g42579 (n_16978, n5961);
  and g42581 (n_16980, n_3695, n_3687);
  and g42582 (n5976, n_3686, n_3696, n_16979, n_16980);
  or g42583 (\asqrt[32] , n6347, n6351, n6356, n6345);
  and g42587 (n6736, n_16984, n_4458, n_4457, n_4201);
  not g42588 (n_16984, n6733);
  and g42589 (n_16985, n_4472, n_4219);
  and g42590 (n_16986, n_4201, n_4199);
  and g42591 (n6761, n_4200, n_4473, n_16985, n_16986);
  and g42592 (n23030, \asqrt[3] , n_14913, n22290, n_14912);
  and g42593 (n20857, \asqrt[6] , n_13467, n20145, n_13466);
  and g42594 (n18769, \asqrt[9] , n_12091, n18093, n_12090);
  and g42595 (n16789, \asqrt[12] , n_10787, n16149, n_10786);
  and g42596 (n14917, \asqrt[15] , n_9555, n14313, n_9554);
  and g42597 (n13153, \asqrt[18] , n_8395, n12585, n_8394);
  and g42598 (n11497, \asqrt[21] , n_7307, n10965, n_7306);
  and g42599 (n9949, \asqrt[24] , n_6291, n9453, n_6290);
  and g42600 (n8509, \asqrt[27] , n_5347, n8049, n_5346);
  and g42601 (n1787, \asqrt[48] , n_979, n1579, n_978);
  and g42602 (n2484, \asqrt[45] , n_1426, n_1427, n2240);
  and g42603 (n3288, \asqrt[42] , n_1947, n3008, n_1946);
  and g42604 (n4200, \asqrt[39] , n_2538, n_2539, n3884);
  and g42605 (n5220, \asqrt[36] , n_3203, n4868, n_3202);
  and g42606 (n5587, \asqrt[35] , n_3443, n5224, n_3442);
  and g42607 (n8973, \asqrt[26] , n_5650, n_5651, n8501);
  and g42608 (n10449, \asqrt[23] , n_6618, n_6619, n9941);
  and g42609 (n12033, \asqrt[20] , n_7658, n_7659, n11489);
  and g42610 (n13725, \asqrt[17] , n_8770, n_8771, n13145);
  and g42611 (n15525, \asqrt[14] , n_9954, n_9955, n14909);
  and g42612 (n17433, \asqrt[11] , n_11210, n_11211, n16781);
  and g42613 (n19449, \asqrt[8] , n_12538, n_12539, n18761);
  and g42614 (n21566, \asqrt[5] , n_13938, n_13939, n20849);
  and g42615 (n23781, \asqrt[2] , n_15407, n_15408, n23022);
  and g42616 (n6404, \asqrt[32] , n_3970, n_3968, n6007);
  and g42617 (n6416, \asqrt[32] , n_3978, n_3979, n6016);
  and g42618 (n6428, \asqrt[32] , n_3987, n6028, n_3986);
  and g42619 (n6036, \asqrt[33] , n_3730, n_3731, n5648);
  and g42620 (n6048, \asqrt[33] , n_3739, n5660, n_3738);
  and g42621 (n6060, \asqrt[33] , n_3746, n_3747, n5672);
  and g42622 (n6072, \asqrt[33] , n_3755, n5684, n_3754);
  and g42623 (n6084, \asqrt[33] , n_3762, n_3763, n5696);
  and g42624 (n6096, \asqrt[33] , n_3771, n5708, n_3770);
  and g42625 (n6108, \asqrt[33] , n_3778, n_3779, n5720);
  and g42626 (n6120, \asqrt[33] , n_3787, n5732, n_3786);
  and g42627 (n6132, \asqrt[33] , n_3794, n_3795, n5744);
  and g42628 (n6144, \asqrt[33] , n_3803, n5756, n_3802);
  and g42629 (n6156, \asqrt[33] , n_3810, n_3811, n5768);
  and g42630 (n6168, \asqrt[33] , n_3819, n5780, n_3818);
  and g42631 (n6180, \asqrt[33] , n_3826, n_3827, n5792);
  and g42632 (n6192, \asqrt[33] , n_3835, n5804, n_3834);
  and g42633 (n6204, \asqrt[33] , n_3842, n_3843, n5816);
  and g42634 (n6216, \asqrt[33] , n_3851, n5828, n_3850);
  and g42635 (n6228, \asqrt[33] , n_3858, n_3859, n5840);
  and g42636 (n6240, \asqrt[33] , n_3867, n5852, n_3866);
  and g42637 (n6252, \asqrt[33] , n_3874, n_3875, n5864);
  and g42638 (n6264, \asqrt[33] , n_3883, n5876, n_3882);
  and g42639 (n6276, \asqrt[33] , n_3890, n_3891, n5888);
  and g42640 (n6288, \asqrt[33] , n_3899, n5900, n_3898);
  and g42641 (n6300, \asqrt[33] , n_3906, n_3907, n5912);
  and g42642 (n6312, \asqrt[33] , n_3915, n5924, n_3914);
  and g42643 (n6324, \asqrt[33] , n_3922, n_3923, n5936);
  and g42644 (n6335, \asqrt[33] , n_3931, n5948, n_3930);
  and g42646 (n_16988, n_3943, n_3935);
  and g42647 (n6356, n_3934, n_3944, n_16987, n_16988);
  and g42648 (n1575, \asqrt[49] , n_842, n_840, n1382);
  and g42649 (n2236, \asqrt[46] , n_1266, n_1267, n2004);
  and g42650 (n3004, \asqrt[43] , n_1763, n2736, n_1762);
  and g42651 (n3880, \asqrt[40] , n_2330, n_2331, n3576);
  and g42652 (n4864, \asqrt[37] , n_2971, n4524, n_2970);
  and g42653 (n6344, n_16989, n_4194, n_4193, n_3945);
  not g42654 (n_16989, n6341);
  and g42655 (n24607, \asqrt[1] , n_15914, n23773, n_15913);
  and g42656 (n22286, \asqrt[4] , n_14418, n21558, n_14417);
  and g42657 (n20141, \asqrt[7] , n_12995, n19441, n_12994);
  and g42658 (n18089, \asqrt[10] , n_11643, n17425, n_11642);
  and g42659 (n16145, \asqrt[13] , n_10363, n15517, n_10362);
  and g42660 (n14309, \asqrt[16] , n_9155, n13717, n_9154);
  and g42661 (n12581, \asqrt[19] , n_8019, n12025, n_8018);
  and g42662 (n10961, \asqrt[22] , n_6955, n10441, n_6954);
  and g42663 (n9449, \asqrt[25] , n_5963, n8965, n_5962);
  and g42664 (n8045, \asqrt[28] , n_5042, n_5040, n7600);
  and g42665 (n_16945, n_4755, n_4737);
  and g42666 (n7179, n_4735, \asqrt[31] , n_4736, n_16945);
  and g42667 (n2000, \asqrt[47] , n_1114, n_1115, n1779);
  and g42668 (n2732, \asqrt[44] , n_1587, n2476, n_1586);
  and g42669 (n3572, \asqrt[41] , n_2130, n_2131, n3280);
  and g42670 (n4520, \asqrt[38] , n_2747, n4192, n_2746);
  and g42671 (n5578, \asqrt[35] , n_3433, n_3435, n5214);
  and g42672 (n5955, \asqrt[34] , n_3681, n_3683, n5582);
  and g42673 (n8497, \asqrt[27] , n_5338, n_5339, n8037);
  and g42674 (n9937, \asqrt[24] , n_6282, n_6283, n9441);
  and g42675 (n11485, \asqrt[21] , n_7298, n_7299, n10953);
  and g42676 (n13141, \asqrt[18] , n_8386, n_8387, n12573);
  and g42677 (n14905, \asqrt[15] , n_9546, n_9547, n14301);
  and g42678 (n16777, \asqrt[12] , n_10778, n_10779, n16137);
  and g42679 (n18757, \asqrt[9] , n_12082, n_12083, n18081);
  and g42680 (n20845, \asqrt[6] , n_13458, n_13459, n20133);
  and g42681 (n23018, \asqrt[3] , n_14904, n_14905, n22278);
  and g42682 (n_16973, n_4219, n_4201);
  and g42683 (n6382, n_4199, \asqrt[33] , n_4200, n_16973);
  and g42684 (n6024, \asqrt[33] , n_3722, n_3720, n5639);
  and g42685 (n5656, \asqrt[34] , n_3482, n_3480, n5283);
  and g42686 (n5668, \asqrt[34] , n_3490, n_3491, n5292);
  and g42687 (n5680, \asqrt[34] , n_3499, n5304, n_3498);
  and g42688 (n5692, \asqrt[34] , n_3506, n_3507, n5316);
  and g42689 (n5704, \asqrt[34] , n_3515, n5328, n_3514);
  and g42690 (n5716, \asqrt[34] , n_3522, n_3523, n5340);
  and g42691 (n5728, \asqrt[34] , n_3531, n5352, n_3530);
  and g42692 (n5740, \asqrt[34] , n_3538, n_3539, n5364);
  and g42693 (n5752, \asqrt[34] , n_3547, n5376, n_3546);
  and g42694 (n5764, \asqrt[34] , n_3554, n_3555, n5388);
  and g42695 (n5776, \asqrt[34] , n_3563, n5400, n_3562);
  and g42696 (n5788, \asqrt[34] , n_3570, n_3571, n5412);
  and g42697 (n5800, \asqrt[34] , n_3579, n5424, n_3578);
  and g42698 (n5812, \asqrt[34] , n_3586, n_3587, n5436);
  and g42699 (n5824, \asqrt[34] , n_3595, n5448, n_3594);
  and g42700 (n5836, \asqrt[34] , n_3602, n_3603, n5460);
  and g42701 (n5848, \asqrt[34] , n_3611, n5472, n_3610);
  and g42702 (n5860, \asqrt[34] , n_3618, n_3619, n5484);
  and g42703 (n5872, \asqrt[34] , n_3627, n5496, n_3626);
  and g42704 (n5884, \asqrt[34] , n_3634, n_3635, n5508);
  and g42705 (n5896, \asqrt[34] , n_3643, n5520, n_3642);
  and g42706 (n5908, \asqrt[34] , n_3650, n_3651, n5532);
  and g42707 (n5920, \asqrt[34] , n_3659, n5544, n_3658);
  and g42708 (n5932, \asqrt[34] , n_3666, n_3667, n5556);
  and g42709 (n5944, \asqrt[34] , n_3675, n5568, n_3674);
  and g42710 (n1775, \asqrt[48] , n_970, n_971, n1567);
  and g42711 (n2472, \asqrt[45] , n_1419, n2228, n_1418);
  and g42712 (n3276, \asqrt[42] , n_1938, n_1939, n2996);
  and g42713 (n4188, \asqrt[39] , n_2531, n3872, n_2530);
  and g42714 (n5210, \asqrt[36] , n_3193, n_3195, n4858);
  and g42715 (n_16992, n_4744, n_4483);
  and g42716 (n_16993, n_4465, n_4463);
  and g42717 (n7166, n_4464, n_4745, n_16992, n_16993);
  and g42718 (n23769, \asqrt[2] , n_15400, n23010, n_15399);
  and g42719 (n21554, \asqrt[5] , n_13931, n20837, n_13930);
  and g42720 (n19437, \asqrt[8] , n_12531, n18749, n_12530);
  and g42721 (n17421, \asqrt[11] , n_11203, n16769, n_11202);
  and g42722 (n15513, \asqrt[14] , n_9947, n14897, n_9946);
  and g42723 (n13713, \asqrt[17] , n_8763, n13133, n_8762);
  and g42724 (n12021, \asqrt[20] , n_7651, n11477, n_7650);
  and g42725 (n10437, \asqrt[23] , n_6611, n9929, n_6610);
  and g42726 (n8961, \asqrt[26] , n_5643, n8489, n_5642);
  and g42727 (n_16994, n_3952, n_3715);
  and g42728 (n_16995, n_3697, n_3695);
  and g42729 (n5989, n_3696, n_3953, n_16994, n_16995);
  and g42730 (n_16996, n_824, n_723);
  and g42731 (n_16997, n_705, n_703);
  and g42732 (n1364, n_704, n_825, n_16996, n_16997);
  and g42733 (n_16761, n_835, n_817);
  and g42734 (n1377, n_815, \asqrt[51] , n_816, n_16761);
  and g42735 (n2224, \asqrt[46] , n_1259, n1992, n_1258);
  and g42736 (n2992, \asqrt[43] , n_1754, n_1755, n2724);
  and g42737 (n3868, \asqrt[40] , n_2323, n3564, n_2322);
  and g42738 (n4854, \asqrt[37] , n_2961, n_2963, n4514);
  and g42739 (n9437, \asqrt[25] , n_5954, n_5955, n8953);
  and g42740 (n10949, \asqrt[22] , n_6946, n_6947, n10429);
  and g42741 (n12569, \asqrt[19] , n_8010, n_8011, n12013);
  and g42742 (n14297, \asqrt[16] , n_9146, n_9147, n13705);
  and g42743 (n16133, \asqrt[13] , n_10354, n_10355, n15505);
  and g42744 (n18077, \asqrt[10] , n_11634, n_11635, n17413);
  and g42745 (n20129, \asqrt[7] , n_12986, n_12987, n19429);
  and g42746 (n22274, \asqrt[4] , n_14409, n_14410, n21546);
  and g42747 (n24138, \asqrt[1] , n_15905, n_15906, n23761);
  and g42748 (n_16987, n_3963, n_3945);
  and g42749 (n6002, n_3943, \asqrt[34] , n_3944, n_16987);
  and g42750 (n5300, \asqrt[35] , n_3250, n_3248, n4939);
  and g42751 (n5312, \asqrt[35] , n_3258, n_3259, n4948);
  and g42752 (n5324, \asqrt[35] , n_3267, n4960, n_3266);
  and g42753 (n5336, \asqrt[35] , n_3274, n_3275, n4972);
  and g42754 (n5348, \asqrt[35] , n_3283, n4984, n_3282);
  and g42755 (n5360, \asqrt[35] , n_3290, n_3291, n4996);
  and g42756 (n5372, \asqrt[35] , n_3299, n5008, n_3298);
  and g42757 (n5384, \asqrt[35] , n_3306, n_3307, n5020);
  and g42758 (n5396, \asqrt[35] , n_3315, n5032, n_3314);
  and g42759 (n5408, \asqrt[35] , n_3322, n_3323, n5044);
  and g42760 (n5420, \asqrt[35] , n_3331, n5056, n_3330);
  and g42761 (n5432, \asqrt[35] , n_3338, n_3339, n5068);
  and g42762 (n5444, \asqrt[35] , n_3347, n5080, n_3346);
  and g42763 (n5456, \asqrt[35] , n_3354, n_3355, n5092);
  and g42764 (n5468, \asqrt[35] , n_3363, n5104, n_3362);
  and g42765 (n5480, \asqrt[35] , n_3370, n_3371, n5116);
  and g42766 (n5492, \asqrt[35] , n_3379, n5128, n_3378);
  and g42767 (n5504, \asqrt[35] , n_3386, n_3387, n5140);
  and g42768 (n5516, \asqrt[35] , n_3395, n5152, n_3394);
  and g42769 (n5528, \asqrt[35] , n_3402, n_3403, n5164);
  and g42770 (n5540, \asqrt[35] , n_3411, n5176, n_3410);
  and g42771 (n5552, \asqrt[35] , n_3418, n_3419, n5188);
  and g42772 (n5564, \asqrt[35] , n_3427, n5200, n_3426);
  and g42773 (n1988, \asqrt[47] , n_1107, n1767, n_1106);
  and g42774 (n2720, \asqrt[44] , n_1578, n_1579, n2464);
  and g42775 (n3560, \asqrt[41] , n_2123, n3268, n_2122);
  and g42776 (n4510, \asqrt[38] , n_2737, n_2739, n4182);
  and g42777 (n23006, \asqrt[3] , n_14897, n22266, n_14896);
  and g42778 (n20833, \asqrt[6] , n_13451, n20121, n_13450);
  and g42779 (n18745, \asqrt[9] , n_12075, n18069, n_12074);
  and g42780 (n16765, \asqrt[12] , n_10771, n16125, n_10770);
  and g42781 (n14893, \asqrt[15] , n_9539, n14289, n_9538);
  and g42782 (n13129, \asqrt[18] , n_8379, n12561, n_8378);
  and g42783 (n11473, \asqrt[21] , n_7291, n10941, n_7290);
  and g42784 (n9925, \asqrt[24] , n_6275, n9429, n_6274);
  and g42785 (n8485, \asqrt[27] , n_5330, n_5328, n8028);
  and g42786 (n_16930, n_5035, n_5017);
  and g42787 (n7595, n_5015, \asqrt[30] , n_5016, n_16930);
  and g42788 (n_17001, n_3704, n_3475);
  and g42789 (n_17002, n_3457, n_3455);
  and g42790 (n5621, n_3456, n_3705, n_17001, n_17002);
  and g42791 (n_17003, n_3464, n_3243);
  and g42792 (n_17004, n_3225, n_3223);
  and g42793 (n5265, n_3224, n_3465, n_17003, n_17004);
  and g42794 (n1763, \asqrt[48] , n_962, n_960, n1558);
  and g42795 (n2460, \asqrt[45] , n_1410, n_1411, n2216);
  and g42796 (n3264, \asqrt[42] , n_1931, n2984, n_1930);
  and g42797 (n4178, \asqrt[39] , n_2521, n_2523, n3862);
  and g42798 (n5196, \asqrt[36] , n_3187, n4844, n_3186);
  and g42799 (n8949, \asqrt[26] , n_5634, n_5635, n8477);
  and g42800 (n10425, \asqrt[23] , n_6602, n_6603, n9917);
  and g42801 (n12009, \asqrt[20] , n_7642, n_7643, n11465);
  and g42802 (n13701, \asqrt[17] , n_8754, n_8755, n13121);
  and g42803 (n15501, \asqrt[14] , n_9938, n_9939, n14885);
  and g42804 (n17409, \asqrt[11] , n_11194, n_11195, n16757);
  and g42805 (n19425, \asqrt[8] , n_12522, n_12523, n18737);
  and g42806 (n21542, \asqrt[5] , n_13922, n_13923, n20825);
  and g42807 (n23757, \asqrt[2] , n_15391, n_15392, n22998);
  and g42808 (n_16979, n_3715, n_3697);
  and g42809 (n5634, n_3695, \asqrt[35] , n_3696, n_16979);
  and g42810 (n_16961, n_3475, n_3457);
  and g42811 (n5278, n_3455, \asqrt[36] , n_3456, n_16961);
  and g42812 (n4956, \asqrt[36] , n_3026, n_3024, n4607);
  and g42813 (n4968, \asqrt[36] , n_3034, n_3035, n4616);
  and g42814 (n4980, \asqrt[36] , n_3043, n4628, n_3042);
  and g42815 (n4992, \asqrt[36] , n_3050, n_3051, n4640);
  and g42816 (n5004, \asqrt[36] , n_3059, n4652, n_3058);
  and g42817 (n5016, \asqrt[36] , n_3066, n_3067, n4664);
  and g42818 (n5028, \asqrt[36] , n_3075, n4676, n_3074);
  and g42819 (n5040, \asqrt[36] , n_3082, n_3083, n4688);
  and g42820 (n5052, \asqrt[36] , n_3091, n4700, n_3090);
  and g42821 (n5064, \asqrt[36] , n_3098, n_3099, n4712);
  and g42822 (n5076, \asqrt[36] , n_3107, n4724, n_3106);
  and g42823 (n5088, \asqrt[36] , n_3114, n_3115, n4736);
  and g42824 (n5100, \asqrt[36] , n_3123, n4748, n_3122);
  and g42825 (n5112, \asqrt[36] , n_3130, n_3131, n4760);
  and g42826 (n5124, \asqrt[36] , n_3139, n4772, n_3138);
  and g42827 (n5136, \asqrt[36] , n_3146, n_3147, n4784);
  and g42828 (n5148, \asqrt[36] , n_3155, n4796, n_3154);
  and g42829 (n5160, \asqrt[36] , n_3162, n_3163, n4808);
  and g42830 (n5172, \asqrt[36] , n_3171, n4820, n_3170);
  and g42831 (n5184, \asqrt[36] , n_3178, n_3179, n4832);
  and g42832 (n2212, \asqrt[46] , n_1250, n_1251, n1980);
  and g42833 (n2980, \asqrt[43] , n_1747, n2712, n_1746);
  and g42834 (n3858, \asqrt[40] , n_2313, n_2315, n3554);
  and g42835 (n4840, \asqrt[37] , n_2955, n4500, n_2954);
  and g42836 (n_17007, n_5024, n_4755);
  and g42837 (n_17008, n_4737, n_4735);
  and g42838 (n7582, n_4736, n_5025, n_17007, n_17008);
  and g42839 (n24590, \asqrt[1] , n_15898, n23749, n_15897);
  and g42840 (n22262, \asqrt[4] , n_14402, n21534, n_14401);
  and g42841 (n20117, \asqrt[7] , n_12979, n19417, n_12978);
  and g42842 (n18065, \asqrt[10] , n_11627, n17401, n_11626);
  and g42843 (n16121, \asqrt[13] , n_10347, n15493, n_10346);
  and g42844 (n14285, \asqrt[16] , n_9139, n13693, n_9138);
  and g42845 (n12557, \asqrt[19] , n_8003, n12001, n_8002);
  and g42846 (n10937, \asqrt[22] , n_6939, n10417, n_6938);
  and g42847 (n9425, \asqrt[25] , n_5947, n8941, n_5946);
  and g42848 (n_17009, n_3232, n_3019);
  and g42849 (n_17010, n_3001, n_2999);
  and g42850 (n4921, n_3000, n_3233, n_17009, n_17010);
  and g42851 (n1976, \asqrt[47] , n_1098, n_1099, n1755);
  and g42852 (n2708, \asqrt[44] , n_1571, n2452, n_1570);
  and g42853 (n3550, \asqrt[41] , n_2113, n_2115, n3258);
  and g42854 (n4496, \asqrt[38] , n_2731, n4168, n_2730);
  and g42855 (n9913, \asqrt[24] , n_6266, n_6267, n9417);
  and g42856 (n11461, \asqrt[21] , n_7282, n_7283, n10929);
  and g42857 (n13117, \asqrt[18] , n_8370, n_8371, n12549);
  and g42858 (n14881, \asqrt[15] , n_9530, n_9531, n14277);
  and g42859 (n16753, \asqrt[12] , n_10762, n_10763, n16113);
  and g42860 (n18733, \asqrt[9] , n_12066, n_12067, n18057);
  and g42861 (n20821, \asqrt[6] , n_13442, n_13443, n20109);
  and g42862 (n22994, \asqrt[3] , n_14888, n_14889, n22254);
  and g42863 (n_16948, n_3243, n_3225);
  and g42864 (n4934, n_3223, \asqrt[37] , n_3224, n_16948);
  and g42865 (n4624, \asqrt[37] , n_2810, n_2808, n4287);
  and g42866 (n4636, \asqrt[37] , n_2818, n_2819, n4296);
  and g42867 (n4648, \asqrt[37] , n_2827, n4308, n_2826);
  and g42868 (n4660, \asqrt[37] , n_2834, n_2835, n4320);
  and g42869 (n4672, \asqrt[37] , n_2843, n4332, n_2842);
  and g42870 (n4684, \asqrt[37] , n_2850, n_2851, n4344);
  and g42871 (n4696, \asqrt[37] , n_2859, n4356, n_2858);
  and g42872 (n4708, \asqrt[37] , n_2866, n_2867, n4368);
  and g42873 (n4720, \asqrt[37] , n_2875, n4380, n_2874);
  and g42874 (n4732, \asqrt[37] , n_2882, n_2883, n4392);
  and g42875 (n4744, \asqrt[37] , n_2891, n4404, n_2890);
  and g42876 (n4756, \asqrt[37] , n_2898, n_2899, n4416);
  and g42877 (n4768, \asqrt[37] , n_2907, n4428, n_2906);
  and g42878 (n4780, \asqrt[37] , n_2914, n_2915, n4440);
  and g42879 (n4792, \asqrt[37] , n_2923, n4452, n_2922);
  and g42880 (n4804, \asqrt[37] , n_2930, n_2931, n4464);
  and g42881 (n4816, \asqrt[37] , n_2939, n4476, n_2938);
  and g42882 (n4828, \asqrt[37] , n_2946, n_2947, n4488);
  and g42883 (n_17012, n_944, n_835);
  and g42884 (n_17013, n_817, n_815);
  and g42885 (n1540, n_816, n_945, n_17012, n_17013);
  and g42886 (n_16776, n_955, n_937);
  and g42887 (n1553, n_935, \asqrt[50] , n_936, n_16776);
  and g42888 (n2448, \asqrt[45] , n_1403, n2204, n_1402);
  and g42889 (n3254, \asqrt[42] , n_1921, n_1923, n2974);
  and g42890 (n4164, \asqrt[39] , n_2515, n3848, n_2514);
  and g42891 (n23745, \asqrt[2] , n_15384, n22986, n_15383);
  and g42892 (n21530, \asqrt[5] , n_13915, n20813, n_13914);
  and g42893 (n19413, \asqrt[8] , n_12515, n18725, n_12514);
  and g42894 (n17397, \asqrt[11] , n_11187, n16745, n_11186);
  and g42895 (n15489, \asqrt[14] , n_9931, n14873, n_9930);
  and g42896 (n13689, \asqrt[17] , n_8747, n13109, n_8746);
  and g42897 (n11997, \asqrt[20] , n_7635, n11453, n_7634);
  and g42898 (n10413, \asqrt[23] , n_6595, n9905, n_6594);
  and g42899 (n8937, \asqrt[26] , n_5626, n_5624, n8468);
  and g42900 (n_16918, n_5323, n_5305);
  and g42901 (n8023, n_5303, \asqrt[29] , n_5304, n_16918);
  and g42902 (n_17016, n_3008, n_2803);
  and g42903 (n_17017, n_2785, n_2783);
  and g42904 (n4589, n_2784, n_3009, n_17016, n_17017);
  and g42905 (n2200, \asqrt[46] , n_1243, n1968, n_1242);
  and g42906 (n2970, \asqrt[43] , n_1737, n_1739, n2702);
  and g42907 (n3844, \asqrt[40] , n_2307, n3540, n_2306);
  and g42908 (n9413, \asqrt[25] , n_5938, n_5939, n8929);
  and g42909 (n10925, \asqrt[22] , n_6930, n_6931, n10405);
  and g42910 (n12545, \asqrt[19] , n_7994, n_7995, n11989);
  and g42911 (n14273, \asqrt[16] , n_9130, n_9131, n13681);
  and g42912 (n16109, \asqrt[13] , n_10338, n_10339, n15481);
  and g42913 (n18053, \asqrt[10] , n_11618, n_11619, n17389);
  and g42914 (n20105, \asqrt[7] , n_12970, n_12971, n19405);
  and g42915 (n22250, \asqrt[4] , n_14393, n_14394, n21522);
  and g42916 (n24145, \asqrt[1] , n_15889, n_15890, n23737);
  and g42917 (n_16933, n_3019, n_3001);
  and g42918 (n4602, n_2999, \asqrt[38] , n_3000, n_16933);
  and g42919 (n4304, \asqrt[38] , n_2602, n_2600, n3979);
  and g42920 (n4316, \asqrt[38] , n_2610, n_2611, n3988);
  and g42921 (n4328, \asqrt[38] , n_2619, n4000, n_2618);
  and g42922 (n4340, \asqrt[38] , n_2626, n_2627, n4012);
  and g42923 (n4352, \asqrt[38] , n_2635, n4024, n_2634);
  and g42924 (n4364, \asqrt[38] , n_2642, n_2643, n4036);
  and g42925 (n4376, \asqrt[38] , n_2651, n4048, n_2650);
  and g42926 (n4388, \asqrt[38] , n_2658, n_2659, n4060);
  and g42927 (n4400, \asqrt[38] , n_2667, n4072, n_2666);
  and g42928 (n4412, \asqrt[38] , n_2674, n_2675, n4084);
  and g42929 (n4424, \asqrt[38] , n_2683, n4096, n_2682);
  and g42930 (n4436, \asqrt[38] , n_2690, n_2691, n4108);
  and g42931 (n4448, \asqrt[38] , n_2699, n4120, n_2698);
  and g42932 (n4460, \asqrt[38] , n_2706, n_2707, n4132);
  and g42933 (n4472, \asqrt[38] , n_2715, n4144, n_2714);
  and g42934 (n4484, \asqrt[38] , n_2722, n_2723, n4156);
  and g42935 (n1964, \asqrt[47] , n_1090, n_1088, n1746);
  and g42936 (n2698, \asqrt[44] , n_1561, n_1563, n2442);
  and g42937 (n3536, \asqrt[41] , n_2107, n3244, n_2106);
  and g42938 (n_17019, n_5312, n_5035);
  and g42939 (n_17020, n_5017, n_5015);
  and g42940 (n8010, n_5016, n_5313, n_17019, n_17020);
  and g42941 (n22982, \asqrt[3] , n_14881, n22242, n_14880);
  and g42942 (n20809, \asqrt[6] , n_13435, n20097, n_13434);
  and g42943 (n18721, \asqrt[9] , n_12059, n18045, n_12058);
  and g42944 (n16741, \asqrt[12] , n_10755, n16101, n_10754);
  and g42945 (n14869, \asqrt[15] , n_9523, n14265, n_9522);
  and g42946 (n13105, \asqrt[18] , n_8363, n12537, n_8362);
  and g42947 (n11449, \asqrt[21] , n_7275, n10917, n_7274);
  and g42948 (n9901, \asqrt[24] , n_6259, n9405, n_6258);
  and g42949 (n_17021, n_2792, n_2595);
  and g42950 (n_17022, n_2577, n_2575);
  and g42951 (n4269, n_2576, n_2793, n_17021, n_17022);
  and g42952 (n2438, \asqrt[45] , n_1393, n_1395, n2194);
  and g42953 (n3240, \asqrt[42] , n_1915, n2960, n_1914);
  and g42954 (n4152, \asqrt[39] , n_2506, n_2507, n3836);
  and g42955 (n10401, \asqrt[23] , n_6586, n_6587, n9893);
  and g42956 (n11985, \asqrt[20] , n_7626, n_7627, n11441);
  and g42957 (n13677, \asqrt[17] , n_8738, n_8739, n13097);
  and g42958 (n15477, \asqrt[14] , n_9922, n_9923, n14861);
  and g42959 (n17385, \asqrt[11] , n_11178, n_11179, n16733);
  and g42960 (n19401, \asqrt[8] , n_12506, n_12507, n18713);
  and g42961 (n21518, \asqrt[5] , n_13906, n_13907, n20801);
  and g42962 (n23733, \asqrt[2] , n_15375, n_15376, n22974);
  and g42963 (n_16921, n_2803, n_2785);
  and g42964 (n4282, n_2783, \asqrt[39] , n_2784, n_16921);
  and g42965 (n3996, \asqrt[39] , n_2402, n_2400, n3683);
  and g42966 (n4008, \asqrt[39] , n_2410, n_2411, n3692);
  and g42967 (n4020, \asqrt[39] , n_2419, n3704, n_2418);
  and g42968 (n4032, \asqrt[39] , n_2426, n_2427, n3716);
  and g42969 (n4044, \asqrt[39] , n_2435, n3728, n_2434);
  and g42970 (n4056, \asqrt[39] , n_2442, n_2443, n3740);
  and g42971 (n4068, \asqrt[39] , n_2451, n3752, n_2450);
  and g42972 (n4080, \asqrt[39] , n_2458, n_2459, n3764);
  and g42973 (n4092, \asqrt[39] , n_2467, n3776, n_2466);
  and g42974 (n4104, \asqrt[39] , n_2474, n_2475, n3788);
  and g42975 (n4116, \asqrt[39] , n_2483, n3800, n_2482);
  and g42976 (n4128, \asqrt[39] , n_2490, n_2491, n3812);
  and g42977 (n4140, \asqrt[39] , n_2499, n3824, n_2498);
  and g42978 (n2190, \asqrt[46] , n_1233, n_1235, n1958);
  and g42979 (n2956, \asqrt[43] , n_1731, n2688, n_1730);
  and g42980 (n3832, \asqrt[40] , n_2298, n_2299, n3528);
  and g42981 (n24573, \asqrt[1] , n_15882, n23725, n_15881);
  and g42982 (n22238, \asqrt[4] , n_14386, n21510, n_14385);
  and g42983 (n20093, \asqrt[7] , n_12963, n19393, n_12962);
  and g42984 (n18041, \asqrt[10] , n_11611, n17377, n_11610);
  and g42985 (n16097, \asqrt[13] , n_10331, n15469, n_10330);
  and g42986 (n14261, \asqrt[16] , n_9123, n13669, n_9122);
  and g42987 (n12533, \asqrt[19] , n_7987, n11977, n_7986);
  and g42988 (n10913, \asqrt[22] , n_6923, n10393, n_6922);
  and g42989 (n9401, \asqrt[25] , n_5930, n_5928, n8920);
  and g42990 (n_16903, n_5619, n_5601);
  and g42991 (n8463, n_5599, \asqrt[28] , n_5600, n_16903);
  and g42992 (n_17025, n_2584, n_2395);
  and g42993 (n_17026, n_2377, n_2375);
  and g42994 (n3961, n_2376, n_2585, n_17025, n_17026);
  and g42995 (n_17027, n_1072, n_955);
  and g42996 (n_17028, n_937, n_935);
  and g42997 (n1732, n_936, n_1073, n_17027, n_17028);
  and g42998 (n_16788, n_1083, n_1065);
  and g42999 (n1741, n_1063, \asqrt[49] , n_1064, n_16788);
  and g43000 (n1954, n_17030, \asqrt[47] , n_1079, n_1078);
  not g43001 (n_17030, n1727);
  and g43002 (n2684, \asqrt[44] , n_1555, n2428, n_1554);
  and g43003 (n3524, \asqrt[41] , n_2098, n_2099, n3232);
  and g43004 (n9889, \asqrt[24] , n_6250, n_6251, n9393);
  and g43005 (n11437, \asqrt[21] , n_7266, n_7267, n10905);
  and g43006 (n13093, \asqrt[18] , n_8354, n_8355, n12525);
  and g43007 (n14857, \asqrt[15] , n_9514, n_9515, n14253);
  and g43008 (n16729, \asqrt[12] , n_10746, n_10747, n16089);
  and g43009 (n18709, \asqrt[9] , n_12050, n_12051, n18033);
  and g43010 (n20797, \asqrt[6] , n_13426, n_13427, n20085);
  and g43011 (n22970, \asqrt[3] , n_14872, n_14873, n22230);
  and g43012 (n_16909, n_2595, n_2577);
  and g43013 (n3974, n_2575, \asqrt[40] , n_2576, n_16909);
  and g43014 (n3700, \asqrt[40] , n_2210, n_2208, n3399);
  and g43015 (n3712, \asqrt[40] , n_2218, n_2219, n3408);
  and g43016 (n3724, \asqrt[40] , n_2227, n3420, n_2226);
  and g43017 (n3736, \asqrt[40] , n_2234, n_2235, n3432);
  and g43018 (n3748, \asqrt[40] , n_2243, n3444, n_2242);
  and g43019 (n3760, \asqrt[40] , n_2250, n_2251, n3456);
  and g43020 (n3772, \asqrt[40] , n_2259, n3468, n_2258);
  and g43021 (n3784, \asqrt[40] , n_2266, n_2267, n3480);
  and g43022 (n3796, \asqrt[40] , n_2275, n3492, n_2274);
  and g43023 (n3808, \asqrt[40] , n_2282, n_2283, n3504);
  and g43024 (n3820, \asqrt[40] , n_2291, n3516, n_2290);
  and g43025 (n2424, \asqrt[45] , n_1387, n2180, n_1386);
  and g43026 (n3228, \asqrt[42] , n_1906, n_1907, n2948);
  and g43027 (n_17032, n_5608, n_5323);
  and g43028 (n_17033, n_5305, n_5303);
  and g43029 (n8450, n_5304, n_5609, n_17032, n_17033);
  and g43030 (n23721, \asqrt[2] , n_15368, n22962, n_15367);
  and g43031 (n21506, \asqrt[5] , n_13899, n20789, n_13898);
  and g43032 (n19389, \asqrt[8] , n_12499, n18701, n_12498);
  and g43033 (n17373, \asqrt[11] , n_11171, n16721, n_11170);
  and g43034 (n15465, \asqrt[14] , n_9915, n14849, n_9914);
  and g43035 (n13665, \asqrt[17] , n_8731, n13085, n_8730);
  and g43036 (n11973, \asqrt[20] , n_7619, n11429, n_7618);
  and g43037 (n10389, \asqrt[23] , n_6579, n9881, n_6578);
  and g43038 (n_17034, n_2384, n_2203);
  and g43039 (n_17035, n_2185, n_2183);
  and g43040 (n3665, n_2184, n_2385, n_17034, n_17035);
  and g43041 (n2176, \asqrt[46] , n_1226, n_1224, n1946);
  and g43042 (n2944, \asqrt[43] , n_1722, n_1723, n2676);
  and g43043 (n10901, \asqrt[22] , n_6914, n_6915, n10381);
  and g43044 (n12521, \asqrt[19] , n_7978, n_7979, n11965);
  and g43045 (n14249, \asqrt[16] , n_9114, n_9115, n13657);
  and g43046 (n16085, \asqrt[13] , n_10322, n_10323, n15457);
  and g43047 (n18029, \asqrt[10] , n_11602, n_11603, n17365);
  and g43048 (n20081, \asqrt[7] , n_12954, n_12955, n19381);
  and g43049 (n22226, \asqrt[4] , n_14377, n_14378, n21498);
  and g43050 (n24152, \asqrt[1] , n_15873, n_15874, n23713);
  and g43051 (n_16894, n_2395, n_2377);
  and g43052 (n3678, n_2375, \asqrt[41] , n_2376, n_16894);
  and g43053 (n3416, \asqrt[41] , n_2026, n_2024, n3127);
  and g43054 (n3428, \asqrt[41] , n_2034, n_2035, n3136);
  and g43055 (n3440, \asqrt[41] , n_2043, n3148, n_2042);
  and g43056 (n3452, \asqrt[41] , n_2050, n_2051, n3160);
  and g43057 (n3464, \asqrt[41] , n_2059, n3172, n_2058);
  and g43058 (n3476, \asqrt[41] , n_2066, n_2067, n3184);
  and g43059 (n3488, \asqrt[41] , n_2075, n3196, n_2074);
  and g43060 (n3500, \asqrt[41] , n_2082, n_2083, n3208);
  and g43061 (n3512, \asqrt[41] , n_2091, n3220, n_2090);
  and g43062 (n2672, \asqrt[44] , n_1546, n_1547, n2416);
  and g43063 (n22958, \asqrt[3] , n_14865, n22218, n_14864);
  and g43064 (n20785, \asqrt[6] , n_13419, n20073, n_13418);
  and g43065 (n18697, \asqrt[9] , n_12043, n18021, n_12042);
  and g43066 (n16717, \asqrt[12] , n_10739, n16077, n_10738);
  and g43067 (n14845, \asqrt[15] , n_9507, n14241, n_9506);
  and g43068 (n13081, \asqrt[18] , n_8347, n12513, n_8346);
  and g43069 (n11425, \asqrt[21] , n_7259, n10893, n_7258);
  and g43070 (n9877, \asqrt[24] , n_6242, n_6240, n9384);
  and g43071 (n_16891, n_5923, n_5905);
  and g43072 (n8915, n_5903, \asqrt[27] , n_5904, n_16891);
  and g43073 (n_17038, n_2192, n_2019);
  and g43074 (n_17039, n_2001, n_1999);
  and g43075 (n3381, n_2000, n_2193, n_17038, n_17039);
  and g43076 (n2412, \asqrt[45] , n_1378, n_1379, n2168);
  and g43077 (n3216, \asqrt[42] , n_1899, n2936, n_1898);
  and g43078 (n10377, \asqrt[23] , n_6570, n_6571, n9869);
  and g43079 (n11961, \asqrt[20] , n_7610, n_7611, n11417);
  and g43080 (n13653, \asqrt[17] , n_8722, n_8723, n13073);
  and g43081 (n15453, \asqrt[14] , n_9906, n_9907, n14837);
  and g43082 (n17361, \asqrt[11] , n_11162, n_11163, n16709);
  and g43083 (n19377, \asqrt[8] , n_12490, n_12491, n18689);
  and g43084 (n21494, \asqrt[5] , n_13890, n_13891, n20777);
  and g43085 (n23709, \asqrt[2] , n_15359, n_15360, n22950);
  and g43086 (n_16882, n_2203, n_2185);
  and g43087 (n3394, n_2183, \asqrt[42] , n_2184, n_16882);
  and g43088 (n3144, \asqrt[42] , n_1850, n_1848, n2867);
  and g43089 (n3156, \asqrt[42] , n_1858, n_1859, n2876);
  and g43090 (n3168, \asqrt[42] , n_1867, n2888, n_1866);
  and g43091 (n3180, \asqrt[42] , n_1874, n_1875, n2900);
  and g43092 (n3192, \asqrt[42] , n_1883, n2912, n_1882);
  and g43093 (n3204, \asqrt[42] , n_1890, n_1891, n2924);
  and g43094 (n_17041, n_1208, n_1083);
  and g43095 (n_17042, n_1065, n_1063);
  and g43096 (n1928, n_1064, n_1209, n_17041, n_17042);
  and g43097 (n_16800, n_1219, n_1201);
  and g43098 (n1941, n_1199, \asqrt[48] , n_1200, n_16800);
  and g43099 (n2932, \asqrt[43] , n_1715, n2664, n_1714);
  and g43100 (n_17044, n_5912, n_5619);
  and g43101 (n_17045, n_5601, n_5599);
  and g43102 (n8902, n_5600, n_5913, n_17044, n_17045);
  and g43103 (n24556, \asqrt[1] , n_15866, n23701, n_15865);
  and g43104 (n22214, \asqrt[4] , n_14370, n21486, n_14369);
  and g43105 (n20069, \asqrt[7] , n_12947, n19369, n_12946);
  and g43106 (n18017, \asqrt[10] , n_11595, n17353, n_11594);
  and g43107 (n16073, \asqrt[13] , n_10315, n15445, n_10314);
  and g43108 (n14237, \asqrt[16] , n_9107, n13645, n_9106);
  and g43109 (n12509, \asqrt[19] , n_7971, n11953, n_7970);
  and g43110 (n10889, \asqrt[22] , n_6907, n10369, n_6906);
  and g43111 (n_17046, n_2008, n_1843);
  and g43112 (n_17047, n_1825, n_1823);
  and g43113 (n3109, n_1824, n_2009, n_17046, n_17047);
  and g43114 (n2660, \asqrt[44] , n_1539, n2404, n_1538);
  and g43115 (n11413, \asqrt[21] , n_7250, n_7251, n10881);
  and g43116 (n13069, \asqrt[18] , n_8338, n_8339, n12501);
  and g43117 (n14833, \asqrt[15] , n_9498, n_9499, n14229);
  and g43118 (n16705, \asqrt[12] , n_10730, n_10731, n16065);
  and g43119 (n18685, \asqrt[9] , n_12034, n_12035, n18009);
  and g43120 (n20773, \asqrt[6] , n_13410, n_13411, n20061);
  and g43121 (n22946, \asqrt[3] , n_14856, n_14857, n22206);
  and g43122 (n_16867, n_2019, n_2001);
  and g43123 (n3122, n_1999, \asqrt[43] , n_2000, n_16867);
  and g43124 (n2884, \asqrt[43] , n_1682, n_1680, n2619);
  and g43125 (n2896, \asqrt[43] , n_1690, n_1691, n2628);
  and g43126 (n2908, \asqrt[43] , n_1699, n2640, n_1698);
  and g43127 (n2920, \asqrt[43] , n_1706, n_1707, n2652);
  and g43128 (n2400, \asqrt[45] , n_1370, n_1368, n2159);
  and g43129 (n23697, \asqrt[2] , n_15352, n22938, n_15351);
  and g43130 (n21482, \asqrt[5] , n_13883, n20765, n_13882);
  and g43131 (n19365, \asqrt[8] , n_12483, n18677, n_12482);
  and g43132 (n17349, \asqrt[11] , n_11155, n16697, n_11154);
  and g43133 (n15441, \asqrt[14] , n_9899, n14825, n_9898);
  and g43134 (n13641, \asqrt[17] , n_8715, n13061, n_8714);
  and g43135 (n11949, \asqrt[20] , n_7603, n11405, n_7602);
  and g43136 (n10365, \asqrt[23] , n_6562, n_6560, n9860);
  and g43137 (n_16879, n_6235, n_6217);
  and g43138 (n9379, n_6215, \asqrt[26] , n_6216, n_16879);
  and g43139 (n_17050, n_1832, n_1675);
  and g43140 (n_17051, n_1657, n_1655);
  and g43141 (n2849, n_1656, n_1833, n_17050, n_17051);
  and g43142 (n10877, \asqrt[22] , n_6898, n_6899, n10357);
  and g43143 (n12497, \asqrt[19] , n_7962, n_7963, n11941);
  and g43144 (n14225, \asqrt[16] , n_9098, n_9099, n13633);
  and g43145 (n16061, \asqrt[13] , n_10306, n_10307, n15433);
  and g43146 (n18005, \asqrt[10] , n_11586, n_11587, n17341);
  and g43147 (n20057, \asqrt[7] , n_12938, n_12939, n19357);
  and g43148 (n22202, \asqrt[4] , n_14361, n_14362, n21474);
  and g43149 (n24159, \asqrt[1] , n_15857, n_15858, n23689);
  and g43150 (n_16855, n_1843, n_1825);
  and g43151 (n2862, n_1823, \asqrt[44] , n_1824, n_16855);
  and g43152 (n2636, \asqrt[44] , n_1522, n_1520, n2383);
  and g43153 (n2648, \asqrt[44] , n_1530, n_1531, n2392);
  and g43154 (n_17053, n_6224, n_5923);
  and g43155 (n_17054, n_5905, n_5903);
  and g43156 (n9366, n_5904, n_6225, n_17053, n_17054);
  and g43157 (n22934, \asqrt[3] , n_14849, n22194, n_14848);
  and g43158 (n20761, \asqrt[6] , n_13403, n20049, n_13402);
  and g43159 (n18673, \asqrt[9] , n_12027, n17997, n_12026);
  and g43160 (n16693, \asqrt[12] , n_10723, n16053, n_10722);
  and g43161 (n14821, \asqrt[15] , n_9491, n14217, n_9490);
  and g43162 (n13057, \asqrt[18] , n_8331, n12489, n_8330);
  and g43163 (n11401, \asqrt[21] , n_7243, n10869, n_7242);
  and g43164 (n_17055, n_1664, n_1515);
  and g43165 (n_17056, n_1497, n_1495);
  and g43166 (n2601, n_1496, n_1665, n_17055, n_17056);
  and g43167 (n_17057, n_1352, n_1219);
  and g43168 (n_17058, n_1201, n_1199);
  and g43169 (n2141, n_1200, n_1353, n_17057, n_17058);
  and g43170 (n_16816, n_1363, n_1345);
  and g43171 (n2154, n_1343, \asqrt[47] , n_1344, n_16816);
  and g43172 (n11937, \asqrt[20] , n_7594, n_7595, n11393);
  and g43173 (n13629, \asqrt[17] , n_8706, n_8707, n13049);
  and g43174 (n15429, \asqrt[14] , n_9890, n_9891, n14813);
  and g43175 (n17337, \asqrt[11] , n_11146, n_11147, n16685);
  and g43176 (n19353, \asqrt[8] , n_12474, n_12475, n18665);
  and g43177 (n21470, \asqrt[5] , n_13874, n_13875, n20753);
  and g43178 (n23685, \asqrt[2] , n_15343, n_15344, n22926);
  and g43179 (n_16843, n_1675, n_1657);
  and g43180 (n2614, n_1655, \asqrt[45] , n_1656, n_16843);
  and g43181 (n24539, \asqrt[1] , n_15850, n23677, n_15849);
  and g43182 (n22190, \asqrt[4] , n_14354, n21462, n_14353);
  and g43183 (n20045, \asqrt[7] , n_12931, n19345, n_12930);
  and g43184 (n17993, \asqrt[10] , n_11579, n17329, n_11578);
  and g43185 (n16049, \asqrt[13] , n_10299, n15421, n_10298);
  and g43186 (n14213, \asqrt[16] , n_9091, n13621, n_9090);
  and g43187 (n12485, \asqrt[19] , n_7955, n11929, n_7954);
  and g43188 (n10865, \asqrt[22] , n_6890, n_6888, n10348);
  and g43189 (n_16864, n_6555, n_6537);
  and g43190 (n9855, n_6535, \asqrt[25] , n_6536, n_16864);
  and g43191 (n_17062, n_1504, n_1363);
  and g43192 (n_17063, n_1345, n_1343);
  and g43193 (n2365, n_1344, n_1505, n_17062, n_17063);
  and g43194 (n11389, \asqrt[21] , n_7234, n_7235, n10857);
  and g43195 (n13045, \asqrt[18] , n_8322, n_8323, n12477);
  and g43196 (n14809, \asqrt[15] , n_9482, n_9483, n14205);
  and g43197 (n16681, \asqrt[12] , n_10714, n_10715, n16041);
  and g43198 (n18661, \asqrt[9] , n_12018, n_12019, n17985);
  and g43199 (n20749, \asqrt[6] , n_13394, n_13395, n20037);
  and g43200 (n22922, \asqrt[3] , n_14840, n_14841, n22182);
  and g43201 (n_16828, n_1515, n_1497);
  and g43202 (n2378, n_1495, \asqrt[46] , n_1496, n_16828);
  and g43203 (n_17065, n_6544, n_6235);
  and g43204 (n_17066, n_6217, n_6215);
  and g43205 (n9842, n_6216, n_6545, n_17065, n_17066);
  and g43206 (n23673, \asqrt[2] , n_15336, n22914, n_15335);
  and g43207 (n21458, \asqrt[5] , n_13867, n20741, n_13866);
  and g43208 (n19341, \asqrt[8] , n_12467, n18653, n_12466);
  and g43209 (n17325, \asqrt[11] , n_11139, n16673, n_11138);
  and g43210 (n15417, \asqrt[14] , n_9883, n14801, n_9882);
  and g43211 (n13617, \asqrt[17] , n_8699, n13037, n_8698);
  and g43212 (n11925, \asqrt[20] , n_7587, n11381, n_7586);
  and g43213 (n12473, \asqrt[19] , n_7946, n_7947, n11917);
  and g43214 (n14201, \asqrt[16] , n_9082, n_9083, n13609);
  and g43215 (n16037, \asqrt[13] , n_10290, n_10291, n15409);
  and g43216 (n17981, \asqrt[10] , n_11570, n_11571, n17317);
  and g43217 (n20033, \asqrt[7] , n_12922, n_12923, n19333);
  and g43218 (n22178, \asqrt[4] , n_14345, n_14346, n21450);
  and g43219 (n24166, \asqrt[1] , n_15841, n_15842, n23665);
  and g43220 (n22910, \asqrt[3] , n_14833, n22170, n_14832);
  and g43221 (n20737, \asqrt[6] , n_13387, n20025, n_13386);
  and g43222 (n18649, \asqrt[9] , n_12011, n17973, n_12010);
  and g43223 (n16669, \asqrt[12] , n_10707, n16029, n_10706);
  and g43224 (n14797, \asqrt[15] , n_9475, n14193, n_9474);
  and g43225 (n13033, \asqrt[18] , n_8315, n12465, n_8314);
  and g43226 (n11377, \asqrt[21] , n_7226, n_7224, n10848);
  and g43227 (n_16852, n_6883, n_6865);
  and g43228 (n10343, n_6863, \asqrt[24] , n_6864, n_16852);
  and g43229 (n11913, \asqrt[20] , n_7578, n_7579, n11369);
  and g43230 (n13605, \asqrt[17] , n_8690, n_8691, n13025);
  and g43231 (n15405, \asqrt[14] , n_9874, n_9875, n14789);
  and g43232 (n17313, \asqrt[11] , n_11130, n_11131, n16661);
  and g43233 (n19329, \asqrt[8] , n_12458, n_12459, n18641);
  and g43234 (n21446, \asqrt[5] , n_13858, n_13859, n20729);
  and g43235 (n23661, \asqrt[2] , n_15327, n_15328, n22902);
  and g43236 (n_17068, n_6872, n_6555);
  and g43237 (n_17069, n_6537, n_6535);
  and g43238 (n10330, n_6536, n_6873, n_17068, n_17069);
  and g43239 (n24522, \asqrt[1] , n_15834, n23653, n_15833);
  and g43240 (n22166, \asqrt[4] , n_14338, n21438, n_14337);
  and g43241 (n20021, \asqrt[7] , n_12915, n19321, n_12914);
  and g43242 (n17969, \asqrt[10] , n_11563, n17305, n_11562);
  and g43243 (n16025, \asqrt[13] , n_10283, n15397, n_10282);
  and g43244 (n14189, \asqrt[16] , n_9075, n13597, n_9074);
  and g43245 (n12461, \asqrt[19] , n_7939, n11905, n_7938);
  and g43246 (n13021, \asqrt[18] , n_8306, n_8307, n12453);
  and g43247 (n14785, \asqrt[15] , n_9466, n_9467, n14181);
  and g43248 (n16657, \asqrt[12] , n_10698, n_10699, n16017);
  and g43249 (n18637, \asqrt[9] , n_12002, n_12003, n17961);
  and g43250 (n20725, \asqrt[6] , n_13378, n_13379, n20013);
  and g43251 (n22898, \asqrt[3] , n_14824, n_14825, n22158);
  and g43252 (n23649, \asqrt[2] , n_15320, n22890, n_15319);
  and g43253 (n21434, \asqrt[5] , n_13851, n20717, n_13850);
  and g43254 (n19317, \asqrt[8] , n_12451, n18629, n_12450);
  and g43255 (n17301, \asqrt[11] , n_11123, n16649, n_11122);
  and g43256 (n15393, \asqrt[14] , n_9867, n14777, n_9866);
  and g43257 (n13593, \asqrt[17] , n_8683, n13013, n_8682);
  and g43258 (n11901, \asqrt[20] , n_7570, n_7568, n11360);
  and g43259 (n_16837, n_7219, n_7201);
  and g43260 (n10843, n_7199, \asqrt[23] , n_7200, n_16837);
  and g43261 (n12449, \asqrt[19] , n_7930, n_7931, n11893);
  and g43262 (n14177, \asqrt[16] , n_9066, n_9067, n13585);
  and g43263 (n16013, \asqrt[13] , n_10274, n_10275, n15385);
  and g43264 (n17957, \asqrt[10] , n_11554, n_11555, n17293);
  and g43265 (n20009, \asqrt[7] , n_12906, n_12907, n19309);
  and g43266 (n22154, \asqrt[4] , n_14329, n_14330, n21426);
  and g43267 (n24173, \asqrt[1] , n_15825, n_15826, n23641);
  and g43268 (n_17071, n_7208, n_6883);
  and g43269 (n_17072, n_6865, n_6863);
  and g43270 (n10830, n_6864, n_7209, n_17071, n_17072);
  and g43271 (n22886, \asqrt[3] , n_14817, n22146, n_14816);
  and g43272 (n20713, \asqrt[6] , n_13371, n20001, n_13370);
  and g43273 (n18625, \asqrt[9] , n_11995, n17949, n_11994);
  and g43274 (n16645, \asqrt[12] , n_10691, n16005, n_10690);
  and g43275 (n14773, \asqrt[15] , n_9459, n14169, n_9458);
  and g43276 (n13009, \asqrt[18] , n_8299, n12441, n_8298);
  and g43277 (n13581, \asqrt[17] , n_8674, n_8675, n13001);
  and g43278 (n15381, \asqrt[14] , n_9858, n_9859, n14765);
  and g43279 (n17289, \asqrt[11] , n_11114, n_11115, n16637);
  and g43280 (n19305, \asqrt[8] , n_12442, n_12443, n18617);
  and g43281 (n21422, \asqrt[5] , n_13842, n_13843, n20705);
  and g43282 (n23637, \asqrt[2] , n_15311, n_15312, n22878);
  and g43283 (n24505, \asqrt[1] , n_15818, n23629, n_15817);
  and g43284 (n22142, \asqrt[4] , n_14322, n21414, n_14321);
  and g43285 (n19997, \asqrt[7] , n_12899, n19297, n_12898);
  and g43286 (n17945, \asqrt[10] , n_11547, n17281, n_11546);
  and g43287 (n16001, \asqrt[13] , n_10267, n15373, n_10266);
  and g43288 (n14165, \asqrt[16] , n_9059, n13573, n_9058);
  and g43289 (n12437, \asqrt[19] , n_7922, n_7920, n11884);
  and g43290 (n_16825, n_7563, n_7545);
  and g43291 (n11355, n_7543, \asqrt[22] , n_7544, n_16825);
  and g43292 (n12997, \asqrt[18] , n_8290, n_8291, n12429);
  and g43293 (n14761, \asqrt[15] , n_9450, n_9451, n14157);
  and g43294 (n16633, \asqrt[12] , n_10682, n_10683, n15993);
  and g43295 (n18613, \asqrt[9] , n_11986, n_11987, n17937);
  and g43296 (n20701, \asqrt[6] , n_13362, n_13363, n19989);
  and g43297 (n22874, \asqrt[3] , n_14808, n_14809, n22134);
  and g43298 (n_17074, n_7552, n_7219);
  and g43299 (n_17075, n_7201, n_7199);
  and g43300 (n11342, n_7200, n_7553, n_17074, n_17075);
  and g43301 (n23625, \asqrt[2] , n_15304, n22866, n_15303);
  and g43302 (n21410, \asqrt[5] , n_13835, n20693, n_13834);
  and g43303 (n19293, \asqrt[8] , n_12435, n18605, n_12434);
  and g43304 (n17277, \asqrt[11] , n_11107, n16625, n_11106);
  and g43305 (n15369, \asqrt[14] , n_9851, n14753, n_9850);
  and g43306 (n13569, \asqrt[17] , n_8667, n12989, n_8666);
  and g43307 (n14153, \asqrt[16] , n_9050, n_9051, n13561);
  and g43308 (n15989, \asqrt[13] , n_10258, n_10259, n15361);
  and g43309 (n17933, \asqrt[10] , n_11538, n_11539, n17269);
  and g43310 (n19985, \asqrt[7] , n_12890, n_12891, n19285);
  and g43311 (n22130, \asqrt[4] , n_14313, n_14314, n21402);
  and g43312 (n24180, \asqrt[1] , n_15809, n_15810, n23617);
  and g43313 (n22862, \asqrt[3] , n_14801, n22122, n_14800);
  and g43314 (n20689, \asqrt[6] , n_13355, n19977, n_13354);
  and g43315 (n18601, \asqrt[9] , n_11979, n17925, n_11978);
  and g43316 (n16621, \asqrt[12] , n_10675, n15981, n_10674);
  and g43317 (n14749, \asqrt[15] , n_9443, n14145, n_9442);
  and g43318 (n12985, \asqrt[18] , n_8282, n_8280, n12420);
  and g43319 (n_16813, n_7915, n_7897);
  and g43320 (n11879, n_7895, \asqrt[21] , n_7896, n_16813);
  and g43321 (n13557, \asqrt[17] , n_8658, n_8659, n12977);
  and g43322 (n15357, \asqrt[14] , n_9842, n_9843, n14741);
  and g43323 (n17265, \asqrt[11] , n_11098, n_11099, n16613);
  and g43324 (n19281, \asqrt[8] , n_12426, n_12427, n18593);
  and g43325 (n21398, \asqrt[5] , n_13826, n_13827, n20681);
  and g43326 (n23613, \asqrt[2] , n_15295, n_15296, n22854);
  and g43327 (n_17077, n_7904, n_7563);
  and g43328 (n_17078, n_7545, n_7543);
  and g43329 (n11866, n_7544, n_7905, n_17077, n_17078);
  and g43330 (n24488, \asqrt[1] , n_15802, n23605, n_15801);
  and g43331 (n22118, \asqrt[4] , n_14306, n21390, n_14305);
  and g43332 (n19973, \asqrt[7] , n_12883, n19273, n_12882);
  and g43333 (n17921, \asqrt[10] , n_11531, n17257, n_11530);
  and g43334 (n15977, \asqrt[13] , n_10251, n15349, n_10250);
  and g43335 (n14141, \asqrt[16] , n_9043, n13549, n_9042);
  and g43336 (n14737, \asqrt[15] , n_9434, n_9435, n14133);
  and g43337 (n16609, \asqrt[12] , n_10666, n_10667, n15969);
  and g43338 (n18589, \asqrt[9] , n_11970, n_11971, n17913);
  and g43339 (n20677, \asqrt[6] , n_13346, n_13347, n19965);
  and g43340 (n22850, \asqrt[3] , n_14792, n_14793, n22110);
  and g43341 (n23601, \asqrt[2] , n_15288, n22842, n_15287);
  and g43342 (n21386, \asqrt[5] , n_13819, n20669, n_13818);
  and g43343 (n19269, \asqrt[8] , n_12419, n18581, n_12418);
  and g43344 (n17253, \asqrt[11] , n_11091, n16601, n_11090);
  and g43345 (n15345, \asqrt[14] , n_9835, n14729, n_9834);
  and g43346 (n13545, \asqrt[17] , n_8650, n_8648, n12968);
  and g43347 (n_16797, n_8275, n_8257);
  and g43348 (n12415, n_8255, \asqrt[20] , n_8256, n_16797);
  and g43349 (n14129, \asqrt[16] , n_9034, n_9035, n13537);
  and g43350 (n15965, \asqrt[13] , n_10242, n_10243, n15337);
  and g43351 (n17909, \asqrt[10] , n_11522, n_11523, n17245);
  and g43352 (n19961, \asqrt[7] , n_12874, n_12875, n19261);
  and g43353 (n22106, \asqrt[4] , n_14297, n_14298, n21378);
  and g43354 (n24187, \asqrt[1] , n_15793, n_15794, n23593);
  and g43355 (n_17080, n_8264, n_7915);
  and g43356 (n_17081, n_7897, n_7895);
  and g43357 (n12402, n_7896, n_8265, n_17080, n_17081);
  and g43358 (n22838, \asqrt[3] , n_14785, n22098, n_14784);
  and g43359 (n20665, \asqrt[6] , n_13339, n19953, n_13338);
  and g43360 (n18577, \asqrt[9] , n_11963, n17901, n_11962);
  and g43361 (n16597, \asqrt[12] , n_10659, n15957, n_10658);
  and g43362 (n14725, \asqrt[15] , n_9427, n14121, n_9426);
  and g43363 (n15333, \asqrt[14] , n_9826, n_9827, n14717);
  and g43364 (n17241, \asqrt[11] , n_11082, n_11083, n16589);
  and g43365 (n19257, \asqrt[8] , n_12410, n_12411, n18569);
  and g43366 (n21374, \asqrt[5] , n_13810, n_13811, n20657);
  and g43367 (n23589, \asqrt[2] , n_15279, n_15280, n22830);
  and g43368 (n24471, \asqrt[1] , n_15786, n23581, n_15785);
  and g43369 (n22094, \asqrt[4] , n_14290, n21366, n_14289);
  and g43370 (n19949, \asqrt[7] , n_12867, n19249, n_12866);
  and g43371 (n17897, \asqrt[10] , n_11515, n17233, n_11514);
  and g43372 (n15953, \asqrt[13] , n_10235, n15325, n_10234);
  and g43373 (n14117, \asqrt[16] , n_9026, n_9024, n13528);
  and g43374 (n_16785, n_8643, n_8625);
  and g43375 (n12963, n_8623, \asqrt[19] , n_8624, n_16785);
  and g43376 (n14713, \asqrt[15] , n_9418, n_9419, n14109);
  and g43377 (n16585, \asqrt[12] , n_10650, n_10651, n15945);
  and g43378 (n18565, \asqrt[9] , n_11954, n_11955, n17889);
  and g43379 (n20653, \asqrt[6] , n_13330, n_13331, n19941);
  and g43380 (n22826, \asqrt[3] , n_14776, n_14777, n22086);
  and g43381 (n_17083, n_8632, n_8275);
  and g43382 (n_17084, n_8257, n_8255);
  and g43383 (n12950, n_8256, n_8633, n_17083, n_17084);
  and g43384 (n23577, \asqrt[2] , n_15272, n22818, n_15271);
  and g43385 (n21362, \asqrt[5] , n_13803, n20645, n_13802);
  and g43386 (n19245, \asqrt[8] , n_12403, n18557, n_12402);
  and g43387 (n17229, \asqrt[11] , n_11075, n16577, n_11074);
  and g43388 (n15321, \asqrt[14] , n_9819, n14705, n_9818);
  and g43389 (n15941, \asqrt[13] , n_10226, n_10227, n15313);
  and g43390 (n17885, \asqrt[10] , n_11506, n_11507, n17221);
  and g43391 (n19937, \asqrt[7] , n_12858, n_12859, n19237);
  and g43392 (n22082, \asqrt[4] , n_14281, n_14282, n21354);
  and g43393 (n24194, \asqrt[1] , n_15777, n_15778, n23569);
  and g43394 (n22814, \asqrt[3] , n_14769, n22074, n_14768);
  and g43395 (n20641, \asqrt[6] , n_13323, n19929, n_13322);
  and g43396 (n18553, \asqrt[9] , n_11947, n17877, n_11946);
  and g43397 (n16573, \asqrt[12] , n_10643, n15933, n_10642);
  and g43398 (n14701, \asqrt[15] , n_9410, n_9408, n14100);
  and g43399 (n_16770, n_9019, n_9001);
  and g43400 (n13523, n_8999, \asqrt[18] , n_9000, n_16770);
  and g43401 (n15309, \asqrt[14] , n_9810, n_9811, n14693);
  and g43402 (n17217, \asqrt[11] , n_11066, n_11067, n16565);
  and g43403 (n19233, \asqrt[8] , n_12394, n_12395, n18545);
  and g43404 (n21350, \asqrt[5] , n_13794, n_13795, n20633);
  and g43405 (n23565, \asqrt[2] , n_15263, n_15264, n22806);
  and g43406 (n_17086, n_9008, n_8643);
  and g43407 (n_17087, n_8625, n_8623);
  and g43408 (n13510, n_8624, n_9009, n_17086, n_17087);
  and g43409 (n24454, \asqrt[1] , n_15770, n23557, n_15769);
  and g43410 (n22070, \asqrt[4] , n_14274, n21342, n_14273);
  and g43411 (n19925, \asqrt[7] , n_12851, n19225, n_12850);
  and g43412 (n17873, \asqrt[10] , n_11499, n17209, n_11498);
  and g43413 (n15929, \asqrt[13] , n_10219, n15301, n_10218);
  and g43414 (n16561, \asqrt[12] , n_10634, n_10635, n15921);
  and g43415 (n18541, \asqrt[9] , n_11938, n_11939, n17865);
  and g43416 (n20629, \asqrt[6] , n_13314, n_13315, n19917);
  and g43417 (n22802, \asqrt[3] , n_14760, n_14761, n22062);
  and g43418 (n23553, \asqrt[2] , n_15256, n22794, n_15255);
  and g43419 (n21338, \asqrt[5] , n_13787, n20621, n_13786);
  and g43420 (n19221, \asqrt[8] , n_12387, n18533, n_12386);
  and g43421 (n17205, \asqrt[11] , n_11059, n16553, n_11058);
  and g43422 (n15297, \asqrt[14] , n_9802, n_9800, n14684);
  and g43423 (n_16758, n_9403, n_9385);
  and g43424 (n14095, n_9383, \asqrt[17] , n_9384, n_16758);
  and g43425 (n15917, \asqrt[13] , n_10210, n_10211, n15289);
  and g43426 (n17861, \asqrt[10] , n_11490, n_11491, n17197);
  and g43427 (n19913, \asqrt[7] , n_12842, n_12843, n19213);
  and g43428 (n22058, \asqrt[4] , n_14265, n_14266, n21330);
  and g43429 (n24201, \asqrt[1] , n_15761, n_15762, n23545);
  and g43430 (n_17089, n_9392, n_9019);
  and g43431 (n_17090, n_9001, n_8999);
  and g43432 (n14082, n_9000, n_9393, n_17089, n_17090);
  and g43433 (n22790, \asqrt[3] , n_14753, n22050, n_14752);
  and g43434 (n20617, \asqrt[6] , n_13307, n19905, n_13306);
  and g43435 (n18529, \asqrt[9] , n_11931, n17853, n_11930);
  and g43436 (n16549, \asqrt[12] , n_10627, n15909, n_10626);
  and g43437 (n17193, \asqrt[11] , n_11050, n_11051, n16541);
  and g43438 (n19209, \asqrt[8] , n_12378, n_12379, n18521);
  and g43439 (n21326, \asqrt[5] , n_13778, n_13779, n20609);
  and g43440 (n23541, \asqrt[2] , n_15247, n_15248, n22782);
  and g43441 (n24437, \asqrt[1] , n_15754, n23533, n_15753);
  and g43442 (n22046, \asqrt[4] , n_14258, n21318, n_14257);
  and g43443 (n19901, \asqrt[7] , n_12835, n19201, n_12834);
  and g43444 (n17849, \asqrt[10] , n_11483, n17185, n_11482);
  and g43445 (n15905, \asqrt[13] , n_10202, n_10200, n15280);
  and g43446 (n_16746, n_9795, n_9777);
  and g43447 (n14679, n_9775, \asqrt[16] , n_9776, n_16746);
  and g43448 (n16537, \asqrt[12] , n_10618, n_10619, n15897);
  and g43449 (n18517, \asqrt[9] , n_11922, n_11923, n17841);
  and g43450 (n20605, \asqrt[6] , n_13298, n_13299, n19893);
  and g43451 (n22778, \asqrt[3] , n_14744, n_14745, n22038);
  and g43452 (n_17092, n_9784, n_9403);
  and g43453 (n_17093, n_9385, n_9383);
  and g43454 (n14666, n_9384, n_9785, n_17092, n_17093);
  and g43455 (n23529, \asqrt[2] , n_15240, n22770, n_15239);
  and g43456 (n21314, \asqrt[5] , n_13771, n20597, n_13770);
  and g43457 (n19197, \asqrt[8] , n_12371, n18509, n_12370);
  and g43458 (n17181, \asqrt[11] , n_11043, n16529, n_11042);
  and g43459 (n17837, \asqrt[10] , n_11474, n_11475, n17173);
  and g43460 (n19889, \asqrt[7] , n_12826, n_12827, n19189);
  and g43461 (n22034, \asqrt[4] , n_14249, n_14250, n21306);
  and g43462 (n24208, \asqrt[1] , n_15745, n_15746, n23521);
  and g43463 (n22766, \asqrt[3] , n_14737, n22026, n_14736);
  and g43464 (n20593, \asqrt[6] , n_13291, n19881, n_13290);
  and g43465 (n18505, \asqrt[9] , n_11915, n17829, n_11914);
  and g43466 (n16525, \asqrt[12] , n_10610, n_10608, n15888);
  and g43467 (n_16731, n_10195, n_10177);
  and g43468 (n15275, n_10175, \asqrt[15] , n_10176, n_16731);
  and g43469 (n17169, \asqrt[11] , n_11034, n_11035, n16517);
  and g43470 (n19185, \asqrt[8] , n_12362, n_12363, n18497);
  and g43471 (n21302, \asqrt[5] , n_13762, n_13763, n20585);
  and g43472 (n23517, \asqrt[2] , n_15231, n_15232, n22758);
  and g43473 (n_17095, n_10184, n_9795);
  and g43474 (n_17096, n_9777, n_9775);
  and g43475 (n15262, n_9776, n_10185, n_17095, n_17096);
  and g43476 (n24420, \asqrt[1] , n_15738, n23509, n_15737);
  and g43477 (n22022, \asqrt[4] , n_14242, n21294, n_14241);
  and g43478 (n19877, \asqrt[7] , n_12819, n19177, n_12818);
  and g43479 (n17825, \asqrt[10] , n_11467, n17161, n_11466);
  and g43480 (n18493, \asqrt[9] , n_11906, n_11907, n17817);
  and g43481 (n20581, \asqrt[6] , n_13282, n_13283, n19869);
  and g43482 (n22754, \asqrt[3] , n_14728, n_14729, n22014);
  and g43483 (n23505, \asqrt[2] , n_15224, n22746, n_15223);
  and g43484 (n21290, \asqrt[5] , n_13755, n20573, n_13754);
  and g43485 (n19173, \asqrt[8] , n_12355, n18485, n_12354);
  and g43486 (n17157, \asqrt[11] , n_11026, n_11024, n16508);
  and g43487 (n_16719, n_10603, n_10585);
  and g43488 (n15883, n_10583, \asqrt[14] , n_10584, n_16719);
  and g43489 (n17813, \asqrt[10] , n_11458, n_11459, n17149);
  and g43490 (n19865, \asqrt[7] , n_12810, n_12811, n19165);
  and g43491 (n22010, \asqrt[4] , n_14233, n_14234, n21282);
  and g43492 (n24215, \asqrt[1] , n_15729, n_15730, n23497);
  and g43493 (n_17098, n_10592, n_10195);
  and g43494 (n_17099, n_10177, n_10175);
  and g43495 (n15870, n_10176, n_10593, n_17098, n_17099);
  and g43496 (n22742, \asqrt[3] , n_14721, n22002, n_14720);
  and g43497 (n20569, \asqrt[6] , n_13275, n19857, n_13274);
  and g43498 (n18481, \asqrt[9] , n_11899, n17805, n_11898);
  and g43499 (n19161, \asqrt[8] , n_12346, n_12347, n18473);
  and g43500 (n21278, \asqrt[5] , n_13746, n_13747, n20561);
  and g43501 (n23493, \asqrt[2] , n_15215, n_15216, n22734);
  and g43502 (n24403, \asqrt[1] , n_15722, n23485, n_15721);
  and g43503 (n21998, \asqrt[4] , n_14226, n21270, n_14225);
  and g43504 (n19853, \asqrt[7] , n_12803, n19153, n_12802);
  and g43505 (n17801, \asqrt[10] , n_11450, n_11448, n17140);
  and g43506 (n_16707, n_11019, n_11001);
  and g43507 (n16503, n_10999, \asqrt[13] , n_11000, n_16707);
  and g43508 (n18469, \asqrt[9] , n_11890, n_11891, n17793);
  and g43509 (n20557, \asqrt[6] , n_13266, n_13267, n19845);
  and g43510 (n22730, \asqrt[3] , n_14712, n_14713, n21990);
  and g43511 (n_17101, n_11008, n_10603);
  and g43512 (n_17102, n_10585, n_10583);
  and g43513 (n16490, n_10584, n_11009, n_17101, n_17102);
  and g43514 (n23481, \asqrt[2] , n_15208, n22722, n_15207);
  and g43515 (n21266, \asqrt[5] , n_13739, n20549, n_13738);
  and g43516 (n19149, \asqrt[8] , n_12339, n18461, n_12338);
  and g43517 (n19841, \asqrt[7] , n_12794, n_12795, n19141);
  and g43518 (n21986, \asqrt[4] , n_14217, n_14218, n21258);
  and g43519 (n24222, \asqrt[1] , n_15713, n_15714, n23473);
  and g43520 (n22718, \asqrt[3] , n_14705, n21978, n_14704);
  and g43521 (n20545, \asqrt[6] , n_13259, n19833, n_13258);
  and g43522 (n18457, \asqrt[9] , n_11882, n_11880, n17784);
  and g43523 (n_16692, n_11443, n_11425);
  and g43524 (n17135, n_11423, \asqrt[12] , n_11424, n_16692);
  and g43525 (n19137, \asqrt[8] , n_12330, n_12331, n18449);
  and g43526 (n21254, \asqrt[5] , n_13730, n_13731, n20537);
  and g43527 (n23469, \asqrt[2] , n_15199, n_15200, n22710);
  and g43528 (n_17104, n_11432, n_11019);
  and g43529 (n_17105, n_11001, n_10999);
  and g43530 (n17122, n_11000, n_11433, n_17104, n_17105);
  and g43531 (n24386, \asqrt[1] , n_15706, n23461, n_15705);
  and g43532 (n21974, \asqrt[4] , n_14210, n21246, n_14209);
  and g43533 (n19829, \asqrt[7] , n_12787, n19129, n_12786);
  and g43534 (n20533, \asqrt[6] , n_13250, n_13251, n19821);
  and g43535 (n22706, \asqrt[3] , n_14696, n_14697, n21966);
  and g43536 (n23457, \asqrt[2] , n_15192, n22698, n_15191);
  and g43537 (n21242, \asqrt[5] , n_13723, n20525, n_13722);
  and g43538 (n19125, \asqrt[8] , n_12322, n_12320, n18440);
  and g43539 (n_16680, n_11875, n_11857);
  and g43540 (n17779, n_11855, \asqrt[11] , n_11856, n_16680);
  and g43541 (n19817, \asqrt[7] , n_12778, n_12779, n19117);
  and g43542 (n21962, \asqrt[4] , n_14201, n_14202, n21234);
  and g43543 (n24229, \asqrt[1] , n_15697, n_15698, n23449);
  and g43544 (n_17107, n_11864, n_11443);
  and g43545 (n_17108, n_11425, n_11423);
  and g43546 (n17766, n_11424, n_11865, n_17107, n_17108);
  and g43547 (n22694, \asqrt[3] , n_14689, n21954, n_14688);
  and g43548 (n20521, \asqrt[6] , n_13243, n19809, n_13242);
  and g43549 (n21230, \asqrt[5] , n_13714, n_13715, n20513);
  and g43550 (n23445, \asqrt[2] , n_15183, n_15184, n22686);
  and g43551 (n24369, \asqrt[1] , n_15690, n23437, n_15689);
  and g43552 (n21950, \asqrt[4] , n_14194, n21222, n_14193);
  and g43553 (n19805, \asqrt[7] , n_12770, n_12768, n19108);
  and g43554 (n_16665, n_12315, n_12297);
  and g43555 (n18435, n_12295, \asqrt[10] , n_12296, n_16665);
  and g43556 (n20509, \asqrt[6] , n_13234, n_13235, n19797);
  and g43557 (n22682, \asqrt[3] , n_14680, n_14681, n21942);
  and g43558 (n_17110, n_12304, n_11875);
  and g43559 (n_17111, n_11857, n_11855);
  and g43560 (n18422, n_11856, n_12305, n_17110, n_17111);
  and g43561 (n23433, \asqrt[2] , n_15176, n22674, n_15175);
  and g43562 (n21218, \asqrt[5] , n_13707, n20501, n_13706);
  and g43563 (n21938, \asqrt[4] , n_14185, n_14186, n21210);
  and g43564 (n24236, \asqrt[1] , n_15681, n_15682, n23425);
  and g43565 (n22670, \asqrt[3] , n_14673, n21930, n_14672);
  and g43566 (n20497, \asqrt[6] , n_13226, n_13224, n19788);
  and g43567 (n_16653, n_12763, n_12745);
  and g43568 (n19103, n_12743, \asqrt[9] , n_12744, n_16653);
  and g43569 (n21206, \asqrt[5] , n_13698, n_13699, n20489);
  and g43570 (n23421, \asqrt[2] , n_15167, n_15168, n22662);
  and g43571 (n_17113, n_12752, n_12315);
  and g43572 (n_17114, n_12297, n_12295);
  and g43573 (n19090, n_12296, n_12753, n_17113, n_17114);
  and g43574 (n24352, \asqrt[1] , n_15674, n23413, n_15673);
  and g43575 (n21926, \asqrt[4] , n_14178, n21198, n_14177);
  and g43576 (n22658, \asqrt[3] , n_14664, n_14665, n21918);
  and g43577 (n23409, \asqrt[2] , n_15160, n22650, n_15159);
  and g43578 (n21194, \asqrt[5] , n_13690, n_13688, n20480);
  and g43579 (n_16645, n_13219, n_13201);
  and g43580 (n19783, n_13199, \asqrt[8] , n_13200, n_16645);
  and g43581 (n21914, \asqrt[4] , n_14169, n_14170, n21186);
  and g43582 (n24243, \asqrt[1] , n_15665, n_15666, n23401);
  and g43583 (n_17116, n_13208, n_12763);
  and g43584 (n_17117, n_12745, n_12743);
  and g43585 (n19770, n_12744, n_13209, n_17116, n_17117);
  and g43586 (n22646, \asqrt[3] , n_14657, n21906, n_14656);
  and g43587 (n23397, \asqrt[2] , n_15151, n_15152, n22638);
  and g43588 (n24335, \asqrt[1] , n_15658, n23389, n_15657);
  and g43589 (n21902, \asqrt[4] , n_14161, n_14159, n21177);
  and g43590 (n_17118, n_13683, n_13665);
  and g43591 (n20475, n_13663, \asqrt[7] , n_13664, n_17118);
  and g43592 (n22634, \asqrt[3] , n_14648, n_14649, n21894);
  and g43593 (n_17119, n_13672, n_13219);
  and g43594 (n_17120, n_13201, n_13199);
  and g43595 (n20462, n_13200, n_13673, n_17119, n_17120);
  and g43596 (n23385, \asqrt[2] , n_15144, n22626, n_15143);
  and g43597 (n24250, \asqrt[1] , n_15649, n_15650, n23377);
  and g43598 (n22622, \asqrt[3] , n_14640, n_14638, n21885);
  and g43599 (n21172, n_14154, n_14135, \asqrt[6] , n_14136);
  and g43600 (n23373, \asqrt[2] , n_15135, n_15136, n22614);
  and g43601 (n_17121, n_14143, n_13683);
  and g43602 (n_17122, n_13665, n_13663);
  and g43603 (n21160, n_13664, n_14144, n_17121, n_17122);
  and g43604 (n24318, \asqrt[1] , n_15642, n23365, n_15641);
  and g43605 (n23361, \asqrt[2] , n_15127, n_15125, n22605);
  and g43606 (n21880, n_14633, n_14614, \asqrt[5] , n_14615);
  and g43607 (n24254, \asqrt[1] , n_15633, n_15634, n23353);
  and g43608 (n_17123, n_14622, n_14154);
  and g43609 (n21868, n_14135, n_14136, n_14623, n_17123);
  and g43610 (n24301, \asqrt[1] , n_15625, n_15623, n23344);
  and g43611 (n22600, n_15120, n_15101, \asqrt[4] , n_15102);
  and g43612 (n_17124, n_15109, n_14633);
  and g43613 (n22588, n_14614, n_14615, n_15110, n_17124);
  and g43614 (n23339, n_17125, n_15596, \asqrt[3] , n_15597);
  not g43615 (n_17125, n23303);
  and g43616 (n_17126, n_15607, n_15120);
  and g43617 (n23327, n_15101, n_15102, n_15608, n_17126);
  and g43618 (n24268, n_16194, n_16099, \asqrt[2] , n_16100);
  and g43619 (n24280, n_16194, n_16099, \a[2] , n_16100);
endmodule

