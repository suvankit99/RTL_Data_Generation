
module c2670(N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19,
     N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34,
     N35, N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53,
     N54, N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68,
     N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85,
     N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100,
     N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, N113,
     N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126,
     N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139,
     N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241,
     N246, N253, N256, N259, N262, N263, N266, N269, N272, N275, N278,
     N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, N316,
     N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349,
     N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I,
     N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I,
     N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I,
     N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I,
     N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I,
     N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I,
     N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I,
     N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I,
     N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I,
     N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, N401,
     N419, N420, N456, N457, N458, N487, N488, N489, N490, N491, N492,
     N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, N1277,
     N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969,
     N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022,
     N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925,
     N2970, N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809,
     N3851, N3875, N3881, N3882, N143_O, N144_O, N145_O, N146_O,
     N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, N154_O,
     N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O,
     N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O,
     N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O,
     N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O,
     N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O,
     N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O,
     N203_O, N204_O, N205_O, N206_O, N207_O, N208_O, N209_O, N210_O,
     N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, N217_O, N218_O);
  input N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20,
       N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35,
       N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54,
       N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
       N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86,
       N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100,
       N101, N102, N103, N104, N105, N106, N107, N108, N111, N112,
       N113, N114, N115, N116, N117, N118, N119, N120, N123, N124,
       N125, N126, N127, N128, N129, N130, N131, N132, N135, N136,
       N137, N138, N139, N140, N141, N142, N219, N224, N227, N230,
       N231, N234, N237, N241, N246, N253, N256, N259, N262, N263,
       N266, N269, N272, N275, N278, N281, N284, N287, N290, N294,
       N297, N301, N305, N309, N313, N316, N319, N322, N325, N328,
       N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I,
       N144_I, N145_I, N146_I, N147_I, N148_I, N149_I, N150_I, N151_I,
       N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, N159_I,
       N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I,
       N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I,
       N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I,
       N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, N190_I, N191_I,
       N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, N199_I,
       N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I,
       N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I,
       N216_I, N217_I, N218_I;
  output N398, N400, N401, N419, N420, N456, N457, N458, N487, N488,
       N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026,
       N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818,
       N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014,
       N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496,
       N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546,
       N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O,
       N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O,
       N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O,
       N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O,
       N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O,
       N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O,
       N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, N190_O, N191_O,
       N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O,
       N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O,
       N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O,
       N216_O, N217_O, N218_O;
  wire N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20,
       N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35,
       N36, N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54,
       N55, N56, N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
       N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N85, N86,
       N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N99, N100,
       N101, N102, N103, N104, N105, N106, N107, N108, N111, N112,
       N113, N114, N115, N116, N117, N118, N119, N120, N123, N124,
       N125, N126, N127, N128, N129, N130, N131, N132, N135, N136,
       N137, N138, N139, N140, N141, N142, N219, N224, N227, N230,
       N231, N234, N237, N241, N246, N253, N256, N259, N262, N263,
       N266, N269, N272, N275, N278, N281, N284, N287, N290, N294,
       N297, N301, N305, N309, N313, N316, N319, N322, N325, N328,
       N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I,
       N144_I, N145_I, N146_I, N147_I, N148_I, N149_I, N150_I, N151_I,
       N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, N159_I,
       N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I,
       N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I,
       N176_I, N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I,
       N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, N190_I, N191_I,
       N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, N199_I,
       N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I,
       N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I,
       N216_I, N217_I, N218_I;
  wire N398, N400, N401, N419, N420, N456, N457, N458, N487, N488,
       N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026,
       N1028, N1029, N1269, N1277, N1448, N1726, N1816, N1817, N1818,
       N1819, N1820, N1821, N1969, N1970, N1971, N2010, N2012, N2014,
       N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, N2496,
       N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546,
       N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O,
       N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O,
       N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O,
       N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O,
       N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O,
       N176_O, N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O,
       N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, N190_O, N191_O,
       N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, N199_O,
       N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O,
       N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O,
       N216_O, N217_O, N218_O;
  wire N405, N408, N425, N485, N486, N495, N533, N537;
  wire N543, N544, N547, N574, N578, N606, N607, N608;
  wire N609, N610, N611, N612, N650, N651, N655, N659;
  wire N663, N667, N671, N675, N679, N683, N687, N705;
  wire N711, N715, N719, N723, N727, N730, N733, N734;
  wire N800, N900, N901, N902, N903, N904, N905, N998;
  wire N999, N1027, N1032, N1033, N1042, N1053, N1064, N1065;
  wire N1066, N1067, N1068, N1069, N1097, N1098, N1099, N1100;
  wire N1101, N1102, N1113, N1124, N1125, N1126, N1127, N1128;
  wire N1129, N1133, N1137, N1141, N1168, N1169, N1170, N1171;
  wire N1172, N1173, N1185, N1200, N1216, N1275, N1276, N1302;
  wire N1351, N1352, N1353, N1354, N1355, N1395, N1396, N1397;
  wire N1398, N1399, N1422, N1423, N1424, N1425, N1426, N1427;
  wire N1440, N1441, N1449, N1450, N1451, N1452, N1453, N1454;
  wire N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462;
  wire N1463, N1464, N1465, N1466, N1467, N1468, N1469, N1470;
  wire N1471, N1472, N1473, N1474, N1475, N1476, N1477, N1478;
  wire N1479, N1480, N1481, N1482, N1483, N1484, N1485, N1486;
  wire N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494;
  wire N1495, N1496, N1499, N1502, N1506, N1510, N1529, N1530;
  wire N1531, N1532, N1533, N1534, N1535, N1536, N1537, N1538;
  wire N1539, N1540, N1541, N1542, N1543, N1544, N1545, N1546;
  wire N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1557;
  wire N1561, N1564, N1565, N1566, N1567, N1568, N1569, N1570;
  wire N1571, N1578, N1581, N1582, N1585, N1588, N1596, N1600;
  wire N1606, N1637, N1642, N1647, N1651, N1656, N1676, N1681;
  wire N1686, N1690, N1708, N1770, N1773, N1776, N1784, N1785;
  wire N1795, N1798, N1807, N1808, N1809, N1810, N1811, N1813;
  wire N1814, N1815, N1822, N1823, N1827, N1830, N1831, N1832;
  wire N1833, N1836, N1885, N1888, N1894, N1908, N1909, N1910;
  wire N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918;
  wire N1919, N1928, N1929, N1930, N1931, N1932, N1933, N1934;
  wire N1935, N1939, N1940, N1941, N2028, N2030, N2031, N2032;
  wire N2033, N2034, N2040, N2042, N2043, N2046, N2049, N2052;
  wire N2055, N2058, N2061, N2064, N2067, N2070, N2073, N2076;
  wire N2079, N2095, N2098, N2101, N2104, N2107, N2110, N2113;
  wire N2119, N2120, N2125, N2126, N2127, N2128, N2144, N2147;
  wire N2150, N2153, N2154, N2155, N2156, N2157, N2158, N2171;
  wire N2172, N2173, N2174, N2176, N2177, N2178, N2219, N2236;
  wire N2237, N2250, N2291, N2294, N2297, N2298, N2300, N2301;
  wire N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309;
  wire N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317;
  wire N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325;
  wire N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333;
  wire N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2354;
  wire N2355, N2356, N2357, N2358, N2359, N2386, N2400, N2406;
  wire N2407, N2408, N2409, N2410, N2411, N2412, N2413, N2414;
  wire N2415, N2416, N2417, N2421, N2425, N2428, N2429, N2430;
  wire N2431, N2432, N2433, N2453, N2469, N2484, N2487, N2490;
  wire N2493, N2503, N2504, N2528, N2531, N2534, N2579, N2607;
  wire N2608, N2609, N2610, N2611, N2612, N2613, N2618, N2619;
  wire N2652, N2663, N2664, N2681, N2684, N2693, N2694, N2703;
  wire N2707, N2708, N2719, N2720, N2743, N2747, N2760, N2771;
  wire N2772, N2773, N2774, N2781, N2782, N2789, N2790, N2791;
  wire N2792, N2793, N2796, N2800, N2826, N2837, N2839, N2840;
  wire N2841, N2874, N2877, N2880, N2881, N2888, N2894, N2895;
  wire N2896, N2897, N2898, N2899, N2900, N2901, N2938, N2939;
  wire N2963, N2972, N2975, N2978, N2981, N2984, N2985, N2986;
  wire N2989, N2992, N3007, N3028, N3035, N3036, N3037, N3047;
  wire N3048, N3049, N3053, N3054, N3055, N3056, N3057, N3058;
  wire N3059, N3060, N3072, N3073, N3076, N3088, N3091, N3137;
  wire N3140, N3143, N3146, N3149, N3152, N3175, N3176, N3180;
  wire N3187, N3191, N3192, N3193, N3194, N3195, N3196, N3197;
  wire N3215, N3216, N3217, N3222, N3223, N3238, N3281, N3282;
  wire N3283, N3284, N3286, N3288, N3289, N3291, N3293, N3296;
  wire N3299, N3301, N3315, N3318, N3321, N3333, N3334, N3335;
  wire N3400, N3401, N3402, N3403, N3404, N3405, N3410, N3450;
  wire N3453, N3478, N3479, N3480, N3481, N3482, N3483, N3484;
  wire N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492;
  wire N3493, N3522, N3525, N3551, N3552, N3553, N3554, N3555;
  wire N3556, N3557, N3559, N3592, N3593, N3594, N3595, N3596;
  wire N3597, N3598, N3599, N3603, N3608, N3612, N3615, N3616;
  wire N3622, N3629, N3630, N3667, N3668, N3669, N3670, N3691;
  wire N3692, N3693, N3694, N3695, N3721, N3722, N3723, N3726;
  wire N3727, N3728, N3729, N3730, N3731, N3732, N3733, N3734;
  wire N3735, N3736, N3750, N3753, N3754, N3758, N3761, N3762;
  wire N3778, N3779, N3802, N3805, N3807, N3808, N3817, N3818;
  wire N3819, N3823, N3826, N3834, N3835, N3838, N3876, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399;
  assign N218_O = N218_I;
  assign N217_O = N217_I;
  assign N216_O = N216_I;
  assign N215_O = N215_I;
//   assign N214_O = N214_I;
  assign N213_O = N213_I;
  assign N212_O = N212_I;
  assign N211_O = N211_I;
  assign N210_O = N210_I;
  assign N209_O = N209_I;
  assign N208_O = N208_I;
  assign N207_O = N207_I;
  assign N206_O = N206_I;
  assign N205_O = N205_I;
//   assign N204_O = N204_I;
  assign N203_O = N203_I;
  assign N202_O = N202_I;
  assign N201_O = N201_I;
  assign N200_O = N200_I;
  assign N199_O = N199_I;
  assign N198_O = N198_I;
  assign N197_O = N197_I;
  assign N196_O = N196_I;
//   assign N195_O = N195_I;
  assign N194_O = N194_I;
  assign N193_O = N193_I;
  assign N192_O = N192_I;
  assign N191_O = N191_I;
  assign N190_O = N190_I;
  assign N189_O = N189_I;
  assign N188_O = N188_I;
  assign N187_O = N187_I;
  assign N186_O = N186_I;
  assign N185_O = N185_I;
  assign N184_O = N184_I;
  assign N183_O = N183_I;
  assign N182_O = N182_I;
  assign N181_O = N181_I;
  assign N180_O = N180_I;
  assign N179_O = N179_I;
  assign N178_O = N178_I;
  assign N177_O = N177_I;
  assign N176_O = N176_I;
  assign N175_O = N175_I;
  assign N174_O = N174_I;
  assign N173_O = N173_I;
  assign N172_O = N172_I;
  assign N171_O = N171_I;
  assign N170_O = N170_I;
//   assign N169_O = N169_I;
  assign N168_O = N168_I;
//   assign N167_O = N167_I;
  assign N166_O = N166_I;
  assign N165_O = N165_I;
  assign N164_O = N164_I;
  assign N163_O = N163_I;
  assign N162_O = N162_I;
  assign N161_O = N161_I;
  assign N160_O = N160_I;
  assign N159_O = N159_I;
  assign N158_O = N158_I;
  assign N157_O = N157_I;
//   assign N156_O = N156_I;
  assign N155_O = N155_I;
  assign N154_O = N154_I;
  assign N153_O = N153_I;
  assign N152_O = N152_I;
//   assign N151_O = N151_I;
  assign N150_O = N150_I;
  assign N149_O = N149_I;
  assign N148_O = N148_I;
  assign N147_O = N147_I;
//   assign N146_O = N146_I;
  assign N145_O = N145_I;
  assign N144_O = N144_I;
  assign N143_O = N143_I;
//   assign N3875 = 1'b0;
//   assign N3804 = N3803;
  assign N2644 = N2643;
  assign N2390 = N2389;
  assign N2388 = N2387;
  assign N805 = N219;
  assign N458 = N290;
  assign N457 = N290;
  assign N456 = N290;
  assign N420 = N253;
  assign N419 = N253;
  assign N401 = N219;
  assign N400 = N219;
  assign N398 = N219;
  and AND2_4 (N405, N1, N3);
  and AND2_32 (N543, N11, N246);
  and AND2_53 (N651, N7, N237);
  and AND2_104 (N1026, N94, N219);
  and AND2_105 (N1027, N325, N651);
  and AND2_110 (N1277, N547, N544);
  and AND2_119 (N1069, N11, N537);
  and AND2_134 (N1128, N319, N322);
  and AND2_189 (N1275, N325, N1032);
  and AND2_190 (N1276, N231, N1033);
  and AND2_237 (N1474, N1042, N234);
  and AND2_256 (N1493, N1102, N1113);
  and AND2_257 (N1494, N319, N1113);
  and AND2_258 (N1495, N1102, N322);
  and AND2_291 (N1544, N19, N1173);
  and AND2_292 (N1545, N4, N1173);
  and AND2_293 (N1546, N20, N1173);
  and AND2_294 (N1547, N5, N1173);
  and AND2_295 (N1548, N21, N1173);
  and AND2_296 (N1549, N22, N1173);
  and AND2_297 (N1550, N23, N1173);
  and AND2_298 (N1551, N6, N1173);
  and AND2_299 (N1552, N24, N1173);
  and AND2_303 (N1564, N25, N1200);
  and AND2_304 (N1565, N32, N1200);
  and AND2_305 (N1566, N26, N1200);
  and AND2_306 (N1567, N33, N1200);
  and AND2_307 (N1568, N27, N1200);
  and AND2_308 (N1569, N34, N1200);
  and AND2_309 (N1570, N35, N1200);
  and AND2_310 (N1571, N28, N1200);
  and AND2_322 (N1726, N1449, N1450);
  and AND2_361 (N1813, N1596, N241);
  and AND2_362 (N1814, N1606, N241);
  and AND2_363 (N1815, N1600, N241);
  and AND2_374 (N1830, N1600, N537);
  and AND2_375 (N1831, N1606, N537);
  and AND2_376 (N1832, N2014, N246);
  and AND2_390 (N1894, N1637, N425);
  and AND2_394 (N1910, N1600, N16);
  and AND2_395 (N1911, N1606, N16);
  and AND2_396 (N1912, N2010, N16);
  and AND2_397 (N1913, N2012, N16);
  and AND2_398 (N1914, N2014, N16);
  and AND2_399 (N1915, N2016, N16);
  and AND2_400 (N1916, N2018, N16);
  and AND2_401 (N1917, N2020, N16);
  and AND2_402 (N1918, N2022, N16);
  and AND2_404 (N1928, N1676, N29);
  and AND2_405 (N1929, N1681, N29);
  and AND2_406 (N1930, N1686, N29);
  and AND2_407 (N1931, N1690, N29);
  and AND2_408 (N1932, N1637, N29);
  and AND2_409 (N1933, N1642, N29);
  and AND2_410 (N1934, N1647, N29);
  and AND2_411 (N1935, N1651, N29);
  and AND2_467 (N2125, N1596, N537);
  and AND2_468 (N2126, N2012, N246);
  and AND2_469 (N2127, N2010, N537);
  and AND2_476 (N2153, N727, N1885);
  and AND2_477 (N2154, N1885, N1651);
  and AND2_478 (N2155, N730, N1888);
  and AND2_479 (N2156, N1888, N1656);
  and AND2_559 (N2358, N2120, N533);
  and AND2_573 (N2386, N2120, N246);
  and AND2_653 (N2607, N2022, N2359);
  and AND2_654 (N2608, N1676, N2359);
  and AND2_655 (N2609, N1681, N2359);
  and AND2_656 (N2610, N1686, N2359);
  and AND2_657 (N2611, N2014, N2113);
  and AND2_658 (N2612, N2016, N2113);
  and AND2_748 (N2789, N2014, N2359);
  and AND2_749 (N2790, N2016, N2359);
  and AND2_750 (N2791, N2018, N2359);
  and AND2_751 (N2792, N2020, N2359);
  and AND2_761 (N2925, N2743, N14);
  and AND2_784 (N2894, N2607, N2250);
  and AND2_785 (N2895, N2608, N2250);
  and AND2_786 (N2896, N2609, N2250);
  and AND2_787 (N2897, N2610, N2250);
  and AND2_790 (N2900, N2791, N8);
  and AND2_791 (N2901, N2792, N8);
  and AND2_811 (N2984, N2898, N8);
  and AND2_812 (N2985, N2899, N8);
  and AND2_820 (N3007, N574, N2359);
  and AND2_832 (N3035, N578, N2359);
  and AND2_833 (N3036, N655, N2359);
  and AND2_834 (N3037, N659, N2359);
  and AND2_844 (N3053, N663, N2359);
  and AND2_845 (N3054, N667, N2359);
  and AND2_846 (N3055, N671, N2359);
  and AND2_847 (N3056, N675, N2359);
  and AND2_848 (N3057, N679, N2359);
  and AND2_849 (N3058, N683, N2359);
  and AND2_850 (N3059, N687, N2359);
  and AND2_851 (N3060, N705, N2359);
  and AND2_871 (N3137, N3055, N8);
  and AND2_872 (N3140, N3056, N8);
  and AND2_873 (N3143, N3057, N2250);
  and AND2_874 (N3146, N3058, N2250);
  and AND2_875 (N3149, N3059, N2250);
  and AND2_876 (N3152, N3060, N2250);
  and AND2_898 (N3197, N687, N2113);
  and AND2_900 (N3215, N705, N2113);
  and AND2_901 (N3216, N711, N2113);
  and AND2_902 (N3217, N715, N2113);
  and AND2_906 (N3222, N719, N2113);
  and AND2_907 (N3223, N723, N2113);
  and AND2_931 (N3291, N3152, N2981);
  and AND2_932 (N3293, N3149, N2978);
  and AND2_934 (N3296, N2972, N3143);
  and AND2_935 (N3299, N3140, N2989);
  and AND2_936 (N3301, N3137, N2986);
  and AND2_993 (N3450, N3334, N8);
  and AND2_994 (N3453, N3335, N8);
  and AND2_997 (N3478, N3400, N533);
  and AND2_998 (N3479, N3318, N2128);
  and AND2_999 (N3480, N3315, N1827);
  and AND2_1050 (N3559, N3450, N3088);
  and AND2_1071 (N3671, N3551, N800);
  and AND2_1118 (N3732, N3603, N3293);
  and AND2_1121 (N3735, N3616, N3301);
  and AND2_1135 (N3753, N3722, N246);
  and AND2_1144 (N3778, N3723, N3480);
  and AND2_1147 (N3809, N3750, N800);
  and AND2_1174 (N3835, N3818, N3823);
  and AND2_1177 (N3838, N3762, N3834);
  and AND3_22 (N495, N2, N15, N237);
  and AND3_114 (N1064, N80, N227, N234);
  and AND3_115 (N1065, N68, N227, N234);
  and AND3_116 (N1066, N79, N227, N234);
  and AND3_117 (N1067, N78, N227, N234);
  and AND3_118 (N1068, N77, N227, N234);
  and AND3_123 (N1097, N76, N227, N234);
  and AND3_124 (N1098, N75, N227, N234);
  and AND3_125 (N1099, N74, N227, N234);
  and AND3_126 (N1100, N73, N227, N234);
  and AND3_127 (N1101, N72, N227, N234);
  and AND3_130 (N1124, N114, N319, N322);
  and AND3_131 (N1125, N113, N319, N322);
  and AND3_132 (N1126, N112, N319, N322);
  and AND3_133 (N1127, N111, N319, N322);
  and AND3_146 (N1168, N118, N319, N322);
  and AND3_147 (N1169, N107, N319, N322);
  and AND3_148 (N1170, N117, N319, N322);
  and AND3_149 (N1171, N116, N319, N322);
  and AND3_150 (N1172, N115, N319, N322);
  and AND3_214 (N1451, N93, N1042, N1053);
  and AND3_215 (N1452, N55, N227, N1053);
  and AND3_216 (N1453, N67, N1042, N234);
  and AND3_217 (N1454, N81, N1042, N1053);
  and AND3_218 (N1455, N43, N227, N1053);
  and AND3_219 (N1456, N56, N1042, N234);
  and AND3_220 (N1457, N92, N1042, N1053);
  and AND3_221 (N1458, N54, N227, N1053);
  and AND3_222 (N1459, N66, N1042, N234);
  and AND3_223 (N1460, N91, N1042, N1053);
  and AND3_224 (N1461, N53, N227, N1053);
  and AND3_225 (N1462, N65, N1042, N234);
  and AND3_226 (N1463, N90, N1042, N1053);
  and AND3_227 (N1464, N52, N227, N1053);
  and AND3_228 (N1465, N64, N1042, N234);
  and AND3_229 (N1466, N89, N1042, N1053);
  and AND3_230 (N1467, N51, N227, N1053);
  and AND3_231 (N1468, N63, N1042, N234);
  and AND3_232 (N1469, N88, N1042, N1053);
  and AND3_233 (N1470, N50, N227, N1053);
  and AND3_234 (N1471, N62, N1042, N234);
  and AND3_235 (N1472, N87, N1042, N1053);
  and AND3_236 (N1473, N49, N227, N1053);
  and AND3_238 (N1475, N86, N1042, N1053);
  and AND3_239 (N1476, N48, N227, N1053);
  and AND3_240 (N1477, N61, N1042, N234);
  and AND3_241 (N1478, N85, N1042, N1053);
  and AND3_242 (N1479, N47, N227, N1053);
  and AND3_243 (N1480, N60, N1042, N234);
  and AND3_244 (N1481, N138, N1102, N1113);
  and AND3_245 (N1482, N102, N319, N1113);
  and AND3_246 (N1483, N126, N1102, N322);
  and AND3_247 (N1484, N137, N1102, N1113);
  and AND3_248 (N1485, N101, N319, N1113);
  and AND3_249 (N1486, N125, N1102, N322);
  and AND3_250 (N1487, N136, N1102, N1113);
  and AND3_251 (N1488, N100, N319, N1113);
  and AND3_252 (N1489, N124, N1102, N322);
  and AND3_253 (N1490, N135, N1102, N1113);
  and AND3_254 (N1491, N99, N319, N1113);
  and AND3_255 (N1492, N123, N1102, N322);
  and AND3_276 (N1529, N142, N1102, N1113);
  and AND3_277 (N1530, N106, N319, N1113);
  and AND3_278 (N1531, N130, N1102, N322);
  and AND3_279 (N1532, N131, N1102, N1113);
  and AND3_280 (N1533, N95, N319, N1113);
  and AND3_281 (N1534, N119, N1102, N322);
  and AND3_282 (N1535, N141, N1102, N1113);
  and AND3_283 (N1536, N105, N319, N1113);
  and AND3_284 (N1537, N129, N1102, N322);
  and AND3_285 (N1538, N140, N1102, N1113);
  and AND3_286 (N1539, N104, N319, N1113);
  and AND3_287 (N1540, N128, N1102, N322);
  and AND3_288 (N1541, N139, N1102, N1113);
  and AND3_289 (N1542, N103, N319, N1113);
  and AND3_290 (N1543, N127, N1102, N322);
  and AND3_350 (N1784, N1133, N1129, N1137);
  and AND3_351 (N1785, N1499, N1496, N1137);
  and AND3_392 (N1908, N1496, N1133, N1776);
  and AND3_393 (N1909, N1129, N1499, N1776);
  and AND3_439 (N2032, N1506, N1502, N1510);
  and AND3_440 (N2033, N1773, N1770, N1510);
  and AND3_444 (N2042, N1557, N1553, N1561);
  and AND3_445 (N2043, N1798, N1795, N1561);
  and AND3_464 (N2113, N1816, N1894, N40);
  and AND3_480 (N2157, N1770, N1506, N2028);
  and AND3_481 (N2158, N1502, N1773, N2028);
  and AND3_488 (N2177, N1795, N1557, N2040);
  and AND3_489 (N2178, N1553, N1798, N2040);
  and AND3_507 (N2250, N40, N1816, N2119);
  and AND3_769 (N2839, N2421, N2417, N2425);
  and AND3_770 (N2840, N2684, N2681, N2425);
  and AND3_802 (N2938, N2681, N2421, N2837);
  and AND3_803 (N2939, N2417, N2684, N2837);
  and AND3_892 (N3191, N2796, N2613, N2800);
  and AND3_893 (N3192, N2992, N2793, N2800);
  and AND3_894 (N3193, N2613, N2120, N2796);
  and AND3_895 (N3194, N2793, N2469, N2796);
  and AND3_924 (N3281, N2793, N2796, N3187);
  and AND3_925 (N3282, N2613, N2992, N3187);
  and AND3_926 (N3283, N2469, N2613, N2992);
  and AND3_927 (N3284, N2120, N2793, N2992);
  and AND3_1171 (N3826, N3727, N3819, N2841);
  and AND3_1191 (N3881, N3826, N3876, N1726);
  and AND4_12 (N485, N309, N305, N301, N297);
  and AND4_33 (N544, N132, N82, N96, N44);
  and AND4_34 (N547, N120, N57, N108, N69);
  and AND4_370 (N1822, N237, N224, N36, N1726);
  and AND4_371 (N1823, N237, N224, N1726, N486);
  and AND4_1117 (N3731, N3608, N3615, N3612, N3603);
  and AND4_1120 (N3734, N3612, N3603, N3296, N3608);
  and AND4_1155 (N3807, N3754, N3616, N3559, N3622);
  nand NAND2_96 (N900, N331, N606);
  nand NAND2_97 (N901, N328, N607);
  nand NAND2_98 (N902, N337, N608);
  nand NAND2_99 (N903, N334, N609);
  nand NAND2_100 (N904, N343, N610);
  nand NAND2_101 (N905, N340, N611);
  nand NAND2_102 (N998, N349, N733);
  nand NAND2_103 (N999, N346, N734);
  nand NAND2_107 (N1029, N231, N651);
  nand NAND2_135 (N1129, N900, N901);
  nand NAND2_136 (N1133, N902, N903);
  nand NAND2_137 (N1137, N904, N905);
  nand NAND2_139 (N1141, N263, N612);
  nand NAND2_154 (N1185, N294, N650);
  nand NAND2_169 (N1216, N998, N999);
  nand NAND2_193 (N1351, N352, N655);
  nand NAND2_194 (N1352, N266, N663);
  nand NAND2_195 (N1353, N269, N659);
  nand NAND2_196 (N1354, N272, N671);
  nand NAND2_197 (N1355, N275, N667);
  nand NAND2_198 (N1395, N355, N705);
  nand NAND2_199 (N1396, N297, N715);
  nand NAND2_200 (N1397, N301, N711);
  nand NAND2_201 (N1398, N305, N723);
  nand NAND2_202 (N1399, N309, N719);
  nand NAND2_203 (N1422, N256, N578);
  nand NAND2_204 (N1423, N259, N574);
  nand NAND2_205 (N1424, N278, N679);
  nand NAND2_206 (N1425, N281, N675);
  nand NAND2_207 (N1426, N284, N687);
  nand NAND2_208 (N1427, N287, N683);
  nand NAND2_209 (N1440, N313, N730);
  nand NAND2_210 (N1441, N316, N727);
  nand NAND2_261 (N1502, N1351, N1141);
  nand NAND2_262 (N1506, N1352, N1353);
  nand NAND2_263 (N1510, N1354, N1355);
  nand NAND2_300 (N1553, N1395, N1185);
  nand NAND2_301 (N1557, N1396, N1397);
  nand NAND2_302 (N1561, N1398, N1399);
  nand NAND2_317 (N1578, N1422, N1423);
  nand NAND2_319 (N1582, N1426, N1427);
  nand NAND2_320 (N1585, N1424, N1425);
  nand NAND2_321 (N1588, N1440, N1441);
  nand NAND2_358 (N1809, N1578, N1581);
  nand NAND2_387 (N1885, N727, N1651);
  nand NAND2_388 (N1888, N730, N1656);
  nand NAND2_413 (N1939, N1216, N1808);
  nand NAND2_414 (N1940, N1585, N1810);
  nand NAND2_415 (N1941, N1582, N1811);
  nand NAND2_446 (N2046, N1939, N1809);
  nand NAND2_447 (N2049, N1940, N1941);
  nand NAND2_466 (N2120, N408, N1827);
  nand NAND2_483 (N2172, N1676, N1919);
  nand NAND2_502 (N2219, N2031, N2030);
  nand NAND2_516 (N2302, N2052, N256);
  nand NAND2_518 (N2304, N2055, N259);
  nand NAND2_520 (N2306, N2058, N263);
  nand NAND2_522 (N2308, N2061, N266);
  nand NAND2_524 (N2310, N2064, N269);
  nand NAND2_526 (N2312, N2067, N272);
  nand NAND2_528 (N2314, N2070, N275);
  nand NAND2_530 (N2316, N2073, N278);
  nand NAND2_532 (N2318, N2076, N281);
  nand NAND2_534 (N2320, N2079, N284);
  nand NAND2_536 (N2322, N1708, N2171);
  nand NAND2_537 (N2323, N1681, N2173);
  nand NAND2_538 (N2324, N1686, N2174);
  nand NAND2_539 (N2325, N1690, N1818);
  nand NAND2_540 (N2326, N1637, N2176);
  nand NAND2_543 (N2329, N2095, N287);
  nand NAND2_545 (N2331, N2098, N294);
  nand NAND2_547 (N2333, N2101, N297);
  nand NAND2_549 (N2335, N2104, N301);
  nand NAND2_551 (N2337, N2107, N305);
  nand NAND2_553 (N2339, N2110, N309);
  nand NAND2_555 (N2354, N1642, N1817);
  nand NAND2_556 (N2355, N1647, N1816);
  nand NAND2_557 (N2356, N1651, N2236);
  nand NAND2_558 (N2357, N1656, N2237);
  nand NAND2_580 (N2400, N2219, N2300);
  nand NAND2_583 (N2407, N574, N2303);
  nand NAND2_584 (N2408, N578, N2305);
  nand NAND2_585 (N2409, N655, N2307);
  nand NAND2_586 (N2410, N659, N2309);
  nand NAND2_587 (N2411, N663, N2311);
  nand NAND2_588 (N2412, N667, N2313);
  nand NAND2_589 (N2413, N671, N2315);
  nand NAND2_590 (N2414, N675, N2317);
  nand NAND2_591 (N2415, N679, N2319);
  nand NAND2_592 (N2416, N683, N2321);
  nand NAND2_593 (N2417, N2322, N2172);
  nand NAND2_594 (N2421, N2323, N2324);
  nand NAND2_595 (N2425, N2325, N2326);
  nand NAND2_596 (N2428, N687, N2330);
  nand NAND2_597 (N2429, N705, N2332);
  nand NAND2_598 (N2430, N711, N2334);
  nand NAND2_599 (N2431, N715, N2336);
  nand NAND2_600 (N2432, N719, N2338);
  nand NAND2_601 (N2433, N723, N2340);
  nand NAND2_609 (N2453, N1606, N1836);
  nand NAND2_620 (N2484, N2298, N2297);
  nand NAND2_621 (N2487, N2356, N2357);
  nand NAND2_622 (N2490, N2354, N2355);
  nand NAND2_623 (N2493, N2328, N2327);
  nand NAND2_625 (N2503, N1833, N1600);
  nand NAND2_626 (N2504, N1836, N1596);
  nand NAND2_630 (N2528, N2046, N2406);
  nand NAND2_651 (N2579, N1600, N1827);
  nand NAND2_659 (N2613, N2503, N2504);
  nand NAND2_661 (N2618, N2128, N1606);
  nand NAND2_662 (N2619, N1821, N2014);
  nand NAND2_680 (N2652, N2528, N2400);
  nand NAND2_685 (N2664, N2484, N2301);
  nand NAND2_707 (N2694, N2493, N1807);
  nand NAND2_716 (N2703, N2579, N2453);
  nand NAND2_722 (N2719, N1827, N2010);
  nand NAND2_723 (N2720, N1820, N2012);
  nand NAND2_728 (N2747, N2049, N2663);
  nand NAND2_733 (N2760, N1588, N2693);
  nand NAND2_736 (N2771, N1819, N2018);
  nand NAND2_737 (N2772, N2144, N2016);
  nand NAND2_738 (N2773, N2147, N2022);
  nand NAND2_739 (N2774, N2150, N2020);
  nand NAND2_744 (N2781, N2490, N2707);
  nand NAND2_745 (N2782, N2487, N2708);
  nand NAND2_753 (N2796, N2719, N2618);
  nand NAND2_754 (N2800, N2619, N2720);
  nand NAND2_763 (N2826, N2747, N2664);
  nand NAND2_771 (N2841, N2760, N2694);
  nand NAND2_776 (N2874, N2773, N2774);
  nand NAND2_777 (N2877, N2771, N2772);
  nand NAND2_779 (N2881, N2703, N2120);
  nand NAND2_782 (N2888, N2781, N2782);
  nand NAND2_783 (N2891, N2534, N2531);
  nand NAND2_804 (N2963, N2469, N2880);
  nand NAND2_865 (N3076, N2881, N2963);
  nand NAND2_883 (N3175, N2877, N3072);
  nand NAND2_884 (N3176, N2874, N3073);
  nand NAND2_887 (N3180, N3048, N3047);
  nand NAND2_896 (N3195, N3076, N1833);
  nand NAND2_910 (N3238, N3175, N3176);
  nand NAND2_928 (N3286, N1596, N3196);
  nand NAND2_930 (N3289, N3180, N3049);
  nand NAND2_971 (N3400, N3195, N3286);
  nand NAND2_979 (N3410, N2888, N3333);
  nand NAND2_1000 (N3481, N3410, N3289);
  nand NAND2_1002 (N3483, N3152, N2897);
  nand NAND2_1004 (N3485, N3149, N2896);
  nand NAND2_1006 (N3487, N3146, N2895);
  nand NAND2_1008 (N3489, N3143, N2894);
  nand NAND2_1010 (N3491, N3140, N2901);
  nand NAND2_1012 (N3493, N3137, N2900);
  nand NAND2_1033 (N3522, N3402, N3401);
  nand NAND2_1034 (N3525, N3404, N3403);
  nand NAND2_1043 (N3552, N2981, N3482);
  nand NAND2_1044 (N3553, N2978, N3484);
  nand NAND2_1045 (N3554, N2975, N3486);
  nand NAND2_1046 (N3555, N2972, N3488);
  nand NAND2_1047 (N3556, N2989, N3490);
  nand NAND2_1048 (N3557, N2986, N3492);
  nand NAND2_1064 (N3593, N3522, N3405);
  nand NAND2_1066 (N3595, N3525, N3405);
  nand NAND2_1068 (N3597, N3318, N2010);
  nand NAND2_1069 (N3598, N3315, N1606);
  nand NAND2_1072 (N3603, N3552, N3483);
  nand NAND2_1073 (N3608, N3553, N3485);
  nand NAND2_1074 (N3612, N3554, N3487);
  nand NAND2_1075 (N3615, N3555, N3489);
  nand NAND2_1076 (N3616, N3556, N3491);
  nand NAND2_1077 (N3622, N3557, N3493);
  nand NAND2_1079 (N3630, N3321, N2012);
  nand NAND2_1092 (N3667, N3238, N3592);
  nand NAND2_1093 (N3668, N3238, N3594);
  nand NAND2_1094 (N3669, N2128, N3596);
  nand NAND2_1095 (N3670, N1827, N3599);
  nand NAND2_1098 (N3692, N3453, N2985);
  nand NAND2_1100 (N3694, N3450, N2984);
  nand NAND2_1101 (N3695, N1821, N3629);
  nand NAND2_1109 (N3721, N3667, N3593);
  nand NAND2_1110 (N3722, N3668, N3595);
  nand NAND2_1111 (N3723, N3669, N3597);
  nand NAND2_1112 (N3726, N3670, N3598);
  nand NAND2_1114 (N3728, N3091, N3691);
  nand NAND2_1115 (N3729, N3088, N3693);
  nand NAND2_1116 (N3730, N3695, N3630);
  nand NAND2_1136 (N3754, N3728, N3692);
  nand NAND2_1137 (N3758, N3729, N3694);
  nand NAND2_1165 (N3818, N3805, N3761);
  nor NOR2_437 (N2030, N1908, N1784);
  nor NOR2_438 (N2031, N1909, N1785);
  nor NOR2_512 (N2297, N2157, N2032);
  nor NOR2_513 (N2298, N2158, N2033);
  nor NOR2_541 (N2327, N2177, N2042);
  nor NOR2_542 (N2328, N2178, N2043);
  nor NOR2_840 (N3047, N2938, N2839);
  nor NOR2_841 (N3048, N2939, N2840);
  nor NOR2_972 (N3401, N3281, N3191);
  nor NOR2_973 (N3402, N3282, N3192);
  nor NOR2_974 (N3403, N3283, N3193);
  nor NOR2_975 (N3404, N3284, N3194);
  not NOT1_5 (N408, N230);
  not NOT1_8 (N425, N262);
  not NOT1_13 (N486, N405);
  not NOT1_14 (N487, N44);
  not NOT1_15 (N488, N132);
  not NOT1_16 (N489, N82);
  not NOT1_17 (N490, N96);
  not NOT1_18 (N491, N69);
  not NOT1_19 (N492, N120);
  not NOT1_20 (N493, N57);
  not NOT1_21 (N494, N108);
  not NOT1_30 (N533, N241);
  not NOT1_31 (N537, N246);
  not NOT1_37 (N574, N256);
  not NOT1_38 (N578, N259);
  not NOT1_41 (N606, N328);
  not NOT1_42 (N607, N331);
  not NOT1_43 (N608, N334);
  not NOT1_44 (N609, N337);
  not NOT1_45 (N610, N340);
  not NOT1_46 (N611, N343);
  not NOT1_47 (N612, N352);
  not NOT1_52 (N650, N355);
  not NOT1_54 (N655, N263);
  not NOT1_55 (N659, N266);
  not NOT1_56 (N663, N269);
  not NOT1_57 (N667, N272);
  not NOT1_58 (N671, N275);
  not NOT1_59 (N675, N278);
  not NOT1_60 (N679, N281);
  not NOT1_61 (N683, N284);
  not NOT1_62 (N687, N287);
  not NOT1_65 (N705, N294);
  not NOT1_66 (N711, N297);
  not NOT1_67 (N715, N301);
  not NOT1_68 (N719, N305);
  not NOT1_69 (N723, N309);
  not NOT1_70 (N727, N313);
  not NOT1_71 (N730, N316);
  not NOT1_72 (N733, N346);
  not NOT1_73 (N734, N349);
  not NOT1_92 (N792, N485);
  not NOT1_93 (N799, N495);
  not NOT1_94 (N800, N37);
  not NOT1_106 (N1028, N651);
  not NOT1_108 (N1032, N544);
  not NOT1_109 (N1033, N547);
  not NOT1_112 (N1042, N227);
  not NOT1_113 (N1053, N234);
  not NOT1_128 (N1102, N319);
  not NOT1_129 (N1113, N322);
  not NOT1_151 (N1173, N16);
  not NOT1_161 (N1200, N29);
  not NOT1_188 (N1269, N1027);
  not NOT1_211 (N1448, N1277);
  not NOT1_212 (N1449, N1275);
  not NOT1_213 (N1450, N1276);
  not NOT1_259 (N1496, N1129);
  not NOT1_260 (N1499, N1133);
  not NOT1_318 (N1581, N1216);
  not NOT1_344 (N1770, N1502);
  not NOT1_345 (N1773, N1506);
  not NOT1_346 (N1776, N1137);
  not NOT1_352 (N1795, N1553);
  not NOT1_353 (N1798, N1557);
  not NOT1_356 (N1807, N1588);
  not NOT1_357 (N1808, N1578);
  not NOT1_359 (N1810, N1582);
  not NOT1_360 (N1811, N1585);
  not NOT1_364 (N1816, N1642);
  not NOT1_365 (N1817, N1647);
  not NOT1_366 (N1818, N1637);
  not NOT1_367 (N1819, N2016);
  not NOT1_368 (N1820, N2014);
  not NOT1_369 (N1821, N2012);
  not NOT1_373 (N1827, N1606);
  not NOT1_377 (N1833, N1596);
  not NOT1_378 (N1836, N1600);
  not NOT1_403 (N1919, N1708);
  not NOT1_426 (N1970, N1822);
  not NOT1_427 (N1971, N1823);
  not NOT1_435 (N2028, N1510);
  not NOT1_442 (N2040, N1561);
  not NOT1_465 (N2119, N1894);
  not NOT1_470 (N2128, N2010);
  not NOT1_473 (N2144, N2018);
  not NOT1_474 (N2147, N2020);
  not NOT1_475 (N2150, N2022);
  not NOT1_482 (N2171, N1676);
  not NOT1_484 (N2173, N1686);
  not NOT1_485 (N2174, N1681);
  not NOT1_487 (N2176, N1690);
  not NOT1_505 (N2236, N1656);
  not NOT1_506 (N2237, N1651);
  not NOT1_514 (N2300, N2046);
  not NOT1_515 (N2301, N2049);
  not NOT1_517 (N2303, N2052);
  not NOT1_519 (N2305, N2055);
  not NOT1_521 (N2307, N2058);
  not NOT1_523 (N2309, N2061);
  not NOT1_525 (N2311, N2064);
  not NOT1_527 (N2313, N2067);
  not NOT1_529 (N2315, N2070);
  not NOT1_531 (N2317, N2073);
  not NOT1_533 (N2319, N2076);
  not NOT1_535 (N2321, N2079);
  not NOT1_544 (N2330, N2095);
  not NOT1_546 (N2332, N2098);
  not NOT1_548 (N2334, N2101);
  not NOT1_550 (N2336, N2104);
  not NOT1_552 (N2338, N2107);
  not NOT1_554 (N2340, N2110);
  not NOT1_560 (N2359, N2113);
  not NOT1_582 (N2406, N2219);
  not NOT1_615 (N2469, N2120);
  not NOT1_631 (N2531, N2291);
  not NOT1_632 (N2534, N2294);
  not NOT1_684 (N2663, N2484);
  not NOT1_702 (N2681, N2417);
  not NOT1_703 (N2684, N2421);
  not NOT1_706 (N2693, N2493);
  not NOT1_718 (N2707, N2487);
  not NOT1_719 (N2708, N2490);
  not NOT1_727 (N2743, N2652);
  not NOT1_752 (N2793, N2613);
  not NOT1_767 (N2837, N2425);
  not NOT1_778 (N2880, N2703);
  not NOT1_805 (N2970, N2841);
  not NOT1_806 (N2971, N2826);
  not NOT1_807 (N2972, N2894);
  not NOT1_808 (N2975, N2895);
  not NOT1_809 (N2978, N2896);
  not NOT1_810 (N2981, N2897);
  not NOT1_813 (N2986, N2900);
  not NOT1_814 (N2989, N2901);
  not NOT1_815 (N2992, N2796);
  not NOT1_829 (N3028, N2925);
  not NOT1_842 (N3049, N2888);
  not NOT1_861 (N3072, N2874);
  not NOT1_862 (N3073, N2877);
  not NOT1_866 (N3079, N3038);
  not NOT1_867 (N3088, N2984);
  not NOT1_868 (N3091, N2985);
  not NOT1_888 (N3187, N2800);
  not NOT1_897 (N3196, N3076);
  not NOT1_950 (N3333, N3180);
  not NOT1_976 (N3405, N3238);
  not NOT1_1001 (N3482, N3152);
  not NOT1_1003 (N3484, N3149);
  not NOT1_1005 (N3486, N3146);
  not NOT1_1007 (N3488, N3143);
  not NOT1_1009 (N3490, N3140);
  not NOT1_1011 (N3492, N3137);
  not NOT1_1042 (N3551, N3481);
  not NOT1_1063 (N3592, N3522);
  not NOT1_1065 (N3594, N3525);
  not NOT1_1067 (N3596, N3318);
  not NOT1_1070 (N3599, N3315);
  not NOT1_1078 (N3629, N3321);
  not NOT1_1097 (N3691, N3453);
  not NOT1_1099 (N3693, N3450);
  not NOT1_1113 (N3727, N3671);
  not NOT1_1134 (N3750, N3721);
  not NOT1_1138 (N3761, N3731);
  not NOT1_1153 (N3805, N3762);
  not NOT1_1166 (N3819, N3809);
  not NOT1_1173 (N3834, N3823);
  not NOT1_1193 (N3882, N3881);
  or OR2_192 (N1302, N1069, N543);
  or OR2_425 (N1969, N533, N1815);
  or OR2_441 (N2034, N1571, N1935);
  or OR2_448 (N2052, N1544, N1910);
  or OR2_449 (N2055, N1545, N1911);
  or OR2_450 (N2058, N1546, N1912);
  or OR2_451 (N2061, N1547, N1913);
  or OR2_452 (N2064, N1548, N1914);
  or OR2_453 (N2067, N1549, N1915);
  or OR2_454 (N2070, N1550, N1916);
  or OR2_455 (N2073, N1551, N1917);
  or OR2_456 (N2076, N1552, N1918);
  or OR2_457 (N2079, N1564, N1928);
  or OR2_458 (N2095, N1565, N1929);
  or OR2_459 (N2098, N1566, N1930);
  or OR2_460 (N2101, N1567, N1931);
  or OR2_461 (N2104, N1568, N1932);
  or OR2_462 (N2107, N1569, N1933);
  or OR2_463 (N2110, N1570, N1934);
  or OR2_508 (N2387, N1831, N2126);
  or OR2_509 (N2389, N2127, N1832);
  or OR2_510 (N2291, N2153, N2154);
  or OR2_511 (N2294, N2155, N2156);
  or OR2_624 (N2496, N2358, N1814);
  or OR2_629 (N2643, N1830, N2386);
  or OR2_788 (N2898, N2789, N2611);
  or OR2_789 (N2899, N2790, N2612);
  or OR2_929 (N3288, N3197, N3007);
  or OR2_944 (N3315, N3215, N3035);
  or OR2_945 (N3318, N3216, N3036);
  or OR2_946 (N3321, N3217, N3037);
  or OR2_951 (N3334, N3222, N3053);
  or OR2_952 (N3335, N3223, N3054);
  or OR2_1041 (N3546, N3478, N1813);
  or OR2_1146 (N3803, N2125, N3753);
  or OR2_1179 (N3851, N3838, N3835);
  or OR3_1150 (N3802, N3479, N3778, N3779);
  or OR4_323 (N1596, N1451, N1452, N1453, N1064);
  or OR4_324 (N1600, N1454, N1455, N1456, N1065);
  or OR4_325 (N1606, N1457, N1458, N1459, N1066);
  or OR4_326 (N2010, N1460, N1461, N1462, N1067);
  or OR4_327 (N2012, N1463, N1464, N1465, N1068);
  or OR4_328 (N2014, N1466, N1467, N1468, N1097);
  or OR4_329 (N2016, N1469, N1470, N1471, N1098);
  or OR4_330 (N2018, N1472, N1473, N1474, N1099);
  or OR4_331 (N2020, N1475, N1476, N1477, N1100);
  or OR4_332 (N2022, N1478, N1479, N1480, N1101);
  or OR4_333 (N1637, N1481, N1482, N1483, N1124);
  or OR4_334 (N1642, N1484, N1485, N1486, N1125);
  or OR4_335 (N1647, N1487, N1488, N1489, N1126);
  or OR4_336 (N1651, N1490, N1491, N1492, N1127);
  or OR4_337 (N1656, N1493, N1494, N1495, N1128);
  or OR4_338 (N1676, N1532, N1533, N1534, N1169);
  or OR4_339 (N1681, N1535, N1536, N1537, N1170);
  or OR4_340 (N1686, N1538, N1539, N1540, N1171);
  or OR4_341 (N1690, N1541, N1542, N1543, N1172);
  or OR4_342 (N1708, N1529, N1530, N1531, N1168);
  or OR4_1139 (N3762, N3291, N3732, N3733, N3734);
  and g2 (N3876, N2826, N3028);
  and g3 (n_374, N2320, N2416, N2318);
  and g4 (n_375, N2415, N2316, N2414);
  and g5 (n_376, N2314, N2413);
  and g6 (n_377, N2312, N2412);
  and g7 (n_378, N2310, N2411);
  and g8 (n_379, N2308, N2410);
  and g9 (n_380, N2306, N2409);
  and g10 (n_381, N2304, N2408);
  and g11 (n_382, N2302, N2407);
  and g12 (n_383, N2034, N2339);
  and g13 (n_384, N2433, N2337);
  and g14 (n_385, N2432, N2335);
  and g15 (n_386, N2431, N2333);
  and g16 (n_387, N2430, N2331);
  and g17 (n_388, N2429, N2329);
  and g18 (n_389, N2428, N1302);
  and g19 (n_390, n_374, n_375, n_376, n_377);
  and g20 (n_391, n_378, n_379, n_380, n_381);
  and g21 (n_392, n_382, n_383, n_384, n_385);
  and g22 (n_393, n_386, n_387, n_388, n_389);
  and g23 (N3038, n_390, n_391, n_392, n_393);
  or g24 (n_394, N3299, N3735);
  or g25 (n_395, N3736, N3807);
  or g26 (N3823, N3808, N3817, n_394, n_395);
  and g27 (N3733, N3608, N3603, N3146, N2975);
  and g28 (N3736, N3622, N3616, N3453, N3091);
  and g29 (n_396, N3758, N3754);
  and g30 (n_397, N3616, N3321);
  and g31 (N3808, N1821, N3622, n_396, n_397);
  and g32 (n_398, N3622, N3730);
  and g33 (n_399, N3754, N3616);
  and g34 (N3817, N3758, N3802, n_398, n_399);
  and g35 (N3779, N3726, N3723, N3288, N1836);
endmodule

