
module adder(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] ,
     \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14]
     , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
     \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
     \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
     \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
     \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
     \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
     \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
     \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
     \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
     \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
     \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
     \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
     \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105]
     , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] ,
     \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
     \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
     \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] ,
     \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] ,
     \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
     \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
     \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] ,
     \b[32] , \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] ,
     \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] , \b[45] ,
     \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
     \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
     \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] ,
     \b[67] , \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] ,
     \b[74] , \b[75] , \b[76] , \b[77] , \b[78] , \b[79] , \b[80] ,
     \b[81] , \b[82] , \b[83] , \b[84] , \b[85] , \b[86] , \b[87] ,
     \b[88] , \b[89] , \b[90] , \b[91] , \b[92] , \b[93] , \b[94] ,
     \b[95] , \b[96] , \b[97] , \b[98] , \b[99] , \b[100] , \b[101] ,
     \b[102] , \b[103] , \b[104] , \b[105] , \b[106] , \b[107] ,
     \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
     \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] ,
     \b[120] , \b[121] , \b[122] , \b[123] , \b[124] , \b[125] ,
     \b[126] , \b[127] , \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5]
     , \f[6] , \f[7] , \f[8] , \f[9] , \f[10] , \f[11] , \f[12] ,
     \f[13] , \f[14] , \f[15] , \f[16] , \f[17] , \f[18] , \f[19] ,
     \f[20] , \f[21] , \f[22] , \f[23] , \f[24] , \f[25] , \f[26] ,
     \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] , \f[33] ,
     \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
     \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
     \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] ,
     \f[55] , \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] ,
     \f[62] , \f[63] , \f[64] , \f[65] , \f[66] , \f[67] , \f[68] ,
     \f[69] , \f[70] , \f[71] , \f[72] , \f[73] , \f[74] , \f[75] ,
     \f[76] , \f[77] , \f[78] , \f[79] , \f[80] , \f[81] , \f[82] ,
     \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] , \f[89] ,
     \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
     \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
     \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
     \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] ,
     \f[116] , \f[117] , \f[118] , \f[119] , \f[120] , \f[121] ,
     \f[122] , \f[123] , \f[124] , \f[125] , \f[126] , \f[127] , cOut);
//   input \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
       \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
       \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
       \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
       \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
       \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] ,
       \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
       \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
       \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] ,
       \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1]
       , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9]
       , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
       \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] ,
       \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] ,
       \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] , \b[37] ,
       \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
       \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
       \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] ,
       \b[59] , \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] ,
       \b[66] , \b[67] , \b[68] , \b[69] , \b[70] , \b[71] , \b[72] ,
       \b[73] , \b[74] , \b[75] , \b[76] , \b[77] , \b[78] , \b[79] ,
       \b[80] , \b[81] , \b[82] , \b[83] , \b[84] , \b[85] , \b[86] ,
       \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] , \b[93] ,
       \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] , \b[100] ,
       \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
       \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] ,
       \b[113] , \b[114] , \b[115] , \b[116] , \b[117] , \b[118] ,
       \b[119] , \b[120] , \b[121] , \b[122] , \b[123] , \b[124] ,
       \b[125] , \b[126] , \b[127] ;
//   output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7]
       , \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] ,
       \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] ,
       \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] ,
       \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] ,
       \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] ,
       \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] ,
       \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
       \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
       \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] ,
       \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] ,
       \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] ,
       \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] ,
       \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] ,
       \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] ,
       \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
       \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
       \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] ,
       \f[123] , \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
       \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] ,
       \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] ,
       \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] ,
       \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] ,
       \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] ,
       \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] ,
       \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
       \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
       \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] ,
       \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] ,
       \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] ,
       \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] ,
       \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] ,
       \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] ,
       \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
       \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
       \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] ,
       \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1]
       , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9]
       , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
       \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] ,
       \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] ,
       \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] , \b[37] ,
       \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
       \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
       \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] ,
       \b[59] , \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] ,
       \b[66] , \b[67] , \b[68] , \b[69] , \b[70] , \b[71] , \b[72] ,
       \b[73] , \b[74] , \b[75] , \b[76] , \b[77] , \b[78] , \b[79] ,
       \b[80] , \b[81] , \b[82] , \b[83] , \b[84] , \b[85] , \b[86] ,
       \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] , \b[93] ,
       \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] , \b[100] ,
       \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
       \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] ,
       \b[113] , \b[114] , \b[115] , \b[116] , \b[117] , \b[118] ,
       \b[119] , \b[120] , \b[121] , \b[122] , \b[123] , \b[124] ,
       \b[125] , \b[126] , \b[127] ;
  wire \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
       \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] ,
       \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] ,
       \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] ,
       \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] ,
       \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] ,
       \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] ,
       \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
       \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
       \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] ,
       \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] ,
       \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] ,
       \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] ,
       \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] ,
       \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] ,
       \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
       \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
       \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] ,
       \f[123] , \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire n386, n387, n389, n390, n391, n392, n393, n394;
  wire n396, n397, n398, n399, n400, n401, n402, n404;
  wire n405, n406, n407, n408, n409, n410, n412, n413;
  wire n414, n415, n416, n417, n418, n420, n421, n422;
  wire n423, n424, n425, n426, n428, n429, n430, n431;
  wire n432, n433, n434, n436, n437, n438, n439, n440;
  wire n441, n442, n444, n445, n446, n447, n448, n449;
  wire n450, n452, n453, n454, n455, n456, n457, n458;
  wire n460, n461, n462, n463, n464, n465, n466, n468;
  wire n469, n470, n471, n472, n473, n474, n476, n477;
  wire n478, n479, n480, n481, n482, n484, n485, n486;
  wire n487, n488, n489, n490, n492, n493, n494, n495;
  wire n496, n497, n498, n500, n501, n502, n503, n504;
  wire n505, n506, n508, n509, n510, n511, n512, n513;
  wire n514, n516, n517, n518, n519, n520, n521, n522;
  wire n524, n525, n526, n527, n528, n529, n530, n532;
  wire n533, n534, n535, n536, n537, n538, n540, n541;
  wire n542, n543, n544, n545, n546, n548, n549, n550;
  wire n551, n552, n553, n554, n556, n557, n558, n559;
  wire n560, n561, n562, n564, n565, n566, n567, n568;
  wire n569, n570, n572, n573, n574, n575, n576, n577;
  wire n578, n580, n581, n582, n583, n584, n585, n586;
  wire n588, n589, n590, n591, n592, n593, n594, n596;
  wire n597, n598, n599, n600, n601, n602, n604, n605;
  wire n606, n607, n608, n609, n610, n612, n613, n614;
  wire n615, n616, n617, n618, n620, n621, n622, n623;
  wire n624, n625, n626, n628, n629, n630, n631, n632;
  wire n633, n634, n636, n637, n638, n639, n640, n641;
  wire n642, n644, n645, n646, n647, n648, n649, n650;
  wire n652, n653, n654, n655, n656, n657, n658, n660;
  wire n661, n662, n663, n664, n665, n666, n668, n669;
  wire n670, n671, n672, n673, n674, n676, n677, n678;
  wire n679, n680, n681, n682, n684, n685, n686, n687;
  wire n688, n689, n690, n692, n693, n694, n695, n696;
  wire n697, n698, n700, n701, n702, n703, n704, n705;
  wire n706, n708, n709, n710, n711, n712, n713, n714;
  wire n716, n717, n718, n719, n720, n721, n722, n724;
  wire n725, n726, n727, n728, n729, n730, n732, n733;
  wire n734, n735, n736, n737, n738, n740, n741, n742;
  wire n743, n744, n745, n746, n748, n749, n750, n751;
  wire n752, n753, n754, n756, n757, n758, n759, n760;
  wire n761, n762, n764, n765, n766, n767, n768, n769;
  wire n770, n772, n773, n774, n775, n776, n777, n778;
  wire n780, n781, n782, n783, n784, n785, n786, n788;
  wire n789, n790, n791, n792, n793, n794, n796, n797;
  wire n798, n799, n800, n801, n802, n804, n805, n806;
  wire n807, n808, n809, n810, n812, n813, n814, n815;
  wire n816, n817, n818, n820, n821, n822, n823, n824;
  wire n825, n826, n828, n829, n830, n831, n832, n833;
  wire n834, n836, n837, n838, n839, n840, n841, n842;
  wire n844, n845, n846, n847, n848, n849, n850, n852;
  wire n853, n854, n855, n856, n857, n858, n860, n861;
  wire n862, n863, n864, n865, n866, n868, n869, n870;
  wire n871, n872, n873, n874, n876, n877, n878, n879;
  wire n880, n881, n882, n884, n885, n886, n887, n888;
  wire n889, n890, n892, n893, n894, n895, n896, n897;
  wire n898, n900, n901, n902, n903, n904, n905, n906;
  wire n908, n909, n910, n911, n912, n913, n914, n916;
  wire n917, n918, n919, n920, n921, n922, n924, n925;
  wire n926, n927, n928, n929, n930, n932, n933, n934;
  wire n935, n936, n937, n938, n940, n941, n942, n943;
  wire n944, n945, n946, n948, n949, n950, n951, n952;
  wire n953, n954, n956, n957, n958, n959, n960, n961;
  wire n962, n964, n965, n966, n967, n968, n969, n970;
  wire n972, n973, n974, n975, n976, n977, n978, n980;
  wire n981, n982, n983, n984, n985, n986, n988, n989;
  wire n990, n991, n992, n993, n994, n996, n997, n998;
  wire n999, n1000, n1001, n1002, n1004, n1005, n1006, n1007;
  wire n1008, n1009, n1010, n1012, n1013, n1014, n1015, n1016;
  wire n1017, n1018, n1020, n1021, n1022, n1023, n1024, n1025;
  wire n1026, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  wire n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1044;
  wire n1045, n1046, n1047, n1048, n1049, n1050, n1052, n1053;
  wire n1054, n1055, n1056, n1057, n1058, n1060, n1061, n1062;
  wire n1063, n1064, n1065, n1066, n1068, n1069, n1070, n1071;
  wire n1072, n1073, n1074, n1076, n1077, n1078, n1079, n1080;
  wire n1081, n1082, n1084, n1085, n1086, n1087, n1088, n1089;
  wire n1090, n1092, n1093, n1094, n1095, n1096, n1097, n1098;
  wire n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1108;
  wire n1109, n1110, n1111, n1112, n1113, n1114, n1116, n1117;
  wire n1118, n1119, n1120, n1121, n1122, n1124, n1125, n1126;
  wire n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1135;
  wire n1136, n1137, n1138, n1140, n1141, n1142, n1143, n1144;
  wire n1145, n1146, n1148, n1149, n1150, n1151, n1152, n1153;
  wire n1154, n1156, n1157, n1158, n1159, n1160, n1161, n1162;
  wire n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1172;
  wire n1173, n1174, n1175, n1176, n1177, n1178, n1180, n1181;
  wire n1182, n1183, n1184, n1185, n1186, n1188, n1189, n1190;
  wire n1191, n1192, n1193, n1194, n1196, n1197, n1198, n1199;
  wire n1200, n1201, n1202, n1204, n1205, n1206, n1207, n1208;
  wire n1209, n1210, n1212, n1213, n1214, n1215, n1216, n1217;
  wire n1218, n1220, n1221, n1222, n1223, n1224, n1225, n1226;
  wire n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1236;
  wire n1237, n1238, n1239, n1240, n1241, n1242, n1244, n1245;
  wire n1246, n1247, n1248, n1249, n1250, n1252, n1253, n1254;
  wire n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263;
  wire n1264, n1265, n1266, n1268, n1269, n1270, n1271, n1272;
  wire n1273, n1274, n1276, n1277, n1278, n1279, n1280, n1281;
  wire n1282, n1284, n1285, n1286, n1287, n1288, n1289, n1290;
  wire n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1300;
  wire n1301, n1302, n1303, n1304, n1305, n1306, n1308, n1309;
  wire n1310, n1311, n1312, n1313, n1314, n1316, n1317, n1318;
  wire n1319, n1320, n1321, n1322, n1324, n1325, n1326, n1327;
  wire n1328, n1329, n1330, n1332, n1333, n1334, n1335, n1336;
  wire n1337, n1338, n1340, n1341, n1342, n1343, n1344, n1345;
  wire n1346, n1348, n1349, n1350, n1351, n1352, n1353, n1354;
  wire n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1364;
  wire n1365, n1366, n1367, n1368, n1369, n1370, n1372, n1373;
  wire n1374, n1375, n1376, n1377, n1378, n1380, n1381, n1382;
  wire n1383, n1384, n1385, n1386, n1388, n1389, n1390, n1391;
  wire n1392, n1393, n1394, n1396, n1397, n1398, n1399, n1400;
  wire n1401, n1402, n1404, n_3, n_4, n_7, n_8, n_9;
  wire n_10, n_11, n_12, n_13, n_16, n_17, n_18, n_19;
  wire n_20, n_21, n_22, n_23, n_24, n_27, n_28, n_29;
  wire n_30, n_31, n_32, n_33, n_34, n_35, n_38, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_49;
  wire n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_115, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_123, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_192, n_193, n_194, n_195;
  wire n_196, n_197, n_198, n_199, n_200, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_280, n_281, n_282, n_283;
  wire n_284, n_285, n_286, n_287, n_288, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_387, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_467, n_468, n_469;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_511, n_512, n_513, n_514, n_515, n_516, n_517;
  wire n_518, n_519, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_566, n_567;
  wire n_568, n_569, n_570, n_571, n_572, n_573, n_574, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595;
  wire n_596, n_599, n_600, n_601, n_602, n_603, n_604, n_605;
  wire n_606, n_607, n_610, n_611, n_612, n_613, n_614, n_615;
  wire n_616, n_617, n_618, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_632, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_643, n_644, n_645;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_654, n_655;
  wire n_656, n_657, n_658, n_659, n_660, n_661, n_662, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_694, n_695, n_698, n_699, n_700, n_701, n_702, n_703;
  wire n_704, n_705, n_706, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_731, n_732, n_733;
  wire n_734, n_735, n_736, n_737, n_738, n_739, n_742, n_743;
  wire n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_775, n_776, n_777, n_778, n_779, n_780, n_781;
  wire n_782, n_783, n_786, n_787, n_788, n_789, n_790, n_791;
  wire n_792, n_793, n_794, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_808, n_809, n_810, n_811;
  wire n_812, n_813, n_814, n_815, n_816, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_830, n_831;
  wire n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_841;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_860, n_863, n_864, n_865, n_866, n_867, n_868, n_869;
  wire n_870, n_871, n_874, n_875, n_876, n_877, n_878, n_879;
  wire n_880, n_881, n_882, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_896, n_897, n_898, n_899;
  wire n_900, n_901, n_902, n_903, n_904, n_907, n_908, n_909;
  wire n_910, n_911, n_912, n_913, n_914, n_915, n_918, n_919;
  wire n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937;
  wire n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947;
  wire n_948, n_951, n_952, n_953, n_954, n_955, n_956, n_957;
  wire n_958, n_959, n_962, n_963, n_964, n_965, n_966, n_967;
  wire n_968, n_969, n_970, n_973, n_974, n_975, n_976, n_977;
  wire n_978, n_979, n_980, n_981, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_995, n_996, n_997;
  wire n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1006, n_1007;
  wire n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1017;
  wire n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1036, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045;
  wire n_1046, n_1047, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055;
  wire n_1056, n_1057, n_1058, n_1061, n_1062, n_1063, n_1064, n_1065;
  wire n_1066, n_1067, n_1068, n_1069, n_1072, n_1073, n_1074, n_1075;
  wire n_1076, n_1077, n_1078, n_1079, n_1080, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1094, n_1095;
  wire n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1105;
  wire n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113;
  wire n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123;
  wire n_1124, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133;
  wire n_1134, n_1135, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143;
  wire n_1144, n_1145, n_1146, n_1149, n_1150, n_1151, n_1152, n_1153;
  wire n_1154, n_1155, n_1156, n_1157, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1182, n_1183;
  wire n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1193;
  wire n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231;
  wire n_1232, n_1233, n_1234, n_1237, n_1238, n_1239, n_1240, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1259, n_1260, n_1261;
  wire n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1281;
  wire n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1300, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319;
  wire n_1320, n_1321, n_1322, n_1325, n_1326, n_1327, n_1328, n_1329;
  wire n_1330, n_1331, n_1332, n_1333, n_1336, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1342, n_1343, n_1344, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1358, n_1359;
  wire n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1369;
  wire n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1388, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398;
  not g1 (n_3, \b[0] );
  and g2 (n386, \a[0] , n_3);
  not g3 (n_4, \a[0] );
  and g4 (n387, n_4, \b[0] );
  or g5 (\f[0] , n386, n387);
  and g6 (n389, \a[0] , \b[0] );
  not g7 (n_7, \a[1] );
  not g8 (n_8, \b[1] );
  and g9 (n390, n_7, n_8);
  and g10 (n391, \a[1] , \b[1] );
  not g11 (n_9, n390);
  not g12 (n_10, n391);
  and g13 (n392, n_9, n_10);
  not g14 (n_11, n392);
  and g15 (n393, n389, n_11);
  not g16 (n_12, n389);
  and g17 (n394, n_12, n392);
  or g18 (\f[1] , n393, n394);
  and g19 (n396, n389, n_9);
  not g20 (n_13, n396);
  and g21 (n397, n_10, n_13);
  not g22 (n_16, \a[2] );
  not g23 (n_17, \b[2] );
  and g24 (n398, n_16, n_17);
  and g25 (n399, \a[2] , \b[2] );
  not g26 (n_18, n398);
  not g27 (n_19, n399);
  and g28 (n400, n_18, n_19);
  not g29 (n_20, n400);
  and g30 (n401, n397, n_20);
  not g31 (n_21, n397);
  and g32 (n402, n_21, n400);
  not g33 (n_22, n401);
  not g34 (n_23, n402);
  and g35 (\f[2] , n_22, n_23);
  and g36 (n404, n_21, n_18);
  not g37 (n_24, n404);
  and g38 (n405, n_19, n_24);
  not g39 (n_27, \a[3] );
  not g40 (n_28, \b[3] );
  and g41 (n406, n_27, n_28);
  and g42 (n407, \a[3] , \b[3] );
  not g43 (n_29, n406);
  not g44 (n_30, n407);
  and g45 (n408, n_29, n_30);
  not g46 (n_31, n408);
  and g47 (n409, n405, n_31);
  not g48 (n_32, n405);
  and g49 (n410, n_32, n408);
  not g50 (n_33, n409);
  not g51 (n_34, n410);
  and g52 (\f[3] , n_33, n_34);
  and g53 (n412, n_32, n_29);
  not g54 (n_35, n412);
  and g55 (n413, n_30, n_35);
  not g56 (n_38, \a[4] );
  not g57 (n_39, \b[4] );
  and g58 (n414, n_38, n_39);
  and g59 (n415, \a[4] , \b[4] );
  not g60 (n_40, n414);
  not g61 (n_41, n415);
  and g62 (n416, n_40, n_41);
  not g63 (n_42, n416);
  and g64 (n417, n413, n_42);
  not g65 (n_43, n413);
  and g66 (n418, n_43, n416);
  not g67 (n_44, n417);
  not g68 (n_45, n418);
  and g69 (\f[4] , n_44, n_45);
  and g70 (n420, n_43, n_40);
  not g71 (n_46, n420);
  and g72 (n421, n_41, n_46);
  not g73 (n_49, \a[5] );
  not g74 (n_50, \b[5] );
  and g75 (n422, n_49, n_50);
  and g76 (n423, \a[5] , \b[5] );
  not g77 (n_51, n422);
  not g78 (n_52, n423);
  and g79 (n424, n_51, n_52);
  not g80 (n_53, n424);
  and g81 (n425, n421, n_53);
  not g82 (n_54, n421);
  and g83 (n426, n_54, n424);
  not g84 (n_55, n425);
  not g85 (n_56, n426);
  and g86 (\f[5] , n_55, n_56);
  and g87 (n428, n_54, n_51);
  not g88 (n_57, n428);
  and g89 (n429, n_52, n_57);
  not g90 (n_60, \a[6] );
  not g91 (n_61, \b[6] );
  and g92 (n430, n_60, n_61);
  and g93 (n431, \a[6] , \b[6] );
  not g94 (n_62, n430);
  not g95 (n_63, n431);
  and g96 (n432, n_62, n_63);
  not g97 (n_64, n432);
  and g98 (n433, n429, n_64);
  not g99 (n_65, n429);
  and g100 (n434, n_65, n432);
  not g101 (n_66, n433);
  not g102 (n_67, n434);
  and g103 (\f[6] , n_66, n_67);
  and g104 (n436, n_65, n_62);
  not g105 (n_68, n436);
  and g106 (n437, n_63, n_68);
  not g107 (n_71, \a[7] );
  not g108 (n_72, \b[7] );
  and g109 (n438, n_71, n_72);
  and g110 (n439, \a[7] , \b[7] );
  not g111 (n_73, n438);
  not g112 (n_74, n439);
  and g113 (n440, n_73, n_74);
  not g114 (n_75, n440);
  and g115 (n441, n437, n_75);
  not g116 (n_76, n437);
  and g117 (n442, n_76, n440);
  not g118 (n_77, n441);
  not g119 (n_78, n442);
  and g120 (\f[7] , n_77, n_78);
  and g121 (n444, n_76, n_73);
  not g122 (n_79, n444);
  and g123 (n445, n_74, n_79);
  not g124 (n_82, \a[8] );
  not g125 (n_83, \b[8] );
  and g126 (n446, n_82, n_83);
  and g127 (n447, \a[8] , \b[8] );
  not g128 (n_84, n446);
  not g129 (n_85, n447);
  and g130 (n448, n_84, n_85);
  not g131 (n_86, n448);
  and g132 (n449, n445, n_86);
  not g133 (n_87, n445);
  and g134 (n450, n_87, n448);
  not g135 (n_88, n449);
  not g136 (n_89, n450);
  and g137 (\f[8] , n_88, n_89);
  and g138 (n452, n_87, n_84);
  not g139 (n_90, n452);
  and g140 (n453, n_85, n_90);
  not g141 (n_93, \a[9] );
  not g142 (n_94, \b[9] );
  and g143 (n454, n_93, n_94);
  and g144 (n455, \a[9] , \b[9] );
  not g145 (n_95, n454);
  not g146 (n_96, n455);
  and g147 (n456, n_95, n_96);
  not g148 (n_97, n456);
  and g149 (n457, n453, n_97);
  not g150 (n_98, n453);
  and g151 (n458, n_98, n456);
  not g152 (n_99, n457);
  not g153 (n_100, n458);
  and g154 (\f[9] , n_99, n_100);
  and g155 (n460, n_98, n_95);
  not g156 (n_101, n460);
  and g157 (n461, n_96, n_101);
  not g158 (n_104, \a[10] );
  not g159 (n_105, \b[10] );
  and g160 (n462, n_104, n_105);
  and g161 (n463, \a[10] , \b[10] );
  not g162 (n_106, n462);
  not g163 (n_107, n463);
  and g164 (n464, n_106, n_107);
  not g165 (n_108, n464);
  and g166 (n465, n461, n_108);
  not g167 (n_109, n461);
  and g168 (n466, n_109, n464);
  not g169 (n_110, n465);
  not g170 (n_111, n466);
  and g171 (\f[10] , n_110, n_111);
  and g172 (n468, n_109, n_106);
  not g173 (n_112, n468);
  and g174 (n469, n_107, n_112);
  not g175 (n_115, \a[11] );
  not g176 (n_116, \b[11] );
  and g177 (n470, n_115, n_116);
  and g178 (n471, \a[11] , \b[11] );
  not g179 (n_117, n470);
  not g180 (n_118, n471);
  and g181 (n472, n_117, n_118);
  not g182 (n_119, n472);
  and g183 (n473, n469, n_119);
  not g184 (n_120, n469);
  and g185 (n474, n_120, n472);
  not g186 (n_121, n473);
  not g187 (n_122, n474);
  and g188 (\f[11] , n_121, n_122);
  and g189 (n476, n_120, n_117);
  not g190 (n_123, n476);
  and g191 (n477, n_118, n_123);
  not g192 (n_126, \a[12] );
  not g193 (n_127, \b[12] );
  and g194 (n478, n_126, n_127);
  and g195 (n479, \a[12] , \b[12] );
  not g196 (n_128, n478);
  not g197 (n_129, n479);
  and g198 (n480, n_128, n_129);
  not g199 (n_130, n480);
  and g200 (n481, n477, n_130);
  not g201 (n_131, n477);
  and g202 (n482, n_131, n480);
  not g203 (n_132, n481);
  not g204 (n_133, n482);
  and g205 (\f[12] , n_132, n_133);
  and g206 (n484, n_131, n_128);
  not g207 (n_134, n484);
  and g208 (n485, n_129, n_134);
  not g209 (n_137, \a[13] );
  not g210 (n_138, \b[13] );
  and g211 (n486, n_137, n_138);
  and g212 (n487, \a[13] , \b[13] );
  not g213 (n_139, n486);
  not g214 (n_140, n487);
  and g215 (n488, n_139, n_140);
  not g216 (n_141, n488);
  and g217 (n489, n485, n_141);
  not g218 (n_142, n485);
  and g219 (n490, n_142, n488);
  not g220 (n_143, n489);
  not g221 (n_144, n490);
  and g222 (\f[13] , n_143, n_144);
  and g223 (n492, n_142, n_139);
  not g224 (n_145, n492);
  and g225 (n493, n_140, n_145);
  not g226 (n_148, \a[14] );
  not g227 (n_149, \b[14] );
  and g228 (n494, n_148, n_149);
  and g229 (n495, \a[14] , \b[14] );
  not g230 (n_150, n494);
  not g231 (n_151, n495);
  and g232 (n496, n_150, n_151);
  not g233 (n_152, n496);
  and g234 (n497, n493, n_152);
  not g235 (n_153, n493);
  and g236 (n498, n_153, n496);
  not g237 (n_154, n497);
  not g238 (n_155, n498);
  and g239 (\f[14] , n_154, n_155);
  and g240 (n500, n_153, n_150);
  not g241 (n_156, n500);
  and g242 (n501, n_151, n_156);
  not g243 (n_159, \a[15] );
  not g244 (n_160, \b[15] );
  and g245 (n502, n_159, n_160);
  and g246 (n503, \a[15] , \b[15] );
  not g247 (n_161, n502);
  not g248 (n_162, n503);
  and g249 (n504, n_161, n_162);
  not g250 (n_163, n504);
  and g251 (n505, n501, n_163);
  not g252 (n_164, n501);
  and g253 (n506, n_164, n504);
  not g254 (n_165, n505);
  not g255 (n_166, n506);
  and g256 (\f[15] , n_165, n_166);
  and g257 (n508, n_164, n_161);
  not g258 (n_167, n508);
  and g259 (n509, n_162, n_167);
  not g260 (n_170, \a[16] );
  not g261 (n_171, \b[16] );
  and g262 (n510, n_170, n_171);
  and g263 (n511, \a[16] , \b[16] );
  not g264 (n_172, n510);
  not g265 (n_173, n511);
  and g266 (n512, n_172, n_173);
  not g267 (n_174, n512);
  and g268 (n513, n509, n_174);
  not g269 (n_175, n509);
  and g270 (n514, n_175, n512);
  not g271 (n_176, n513);
  not g272 (n_177, n514);
  and g273 (\f[16] , n_176, n_177);
  and g274 (n516, n_175, n_172);
  not g275 (n_178, n516);
  and g276 (n517, n_173, n_178);
  not g277 (n_181, \a[17] );
  not g278 (n_182, \b[17] );
  and g279 (n518, n_181, n_182);
  and g280 (n519, \a[17] , \b[17] );
  not g281 (n_183, n518);
  not g282 (n_184, n519);
  and g283 (n520, n_183, n_184);
  not g284 (n_185, n520);
  and g285 (n521, n517, n_185);
  not g286 (n_186, n517);
  and g287 (n522, n_186, n520);
  not g288 (n_187, n521);
  not g289 (n_188, n522);
  and g290 (\f[17] , n_187, n_188);
  and g291 (n524, n_186, n_183);
  not g292 (n_189, n524);
  and g293 (n525, n_184, n_189);
  not g294 (n_192, \a[18] );
  not g295 (n_193, \b[18] );
  and g296 (n526, n_192, n_193);
  and g297 (n527, \a[18] , \b[18] );
  not g298 (n_194, n526);
  not g299 (n_195, n527);
  and g300 (n528, n_194, n_195);
  not g301 (n_196, n528);
  and g302 (n529, n525, n_196);
  not g303 (n_197, n525);
  and g304 (n530, n_197, n528);
  not g305 (n_198, n529);
  not g306 (n_199, n530);
  and g307 (\f[18] , n_198, n_199);
  and g308 (n532, n_197, n_194);
  not g309 (n_200, n532);
  and g310 (n533, n_195, n_200);
  not g311 (n_203, \a[19] );
  not g312 (n_204, \b[19] );
  and g313 (n534, n_203, n_204);
  and g314 (n535, \a[19] , \b[19] );
  not g315 (n_205, n534);
  not g316 (n_206, n535);
  and g317 (n536, n_205, n_206);
  not g318 (n_207, n536);
  and g319 (n537, n533, n_207);
  not g320 (n_208, n533);
  and g321 (n538, n_208, n536);
  not g322 (n_209, n537);
  not g323 (n_210, n538);
  and g324 (\f[19] , n_209, n_210);
  and g325 (n540, n_208, n_205);
  not g326 (n_211, n540);
  and g327 (n541, n_206, n_211);
  not g328 (n_214, \a[20] );
  not g329 (n_215, \b[20] );
  and g330 (n542, n_214, n_215);
  and g331 (n543, \a[20] , \b[20] );
  not g332 (n_216, n542);
  not g333 (n_217, n543);
  and g334 (n544, n_216, n_217);
  not g335 (n_218, n544);
  and g336 (n545, n541, n_218);
  not g337 (n_219, n541);
  and g338 (n546, n_219, n544);
  not g339 (n_220, n545);
  not g340 (n_221, n546);
  and g341 (\f[20] , n_220, n_221);
  and g342 (n548, n_219, n_216);
  not g343 (n_222, n548);
  and g344 (n549, n_217, n_222);
  not g345 (n_225, \a[21] );
  not g346 (n_226, \b[21] );
  and g347 (n550, n_225, n_226);
  and g348 (n551, \a[21] , \b[21] );
  not g349 (n_227, n550);
  not g350 (n_228, n551);
  and g351 (n552, n_227, n_228);
  not g352 (n_229, n552);
  and g353 (n553, n549, n_229);
  not g354 (n_230, n549);
  and g355 (n554, n_230, n552);
  not g356 (n_231, n553);
  not g357 (n_232, n554);
  and g358 (\f[21] , n_231, n_232);
  and g359 (n556, n_230, n_227);
  not g360 (n_233, n556);
  and g361 (n557, n_228, n_233);
  not g362 (n_236, \a[22] );
  not g363 (n_237, \b[22] );
  and g364 (n558, n_236, n_237);
  and g365 (n559, \a[22] , \b[22] );
  not g366 (n_238, n558);
  not g367 (n_239, n559);
  and g368 (n560, n_238, n_239);
  not g369 (n_240, n560);
  and g370 (n561, n557, n_240);
  not g371 (n_241, n557);
  and g372 (n562, n_241, n560);
  not g373 (n_242, n561);
  not g374 (n_243, n562);
  and g375 (\f[22] , n_242, n_243);
  and g376 (n564, n_241, n_238);
  not g377 (n_244, n564);
  and g378 (n565, n_239, n_244);
  not g379 (n_247, \a[23] );
  not g380 (n_248, \b[23] );
  and g381 (n566, n_247, n_248);
  and g382 (n567, \a[23] , \b[23] );
  not g383 (n_249, n566);
  not g384 (n_250, n567);
  and g385 (n568, n_249, n_250);
  not g386 (n_251, n568);
  and g387 (n569, n565, n_251);
  not g388 (n_252, n565);
  and g389 (n570, n_252, n568);
  not g390 (n_253, n569);
  not g391 (n_254, n570);
  and g392 (\f[23] , n_253, n_254);
  and g393 (n572, n_252, n_249);
  not g394 (n_255, n572);
  and g395 (n573, n_250, n_255);
  not g396 (n_258, \a[24] );
  not g397 (n_259, \b[24] );
  and g398 (n574, n_258, n_259);
  and g399 (n575, \a[24] , \b[24] );
  not g400 (n_260, n574);
  not g401 (n_261, n575);
  and g402 (n576, n_260, n_261);
  not g403 (n_262, n576);
  and g404 (n577, n573, n_262);
  not g405 (n_263, n573);
  and g406 (n578, n_263, n576);
  not g407 (n_264, n577);
  not g408 (n_265, n578);
  and g409 (\f[24] , n_264, n_265);
  and g410 (n580, n_263, n_260);
  not g411 (n_266, n580);
  and g412 (n581, n_261, n_266);
  not g413 (n_269, \a[25] );
  not g414 (n_270, \b[25] );
  and g415 (n582, n_269, n_270);
  and g416 (n583, \a[25] , \b[25] );
  not g417 (n_271, n582);
  not g418 (n_272, n583);
  and g419 (n584, n_271, n_272);
  not g420 (n_273, n584);
  and g421 (n585, n581, n_273);
  not g422 (n_274, n581);
  and g423 (n586, n_274, n584);
  not g424 (n_275, n585);
  not g425 (n_276, n586);
  and g426 (\f[25] , n_275, n_276);
  and g427 (n588, n_274, n_271);
  not g428 (n_277, n588);
  and g429 (n589, n_272, n_277);
  not g430 (n_280, \a[26] );
  not g431 (n_281, \b[26] );
  and g432 (n590, n_280, n_281);
  and g433 (n591, \a[26] , \b[26] );
  not g434 (n_282, n590);
  not g435 (n_283, n591);
  and g436 (n592, n_282, n_283);
  not g437 (n_284, n592);
  and g438 (n593, n589, n_284);
  not g439 (n_285, n589);
  and g440 (n594, n_285, n592);
  not g441 (n_286, n593);
  not g442 (n_287, n594);
  and g443 (\f[26] , n_286, n_287);
  and g444 (n596, n_285, n_282);
  not g445 (n_288, n596);
  and g446 (n597, n_283, n_288);
  not g447 (n_291, \a[27] );
  not g448 (n_292, \b[27] );
  and g449 (n598, n_291, n_292);
  and g450 (n599, \a[27] , \b[27] );
  not g451 (n_293, n598);
  not g452 (n_294, n599);
  and g453 (n600, n_293, n_294);
  not g454 (n_295, n600);
  and g455 (n601, n597, n_295);
  not g456 (n_296, n597);
  and g457 (n602, n_296, n600);
  not g458 (n_297, n601);
  not g459 (n_298, n602);
  and g460 (\f[27] , n_297, n_298);
  and g461 (n604, n_296, n_293);
  not g462 (n_299, n604);
  and g463 (n605, n_294, n_299);
  not g464 (n_302, \a[28] );
  not g465 (n_303, \b[28] );
  and g466 (n606, n_302, n_303);
  and g467 (n607, \a[28] , \b[28] );
  not g468 (n_304, n606);
  not g469 (n_305, n607);
  and g470 (n608, n_304, n_305);
  not g471 (n_306, n608);
  and g472 (n609, n605, n_306);
  not g473 (n_307, n605);
  and g474 (n610, n_307, n608);
  not g475 (n_308, n609);
  not g476 (n_309, n610);
  and g477 (\f[28] , n_308, n_309);
  and g478 (n612, n_307, n_304);
  not g479 (n_310, n612);
  and g480 (n613, n_305, n_310);
  not g481 (n_313, \a[29] );
  not g482 (n_314, \b[29] );
  and g483 (n614, n_313, n_314);
  and g484 (n615, \a[29] , \b[29] );
  not g485 (n_315, n614);
  not g486 (n_316, n615);
  and g487 (n616, n_315, n_316);
  not g488 (n_317, n616);
  and g489 (n617, n613, n_317);
  not g490 (n_318, n613);
  and g491 (n618, n_318, n616);
  not g492 (n_319, n617);
  not g493 (n_320, n618);
  and g494 (\f[29] , n_319, n_320);
  and g495 (n620, n_318, n_315);
  not g496 (n_321, n620);
  and g497 (n621, n_316, n_321);
  not g498 (n_324, \a[30] );
  not g499 (n_325, \b[30] );
  and g500 (n622, n_324, n_325);
  and g501 (n623, \a[30] , \b[30] );
  not g502 (n_326, n622);
  not g503 (n_327, n623);
  and g504 (n624, n_326, n_327);
  not g505 (n_328, n624);
  and g506 (n625, n621, n_328);
  not g507 (n_329, n621);
  and g508 (n626, n_329, n624);
  not g509 (n_330, n625);
  not g510 (n_331, n626);
  and g511 (\f[30] , n_330, n_331);
  and g512 (n628, n_329, n_326);
  not g513 (n_332, n628);
  and g514 (n629, n_327, n_332);
  not g515 (n_335, \a[31] );
  not g516 (n_336, \b[31] );
  and g517 (n630, n_335, n_336);
  and g518 (n631, \a[31] , \b[31] );
  not g519 (n_337, n630);
  not g520 (n_338, n631);
  and g521 (n632, n_337, n_338);
  not g522 (n_339, n632);
  and g523 (n633, n629, n_339);
  not g524 (n_340, n629);
  and g525 (n634, n_340, n632);
  not g526 (n_341, n633);
  not g527 (n_342, n634);
  and g528 (\f[31] , n_341, n_342);
  and g529 (n636, n_340, n_337);
  not g530 (n_343, n636);
  and g531 (n637, n_338, n_343);
  not g532 (n_346, \a[32] );
  not g533 (n_347, \b[32] );
  and g534 (n638, n_346, n_347);
  and g535 (n639, \a[32] , \b[32] );
  not g536 (n_348, n638);
  not g537 (n_349, n639);
  and g538 (n640, n_348, n_349);
  not g539 (n_350, n640);
  and g540 (n641, n637, n_350);
  not g541 (n_351, n637);
  and g542 (n642, n_351, n640);
  not g543 (n_352, n641);
  not g544 (n_353, n642);
  and g545 (\f[32] , n_352, n_353);
  and g546 (n644, n_351, n_348);
  not g547 (n_354, n644);
  and g548 (n645, n_349, n_354);
  not g549 (n_357, \a[33] );
  not g550 (n_358, \b[33] );
  and g551 (n646, n_357, n_358);
  and g552 (n647, \a[33] , \b[33] );
  not g553 (n_359, n646);
  not g554 (n_360, n647);
  and g555 (n648, n_359, n_360);
  not g556 (n_361, n648);
  and g557 (n649, n645, n_361);
  not g558 (n_362, n645);
  and g559 (n650, n_362, n648);
  not g560 (n_363, n649);
  not g561 (n_364, n650);
  and g562 (\f[33] , n_363, n_364);
  and g563 (n652, n_362, n_359);
  not g564 (n_365, n652);
  and g565 (n653, n_360, n_365);
  not g566 (n_368, \a[34] );
  not g567 (n_369, \b[34] );
  and g568 (n654, n_368, n_369);
  and g569 (n655, \a[34] , \b[34] );
  not g570 (n_370, n654);
  not g571 (n_371, n655);
  and g572 (n656, n_370, n_371);
  not g573 (n_372, n656);
  and g574 (n657, n653, n_372);
  not g575 (n_373, n653);
  and g576 (n658, n_373, n656);
  not g577 (n_374, n657);
  not g578 (n_375, n658);
  and g579 (\f[34] , n_374, n_375);
  and g580 (n660, n_373, n_370);
  not g581 (n_376, n660);
  and g582 (n661, n_371, n_376);
  not g583 (n_379, \a[35] );
  not g584 (n_380, \b[35] );
  and g585 (n662, n_379, n_380);
  and g586 (n663, \a[35] , \b[35] );
  not g587 (n_381, n662);
  not g588 (n_382, n663);
  and g589 (n664, n_381, n_382);
  not g590 (n_383, n664);
  and g591 (n665, n661, n_383);
  not g592 (n_384, n661);
  and g593 (n666, n_384, n664);
  not g594 (n_385, n665);
  not g595 (n_386, n666);
  and g596 (\f[35] , n_385, n_386);
  and g597 (n668, n_384, n_381);
  not g598 (n_387, n668);
  and g599 (n669, n_382, n_387);
  not g600 (n_390, \a[36] );
  not g601 (n_391, \b[36] );
  and g602 (n670, n_390, n_391);
  and g603 (n671, \a[36] , \b[36] );
  not g604 (n_392, n670);
  not g605 (n_393, n671);
  and g606 (n672, n_392, n_393);
  not g607 (n_394, n672);
  and g608 (n673, n669, n_394);
  not g609 (n_395, n669);
  and g610 (n674, n_395, n672);
  not g611 (n_396, n673);
  not g612 (n_397, n674);
  and g613 (\f[36] , n_396, n_397);
  and g614 (n676, n_395, n_392);
  not g615 (n_398, n676);
  and g616 (n677, n_393, n_398);
  not g617 (n_401, \a[37] );
  not g618 (n_402, \b[37] );
  and g619 (n678, n_401, n_402);
  and g620 (n679, \a[37] , \b[37] );
  not g621 (n_403, n678);
  not g622 (n_404, n679);
  and g623 (n680, n_403, n_404);
  not g624 (n_405, n680);
  and g625 (n681, n677, n_405);
  not g626 (n_406, n677);
  and g627 (n682, n_406, n680);
  not g628 (n_407, n681);
  not g629 (n_408, n682);
  and g630 (\f[37] , n_407, n_408);
  and g631 (n684, n_406, n_403);
  not g632 (n_409, n684);
  and g633 (n685, n_404, n_409);
  not g634 (n_412, \a[38] );
  not g635 (n_413, \b[38] );
  and g636 (n686, n_412, n_413);
  and g637 (n687, \a[38] , \b[38] );
  not g638 (n_414, n686);
  not g639 (n_415, n687);
  and g640 (n688, n_414, n_415);
  not g641 (n_416, n688);
  and g642 (n689, n685, n_416);
  not g643 (n_417, n685);
  and g644 (n690, n_417, n688);
  not g645 (n_418, n689);
  not g646 (n_419, n690);
  and g647 (\f[38] , n_418, n_419);
  and g648 (n692, n_417, n_414);
  not g649 (n_420, n692);
  and g650 (n693, n_415, n_420);
  not g651 (n_423, \a[39] );
  not g652 (n_424, \b[39] );
  and g653 (n694, n_423, n_424);
  and g654 (n695, \a[39] , \b[39] );
  not g655 (n_425, n694);
  not g656 (n_426, n695);
  and g657 (n696, n_425, n_426);
  not g658 (n_427, n696);
  and g659 (n697, n693, n_427);
  not g660 (n_428, n693);
  and g661 (n698, n_428, n696);
  not g662 (n_429, n697);
  not g663 (n_430, n698);
  and g664 (\f[39] , n_429, n_430);
  and g665 (n700, n_428, n_425);
  not g666 (n_431, n700);
  and g667 (n701, n_426, n_431);
  not g668 (n_434, \a[40] );
  not g669 (n_435, \b[40] );
  and g670 (n702, n_434, n_435);
  and g671 (n703, \a[40] , \b[40] );
  not g672 (n_436, n702);
  not g673 (n_437, n703);
  and g674 (n704, n_436, n_437);
  not g675 (n_438, n704);
  and g676 (n705, n701, n_438);
  not g677 (n_439, n701);
  and g678 (n706, n_439, n704);
  not g679 (n_440, n705);
  not g680 (n_441, n706);
  and g681 (\f[40] , n_440, n_441);
  and g682 (n708, n_439, n_436);
  not g683 (n_442, n708);
  and g684 (n709, n_437, n_442);
  not g685 (n_445, \a[41] );
  not g686 (n_446, \b[41] );
  and g687 (n710, n_445, n_446);
  and g688 (n711, \a[41] , \b[41] );
  not g689 (n_447, n710);
  not g690 (n_448, n711);
  and g691 (n712, n_447, n_448);
  not g692 (n_449, n712);
  and g693 (n713, n709, n_449);
  not g694 (n_450, n709);
  and g695 (n714, n_450, n712);
  not g696 (n_451, n713);
  not g697 (n_452, n714);
  and g698 (\f[41] , n_451, n_452);
  and g699 (n716, n_450, n_447);
  not g700 (n_453, n716);
  and g701 (n717, n_448, n_453);
  not g702 (n_456, \a[42] );
  not g703 (n_457, \b[42] );
  and g704 (n718, n_456, n_457);
  and g705 (n719, \a[42] , \b[42] );
  not g706 (n_458, n718);
  not g707 (n_459, n719);
  and g708 (n720, n_458, n_459);
  not g709 (n_460, n720);
  and g710 (n721, n717, n_460);
  not g711 (n_461, n717);
  and g712 (n722, n_461, n720);
  not g713 (n_462, n721);
  not g714 (n_463, n722);
  and g715 (\f[42] , n_462, n_463);
  and g716 (n724, n_461, n_458);
  not g717 (n_464, n724);
  and g718 (n725, n_459, n_464);
  not g719 (n_467, \a[43] );
  not g720 (n_468, \b[43] );
  and g721 (n726, n_467, n_468);
  and g722 (n727, \a[43] , \b[43] );
  not g723 (n_469, n726);
  not g724 (n_470, n727);
  and g725 (n728, n_469, n_470);
  not g726 (n_471, n728);
  and g727 (n729, n725, n_471);
  not g728 (n_472, n725);
  and g729 (n730, n_472, n728);
  not g730 (n_473, n729);
  not g731 (n_474, n730);
  and g732 (\f[43] , n_473, n_474);
  and g733 (n732, n_472, n_469);
  not g734 (n_475, n732);
  and g735 (n733, n_470, n_475);
  not g736 (n_478, \a[44] );
  not g737 (n_479, \b[44] );
  and g738 (n734, n_478, n_479);
  and g739 (n735, \a[44] , \b[44] );
  not g740 (n_480, n734);
  not g741 (n_481, n735);
  and g742 (n736, n_480, n_481);
  not g743 (n_482, n736);
  and g744 (n737, n733, n_482);
  not g745 (n_483, n733);
  and g746 (n738, n_483, n736);
  not g747 (n_484, n737);
  not g748 (n_485, n738);
  and g749 (\f[44] , n_484, n_485);
  and g750 (n740, n_483, n_480);
  not g751 (n_486, n740);
  and g752 (n741, n_481, n_486);
  not g753 (n_489, \a[45] );
  not g754 (n_490, \b[45] );
  and g755 (n742, n_489, n_490);
  and g756 (n743, \a[45] , \b[45] );
  not g757 (n_491, n742);
  not g758 (n_492, n743);
  and g759 (n744, n_491, n_492);
  not g760 (n_493, n744);
  and g761 (n745, n741, n_493);
  not g762 (n_494, n741);
  and g763 (n746, n_494, n744);
  not g764 (n_495, n745);
  not g765 (n_496, n746);
  and g766 (\f[45] , n_495, n_496);
  and g767 (n748, n_494, n_491);
  not g768 (n_497, n748);
  and g769 (n749, n_492, n_497);
  not g770 (n_500, \a[46] );
  not g771 (n_501, \b[46] );
  and g772 (n750, n_500, n_501);
  and g773 (n751, \a[46] , \b[46] );
  not g774 (n_502, n750);
  not g775 (n_503, n751);
  and g776 (n752, n_502, n_503);
  not g777 (n_504, n752);
  and g778 (n753, n749, n_504);
  not g779 (n_505, n749);
  and g780 (n754, n_505, n752);
  not g781 (n_506, n753);
  not g782 (n_507, n754);
  and g783 (\f[46] , n_506, n_507);
  and g784 (n756, n_505, n_502);
  not g785 (n_508, n756);
  and g786 (n757, n_503, n_508);
  not g787 (n_511, \a[47] );
  not g788 (n_512, \b[47] );
  and g789 (n758, n_511, n_512);
  and g790 (n759, \a[47] , \b[47] );
  not g791 (n_513, n758);
  not g792 (n_514, n759);
  and g793 (n760, n_513, n_514);
  not g794 (n_515, n760);
  and g795 (n761, n757, n_515);
  not g796 (n_516, n757);
  and g797 (n762, n_516, n760);
  not g798 (n_517, n761);
  not g799 (n_518, n762);
  and g800 (\f[47] , n_517, n_518);
  and g801 (n764, n_516, n_513);
  not g802 (n_519, n764);
  and g803 (n765, n_514, n_519);
  not g804 (n_522, \a[48] );
  not g805 (n_523, \b[48] );
  and g806 (n766, n_522, n_523);
  and g807 (n767, \a[48] , \b[48] );
  not g808 (n_524, n766);
  not g809 (n_525, n767);
  and g810 (n768, n_524, n_525);
  not g811 (n_526, n768);
  and g812 (n769, n765, n_526);
  not g813 (n_527, n765);
  and g814 (n770, n_527, n768);
  not g815 (n_528, n769);
  not g816 (n_529, n770);
  and g817 (\f[48] , n_528, n_529);
  and g818 (n772, n_527, n_524);
  not g819 (n_530, n772);
  and g820 (n773, n_525, n_530);
  not g821 (n_533, \a[49] );
  not g822 (n_534, \b[49] );
  and g823 (n774, n_533, n_534);
  and g824 (n775, \a[49] , \b[49] );
  not g825 (n_535, n774);
  not g826 (n_536, n775);
  and g827 (n776, n_535, n_536);
  not g828 (n_537, n776);
  and g829 (n777, n773, n_537);
  not g830 (n_538, n773);
  and g831 (n778, n_538, n776);
  not g832 (n_539, n777);
  not g833 (n_540, n778);
  and g834 (\f[49] , n_539, n_540);
  and g835 (n780, n_538, n_535);
  not g836 (n_541, n780);
  and g837 (n781, n_536, n_541);
  not g838 (n_544, \a[50] );
  not g839 (n_545, \b[50] );
  and g840 (n782, n_544, n_545);
  and g841 (n783, \a[50] , \b[50] );
  not g842 (n_546, n782);
  not g843 (n_547, n783);
  and g844 (n784, n_546, n_547);
  not g845 (n_548, n784);
  and g846 (n785, n781, n_548);
  not g847 (n_549, n781);
  and g848 (n786, n_549, n784);
  not g849 (n_550, n785);
  not g850 (n_551, n786);
  and g851 (\f[50] , n_550, n_551);
  and g852 (n788, n_549, n_546);
  not g853 (n_552, n788);
  and g854 (n789, n_547, n_552);
  not g855 (n_555, \a[51] );
  not g856 (n_556, \b[51] );
  and g857 (n790, n_555, n_556);
  and g858 (n791, \a[51] , \b[51] );
  not g859 (n_557, n790);
  not g860 (n_558, n791);
  and g861 (n792, n_557, n_558);
  not g862 (n_559, n792);
  and g863 (n793, n789, n_559);
  not g864 (n_560, n789);
  and g865 (n794, n_560, n792);
  not g866 (n_561, n793);
  not g867 (n_562, n794);
  and g868 (\f[51] , n_561, n_562);
  and g869 (n796, n_560, n_557);
  not g870 (n_563, n796);
  and g871 (n797, n_558, n_563);
  not g872 (n_566, \a[52] );
  not g873 (n_567, \b[52] );
  and g874 (n798, n_566, n_567);
  and g875 (n799, \a[52] , \b[52] );
  not g876 (n_568, n798);
  not g877 (n_569, n799);
  and g878 (n800, n_568, n_569);
  not g879 (n_570, n800);
  and g880 (n801, n797, n_570);
  not g881 (n_571, n797);
  and g882 (n802, n_571, n800);
  not g883 (n_572, n801);
  not g884 (n_573, n802);
  and g885 (\f[52] , n_572, n_573);
  and g886 (n804, n_571, n_568);
  not g887 (n_574, n804);
  and g888 (n805, n_569, n_574);
  not g889 (n_577, \a[53] );
  not g890 (n_578, \b[53] );
  and g891 (n806, n_577, n_578);
  and g892 (n807, \a[53] , \b[53] );
  not g893 (n_579, n806);
  not g894 (n_580, n807);
  and g895 (n808, n_579, n_580);
  not g896 (n_581, n808);
  and g897 (n809, n805, n_581);
  not g898 (n_582, n805);
  and g899 (n810, n_582, n808);
  not g900 (n_583, n809);
  not g901 (n_584, n810);
  and g902 (\f[53] , n_583, n_584);
  and g903 (n812, n_582, n_579);
  not g904 (n_585, n812);
  and g905 (n813, n_580, n_585);
  not g906 (n_588, \a[54] );
  not g907 (n_589, \b[54] );
  and g908 (n814, n_588, n_589);
  and g909 (n815, \a[54] , \b[54] );
  not g910 (n_590, n814);
  not g911 (n_591, n815);
  and g912 (n816, n_590, n_591);
  not g913 (n_592, n816);
  and g914 (n817, n813, n_592);
  not g915 (n_593, n813);
  and g916 (n818, n_593, n816);
  not g917 (n_594, n817);
  not g918 (n_595, n818);
  and g919 (\f[54] , n_594, n_595);
  and g920 (n820, n_593, n_590);
  not g921 (n_596, n820);
  and g922 (n821, n_591, n_596);
  not g923 (n_599, \a[55] );
  not g924 (n_600, \b[55] );
  and g925 (n822, n_599, n_600);
  and g926 (n823, \a[55] , \b[55] );
  not g927 (n_601, n822);
  not g928 (n_602, n823);
  and g929 (n824, n_601, n_602);
  not g930 (n_603, n824);
  and g931 (n825, n821, n_603);
  not g932 (n_604, n821);
  and g933 (n826, n_604, n824);
  not g934 (n_605, n825);
  not g935 (n_606, n826);
  and g936 (\f[55] , n_605, n_606);
  and g937 (n828, n_604, n_601);
  not g938 (n_607, n828);
  and g939 (n829, n_602, n_607);
  not g940 (n_610, \a[56] );
  not g941 (n_611, \b[56] );
  and g942 (n830, n_610, n_611);
  and g943 (n831, \a[56] , \b[56] );
  not g944 (n_612, n830);
  not g945 (n_613, n831);
  and g946 (n832, n_612, n_613);
  not g947 (n_614, n832);
  and g948 (n833, n829, n_614);
  not g949 (n_615, n829);
  and g950 (n834, n_615, n832);
  not g951 (n_616, n833);
  not g952 (n_617, n834);
  and g953 (\f[56] , n_616, n_617);
  and g954 (n836, n_615, n_612);
  not g955 (n_618, n836);
  and g956 (n837, n_613, n_618);
  not g957 (n_621, \a[57] );
  not g958 (n_622, \b[57] );
  and g959 (n838, n_621, n_622);
  and g960 (n839, \a[57] , \b[57] );
  not g961 (n_623, n838);
  not g962 (n_624, n839);
  and g963 (n840, n_623, n_624);
  not g964 (n_625, n840);
  and g965 (n841, n837, n_625);
  not g966 (n_626, n837);
  and g967 (n842, n_626, n840);
  not g968 (n_627, n841);
  not g969 (n_628, n842);
  and g970 (\f[57] , n_627, n_628);
  and g971 (n844, n_626, n_623);
  not g972 (n_629, n844);
  and g973 (n845, n_624, n_629);
  not g974 (n_632, \a[58] );
  not g975 (n_633, \b[58] );
  and g976 (n846, n_632, n_633);
  and g977 (n847, \a[58] , \b[58] );
  not g978 (n_634, n846);
  not g979 (n_635, n847);
  and g980 (n848, n_634, n_635);
  not g981 (n_636, n848);
  and g982 (n849, n845, n_636);
  not g983 (n_637, n845);
  and g984 (n850, n_637, n848);
  not g985 (n_638, n849);
  not g986 (n_639, n850);
  and g987 (\f[58] , n_638, n_639);
  and g988 (n852, n_637, n_634);
  not g989 (n_640, n852);
  and g990 (n853, n_635, n_640);
  not g991 (n_643, \a[59] );
  not g992 (n_644, \b[59] );
  and g993 (n854, n_643, n_644);
  and g994 (n855, \a[59] , \b[59] );
  not g995 (n_645, n854);
  not g996 (n_646, n855);
  and g997 (n856, n_645, n_646);
  not g998 (n_647, n856);
  and g999 (n857, n853, n_647);
  not g1000 (n_648, n853);
  and g1001 (n858, n_648, n856);
  not g1002 (n_649, n857);
  not g1003 (n_650, n858);
  and g1004 (\f[59] , n_649, n_650);
  and g1005 (n860, n_648, n_645);
  not g1006 (n_651, n860);
  and g1007 (n861, n_646, n_651);
  not g1008 (n_654, \a[60] );
  not g1009 (n_655, \b[60] );
  and g1010 (n862, n_654, n_655);
  and g1011 (n863, \a[60] , \b[60] );
  not g1012 (n_656, n862);
  not g1013 (n_657, n863);
  and g1014 (n864, n_656, n_657);
  not g1015 (n_658, n864);
  and g1016 (n865, n861, n_658);
  not g1017 (n_659, n861);
  and g1018 (n866, n_659, n864);
  not g1019 (n_660, n865);
  not g1020 (n_661, n866);
  and g1021 (\f[60] , n_660, n_661);
  and g1022 (n868, n_659, n_656);
  not g1023 (n_662, n868);
  and g1024 (n869, n_657, n_662);
  not g1025 (n_665, \a[61] );
  not g1026 (n_666, \b[61] );
  and g1027 (n870, n_665, n_666);
  and g1028 (n871, \a[61] , \b[61] );
  not g1029 (n_667, n870);
  not g1030 (n_668, n871);
  and g1031 (n872, n_667, n_668);
  not g1032 (n_669, n872);
  and g1033 (n873, n869, n_669);
  not g1034 (n_670, n869);
  and g1035 (n874, n_670, n872);
  not g1036 (n_671, n873);
  not g1037 (n_672, n874);
  and g1038 (\f[61] , n_671, n_672);
  and g1039 (n876, n_670, n_667);
  not g1040 (n_673, n876);
  and g1041 (n877, n_668, n_673);
  not g1042 (n_676, \a[62] );
  not g1043 (n_677, \b[62] );
  and g1044 (n878, n_676, n_677);
  and g1045 (n879, \a[62] , \b[62] );
  not g1046 (n_678, n878);
  not g1047 (n_679, n879);
  and g1048 (n880, n_678, n_679);
  not g1049 (n_680, n880);
  and g1050 (n881, n877, n_680);
  not g1051 (n_681, n877);
  and g1052 (n882, n_681, n880);
  not g1053 (n_682, n881);
  not g1054 (n_683, n882);
  and g1055 (\f[62] , n_682, n_683);
  and g1056 (n884, n_681, n_678);
  not g1057 (n_684, n884);
  and g1058 (n885, n_679, n_684);
  not g1059 (n_687, \a[63] );
  not g1060 (n_688, \b[63] );
  and g1061 (n886, n_687, n_688);
  and g1062 (n887, \a[63] , \b[63] );
  not g1063 (n_689, n886);
  not g1064 (n_690, n887);
  and g1065 (n888, n_689, n_690);
  not g1066 (n_691, n888);
  and g1067 (n889, n885, n_691);
  not g1068 (n_692, n885);
  and g1069 (n890, n_692, n888);
  not g1070 (n_693, n889);
  not g1071 (n_694, n890);
  and g1072 (\f[63] , n_693, n_694);
  and g1073 (n892, n_692, n_689);
  not g1074 (n_695, n892);
  and g1075 (n893, n_690, n_695);
  not g1076 (n_698, \a[64] );
  not g1077 (n_699, \b[64] );
  and g1078 (n894, n_698, n_699);
  and g1079 (n895, \a[64] , \b[64] );
  not g1080 (n_700, n894);
  not g1081 (n_701, n895);
  and g1082 (n896, n_700, n_701);
  not g1083 (n_702, n896);
  and g1084 (n897, n893, n_702);
  not g1085 (n_703, n893);
  and g1086 (n898, n_703, n896);
  not g1087 (n_704, n897);
  not g1088 (n_705, n898);
  and g1089 (\f[64] , n_704, n_705);
  and g1090 (n900, n_703, n_700);
  not g1091 (n_706, n900);
  and g1092 (n901, n_701, n_706);
  not g1093 (n_709, \a[65] );
  not g1094 (n_710, \b[65] );
  and g1095 (n902, n_709, n_710);
  and g1096 (n903, \a[65] , \b[65] );
  not g1097 (n_711, n902);
  not g1098 (n_712, n903);
  and g1099 (n904, n_711, n_712);
  not g1100 (n_713, n904);
  and g1101 (n905, n901, n_713);
  not g1102 (n_714, n901);
  and g1103 (n906, n_714, n904);
  not g1104 (n_715, n905);
  not g1105 (n_716, n906);
  and g1106 (\f[65] , n_715, n_716);
  and g1107 (n908, n_714, n_711);
  not g1108 (n_717, n908);
  and g1109 (n909, n_712, n_717);
  not g1110 (n_720, \a[66] );
  not g1111 (n_721, \b[66] );
  and g1112 (n910, n_720, n_721);
  and g1113 (n911, \a[66] , \b[66] );
  not g1114 (n_722, n910);
  not g1115 (n_723, n911);
  and g1116 (n912, n_722, n_723);
  not g1117 (n_724, n912);
  and g1118 (n913, n909, n_724);
  not g1119 (n_725, n909);
  and g1120 (n914, n_725, n912);
  not g1121 (n_726, n913);
  not g1122 (n_727, n914);
  and g1123 (\f[66] , n_726, n_727);
  and g1124 (n916, n_725, n_722);
  not g1125 (n_728, n916);
  and g1126 (n917, n_723, n_728);
  not g1127 (n_731, \a[67] );
  not g1128 (n_732, \b[67] );
  and g1129 (n918, n_731, n_732);
  and g1130 (n919, \a[67] , \b[67] );
  not g1131 (n_733, n918);
  not g1132 (n_734, n919);
  and g1133 (n920, n_733, n_734);
  not g1134 (n_735, n920);
  and g1135 (n921, n917, n_735);
  not g1136 (n_736, n917);
  and g1137 (n922, n_736, n920);
  not g1138 (n_737, n921);
  not g1139 (n_738, n922);
  and g1140 (\f[67] , n_737, n_738);
  and g1141 (n924, n_736, n_733);
  not g1142 (n_739, n924);
  and g1143 (n925, n_734, n_739);
  not g1144 (n_742, \a[68] );
  not g1145 (n_743, \b[68] );
  and g1146 (n926, n_742, n_743);
  and g1147 (n927, \a[68] , \b[68] );
  not g1148 (n_744, n926);
  not g1149 (n_745, n927);
  and g1150 (n928, n_744, n_745);
  not g1151 (n_746, n928);
  and g1152 (n929, n925, n_746);
  not g1153 (n_747, n925);
  and g1154 (n930, n_747, n928);
  not g1155 (n_748, n929);
  not g1156 (n_749, n930);
  and g1157 (\f[68] , n_748, n_749);
  and g1158 (n932, n_747, n_744);
  not g1159 (n_750, n932);
  and g1160 (n933, n_745, n_750);
  not g1161 (n_753, \a[69] );
  not g1162 (n_754, \b[69] );
  and g1163 (n934, n_753, n_754);
  and g1164 (n935, \a[69] , \b[69] );
  not g1165 (n_755, n934);
  not g1166 (n_756, n935);
  and g1167 (n936, n_755, n_756);
  not g1168 (n_757, n936);
  and g1169 (n937, n933, n_757);
  not g1170 (n_758, n933);
  and g1171 (n938, n_758, n936);
  not g1172 (n_759, n937);
  not g1173 (n_760, n938);
  and g1174 (\f[69] , n_759, n_760);
  and g1175 (n940, n_758, n_755);
  not g1176 (n_761, n940);
  and g1177 (n941, n_756, n_761);
  not g1178 (n_764, \a[70] );
  not g1179 (n_765, \b[70] );
  and g1180 (n942, n_764, n_765);
  and g1181 (n943, \a[70] , \b[70] );
  not g1182 (n_766, n942);
  not g1183 (n_767, n943);
  and g1184 (n944, n_766, n_767);
  not g1185 (n_768, n944);
  and g1186 (n945, n941, n_768);
  not g1187 (n_769, n941);
  and g1188 (n946, n_769, n944);
  not g1189 (n_770, n945);
  not g1190 (n_771, n946);
  and g1191 (\f[70] , n_770, n_771);
  and g1192 (n948, n_769, n_766);
  not g1193 (n_772, n948);
  and g1194 (n949, n_767, n_772);
  not g1195 (n_775, \a[71] );
  not g1196 (n_776, \b[71] );
  and g1197 (n950, n_775, n_776);
  and g1198 (n951, \a[71] , \b[71] );
  not g1199 (n_777, n950);
  not g1200 (n_778, n951);
  and g1201 (n952, n_777, n_778);
  not g1202 (n_779, n952);
  and g1203 (n953, n949, n_779);
  not g1204 (n_780, n949);
  and g1205 (n954, n_780, n952);
  not g1206 (n_781, n953);
  not g1207 (n_782, n954);
  and g1208 (\f[71] , n_781, n_782);
  and g1209 (n956, n_780, n_777);
  not g1210 (n_783, n956);
  and g1211 (n957, n_778, n_783);
  not g1212 (n_786, \a[72] );
  not g1213 (n_787, \b[72] );
  and g1214 (n958, n_786, n_787);
  and g1215 (n959, \a[72] , \b[72] );
  not g1216 (n_788, n958);
  not g1217 (n_789, n959);
  and g1218 (n960, n_788, n_789);
  not g1219 (n_790, n960);
  and g1220 (n961, n957, n_790);
  not g1221 (n_791, n957);
  and g1222 (n962, n_791, n960);
  not g1223 (n_792, n961);
  not g1224 (n_793, n962);
  and g1225 (\f[72] , n_792, n_793);
  and g1226 (n964, n_791, n_788);
  not g1227 (n_794, n964);
  and g1228 (n965, n_789, n_794);
  not g1229 (n_797, \a[73] );
  not g1230 (n_798, \b[73] );
  and g1231 (n966, n_797, n_798);
  and g1232 (n967, \a[73] , \b[73] );
  not g1233 (n_799, n966);
  not g1234 (n_800, n967);
  and g1235 (n968, n_799, n_800);
  not g1236 (n_801, n968);
  and g1237 (n969, n965, n_801);
  not g1238 (n_802, n965);
  and g1239 (n970, n_802, n968);
  not g1240 (n_803, n969);
  not g1241 (n_804, n970);
  and g1242 (\f[73] , n_803, n_804);
  and g1243 (n972, n_802, n_799);
  not g1244 (n_805, n972);
  and g1245 (n973, n_800, n_805);
  not g1246 (n_808, \a[74] );
  not g1247 (n_809, \b[74] );
  and g1248 (n974, n_808, n_809);
  and g1249 (n975, \a[74] , \b[74] );
  not g1250 (n_810, n974);
  not g1251 (n_811, n975);
  and g1252 (n976, n_810, n_811);
  not g1253 (n_812, n976);
  and g1254 (n977, n973, n_812);
  not g1255 (n_813, n973);
  and g1256 (n978, n_813, n976);
  not g1257 (n_814, n977);
  not g1258 (n_815, n978);
  and g1259 (\f[74] , n_814, n_815);
  and g1260 (n980, n_813, n_810);
  not g1261 (n_816, n980);
  and g1262 (n981, n_811, n_816);
  not g1263 (n_819, \a[75] );
  not g1264 (n_820, \b[75] );
  and g1265 (n982, n_819, n_820);
  and g1266 (n983, \a[75] , \b[75] );
  not g1267 (n_821, n982);
  not g1268 (n_822, n983);
  and g1269 (n984, n_821, n_822);
  not g1270 (n_823, n984);
  and g1271 (n985, n981, n_823);
  not g1272 (n_824, n981);
  and g1273 (n986, n_824, n984);
  not g1274 (n_825, n985);
  not g1275 (n_826, n986);
  and g1276 (\f[75] , n_825, n_826);
  and g1277 (n988, n_824, n_821);
  not g1278 (n_827, n988);
  and g1279 (n989, n_822, n_827);
  not g1280 (n_830, \a[76] );
  not g1281 (n_831, \b[76] );
  and g1282 (n990, n_830, n_831);
  and g1283 (n991, \a[76] , \b[76] );
  not g1284 (n_832, n990);
  not g1285 (n_833, n991);
  and g1286 (n992, n_832, n_833);
  not g1287 (n_834, n992);
  and g1288 (n993, n989, n_834);
  not g1289 (n_835, n989);
  and g1290 (n994, n_835, n992);
  not g1291 (n_836, n993);
  not g1292 (n_837, n994);
  and g1293 (\f[76] , n_836, n_837);
  and g1294 (n996, n_835, n_832);
  not g1295 (n_838, n996);
  and g1296 (n997, n_833, n_838);
  not g1297 (n_841, \a[77] );
  not g1298 (n_842, \b[77] );
  and g1299 (n998, n_841, n_842);
  and g1300 (n999, \a[77] , \b[77] );
  not g1301 (n_843, n998);
  not g1302 (n_844, n999);
  and g1303 (n1000, n_843, n_844);
  not g1304 (n_845, n1000);
  and g1305 (n1001, n997, n_845);
  not g1306 (n_846, n997);
  and g1307 (n1002, n_846, n1000);
  not g1308 (n_847, n1001);
  not g1309 (n_848, n1002);
  and g1310 (\f[77] , n_847, n_848);
  and g1311 (n1004, n_846, n_843);
  not g1312 (n_849, n1004);
  and g1313 (n1005, n_844, n_849);
  not g1314 (n_852, \a[78] );
  not g1315 (n_853, \b[78] );
  and g1316 (n1006, n_852, n_853);
  and g1317 (n1007, \a[78] , \b[78] );
  not g1318 (n_854, n1006);
  not g1319 (n_855, n1007);
  and g1320 (n1008, n_854, n_855);
  not g1321 (n_856, n1008);
  and g1322 (n1009, n1005, n_856);
  not g1323 (n_857, n1005);
  and g1324 (n1010, n_857, n1008);
  not g1325 (n_858, n1009);
  not g1326 (n_859, n1010);
  and g1327 (\f[78] , n_858, n_859);
  and g1328 (n1012, n_857, n_854);
  not g1329 (n_860, n1012);
  and g1330 (n1013, n_855, n_860);
  not g1331 (n_863, \a[79] );
  not g1332 (n_864, \b[79] );
  and g1333 (n1014, n_863, n_864);
  and g1334 (n1015, \a[79] , \b[79] );
  not g1335 (n_865, n1014);
  not g1336 (n_866, n1015);
  and g1337 (n1016, n_865, n_866);
  not g1338 (n_867, n1016);
  and g1339 (n1017, n1013, n_867);
  not g1340 (n_868, n1013);
  and g1341 (n1018, n_868, n1016);
  not g1342 (n_869, n1017);
  not g1343 (n_870, n1018);
  and g1344 (\f[79] , n_869, n_870);
  and g1345 (n1020, n_868, n_865);
  not g1346 (n_871, n1020);
  and g1347 (n1021, n_866, n_871);
  not g1348 (n_874, \a[80] );
  not g1349 (n_875, \b[80] );
  and g1350 (n1022, n_874, n_875);
  and g1351 (n1023, \a[80] , \b[80] );
  not g1352 (n_876, n1022);
  not g1353 (n_877, n1023);
  and g1354 (n1024, n_876, n_877);
  not g1355 (n_878, n1024);
  and g1356 (n1025, n1021, n_878);
  not g1357 (n_879, n1021);
  and g1358 (n1026, n_879, n1024);
  not g1359 (n_880, n1025);
  not g1360 (n_881, n1026);
  and g1361 (\f[80] , n_880, n_881);
  and g1362 (n1028, n_879, n_876);
  not g1363 (n_882, n1028);
  and g1364 (n1029, n_877, n_882);
  not g1365 (n_885, \a[81] );
  not g1366 (n_886, \b[81] );
  and g1367 (n1030, n_885, n_886);
  and g1368 (n1031, \a[81] , \b[81] );
  not g1369 (n_887, n1030);
  not g1370 (n_888, n1031);
  and g1371 (n1032, n_887, n_888);
  not g1372 (n_889, n1032);
  and g1373 (n1033, n1029, n_889);
  not g1374 (n_890, n1029);
  and g1375 (n1034, n_890, n1032);
  not g1376 (n_891, n1033);
  not g1377 (n_892, n1034);
  and g1378 (\f[81] , n_891, n_892);
  and g1379 (n1036, n_890, n_887);
  not g1380 (n_893, n1036);
  and g1381 (n1037, n_888, n_893);
  not g1382 (n_896, \a[82] );
  not g1383 (n_897, \b[82] );
  and g1384 (n1038, n_896, n_897);
  and g1385 (n1039, \a[82] , \b[82] );
  not g1386 (n_898, n1038);
  not g1387 (n_899, n1039);
  and g1388 (n1040, n_898, n_899);
  not g1389 (n_900, n1040);
  and g1390 (n1041, n1037, n_900);
  not g1391 (n_901, n1037);
  and g1392 (n1042, n_901, n1040);
  not g1393 (n_902, n1041);
  not g1394 (n_903, n1042);
  and g1395 (\f[82] , n_902, n_903);
  and g1396 (n1044, n_901, n_898);
  not g1397 (n_904, n1044);
  and g1398 (n1045, n_899, n_904);
  not g1399 (n_907, \a[83] );
  not g1400 (n_908, \b[83] );
  and g1401 (n1046, n_907, n_908);
  and g1402 (n1047, \a[83] , \b[83] );
  not g1403 (n_909, n1046);
  not g1404 (n_910, n1047);
  and g1405 (n1048, n_909, n_910);
  not g1406 (n_911, n1048);
  and g1407 (n1049, n1045, n_911);
  not g1408 (n_912, n1045);
  and g1409 (n1050, n_912, n1048);
  not g1410 (n_913, n1049);
  not g1411 (n_914, n1050);
  and g1412 (\f[83] , n_913, n_914);
  and g1413 (n1052, n_912, n_909);
  not g1414 (n_915, n1052);
  and g1415 (n1053, n_910, n_915);
  not g1416 (n_918, \a[84] );
  not g1417 (n_919, \b[84] );
  and g1418 (n1054, n_918, n_919);
  and g1419 (n1055, \a[84] , \b[84] );
  not g1420 (n_920, n1054);
  not g1421 (n_921, n1055);
  and g1422 (n1056, n_920, n_921);
  not g1423 (n_922, n1056);
  and g1424 (n1057, n1053, n_922);
  not g1425 (n_923, n1053);
  and g1426 (n1058, n_923, n1056);
  not g1427 (n_924, n1057);
  not g1428 (n_925, n1058);
  and g1429 (\f[84] , n_924, n_925);
  and g1430 (n1060, n_923, n_920);
  not g1431 (n_926, n1060);
  and g1432 (n1061, n_921, n_926);
  not g1433 (n_929, \a[85] );
  not g1434 (n_930, \b[85] );
  and g1435 (n1062, n_929, n_930);
  and g1436 (n1063, \a[85] , \b[85] );
  not g1437 (n_931, n1062);
  not g1438 (n_932, n1063);
  and g1439 (n1064, n_931, n_932);
  not g1440 (n_933, n1064);
  and g1441 (n1065, n1061, n_933);
  not g1442 (n_934, n1061);
  and g1443 (n1066, n_934, n1064);
  not g1444 (n_935, n1065);
  not g1445 (n_936, n1066);
  and g1446 (\f[85] , n_935, n_936);
  and g1447 (n1068, n_934, n_931);
  not g1448 (n_937, n1068);
  and g1449 (n1069, n_932, n_937);
  not g1450 (n_940, \a[86] );
  not g1451 (n_941, \b[86] );
  and g1452 (n1070, n_940, n_941);
  and g1453 (n1071, \a[86] , \b[86] );
  not g1454 (n_942, n1070);
  not g1455 (n_943, n1071);
  and g1456 (n1072, n_942, n_943);
  not g1457 (n_944, n1072);
  and g1458 (n1073, n1069, n_944);
  not g1459 (n_945, n1069);
  and g1460 (n1074, n_945, n1072);
  not g1461 (n_946, n1073);
  not g1462 (n_947, n1074);
  and g1463 (\f[86] , n_946, n_947);
  and g1464 (n1076, n_945, n_942);
  not g1465 (n_948, n1076);
  and g1466 (n1077, n_943, n_948);
  not g1467 (n_951, \a[87] );
  not g1468 (n_952, \b[87] );
  and g1469 (n1078, n_951, n_952);
  and g1470 (n1079, \a[87] , \b[87] );
  not g1471 (n_953, n1078);
  not g1472 (n_954, n1079);
  and g1473 (n1080, n_953, n_954);
  not g1474 (n_955, n1080);
  and g1475 (n1081, n1077, n_955);
  not g1476 (n_956, n1077);
  and g1477 (n1082, n_956, n1080);
  not g1478 (n_957, n1081);
  not g1479 (n_958, n1082);
  and g1480 (\f[87] , n_957, n_958);
  and g1481 (n1084, n_956, n_953);
  not g1482 (n_959, n1084);
  and g1483 (n1085, n_954, n_959);
  not g1484 (n_962, \a[88] );
  not g1485 (n_963, \b[88] );
  and g1486 (n1086, n_962, n_963);
  and g1487 (n1087, \a[88] , \b[88] );
  not g1488 (n_964, n1086);
  not g1489 (n_965, n1087);
  and g1490 (n1088, n_964, n_965);
  not g1491 (n_966, n1088);
  and g1492 (n1089, n1085, n_966);
  not g1493 (n_967, n1085);
  and g1494 (n1090, n_967, n1088);
  not g1495 (n_968, n1089);
  not g1496 (n_969, n1090);
  and g1497 (\f[88] , n_968, n_969);
  and g1498 (n1092, n_967, n_964);
  not g1499 (n_970, n1092);
  and g1500 (n1093, n_965, n_970);
  not g1501 (n_973, \a[89] );
  not g1502 (n_974, \b[89] );
  and g1503 (n1094, n_973, n_974);
  and g1504 (n1095, \a[89] , \b[89] );
  not g1505 (n_975, n1094);
  not g1506 (n_976, n1095);
  and g1507 (n1096, n_975, n_976);
  not g1508 (n_977, n1096);
  and g1509 (n1097, n1093, n_977);
  not g1510 (n_978, n1093);
  and g1511 (n1098, n_978, n1096);
  not g1512 (n_979, n1097);
  not g1513 (n_980, n1098);
  and g1514 (\f[89] , n_979, n_980);
  and g1515 (n1100, n_978, n_975);
  not g1516 (n_981, n1100);
  and g1517 (n1101, n_976, n_981);
  not g1518 (n_984, \a[90] );
  not g1519 (n_985, \b[90] );
  and g1520 (n1102, n_984, n_985);
  and g1521 (n1103, \a[90] , \b[90] );
  not g1522 (n_986, n1102);
  not g1523 (n_987, n1103);
  and g1524 (n1104, n_986, n_987);
  not g1525 (n_988, n1104);
  and g1526 (n1105, n1101, n_988);
  not g1527 (n_989, n1101);
  and g1528 (n1106, n_989, n1104);
  not g1529 (n_990, n1105);
  not g1530 (n_991, n1106);
  and g1531 (\f[90] , n_990, n_991);
  and g1532 (n1108, n_989, n_986);
  not g1533 (n_992, n1108);
  and g1534 (n1109, n_987, n_992);
  not g1535 (n_995, \a[91] );
  not g1536 (n_996, \b[91] );
  and g1537 (n1110, n_995, n_996);
  and g1538 (n1111, \a[91] , \b[91] );
  not g1539 (n_997, n1110);
  not g1540 (n_998, n1111);
  and g1541 (n1112, n_997, n_998);
  not g1542 (n_999, n1112);
  and g1543 (n1113, n1109, n_999);
  not g1544 (n_1000, n1109);
  and g1545 (n1114, n_1000, n1112);
  not g1546 (n_1001, n1113);
  not g1547 (n_1002, n1114);
  and g1548 (\f[91] , n_1001, n_1002);
  and g1549 (n1116, n_1000, n_997);
  not g1550 (n_1003, n1116);
  and g1551 (n1117, n_998, n_1003);
  not g1552 (n_1006, \a[92] );
  not g1553 (n_1007, \b[92] );
  and g1554 (n1118, n_1006, n_1007);
  and g1555 (n1119, \a[92] , \b[92] );
  not g1556 (n_1008, n1118);
  not g1557 (n_1009, n1119);
  and g1558 (n1120, n_1008, n_1009);
  not g1559 (n_1010, n1120);
  and g1560 (n1121, n1117, n_1010);
  not g1561 (n_1011, n1117);
  and g1562 (n1122, n_1011, n1120);
  not g1563 (n_1012, n1121);
  not g1564 (n_1013, n1122);
  and g1565 (\f[92] , n_1012, n_1013);
  and g1566 (n1124, n_1011, n_1008);
  not g1567 (n_1014, n1124);
  and g1568 (n1125, n_1009, n_1014);
  not g1569 (n_1017, \a[93] );
  not g1570 (n_1018, \b[93] );
  and g1571 (n1126, n_1017, n_1018);
  and g1572 (n1127, \a[93] , \b[93] );
  not g1573 (n_1019, n1126);
  not g1574 (n_1020, n1127);
  and g1575 (n1128, n_1019, n_1020);
  not g1576 (n_1021, n1128);
  and g1577 (n1129, n1125, n_1021);
  not g1578 (n_1022, n1125);
  and g1579 (n1130, n_1022, n1128);
  not g1580 (n_1023, n1129);
  not g1581 (n_1024, n1130);
  and g1582 (\f[93] , n_1023, n_1024);
  and g1583 (n1132, n_1022, n_1019);
  not g1584 (n_1025, n1132);
  and g1585 (n1133, n_1020, n_1025);
  not g1586 (n_1028, \a[94] );
  not g1587 (n_1029, \b[94] );
  and g1588 (n1134, n_1028, n_1029);
  and g1589 (n1135, \a[94] , \b[94] );
  not g1590 (n_1030, n1134);
  not g1591 (n_1031, n1135);
  and g1592 (n1136, n_1030, n_1031);
  not g1593 (n_1032, n1136);
  and g1594 (n1137, n1133, n_1032);
  not g1595 (n_1033, n1133);
  and g1596 (n1138, n_1033, n1136);
  not g1597 (n_1034, n1137);
  not g1598 (n_1035, n1138);
  and g1599 (\f[94] , n_1034, n_1035);
  and g1600 (n1140, n_1033, n_1030);
  not g1601 (n_1036, n1140);
  and g1602 (n1141, n_1031, n_1036);
  not g1603 (n_1039, \a[95] );
  not g1604 (n_1040, \b[95] );
  and g1605 (n1142, n_1039, n_1040);
  and g1606 (n1143, \a[95] , \b[95] );
  not g1607 (n_1041, n1142);
  not g1608 (n_1042, n1143);
  and g1609 (n1144, n_1041, n_1042);
  not g1610 (n_1043, n1144);
  and g1611 (n1145, n1141, n_1043);
  not g1612 (n_1044, n1141);
  and g1613 (n1146, n_1044, n1144);
  not g1614 (n_1045, n1145);
  not g1615 (n_1046, n1146);
  and g1616 (\f[95] , n_1045, n_1046);
  and g1617 (n1148, n_1044, n_1041);
  not g1618 (n_1047, n1148);
  and g1619 (n1149, n_1042, n_1047);
  not g1620 (n_1050, \a[96] );
  not g1621 (n_1051, \b[96] );
  and g1622 (n1150, n_1050, n_1051);
  and g1623 (n1151, \a[96] , \b[96] );
  not g1624 (n_1052, n1150);
  not g1625 (n_1053, n1151);
  and g1626 (n1152, n_1052, n_1053);
  not g1627 (n_1054, n1152);
  and g1628 (n1153, n1149, n_1054);
  not g1629 (n_1055, n1149);
  and g1630 (n1154, n_1055, n1152);
  not g1631 (n_1056, n1153);
  not g1632 (n_1057, n1154);
  and g1633 (\f[96] , n_1056, n_1057);
  and g1634 (n1156, n_1055, n_1052);
  not g1635 (n_1058, n1156);
  and g1636 (n1157, n_1053, n_1058);
  not g1637 (n_1061, \a[97] );
  not g1638 (n_1062, \b[97] );
  and g1639 (n1158, n_1061, n_1062);
  and g1640 (n1159, \a[97] , \b[97] );
  not g1641 (n_1063, n1158);
  not g1642 (n_1064, n1159);
  and g1643 (n1160, n_1063, n_1064);
  not g1644 (n_1065, n1160);
  and g1645 (n1161, n1157, n_1065);
  not g1646 (n_1066, n1157);
  and g1647 (n1162, n_1066, n1160);
  not g1648 (n_1067, n1161);
  not g1649 (n_1068, n1162);
  and g1650 (\f[97] , n_1067, n_1068);
  and g1651 (n1164, n_1066, n_1063);
  not g1652 (n_1069, n1164);
  and g1653 (n1165, n_1064, n_1069);
  not g1654 (n_1072, \a[98] );
  not g1655 (n_1073, \b[98] );
  and g1656 (n1166, n_1072, n_1073);
  and g1657 (n1167, \a[98] , \b[98] );
  not g1658 (n_1074, n1166);
  not g1659 (n_1075, n1167);
  and g1660 (n1168, n_1074, n_1075);
  not g1661 (n_1076, n1168);
  and g1662 (n1169, n1165, n_1076);
  not g1663 (n_1077, n1165);
  and g1664 (n1170, n_1077, n1168);
  not g1665 (n_1078, n1169);
  not g1666 (n_1079, n1170);
  and g1667 (\f[98] , n_1078, n_1079);
  and g1668 (n1172, n_1077, n_1074);
  not g1669 (n_1080, n1172);
  and g1670 (n1173, n_1075, n_1080);
  not g1671 (n_1083, \a[99] );
  not g1672 (n_1084, \b[99] );
  and g1673 (n1174, n_1083, n_1084);
  and g1674 (n1175, \a[99] , \b[99] );
  not g1675 (n_1085, n1174);
  not g1676 (n_1086, n1175);
  and g1677 (n1176, n_1085, n_1086);
  not g1678 (n_1087, n1176);
  and g1679 (n1177, n1173, n_1087);
  not g1680 (n_1088, n1173);
  and g1681 (n1178, n_1088, n1176);
  not g1682 (n_1089, n1177);
  not g1683 (n_1090, n1178);
  and g1684 (\f[99] , n_1089, n_1090);
  and g1685 (n1180, n_1088, n_1085);
  not g1686 (n_1091, n1180);
  and g1687 (n1181, n_1086, n_1091);
  not g1688 (n_1094, \a[100] );
  not g1689 (n_1095, \b[100] );
  and g1690 (n1182, n_1094, n_1095);
  and g1691 (n1183, \a[100] , \b[100] );
  not g1692 (n_1096, n1182);
  not g1693 (n_1097, n1183);
  and g1694 (n1184, n_1096, n_1097);
  not g1695 (n_1098, n1184);
  and g1696 (n1185, n1181, n_1098);
  not g1697 (n_1099, n1181);
  and g1698 (n1186, n_1099, n1184);
  not g1699 (n_1100, n1185);
  not g1700 (n_1101, n1186);
  and g1701 (\f[100] , n_1100, n_1101);
  and g1702 (n1188, n_1099, n_1096);
  not g1703 (n_1102, n1188);
  and g1704 (n1189, n_1097, n_1102);
  not g1705 (n_1105, \a[101] );
  not g1706 (n_1106, \b[101] );
  and g1707 (n1190, n_1105, n_1106);
  and g1708 (n1191, \a[101] , \b[101] );
  not g1709 (n_1107, n1190);
  not g1710 (n_1108, n1191);
  and g1711 (n1192, n_1107, n_1108);
  not g1712 (n_1109, n1192);
  and g1713 (n1193, n1189, n_1109);
  not g1714 (n_1110, n1189);
  and g1715 (n1194, n_1110, n1192);
  not g1716 (n_1111, n1193);
  not g1717 (n_1112, n1194);
  and g1718 (\f[101] , n_1111, n_1112);
  and g1719 (n1196, n_1110, n_1107);
  not g1720 (n_1113, n1196);
  and g1721 (n1197, n_1108, n_1113);
  not g1722 (n_1116, \a[102] );
  not g1723 (n_1117, \b[102] );
  and g1724 (n1198, n_1116, n_1117);
  and g1725 (n1199, \a[102] , \b[102] );
  not g1726 (n_1118, n1198);
  not g1727 (n_1119, n1199);
  and g1728 (n1200, n_1118, n_1119);
  not g1729 (n_1120, n1200);
  and g1730 (n1201, n1197, n_1120);
  not g1731 (n_1121, n1197);
  and g1732 (n1202, n_1121, n1200);
  not g1733 (n_1122, n1201);
  not g1734 (n_1123, n1202);
  and g1735 (\f[102] , n_1122, n_1123);
  and g1736 (n1204, n_1121, n_1118);
  not g1737 (n_1124, n1204);
  and g1738 (n1205, n_1119, n_1124);
  not g1739 (n_1127, \a[103] );
  not g1740 (n_1128, \b[103] );
  and g1741 (n1206, n_1127, n_1128);
  and g1742 (n1207, \a[103] , \b[103] );
  not g1743 (n_1129, n1206);
  not g1744 (n_1130, n1207);
  and g1745 (n1208, n_1129, n_1130);
  not g1746 (n_1131, n1208);
  and g1747 (n1209, n1205, n_1131);
  not g1748 (n_1132, n1205);
  and g1749 (n1210, n_1132, n1208);
  not g1750 (n_1133, n1209);
  not g1751 (n_1134, n1210);
  and g1752 (\f[103] , n_1133, n_1134);
  and g1753 (n1212, n_1132, n_1129);
  not g1754 (n_1135, n1212);
  and g1755 (n1213, n_1130, n_1135);
  not g1756 (n_1138, \a[104] );
  not g1757 (n_1139, \b[104] );
  and g1758 (n1214, n_1138, n_1139);
  and g1759 (n1215, \a[104] , \b[104] );
  not g1760 (n_1140, n1214);
  not g1761 (n_1141, n1215);
  and g1762 (n1216, n_1140, n_1141);
  not g1763 (n_1142, n1216);
  and g1764 (n1217, n1213, n_1142);
  not g1765 (n_1143, n1213);
  and g1766 (n1218, n_1143, n1216);
  not g1767 (n_1144, n1217);
  not g1768 (n_1145, n1218);
  and g1769 (\f[104] , n_1144, n_1145);
  and g1770 (n1220, n_1143, n_1140);
  not g1771 (n_1146, n1220);
  and g1772 (n1221, n_1141, n_1146);
  not g1773 (n_1149, \a[105] );
  not g1774 (n_1150, \b[105] );
  and g1775 (n1222, n_1149, n_1150);
  and g1776 (n1223, \a[105] , \b[105] );
  not g1777 (n_1151, n1222);
  not g1778 (n_1152, n1223);
  and g1779 (n1224, n_1151, n_1152);
  not g1780 (n_1153, n1224);
  and g1781 (n1225, n1221, n_1153);
  not g1782 (n_1154, n1221);
  and g1783 (n1226, n_1154, n1224);
  not g1784 (n_1155, n1225);
  not g1785 (n_1156, n1226);
  and g1786 (\f[105] , n_1155, n_1156);
  and g1787 (n1228, n_1154, n_1151);
  not g1788 (n_1157, n1228);
  and g1789 (n1229, n_1152, n_1157);
  not g1790 (n_1160, \a[106] );
  not g1791 (n_1161, \b[106] );
  and g1792 (n1230, n_1160, n_1161);
  and g1793 (n1231, \a[106] , \b[106] );
  not g1794 (n_1162, n1230);
  not g1795 (n_1163, n1231);
  and g1796 (n1232, n_1162, n_1163);
  not g1797 (n_1164, n1232);
  and g1798 (n1233, n1229, n_1164);
  not g1799 (n_1165, n1229);
  and g1800 (n1234, n_1165, n1232);
  not g1801 (n_1166, n1233);
  not g1802 (n_1167, n1234);
  and g1803 (\f[106] , n_1166, n_1167);
  and g1804 (n1236, n_1165, n_1162);
  not g1805 (n_1168, n1236);
  and g1806 (n1237, n_1163, n_1168);
  not g1807 (n_1171, \a[107] );
  not g1808 (n_1172, \b[107] );
  and g1809 (n1238, n_1171, n_1172);
  and g1810 (n1239, \a[107] , \b[107] );
  not g1811 (n_1173, n1238);
  not g1812 (n_1174, n1239);
  and g1813 (n1240, n_1173, n_1174);
  not g1814 (n_1175, n1240);
  and g1815 (n1241, n1237, n_1175);
  not g1816 (n_1176, n1237);
  and g1817 (n1242, n_1176, n1240);
  not g1818 (n_1177, n1241);
  not g1819 (n_1178, n1242);
  and g1820 (\f[107] , n_1177, n_1178);
  and g1821 (n1244, n_1176, n_1173);
  not g1822 (n_1179, n1244);
  and g1823 (n1245, n_1174, n_1179);
  not g1824 (n_1182, \a[108] );
  not g1825 (n_1183, \b[108] );
  and g1826 (n1246, n_1182, n_1183);
  and g1827 (n1247, \a[108] , \b[108] );
  not g1828 (n_1184, n1246);
  not g1829 (n_1185, n1247);
  and g1830 (n1248, n_1184, n_1185);
  not g1831 (n_1186, n1248);
  and g1832 (n1249, n1245, n_1186);
  not g1833 (n_1187, n1245);
  and g1834 (n1250, n_1187, n1248);
  not g1835 (n_1188, n1249);
  not g1836 (n_1189, n1250);
  and g1837 (\f[108] , n_1188, n_1189);
  and g1838 (n1252, n_1187, n_1184);
  not g1839 (n_1190, n1252);
  and g1840 (n1253, n_1185, n_1190);
  not g1841 (n_1193, \a[109] );
  not g1842 (n_1194, \b[109] );
  and g1843 (n1254, n_1193, n_1194);
  and g1844 (n1255, \a[109] , \b[109] );
  not g1845 (n_1195, n1254);
  not g1846 (n_1196, n1255);
  and g1847 (n1256, n_1195, n_1196);
  not g1848 (n_1197, n1256);
  and g1849 (n1257, n1253, n_1197);
  not g1850 (n_1198, n1253);
  and g1851 (n1258, n_1198, n1256);
  not g1852 (n_1199, n1257);
  not g1853 (n_1200, n1258);
  and g1854 (\f[109] , n_1199, n_1200);
  and g1855 (n1260, n_1198, n_1195);
  not g1856 (n_1201, n1260);
  and g1857 (n1261, n_1196, n_1201);
  not g1858 (n_1204, \a[110] );
  not g1859 (n_1205, \b[110] );
  and g1860 (n1262, n_1204, n_1205);
  and g1861 (n1263, \a[110] , \b[110] );
  not g1862 (n_1206, n1262);
  not g1863 (n_1207, n1263);
  and g1864 (n1264, n_1206, n_1207);
  not g1865 (n_1208, n1264);
  and g1866 (n1265, n1261, n_1208);
  not g1867 (n_1209, n1261);
  and g1868 (n1266, n_1209, n1264);
  not g1869 (n_1210, n1265);
  not g1870 (n_1211, n1266);
  and g1871 (\f[110] , n_1210, n_1211);
  and g1872 (n1268, n_1209, n_1206);
  not g1873 (n_1212, n1268);
  and g1874 (n1269, n_1207, n_1212);
  not g1875 (n_1215, \a[111] );
  not g1876 (n_1216, \b[111] );
  and g1877 (n1270, n_1215, n_1216);
  and g1878 (n1271, \a[111] , \b[111] );
  not g1879 (n_1217, n1270);
  not g1880 (n_1218, n1271);
  and g1881 (n1272, n_1217, n_1218);
  not g1882 (n_1219, n1272);
  and g1883 (n1273, n1269, n_1219);
  not g1884 (n_1220, n1269);
  and g1885 (n1274, n_1220, n1272);
  not g1886 (n_1221, n1273);
  not g1887 (n_1222, n1274);
  and g1888 (\f[111] , n_1221, n_1222);
  and g1889 (n1276, n_1220, n_1217);
  not g1890 (n_1223, n1276);
  and g1891 (n1277, n_1218, n_1223);
  not g1892 (n_1226, \a[112] );
  not g1893 (n_1227, \b[112] );
  and g1894 (n1278, n_1226, n_1227);
  and g1895 (n1279, \a[112] , \b[112] );
  not g1896 (n_1228, n1278);
  not g1897 (n_1229, n1279);
  and g1898 (n1280, n_1228, n_1229);
  not g1899 (n_1230, n1280);
  and g1900 (n1281, n1277, n_1230);
  not g1901 (n_1231, n1277);
  and g1902 (n1282, n_1231, n1280);
  not g1903 (n_1232, n1281);
  not g1904 (n_1233, n1282);
  and g1905 (\f[112] , n_1232, n_1233);
  and g1906 (n1284, n_1231, n_1228);
  not g1907 (n_1234, n1284);
  and g1908 (n1285, n_1229, n_1234);
  not g1909 (n_1237, \a[113] );
  not g1910 (n_1238, \b[113] );
  and g1911 (n1286, n_1237, n_1238);
  and g1912 (n1287, \a[113] , \b[113] );
  not g1913 (n_1239, n1286);
  not g1914 (n_1240, n1287);
  and g1915 (n1288, n_1239, n_1240);
  not g1916 (n_1241, n1288);
  and g1917 (n1289, n1285, n_1241);
  not g1918 (n_1242, n1285);
  and g1919 (n1290, n_1242, n1288);
  not g1920 (n_1243, n1289);
  not g1921 (n_1244, n1290);
  and g1922 (\f[113] , n_1243, n_1244);
  and g1923 (n1292, n_1242, n_1239);
  not g1924 (n_1245, n1292);
  and g1925 (n1293, n_1240, n_1245);
  not g1926 (n_1248, \a[114] );
  not g1927 (n_1249, \b[114] );
  and g1928 (n1294, n_1248, n_1249);
  and g1929 (n1295, \a[114] , \b[114] );
  not g1930 (n_1250, n1294);
  not g1931 (n_1251, n1295);
  and g1932 (n1296, n_1250, n_1251);
  not g1933 (n_1252, n1296);
  and g1934 (n1297, n1293, n_1252);
  not g1935 (n_1253, n1293);
  and g1936 (n1298, n_1253, n1296);
  not g1937 (n_1254, n1297);
  not g1938 (n_1255, n1298);
  and g1939 (\f[114] , n_1254, n_1255);
  and g1940 (n1300, n_1253, n_1250);
  not g1941 (n_1256, n1300);
  and g1942 (n1301, n_1251, n_1256);
  not g1943 (n_1259, \a[115] );
  not g1944 (n_1260, \b[115] );
  and g1945 (n1302, n_1259, n_1260);
  and g1946 (n1303, \a[115] , \b[115] );
  not g1947 (n_1261, n1302);
  not g1948 (n_1262, n1303);
  and g1949 (n1304, n_1261, n_1262);
  not g1950 (n_1263, n1304);
  and g1951 (n1305, n1301, n_1263);
  not g1952 (n_1264, n1301);
  and g1953 (n1306, n_1264, n1304);
  not g1954 (n_1265, n1305);
  not g1955 (n_1266, n1306);
  and g1956 (\f[115] , n_1265, n_1266);
  and g1957 (n1308, n_1264, n_1261);
  not g1958 (n_1267, n1308);
  and g1959 (n1309, n_1262, n_1267);
  not g1960 (n_1270, \a[116] );
  not g1961 (n_1271, \b[116] );
  and g1962 (n1310, n_1270, n_1271);
  and g1963 (n1311, \a[116] , \b[116] );
  not g1964 (n_1272, n1310);
  not g1965 (n_1273, n1311);
  and g1966 (n1312, n_1272, n_1273);
  not g1967 (n_1274, n1312);
  and g1968 (n1313, n1309, n_1274);
  not g1969 (n_1275, n1309);
  and g1970 (n1314, n_1275, n1312);
  not g1971 (n_1276, n1313);
  not g1972 (n_1277, n1314);
  and g1973 (\f[116] , n_1276, n_1277);
  and g1974 (n1316, n_1275, n_1272);
  not g1975 (n_1278, n1316);
  and g1976 (n1317, n_1273, n_1278);
  not g1977 (n_1281, \a[117] );
  not g1978 (n_1282, \b[117] );
  and g1979 (n1318, n_1281, n_1282);
  and g1980 (n1319, \a[117] , \b[117] );
  not g1981 (n_1283, n1318);
  not g1982 (n_1284, n1319);
  and g1983 (n1320, n_1283, n_1284);
  not g1984 (n_1285, n1320);
  and g1985 (n1321, n1317, n_1285);
  not g1986 (n_1286, n1317);
  and g1987 (n1322, n_1286, n1320);
  not g1988 (n_1287, n1321);
  not g1989 (n_1288, n1322);
  and g1990 (\f[117] , n_1287, n_1288);
  and g1991 (n1324, n_1286, n_1283);
  not g1992 (n_1289, n1324);
  and g1993 (n1325, n_1284, n_1289);
  not g1994 (n_1292, \a[118] );
  not g1995 (n_1293, \b[118] );
  and g1996 (n1326, n_1292, n_1293);
  and g1997 (n1327, \a[118] , \b[118] );
  not g1998 (n_1294, n1326);
  not g1999 (n_1295, n1327);
  and g2000 (n1328, n_1294, n_1295);
  not g2001 (n_1296, n1328);
  and g2002 (n1329, n1325, n_1296);
  not g2003 (n_1297, n1325);
  and g2004 (n1330, n_1297, n1328);
  not g2005 (n_1298, n1329);
  not g2006 (n_1299, n1330);
  and g2007 (\f[118] , n_1298, n_1299);
  and g2008 (n1332, n_1297, n_1294);
  not g2009 (n_1300, n1332);
  and g2010 (n1333, n_1295, n_1300);
  not g2011 (n_1303, \a[119] );
  not g2012 (n_1304, \b[119] );
  and g2013 (n1334, n_1303, n_1304);
  and g2014 (n1335, \a[119] , \b[119] );
  not g2015 (n_1305, n1334);
  not g2016 (n_1306, n1335);
  and g2017 (n1336, n_1305, n_1306);
  not g2018 (n_1307, n1336);
  and g2019 (n1337, n1333, n_1307);
  not g2020 (n_1308, n1333);
  and g2021 (n1338, n_1308, n1336);
  not g2022 (n_1309, n1337);
  not g2023 (n_1310, n1338);
  and g2024 (\f[119] , n_1309, n_1310);
  and g2025 (n1340, n_1308, n_1305);
  not g2026 (n_1311, n1340);
  and g2027 (n1341, n_1306, n_1311);
  not g2028 (n_1314, \a[120] );
  not g2029 (n_1315, \b[120] );
  and g2030 (n1342, n_1314, n_1315);
  and g2031 (n1343, \a[120] , \b[120] );
  not g2032 (n_1316, n1342);
  not g2033 (n_1317, n1343);
  and g2034 (n1344, n_1316, n_1317);
  not g2035 (n_1318, n1344);
  and g2036 (n1345, n1341, n_1318);
  not g2037 (n_1319, n1341);
  and g2038 (n1346, n_1319, n1344);
  not g2039 (n_1320, n1345);
  not g2040 (n_1321, n1346);
  and g2041 (\f[120] , n_1320, n_1321);
  and g2042 (n1348, n_1319, n_1316);
  not g2043 (n_1322, n1348);
  and g2044 (n1349, n_1317, n_1322);
  not g2045 (n_1325, \a[121] );
  not g2046 (n_1326, \b[121] );
  and g2047 (n1350, n_1325, n_1326);
  and g2048 (n1351, \a[121] , \b[121] );
  not g2049 (n_1327, n1350);
  not g2050 (n_1328, n1351);
  and g2051 (n1352, n_1327, n_1328);
  not g2052 (n_1329, n1352);
  and g2053 (n1353, n1349, n_1329);
  not g2054 (n_1330, n1349);
  and g2055 (n1354, n_1330, n1352);
  not g2056 (n_1331, n1353);
  not g2057 (n_1332, n1354);
  and g2058 (\f[121] , n_1331, n_1332);
  and g2059 (n1356, n_1330, n_1327);
  not g2060 (n_1333, n1356);
  and g2061 (n1357, n_1328, n_1333);
  not g2062 (n_1336, \a[122] );
  not g2063 (n_1337, \b[122] );
  and g2064 (n1358, n_1336, n_1337);
  and g2065 (n1359, \a[122] , \b[122] );
  not g2066 (n_1338, n1358);
  not g2067 (n_1339, n1359);
  and g2068 (n1360, n_1338, n_1339);
  not g2069 (n_1340, n1360);
  and g2070 (n1361, n1357, n_1340);
  not g2071 (n_1341, n1357);
  and g2072 (n1362, n_1341, n1360);
  not g2073 (n_1342, n1361);
  not g2074 (n_1343, n1362);
  and g2075 (\f[122] , n_1342, n_1343);
  and g2076 (n1364, n_1341, n_1338);
  not g2077 (n_1344, n1364);
  and g2078 (n1365, n_1339, n_1344);
  not g2079 (n_1347, \a[123] );
  not g2080 (n_1348, \b[123] );
  and g2081 (n1366, n_1347, n_1348);
  and g2082 (n1367, \a[123] , \b[123] );
  not g2083 (n_1349, n1366);
  not g2084 (n_1350, n1367);
  and g2085 (n1368, n_1349, n_1350);
  not g2086 (n_1351, n1368);
  and g2087 (n1369, n1365, n_1351);
  not g2088 (n_1352, n1365);
  and g2089 (n1370, n_1352, n1368);
  not g2090 (n_1353, n1369);
  not g2091 (n_1354, n1370);
  and g2092 (\f[123] , n_1353, n_1354);
  and g2093 (n1372, n_1352, n_1349);
  not g2094 (n_1355, n1372);
  and g2095 (n1373, n_1350, n_1355);
  not g2096 (n_1358, \a[124] );
  not g2097 (n_1359, \b[124] );
  and g2098 (n1374, n_1358, n_1359);
  and g2099 (n1375, \a[124] , \b[124] );
  not g2100 (n_1360, n1374);
  not g2101 (n_1361, n1375);
  and g2102 (n1376, n_1360, n_1361);
  not g2103 (n_1362, n1376);
  and g2104 (n1377, n1373, n_1362);
  not g2105 (n_1363, n1373);
  and g2106 (n1378, n_1363, n1376);
  not g2107 (n_1364, n1377);
  not g2108 (n_1365, n1378);
  and g2109 (\f[124] , n_1364, n_1365);
  and g2110 (n1380, n_1363, n_1360);
  not g2111 (n_1366, n1380);
  and g2112 (n1381, n_1361, n_1366);
  not g2113 (n_1369, \a[125] );
  not g2114 (n_1370, \b[125] );
  and g2115 (n1382, n_1369, n_1370);
  and g2116 (n1383, \a[125] , \b[125] );
  not g2117 (n_1371, n1382);
  not g2118 (n_1372, n1383);
  and g2119 (n1384, n_1371, n_1372);
  not g2120 (n_1373, n1384);
  and g2121 (n1385, n1381, n_1373);
  not g2122 (n_1374, n1381);
  and g2123 (n1386, n_1374, n1384);
  not g2124 (n_1375, n1385);
  not g2125 (n_1376, n1386);
  and g2126 (\f[125] , n_1375, n_1376);
  and g2127 (n1388, n_1374, n_1371);
  not g2128 (n_1377, n1388);
  and g2129 (n1389, n_1372, n_1377);
  not g2130 (n_1380, \a[126] );
  not g2131 (n_1381, \b[126] );
  and g2132 (n1390, n_1380, n_1381);
  and g2133 (n1391, \a[126] , \b[126] );
  not g2134 (n_1382, n1390);
  not g2135 (n_1383, n1391);
  and g2136 (n1392, n_1382, n_1383);
  not g2137 (n_1384, n1392);
  and g2138 (n1393, n1389, n_1384);
  not g2139 (n_1385, n1389);
  and g2140 (n1394, n_1385, n1392);
  not g2141 (n_1386, n1393);
  not g2142 (n_1387, n1394);
  and g2143 (\f[126] , n_1386, n_1387);
  and g2144 (n1396, n_1385, n_1382);
  not g2145 (n_1388, n1396);
  and g2146 (n1397, n_1383, n_1388);
  not g2147 (n_1391, \a[127] );
  not g2148 (n_1392, \b[127] );
  and g2149 (n1398, n_1391, n_1392);
  and g2150 (n1399, \a[127] , \b[127] );
  not g2151 (n_1393, n1398);
  not g2152 (n_1394, n1399);
  and g2153 (n1400, n_1393, n_1394);
  not g2154 (n_1395, n1400);
  and g2155 (n1401, n1397, n_1395);
  not g2156 (n_1396, n1397);
  and g2157 (n1402, n_1396, n1400);
  not g2158 (n_1397, n1401);
  not g2159 (n_1398, n1402);
  and g2160 (\f[127] , n_1397, n_1398);
  and g2161 (n1404, n_1396, n_1393);
  or g2162 (cOut, n1399, n1404);
endmodule

