//# 62 inputs
//# 152 outputs
//# 638 D-type flipflops
//# 5378 inverters
//# 2573 gates (1114 ANDs + 849 NANDs + 512 ORs + 98 NORs)

mmodule dff(CK,q,d);
input CK,d;
output reg q;
always @ (negedge CK)
q<=d;
endmodule


module s13207a(GND,VDD,CK,g1,g10,g1000,g1006,g1008,g1015,g1016,g1017,g1080,g11,
  g1193,
  g1194,g1195,g1196,g1197,g1198,g1201,g1202,g1203,g1205,g1206,g1234,g1246,
  g1553,g1554,g1724,g1783,g1798,g1804,g1810,g1817,g1824,g1829,g1870,g1871,
  g1894,g1911,g1944,g206,g21,g22,g23,g24,g25,g26,g2662,g27,g28,g2844,g2888,g29,
  g291,g30,g3077,g3096,g31,g3130,g3159,g3191,g32,g37,g372,g3829,g3854,g3856,
  g3857,g3859,g3860,g41,g42,g4267,g43,g4316,g4370,g4371,g4372,g4373,g44,g45,
  g453,g4655,g4657,g4660,g4661,g4663,g4664,g49,g5143,g5164,g534,g5571,g5669,
  g5678,g5682,g5684,g5687,g5729,g594,g6207,g6212,g6223,g6236,g6269,g6288,g6289,
  g6290,g6291,g6292,g6293,g6294,g6295,g6296,g6297,g6298,g6299,g6300,g6301,
  g6302,g6303,g6304,g6305,g6306,g6307,g6308,g633,g634,g635,g6376,g6425,g645,
  g647,g648,g6648,g6653,g6675,g6849,g6850,g6895,g690,g6909,g694,g698,g702,
  g7048,g7063,g7103,g722,g723,g7283,g7284,g7285,g7286,g7287,g7288,g7289,g7290,
  g7291,g7292,g7293,g7294,g7295,g7298,g7423,g7424,g7425,g7474,g7504,g7505,
  g7506,g7507,g7508,g751,g7514,g752,g753,g754,g755,g756,g757,g7729,g7730,g7731,
  g7732,g7763,g781,g785,g786,g795,g8216,g8217,g8218,g8219,g8234,g8661,g8663,
  g8872,g8958,g9,g9128,g9132,g9204,g9280,g929,g9297,g9299,g9305,g9308,g9310,
  g9312,g9314,g9378,g941,g955,g962);
input GND,VDD,CK,g43,g49,g633,g634,g635,g645,g647,g648,g690,g694,g698,g702,
  g722,g723,g751,
  g752,g753,g754,g755,g756,g757,g781,g941,g962,g1000,g1008,g1016,g1080,g1234,
  g1553,g1554,g786,g1206,g929,g955,g795,g1194,g1198,g1202,g24,g1203,g1196,g29,
  g22,g28,g10,g23,g37,g26,g1,g27,g42,g11,g32,g41,g31,g45,g9,g44,g21,g30,g25;
output g206,g291,g372,g453,g534,g594,g785,g1006,g1015,g1017,g1246,g1724,g1783,
  g1798,g1804,g1810,g1817,g1824,g1829,g1870,g1871,g1894,g1911,g1944,g2662,
  g2844,g2888,g3077,g3096,g3130,g3159,g3191,g3829,g3859,g3860,g4267,g4316,
  g4370,g4371,g4372,g4373,g4655,g4657,g4660,g4661,g4663,g4664,g5143,g5164,
  g5571,g5669,g5678,g5682,g5684,g5687,g5729,g6207,g6212,g6223,g6236,g6269,
  g6425,g6648,g6653,g6675,g6849,g6850,g6895,g6909,g7048,g7063,g7103,g7283,
  g7284,g7285,g7286,g7287,g7288,g7289,g7290,g7291,g7292,g7293,g7294,g7295,
  g7298,g7423,g7424,g7425,g7474,g7504,g7505,g7506,g7507,g7508,g7514,g7729,
  g7730,g7731,g7732,g8216,g8217,g8218,g8219,g8234,g8661,g8663,g8872,g8958,
  g9128,g9132,g9204,g9280,g9297,g9299,g9305,g9308,g9310,g9312,g9314,g9378,
  g7763,g1205,g3856,g3857,g3854,g1193,g1197,g1201,g6294,g6376,g1195,g6300,
  g6292,g6298,g6291,g6293,g6304,g6296,g6289,g6297,g6306,g6290,g6303,g6305,
  g6302,g6308,g6288,g6307,g6299,g6301,g6295;

  wire g397,g4635,g1271,g5176,g312,g4618,g273,g4611,g452,g449,g948,g8664,g629,
    g6827,g207,g5733,g1541,g7778,g1153,g6856,g940,g5735,g976,g8864,g498,g9111,
    g314,g4620,g1092,g7520,g454,g4639,g196,g5731,g535,g3844,g292,g4613,g772,
    g6846,g1375,g6869,g689,g6371,g183,g6309,g359,g6336,g1384,g6881,g1339,g6865,
    g20,g6386,g1424,g3862,g767,g6841,g393,g4631,g1077,g7767,g1231,g1236,g294,
    g4615,g1477,g9036,g4,g9372,g608,g6806,g1204,g465,g6352,g774,g6848,g921,
    g916,g1304,g1312,g243,g6318,g1499,g7772,g80,g6778,g1444,g5185,g1269,g5740,
    g600,g6807,g423,g9105,g771,g6845,g803,g7757,g843,g2647,g315,g4621,g455,
    g4640,g906,g901,g622,g6821,g891,g3855,g1014,g1012,g984,g9133,g117,g5153,
    g137,g5150,g527,g9110,g1513,g1524,g278,g6323,g1378,g6880,g718,g7753,g598,
    g6797,g1182,g1160,g1288,g7527,g1382,g6888,g179,g5159,g624,g6831,g48,g9362,
    g362,g9093,g878,g890,g270,g9092,g763,g6836,g710,g7751,g730,g7754,g295,
    g4616,g1037,g7519,g1102,g6855,g483,g6356,g775,g7759,g621,g6819,g1364,g6878,
    g1454,g5187,g1296,g7304,g5,g9373,g1532,g7781,g587,g3852,g741,g9386,g13,
    g7308,g606,g6804,g6851,g52,g6781,g646,g4652,g1412,g5745,g327,g6332,g1189,
    g6392,g1389,g4658,g1029,g2654,g1371,g6868,g1429,g2671,g398,g4636,g985,
    g7515,g354,g4624,g619,g6817,g113,g5148,g133,g5149,g180,g5158,g1138,g7524,
    g1309,g1308,g889,g7101,g390,g6341,g625,g6823,g417,g9103,g681,g7748,g437,
    g6348,g351,g9100,g1200,g109,g6785,g1049,g8673,g1098,g6854,g200,g199,g240,
    g6317,g479,g4649,g126,g6789,g596,g6795,g1268,g5175,g222,g6313,g420,g9104,
    g3,g9360,g58,g7734,g172,g1270,g387,g6340,g840,g2648,g365,g9094,g1486,g8226,
    g1504,g7773,g1185,g1155,g1385,g6883,g583,g3851,g822,g7512,g1025,g8871,g969,
    g966,g768,g6842,g174,g7737,g685,g7749,g1087,g6853,g355,g4625,g911,g1226,
    g6859,g99,g6783,g1045,g8224,g1173,g7526,g1373,g6871,g186,g3830,g760,g6833,
    g959,g5169,g1369,g6875,g1007,g8867,g1459,g3863,g758,g6840,g480,g6355,g396,
    g4634,g612,g6811,g38,g5746,g632,g6830,g1415,g5180,g1227,g7108,g246,g6319,
    g3840,g517,g4651,g118,g6787,g138,g6792,g16,g1404,g284,g9086,g142,g6793,
    g219,g6312,g426,g9106,g1388,g6882,g806,g7510,g846,g2646,g1428,g2672,g579,
    g3850,g1030,g7518,g614,g6812,g1430,g4666,g1247,g6380,g669,g7745,g110,g130,
    g6790,g225,g6314,g281,g9085,g819,g7761,g6385,g611,g6810,g631,g6829,g1217,
    g6377,g104,g6784,g1365,g6867,g825,g7513,g1333,g6863,g474,g4644,g1396,g4662,
    g141,g5151,g1509,g7774,g766,g6839,g1018,g8869,g588,g9031,g1467,g8875,g317,
    g4623,g457,g4642,g486,g6357,g471,g6354,g1381,g6887,g513,g9116,g1397,g6389,
    g533,g530,g1021,g8870,g1421,g5179,g952,g8668,g1263,g5737,g580,g6368,g615,
    g6813,g1257,g5738,g46,g8955,g402,g6343,g998,g1005,g1041,g7765,g297,g6324,
    g954,g8670,g105,g145,g5152,g212,g4601,g1368,g6874,g232,g4606,g990,g7516,
    g475,g4645,g33,g5184,g951,g8667,g799,g7756,g812,g7758,g567,g6367,g313,
    g4619,g333,g6334,g168,g7742,g214,g4603,g234,g4608,g652,g1126,g8674,g1400,
    g6390,g1326,g7306,g92,g6794,g309,g6328,g211,g4600,g834,g2650,g231,g4605,
    g557,g6366,g1383,g6889,g1220,g6378,g158,g7740,g627,g6825,g661,g7743,g77,
    g6777,g831,g2651,g1327,g7307,g293,g4614,g1146,g1612,g89,g150,g7738,g773,
    g6847,g859,g8221,g1240,g1235,g518,g6361,g1472,g8960,g1443,g4667,g436,g4638,
    g405,g6344,g1034,g8957,g1147,g374,g4627,g98,g5146,g563,g9029,g510,g9115,
    g3842,g215,g4604,g235,g4609,g1013,g6,g9374,g55,g7733,g1317,g5743,g504,
    g9113,g665,g7744,g544,g6365,g371,g368,g62,g7509,g792,g5162,g468,g6353,g815,
    g7760,g1460,g4668,g553,g9028,g623,g6822,g501,g9112,g1190,g8677,g1390,g4659,
    g74,g6776,g1156,g1081,g318,g6329,g458,g4643,g342,g9097,g1250,g7111,g1163,
    g2655,g1363,g6877,g1432,g5183,g1053,g8873,g252,g6321,g330,g6333,g264,g9090,
    g1157,g1357,g8675,g375,g4628,g68,g6774,g852,g2644,g261,g9089,g516,g4650,
    g536,g6363,g979,g7104,g778,g7296,g3832,g1292,g7302,g290,g287,g1084,g7106,
    g1439,g5182,g770,g6844,g1276,g6384,g7102,g1004,g7105,g1403,g93,g5145,g2,
    g9361,g3836,g560,g6370,g1224,g6857,g1320,g7114,g617,g6815,g316,g4622,g336,
    g9095,g933,g5166,g456,g4641,g345,g9098,g628,g6826,g8,g9376,g887,g7099,g789,
    g7297,g173,g7736,g550,g9027,g255,g9087,g949,g8665,g1244,g2659,g620,g6818,
    g1435,g5181,g477,g4647,g926,g3838,g855,g8220,g1214,g5736,g1110,g7299,g1310,
    g296,g4617,g972,g2653,g1402,g6391,g896,g613,g6820,g566,g3848,g1394,g6388,
    g1489,g7770,g883,g47,g9389,g971,g5171,g609,g6808,g103,g5157,g1254,g6381,
    g556,g3847,g1409,g5178,g626,g6824,g1229,g7110,g782,g5734,g237,g6316,g942,
    g2652,g228,g6315,g706,g7750,g746,g8956,g1462,g8678,g963,g7764,g129,g5156,
    g837,g2649,g599,g6798,g1192,g1191,g828,g7762,g1392,g6387,g492,g6359,g95,
    g94,g944,g6372,g195,g3831,g1431,g2673,g1252,g2661,g356,g6335,g953,g8669,
    g1176,g5172,g1376,g6890,g1405,g5744,g1225,g6858,g1073,g9145,g1324,g7118,
    g1069,g9134,g443,g9101,g1377,g6891,g377,g4630,g618,g6816,g602,g6800,g213,
    g4602,g233,g4607,g1199,g6375,g1399,g3861,g83,g6779,g888,g7100,g573,g9033,
    g399,g6342,g1245,g507,g9114,g547,g9026,g108,g5147,g610,g6809,g630,g6828,
    g1207,g5173,g249,g6320,g65,g4598,g936,g5168,g478,g4648,g604,g6802,g945,
    g5170,g1114,g7521,g100,g429,g9107,g809,g7511,g849,g2645,g1408,g5177,g1336,
    g6864,g601,g6799,g122,g6788,g1065,g9117,g1122,g8225,g1228,g7109,g495,g6360,
    g1322,g7116,g1230,g7300,g1033,g9034,g267,g9091,g6374,g1395,g1393,g373,
    g4626,g274,g4612,g1266,g5739,g714,g7752,g734,g7755,g1142,g8874,g1342,g7119,
    g769,g6843,g6852,g1481,g7769,g1097,g543,g3846,g1154,g1354,g7768,g489,g6358,
    g874,g4654,g121,g5154,g591,g9032,g616,g6814,g1267,g4656,g1311,g605,g6803,
    g182,g5161,g1401,g950,g8666,g1329,g2663,g408,g6345,g871,g5167,g759,g6832,
    g146,g7735,g202,g5732,g440,g6349,g476,g4646,g184,g6310,g1149,g7525,g1398,
    g210,g3834,g394,g4632,g86,g6780,g570,g9030,g275,g6322,g303,g6326,g125,
    g5155,g181,g5160,g6393,g595,g576,g1319,g7113,g863,g8222,g1211,g5174,g8223,
    g1186,g1386,g6884,g875,g5165,g1170,g1370,g6876,g201,g1325,g7305,g1280,
    g7112,g1106,g7107,g1061,g9035,g1387,g6885,g762,g6835,g1461,g4669,g378,
    g6337,g1514,g7775,g1345,g7528,g6373,g1391,g185,g4599,g1307,g3858,g1159,
    g1223,g6379,g446,g9102,g1416,g4665,g395,g4633,g764,g6837,g1251,g6860,g216,
    g6311,g236,g4610,g205,g3835,g540,g6364,g3849,g1537,g7777,g727,g8228,g999,
    g8865,g761,g6834,g1272,g6383,g1243,g2660,g1328,g7309,g1130,g7522,g1330,
    g6862,g114,g6786,g134,g6791,g1166,g1167,g524,g9109,g1366,g6866,g348,g9099,
    g1148,g1348,g7529,g1260,g6382,g7,g9375,g258,g9088,g521,g6362,g300,g6325,
    g765,g6838,g1118,g7766,g1318,g6861,g1367,g6873,g677,g7747,g376,g4629,g1057,
    g8959,g973,g8672,g2664,g1549,g7780,g1321,g7115,g1253,g5741,g1519,g8227,
    g584,g6369,g539,g3845,g324,g6331,g432,g9108,g1158,g321,g6330,g414,g6347,
    g1374,g6872,g6782,g1284,g7301,g1545,g7779,g1380,g6886,g673,g7746,g607,
    g6805,g306,g6327,g943,g8671,g162,g7741,g411,g6346,g866,g5163,g1300,g7303,
    g384,g6339,g339,g9096,g459,g6350,g1323,g7117,g381,g6338,g1528,g7776,g1351,
    g7530,g597,g6796,g1372,g6870,g154,g7739,g435,g4637,g970,g1134,g7523,g995,
    g7517,g190,g1313,g5742,g603,g6801,g1494,g7771,g462,g6351,g1360,g8676,g1450,
    g5186,g187,g5730,g1179,g1379,g6879,g12,g8662,g71,g6775,g1658,g1777,I9325,
    g4242,I7758,g2605,g5652,I10135,I13502,g7135,I12558,g3880,g2965,I12382,
    I15824,g9157,g5843,g5367,I6112,g7189,I13109,g8970,I15414,I6267,g6062,
    I10675,I16126,g9354,I10519,g5242,I15181,g8734,I11443,g6038,I12436,g6635,
    g5662,g2547,I6371,I7365,g3061,I10154,g5109,g1611,I11278,g5780,g7171,g7071,
    I14154,g7558,I12274,g6672,I14451,g5834,I10525,g5971,I10587,g3978,g3160,
    I6676,g1603,g3612,I7082,I8520,g3652,g2892,g2266,I13469,g7123,I12346,g6737,
    I9636,g4802,I14637,g8012,I12235,g1799,I5657,g3935,I7602,I5933,g9207,g9197,
    I13039,g6961,I15426,g8895,g5598,g4938,g1674,g7281,I13277,g3982,g3192,I8913,
    I15190,g8685,g2945,g2364,g5121,I9515,g3128,I6839,g3629,g2424,I13323,g5670,
    I10157,I11815,g6169,I12397,I6849,I15654,g8789,g8564,g3542,I12292,g6657,
    I11221,g2709,g1747,I11677,g6076,I11503,I8859,I8829,g4029,I15546,g9007,
    g1680,I5515,I15211,g8808,g2340,I12409,g6398,I8880,I14106,g7138,I12996,
    I6703,g1983,g5938,g5412,g8771,g2478,g5813,I10472,g7338,I13432,g2907,g2289,
    g1744,g9215,I15921,I12915,I12433,I12635,g6509,I13359,g1802,I10439,g5214,
    g2959,g1926,I14728,g8152,I8733,g3996,I14439,g8063,g2517,I6348,g4010,g3097,
    I7662,g3642,I9446,g3926,I8974,g3871,I10277,g5519,I9929,I15732,g1558,I5435,
    I7290,g2936,g2876,g2231,I16058,I11884,g6091,I9145,g4264,I6468,g1917,g5606,
    g4748,I8796,g3934,I14148,I14349,g7588,I11410,g5845,I12164,g5847,g695,I5392,
    g6708,g6250,I13410,g7274,I15625,g9000,g6520,I11704,g1901,I5781,g6219,
    I10998,g6640,I11908,I8980,g4535,g3902,I7495,I12891,g6950,I11479,g6201,
    I11666,g5772,I10190,g2915,I6643,I13666,g7238,g6252,g5418,I12307,I8357,
    g7049,I12813,g3512,g1616,I13478,g7126,g5586,g6958,I12675,I15943,g9214,
    I8769,I6716,g1721,I11455,I8916,I5981,I8177,g2810,I7847,g3798,I16055,g9291,
    g9336,I16084,g2310,I6087,g7715,I14022,g1600,g1574,g1864,g4566,g2902,I11556,
    g6065,g7098,g6525,I5997,I12358,g7498,I13672,I6460,I12108,g5939,g6765,g3529,
    g2323,I15391,I6198,g4693,I13580,g7208,g4134,g3676,g3649,I14139,g7548,I9416,
    g4273,I12283,g6692,g8482,g8094,g5525,g4934,I7356,g5645,I5353,g3833,g2402,
    I7950,g2774,g2824,g1688,g1580,g2236,I5969,g7584,I13897,g4555,g2894,g9065,
    I15589,I9642,g4788,g7539,I13797,I15411,g8897,I15527,g9020,I10415,g5397,
    I13084,g9322,g9313,g3964,g4792,I9111,g9230,I15950,g6225,I11014,I8781,g3932,
    I8898,g4089,g6073,g5384,g2877,g2232,I12259,g1736,I5577,I12091,g5988,I8778,
    g5607,I15513,g7162,I13060,g7268,I13244,g7019,I12771,I11740,g6136,g7362,
    I9600,I13740,g7364,I9654,I15894,g9195,I11299,I7723,g3052,g4113,g6069,
    I10690,g2556,g1889,I7101,I5901,g2222,I5939,I13676,g7256,I15678,I8291,
    I13373,g7270,g2928,g2326,g4202,I14783,I7605,g2752,I15714,g9077,g5587,g2930,
    g2328,I15315,g8738,I11800,g6164,I5754,g4908,g4088,I11458,g6206,g5639,g5311,
    g2899,g2272,I15871,g4094,I7905,I11936,g5918,g3872,g2954,I15202,g8797,I7132,
    g4567,g2903,g7728,I14055,g7486,I13646,g3843,I7332,g3989,g3131,I6186,I14061,
    I9612,g4776,I10608,g5701,I9648,g8762,g8585,I13692,I15978,g9235,I14115,
    g7563,g7185,I13099,I9081,I7041,g2401,I12418,I9935,g4812,g4593,g2939,I11964,
    g3549,g2404,I7305,g3971,I7688,g7070,g6562,g2295,I14052,g7494,g2237,I5972,
    g7470,g7253,I15741,g9083,g8657,I14763,I12214,I13550,I9666,I6574,I8215,
    g3577,g6898,I12567,g1838,g5591,g4841,g6900,I12571,I14445,I8886,g4308,g5832,
    I14813,g8640,g1795,I5649,I12262,g1737,g2394,I6270,g9248,g1809,I10973,g5726,
    I14798,g8605,g6245,g5690,g4360,I8333,I7368,g3018,g9255,I15985,g9081,I15635,
    I12948,g6919,I13909,g7339,I15735,g9078,g4521,g2866,I14184,g7726,g1672,
    I14674,g7788,g8464,g8039,I11200,I12702,g6497,g2557,g4050,g3080,I8838,
    I12757,g6577,I15681,g2966,g1856,g5794,I10421,I5889,g1643,I11569,g6279,
    g7131,g6976,I11359,g2471,I6309,g7006,I12748,g7331,I13413,I15196,g8778,
    I6636,g1704,I14732,g8155,g2242,I10962,g3909,I7520,I11747,g6123,I12564,
    g6720,g8563,I14662,g2948,g2366,I11242,g6183,I14169,I12328,I12903,g3519,
    g2185,I10761,g5302,I13347,I7856,g3805,I7734,g2595,g2955,g7487,I13649,g5628,
    g1742,g6088,I10708,I12427,g5515,g4923,g6764,g6488,I11652,I8889,g4777,I9084,
    I10400,g5201,g5100,I9484,I9512,g3985,I13807,g7320,I11974,g5956,I12062,
    I14400,g7677,g2350,I6166,I15726,I14136,g9218,I15930,I9823,g5138,I16052,
    g2038,g4882,g4069,I14214,g7576,I12933,g7018,I9366,g4350,g7226,g6937,I11230,
    g6140,I11293,g5824,I10207,g5075,I13293,g7159,I12508,g6593,I11638,I12529,
    I6446,g1812,I8748,I5356,I14005,g7434,g7045,g6490,I11416,g5829,I10538,g5255,
    I6003,I9148,g4354,I13416,g7165,I5795,g9129,I15765,g2769,g7173,g6980,g9329,
    g9317,I11269,g7091,g7491,I13653,I12481,I7383,g2918,g3341,I6936,I5839,g6650,
    g6213,g7169,I13075,I13281,g1572,I15379,I6695,g2246,g4541,g2883,g7059,g6538,
    g7920,I14282,g7578,I13879,g6008,I11835,g6181,g3691,I7195,g5621,g7459,
    I13617,g9221,I15937,I12205,I9463,g3942,g7718,I14031,I14172,g4153,I8024,
    g4680,I8945,g3650,I10773,g4353,g3665,I11586,g6256,I12912,I11335,I14100,
    g7580,I6223,g8038,g7694,g6768,I12173,g4306,g7582,I13891,g6594,I11796,g1961,
    g3879,g2963,I9129,g7261,I13225,I14683,g7825,g3962,I9579,g7793,I14234,g3158,
    I6853,g3659,g2293,I12289,g5648,I6416,g1794,g3506,g1781,g7015,I12763,I12592,
    g4558,g2897,g9068,I15598,I7126,g2494,I5926,I7400,g3075,g3968,I7326,g2940,
    I6115,I6251,g2921,g2312,I10684,I12532,g6122,I10752,I10882,g5600,g6228,
    I11021,g3587,g1964,I11275,g5768,I9457,g3940,g8918,I15340,I16180,g9387,
    g6230,I11025,g7246,I13196,g8967,I15405,I13746,g7311,I13493,g7132,I9393,
    g4266,g4511,g2841,I15660,g9062,g2895,g2268,g6033,g2837,g1780,g7721,g7344,
    g5839,I10532,I9834,g4782,g4092,I7899,I13035,g6964,I7712,I12731,g6579,
    I11806,g6275,I8715,g3465,g4574,g3466,g6096,g5317,g6496,I11662,g1679,I5512,
    I8097,g3237,g5278,I9794,I12406,g7502,I13682,I15550,g9008,g9198,g9187,g3545,
    g2344,I8354,g738,I5404,g6195,I10940,g5618,g5015,g6137,I10776,I12544,I9555,
    g1831,I11338,g3591,g1789,I7299,g4580,g2919,g9241,I15971,I7588,g2584,g3853,
    I7362,I14725,g8145,g7188,I13106,I10592,g2842,g2209,I9938,g4878,I10758,
    g1805,I5667,g1916,g5693,I10204,g7216,I13152,g1749,g2298,I6072,I14082,
    I12448,g2392,I13193,g7007,g2485,I11362,g5821,g7028,I13362,g7265,g3931,
    I7592,I8218,g3002,I15773,g9126,I6629,g2052,I8784,g7247,I13199,I5654,I6130,
    g4076,I7859,g9319,g9309,g5489,g2941,g2349,I9606,g4687,I11353,g3905,I13475,
    g7125,I14848,g8625,g6255,I11066,I12316,I10804,g5526,I6800,g2016,I9687,
    g4822,g3630,I7095,g6481,I11641,I14804,I14094,I8868,g5113,I9499,I12008,
    g6097,g5345,I11437,g5801,I15839,g9168,g2520,g9209,g2640,g1584,g9211,I15909,
    I11389,g4285,I8233,I8727,g3944,g9186,I15836,I5679,g4500,g2832,I16176,g6960,
    I12681,I15965,g9219,I7944,g3774,g1579,g703,g1869,g4960,I13356,I11347,g5761,
    g2958,g2377,g7224,I15492,I5831,g2376,I6226,g5494,I9918,g3750,g2177,I9570,
    g4696,I10406,g5203,I9341,g4251,g5719,g1752,I14406,g7681,g3973,I9525,g4413,
    I11781,g6284,I12768,g6718,I15619,g8998,g9370,I16138,I9645,g4900,I15557,
    g9010,g2829,g1785,g9125,I15753,g4024,I11236,g6148,g2286,I6042,I12220,
    I14145,g7066,I12839,I10500,g5234,I16168,g9381,g7589,I13912,I6090,g2911,
    g2292,g4795,I9116,I8932,g4096,I5422,g7466,I13622,g4809,g6267,I11086,I11263,
    g3969,I14049,g7493,I16006,I11821,g6170,I12881,g6478,g1786,g7365,I13509,
    I12810,I7347,g2985,I15641,g2270,I6015,g4477,I8517,g7448,I13605,I13063,
    g6973,g7711,I14012,g4523,g2868,g6676,I11984,I11790,g6282,I11206,I13264,
    g7061,I6148,g7055,g6517,I14436,I8844,g3666,g2134,I9158,g4256,I13137,g7027,
    g2225,I5948,g6129,g7455,I13613,I11314,g6761,I12154,g2073,g7133,I12983,
    I7697,I15708,g7333,I13419,I13873,g7342,g9306,I16036,I12355,g1770,I14193,
    g5521,g4929,I15388,I12361,I8817,g3648,g3875,g2324,g3530,g4232,g7196,I13122,
    g4742,I9064,g9061,I15577,I15601,g8992,g4104,I7925,I10605,g5440,I11422,
    g5842,g6592,g3655,g1844,I15187,g8682,I14273,g7631,I11209,g6139,I13422,
    g7586,I13209,g6912,g2540,I9615,g4739,g6221,I11004,I12003,g6202,g8765,g8524,
    g7538,I13794,I13834,I6463,g1769,I10463,g5220,g9324,I14211,I15495,g5724,
    g4969,I6229,I14463,g8072,I12779,g6740,I9663,g6703,I12041,I13707,g4926,
    g9212,g9200,g9189,g5627,g7614,g3884,I7417,g3839,I7320,g2287,I6045,g7067,
    g6658,g8974,I7317,g2893,g5658,I15791,g9140,g7418,I13533,g6624,I11864,g7467,
    g7236,g6953,g6745,I6118,I14795,g8604,I14454,g5835,I10528,I13302,I8754,
    g6068,I10687,g1888,I6872,g4044,g6468,I11622,I12945,I9591,g4710,g4444,I8452,
    g1787,I6652,I11607,g5767,I6057,I12826,g6441,I12999,g7029,I11320,g5797,
    I15666,g9070,I13320,g7139,I6457,g1886,I13659,g1675,g6677,I11987,g7058,
    I13274,g6917,I7775,g3705,g5611,g8324,I14573,g4572,g2909,I7922,g3462,g2898,
    g2271,I15478,g8910,g2900,g2273,I12469,I12672,g6473,I7581,I15711,g4543,
    g2885,g5208,I11464,g5799,I10436,I13565,g7181,g4778,I6834,g9307,g9300,g2510,
    g639,I5374,g2245,g6149,I10810,g3988,I6686,I11374,g5674,g5042,g8177,I14410,
    g3693,I11034,g5644,g9223,I14163,g7533,g2291,g7438,I12415,I15580,g8985,
    I12331,g6704,g5541,g4814,g3548,g1684,g1745,g6198,g5335,g1639,I11515,I10541,
    g5256,I6121,g7263,I13231,g2207,I5920,I9585,g5680,g5101,I12897,g6962,g6569,
    I12961,g6921,g4301,I9630,g4867,I14789,g8544,g2259,g4014,I7769,I7079,g2532,
    I12505,g6612,g9315,I16061,g1808,g4885,g4070,I13635,g7243,I10289,g8199,
    I14424,g9047,I15543,g5802,I10445,I8895,g2923,I6657,I12717,g6543,g1707,
    I14325,g7713,I10829,g5224,g8781,I10535,g5254,I5389,I5706,g8898,I15308,
    g4903,g4084,g7562,I13858,I15178,g8753,I10946,g5563,I15003,g6524,I11710,
    I14828,g8639,g6644,g6208,g8510,I14643,I13164,g7086,I5371,g7723,I14042,
    I14121,g7587,g2215,I15953,I11284,g2886,g2240,g3908,I7517,I13335,g2843,
    g7336,g9057,g4036,g6152,I10815,g6258,g5427,I11383,I12325,g1575,g1865,I8483,
    g3641,I12472,g3567,g2407,I15417,g8893,g1715,I5559,g2314,I6099,I9440,I14291,
    g7680,g6632,g4335,I9123,g4455,I15334,g8800,I14124,g2870,g5492,g4919,I12148,
    g4382,I8373,g1833,g5128,I13537,g7152,g5574,I8790,g4020,g6211,g2825,I6553,
    I6434,g6186,I10919,I11485,I12646,g6493,g7585,I13900,g9017,I15475,g4931,
    I15762,g9039,I12343,g6731,g4805,I9136,g6975,I12712,g4916,g4022,I7785,g3965,
    I7676,I5963,g6599,I11809,g1896,g7441,I15423,g8894,g6026,I9528,g4006,g6426,
    I11559,I6860,g3264,I6900,I7053,g2452,I6341,I10506,g5236,g5580,g9234,I15956,
    I10028,g4825,g6614,I11838,I14028,g7501,g3933,I8904,g4126,g9330,I11302,
    I12334,g3521,g4560,I8446,g3014,g3050,I6788,I7115,g9201,g9006,I10265,g2943,
    g2362,g6984,I12725,g7168,I13072,g6939,I7731,g6287,I12412,g6404,I8841,g3979,
    g5623,I14187,g6083,I10702,g6649,I5957,g2887,g2241,g4873,I9217,I8811,g7531,
    I13773,g4095,I7908,g5076,I8763,g3947,g4037,g2845,g6483,I11645,I12229,g6659,
    I9884,g4868,g2934,g5476,g4907,g4653,I8874,I6358,g4102,I7919,g6636,I11900,
    I15568,g8981,I15747,g9042,I5865,g9213,I15915,g6106,I9651,g4579,I10649,
    g5657,I12011,I11245,I5715,I13695,g5871,I10558,g3878,g2962,g8008,g7559,
    g4719,I9021,I12241,I14073,I6587,g1708,g3777,g2170,g7411,g7202,I9372,I10491,
    g5231,I15814,g9154,I7308,I16116,g9350,I11488,I11522,g2096,I9618,I12582,
    g5285,g6461,g8768,I13663,g7235,g3882,g2970,g2496,I7626,g3632,g4917,I15974,
    I6615,g6756,I12141,g8972,I15420,I10770,g5441,I12310,g6723,g1897,g6622,
    I11858,I13628,I8757,g3921,g6027,g7992,g7557,g4265,g3611,g6427,I11562,g2137,
    g2891,g2265,I9678,I15638,g8978,g9366,g2913,g2307,I12379,g5139,I9543,I9837,
    g6904,I12958,g6920,g9056,I15562,g8065,I14338,I8315,g6446,I11591,g3981,
    I7706,g5024,I9360,g6514,I11696,I6239,g3674,I7164,g2807,g1782,I5362,g3841,
    I11326,g5819,g4892,g5795,I10424,I10268,g8917,g6403,I13326,g7176,g5809,
    I10460,I5419,I9804,I10262,g5551,I7683,g2573,g3997,I12742,g6590,I12394,
    I15510,g8969,I11040,g5299,I11948,g5897,g6763,I12158,I7778,g3019,I16142,
    I11500,I5410,g4296,g3790,g3238,I6894,I9621,g4732,g5477,g9260,I15990,g5523,
    g6469,I10719,g5559,g6637,I11903,g5643,I10128,I15014,g8607,g1801,g4553,
    g9063,I15583,I11248,I15586,g8987,I15007,g8627,g4303,I14718,g8068,g3802,
    g1832,g7688,g7406,I11404,I11008,g2481,I6317,g8913,I15329,g1748,g2692,g1671,
    g4012,I7765,I12445,I10283,I9974,g5099,g2497,I12690,g6467,g2354,I6178,
    I16165,g9377,g2960,g2381,g4706,I9005,I9567,I7526,I5897,g8179,I10247,g5266,
    g3901,I7492,g7000,g7137,I15720,g9053,g9318,g9304,g9367,I16129,I11933,
    I12968,I8935,g4005,I5425,I7800,g6251,I11060,I11272,I12304,g6642,I11912,
    I11851,g6277,g3511,g5754,g5403,I15565,g9261,I14151,I14388,g7605,I7850,
    g2795,g9193,g9181,g3092,I6826,I14777,g8511,g3492,I6970,g4281,g2562,I12493,
    g5613,I14251,g7541,g3574,g1771,g3864,g8342,g8856,g2267,I6006,I6093,g6654,
    I11942,g5444,g5074,g5269,I9791,I7702,g3062,I15684,g9067,g8481,I12128,g1578,
    g699,g1868,I5747,g4257,g3761,I10032,g1718,I5562,I14208,I12511,g4684,I8949,
    I9050,g3881,I11452,g6071,g6595,I8832,I5682,I5766,I11047,g5653,I13574,g7205,
    g2329,I6440,g1806,g7023,g9121,g4963,g4328,g2761,g1820,I5801,g9321,g9311,
    I15394,I13544,g1582,I11311,g5760,g7359,I13311,g2828,g1980,I12298,g6697,
    I6323,g7546,g1793,I7561,I10766,g2727,g4808,g6978,I11832,g7161,I13057,I5416,
    g5144,g6243,I11050,g7361,I13499,I15193,g8774,I13051,g6967,g6969,g2746,
    I12737,g6460,g2221,I5936,g3076,g7127,g6974,g8783,g7327,I13403,I12232,g6662,
    g1664,I6151,g2703,I14433,I8823,g5014,I9344,g6130,g7146,g6998,g6542,I11718,
    I11317,g7346,I13454,g7633,I13962,I5565,I11350,g5763,g2953,I7970,g3557,
    I13350,g7223,g8901,g2932,I9271,g4263,g3651,I7129,I13341,I14822,g2624,g1569,
    g2373,I15222,g8834,I12271,g3285,g1689,g6966,g8761,I10451,g5216,g5223,
    I13846,g3500,g8172,I14067,I5407,I13731,I5868,g2927,g2677,I14130,I9660,
    g5679,I10172,I11413,I5718,I13704,I10976,I5535,g4584,g6568,g4539,g2881,
    g8746,I14442,g4677,g5831,I10516,g2149,I5894,I6163,I12499,g6597,g7043,g9141,
    I9672,g5576,g6736,I9132,g4284,I6143,I9209,g4349,I12936,I7987,g3528,g5805,
    I10448,g5916,g5022,g4438,g2699,g4019,g6090,g5529,g4362,I11929,g6190,I12989,
    g6932,I6805,g7034,g5749,g5207,I11656,I12340,I14825,g8651,g3523,I14370,
    g7603,I11425,I12722,g6611,g7565,I13865,g2961,I5664,g3643,g2453,I12924,
    g6983,I13583,g7252,I5984,g1564,g642,g7147,I16122,g9353,I10151,g5007,g7347,
    I13457,I15516,g8977,I9558,g4597,g5798,I10433,g7555,g1826,g6663,g7545,
    I10807,I14996,I11371,I8989,g4537,I13779,g3634,I7107,I8193,g3547,g6155,
    I10826,I14844,g8641,I12424,I11392,I11787,g6273,I14394,g7536,I12753,g6445,
    g8866,I15184,g7210,I13144,g3499,I8971,g4464,I12145,g1638,g5796,I7738,g3038,
    g5873,g7164,g5037,I15723,I12199,g6475,g7013,I16049,g5437,g5041,I11827,
    g6231,g7413,I13524,I13743,g7454,g5028,I14420,g7554,I15208,g8810,g2818,
    g1792,g6063,I10678,g6628,g2867,g3754,g2543,g4698,g8198,g8747,g8545,g4025,
    I7792,I14318,g7657,I10236,I12696,g6503,I16148,I14227,g7552,I5689,I7959,
    g2793,g1758,g1589,I14025,g7500,g3578,I11803,g6280,g2470,g9069,I12939,
    I11132,g5917,g7317,I13383,I14058,g7544,g6254,I5428,g6118,g5549,g6167,
    I10862,I11281,g1571,g3983,I11428,g9180,I12487,g7601,g7450,I15607,g8994,
    g9380,g9379,I7389,I9396,g1711,I5555,g2274,g6652,I12161,g4678,g3712,g1952,
    g7855,I12400,I15530,g5786,I10403,I7749,g1827,g2614,g1562,I15484,I14196,
    I11506,I8820,g5364,g5124,g8980,g2325,g2821,I10377,g5188,g1774,I5616,I12708,
    g6482,g7581,I13888,I10739,g5572,g4087,I7882,g4105,I7928,I9076,g5054,g4457,
    I12373,g4801,I9126,I9889,g4819,I14739,g8173,g2348,g3961,g7060,I11890,g6135,
    g1803,g7460,g7172,I6160,g5725,g4465,I11482,g6117,g6598,g3927,I7584,I5609,
    I12244,g6098,I13710,g7340,g2636,I14088,I6767,I11290,g4226,g8386,g8014,
    I5883,g2106,g8975,I15429,g3946,g2306,I6075,I15408,g8896,g8976,g6625,I11867,
    g1662,g2790,g7937,I14285,I7762,g3029,g6607,g6232,I11031,I11778,g6180,g3903,
    I7498,I15690,I12068,I10427,g5210,g7479,I16026,I9850,I10366,g5715,g6253,
    g6938,I14427,g7835,I5466,I13314,I8360,g3513,I9139,g4364,g7190,I13112,g2622,
    g1568,I11945,g5874,I12337,g6724,I5365,I5861,I11356,g7221,g1816,I9639,I8721,
    I13679,I11380,g5822,g5202,g5787,g4007,I7752,g2904,I14403,g7679,g7156,
    I13042,I10582,g6552,I11722,g7356,I13484,g4920,g6606,I11824,g4578,g2917,
    I11090,g2873,I11998,I14657,I7296,I11233,g6147,g2514,g4718,I9018,g8483,
    I8962,I7064,g2458,I11672,g1847,g4803,g9075,g7242,g3743,g2403,g8636,g1685,
    I5528,g2145,g6687,g2345,g2208,g7704,I14001,g4582,g2922,g3916,I7545,g9323,
    g6586,g8790,g2695,g4015,g2637,g1581,I11449,I12918,I10183,g8061,I14330,
    I10292,g8971,I14127,g7594,g7163,I7640,I11897,g6141,I6078,I11961,g7032,
    g2536,I9493,g7354,g8756,g1757,g5309,g7432,I13559,I10786,I12451,g2359,I8907,
    g3560,g2361,g9351,I16103,g2223,I5942,I7844,g3784,I15982,g9236,g5808,I10457,
    g636,I6680,g6645,I11917,I16040,g9285,g4721,I9025,I14103,I11212,g6146,I5852,
    g5759,I10350,g8514,g8040,g3873,g2956,g3095,I6831,g3495,g3653,g2459,I8180,
    I12322,g6751,I14381,g2522,I14181,g7725,g7157,I13045,g2642,g1588,g3936,
    g7357,I13487,g3579,g1929,g3869,I12687,I8853,g4034,I11955,I11401,g6506,
    I11680,g1751,I5847,I12561,g6449,I16183,g9388,g5604,I12295,g6693,g3917,
    I7548,g4670,g1585,g724,g4689,I8966,g6587,I15522,g9018,I15663,g9066,I14190,
    g4279,g6111,g5453,I14448,I11260,g5833,I10522,I7814,g7245,I15959,g4028,
    I7797,g2880,g2234,I7350,g2971,I6864,g2528,I11971,g6179,g4030,g8016,I14311,
    g8757,g5584,g1673,g7712,I15776,I15553,g9009,I13369,I6021,g4564,I8665,
    I11368,g8642,I12364,g6714,g3770,g2551,g5268,I9788,I9014,g5362,I10497,g5233,
    I15536,g9004,g1772,I11467,g4806,g6591,I15702,g9064,I13850,g7328,I12367,
    I5817,g2982,g1848,g3532,I7967,g2787,I14205,g1743,I12430,g2128,g2629,g6020,
    I6127,I10987,g5609,g6702,I5605,I10250,I14076,I8742,g6507,I11683,I8277,
    g1011,I5413,I13228,g6892,I15729,I12253,g6729,I11011,I5751,g5086,I9460,
    g8880,I15218,g3189,I13716,g7475,I13631,I16072,g9303,g3990,g2554,I6376,
    I9681,g4589,I10969,I15672,g7627,I13956,g3888,I15062,g8632,g6905,I12586,
    I13308,g3787,g1842,g8017,g7692,I11880,I15933,g9210,I13758,g5470,g4899,
    I10569,g3956,g5025,I9363,g6515,g6125,I11627,g6630,g4571,g2908,g3675,I7167,
    I12976,g6928,g1573,g1863,I11227,g7021,I13940,I11958,g7039,I9422,I8351,
    I14489,g3811,g2285,g7439,I12643,g6501,I5368,I11386,g5764,I5772,g2490,I6326,
    I6024,I5531,I12669,g6477,g7583,I13894,g7702,I13997,g4196,I10169,I6795,
    g1683,I10503,g5235,g3684,g2180,g3639,g5006,I9333,g3338,I15010,g3963,I7672,
    I15574,g8983,g4538,g2148,I15205,g8809,I6431,g4780,I9089,g1857,I7788,g9050,
    I10177,g5766,I10373,g5087,g1976,I15912,I9095,g4283,I10442,g3808,g7276,
    g5487,I9907,I14315,g7676,g1970,I11793,g6188,I13428,g7167,g3707,g2226,
    I11296,I14819,g8647,I8901,g2698,g4018,I14202,g7708,I8172,g3524,I14257,
    g7716,g4713,g2964,g7495,I16020,g9264,I16161,I7392,g3230,g5755,I15592,g8989,
    I15756,I13761,I14070,g7714,g3957,g6617,I9752,g4705,g4093,I7902,g8512,I8282,
    g3515,I16046,g9288,g1760,g4493,I8543,I11926,I12496,I13822,g3865,g2944,
    I10384,g5193,g6655,g5445,g5059,g3604,I13317,g7211,g5491,g4918,g3498,g7550,
    g7593,g4381,g8649,I14743,g6010,I7302,I11129,g2872,I6590,g1924,I9633,g4685,
    I8952,g4197,I10801,g5463,g6410,I11533,g2734,g4021,I9336,g6968,I14801,g8608,
    g1779,g2057,I12124,I12678,g6516,I12523,I6571,g7120,I9419,I12388,g2457,
    g5578,g5868,I10555,I13388,g2989,g1843,g3539,g3896,I7473,g6143,g5459,I14019,
    g7480,g2393,g5718,I12460,g6674,g7022,I11323,g1977,g7145,g7534,I13299,
    I14695,g7277,I13267,g2834,I6564,I6723,g7220,I14334,g5582,g8902,g6278,g8463,
    g2686,g1667,g7789,I14224,g5261,g2007,I15770,g5793,I10418,I12065,I8202,
    g9332,g6618,g6003,g1665,I10796,I13728,g4562,g6235,I9347,g9199,I16107,I7911,
    g2767,g5218,I8094,g2976,I14457,g8093,g6566,I8808,I13737,g7446,I5359,g8986,
    I13329,I8190,g6134,g5428,g8619,g7547,I13825,I11329,I8264,g5246,I9760,g2625,
    g1570,I8730,g3086,g1852,g2253,g2938,g2347,g3728,g2202,g7433,I13261,g7041,
    g5748,g6555,I11729,g3546,I6946,g1887,I10256,g5401,I12247,I11512,g1732,
    I9675,g4807,I13512,g2969,I5383,I10280,g5488,I14085,g4585,g2925,g6621,
    I11855,g3897,g4041,I11266,g7078,g6683,I13438,I7377,I13831,g7322,I6036,
    I14157,I12277,g6681,g4673,I8928,I10949,I9684,g4813,g7035,g7134,I15803,
    g9148,I7287,g2561,g6094,I10716,I14231,g7566,g4779,I8922,g1565,g649,I8724,
    g5671,I10160,I12782,g6463,I13722,g7442,I16090,g3635,g1949,I13924,I5633,
    g1681,I7781,I6422,g4890,g4075,I12352,g6752,g7280,g2525,I6354,g3801,I7262,
    g7834,I13271,I6419,I8835,g3954,g5826,g6572,g8606,I12170,g4011,I11461,g9076,
    I15622,I5732,g6264,g7310,I13031,g5638,I11407,g2879,I6597,g7025,I11736,
    I11887,I16151,I7344,g2382,g8633,I8799,g3951,g1655,g6050,I12167,g2506,I6437,
    g1784,g6944,I6302,g3091,I13843,g7326,g9267,g3491,g1800,g4080,I7867,g7577,
    g4573,I11764,g6056,g5758,I10347,I13764,I12088,I11365,g2275,g2311,I9539,
    I10896,I13365,g7267,g5466,I10243,g5026,g5624,g7590,I13915,g9184,I15830,
    I13869,g2615,g1563,g4569,g2906,g3920,I12022,g3868,g2174,I11194,I12202,
    I8802,g6224,g2374,I6220,g5448,g5137,g1922,I9162,g4272,g7556,I13161,g7080,
    g5708,g5055,I12313,g6730,I12376,I6733,g5471,g5827,g6585,I12517,I15651,
    g3582,g2284,I5914,g7095,g7064,I12829,g2239,I5978,I7314,g2916,I10180,g9368,
    g1597,g5846,g2380,I6242,I13258,g6907,I12900,g6947,I7870,g2827,g4122,g2184,
    I12466,g5396,g4692,I5636,I12268,I6054,g2020,I5855,I10930,I11043,I6454,
    I12101,I6770,g1590,I11978,g7033,I13861,g8111,I14374,I10387,g4000,I10694,
    I7981,I10965,g6997,g2794,I11069,I15687,I6532,g1694,g9298,g2931,I6669,g3721,
    I7211,g6238,g5027,I13810,g7312,g8174,I15717,g9051,g5467,g4891,g4462,g7194,
    I13118,g7332,I9425,g655,g2905,I6012,g6744,I14064,g8284,I14531,g2628,g3502,
    g7905,I6189,g2630,g5493,g8180,g7719,I14279,g7700,I8739,g4924,I5775,g7966,
    g2100,I7623,I10469,g5222,I11967,I11994,g7471,g7233,g9044,g1942,I6029,g4023,
    I8736,g4008,I10286,I5548,I9669,I15433,g8911,I10552,I6956,g1907,g6901,
    I14039,g7449,g4588,g2929,g5872,g5685,I10186,g5197,I13425,g7166,g4311,g6511,
    I11693,I5398,I15811,g9151,I12454,g6581,g2973,g1854,I5676,g3430,I8910,g4051,
    g3093,g6092,I13918,g9233,I8871,g7150,g6952,I14677,g7791,g7350,I13466,
    I12463,I13444,g7282,g4146,I8011,g7009,I8814,I10937,g5560,I6963,g658,I6109,
    I6791,g1967,g4103,g6721,I8268,I7807,g3910,I7523,I12238,I14178,g2804,I8983,
    g1912,g5631,g7836,I14260,g5723,I9034,g4259,g6772,g3837,g7697,g2351,I6428,
    g3967,I12176,g6510,g8750,I10479,g5227,I12699,g8973,I9369,g7229,g6623,
    I11861,g7993,I14298,I7255,g1955,g5287,I14015,g7440,I9407,I12538,I13656,
    g7228,g3589,I7061,g7699,g5788,g4443,I8449,I13353,g7231,I8477,g9178,I16158,
    g7031,g4116,I12484,I5954,g2884,g2238,I7386,g3048,I6784,I7811,I9582,g4694,
    I8205,g6651,g9182,I5432,g4565,g2901,I14792,g9382,g9217,g8882,g3919,g2372,
    I6214,g7248,I5568,I7341,g2618,g1566,g9355,g2235,I5966,g2343,I10780,I12439,
    g4697,I8986,I11344,g4914,g8178,g2282,I7112,g2546,g1778,g5058,I12385,g4596,
    g3911,g6024,g4013,I12256,g3780,g5129,I12111,g2334,I8273,I12349,g6742,g5722,
    g2548,I7293,I12906,g6918,g8899,g2495,I13023,g7040,g1661,I7329,g2920,I11224,
    g2555,I11028,I11308,g1796,g6711,I15675,I10259,g6523,I11707,I9502,g3972,
    g3994,g4536,I15696,g9208,g9302,g9281,I8862,g6205,I14397,g9074,g2621,g1567,
    I8712,g2712,g1686,I6728,g1959,g5474,g4904,g1646,I8718,I7746,g6634,I11894,
    I13816,g8235,I14492,g2313,I6096,I12120,I5471,g6104,I14964,g8406,I11239,
    I15504,I12138,g4922,g4111,g5439,I13752,g7315,g5844,g2290,g5480,g4913,I6425,
    g1811,g5713,g4581,g3700,I7953,g6754,I12135,g1583,g5569,I8706,I9564,g4703,
    I11669,I13669,g7240,g8792,g5779,g6613,g3950,g4784,g5417,I9053,g5800,I9910,
    g4681,g5688,I10193,I15533,g9002,g2384,I5478,I14747,g8175,I5475,I7716,
    I12457,g4079,I7864,I11525,g6034,g7177,g3562,I7044,I9609,g2264,g6712,g7405,
    I13518,I8919,I6305,g3631,I7098,g7829,g2360,g2933,I6673,g3723,I12609,g6571,
    I13290,I14166,I7198,g2509,g5294,g5000,I5646,g7705,I14807,g8603,g2641,g1587,
    I14974,g8442,I10639,g4501,g2801,g6263,I12684,g3605,g1938,g2996,g1828,I9466,
    g3943,I10353,I15845,I12921,g6993,I13713,g7341,I13250,I8805,g3976,g5468,
    g4195,g1925,g8776,g2724,g1814,g7225,g6936,g7610,I15501,g6014,I10614,I14416,
    g7727,g2379,I13610,g7227,I16145,I12526,g4704,I9001,g6963,g6660,g6946,
    I12649,I13255,g7057,g2878,g2233,I13189,g7002,I7644,g7259,g7124,g6896,
    I12973,g6927,g5608,g4245,I6051,g6903,g2777,g1797,I16009,I10579,g5433,I9774,
    g4250,g2882,I11686,I11939,g6015,I16017,I13460,g4032,I6018,g7275,g7206,
    I13134,I6578,I6868,g6036,I10643,g6913,g1933,I16132,g9356,g5215,I15498,
    g1987,I5842,g4568,g3013,g5665,g5051,I11332,I16043,g3531,g5127,g2674,I11191,
    I11473,g9363,g1776,I7599,I15924,g6767,g4357,g3679,I12286,g5633,g4895,
    I11218,g6161,I5975,g2332,I10430,g5211,I13837,g7324,I7371,g2680,I14430,
    g2353,g4426,g4120,g9183,g6760,g9080,g5696,g1945,I12652,I12265,g1738,g3074,
    I10253,I13305,g3992,I14035,I15199,g5258,g6087,I8793,g3588,I11470,g6095,
    g5240,g5072,g7360,g8799,I14142,g7551,g5472,I9892,g4489,I12490,g7207,I14816,
    g6037,I10646,g3573,I5789,g6102,g8541,g2511,I12478,g1876,g6735,g6064,I11494,
    I13595,g7488,g2092,g5434,g5112,I11037,g7592,g7532,I12131,I13782,g6246,
    g8802,I11419,g1818,g9019,I15481,I7374,g7951,I14288,g3828,I15225,g8689,
    g9072,I10475,I9301,g4295,I12930,I7145,g2501,I5945,I8787,g4475,g3818,g5596,
    g1663,g7870,I14270,g5013,I5709,I14646,I15648,I11215,g2480,g2623,g6725,
    g5706,g5820,I10485,I7359,g2871,g9185,I15833,I7875,g7151,I15657,g9059,g9385,
    I16173,I15068,g8638,I14175,g1877,g5828,g6553,I11725,I15604,I13927,I8745,
    g3929,g2375,g6565,g3220,I15337,I6217,g6012,g1556,g7068,g3779,g4583,g2924,
    g5753,I6039,g6189,g4909,I13749,g7313,g7887,g7122,g3977,I12535,I6048,g5241,
    g5581,I14264,g7698,I9531,g4463,I5911,I6711,g1726,I11440,g8968,I6254,g5060,
    g7352,I11305,g5807,g9331,g6956,g5460,g5597,I11254,I13562,I11981,g6285,
    g4561,g3051,I6333,I9505,g4300,g6664,I15705,g5784,I10397,g4004,g8584,I15918,
    I16033,I10274,I8865,g7496,g4527,g3999,I8856,I7595,g3633,I7104,I6471,I12993,
    g2477,g2643,g6684,g6639,g5668,I11341,g8991,I6509,g4503,I8565,g5840,I7978,
    g2205,g6773,g5190,g4925,g4114,g3732,g2533,g1557,g2634,g3753,I9573,g4701,
    g9045,I15539,g5213,I5401,I14614,g7832,g7266,I13238,g7904,g2104,I5879,I7635,
    I9594,I16023,I7629,g6759,g5524,I13009,g6935,g1948,I15065,g7142,I13012,
    g2926,g9369,I16135,I10565,g5402,g6957,g7255,I8766,g2816,I5380,I14810,g3316,
    I6930,I15571,I11476,g6194,I11596,I7554,g7097,g7497,g5577,g2044,g6604,
    I11818,g5810,I13570,g7198,g6498,g2269,g1773,I8486,I10409,g5204,g4547,g5053,
    I12370,g3987,g3533,g2397,g2862,I15631,g9003,g6682,I9250,g6173,g2039,g9227,
    I15947,g3870,g4838,I6764,g1918,I13241,I9597,g4738,g8754,g6019,I13185,g7020,
    I13092,g7047,I6663,I12514,g6605,g7141,g7129,g8982,g1822,g7329,I13407,g4035,
    I6451,g2946,g2365,I12421,g6486,I14109,g4482,I7964,g3488,g5626,I13921,g3960,
    I9588,I11648,I8105,g3339,I8883,I12098,g9188,I15842,I13157,g9071,g3922,
    g9237,g9216,I12541,g4915,g6156,g6070,g1895,g6897,g1837,I13577,g7186,g6025,
    g7596,g5683,g6755,g4800,g2288,I7118,g2484,g2505,I14091,I6248,g6556,I15669,
    g1768,g7564,I9103,g4374,g7143,g3739,g1698,I6368,I6646,g9171,g3783,g1788,
    g3995,I7728,g3937,g8903,g3079,g5782,I10393,g4002,I10390,g5195,I13906,g7358,
    I13284,g6131,I9443,I7323,g2947,g7149,g2798,g7349,I13463,g7279,g3390,I6949,
    g6766,I10705,I14413,I6856,g4590,g5243,g3501,I13126,I14112,I14267,I15927,
    g2632,g1576,g4297,I8261,g4556,g5084,g5603,g1941,I5812,I6474,g3923,g4317,
    I6443,g7241,I5923,I12760,g6685,g4928,g4119,g6226,g4930,g4121,g8916,g2869,
    g2224,I15610,g8995,g5513,g9048,I5552,g4811,g2389,I7655,I11446,g9060,g2309,
    g9333,g7319,I14904,g8629,g3918,g1958,I6000,I11434,I13472,I13876,g6007,
    I12927,g7014,g9196,g7717,g6059,I12475,g5616,g3568,g1935,g7128,I14712,I6192,
    g6457,I5960,g5200,I13147,g3912,g7686,I7888,g2454,I6294,g2826,g2770,g2210,
    I12250,I10509,g5237,g4557,g2896,I10369,g7599,I15595,g1974,I10933,g8801,
    I10617,g4071,g8752,g6227,I11018,I14851,g8630,I8161,I12965,I8428,I11055,
    I7691,I15160,g8631,I13813,g7314,g8042,g5114,I14623,g6257,g8786,g5120,g6656,
    g9177,g2706,g1821,I8826,g7483,g9194,g3941,I6183,I6608,I10574,g5426,g2371,
    g4200,g1807,I11732,g5617,g8770,g6502,g7710,g5789,I10412,g4009,I16119,g7790,
    g5516,g8990,g6940,I12639,I8308,g7187,I13103,I7311,g5987,g1849,g3778,g7343,
    I5377,g4198,I11491,I9840,g4702,g3735,g6216,g3084,I14305,g6028,I14780,g6646,
    g6671,I14276,g2639,g7046,I12806,g5825,g2216,g2383,g4229,I8140,g5707,g3949,
    I6084,I15693,g9301,I9177,g8029,I7380,g3461,g7345,I13451,g8787,g9282,I7832,
    g2768,I10271,I14160,g3526,I15382,g3998,g5709,g6741,I12117,g8988,I6820,
    g3603,g5478,g7030,I12909,g4921,I7353,g9165,g2957,I8196,g3654,I7931,g2780,
    g1923,g6108,g5435,I11251,g5517,g4258,g5482,g1701,I5545,I12520,g4327,g8684,
    g3583,g4078,g2863,I8775,g8791,I8480,g2498,g6217,g5649,g6758,g6589,I7204,
    I15616,g8997,g2833,I6561,g7251,I13203,g1830,g3952,I7651,g7811,I14238,I8994,
    I10046,g4840,I14046,g7492,g6048,I11991,g2539,I6363,g3561,g9058,I13515,
    g8759,I13882,I12059,g5841,g7271,g1825,g3527,I15385,g6133,g7709,g3647,g5052,
    g2162,I7973,g3071,I6009,I12193,I12629,g3764,g4085,I7878,I7029,g5002,I8847,
    g7595,I13930,I12280,g3503,g3970,I11714,I13441,I12211,I11689,I5670,g1943,
    g1878,I12776,g6739,I13725,g7437,g2728,g2256,g2486,g6018,g7414,I13435,g7170,
    g1934,I11197,I7648,I16154,g3819,g4031,I7804,g7130,g3617,g6093,I11744,g6120,
    g7542,g7330,I11659,I12151,I12319,g5785,g6934,g7355,I8101,g3259,g7783,g3771,
    g1853,I11848,g6159,I9782,g4720,I11398,g5823,I6060,g4286,I10482,g5228,g6700,
    g6244,g6397,I8751,g3892,I9627,g2131,g2006,g2331,g4733,I10545,I13332,g4270,
    g2635,I12659,g8881,g8683,g2105,I7667,g3945,g5452,I12025,g2487,g4358,I9603,
    I14786,g3991,g7090,g4798,I10356,g5711,g8883,g7366,I15519,g5071,g3078,g3340,
    g2474,I10380,g5705,g7056,g6631,g4540,g3590,g5672,I12044,I12085,g7456,g7174,
    I13048,I13767,g3959,g1815,g6101,g7148,I13028,g9161,g7348,g3517,g2283,g3082,
    g9383,I8772,g9220,g9205,g7155,I13481,I12301,g3876,g8131,I14378,g2091,g7273,
    g1960,g5814,g7260,I9576,g3225,I9561,g4695,g8766,g5038,I5395,g3955,I6033,
    g6504,g9358,g7197,g7463,g7239,g5009,g4344,I6286,g7792,g9073,I6299,g8984,
    g4898,g7264,g9127,I15759,I9258,g3516,g5769,I11951,g8755,g5836,g4510,g2840,
    I13234,g7720,I12942,g7367,I12632,I15699,g1676,g2015,g3640,I11431,g3124,
    I12187,I6157,I12403,g6769,I12547,I5989,g7549,I8977,g8999,g1727,g3877,g5212,
    I5692,g8602,g5194,I12226,I13979,g8407,g8013,I7885,g6616,g3657,g4112,g2721,
    g6505,g8868,g7543,g6011,g1746,I14097,g8767,g9043,g3556,I7036,I10343,g5704,
    g3928,g8582,I15738,g6074,g3930,g2502,I6337,g9316,I13541,g7209,g4886,g5716,
    g8015,g7689,I14460,g4879,g5462,g2689,g1670,g6573,I11920,I12980,g6929,I8760,
    g3563,g5205,g6713,g1677,I7658,I12888,g6948,I13828,g7321,I14133,g7574,g691,
    g1866,g2700,I7755,g5475,I7335,I13344,g5537,g4594,g2183,g1855,I12442,I13903,
    g4837,I13173,g7089,g5192,g5085,g3555,I12190,g3966,g2910,g2638,g4065,I7838,
    I14857,g9206,g3677,I14925,g8381,g3948,g4125,g2308,I6081,g7017,g7560,I13755,
    I14009,I7680,g7691,g5642,I13506,g4033,g7087,I14603,g7827,g5520,g1577,g1867,
    I9310,g4268,I7558,I10681,g5686,g5812,I10914,g7158,I6195,g6459,I13490,g6220,
    I11001,I13698,I5386,I15324,I16100,g9338,I12208,g3769,I6952,I14722,I10512,
    g5286,g4714,g1975,I9142,g6977,I7551,g1813,g5538,g6588,g9079,I10842,g2396,
    g3812,I10548,g5260,g6051,g3993,I13770,I9657,g6925,g8793,I6517,g3822,g5610,
    g9005,g5073,g5473,g4081,g6945,I13819,g1872,I9520,g7180,g6103,g7591,g2467,
    g4302,I11395,g5469,g4688,g6696,I9785,g4747,g7420,I11633,I12894,I13701,
    g5206,I13719,g7334,g6508,g6072,g6115,g7678,g1756,I6245,g6274,g8780,I7947,
    g9337,g6009,g5199,g1904,g5747,g5781,g4001,g8018,g8067,I14342,g2263,I13247,
    g6906,I12986,g6931,g8900,g6955,g7054,I11701,g8493,g8041,g5238,g3085,g2781,
    g3485,g1652,g1695,g1637,g4592,g5344,I9819,g6210,g2631,g1586,g4746,I12877,
    g8181,g6596,g2817,g9357,I8998,I12196,g6471,I13140,g6954,I9350,g8421,g5088,
    g4932,g6626,g9082,I9009,g4591,I6959,g3520,g3219,g1687,g2479,g1750,g8076,
    g3958,g7351,g6601,I12866,g8562,g4968,g4576,I15940,I13447,I14709,g6922,
    I5763,I11773,I14680,g6647,g7262,I14199,g3974,g8751,I12223,g2743,g3610,
    g2890,g5245,g5196,g7092,g7701,I15962,g2011,g5806,g3980,g6996,I13776,g4524,
    I12391,g7024,g3540,g9162,g4781,g2074,I5872,I11497,I12885,g7318,g2992,g6165,
    g4577,g2914,g5545,g6686,g3287,I6911,g8772,g1649,I15613,g8996,g4711,g8743,
    g5395,g3898,g4026,g4274,g3510,g6032,g6432,I10454,g7782,g7094,g1823,I13734,
    g4544,I11203,I5542,g7088,g3692,g3694,g8583,g4106,I15507,I7564,g6661,g9320,
    g5481,I12655,g6458,I11377,g5811,g5479,g7160,I13054,I13496,g7179,g4027,
    I5908,g7050,I7632,g6933,g5259,I11870,g5818,I14079,g7579,g6924,g4003,g4676,
    I9496,g3825,g5267,g2161,I8084,g3706,I12502,g4191,g8760,g3008,I8850,g2665,
    g6237,I9845,I10125,g5253,g2327,I6124,g3768,I10783,g5542,g6894,g7269,I13547,
    g4307,g2999,g2346,I6154,g2633,g9244,I10561,g5265,I14687,g5710,I12217,g2157,
    I10295,I15784,g4299,I15628,g9340,g7254,g5592,g7810,g6075,g4016,I12038,
    I6887,g4522,g4115,I7956,g2363,g4552,g1909,g7353,g6603,g7499,g3496,I6974,
    I8877,I7338,g2316,g6283,g5677,I10166,g7335,g3891,I8925,g3913,g3505,g4595,
    g2942,I12666,g6476,g7722,g4341,g4017,g3504,g5198,g4691,g4935,g8993,g1860,
    g8443,g6004,g7826,I11923,g4130,g4542,g3815,g7693,I13088,g9222,g7837,g3497,
    I13885,g9174,I8892,g1879,g4554,g9239,I14668,g7787,g5717,g6949,g7232,I11287,
    g7036,g7561,g5244,I10488,g5230,g9294,g5209,g7476,I8709,g7652,g5264,g3429,
    g4280,I13296,g4512,g2460,I13338,I13287,g2784,g4056,g6959,g5751,g8779,g2937,
    g5752,I13527,g7217,g2668,g8775,g3746,g5083,g7838,g7703,g5566,g8581,g6286,
    g5219,g7077,g5790,g4728,g3953,g5061,g7695,I14294,g7553,g8784,g5461,I13131,
    g7426,g5756,g6035,I11257,g5622,g6276,g5115,g7415,g4057,g3866,g7258,g3716,
    g5514,I6291,g4236,g5191,g8156,g3398,g6110,g7044,g9001,g7983,g7008,g1666,
    g4253,g6643,g5016,g5757,g3644,g8363,I10494,g5232,g7833,g5522,I10466,g2626,
    g3867,g6222,g5654,g5698,g3975,g4586,g6899,g2683,g6930,g6602,g6472,g4570,
    I15645,g4525,g7178,g2782,g5612,I13066,g2627,I14118,I9624,g7443,g6089,g7422,
    g1555,g3680,I13854,g3187,g7625,g6242,g7537,g9252,g4587,g5221,g4275,g8979,
    g3904,g3514,g7037,g6150,g1908,g2276,g9339,g4545,g2616,g5490,g7696,g3359,
    g7436,g2764,g7042,g6262,g4559,g4249,g3757,g6229,g5229,g5217,g3522,g3047,
    g8059,g6281,g3874,g6951,g2521,g2617,g7608,g7412,g7121,g6462,g6215,g8925,
    g7429,g7212,g9144,g9123,g9344,g4123,g8320,I8431,g9259,g8277,I8005,g4351,
    g8299,g6941,g6582,g4410,g8892,g8681,I7994,g5552,g4832,g8945,g6431,g4172,
    I8057,I8058,g7272,g8709,g6176,g6005,g5557,g4343,g8078,g7634,g8340,g6405,
    g4282,g7604,g1714,g5570,g1759,g8690,g4334,g8876,g8769,g6733,g3613,g4804,
    g8915,g8794,g8239,g7419,g7230,g8310,g4494,I8546,I8547,g8824,g8877,g8773,
    g6399,I9330,g9142,g9124,g8928,g5020,g4933,g4320,g8930,I8114,g8064,g4158,
    g4724,g4038,g6440,g4379,g8295,g8237,g6923,g6570,I9222,g8844,I8594,I9166,
    g8089,g7658,g8731,g4271,g5511,g8071,g7540,g8705,g4799,I8033,g8948,g5969,
    g5564,g7602,g6627,g5123,g4132,I8496,g4238,I8157,g8814,g6408,g8150,g4744,
    g3525,g8438,g6972,g5661,g7222,g8836,g4901,g4288,I9261,g6433,g8229,g9349,
    g8822,g6395,g8921,g4417,g5334,g4887,g5548,g4826,g4403,g6266,g8837,g6705,
    g8062,g8620,g8462,g9119,g9049,I8001,g9258,I8401,g4175,g4375,g5313,g4820,
    g6726,g6154,g8842,g7609,g8298,g5094,g9274,g4139,I8000,g4384,g4517,g8854,
    g8941,g4424,g6979,g5095,g5593,g4110,g6112,g5673,g4077,g6001,g5540,g6401,
    g8708,g7575,g5050,g1725,g6727,g8405,g4099,g4304,g8829,g8286,g8798,g8733,
    g8270,g8610,g9345,g4269,I8209,I8524,g8069,g4712,g4276,g6124,g9159,g9138,
    g9359,g8377,g7093,g6673,g4729,g4059,g4961,g9016,g8904,g8287,I8186,g5132,
    I9534,I9535,g8849,I7995,g9251,g4414,I8412,I8413,g3313,g4187,g8291,g3094,
    g1898,g4436,g6142,g4160,g7435,g4378,g4135,g5092,g4182,I8071,I8072,I8240,
    g9272,g8259,g5714,g8088,g8852,g8923,I8461,g6734,g4422,g8701,g9328,g6465,
    g4216,g9130,g9054,g2972,I8046,g8951,g8785,g8314,g4437,g8825,g8650,g1728,
    g8336,g6061,g5257,g8943,g6046,I8115,I8642,g8322,I10597,g8934,g9348,g6145,
    g4054,g3767,g4454,g5077,g4532,I8617,I8618,g6107,g8845,I9202,g8337,g4412,
    g5104,g6757,g9279,g4389,I8612,g6416,I8417,g9118,g9046,g4787,g6047,g8266,
    g6447,g4956,g2979,g1733,g5044,g8081,g8815,g7183,g6132,g4169,g8692,g8726,
    g4138,g4109,g4791,g4707,g4062,g6417,I8090,I8490,g4201,I8108,I8109,g8267,
    g8312,g6629,g6023,g4957,g4049,I8456,I8529,g8293,g8329,g4469,g4889,g4098,
    g6554,g5762,g8828,g8830,g8727,g5436,g6719,I8063,g8703,g8932,g6166,g8624,
    g8953,g8758,g4052,g7687,g4452,g3760,g6456,g6116,g7444,g9158,g9137,g5036,
    g4086,g4179,g4486,I8528,g8716,g7428,g4504,I8568,I8569,g4185,g9275,g4385,
    g8848,g5579,g4090,g4425,g2386,g5442,g4679,g6057,g4131,g8319,I8552,g8258,
    g6971,g6424,g8717,g7597,g7316,g7079,g8274,g4445,I8455,g4091,g4491,g8325,
    g8821,I8052,I8053,g5029,g4369,g8280,g8939,g4407,g4227,g8306,g4793,g3887,
    g8461,g8622,g4246,g3226,g8403,g8841,g5049,I8020,g8695,g8307,g9278,g4388,
    g8359,g9143,g9122,g9343,g7626,g8858,g4430,I8436,I8437,g9334,g8315,g4239,
    g6239,g5314,g5019,g2935,g7683,g4876,g8654,g6420,g4108,g4883,I8040,g4066,
    g8272,g4466,I8491,g8909,g8612,g6204,g4365,g4048,g8935,g5425,g4448,I8460,
    g4072,g8328,g4133,g4333,g8542,g8330,g4396,g9160,g9139,g6040,g5105,g7616,
    g4163,g4067,I8143,g3049,g8090,g6151,g8823,g5045,g5091,g4181,g8456,g9271,
    g4397,g8851,g4421,g8698,g8260,g6172,g9238,g8720,g4101,g8318,g8652,g8843,
    I8593,g8457,g1753,g8686,g4529,g8321,g6908,g4168,g6567,g6265,g4368,g8938,
    g8813,g5030,g4058,g3656,g4743,g3518,g8740,g6965,g6489,g4411,g8687,g6160,
    g1919,g4074,g5108,g6641,g6770,g3678,g5066,g8860,g8341,g8710,g9384,g8645,
    g8691,g5048,g9024,g8884,g8879,g8782,g8154,g8962,g8890,g6249,g1739,g8275,
    g8311,g4400,g3614,g6541,g6144,I8574,g5018,g5067,g5093,g9273,g4147,g4383,
    g4220,g8380,g8832,g4176,g4514,g8853,g7081,g4423,g3188,g5700,g4361,g8931,
    g4127,g4451,g6574,g5984,g7038,g6466,g8628,g8300,g9014,g8906,g7010,g5817,
    g4472,g8440,I8523,g5585,g4741,I8643,g6175,g4332,g5614,g8323,g9335,g4870,
    g4434,I8014,I8015,I8551,g9022,g8887,g4255,g8151,g8648,g6470,g5458,g4686,
    g3509,I8613,g8839,g9037,g8965,g4936,g4117,g8278,g7192,g7026,g8282,g5080,
    g5573,g3011,g8693,g8334,g6044,g6717,g6444,g8621,g4937,g4309,g8313,g4235,
    g4190,g4390,g5126,g9012,g8908,I8288,g4356,g9371,g9352,g6414,g8264,I8041,
    g8933,g7016,g4053,g5588,g3028,g4453,I8495,g6182,g8724,g8379,g7199,g7003,
    g6916,g6022,g5595,g8878,g8777,g6422,g8289,g8835,g8271,g8611,g5043,I8296,
    g6437,g5443,g5116,g8238,g5034,g8332,g4497,g8153,g8744,g7215,g6042,I8029,
    g8804,g6054,g4526,g6615,g2889,g7136,g5117,g8714,g9025,g8889,g4243,g1690,
    g6412,g6688,g6990,g8262,g6171,g5363,g8736,g6429,g6716,g9131,g9055,g8623,
    g7690,g7096,g8722,g7195,g5937,g5562,g5079,g4546,g5141,g8285,g9226,g6109,
    g4224,I8127,g8384,g8339,I8299,g8838,I8019,g8737,g4906,g4789,g2751,g6049,
    g8077,g8643,g6715,g5681,g5032,g5432,g3233,g3358,g9015,g8905,g8742,g8304,
    g8926,g6162,g6268,g7001,g3722,g8273,g6419,g6052,g8269,g4959,I8006,g4435,
    g4690,g4082,g8712,g8543,g8729,g8961,g8885,g9247,g8927,I8045,g5894,g8660,
    g8147,g8946,g7503,g6006,g5575,g3260,g3221,g8513,g6406,g3190,g6105,g4877,
    g8378,g6487,g5750,g8335,g8831,g8288,g8382,g5484,g5096,g8749,g4785,g1678,
    g6045,g5583,g1775,g5712,g8947,g6407,g6578,g6218,g4194,I8089,g8653,g4394,
    g8302,g6600,g8719,g3986,g6415,g5970,g5605,I8028,g8265,g4955,g4254,g4150,
    g2949,g9021,g8886,g8296,g4409,g8725,g6689,g6698,g5547,g1819,g7427,I8589,
    g6428,g6430,g8281,g5078,g6638,g8297,g5082,g8745,g8338,g8963,g8891,g2986,
    g7416,g7140,g8309,I8418,g6448,g6055,g5239,g7654,g4142,g4192,g4392,g6196,
    g4927,g5615,g6396,g8715,g7363,g8833,g6706,g7417,g7144,g8146,g9011,g6418,
    g6994,g3658,g6926,g8268,g5064,g8362,g4958,I8064,g4376,g5070,g1913,g6021,
    g5594,g6421,g8728,g8730,g4225,g8385,g4073,g4796,g8070,g5089,g4473,g4912,
    g4124,g4377,g8331,g9023,g8888,g4287,I8237,g4483,g8087,g8305,g4199,g5438,
    g6041,g5189,g8748,g9327,g4797,g3893,g9146,g9135,g9346,g1834,I8573,g6168,
    g6058,g5561,g7193,g6911,g6743,g8283,g9240,g7682,g8920,g8459,g6411,g8718,
    g7598,g3222,g8261,g6474,g6203,g8637,g6992,g6610,g6694,g4314,I8400,g9147,
    g9136,g5062,g9347,g4228,g8721,g7606,g4408,g9013,g8907,g5298,g4399,g8940,
    I8588,g4230,g6400,g4433,g4427,g5031,g7607,g7325,g8826,g4395,g8741,g5005,
    g6423,g5765,g8609,g7828,g8308,g7615,g3229,g8066,I8034,g4342,g6999,g6633,
    g8711,g5069,g4097,g5343,g8455,g4154,g8827,g8333,g6732,g8846,g6753,g4155,
    g4783,g6043,g4312,g7628,g6434,g8290,g4129,g8256,g4830,g8816,g6914,g6013,
    g5589,g6413,g8700,g7323,g8263,g8950,g4068,I8079,g8723,g8257,g8817,g8301,
    g6060,g4699,g6178,g4398,g5008,g7278,g6995,g6435,g8441,g6699,I8432,g9084,
    g8964,g5830,g5065,g5122,g4319,g4352,g5033,g8458,g4186,g9276,g4386,g5518,
    g8074,g6053,g4083,g8080,g8713,g5142,g6157,g5081,g9120,g9052,I8078,g9277,
    g4387,g8688,g8857,g5783,g7724,g7337,g6121,g8326,g4145,g4391,g5001,g4107,
    g6436,g4159,g8383,g8924,g7611,g4507,g8634,g5483,g4315,g4047,g8361,g4474,
    g6707,g5140,g4166,g8327,g6039,g5068,g6439,g8303,g8696,g8732,g3286,g8944,
    g5699,g7600,g4128,g3081,g1682,g8316,g6970,g5035,g5119,g8697,g8914,g8795,
    g4902,g7175,g6893,g5599,g4745,g4490,g4823,g8820,g4366,g8936,g6771,g8317,
    g5125,g7184,g6138,g4355,g8922,g6738,g8060,g7535,g5106,g6991,g5689,g8460,
    g9038,g8966,g8739,g4055,g4118,g4167,g2783,g4367,g4872,g4549,g8937,g8079,
    g8294,g5046,g8840,g4193,g4393,g6915,g8942,g2912,g5107,g8704,g6002,g5539,
    g6402,g8954,g8763,g6762,g4740,g3258,g5047,g8912,g8796,g6464,g6177,g8929,
    g6728,g7447,g8626,g3984,g5017,g4219,g7182,g6902,g6394,g4962,g6580,g8735,
    g8075,g8949,g7632,g7445,g7653,g8292,g2952,g6438,g4829,g3314,g5090,g8646,
    g6409,g4180,g9270,g4380,g8439,g4420,g4794,g8702,g8919,g8952,g8788,g8276,
    g5063,g4100,g8404,g5118,g8764,g8231,g5057,g3939,g3925,g3915,g3907,I14941,
    g8699,I8225,I15250,I9107,g2214,g8707,g8082,I9047,g6270,I14484,I15055,
    I15051,I15052,I15053,I15054,I15111,g4824,g3315,g8656,I14985,I15019,I15018,
    g3083,g8850,g5040,g3900,g3895,g3890,g4363,g4790,g4786,I15102,I15098,I15099,
    I15100,I15101,g2229,I14771,I15231,I14959,I14960,g8009,I14302,I14951,I14952,
    I15085,g4810,I14759,I15243,I15239,I15240,I15241,I15242,I14758,g4736,I9044,
    g8658,I14990,g4737,g8176,g6452,g2206,g8862,I15169,g8360,g7421,g4318,I15084,
    I15110,g8812,I15254,g2230,I15230,I15265,I15261,I15262,I15263,I15264,I9099,
    I13553,g8819,I14767,g3541,g8811,I15297,I15298,I15041,g5558,I15275,g3602,
    g7062,I14766,I15165,g2014,I15253,I14754,I15175,I15021,I15017,I15020,I15073,
    I15274,g6209,I15292,g8805,g7784,I14219,I14366,I15109,I15283,g6710,I6209,
    g8706,I14980,g8232,I14942,I15040,I15252,I14969,g2213,g3012,g8128,g6910,
    I11603,g6193,g6197,g5556,I15072,I14496,I15152,g8863,I15400,I9029,I15113,
    I15112,g4734,I9038,I14480,I6208,I14468,g8523,g5021,g8694,I15229,I14479,
    I15228,g2995,g8818,I15232,g8680,g8855,I14772,g8847,I14970,g8861,I15031,
    g4735,I9041,g8679,g2262,I15043,I7232,I7233,g4727,g8236,I15284,I15285,
    I14834,I15086,I15082,I15083,g8279,g8613,g8806,g2367,g2352,g2378,g2330,
    I15042,g8859,g7083,I13220,I15030,g6259,g6185,I14933,I15075,I15071,I15074,
    I15276,g8807,g7191,I15272,I15273,g8803,I15251,g3129,g4237,I14932,g6119,
    g8091,g6184,g6174,g6214,g8655,g5546,I14831,I14753,g2368,I5757,I8363,g8230,
    I15290,I15291,I15033,I15029,I15032,g8233,I8224,g2315,g2385,g2294,g2395,
    g2043,I14495,g5555,I14467,I15147,g6153,I15172,g4835,I15044,g8659,I14485,
    I15888,g9192,I15887,I7466,I10092,g4881,I5521,I5519,g4528,I8606,I8607,g5625,
    I7538,I11143,I11142,I7467,g4839,I10906,I12575,I7181,I7179,I11178,I11179,
    I7421,I9548,I9549,I12597,I12598,g4548,I8636,I8637,I15855,I11110,I11108,
    I11177,I6524,I6522,I8510,I8245,I8243,g4313,I11186,I11184,I13685,g7237,
    I6258,I6257,I10889,I10890,I13800,I15819,I15817,I15818,I5600,I5598,I11185,
    I9978,g4880,I9243,g4305,I9241,I6274,I6273,g5284,I10745,I10743,I9746,I9747,
    I9234,g4310,I9233,I6170,I13587,g7234,I6939,g2051,I11117,I11115,g3232,I7531,
    g3938,I7610,I7611,I7505,I7503,I7011,g2333,I7009,I11123,I11122,I11751,
    I11750,g6701,I12032,I12033,I9195,I9196,I13639,g7257,I13638,I10329,I10327,
    I10981,I10982,I6904,g7069,I10328,I10314,I10315,I7480,I7478,I11841,g6158,
    I7569,I7567,I9964,I9963,I7010,g3681,I13786,I13787,I6757,I12051,I6940,I6941,
    I11116,I11615,I11614,I9057,I10991,g5632,I9547,I8255,I8253,g4492,I8537,
    I8538,I7423,I11165,I11163,I6234,I6232,I10744,g5550,I9979,I9980,I10849,
    I10847,I9242,g4476,I8511,I8512,I10790,I10791,I10848,g4871,I7240,I7239,
    g5567,I10361,I10359,I7443,I13600,g7244,I13598,I9691,I10992,I10993,g4231,
    I11137,I11135,I7533,I11873,g6187,I12552,I12550,I9985,g4836,I12870,I12871,
    g9191,I15856,I15857,I6843,I6842,I8119,I8152,I8150,I7460,I7459,I14473,
    I14472,I10789,g5512,I7937,I11136,I7479,I6813,I5599,I10000,I10001,I6740,
    I6739,g4513,I8582,I8583,I11164,I8939,I8938,I13214,I13215,I7156,I8940,
    I11575,I11574,I6997,I6998,I8635,g4831,I11109,I12551,I11102,I11103,I9151,
    g3883,I7453,I7452,I10874,I10875,I7568,I7157,g4869,I8536,I9278,I9276,I7149,
    I7150,I6275,I9235,I10980,I9693,I13640,I10899,I5506,I5507,I11757,g5056,
    g5039,g5023,g6695,I12016,I12017,I7187,I7188,I5520,I10835,I10836,I13397,
    I13395,I6905,I8328,I8326,I6523,I9965,I6750,I13213,g7065,g7082,I10224,
    I10225,I9070,I9071,I10061,g4910,I10060,I7616,g3889,I7437,I7438,I10360,
    I8166,g3231,I8164,I7215,I7216,g4575,I8679,I8680,I15863,I15862,I13396,
    I14246,I14244,I7277,I10071,g4954,I6172,I7617,I12576,I12577,I9153,I13377,
    I13378,I6134,I6133,I12080,I12078,I7892,I7891,I8393,I8392,g1910,I13785,
    I12031,I9476,I9477,I6171,I7140,I7138,I8121,I6202,I6201,I7086,I7087,I12869,
    I6776,I6774,I8605,I7214,I9475,I13003,I13002,I6996,I9692,I6878,I6876,I7180,
    I8659,I8658,I8133,I8134,I12079,I11752,I12596,g5590,I10888,I6103,I6104,
    g4502,I8559,I8560,I10039,I10040,I11149,I8558,I11842,I11843,I7148,I9947,
    I9948,I7436,I12015,I10900,I10901,I9058,I9059,I9946,g4905,I10625,I6135,
    g6559,I6758,I6759,g9202,I15881,I15882,I9182,I9181,I9382,I9381,I10197,
    I10196,I6500,I6499,I10855,I10854,I8151,I13376,I11096,I11094,I10867,I10866,
    I5505,I13802,I10313,g5305,I10819,I10818,I10306,I10307,I11549,g9179,I7085,
    I7485,I6102,I8132,I13686,I13687,I10094,I6203,g4700,I10019,I10017,I10018,
    I11150,I11151,I7270,I7268,I9999,I7609,I9171,g4244,I9169,I10923,I7069,I7068,
    I10300,I10298,I7540,I13004,I10198,I9745,I12853,I12854,I7173,I7174,g9190,
    I15880,I11080,I11078,I6916,I5696,I5695,I7510,I12852,I8503,I8504,I10305,
    I10062,I8678,I7070,I6752,I6917,I5620,I5621,I7241,I5697,I12053,I6233,I10335,
    I10334,I15898,I15899,I14839,I14837,I15897,g9203,I14838,I9069,I10820,g6680,
    g8073,g8092,I11171,I11170,g4893,I10038,I6775,I11079,g5697,I10143,I10142,
    I13599,I10010,I10011,I15850,I15848,I8339,I8338,I9768,I9769,I10093,I11158,
    I11156,I10321,I10322,I11144,I9767,g6722,I10223,I11172,I6539,I6538,I10320,
    I13017,I13016,I11550,I11551,I10953,g5565,I10952,I9170,I7468,I11095,I9826,
    I8660,I10908,I7576,I7574,g4294,I8244,I12052,I9827,I11124,I9152,I13801,
    I8340,I9194,I10834,g5568,I7893,I7186,I11875,I9277,I7444,I7445,I9994,I9992,
    I6751,I7939,I10336,I13018,I7461,I8956,I8955,I6741,I12180,I12181,I13589,
    I13588,g3924,I6066,I6064,I12833,I12834,I11616,I10873,I8957,I7158,I11101,
    I11874,I12832,I10073,I14474,I9828,I8502,g3914,I7532,I12951,I8470,I7512,
    I15889,I9183,I9383,I14245,I7279,I7938,I10144,I8581,I5619,g8644,g4563,
    I10868,I11157,I11576,I10954,I6924,I6923,g6709,I10072,g3894,I10924,I10925,
    I7172,I8165,I9954,I9953,I15864,I10856,I11758,I11759,g5310,g4298,I8254,
    I7575,I9986,I9987,I8120,I6259,g4252,g3906,I7504,I10907,g4911,I7278,I7618,
    I6540,I9993,I7511,I6501,I7139,I7539,I8394,I12952,I12953,g3899,g6163,I12179,
    g4821,I10009,I10627,I8327,I10626,I8472,I15849,I6925,I9955,I10299,I6906,
    g5291,I10080,I10078,I7269,I6877,I7486,I7487,I6844,I7422,g3886,I6814,I10079,
    I6918,g5312,g4359,I7429,I7430,I7454,g4894,g4888,g4884,I7428,g4456,I8471,
    I6065,I6815,g3885,g3310,g8635;

  dff DFF_0(CK,g397,g4635);
  dff DFF_1(CK,g1271,g5176);
  dff DFF_2(CK,g312,g4618);
  dff DFF_3(CK,g273,g4611);
  dff DFF_4(CK,g452,g449);
  dff DFF_5(CK,g948,g8664);
  dff DFF_6(CK,g629,g6827);
  dff DFF_7(CK,g207,g5733);
  dff DFF_8(CK,g1541,g7778);
  dff DFF_9(CK,g1153,g6856);
  dff DFF_10(CK,g940,g5735);
  dff DFF_11(CK,g976,g8864);
  dff DFF_12(CK,g498,g9111);
  dff DFF_13(CK,g314,g4620);
  dff DFF_14(CK,g1092,g7520);
  dff DFF_15(CK,g454,g4639);
  dff DFF_16(CK,g196,g5731);
  dff DFF_17(CK,g535,g3844);
  dff DFF_18(CK,g292,g4613);
  dff DFF_19(CK,g772,g6846);
  dff DFF_20(CK,g1375,g6869);
  dff DFF_21(CK,g689,g6371);
  dff DFF_22(CK,g183,g6309);
  dff DFF_23(CK,g359,g6336);
  dff DFF_24(CK,g1384,g6881);
  dff DFF_25(CK,g1339,g6865);
  dff DFF_26(CK,g20,g6386);
  dff DFF_27(CK,g1424,g3862);
  dff DFF_28(CK,g767,g6841);
  dff DFF_29(CK,g393,g4631);
  dff DFF_30(CK,g1077,g7767);
  dff DFF_31(CK,g1231,g1236);
  dff DFF_32(CK,g294,g4615);
  dff DFF_33(CK,g1477,g9036);
  dff DFF_34(CK,g4,g9372);
  dff DFF_35(CK,g608,g6806);
  dff DFF_36(CK,g1205,g1204);
  dff DFF_37(CK,g465,g6352);
  dff DFF_38(CK,g774,g6848);
  dff DFF_39(CK,g921,g916);
  dff DFF_40(CK,g1304,g1312);
  dff DFF_41(CK,g243,g6318);
  dff DFF_42(CK,g1499,g7772);
  dff DFF_43(CK,g80,g6778);
  dff DFF_44(CK,g1444,g5185);
  dff DFF_45(CK,g1269,g5740);
  dff DFF_46(CK,g600,g6807);
  dff DFF_47(CK,g423,g9105);
  dff DFF_48(CK,g771,g6845);
  dff DFF_49(CK,g803,g7757);
  dff DFF_50(CK,g843,g2647);
  dff DFF_51(CK,g315,g4621);
  dff DFF_52(CK,g455,g4640);
  dff DFF_53(CK,g906,g901);
  dff DFF_54(CK,g622,g6821);
  dff DFF_55(CK,g891,g3855);
  dff DFF_56(CK,g1014,g1012);
  dff DFF_57(CK,g984,g9133);
  dff DFF_58(CK,g117,g5153);
  dff DFF_59(CK,g137,g5150);
  dff DFF_60(CK,g527,g9110);
  dff DFF_61(CK,g1513,g1524);
  dff DFF_62(CK,g278,g6323);
  dff DFF_63(CK,g1378,g6880);
  dff DFF_64(CK,g718,g7753);
  dff DFF_65(CK,g598,g6797);
  dff DFF_66(CK,g1182,g1160);
  dff DFF_67(CK,g1288,g7527);
  dff DFF_68(CK,g1382,g6888);
  dff DFF_69(CK,g179,g5159);
  dff DFF_70(CK,g624,g6831);
  dff DFF_71(CK,g48,g9362);
  dff DFF_72(CK,g362,g9093);
  dff DFF_73(CK,g878,g890);
  dff DFF_74(CK,g270,g9092);
  dff DFF_75(CK,g763,g6836);
  dff DFF_76(CK,g710,g7751);
  dff DFF_77(CK,g730,g7754);
  dff DFF_78(CK,g295,g4616);
  dff DFF_79(CK,g1037,g7519);
  dff DFF_80(CK,g1102,g6855);
  dff DFF_81(CK,g483,g6356);
  dff DFF_82(CK,g775,g7759);
  dff DFF_83(CK,g621,g6819);
  dff DFF_84(CK,g1364,g6878);
  dff DFF_85(CK,g1454,g5187);
  dff DFF_86(CK,g1296,g7304);
  dff DFF_87(CK,g5,g9373);
  dff DFF_88(CK,g1532,g7781);
  dff DFF_89(CK,g587,g3852);
  dff DFF_90(CK,g741,g9386);
  dff DFF_91(CK,g13,g7308);
  dff DFF_92(CK,g606,g6804);
  dff DFF_93(CK,g1012,g6851);
  dff DFF_94(CK,g52,g6781);
  dff DFF_95(CK,g646,g4652);
  dff DFF_96(CK,g1412,g5745);
  dff DFF_97(CK,g327,g6332);
  dff DFF_98(CK,g1189,g6392);
  dff DFF_99(CK,g1389,g4658);
  dff DFF_100(CK,g1029,g2654);
  dff DFF_101(CK,g1371,g6868);
  dff DFF_102(CK,g1429,g2671);
  dff DFF_103(CK,g398,g4636);
  dff DFF_104(CK,g985,g7515);
  dff DFF_105(CK,g354,g4624);
  dff DFF_106(CK,g619,g6817);
  dff DFF_107(CK,g113,g5148);
  dff DFF_108(CK,g133,g5149);
  dff DFF_109(CK,g180,g5158);
  dff DFF_110(CK,g1138,g7524);
  dff DFF_111(CK,g1309,g1308);
  dff DFF_112(CK,g889,g7101);
  dff DFF_113(CK,g390,g6341);
  dff DFF_114(CK,g625,g6823);
  dff DFF_115(CK,g417,g9103);
  dff DFF_116(CK,g681,g7748);
  dff DFF_117(CK,g437,g6348);
  dff DFF_118(CK,g351,g9100);
  dff DFF_119(CK,g1201,g1200);
  dff DFF_120(CK,g109,g6785);
  dff DFF_121(CK,g1049,g8673);
  dff DFF_122(CK,g1098,g6854);
  dff DFF_123(CK,g200,g199);
  dff DFF_124(CK,g240,g6317);
  dff DFF_125(CK,g479,g4649);
  dff DFF_126(CK,g126,g6789);
  dff DFF_127(CK,g596,g6795);
  dff DFF_128(CK,g1268,g5175);
  dff DFF_129(CK,g222,g6313);
  dff DFF_130(CK,g420,g9104);
  dff DFF_131(CK,g3,g9360);
  dff DFF_132(CK,g58,g7734);
  dff DFF_133(CK,g172,g1270);
  dff DFF_134(CK,g387,g6340);
  dff DFF_135(CK,g840,g2648);
  dff DFF_136(CK,g365,g9094);
  dff DFF_137(CK,g1486,g8226);
  dff DFF_138(CK,g1504,g7773);
  dff DFF_139(CK,g1185,g1155);
  dff DFF_140(CK,g1385,g6883);
  dff DFF_141(CK,g583,g3851);
  dff DFF_142(CK,g822,g7512);
  dff DFF_143(CK,g1025,g8871);
  dff DFF_144(CK,g969,g966);
  dff DFF_145(CK,g768,g6842);
  dff DFF_146(CK,g174,g7737);
  dff DFF_147(CK,g685,g7749);
  dff DFF_148(CK,g1087,g6853);
  dff DFF_149(CK,g355,g4625);
  dff DFF_150(CK,g911,g906);
  dff DFF_151(CK,g1226,g6859);
  dff DFF_152(CK,g99,g6783);
  dff DFF_153(CK,g1045,g8224);
  dff DFF_154(CK,g1173,g7526);
  dff DFF_155(CK,g1373,g6871);
  dff DFF_156(CK,g186,g3830);
  dff DFF_157(CK,g760,g6833);
  dff DFF_158(CK,g959,g5169);
  dff DFF_159(CK,g1369,g6875);
  dff DFF_160(CK,g1007,g8867);
  dff DFF_161(CK,g1459,g3863);
  dff DFF_162(CK,g758,g6840);
  dff DFF_163(CK,g480,g6355);
  dff DFF_164(CK,g396,g4634);
  dff DFF_165(CK,g612,g6811);
  dff DFF_166(CK,g38,g5746);
  dff DFF_167(CK,g632,g6830);
  dff DFF_168(CK,g1415,g5180);
  dff DFF_169(CK,g1227,g7108);
  dff DFF_170(CK,g246,g6319);
  dff DFF_171(CK,g449,g3840);
  dff DFF_172(CK,g517,g4651);
  dff DFF_173(CK,g118,g6787);
  dff DFF_174(CK,g138,g6792);
  dff DFF_175(CK,g16,g1404);
  dff DFF_176(CK,g284,g9086);
  dff DFF_177(CK,g142,g6793);
  dff DFF_178(CK,g219,g6312);
  dff DFF_179(CK,g426,g9106);
  dff DFF_180(CK,g1388,g6882);
  dff DFF_181(CK,g806,g7510);
  dff DFF_182(CK,g846,g2646);
  dff DFF_183(CK,g1428,g2672);
  dff DFF_184(CK,g579,g3850);
  dff DFF_185(CK,g1030,g7518);
  dff DFF_186(CK,g614,g6812);
  dff DFF_187(CK,g1430,g4666);
  dff DFF_188(CK,g1247,g6380);
  dff DFF_189(CK,g669,g7745);
  dff DFF_190(CK,g110,g109);
  dff DFF_191(CK,g130,g6790);
  dff DFF_192(CK,g225,g6314);
  dff DFF_193(CK,g281,g9085);
  dff DFF_194(CK,g819,g7761);
  dff DFF_195(CK,g1308,g6385);
  dff DFF_196(CK,g611,g6810);
  dff DFF_197(CK,g631,g6829);
  dff DFF_198(CK,g1217,g6377);
  dff DFF_199(CK,g104,g6784);
  dff DFF_200(CK,g1365,g6867);
  dff DFF_201(CK,g825,g7513);
  dff DFF_202(CK,g1333,g6863);
  dff DFF_203(CK,g474,g4644);
  dff DFF_204(CK,g1396,g4662);
  dff DFF_205(CK,g141,g5151);
  dff DFF_206(CK,g1509,g7774);
  dff DFF_207(CK,g766,g6839);
  dff DFF_208(CK,g1018,g8869);
  dff DFF_209(CK,g588,g9031);
  dff DFF_210(CK,g1467,g8875);
  dff DFF_211(CK,g317,g4623);
  dff DFF_212(CK,g457,g4642);
  dff DFF_213(CK,g486,g6357);
  dff DFF_214(CK,g471,g6354);
  dff DFF_215(CK,g1381,g6887);
  dff DFF_216(CK,g1197,g1196);
  dff DFF_217(CK,g513,g9116);
  dff DFF_218(CK,g1397,g6389);
  dff DFF_219(CK,g533,g530);
  dff DFF_220(CK,g1021,g8870);
  dff DFF_221(CK,g1421,g5179);
  dff DFF_222(CK,g952,g8668);
  dff DFF_223(CK,g1263,g5737);
  dff DFF_224(CK,g580,g6368);
  dff DFF_225(CK,g615,g6813);
  dff DFF_226(CK,g1257,g5738);
  dff DFF_227(CK,g46,g8955);
  dff DFF_228(CK,g402,g6343);
  dff DFF_229(CK,g998,g1005);
  dff DFF_230(CK,g1041,g7765);
  dff DFF_231(CK,g297,g6324);
  dff DFF_232(CK,g954,g8670);
  dff DFF_233(CK,g105,g104);
  dff DFF_234(CK,g145,g5152);
  dff DFF_235(CK,g212,g4601);
  dff DFF_236(CK,g1368,g6874);
  dff DFF_237(CK,g232,g4606);
  dff DFF_238(CK,g990,g7516);
  dff DFF_239(CK,g475,g4645);
  dff DFF_240(CK,g33,g5184);
  dff DFF_241(CK,g951,g8667);
  dff DFF_242(CK,g799,g7756);
  dff DFF_243(CK,g812,g7758);
  dff DFF_244(CK,g567,g6367);
  dff DFF_245(CK,g313,g4619);
  dff DFF_246(CK,g333,g6334);
  dff DFF_247(CK,g168,g7742);
  dff DFF_248(CK,g214,g4603);
  dff DFF_249(CK,g234,g4608);
  dff DFF_250(CK,g652,g646);
  dff DFF_251(CK,g1126,g8674);
  dff DFF_252(CK,g1400,g6390);
  dff DFF_253(CK,g1326,g7306);
  dff DFF_254(CK,g92,g6794);
  dff DFF_255(CK,g309,g6328);
  dff DFF_256(CK,g211,g4600);
  dff DFF_257(CK,g834,g2650);
  dff DFF_258(CK,g231,g4605);
  dff DFF_259(CK,g557,g6366);
  dff DFF_260(CK,g1383,g6889);
  dff DFF_261(CK,g1220,g6378);
  dff DFF_262(CK,g158,g7740);
  dff DFF_263(CK,g627,g6825);
  dff DFF_264(CK,g661,g7743);
  dff DFF_265(CK,g77,g6777);
  dff DFF_266(CK,g831,g2651);
  dff DFF_267(CK,g1327,g7307);
  dff DFF_268(CK,g293,g4614);
  dff DFF_269(CK,g1146,g1612);
  dff DFF_270(CK,g89,g92);
  dff DFF_271(CK,g150,g7738);
  dff DFF_272(CK,g773,g6847);
  dff DFF_273(CK,g859,g8221);
  dff DFF_274(CK,g1240,g1235);
  dff DFF_275(CK,g518,g6361);
  dff DFF_276(CK,g1472,g8960);
  dff DFF_277(CK,g1443,g4667);
  dff DFF_278(CK,g436,g4638);
  dff DFF_279(CK,g405,g6344);
  dff DFF_280(CK,g1034,g8957);
  dff DFF_281(CK,g1147,g1146);
  dff DFF_282(CK,g374,g4627);
  dff DFF_283(CK,g98,g5146);
  dff DFF_284(CK,g563,g9029);
  dff DFF_285(CK,g510,g9115);
  dff DFF_286(CK,g530,g3842);
  dff DFF_287(CK,g215,g4604);
  dff DFF_288(CK,g235,g4609);
  dff DFF_289(CK,g1013,g1014);
  dff DFF_290(CK,g6,g9374);
  dff DFF_291(CK,g55,g7733);
  dff DFF_292(CK,g1317,g5743);
  dff DFF_293(CK,g504,g9113);
  dff DFF_294(CK,g665,g7744);
  dff DFF_295(CK,g544,g6365);
  dff DFF_296(CK,g371,g368);
  dff DFF_297(CK,g62,g7509);
  dff DFF_298(CK,g792,g5162);
  dff DFF_299(CK,g468,g6353);
  dff DFF_300(CK,g815,g7760);
  dff DFF_301(CK,g1460,g4668);
  dff DFF_302(CK,g553,g9028);
  dff DFF_303(CK,g623,g6822);
  dff DFF_304(CK,g501,g9112);
  dff DFF_305(CK,g1190,g8677);
  dff DFF_306(CK,g1390,g4659);
  dff DFF_307(CK,g74,g6776);
  dff DFF_308(CK,g1156,g1081);
  dff DFF_309(CK,g318,g6329);
  dff DFF_310(CK,g458,g4643);
  dff DFF_311(CK,g342,g9097);
  dff DFF_312(CK,g1250,g7111);
  dff DFF_313(CK,g1163,g2655);
  dff DFF_314(CK,g1363,g6877);
  dff DFF_315(CK,g1432,g5183);
  dff DFF_316(CK,g1053,g8873);
  dff DFF_317(CK,g252,g6321);
  dff DFF_318(CK,g330,g6333);
  dff DFF_319(CK,g264,g9090);
  dff DFF_320(CK,g1157,g1156);
  dff DFF_321(CK,g1357,g8675);
  dff DFF_322(CK,g375,g4628);
  dff DFF_323(CK,g68,g6774);
  dff DFF_324(CK,g852,g2644);
  dff DFF_325(CK,g261,g9089);
  dff DFF_326(CK,g516,g4650);
  dff DFF_327(CK,g536,g6363);
  dff DFF_328(CK,g979,g7104);
  dff DFF_329(CK,g778,g7296);
  dff DFF_330(CK,g199,g3832);
  dff DFF_331(CK,g1292,g7302);
  dff DFF_332(CK,g290,g287);
  dff DFF_333(CK,g1084,g7106);
  dff DFF_334(CK,g1439,g5182);
  dff DFF_335(CK,g770,g6844);
  dff DFF_336(CK,g1276,g6384);
  dff DFF_337(CK,g890,g7102);
  dff DFF_338(CK,g1004,g7105);
  dff DFF_339(CK,g1404,g1403);
  dff DFF_340(CK,g93,g5145);
  dff DFF_341(CK,g2,g9361);
  dff DFF_342(CK,g287,g3836);
  dff DFF_343(CK,g560,g6370);
  dff DFF_344(CK,g1224,g6857);
  dff DFF_345(CK,g1320,g7114);
  dff DFF_346(CK,g617,g6815);
  dff DFF_347(CK,g316,g4622);
  dff DFF_348(CK,g336,g9095);
  dff DFF_349(CK,g933,g5166);
  dff DFF_350(CK,g456,g4641);
  dff DFF_351(CK,g345,g9098);
  dff DFF_352(CK,g628,g6826);
  dff DFF_353(CK,g8,g9376);
  dff DFF_354(CK,g887,g7099);
  dff DFF_355(CK,g789,g7297);
  dff DFF_356(CK,g173,g7736);
  dff DFF_357(CK,g550,g9027);
  dff DFF_358(CK,g255,g9087);
  dff DFF_359(CK,g949,g8665);
  dff DFF_360(CK,g1244,g2659);
  dff DFF_361(CK,g620,g6818);
  dff DFF_362(CK,g1435,g5181);
  dff DFF_363(CK,g477,g4647);
  dff DFF_364(CK,g926,g878);
  dff DFF_365(CK,g368,g3838);
  dff DFF_366(CK,g855,g8220);
  dff DFF_367(CK,g1214,g5736);
  dff DFF_368(CK,g1110,g7299);
  dff DFF_369(CK,g1310,g1309);
  dff DFF_370(CK,g296,g4617);
  dff DFF_371(CK,g972,g2653);
  dff DFF_372(CK,g1402,g6391);
  dff DFF_373(CK,g1236,g1240);
  dff DFF_374(CK,g896,g891);
  dff DFF_375(CK,g613,g6820);
  dff DFF_376(CK,g566,g3848);
  dff DFF_377(CK,g1394,g6388);
  dff DFF_378(CK,g1489,g7770);
  dff DFF_379(CK,g883,g921);
  dff DFF_380(CK,g47,g9389);
  dff DFF_381(CK,g971,g5171);
  dff DFF_382(CK,g609,g6808);
  dff DFF_383(CK,g103,g5157);
  dff DFF_384(CK,g1254,g6381);
  dff DFF_385(CK,g556,g3847);
  dff DFF_386(CK,g1409,g5178);
  dff DFF_387(CK,g626,g6824);
  dff DFF_388(CK,g1229,g7110);
  dff DFF_389(CK,g782,g5734);
  dff DFF_390(CK,g237,g6316);
  dff DFF_391(CK,g942,g2652);
  dff DFF_392(CK,g228,g6315);
  dff DFF_393(CK,g706,g7750);
  dff DFF_394(CK,g746,g8956);
  dff DFF_395(CK,g1462,g8678);
  dff DFF_396(CK,g963,g7764);
  dff DFF_397(CK,g129,g5156);
  dff DFF_398(CK,g837,g2649);
  dff DFF_399(CK,g599,g6798);
  dff DFF_400(CK,g1192,g1191);
  dff DFF_401(CK,g828,g7762);
  dff DFF_402(CK,g1392,g6387);
  dff DFF_403(CK,g492,g6359);
  dff DFF_404(CK,g95,g94);
  dff DFF_405(CK,g944,g6372);
  dff DFF_406(CK,g195,g3831);
  dff DFF_407(CK,g1431,g2673);
  dff DFF_408(CK,g1252,g2661);
  dff DFF_409(CK,g356,g6335);
  dff DFF_410(CK,g953,g8669);
  dff DFF_411(CK,g1176,g5172);
  dff DFF_412(CK,g1376,g6890);
  dff DFF_413(CK,g1005,g1004);
  dff DFF_414(CK,g1405,g5744);
  dff DFF_415(CK,g901,g896);
  dff DFF_416(CK,g1270,g1271);
  dff DFF_417(CK,g1225,g6858);
  dff DFF_418(CK,g1073,g9145);
  dff DFF_419(CK,g1324,g7118);
  dff DFF_420(CK,g1069,g9134);
  dff DFF_421(CK,g443,g9101);
  dff DFF_422(CK,g1377,g6891);
  dff DFF_423(CK,g377,g4630);
  dff DFF_424(CK,g618,g6816);
  dff DFF_425(CK,g602,g6800);
  dff DFF_426(CK,g213,g4602);
  dff DFF_427(CK,g233,g4607);
  dff DFF_428(CK,g1199,g6375);
  dff DFF_429(CK,g1399,g3861);
  dff DFF_430(CK,g83,g6779);
  dff DFF_431(CK,g888,g7100);
  dff DFF_432(CK,g573,g9033);
  dff DFF_433(CK,g399,g6342);
  dff DFF_434(CK,g1245,g1244);
  dff DFF_435(CK,g507,g9114);
  dff DFF_436(CK,g547,g9026);
  dff DFF_437(CK,g108,g5147);
  dff DFF_438(CK,g610,g6809);
  dff DFF_439(CK,g630,g6828);
  dff DFF_440(CK,g1207,g5173);
  dff DFF_441(CK,g249,g6320);
  dff DFF_442(CK,g65,g4598);
  dff DFF_443(CK,g916,g911);
  dff DFF_444(CK,g936,g5168);
  dff DFF_445(CK,g478,g4648);
  dff DFF_446(CK,g604,g6802);
  dff DFF_447(CK,g945,g5170);
  dff DFF_448(CK,g1114,g7521);
  dff DFF_449(CK,g100,g99);
  dff DFF_450(CK,g429,g9107);
  dff DFF_451(CK,g809,g7511);
  dff DFF_452(CK,g849,g2645);
  dff DFF_453(CK,g1408,g5177);
  dff DFF_454(CK,g1336,g6864);
  dff DFF_455(CK,g601,g6799);
  dff DFF_456(CK,g122,g6788);
  dff DFF_457(CK,g1065,g9117);
  dff DFF_458(CK,g1122,g8225);
  dff DFF_459(CK,g1228,g7109);
  dff DFF_460(CK,g495,g6360);
  dff DFF_461(CK,g1322,g7116);
  dff DFF_462(CK,g1230,g7300);
  dff DFF_463(CK,g1033,g9034);
  dff DFF_464(CK,g267,g9091);
  dff DFF_465(CK,g1195,g6374);
  dff DFF_466(CK,g1395,g1393);
  dff DFF_467(CK,g373,g4626);
  dff DFF_468(CK,g274,g4612);
  dff DFF_469(CK,g1266,g5739);
  dff DFF_470(CK,g714,g7752);
  dff DFF_471(CK,g734,g7755);
  dff DFF_472(CK,g1142,g8874);
  dff DFF_473(CK,g1342,g7119);
  dff DFF_474(CK,g769,g6843);
  dff DFF_475(CK,g1081,g6852);
  dff DFF_476(CK,g1481,g7769);
  dff DFF_477(CK,g1097,g1185);
  dff DFF_478(CK,g543,g3846);
  dff DFF_479(CK,g1154,g1153);
  dff DFF_480(CK,g1354,g7768);
  dff DFF_481(CK,g489,g6358);
  dff DFF_482(CK,g874,g4654);
  dff DFF_483(CK,g121,g5154);
  dff DFF_484(CK,g591,g9032);
  dff DFF_485(CK,g616,g6814);
  dff DFF_486(CK,g1267,g4656);
  dff DFF_487(CK,g1312,g1311);
  dff DFF_488(CK,g605,g6803);
  dff DFF_489(CK,g182,g5161);
  dff DFF_490(CK,g1401,g1399);
  dff DFF_491(CK,g950,g8666);
  dff DFF_492(CK,g1329,g2663);
  dff DFF_493(CK,g408,g6345);
  dff DFF_494(CK,g871,g5167);
  dff DFF_495(CK,g759,g6832);
  dff DFF_496(CK,g146,g7735);
  dff DFF_497(CK,g202,g5732);
  dff DFF_498(CK,g440,g6349);
  dff DFF_499(CK,g476,g4646);
  dff DFF_500(CK,g184,g6310);
  dff DFF_501(CK,g1149,g7525);
  dff DFF_502(CK,g1398,g1396);
  dff DFF_503(CK,g210,g3834);
  dff DFF_504(CK,g394,g4632);
  dff DFF_505(CK,g86,g6780);
  dff DFF_506(CK,g570,g9030);
  dff DFF_507(CK,g275,g6322);
  dff DFF_508(CK,g303,g6326);
  dff DFF_509(CK,g125,g5155);
  dff DFF_510(CK,g181,g5160);
  dff DFF_511(CK,g1524,g6393);
  dff DFF_512(CK,g595,g576);
  dff DFF_513(CK,g1319,g7113);
  dff DFF_514(CK,g863,g8222);
  dff DFF_515(CK,g1211,g5174);
  dff DFF_516(CK,g966,g8223);
  dff DFF_517(CK,g1186,g1182);
  dff DFF_518(CK,g1386,g6884);
  dff DFF_519(CK,g875,g5165);
  dff DFF_520(CK,g1170,g1173);
  dff DFF_521(CK,g1370,g6876);
  dff DFF_522(CK,g201,g200);
  dff DFF_523(CK,g1325,g7305);
  dff DFF_524(CK,g1280,g7112);
  dff DFF_525(CK,g1106,g7107);
  dff DFF_526(CK,g1061,g9035);
  dff DFF_527(CK,g1387,g6885);
  dff DFF_528(CK,g762,g6835);
  dff DFF_529(CK,g1461,g4669);
  dff DFF_530(CK,g378,g6337);
  dff DFF_531(CK,g1200,g1199);
  dff DFF_532(CK,g1514,g7775);
  dff DFF_533(CK,g1403,g1402);
  dff DFF_534(CK,g1345,g7528);
  dff DFF_535(CK,g1191,g6373);
  dff DFF_536(CK,g1391,g1390);
  dff DFF_537(CK,g185,g4599);
  dff DFF_538(CK,g1307,g3858);
  dff DFF_539(CK,g1159,g1157);
  dff DFF_540(CK,g1223,g6379);
  dff DFF_541(CK,g446,g9102);
  dff DFF_542(CK,g1416,g4665);
  dff DFF_543(CK,g395,g4633);
  dff DFF_544(CK,g764,g6837);
  dff DFF_545(CK,g1251,g6860);
  dff DFF_546(CK,g216,g6311);
  dff DFF_547(CK,g236,g4610);
  dff DFF_548(CK,g205,g3835);
  dff DFF_549(CK,g540,g6364);
  dff DFF_550(CK,g576,g3849);
  dff DFF_551(CK,g1537,g7777);
  dff DFF_552(CK,g727,g8228);
  dff DFF_553(CK,g999,g8865);
  dff DFF_554(CK,g761,g6834);
  dff DFF_555(CK,g1272,g6383);
  dff DFF_556(CK,g1243,g2660);
  dff DFF_557(CK,g1328,g7309);
  dff DFF_558(CK,g1130,g7522);
  dff DFF_559(CK,g1330,g6862);
  dff DFF_560(CK,g114,g6786);
  dff DFF_561(CK,g134,g6791);
  dff DFF_562(CK,g1166,g1167);
  dff DFF_563(CK,g524,g9109);
  dff DFF_564(CK,g1366,g6866);
  dff DFF_565(CK,g348,g9099);
  dff DFF_566(CK,g1148,g1147);
  dff DFF_567(CK,g1348,g7529);
  dff DFF_568(CK,g1155,g1154);
  dff DFF_569(CK,g1260,g6382);
  dff DFF_570(CK,g7,g9375);
  dff DFF_571(CK,g258,g9088);
  dff DFF_572(CK,g521,g6362);
  dff DFF_573(CK,g300,g6325);
  dff DFF_574(CK,g765,g6838);
  dff DFF_575(CK,g1118,g7766);
  dff DFF_576(CK,g1167,g1170);
  dff DFF_577(CK,g1318,g6861);
  dff DFF_578(CK,g1367,g6873);
  dff DFF_579(CK,g677,g7747);
  dff DFF_580(CK,g376,g4629);
  dff DFF_581(CK,g1057,g8959);
  dff DFF_582(CK,g973,g8672);
  dff DFF_583(CK,g1193,g1192);
  dff DFF_584(CK,g1393,g2664);
  dff DFF_585(CK,g1549,g7780);
  dff DFF_586(CK,g1321,g7115);
  dff DFF_587(CK,g1253,g5741);
  dff DFF_588(CK,g1519,g8227);
  dff DFF_589(CK,g584,g6369);
  dff DFF_590(CK,g539,g3845);
  dff DFF_591(CK,g324,g6331);
  dff DFF_592(CK,g432,g9108);
  dff DFF_593(CK,g1158,g1159);
  dff DFF_594(CK,g321,g6330);
  dff DFF_595(CK,g1311,g1310);
  dff DFF_596(CK,g414,g6347);
  dff DFF_597(CK,g1374,g6872);
  dff DFF_598(CK,g94,g6782);
  dff DFF_599(CK,g1284,g7301);
  dff DFF_600(CK,g1545,g7779);
  dff DFF_601(CK,g1380,g6886);
  dff DFF_602(CK,g673,g7746);
  dff DFF_603(CK,g607,g6805);
  dff DFF_604(CK,g306,g6327);
  dff DFF_605(CK,g943,g8671);
  dff DFF_606(CK,g162,g7741);
  dff DFF_607(CK,g411,g6346);
  dff DFF_608(CK,g866,g5163);
  dff DFF_609(CK,g1204,g1203);
  dff DFF_610(CK,g1300,g7303);
  dff DFF_611(CK,g384,g6339);
  dff DFF_612(CK,g339,g9096);
  dff DFF_613(CK,g459,g6350);
  dff DFF_614(CK,g1323,g7117);
  dff DFF_615(CK,g381,g6338);
  dff DFF_616(CK,g1528,g7776);
  dff DFF_617(CK,g1351,g7530);
  dff DFF_618(CK,g597,g6796);
  dff DFF_619(CK,g1372,g6870);
  dff DFF_620(CK,g154,g7739);
  dff DFF_621(CK,g435,g4637);
  dff DFF_622(CK,g970,g963);
  dff DFF_623(CK,g1134,g7523);
  dff DFF_624(CK,g995,g7517);
  dff DFF_625(CK,g190,g201);
  dff DFF_626(CK,g1313,g5742);
  dff DFF_627(CK,g603,g6801);
  dff DFF_628(CK,g1494,g7771);
  dff DFF_629(CK,g462,g6351);
  dff DFF_630(CK,g1160,g1163);
  dff DFF_631(CK,g1360,g8676);
  dff DFF_632(CK,g1450,g5186);
  dff DFF_633(CK,g187,g5730);
  dff DFF_634(CK,g1179,g1186);
  dff DFF_635(CK,g1379,g6879);
  dff DFF_636(CK,g12,g8662);
  dff DFF_637(CK,g71,g6775);
  not NOT_0(g1658,g1313);
  not NOT_1(g1777,g611);
  not NOT_2(I9325,g4242);
  not NOT_3(I7758,g2605);
  not NOT_4(g5652,I10135);
  not NOT_5(I13502,g7135);
  not NOT_6(g6895,I12558);
  not NOT_7(g3880,g2965);
  not NOT_8(g6837,I12382);
  not NOT_9(I15824,g9157);
  not NOT_10(g5843,g5367);
  not NOT_11(I6112,g4);
  not NOT_12(g7189,I13109);
  not NOT_13(g8970,I15414);
  not NOT_14(I6267,g100);
  not NOT_15(g6062,I10675);
  not NOT_16(I16126,g9354);
  not NOT_17(I10519,g5242);
  not NOT_18(I15181,g8734);
  not NOT_19(I11443,g6038);
  not NOT_20(I12436,g6635);
  not NOT_21(I10675,g5662);
  not NOT_22(g2547,I6371);
  not NOT_23(I7365,g3061);
  not NOT_24(I10154,g5109);
  not NOT_25(g1611,g1073);
  not NOT_26(I11278,g5780);
  not NOT_27(g7171,g7071);
  not NOT_28(I14154,g7558);
  not NOT_29(I12274,g6672);
  not NOT_30(g8224,I14451);
  not NOT_31(g5834,I10525);
  not NOT_32(g5971,I10587);
  not NOT_33(g3978,g3160);
  not NOT_34(I6676,g1603);
  not NOT_35(g3612,I7082);
  not NOT_36(I8520,g3652);
  not NOT_37(g2892,g2266);
  not NOT_38(I13469,g7123);
  not NOT_39(I12346,g6737);
  not NOT_40(I9636,g4802);
  not NOT_41(I14637,g8012);
  not NOT_42(g6788,I12235);
  not NOT_43(g1799,I5657);
  not NOT_44(g3935,I7602);
  not NOT_45(I5933,g1158);
  not NOT_46(g9207,g9197);
  not NOT_47(I13039,g6961);
  not NOT_48(I15426,g8895);
  not NOT_49(g5598,g4938);
  not NOT_50(g1674,g1514);
  not NOT_51(g7281,I13277);
  not NOT_52(g3982,g3192);
  not NOT_53(g4666,I8913);
  not NOT_54(I15190,g8685);
  not NOT_55(g2945,g2364);
  not NOT_56(g5121,I9515);
  not NOT_57(g3128,I6839);
  not NOT_58(g3629,g2424);
  not NOT_59(g7297,I13323);
  not NOT_60(g5670,I10157);
  not NOT_61(I11815,g6169);
  not NOT_62(g6842,I12397);
  not NOT_63(g3130,I6849);
  not NOT_64(g9088,I15654);
  not NOT_65(g8789,g8564);
  not NOT_66(g3542,g1777);
  not NOT_67(I12292,g6657);
  not NOT_68(g6298,I11221);
  not NOT_69(g2709,g1747);
  not NOT_70(I11677,g6076);
  not NOT_71(g6392,I11503);
  not NOT_72(g4648,I8859);
  not NOT_73(I8829,g4029);
  not NOT_74(I15546,g9007);
  not NOT_75(g1680,I5515);
  not NOT_76(I15211,g8808);
  not NOT_77(g2340,g1327);
  not NOT_78(I12409,g6398);
  not NOT_79(g4655,I8880);
  not NOT_80(g7745,I14106);
  not NOT_81(g7138,I12996);
  not NOT_82(I6703,g1983);
  not NOT_83(g5938,g5412);
  not NOT_84(g8771,g8564);
  not NOT_85(g2478,g31);
  not NOT_86(g5813,I10472);
  not NOT_87(g7338,I13432);
  not NOT_88(g2907,g2289);
  not NOT_89(g1744,g600);
  not NOT_90(g9215,I15921);
  not NOT_91(g7109,I12915);
  not NOT_92(g6854,I12433);
  not NOT_93(I12635,g6509);
  not NOT_94(g7309,I13359);
  not NOT_95(g1802,g628);
  not NOT_96(I10439,g5214);
  not NOT_97(g2959,g1926);
  not NOT_98(I14728,g8152);
  not NOT_99(I8733,g3996);
  not NOT_100(I14439,g8063);
  not NOT_101(g2517,I6348);
  not NOT_102(g4010,g3097);
  not NOT_103(I7662,g3642);
  not NOT_104(I9446,g3926);
  not NOT_105(I8974,g3871);
  not NOT_106(g5740,I10277);
  not NOT_107(g5519,I9929);
  not NOT_108(g9114,I15732);
  not NOT_109(g1558,I5435);
  not NOT_110(I7290,g2936);
  not NOT_111(g2876,g2231);
  not NOT_112(g9314,I16058);
  not NOT_113(I11884,g6091);
  not NOT_114(I9145,g4264);
  not NOT_115(I6468,g1917);
  not NOT_116(g5606,g4748);
  not NOT_117(I8796,g3934);
  not NOT_118(g7759,I14148);
  not NOT_119(I14349,g7588);
  not NOT_120(I11410,g5845);
  not NOT_121(I12164,g5847);
  not NOT_122(g695,I5392);
  not NOT_123(g6708,g6250);
  not NOT_124(I13410,g7274);
  not NOT_125(I15625,g9000);
  not NOT_126(g6520,I11704);
  not NOT_127(g1901,I5781);
  not NOT_128(g6219,I10998);
  not NOT_129(g6640,I11908);
  not NOT_130(I8980,g4535);
  not NOT_131(g3902,I7495);
  not NOT_132(I12891,g6950);
  not NOT_133(I11479,g6201);
  not NOT_134(I11666,g5772);
  not NOT_135(g5687,I10190);
  not NOT_136(g2915,I6643);
  not NOT_137(I13666,g7238);
  not NOT_138(g6252,g5418);
  not NOT_139(g6812,I12307);
  not NOT_140(g4372,I8357);
  not NOT_141(g7049,I12813);
  not NOT_142(g3512,g1616);
  not NOT_143(I13478,g7126);
  not NOT_144(g5586,g4938);
  not NOT_145(g6958,I12675);
  not NOT_146(I15943,g9214);
  not NOT_147(g4618,I8769);
  not NOT_148(I6716,g1721);
  not NOT_149(g6376,I11455);
  not NOT_150(g4667,I8916);
  not NOT_151(I5981,g459);
  not NOT_152(I8177,g2810);
  not NOT_153(I7847,g3798);
  not NOT_154(I16055,g9291);
  not NOT_155(g9336,I16084);
  not NOT_156(g2310,I6087);
  not NOT_157(g7715,I14022);
  not NOT_158(g1600,g976);
  not NOT_159(g1574,g681);
  not NOT_160(g1864,g162);
  not NOT_161(g4566,g2902);
  not NOT_162(I11556,g6065);
  not NOT_163(g7098,g6525);
  not NOT_164(I5997,g114);
  not NOT_165(g6829,I12358);
  not NOT_166(g7498,I13672);
  not NOT_167(g2663,I6460);
  not NOT_168(I12108,g5939);
  not NOT_169(g6765,I12164);
  not NOT_170(g3529,g2323);
  not NOT_171(g8959,I15391);
  not NOT_172(I6198,g483);
  not NOT_173(g4693,I8974);
  not NOT_174(I13580,g7208);
  not NOT_175(g4134,g3676);
  not NOT_176(g3649,g2424);
  not NOT_177(I14139,g7548);
  not NOT_178(I9416,g4273);
  not NOT_179(I12283,g6692);
  not NOT_180(g8482,g8094);
  not NOT_181(g5525,g4934);
  not NOT_182(g3851,I7356);
  not NOT_183(g5645,g4748);
  not NOT_184(I5353,g3833);
  not NOT_185(g2402,g29);
  not NOT_186(I7950,g2774);
  not NOT_187(g2824,g1688);
  not NOT_188(g1580,g706);
  not NOT_189(g2236,I5969);
  not NOT_190(g7584,I13897);
  not NOT_191(g4555,g2894);
  not NOT_192(g9065,I15589);
  not NOT_193(I9642,g4788);
  not NOT_194(g7539,I13797);
  not NOT_195(I15411,g8897);
  not NOT_196(I15527,g9020);
  not NOT_197(I10415,g5397);
  not NOT_198(I13084,g7071);
  not NOT_199(g9322,g9313);
  not NOT_200(g3964,g3160);
  not NOT_201(g4792,I9111);
  not NOT_202(g9230,I15950);
  not NOT_203(g6225,I11014);
  not NOT_204(I8781,g3932);
  not NOT_205(I8898,g4089);
  not NOT_206(g6073,g5384);
  not NOT_207(g2877,g2232);
  not NOT_208(g6796,I12259);
  not NOT_209(g1736,I5577);
  not NOT_210(I12091,g5988);
  not NOT_211(g4621,I8778);
  not NOT_212(g5607,g4938);
  not NOT_213(g9033,I15513);
  not NOT_214(g7162,I13060);
  not NOT_215(g7268,I13244);
  not NOT_216(g7019,I12771);
  not NOT_217(I11740,g6136);
  not NOT_218(g7362,I13502);
  not NOT_219(g5158,I9600);
  not NOT_220(I13740,g7364);
  not NOT_221(I9654,g4792);
  not NOT_222(I15894,g9195);
  not NOT_223(g6324,I11299);
  not NOT_224(I7723,g3052);
  not NOT_225(g4113,I7950);
  not NOT_226(g6069,I10690);
  not NOT_227(g2556,g1190);
  not NOT_228(g1889,g1018);
  not NOT_229(I7101,g2478);
  not NOT_230(I5901,g52);
  not NOT_231(g2222,I5939);
  not NOT_232(I13676,g7256);
  not NOT_233(g9096,I15678);
  not NOT_234(I8291,g878);
  not NOT_235(I13373,g7270);
  not NOT_236(g2928,g2326);
  not NOT_237(g4202,g2810);
  not NOT_238(g8663,I14783);
  not NOT_239(I7605,g2752);
  not NOT_240(I15714,g9077);
  not NOT_241(g5587,g4938);
  not NOT_242(g2930,g2328);
  not NOT_243(I15315,g8738);
  not NOT_244(I11800,g6164);
  not NOT_245(g1871,I5754);
  not NOT_246(g4908,g4088);
  not NOT_247(g6377,I11458);
  not NOT_248(g6206,g5639);
  not NOT_249(g5311,g4938);
  not NOT_250(g2899,g2272);
  not NOT_251(g9195,I15871);
  not NOT_252(g4094,I7905);
  not NOT_253(I11936,g5918);
  not NOT_254(g3872,g2954);
  not NOT_255(I15202,g8797);
  not NOT_256(g3652,I7132);
  not NOT_257(g4567,g2903);
  not NOT_258(g7728,I14055);
  not NOT_259(g7486,I13646);
  not NOT_260(g3843,I7332);
  not NOT_261(g3989,g3131);
  not NOT_262(I6186,g138);
  not NOT_263(g7730,I14061);
  not NOT_264(I9612,g4776);
  not NOT_265(I10608,g5701);
  not NOT_266(g5174,I9648);
  not NOT_267(g8762,g8585);
  not NOT_268(g7504,I13692);
  not NOT_269(I15978,g9235);
  not NOT_270(I14115,g7563);
  not NOT_271(g7185,I13099);
  not NOT_272(g4776,I9081);
  not NOT_273(I7041,g2401);
  not NOT_274(g6849,I12418);
  not NOT_275(I9935,g4812);
  not NOT_276(g4593,g2939);
  not NOT_277(I11964,g5971);
  not NOT_278(g3549,g2404);
  not NOT_279(g3834,I7305);
  not NOT_280(g3971,I7688);
  not NOT_281(g7070,g6562);
  not NOT_282(g2295,g995);
  not NOT_283(I14052,g7494);
  not NOT_284(g2237,I5972);
  not NOT_285(g7470,g7253);
  not NOT_286(I15741,g9083);
  not NOT_287(g8657,I14763);
  not NOT_288(g6781,I12214);
  not NOT_289(g7425,I13550);
  not NOT_290(g5180,I9666);
  not NOT_291(g2844,I6574);
  not NOT_292(I8215,g3577);
  not NOT_293(g6898,I12567);
  not NOT_294(g1838,g1450);
  not NOT_295(g5591,g4841);
  not NOT_296(g6900,I12571);
  not NOT_297(g8222,I14445);
  not NOT_298(I8886,g4308);
  not NOT_299(g5832,I10519);
  not NOT_300(I14813,g8640);
  not NOT_301(g1795,I5649);
  not NOT_302(g6797,I12262);
  not NOT_303(g1737,g597);
  not NOT_304(g2394,I6270);
  not NOT_305(g9248,I15978);
  not NOT_306(g1809,g759);
  not NOT_307(I10973,g5726);
  not NOT_308(I14798,g8605);
  not NOT_309(g6245,g5690);
  not NOT_310(g4360,I8333);
  not NOT_311(I7368,g3018);
  not NOT_312(g9255,I15985);
  not NOT_313(g9081,I15635);
  not NOT_314(I12948,g6919);
  not NOT_315(I13909,g7339);
  not NOT_316(I15735,g9078);
  not NOT_317(g4521,g2866);
  not NOT_318(I14184,g7726);
  not NOT_319(g1672,g1499);
  not NOT_320(I14674,g7788);
  not NOT_321(g8464,g8039);
  not NOT_322(g6291,I11200);
  not NOT_323(I12702,g6497);
  not NOT_324(g2557,g940);
  not NOT_325(g4050,g3080);
  not NOT_326(g4641,I8838);
  not NOT_327(I11908,g5918);
  not NOT_328(I12757,g6577);
  not NOT_329(g9097,I15681);
  not NOT_330(g2966,g1856);
  not NOT_331(g5794,I10421);
  not NOT_332(I5889,g83);
  not NOT_333(g1643,g1211);
  not NOT_334(I11569,g6279);
  not NOT_335(g7131,g6976);
  not NOT_336(g6344,I11359);
  not NOT_337(g2471,I6309);
  not NOT_338(g7006,I12748);
  not NOT_339(g7331,I13413);
  not NOT_340(I15196,g8778);
  not NOT_341(I6636,g1704);
  not NOT_342(I14732,g8155);
  not NOT_343(g2242,g985);
  not NOT_344(g6207,I10962);
  not NOT_345(g3909,I7520);
  not NOT_346(I11747,g6123);
  not NOT_347(I12564,g6720);
  not NOT_348(g8563,I14662);
  not NOT_349(g2948,g2366);
  not NOT_350(I11242,g6183);
  not NOT_351(g7766,I14169);
  not NOT_352(g6819,I12328);
  not NOT_353(g7105,I12903);
  not NOT_354(g3519,g2185);
  not NOT_355(I10761,g5302);
  not NOT_356(g7305,I13347);
  not NOT_357(I7856,g3805);
  not NOT_358(I7734,g2595);
  not NOT_359(g2955,I6703);
  not NOT_360(g7487,I13649);
  not NOT_361(g5628,g4748);
  not NOT_362(g1742,g1486);
  not NOT_363(g6088,I10708);
  not NOT_364(g6852,I12427);
  not NOT_365(g5515,g4923);
  not NOT_366(I12397,g6764);
  not NOT_367(g6488,I11652);
  not NOT_368(g4658,I8889);
  not NOT_369(g7748,I14115);
  not NOT_370(g4777,I9084);
  not NOT_371(I10400,g5201);
  not NOT_372(g5100,I9484);
  not NOT_373(I9512,g3985);
  not NOT_374(I13807,g7320);
  not NOT_375(I11974,g5956);
  not NOT_376(I12062,g5988);
  not NOT_377(I14400,g7677);
  not NOT_378(g2350,I6166);
  not NOT_379(g9112,I15726);
  not NOT_380(g7755,I14136);
  not NOT_381(g9218,I15930);
  not NOT_382(g1926,g874);
  not NOT_383(I9823,g5138);
  not NOT_384(g9312,I16052);
  not NOT_385(g2038,g809);
  not NOT_386(g4882,g4069);
  not NOT_387(I14214,g7576);
  not NOT_388(I12933,g7018);
  not NOT_389(I9366,g4350);
  not NOT_390(g7226,g6937);
  not NOT_391(I11230,g6140);
  not NOT_392(I11293,g5824);
  not NOT_393(I10207,g5075);
  not NOT_394(I13293,g7159);
  not NOT_395(I12508,g6593);
  not NOT_396(I11638,g5847);
  not NOT_397(g6886,I12529);
  not NOT_398(I6446,g1812);
  not NOT_399(g4611,I8748);
  not NOT_400(g291,I5356);
  not NOT_401(I14005,g7434);
  not NOT_402(g7045,g6490);
  not NOT_403(I11416,g5829);
  not NOT_404(I10538,g5255);
  not NOT_405(I6003,g228);
  not NOT_406(I9148,g4354);
  not NOT_407(I13416,g7165);
  not NOT_408(I5795,g1236);
  not NOT_409(g9129,I15765);
  not NOT_410(g2769,g2424);
  not NOT_411(g7173,g6980);
  not NOT_412(g9329,g9317);
  not NOT_413(g6314,I11269);
  not NOT_414(g7091,g6525);
  not NOT_415(g7491,I13653);
  not NOT_416(g6870,I12481);
  not NOT_417(g3860,I7383);
  not NOT_418(g2918,g2310);
  not NOT_419(g3341,I6936);
  not NOT_420(g1983,I5839);
  not NOT_421(g6825,I12346);
  not NOT_422(g6650,g6213);
  not NOT_423(g7169,I13075);
  not NOT_424(g7283,I13281);
  not NOT_425(g1572,g673);
  not NOT_426(g8955,I15379);
  not NOT_427(I6695,g2246);
  not NOT_428(g4541,g2883);
  not NOT_429(g7059,g6538);
  not NOT_430(g7920,I14282);
  not NOT_431(g7578,I13879);
  not NOT_432(g6008,g5367);
  not NOT_433(I11835,g6181);
  not NOT_434(g3691,I7195);
  not NOT_435(I11014,g5621);
  not NOT_436(g7459,I13617);
  not NOT_437(g9221,I15937);
  not NOT_438(I12205,g6488);
  not NOT_439(I9463,g3942);
  not NOT_440(g7718,I14031);
  not NOT_441(g7767,I14172);
  not NOT_442(g4153,I8024);
  not NOT_443(g4680,I8945);
  not NOT_444(I7688,g3650);
  not NOT_445(g6136,I10773);
  not NOT_446(g4353,g3665);
  not NOT_447(I11586,g6256);
  not NOT_448(I12912,g7006);
  not NOT_449(g6336,I11335);
  not NOT_450(I14100,g7580);
  not NOT_451(I6223,g330);
  not NOT_452(g8038,g7694);
  not NOT_453(g6768,I12173);
  not NOT_454(I8913,g4306);
  not NOT_455(g7582,I13891);
  not NOT_456(g6594,I11796);
  not NOT_457(g1961,g1345);
  not NOT_458(g3879,g2963);
  not NOT_459(g4802,I9129);
  not NOT_460(g7261,I13225);
  not NOT_461(I14683,g7825);
  not NOT_462(g3962,g3131);
  not NOT_463(g5151,I9579);
  not NOT_464(g7793,I14234);
  not NOT_465(g3158,I6853);
  not NOT_466(g3659,g2293);
  not NOT_467(g6806,I12289);
  not NOT_468(g5648,g4748);
  not NOT_469(I6416,g1794);
  not NOT_470(g3506,g1781);
  not NOT_471(g7015,I12763);
  not NOT_472(I12592,g1008);
  not NOT_473(g4558,g2897);
  not NOT_474(g9068,I15598);
  not NOT_475(I7126,g2494);
  not NOT_476(I5926,g297);
  not NOT_477(I7400,g3075);
  not NOT_478(I8859,g3968);
  not NOT_479(I7326,g2940);
  not NOT_480(I6115,g134);
  not NOT_481(I6251,g489);
  not NOT_482(g2921,g2312);
  not NOT_483(g6065,I10684);
  not NOT_484(g6887,I12532);
  not NOT_485(g6122,I10752);
  not NOT_486(I10882,g5600);
  not NOT_487(g6228,I11021);
  not NOT_488(I5754,g966);
  not NOT_489(g3587,g1964);
  not NOT_490(g6322,I11293);
  not NOT_491(I11275,g5768);
  not NOT_492(I9457,g3940);
  not NOT_493(g8918,I15340);
  not NOT_494(I16180,g9387);
  not NOT_495(g6230,I11025);
  not NOT_496(g7246,I13196);
  not NOT_497(g8967,I15405);
  not NOT_498(I13746,g7311);
  not NOT_499(I13493,g7132);
  not NOT_500(I9393,g4266);
  not NOT_501(g4511,g2841);
  not NOT_502(I15660,g9062);
  not NOT_503(g2895,g2268);
  not NOT_504(g6033,g5384);
  not NOT_505(g2837,g1780);
  not NOT_506(g7721,g7344);
  not NOT_507(g5839,I10532);
  not NOT_508(I9834,g4782);
  not NOT_509(g4092,I7899);
  not NOT_510(I13035,g6964);
  not NOT_511(g3985,I7712);
  not NOT_512(I12731,g6579);
  not NOT_513(I11806,g6275);
  not NOT_514(g4600,I8715);
  not NOT_515(I7383,g3465);
  not NOT_516(g4574,g3466);
  not NOT_517(g6096,g5317);
  not NOT_518(g6496,I11662);
  not NOT_519(g1679,I5512);
  not NOT_520(I8097,g3237);
  not NOT_521(g5172,I9642);
  not NOT_522(g5278,I9794);
  not NOT_523(g6845,I12406);
  not NOT_524(g7502,I13682);
  not NOT_525(I15550,g9008);
  not NOT_526(g9198,g9187);
  not NOT_527(g3545,g2344);
  not NOT_528(I8354,g1163);
  not NOT_529(g738,I5404);
  not NOT_530(g6195,I10940);
  not NOT_531(g5618,g5015);
  not NOT_532(g6137,I10776);
  not NOT_533(g6891,I12544);
  not NOT_534(g5143,I9555);
  not NOT_535(g1831,g689);
  not NOT_536(g6337,I11338);
  not NOT_537(g3591,g1789);
  not NOT_538(g3832,I7299);
  not NOT_539(g4580,g2919);
  not NOT_540(g9241,I15971);
  not NOT_541(I7588,g2584);
  not NOT_542(g3853,I7362);
  not NOT_543(I14725,g8145);
  not NOT_544(g7188,I13106);
  not NOT_545(g5988,I10592);
  not NOT_546(g2842,g2209);
  not NOT_547(I9938,g4878);
  not NOT_548(I10758,g5662);
  not NOT_549(g1805,I5667);
  not NOT_550(g6807,I12292);
  not NOT_551(g1916,g775);
  not NOT_552(g5693,I10204);
  not NOT_553(g7216,I13152);
  not NOT_554(g1749,g371);
  not NOT_555(g2298,I6072);
  not NOT_556(I14082,g7539);
  not NOT_557(g6859,I12448);
  not NOT_558(g2392,g11);
  not NOT_559(I13193,g7007);
  not NOT_560(g2485,g62);
  not NOT_561(I11362,g5821);
  not NOT_562(g7028,g6525);
  not NOT_563(I13362,g7265);
  not NOT_564(g3931,I7592);
  not NOT_565(I8218,g3002);
  not NOT_566(I15773,g9126);
  not NOT_567(I6629,g2052);
  not NOT_568(g4623,I8784);
  not NOT_569(g7247,I13199);
  not NOT_570(g1798,I5654);
  not NOT_571(I6130,g560);
  not NOT_572(g4076,I7859);
  not NOT_573(g9319,g9309);
  not NOT_574(I10940,g5489);
  not NOT_575(g2941,g2349);
  not NOT_576(I9606,g4687);
  not NOT_577(g6342,I11353);
  not NOT_578(g3905,g3192);
  not NOT_579(I13475,g7125);
  not NOT_580(g5621,g4748);
  not NOT_581(I14848,g8625);
  not NOT_582(g6255,I11066);
  not NOT_583(g6815,I12316);
  not NOT_584(I10804,g5526);
  not NOT_585(I6800,g2016);
  not NOT_586(I9687,g4822);
  not NOT_587(g3630,I7095);
  not NOT_588(g6481,I11641);
  not NOT_589(I14804,g8563);
  not NOT_590(g7741,I14094);
  not NOT_591(g4651,I8868);
  not NOT_592(g5113,I9499);
  not NOT_593(g6692,I12008);
  not NOT_594(g6097,g5345);
  not NOT_595(I11437,g5801);
  not NOT_596(I15839,g9168);
  not NOT_597(g2520,g41);
  not NOT_598(I15930,g9209);
  not NOT_599(g2640,g1584);
  not NOT_600(g9211,I15909);
  not NOT_601(g6354,I11389);
  not NOT_602(g4285,I8233);
  not NOT_603(I8727,g3944);
  not NOT_604(g9186,I15836);
  not NOT_605(I5679,g911);
  not NOT_606(g4500,g2832);
  not NOT_607(g9386,I16176);
  not NOT_608(g6960,I12681);
  not NOT_609(I15965,g9219);
  not NOT_610(I7944,g3774);
  not NOT_611(g1579,g703);
  not NOT_612(g1869,g74);
  not NOT_613(g7108,I12912);
  not NOT_614(I10135,g4960);
  not NOT_615(g7308,I13356);
  not NOT_616(I11347,g5761);
  not NOT_617(g2958,g2377);
  not NOT_618(I13347,g7224);
  not NOT_619(g9026,I15492);
  not NOT_620(I5831,g1194);
  not NOT_621(g2376,I6226);
  not NOT_622(g5494,I9918);
  not NOT_623(g3750,g2177);
  not NOT_624(I9570,g4696);
  not NOT_625(I10406,g5203);
  not NOT_626(I9341,g4251);
  not NOT_627(I10962,g5719);
  not NOT_628(g1752,g603);
  not NOT_629(I14406,g7681);
  not NOT_630(g3973,g3097);
  not NOT_631(I9525,g4413);
  not NOT_632(I11781,g6284);
  not NOT_633(I12768,g6718);
  not NOT_634(I15619,g8998);
  not NOT_635(g9370,I16138);
  not NOT_636(g1917,I5795);
  not NOT_637(I9645,g4900);
  not NOT_638(I15557,g9010);
  not NOT_639(g2829,g1785);
  not NOT_640(g9125,I15753);
  not NOT_641(g4024,g3160);
  not NOT_642(I11236,g6148);
  not NOT_643(g2286,I6042);
  not NOT_644(g6783,I12220);
  not NOT_645(g7758,I14145);
  not NOT_646(g7066,I12839);
  not NOT_647(I10500,g5234);
  not NOT_648(I16168,g9381);
  not NOT_649(g7589,I13912);
  not NOT_650(I6090,g390);
  not NOT_651(g2911,g2292);
  not NOT_652(g4795,I9116);
  not NOT_653(I8932,g4096);
  not NOT_654(I5422,g1234);
  not NOT_655(g7466,I13622);
  not NOT_656(g4809,I9148);
  not NOT_657(g6267,I11086);
  not NOT_658(g6312,I11263);
  not NOT_659(g3969,g3192);
  not NOT_660(I6166,g480);
  not NOT_661(I14049,g7493);
  not NOT_662(g9280,I16006);
  not NOT_663(I11821,g6170);
  not NOT_664(I12881,g6478);
  not NOT_665(g1786,g623);
  not NOT_666(g7365,I13509);
  not NOT_667(g7048,I12810);
  not NOT_668(I7347,g2985);
  not NOT_669(g9083,I15641);
  not NOT_670(g2270,I6015);
  not NOT_671(g4477,I8517);
  not NOT_672(g7448,I13605);
  not NOT_673(I13063,g6973);
  not NOT_674(g7711,I14012);
  not NOT_675(g4523,g2868);
  not NOT_676(g6676,I11984);
  not NOT_677(I11790,g6282);
  not NOT_678(g6293,I11206);
  not NOT_679(I13264,g7061);
  not NOT_680(I6148,g5);
  not NOT_681(g7055,g6517);
  not NOT_682(g8219,I14436);
  not NOT_683(g4643,I8844);
  not NOT_684(g3666,g2134);
  not NOT_685(I9158,g4256);
  not NOT_686(I13137,g7027);
  not NOT_687(I6348,g1354);
  not NOT_688(g2225,I5948);
  not NOT_689(g6129,I10758);
  not NOT_690(g8640,I14728);
  not NOT_691(g7455,I13613);
  not NOT_692(g6329,I11314);
  not NOT_693(g6761,I12154);
  not NOT_694(g2073,g1254);
  not NOT_695(g5160,I9606);
  not NOT_696(g7133,I12983);
  not NOT_697(I7697,g3052);
  not NOT_698(g9106,I15708);
  not NOT_699(g7333,I13419);
  not NOT_700(I13873,g7342);
  not NOT_701(g9306,I16036);
  not NOT_702(g6828,I12355);
  not NOT_703(g1770,g606);
  not NOT_704(g7774,I14193);
  not NOT_705(g5521,g4929);
  not NOT_706(g8958,I15388);
  not NOT_707(g6830,I12361);
  not NOT_708(g4634,I8817);
  not NOT_709(g3648,g2424);
  not NOT_710(g3875,g2958);
  not NOT_711(g2324,I6115);
  not NOT_712(g3530,g2185);
  not NOT_713(I9111,g4232);
  not NOT_714(g7196,I13122);
  not NOT_715(g4742,I9064);
  not NOT_716(g9061,I15577);
  not NOT_717(I15601,g8992);
  not NOT_718(g9187,I15839);
  not NOT_719(g4104,I7925);
  not NOT_720(I10605,g5440);
  not NOT_721(I11422,g5842);
  not NOT_722(g6592,I11790);
  not NOT_723(g3655,g1844);
  not NOT_724(I15187,g8682);
  not NOT_725(I14273,g7631);
  not NOT_726(I11209,g6139);
  not NOT_727(I13422,g7131);
  not NOT_728(I14106,g7586);
  not NOT_729(I13209,g6912);
  not NOT_730(g2540,g1339);
  not NOT_731(I9615,g4739);
  not NOT_732(g6221,I11004);
  not NOT_733(I12003,g6202);
  not NOT_734(g8765,g8524);
  not NOT_735(g7538,I13794);
  not NOT_736(I13834,g7466);
  not NOT_737(I6463,g1769);
  not NOT_738(I10463,g5220);
  not NOT_739(I16084,g9324);
  not NOT_740(g2177,g1322);
  not NOT_741(g7780,I14211);
  not NOT_742(g9027,I15495);
  not NOT_743(g5724,g4969);
  not NOT_744(g2377,I6229);
  not NOT_745(I14463,g8072);
  not NOT_746(I12779,g6740);
  not NOT_747(g5179,I9663);
  not NOT_748(g6703,I12041);
  not NOT_749(g7509,I13707);
  not NOT_750(g4926,g4202);
  not NOT_751(I15937,g9212);
  not NOT_752(g9200,g9189);
  not NOT_753(I11021,g5627);
  not NOT_754(I14234,g7614);
  not NOT_755(g3884,I7417);
  not NOT_756(g3839,I7320);
  not NOT_757(g2287,I6045);
  not NOT_758(g7018,I12768);
  not NOT_759(g4273,I8215);
  not NOT_760(g7067,g6658);
  not NOT_761(g8974,I15426);
  not NOT_762(I7317,g2893);
  not NOT_763(g5658,g4748);
  not NOT_764(I15791,g9140);
  not NOT_765(g7418,I13533);
  not NOT_766(g6624,I11864);
  not NOT_767(g7467,g7236);
  not NOT_768(g6953,g6745);
  not NOT_769(I6118,g243);
  not NOT_770(I14795,g8604);
  not NOT_771(g8225,I14454);
  not NOT_772(g5835,I10528);
  not NOT_773(g7290,I13302);
  not NOT_774(g4613,I8754);
  not NOT_775(g6068,I10687);
  not NOT_776(g1888,g781);
  not NOT_777(I6872,g2185);
  not NOT_778(g9145,I15791);
  not NOT_779(g4044,g2595);
  not NOT_780(g6468,I11622);
  not NOT_781(I12945,g7066);
  not NOT_782(I9591,g4710);
  not NOT_783(g4444,I8452);
  not NOT_784(g1787,g625);
  not NOT_785(I6652,g2016);
  not NOT_786(I11607,g5767);
  not NOT_787(I6057,g518);
  not NOT_788(I12826,g6441);
  not NOT_789(I12999,g7029);
  not NOT_790(I11320,g5797);
  not NOT_791(I15666,g9070);
  not NOT_792(I13320,g7139);
  not NOT_793(I6457,g1886);
  not NOT_794(g7493,I13659);
  not NOT_795(g1675,g1519);
  not NOT_796(g6677,I11987);
  not NOT_797(g7256,g7058);
  not NOT_798(I13274,g6917);
  not NOT_799(I7775,g3705);
  not NOT_800(g5611,g4969);
  not NOT_801(g8324,I14573);
  not NOT_802(g4572,g2909);
  not NOT_803(I7922,g3462);
  not NOT_804(g2898,g2271);
  not NOT_805(I15478,g8910);
  not NOT_806(g2900,g2273);
  not NOT_807(g6866,I12469);
  not NOT_808(I12672,g6473);
  not NOT_809(I7581,g3612);
  not NOT_810(I13122,g7070);
  not NOT_811(g9107,I15711);
  not NOT_812(g4543,g2885);
  not NOT_813(I10421,g5208);
  not NOT_814(I11464,g6088);
  not NOT_815(g5799,I10436);
  not NOT_816(I13565,g7181);
  not NOT_817(I9794,g4778);
  not NOT_818(I6834,g287);
  not NOT_819(g9307,g9300);
  not NOT_820(g2510,g58);
  not NOT_821(g639,I5374);
  not NOT_822(g2245,g999);
  not NOT_823(g6149,I10810);
  not NOT_824(g3988,g3097);
  not NOT_825(I6686,g2246);
  not NOT_826(g6349,I11374);
  not NOT_827(g5674,g5042);
  not NOT_828(g8177,I14410);
  not NOT_829(g3693,g2424);
  not NOT_830(I11034,g5644);
  not NOT_831(g9223,I15943);
  not NOT_832(I14163,g7533);
  not NOT_833(g2291,I6057);
  not NOT_834(I14012,g7438);
  not NOT_835(I11641,g5918);
  not NOT_836(g6848,I12415);
  not NOT_837(I15580,g8985);
  not NOT_838(I13797,g7502);
  not NOT_839(I12331,g6704);
  not NOT_840(g5541,g4814);
  not NOT_841(g3548,g2185);
  not NOT_842(g1684,g1);
  not NOT_843(g1745,g746);
  not NOT_844(g6198,g5335);
  not NOT_845(g1639,g1207);
  not NOT_846(g2344,I6148);
  not NOT_847(g6855,I12436);
  not NOT_848(g6398,I11515);
  not NOT_849(I10541,g5256);
  not NOT_850(I6121,g321);
  not NOT_851(g7263,I13231);
  not NOT_852(g2207,I5920);
  not NOT_853(g5153,I9585);
  not NOT_854(g5680,g5101);
  not NOT_855(I12897,g6962);
  not NOT_856(I12448,g6569);
  not NOT_857(I12961,g6921);
  not NOT_858(I9515,g4301);
  not NOT_859(I9630,g4867);
  not NOT_860(I14789,g8544);
  not NOT_861(g2259,g1325);
  not NOT_862(g9115,I15735);
  not NOT_863(g4014,I7769);
  not NOT_864(I7079,g2532);
  not NOT_865(I12505,g6612);
  not NOT_866(g9315,I16061);
  not NOT_867(g1808,g629);
  not NOT_868(g4885,g4070);
  not NOT_869(I13635,g7243);
  not NOT_870(g5744,I10289);
  not NOT_871(g8199,I14424);
  not NOT_872(g9047,I15543);
  not NOT_873(g5802,I10445);
  not NOT_874(g4660,I8895);
  not NOT_875(g2923,I6657);
  not NOT_876(I12717,g6543);
  not NOT_877(g1707,g955);
  not NOT_878(I14325,g7713);
  not NOT_879(I10829,g5224);
  not NOT_880(g8781,g8585);
  not NOT_881(I10535,g5254);
  not NOT_882(I5389,g690);
  not NOT_883(I5706,g901);
  not NOT_884(g8898,I15308);
  not NOT_885(g4903,g4084);
  not NOT_886(g7562,I13858);
  not NOT_887(I15178,g8753);
  not NOT_888(I10946,g5563);
  not NOT_889(g8797,I15003);
  not NOT_890(g6524,I11710);
  not NOT_891(I14828,g8639);
  not NOT_892(g6644,g6208);
  not NOT_893(g8510,I14643);
  not NOT_894(I13164,g7086);
  not NOT_895(I5371,g633);
  not NOT_896(g7723,I14042);
  not NOT_897(I14121,g7587);
  not NOT_898(g2215,g1416);
  not NOT_899(I15953,g9215);
  not NOT_900(g6319,I11284);
  not NOT_901(g7101,I12891);
  not NOT_902(g2886,g2240);
  not NOT_903(g3908,I7517);
  not NOT_904(g7301,I13335);
  not NOT_905(I7356,g2843);
  not NOT_906(I13891,g7336);
  not NOT_907(I15654,g9057);
  not NOT_908(g4036,g3192);
  not NOT_909(g6152,I10815);
  not NOT_910(g6258,g5427);
  not NOT_911(g6352,I11383);
  not NOT_912(g6818,I12325);
  not NOT_913(g1575,g685);
  not NOT_914(g1865,g1013);
  not NOT_915(I8483,g3641);
  not NOT_916(g6867,I12472);
  not NOT_917(g3567,g2407);
  not NOT_918(I15417,g8893);
  not NOT_919(g1715,I5559);
  not NOT_920(g2314,I6099);
  not NOT_921(I9440,g4285);
  not NOT_922(I14291,g7680);
  not NOT_923(I12433,g6632);
  not NOT_924(g4335,g3659);
  not NOT_925(I9123,g4455);
  not NOT_926(I15334,g8800);
  not NOT_927(g7751,I14124);
  not NOT_928(g2870,g2225);
  not NOT_929(g5492,g4919);
  not NOT_930(I12148,g5988);
  not NOT_931(I13109,g7059);
  not NOT_932(g4382,I8373);
  not NOT_933(g1833,g770);
  not NOT_934(g5600,g5128);
  not NOT_935(I13537,g7152);
  not NOT_936(g5574,g4969);
  not NOT_937(I8790,g4020);
  not NOT_938(g6211,g5645);
  not NOT_939(g2825,I6553);
  not NOT_940(g2650,I6434);
  not NOT_941(g6186,I10919);
  not NOT_942(g6386,I11485);
  not NOT_943(I12646,g6493);
  not NOT_944(g7585,I13900);
  not NOT_945(g9017,I15475);
  not NOT_946(I9666,g4931);
  not NOT_947(I15762,g9039);
  not NOT_948(I12343,g6731);
  not NOT_949(g4805,I9136);
  not NOT_950(g6975,I12712);
  not NOT_951(g4916,g4202);
  not NOT_952(g4022,I7785);
  not NOT_953(g3965,I7676);
  not NOT_954(I5963,g225);
  not NOT_955(g1584,g738);
  not NOT_956(g6599,I11809);
  not NOT_957(g1896,g86);
  not NOT_958(g7441,I13580);
  not NOT_959(I15423,g8894);
  not NOT_960(g6026,g5384);
  not NOT_961(I9528,g4006);
  not NOT_962(g6426,I11559);
  not NOT_963(I6860,g2185);
  not NOT_964(g3264,I6900);
  not NOT_965(I7053,g2452);
  not NOT_966(I6341,g1351);
  not NOT_967(I10506,g5236);
  not NOT_968(g5580,g4938);
  not NOT_969(I9648,g4795);
  not NOT_970(g9234,I15956);
  not NOT_971(I10028,g4825);
  not NOT_972(g9128,I15762);
  not NOT_973(g6614,I11838);
  not NOT_974(g6370,I11437);
  not NOT_975(I14028,g7501);
  not NOT_976(g3933,g3131);
  not NOT_977(I8904,g4126);
  not NOT_978(g9330,g9319);
  not NOT_979(g6325,I11302);
  not NOT_980(g6821,I12334);
  not NOT_981(g3521,g2185);
  not NOT_982(g4560,g2899);
  not NOT_983(I8446,g3014);
  not NOT_984(g3050,I6788);
  not NOT_985(g3641,I7115);
  not NOT_986(I15909,g9201);
  not NOT_987(I15543,g9006);
  not NOT_988(g5736,I10265);
  not NOT_989(g2943,g2362);
  not NOT_990(g6984,I12725);
  not NOT_991(g7168,I13072);
  not NOT_992(g6939,g6543);
  not NOT_993(g3996,I7731);
  not NOT_994(I11796,g6287);
  not NOT_995(I12412,g6404);
  not NOT_996(I8841,g3979);
  not NOT_997(g5623,g4969);
  not NOT_998(g7772,I14187);
  not NOT_999(g6083,I10702);
  not NOT_1000(g7058,g6649);
  not NOT_1001(I5957,g110);
  not NOT_1002(g2887,g2241);
  not NOT_1003(g4873,I9217);
  not NOT_1004(g4632,I8811);
  not NOT_1005(g7531,I13773);
  not NOT_1006(g4095,I7908);
  not NOT_1007(g5076,I9446);
  not NOT_1008(g8870,I15196);
  not NOT_1009(I8763,g3947);
  not NOT_1010(g4037,g2845);
  not NOT_1011(g6483,I11645);
  not NOT_1012(I12229,g6659);
  not NOT_1013(I9884,g4868);
  not NOT_1014(g2934,I6676);
  not NOT_1015(g5476,g4907);
  not NOT_1016(g7743,I14100);
  not NOT_1017(g4653,I8874);
  not NOT_1018(I6358,g13);
  not NOT_1019(g4102,I7919);
  not NOT_1020(g6636,I11900);
  not NOT_1021(I15568,g8981);
  not NOT_1022(I15747,g9042);
  not NOT_1023(I5865,g1206);
  not NOT_1024(g9213,I15915);
  not NOT_1025(g6106,g5345);
  not NOT_1026(g5175,I9651);
  not NOT_1027(g4579,g2918);
  not NOT_1028(I10649,g5657);
  not NOT_1029(I12011,g5939);
  not NOT_1030(g6306,I11245);
  not NOT_1031(I5715,g896);
  not NOT_1032(g7505,I13695);
  not NOT_1033(g5871,I10558);
  not NOT_1034(g3878,g2962);
  not NOT_1035(g8008,g7559);
  not NOT_1036(g4719,I9021);
  not NOT_1037(g6790,I12241);
  not NOT_1038(g7734,I14073);
  not NOT_1039(I6587,g1708);
  not NOT_1040(g3777,g2170);
  not NOT_1041(g7411,g7202);
  not NOT_1042(I9372,g3902);
  not NOT_1043(I10491,g5231);
  not NOT_1044(I15814,g9154);
  not NOT_1045(g3835,I7308);
  not NOT_1046(I16116,g9350);
  not NOT_1047(g6387,I11488);
  not NOT_1048(I11522,g5847);
  not NOT_1049(g2096,g1226);
  not NOT_1050(I9618,g4742);
  not NOT_1051(I12582,g6745);
  not NOT_1052(g5285,g4841);
  not NOT_1053(g6461,I11607);
  not NOT_1054(g8768,g8585);
  not NOT_1055(I13663,g7235);
  not NOT_1056(g3882,g2970);
  not NOT_1057(g2496,g942);
  not NOT_1058(I7626,g3632);
  not NOT_1059(g4917,g4102);
  not NOT_1060(I15974,g9234);
  not NOT_1061(I6615,g1983);
  not NOT_1062(g6756,I12141);
  not NOT_1063(g8972,I15420);
  not NOT_1064(I10770,g5441);
  not NOT_1065(I12310,g6723);
  not NOT_1066(g1897,g789);
  not NOT_1067(g9090,I15660);
  not NOT_1068(g6622,I11858);
  not NOT_1069(g7474,I13628);
  not NOT_1070(I8757,g3921);
  not NOT_1071(g6027,g5384);
  not NOT_1072(g7992,g7557);
  not NOT_1073(g4265,g3591);
  not NOT_1074(g3611,I7079);
  not NOT_1075(g6427,I11562);
  not NOT_1076(g2137,I5889);
  not NOT_1077(g2891,g2265);
  not NOT_1078(g5184,I9678);
  not NOT_1079(I15638,g8978);
  not NOT_1080(g9366,I16126);
  not NOT_1081(g2913,g2307);
  not NOT_1082(I12379,g6768);
  not NOT_1083(g5139,I9543);
  not NOT_1084(g5384,I9837);
  not NOT_1085(g6904,g6426);
  not NOT_1086(I12958,g6920);
  not NOT_1087(g9056,I15562);
  not NOT_1088(g8065,I14338);
  not NOT_1089(I8315,g3691);
  not NOT_1090(I8811,g4022);
  not NOT_1091(g6446,I11591);
  not NOT_1092(g8228,I14463);
  not NOT_1093(g3981,I7706);
  not NOT_1094(g5024,I9360);
  not NOT_1095(g6514,I11696);
  not NOT_1096(I6239,g8);
  not NOT_1097(g3674,I7164);
  not NOT_1098(g2807,g1782);
  not NOT_1099(I5362,g3841);
  not NOT_1100(I11326,g5819);
  not NOT_1101(I9555,g4892);
  not NOT_1102(g5795,I10424);
  not NOT_1103(g5737,I10268);
  not NOT_1104(I15391,g8917);
  not NOT_1105(g6403,I11522);
  not NOT_1106(I13326,g7176);
  not NOT_1107(g5809,I10460);
  not NOT_1108(I5419,g1603);
  not NOT_1109(I9804,g5113);
  not NOT_1110(I10262,g5551);
  not NOT_1111(I7683,g2573);
  not NOT_1112(g3997,I7734);
  not NOT_1113(I12742,g6590);
  not NOT_1114(g6345,I11362);
  not NOT_1115(g6841,I12394);
  not NOT_1116(I15510,g8969);
  not NOT_1117(I11040,g5299);
  not NOT_1118(I11948,g5897);
  not NOT_1119(I8874,g3884);
  not NOT_1120(g2266,I6003);
  not NOT_1121(g6763,I12158);
  not NOT_1122(I7778,g3019);
  not NOT_1123(I16142,g9366);
  not NOT_1124(g6391,I11500);
  not NOT_1125(g1006,I5410);
  not NOT_1126(g4296,g3790);
  not NOT_1127(I6853,g2185);
  not NOT_1128(g3238,I6894);
  not NOT_1129(I9621,g4732);
  not NOT_1130(g5477,g4908);
  not NOT_1131(g9260,I15990);
  not NOT_1132(g5523,I9935);
  not NOT_1133(I12681,g6469);
  not NOT_1134(I10719,g5559);
  not NOT_1135(g6637,I11903);
  not NOT_1136(g5643,I10128);
  not NOT_1137(I15014,g8607);
  not NOT_1138(g1801,g618);
  not NOT_1139(g4553,g2891);
  not NOT_1140(g9063,I15583);
  not NOT_1141(g6307,I11248);
  not NOT_1142(I15586,g8987);
  not NOT_1143(I15007,g8627);
  not NOT_1144(I8880,g4303);
  not NOT_1145(I14718,g8068);
  not NOT_1146(g3802,g1832);
  not NOT_1147(g7688,g7406);
  not NOT_1148(g6359,I11404);
  not NOT_1149(g6223,I11008);
  not NOT_1150(g2481,I6317);
  not NOT_1151(g8913,I15329);
  not NOT_1152(g1748,g601);
  not NOT_1153(g2692,g1671);
  not NOT_1154(g4012,I7765);
  not NOT_1155(g6858,I12445);
  not NOT_1156(g5742,I10283);
  not NOT_1157(g5551,I9974);
  not NOT_1158(g5099,g4477);
  not NOT_1159(g2497,g945);
  not NOT_1160(I12690,g6467);
  not NOT_1161(g2354,I6178);
  not NOT_1162(I16165,g9377);
  not NOT_1163(g2960,g2381);
  not NOT_1164(g4706,I9005);
  not NOT_1165(I9567,g4693);
  not NOT_1166(I7526,g2752);
  not NOT_1167(I5897,g173);
  not NOT_1168(I14573,g8179);
  not NOT_1169(I10247,g5266);
  not NOT_1170(g3901,I7492);
  not NOT_1171(g7000,I12742);
  not NOT_1172(I13509,g7137);
  not NOT_1173(I15720,g9053);
  not NOT_1174(g9318,g9304);
  not NOT_1175(g9367,I16129);
  not NOT_1176(I11933,g5847);
  not NOT_1177(g7126,I12968);
  not NOT_1178(I8935,g4005);
  not NOT_1179(I5425,g1245);
  not NOT_1180(g4029,I7800);
  not NOT_1181(g6251,I11060);
  not NOT_1182(g6315,I11272);
  not NOT_1183(g6811,I12304);
  not NOT_1184(g6642,I11912);
  not NOT_1185(g4371,I8354);
  not NOT_1186(I11851,g6277);
  not NOT_1187(g3511,g1616);
  not NOT_1188(g5754,g5403);
  not NOT_1189(g9057,I15565);
  not NOT_1190(I16006,g9261);
  not NOT_1191(g7760,I14151);
  not NOT_1192(I14388,g7605);
  not NOT_1193(I7850,g2795);
  not NOT_1194(g9193,g9181);
  not NOT_1195(g3092,I6826);
  not NOT_1196(I14777,g8511);
  not NOT_1197(g3492,I6970);
  not NOT_1198(g4281,g2562);
  not NOT_1199(g6874,I12493);
  not NOT_1200(g5613,g4748);
  not NOT_1201(I14251,g7541);
  not NOT_1202(g3574,g1771);
  not NOT_1203(g3864,g2943);
  not NOT_1204(g8342,g8008);
  not NOT_1205(I15340,g8856);
  not NOT_1206(g2267,I6006);
  not NOT_1207(g2312,I6093);
  not NOT_1208(g6654,I11942);
  not NOT_1209(g5444,g5074);
  not NOT_1210(g5269,I9791);
  not NOT_1211(I7702,g3062);
  not NOT_1212(I15684,g9067);
  not NOT_1213(g8481,I14637);
  not NOT_1214(I12128,g5897);
  not NOT_1215(g1578,g699);
  not NOT_1216(g1868,I5747);
  not NOT_1217(I9360,g4257);
  not NOT_1218(g2401,g22);
  not NOT_1219(I7919,g3761);
  not NOT_1220(I10032,g1236);
  not NOT_1221(g1718,I5562);
  not NOT_1222(g7779,I14208);
  not NOT_1223(g2293,g888);
  not NOT_1224(g6880,I12511);
  not NOT_1225(g4684,I8949);
  not NOT_1226(I9050,g3881);
  not NOT_1227(I11452,g6071);
  not NOT_1228(g6595,g6083);
  not NOT_1229(g4639,I8832);
  not NOT_1230(I5682,g168);
  not NOT_1231(I5766,g1254);
  not NOT_1232(I11047,g5653);
  not NOT_1233(I13574,g7205);
  not NOT_1234(g2329,I6130);
  not NOT_1235(I6440,g1806);
  not NOT_1236(g7023,I12779);
  not NOT_1237(g9121,I15747);
  not NOT_1238(g4963,g4328);
  not NOT_1239(g2761,g1820);
  not NOT_1240(I5801,g1424);
  not NOT_1241(g9321,g9311);
  not NOT_1242(g8960,I15394);
  not NOT_1243(g7423,I13544);
  not NOT_1244(g1582,g714);
  not NOT_1245(I11912,g5897);
  not NOT_1246(I11311,g5760);
  not NOT_1247(I13912,g7359);
  not NOT_1248(I13311,g7162);
  not NOT_1249(g2828,g1980);
  not NOT_1250(I12298,g6697);
  not NOT_1251(I6323,g1342);
  not NOT_1252(I14061,g7546);
  not NOT_1253(g1793,g626);
  not NOT_1254(I7561,g2562);
  not NOT_1255(g7588,I13909);
  not NOT_1256(I10766,g5674);
  not NOT_1257(g2727,g2424);
  not NOT_1258(g4808,I9145);
  not NOT_1259(g6978,I12717);
  not NOT_1260(g6612,I11832);
  not NOT_1261(g7161,I13057);
  not NOT_1262(g1015,I5416);
  not NOT_1263(g5729,g5144);
  not NOT_1264(g3968,I7683);
  not NOT_1265(g6243,I11050);
  not NOT_1266(g7361,I13499);
  not NOT_1267(I15193,g8774);
  not NOT_1268(I13051,g6967);
  not NOT_1269(I13072,g6969);
  not NOT_1270(g2746,g2259);
  not NOT_1271(I12737,g6460);
  not NOT_1272(g2221,I5936);
  not NOT_1273(g3076,g1831);
  not NOT_1274(g7127,g6974);
  not NOT_1275(g8783,g8524);
  not NOT_1276(g7327,I13403);
  not NOT_1277(I12232,g6662);
  not NOT_1278(g1664,g1462);
  not NOT_1279(I6151,g12);
  not NOT_1280(g1246,I5425);
  not NOT_1281(g2703,g1809);
  not NOT_1282(g8218,I14433);
  not NOT_1283(I8823,g3965);
  not NOT_1284(g5014,I9344);
  not NOT_1285(g206,I5353);
  not NOT_1286(g6328,I11311);
  not NOT_1287(g6130,I10761);
  not NOT_1288(g7146,g6998);
  not NOT_1289(g6542,I11718);
  not NOT_1290(g6330,I11317);
  not NOT_1291(g7346,I13454);
  not NOT_1292(g7633,I13962);
  not NOT_1293(g1721,I5565);
  not NOT_1294(I11350,g5763);
  not NOT_1295(g3871,g2953);
  not NOT_1296(I7970,g3557);
  not NOT_1297(I13350,g7223);
  not NOT_1298(I15475,g8901);
  not NOT_1299(g2932,g2329);
  not NOT_1300(g7103,I12897);
  not NOT_1301(I9271,g4263);
  not NOT_1302(g3651,I7129);
  not NOT_1303(g7303,I13341);
  not NOT_1304(I7925,g2761);
  not NOT_1305(g8676,I14822);
  not NOT_1306(g2624,g1569);
  not NOT_1307(g2953,g2373);
  not NOT_1308(I15222,g8834);
  not NOT_1309(g6800,I12271);
  not NOT_1310(g3285,g1689);
  not NOT_1311(I13152,g6966);
  not NOT_1312(g8761,g8564);
  not NOT_1313(g4604,I8727);
  not NOT_1314(I10451,g5216);
  not NOT_1315(I10472,g5223);
  not NOT_1316(I13846,g7487);
  not NOT_1317(g3500,g1616);
  not NOT_1318(I14451,g8172);
  not NOT_1319(g7732,I14067);
  not NOT_1320(I5407,g4653);
  not NOT_1321(I13731,g7441);
  not NOT_1322(I5920,g219);
  not NOT_1323(I6839,g2185);
  not NOT_1324(I5868,g74);
  not NOT_1325(I7320,g2927);
  not NOT_1326(g2677,g1664);
  not NOT_1327(g7753,I14130);
  not NOT_1328(g5178,I9660);
  not NOT_1329(g5679,I10172);
  not NOT_1330(I11413,g5871);
  not NOT_1331(I5718,g896);
  not NOT_1332(g7508,I13704);
  not NOT_1333(I13413,g7127);
  not NOT_1334(g6213,I10976);
  not NOT_1335(I5535,g48);
  not NOT_1336(g2866,g2221);
  not NOT_1337(g4584,g3466);
  not NOT_1338(I12445,g6568);
  not NOT_1339(g4539,g2881);
  not NOT_1340(g8746,g8524);
  not NOT_1341(g8221,I14442);
  not NOT_1342(g5335,g4677);
  not NOT_1343(g5831,I10516);
  not NOT_1344(g3838,I7317);
  not NOT_1345(g1689,g855);
  not NOT_1346(g2149,I5894);
  not NOT_1347(g2349,I6163);
  not NOT_1348(I12499,g6597);
  not NOT_1349(g7043,g6543);
  not NOT_1350(g9141,g9129);
  not NOT_1351(g5182,I9672);
  not NOT_1352(I10776,g5576);
  not NOT_1353(I12316,g6736);
  not NOT_1354(I9132,g4284);
  not NOT_1355(I6143,g1217);
  not NOT_1356(I9209,g4349);
  not NOT_1357(g7116,I12936);
  not NOT_1358(g1671,g1494);
  not NOT_1359(I7987,g3528);
  not NOT_1360(g5805,I10448);
  not NOT_1361(g5916,g5384);
  not NOT_1362(g5022,g4438);
  not NOT_1363(g2699,g1674);
  not NOT_1364(g4019,I7778);
  not NOT_1365(g6090,g5529);
  not NOT_1366(g4362,g2810);
  not NOT_1367(I11929,g6190);
  not NOT_1368(I12989,g6932);
  not NOT_1369(g3077,I6805);
  not NOT_1370(g7034,g6525);
  not NOT_1371(g5749,g5207);
  not NOT_1372(g6490,I11656);
  not NOT_1373(g6823,I12340);
  not NOT_1374(g7434,I13565);
  not NOT_1375(I14825,g8651);
  not NOT_1376(g3523,g2407);
  not NOT_1377(I14370,g7603);
  not NOT_1378(g6366,I11425);
  not NOT_1379(I12722,g6611);
  not NOT_1380(g7565,I13865);
  not NOT_1381(I7299,g2961);
  not NOT_1382(I5664,g916);
  not NOT_1383(g3643,g2453);
  not NOT_1384(I12924,g6983);
  not NOT_1385(I13583,g7252);
  not NOT_1386(g2241,I5984);
  not NOT_1387(g1564,g642);
  not NOT_1388(g7147,g6904);
  not NOT_1389(I16122,g9353);
  not NOT_1390(I10151,g5007);
  not NOT_1391(I10172,g4873);
  not NOT_1392(g7347,I13457);
  not NOT_1393(I15516,g8977);
  not NOT_1394(I9558,g4597);
  not NOT_1395(g5798,I10433);
  not NOT_1396(I14151,g7555);
  not NOT_1397(g1826,g632);
  not NOT_1398(I12271,g6663);
  not NOT_1399(I14172,g7545);
  not NOT_1400(g6148,I10807);
  not NOT_1401(g6649,I11929);
  not NOT_1402(I14996,g8510);
  not NOT_1403(g6348,I11371);
  not NOT_1404(I8989,g4537);
  not NOT_1405(g8677,I14825);
  not NOT_1406(g7533,I13779);
  not NOT_1407(g3634,I7107);
  not NOT_1408(I8193,g3547);
  not NOT_1409(g6155,I10826);
  not NOT_1410(I14844,g8641);
  not NOT_1411(g6851,I12424);
  not NOT_1412(g6355,I11392);
  not NOT_1413(I11787,g6273);
  not NOT_1414(I14394,g7536);
  not NOT_1415(I12753,g6445);
  not NOT_1416(g8866,I15184);
  not NOT_1417(g7210,I13144);
  not NOT_1418(g2644,I6416);
  not NOT_1419(g3499,g2185);
  not NOT_1420(I8971,g4464);
  not NOT_1421(I12145,g5971);
  not NOT_1422(g1638,g1092);
  not NOT_1423(I11302,g5796);
  not NOT_1424(I7738,g3038);
  not NOT_1425(g5873,g5367);
  not NOT_1426(I13302,g7164);
  not NOT_1427(g5037,g4438);
  not NOT_1428(g9111,I15723);
  not NOT_1429(I12199,g6475);
  not NOT_1430(g7013,I12757);
  not NOT_1431(g9311,I16049);
  not NOT_1432(g5437,g5041);
  not NOT_1433(I11827,g6231);
  not NOT_1434(g5653,g4748);
  not NOT_1435(g7413,I13524);
  not NOT_1436(I13743,g7454);
  not NOT_1437(g3926,I7581);
  not NOT_1438(g5302,g5028);
  not NOT_1439(I14420,g7554);
  not NOT_1440(I15208,g8810);
  not NOT_1441(g2818,g1792);
  not NOT_1442(g6063,I10678);
  not NOT_1443(g4070,I7847);
  not NOT_1444(I12529,g6628);
  not NOT_1445(g2867,g2222);
  not NOT_1446(g3754,g2543);
  not NOT_1447(I9600,g4698);
  not NOT_1448(g8198,g7721);
  not NOT_1449(g8747,g8545);
  not NOT_1450(g4025,I7792);
  not NOT_1451(I14318,g7657);
  not NOT_1452(g5719,I10236);
  not NOT_1453(I12696,g6503);
  not NOT_1454(g9374,I16148);
  not NOT_1455(I14227,g7552);
  not NOT_1456(I5689,g906);
  not NOT_1457(I7959,g2793);
  not NOT_1458(g1758,g1084);
  not NOT_1459(g1589,g746);
  not NOT_1460(I14025,g7500);
  not NOT_1461(I7517,g3578);
  not NOT_1462(I11803,g6280);
  not NOT_1463(I7082,g2470);
  not NOT_1464(g2893,I6615);
  not NOT_1465(I15726,g9069);
  not NOT_1466(g7117,I12939);
  not NOT_1467(g6279,I11132);
  not NOT_1468(g5917,g5412);
  not NOT_1469(g7317,I13383);
  not NOT_1470(I14058,g7544);
  not NOT_1471(g6720,g6254);
  not NOT_1472(I5428,g49);
  not NOT_1473(g6118,g5549);
  not NOT_1474(g6167,I10862);
  not NOT_1475(g6318,I11281);
  not NOT_1476(g1571,g669);
  not NOT_1477(g3983,g2845);
  not NOT_1478(g6367,I11428);
  not NOT_1479(g9180,I15824);
  not NOT_1480(g6872,I12487);
  not NOT_1481(g7601,g7450);
  not NOT_1482(I15607,g8994);
  not NOT_1483(g9380,g9379);
  not NOT_1484(g3862,I7389);
  not NOT_1485(g5042,I9396);
  not NOT_1486(g1711,I5555);
  not NOT_1487(g2274,g782);
  not NOT_1488(g6652,I11936);
  not NOT_1489(I12161,g5971);
  not NOT_1490(g4678,I8935);
  not NOT_1491(g3712,g1952);
  not NOT_1492(g8524,g7855);
  not NOT_1493(g6843,I12400);
  not NOT_1494(I15530,g8972);
  not NOT_1495(g5786,I10403);
  not NOT_1496(g4006,I7749);
  not NOT_1497(g2170,g1229);
  not NOT_1498(g1827,g762);
  not NOT_1499(g2614,g1562);
  not NOT_1500(g9020,I15484);
  not NOT_1501(g7775,I14196);
  not NOT_1502(g5164,I9618);
  not NOT_1503(g6393,I11506);
  not NOT_1504(g4635,I8820);
  not NOT_1505(g5364,g5124);
  not NOT_1506(I15565,g8980);
  not NOT_1507(g2325,I6118);
  not NOT_1508(g2821,g1786);
  not NOT_1509(I12259,g6652);
  not NOT_1510(I10377,g5188);
  not NOT_1511(g1774,I5616);
  not NOT_1512(I12708,g6482);
  not NOT_1513(g7581,I13888);
  not NOT_1514(I11662,g5956);
  not NOT_1515(I10739,g5572);
  not NOT_1516(g4087,I7882);
  not NOT_1517(g4105,I7928);
  not NOT_1518(g8152,I14388);
  not NOT_1519(I9076,g4353);
  not NOT_1520(g5054,g4457);
  not NOT_1521(g6834,I12373);
  not NOT_1522(g4801,I9126);
  not NOT_1523(g8867,I15187);
  not NOT_1524(I9889,g4819);
  not NOT_1525(I14739,g8173);
  not NOT_1526(g2939,g2348);
  not NOT_1527(g3961,g3131);
  not NOT_1528(g7060,g6654);
  not NOT_1529(I11890,g6135);
  not NOT_1530(g1803,g758);
  not NOT_1531(g7460,g7172);
  not NOT_1532(I15641,g9017);
  not NOT_1533(I6160,g324);
  not NOT_1534(g5725,g4841);
  not NOT_1535(g4748,g4465);
  not NOT_1536(I11482,g6117);
  not NOT_1537(g6598,I11806);
  not NOT_1538(g3927,I7584);
  not NOT_1539(I5609,g16);
  not NOT_1540(I11248,g6149);
  not NOT_1541(g1780,g614);
  not NOT_1542(I12244,g6642);
  not NOT_1543(I11710,g6098);
  not NOT_1544(I13710,g7340);
  not NOT_1545(g2636,g1580);
  not NOT_1546(g7739,I14088);
  not NOT_1547(g3014,I6767);
  not NOT_1548(I9651,g4805);
  not NOT_1549(g6321,I11290);
  not NOT_1550(g4226,g3591);
  not NOT_1551(g8386,g8014);
  not NOT_1552(I5883,g80);
  not NOT_1553(g2106,I5883);
  not NOT_1554(g8975,I15429);
  not NOT_1555(g3946,g3097);
  not NOT_1556(g2306,I6075);
  not NOT_1557(I13779,g7406);
  not NOT_1558(g9204,I15894);
  not NOT_1559(I15408,g8896);
  not NOT_1560(I15635,g8976);
  not NOT_1561(g6625,I11867);
  not NOT_1562(g1662,g1412);
  not NOT_1563(g2790,g1793);
  not NOT_1564(g7937,I14285);
  not NOT_1565(I7762,g3029);
  not NOT_1566(I12810,g6607);
  not NOT_1567(g6232,I11031);
  not NOT_1568(I11778,g6180);
  not NOT_1569(g3903,I7498);
  not NOT_1570(g9100,I15690);
  not NOT_1571(I12068,g5847);
  not NOT_1572(I10427,g5210);
  not NOT_1573(g7479,I13635);
  not NOT_1574(g9300,I16026);
  not NOT_1575(g5412,I9850);
  not NOT_1576(I10366,g5715);
  not NOT_1577(g6253,g5403);
  not NOT_1578(g6938,I12635);
  not NOT_1579(I14427,g7835);
  not NOT_1580(I5466,g926);
  not NOT_1581(g6813,I12310);
  not NOT_1582(g7294,I13314);
  not NOT_1583(g4373,I8360);
  not NOT_1584(g3513,g2407);
  not NOT_1585(I9139,g4364);
  not NOT_1586(g6909,I12592);
  not NOT_1587(g7190,I13112);
  not NOT_1588(g2622,g1568);
  not NOT_1589(I11945,g5874);
  not NOT_1590(I12337,g6724);
  not NOT_1591(I5365,g3843);
  not NOT_1592(I5861,g1313);
  not NOT_1593(I11356,g5799);
  not NOT_1594(I13356,g7221);
  not NOT_1595(g1816,g767);
  not NOT_1596(g5171,I9639);
  not NOT_1597(g4602,I8721);
  not NOT_1598(g7501,I13679);
  not NOT_1599(I11380,g5822);
  not NOT_1600(I10403,g5202);
  not NOT_1601(g5787,I10406);
  not NOT_1602(g4007,I7752);
  not NOT_1603(g2904,g2287);
  not NOT_1604(I14403,g7679);
  not NOT_1605(g7156,I13042);
  not NOT_1606(g5956,I10582);
  not NOT_1607(g6552,I11722);
  not NOT_1608(g7356,I13484);
  not NOT_1609(g4920,g4105);
  not NOT_1610(g6606,I11824);
  not NOT_1611(g4578,g2917);
  not NOT_1612(I11090,g1000);
  not NOT_1613(I7928,g2873);
  not NOT_1614(I11998,g5918);
  not NOT_1615(g8544,I14657);
  not NOT_1616(g3831,I7296);
  not NOT_1617(I11233,g6147);
  not NOT_1618(g2514,g1330);
  not NOT_1619(g4718,I9018);
  not NOT_1620(g8483,g8038);
  not NOT_1621(I8962,g4553);
  not NOT_1622(I7064,g2458);
  not NOT_1623(I11672,g5971);
  not NOT_1624(g1847,g765);
  not NOT_1625(I9672,g4803);
  not NOT_1626(I15711,g9075);
  not NOT_1627(I13672,g7242);
  not NOT_1628(I7899,g3743);
  not NOT_1629(g4535,g2876);
  not NOT_1630(g2403,g1176);
  not NOT_1631(g8636,I14718);
  not NOT_1632(g1685,I5528);
  not NOT_1633(g2145,g1296);
  not NOT_1634(g6687,I12003);
  not NOT_1635(g2345,I6151);
  not NOT_1636(g2841,g2208);
  not NOT_1637(I7785,g3029);
  not NOT_1638(g7704,I14001);
  not NOT_1639(g4582,g2922);
  not NOT_1640(g3805,g1752);
  not NOT_1641(g3916,I7545);
  not NOT_1642(g9323,g9315);
  not NOT_1643(g6586,I11778);
  not NOT_1644(g8790,g8585);
  not NOT_1645(g2695,g1672);
  not NOT_1646(g4015,g3160);
  not NOT_1647(g2637,g1581);
  not NOT_1648(I11449,g6068);
  not NOT_1649(I12918,g7013);
  not NOT_1650(g5684,I10183);
  not NOT_1651(g8061,I14330);
  not NOT_1652(g5745,I10292);
  not NOT_1653(I15492,g8971);
  not NOT_1654(g5639,g4748);
  not NOT_1655(I14127,g7594);
  not NOT_1656(g7163,I13063);
  not NOT_1657(g3947,I7640);
  not NOT_1658(I11897,g6141);
  not NOT_1659(g2307,I6078);
  not NOT_1660(I11961,g5988);
  not NOT_1661(g7032,g6525);
  not NOT_1662(g2536,g1354);
  not NOT_1663(g5109,I9493);
  not NOT_1664(I13897,g7354);
  not NOT_1665(g8756,g8564);
  not NOT_1666(g3798,g1757);
  not NOT_1667(g5309,g4969);
  not NOT_1668(g7432,I13559);
  not NOT_1669(g6141,I10786);
  not NOT_1670(g6860,I12451);
  not NOT_1671(g2359,g1397);
  not NOT_1672(g4664,I8907);
  not NOT_1673(I9499,g4382);
  not NOT_1674(g6341,I11350);
  not NOT_1675(I11404,g5834);
  not NOT_1676(g3560,g2361);
  not NOT_1677(g9351,I16103);
  not NOT_1678(g2223,I5942);
  not NOT_1679(I7844,g3784);
  not NOT_1680(I15982,g9236);
  not NOT_1681(g5808,I10457);
  not NOT_1682(g1562,g636);
  not NOT_1683(I6680,g1558);
  not NOT_1684(g6645,I11917);
  not NOT_1685(I16040,g9285);
  not NOT_1686(g4721,I9025);
  not NOT_1687(I14103,g7584);
  not NOT_1688(I11212,g6146);
  not NOT_1689(g2016,I5852);
  not NOT_1690(I7731,g3029);
  not NOT_1691(g5759,I10350);
  not NOT_1692(g8514,g8040);
  not NOT_1693(g3873,g2956);
  not NOT_1694(g3632,I7101);
  not NOT_1695(g3095,I6831);
  not NOT_1696(g1817,I5689);
  not NOT_1697(g3495,g1616);
  not NOT_1698(g3653,g2459);
  not NOT_1699(I8180,g3529);
  not NOT_1700(I12322,g6751);
  not NOT_1701(g8145,I14381);
  not NOT_1702(g2522,g1342);
  not NOT_1703(I14181,g7725);
  not NOT_1704(g7157,I13045);
  not NOT_1705(g2642,g1588);
  not NOT_1706(I8832,g3936);
  not NOT_1707(g6879,I12508);
  not NOT_1708(g7357,I13487);
  not NOT_1709(g6607,I11827);
  not NOT_1710(I12532,g6594);
  not NOT_1711(g3579,g1929);
  not NOT_1712(g3869,I7400);
  not NOT_1713(g6962,I12687);
  not NOT_1714(I8853,g4034);
  not NOT_1715(g6659,I11955);
  not NOT_1716(I12158,g5956);
  not NOT_1717(g6358,I11401);
  not NOT_1718(g6506,I11680);
  not NOT_1719(g1751,g452);
  not NOT_1720(I5847,g1360);
  not NOT_1721(I12561,g6449);
  not NOT_1722(I16183,g9388);
  not NOT_1723(g5604,g4969);
  not NOT_1724(I12295,g6693);
  not NOT_1725(g3917,I7548);
  not NOT_1726(g2654,I6446);
  not NOT_1727(I10190,g4670);
  not NOT_1728(g1585,g724);
  not NOT_1729(g4689,I8966);
  not NOT_1730(g6587,I11781);
  not NOT_1731(g9372,I16142);
  not NOT_1732(I15522,g9018);
  not NOT_1733(I15663,g9066);
  not NOT_1734(I14190,g7531);
  not NOT_1735(I9543,g4279);
  not NOT_1736(g6111,g5453);
  not NOT_1737(g8223,I14448);
  not NOT_1738(g6311,I11260);
  not NOT_1739(g5833,I10522);
  not NOT_1740(I7814,g2605);
  not NOT_1741(I13646,g7245);
  not NOT_1742(g9235,I15959);
  not NOT_1743(g4028,I7797);
  not NOT_1744(g2880,g2234);
  not NOT_1745(I7350,g2971);
  not NOT_1746(I6574,g576);
  not NOT_1747(g2595,g1643);
  not NOT_1748(I6864,g2528);
  not NOT_1749(I11971,g6179);
  not NOT_1750(g4030,g3160);
  not NOT_1751(g8016,I14311);
  not NOT_1752(g8757,g8585);
  not NOT_1753(g5584,g4841);
  not NOT_1754(g1673,g1504);
  not NOT_1755(g6374,I11449);
  not NOT_1756(I14211,g7712);
  not NOT_1757(g9134,I15776);
  not NOT_1758(I15553,g9009);
  not NOT_1759(I13369,g7268);
  not NOT_1760(g2272,I6021);
  not NOT_1761(I14088,g7585);
  not NOT_1762(g4564,I8665);
  not NOT_1763(I11368,g5833);
  not NOT_1764(g8642,I14732);
  not NOT_1765(I5562,g1300);
  not NOT_1766(I12364,g6714);
  not NOT_1767(I7769,g3038);
  not NOT_1768(g5162,I9612);
  not NOT_1769(g3770,g2551);
  not NOT_1770(g5268,I9788);
  not NOT_1771(I9014,g3864);
  not NOT_1772(g5362,I9823);
  not NOT_1773(I10497,g5233);
  not NOT_1774(I15536,g9004);
  not NOT_1775(g1772,g607);
  not NOT_1776(g6380,I11467);
  not NOT_1777(I9660,g4806);
  not NOT_1778(g6591,I11787);
  not NOT_1779(I15702,g9064);
  not NOT_1780(I13850,g7328);
  not NOT_1781(g6832,I12367);
  not NOT_1782(I5817,g1081);
  not NOT_1783(g2982,g1848);
  not NOT_1784(g8874,I15208);
  not NOT_1785(g3532,g2407);
  not NOT_1786(I7967,g2787);
  not NOT_1787(g7778,I14205);
  not NOT_1788(g1743,g598);
  not NOT_1789(g2234,I5963);
  not NOT_1790(g6853,I12430);
  not NOT_1791(g2128,g1284);
  not NOT_1792(g4638,I8829);
  not NOT_1793(g2629,g1574);
  not NOT_1794(g6020,g5367);
  not NOT_1795(g2328,I6127);
  not NOT_1796(I10987,g5609);
  not NOT_1797(I12289,g6702);
  not NOT_1798(I5605,g58);
  not NOT_1799(I10250,g5268);
  not NOT_1800(g7735,I14076);
  not NOT_1801(g4609,I8742);
  not NOT_1802(g6507,I11683);
  not NOT_1803(g4308,I8277);
  not NOT_1804(g1011,I5413);
  not NOT_1805(I13228,g6892);
  not NOT_1806(g9113,I15729);
  not NOT_1807(g6794,I12253);
  not NOT_1808(g1856,g774);
  not NOT_1809(I12571,g6729);
  not NOT_1810(g9313,I16055);
  not NOT_1811(I11011,g5693);
  not NOT_1812(I5751,g963);
  not NOT_1813(g5086,I9460);
  not NOT_1814(g8880,I15218);
  not NOT_1815(g3189,I6864);
  not NOT_1816(I13716,g7331);
  not NOT_1817(g5730,I10247);
  not NOT_1818(g7475,I13631);
  not NOT_1819(I16072,g9303);
  not NOT_1820(g3990,g3160);
  not NOT_1821(g2554,I6376);
  not NOT_1822(I14338,g7581);
  not NOT_1823(g5185,I9681);
  not NOT_1824(g4589,g2930);
  not NOT_1825(I10969,g5606);
  not NOT_1826(g9094,I15672);
  not NOT_1827(g7627,I13956);
  not NOT_1828(g3888,g3097);
  not NOT_1829(I15062,g8632);
  not NOT_1830(g6905,I12586);
  not NOT_1831(g3029,g1929);
  not NOT_1832(g7292,I13308);
  not NOT_1833(g3787,g1842);
  not NOT_1834(g8017,g7692);
  not NOT_1835(g6628,I11880);
  not NOT_1836(I15933,g9210);
  not NOT_1837(g7526,I13758);
  not NOT_1838(g5470,g4899);
  not NOT_1839(g5897,I10569);
  not NOT_1840(g3956,g2845);
  not NOT_1841(g5025,I9363);
  not NOT_1842(g6515,g6125);
  not NOT_1843(I11627,g5874);
  not NOT_1844(g6630,I11884);
  not NOT_1845(g4571,g2908);
  not NOT_1846(I12687,g6745);
  not NOT_1847(g3675,I7167);
  not NOT_1848(I12976,g6928);
  not NOT_1849(g1573,g677);
  not NOT_1850(g1863,g68);
  not NOT_1851(g6300,I11227);
  not NOT_1852(I13112,g7021);
  not NOT_1853(g7603,I13940);
  not NOT_1854(I11050,g5335);
  not NOT_1855(I11958,g5874);
  not NOT_1856(g7039,g6543);
  not NOT_1857(I9422,g4360);
  not NOT_1858(I8351,g1160);
  not NOT_1859(g8234,I14489);
  not NOT_1860(g4455,g3811);
  not NOT_1861(g2902,g2285);
  not NOT_1862(g7439,I13574);
  not NOT_1863(I12643,g6501);
  not NOT_1864(I5368,g3853);
  not NOT_1865(I11386,g5764);
  not NOT_1866(g1569,g661);
  not NOT_1867(g453,I5362);
  not NOT_1868(I5772,g1240);
  not NOT_1869(g2490,I6326);
  not NOT_1870(I6024,g544);
  not NOT_1871(I5531,g866);
  not NOT_1872(g2366,I6198);
  not NOT_1873(I12669,g6477);
  not NOT_1874(g7583,I13894);
  not NOT_1875(g7702,I13997);
  not NOT_1876(g4196,I8097);
  not NOT_1877(g5678,I10169);
  not NOT_1878(I6795,g1683);
  not NOT_1879(I10503,g5235);
  not NOT_1880(g3684,g2180);
  not NOT_1881(g3639,g2424);
  not NOT_1882(g4803,I9132);
  not NOT_1883(g6973,I12708);
  not NOT_1884(g5006,I9333);
  not NOT_1885(g3338,g1901);
  not NOT_1886(g8800,I15010);
  not NOT_1887(g3963,I7672);
  not NOT_1888(g9360,I16116);
  not NOT_1889(I15574,g8983);
  not NOT_1890(g4538,g2880);
  not NOT_1891(g1688,I5535);
  not NOT_1892(g2148,g1304);
  not NOT_1893(I15205,g8809);
  not NOT_1894(g2649,I6431);
  not NOT_1895(g4780,I9089);
  not NOT_1896(g1857,g889);
  not NOT_1897(g2348,I6160);
  not NOT_1898(I7788,g2595);
  not NOT_1899(g9050,I15550);
  not NOT_1900(g5682,I10177);
  not NOT_1901(g5766,I10373);
  not NOT_1902(g5087,I9463);
  not NOT_1903(g1976,g1269);
  not NOT_1904(g6969,I12702);
  not NOT_1905(I15912,g9193);
  not NOT_1906(I9095,g4283);
  not NOT_1907(g5801,I10442);
  not NOT_1908(g3808,g1827);
  not NOT_1909(g7276,I13264);
  not NOT_1910(g5487,I9907);
  not NOT_1911(I14315,g7676);
  not NOT_1912(I6643,g1970);
  not NOT_1913(I11793,g6188);
  not NOT_1914(I11428,g5813);
  not NOT_1915(I12424,g6446);
  not NOT_1916(I13428,g7167);
  not NOT_1917(g3707,g2226);
  not NOT_1918(g6323,I11296);
  not NOT_1919(I14819,g8647);
  not NOT_1920(g4662,I8901);
  not NOT_1921(g2698,g1673);
  not NOT_1922(g4018,I7775);
  not NOT_1923(I12558,g6449);
  not NOT_1924(I14202,g7708);
  not NOT_1925(I8172,g3524);
  not NOT_1926(I14257,g7716);
  not NOT_1927(I9579,g4713);
  not NOT_1928(g2964,I6716);
  not NOT_1929(I14055,g7495);
  not NOT_1930(I16020,g9264);
  not NOT_1931(g9379,I16161);
  not NOT_1932(I7392,g3230);
  not NOT_1933(g5755,g5494);
  not NOT_1934(I15592,g8989);
  not NOT_1935(I15756,g9081);
  not NOT_1936(g7527,I13761);
  not NOT_1937(I14070,g7714);
  not NOT_1938(g3957,I7662);
  not NOT_1939(I12544,g6617);
  not NOT_1940(I6099,g584);
  not NOT_1941(I9752,g4705);
  not NOT_1942(g4093,I7902);
  not NOT_1943(g8512,g8094);
  not NOT_1944(I8282,g3515);
  not NOT_1945(I16046,g9288);
  not NOT_1946(g1760,I5605);
  not NOT_1947(g4493,I8543);
  not NOT_1948(g7764,I14163);
  not NOT_1949(g6351,I11380);
  not NOT_1950(g6648,I11926);
  not NOT_1951(g6875,I12496);
  not NOT_1952(g7546,I13822);
  not NOT_1953(g3865,g2944);
  not NOT_1954(I10384,g5193);
  not NOT_1955(g6655,I11945);
  not NOT_1956(g5445,g5059);
  not NOT_1957(g5173,I9645);
  not NOT_1958(I11317,g5787);
  not NOT_1959(g3604,g2407);
  not NOT_1960(I13317,g7211);
  not NOT_1961(g5491,g4918);
  not NOT_1962(g3498,g1616);
  not NOT_1963(I14067,g7550);
  not NOT_1964(I14094,g7593);
  not NOT_1965(g4381,g3466);
  not NOT_1966(g8649,I14743);
  not NOT_1967(g6010,I10608);
  not NOT_1968(g3833,I7302);
  not NOT_1969(I11129,g5418);
  not NOT_1970(g2872,I6590);
  not NOT_1971(g1924,g174);
  not NOT_1972(g5169,I9633);
  not NOT_1973(g4685,I8952);
  not NOT_1974(g4197,g3591);
  not NOT_1975(I10801,g5463);
  not NOT_1976(g6410,I11533);
  not NOT_1977(g7224,I13164);
  not NOT_1978(I7520,g2734);
  not NOT_1979(g4021,g3131);
  not NOT_1980(g5007,I9336);
  not NOT_1981(I13057,g6968);
  not NOT_1982(I14801,g8608);
  not NOT_1983(g2652,I6440);
  not NOT_1984(g1779,g612);
  not NOT_1985(g2057,I5868);
  not NOT_1986(I7640,g3062);
  not NOT_1987(I12124,g5847);
  not NOT_1988(I12678,g6516);
  not NOT_1989(g6884,I12523);
  not NOT_1990(g2843,I6571);
  not NOT_1991(g7120,I12948);
  not NOT_1992(g5059,I9419);
  not NOT_1993(g6839,I12388);
  not NOT_1994(g2457,g24);
  not NOT_1995(g5578,g4841);
  not NOT_1996(g5868,I10555);
  not NOT_1997(g7320,I13388);
  not NOT_1998(g2989,g1843);
  not NOT_1999(g3539,g2424);
  not NOT_2000(g3896,I7473);
  not NOT_2001(I11245,g6143);
  not NOT_2002(g5459,g4882);
  not NOT_2003(I14019,g7480);
  not NOT_2004(g2393,I6267);
  not NOT_2005(g5718,g4841);
  not NOT_2006(I12460,g6674);
  not NOT_2007(I12939,g7022);
  not NOT_2008(I11323,g5808);
  not NOT_2009(g1977,g1357);
  not NOT_2010(I11299,g5786);
  not NOT_2011(I13323,g7145);
  not NOT_2012(I14196,g7534);
  not NOT_2013(I13299,g7163);
  not NOT_2014(I14695,g8016);
  not NOT_2015(g7277,I13267);
  not NOT_2016(g1588,g741);
  not NOT_2017(I11533,g5847);
  not NOT_2018(g2834,I6564);
  not NOT_2019(g2971,I6723);
  not NOT_2020(I13533,g7220);
  not NOT_2021(g8063,I14334);
  not NOT_2022(g5582,g4969);
  not NOT_2023(I15405,g8902);
  not NOT_2024(g6278,I11129);
  not NOT_2025(g8463,g8094);
  not NOT_2026(g2686,g1667);
  not NOT_2027(g6372,I11443);
  not NOT_2028(g7789,I14224);
  not NOT_2029(g5261,g4748);
  not NOT_2030(g3019,g2007);
  not NOT_2031(g9132,I15770);
  not NOT_2032(g5793,I10418);
  not NOT_2033(I12065,g5897);
  not NOT_2034(I8202,g3560);
  not NOT_2035(g9332,g9322);
  not NOT_2036(g6618,g6003);
  not NOT_2037(g1665,g1467);
  not NOT_2038(g6143,I10796);
  not NOT_2039(g7516,I13728);
  not NOT_2040(I7765,g2595);
  not NOT_2041(g6343,I11356);
  not NOT_2042(g4562,g3466);
  not NOT_2043(g6235,I11034);
  not NOT_2044(g5015,I9347);
  not NOT_2045(g3052,g2096);
  not NOT_2046(g9209,g9199);
  not NOT_2047(g9353,I16107);
  not NOT_2048(I7911,g2767);
  not NOT_2049(I10457,g5218);
  not NOT_2050(I8094,g2976);
  not NOT_2051(g7771,I14184);
  not NOT_2052(I14457,g8093);
  not NOT_2053(g6566,I11740);
  not NOT_2054(g4631,I8808);
  not NOT_2055(I13737,g7446);
  not NOT_2056(g372,I5359);
  not NOT_2057(I15583,g8986);
  not NOT_2058(g7299,I13329);
  not NOT_2059(g4257,I8190);
  not NOT_2060(g6693,I12011);
  not NOT_2061(g6134,g5428);
  not NOT_2062(g8619,I14695);
  not NOT_2063(g7547,I13825);
  not NOT_2064(g6334,I11329);
  not NOT_2065(g4301,I8264);
  not NOT_2066(g5246,I9760);
  not NOT_2067(g2625,g1570);
  not NOT_2068(g8872,I15202);
  not NOT_2069(g2232,I5957);
  not NOT_2070(g4605,I8730);
  not NOT_2071(g3086,g1852);
  not NOT_2072(g2253,g1323);
  not NOT_2073(g2938,g2347);
  not NOT_2074(g3728,g2202);
  not NOT_2075(I14001,g7433);
  not NOT_2076(I13261,g7041);
  not NOT_2077(I11880,g5748);
  not NOT_2078(g6555,I11729);
  not NOT_2079(g6804,I12283);
  not NOT_2080(I7473,g3546);
  not NOT_2081(g2909,g2291);
  not NOT_2082(I6946,g1887);
  not NOT_2083(I10256,g5401);
  not NOT_2084(g6792,I12247);
  not NOT_2085(I11512,g5874);
  not NOT_2086(g1732,g1439);
  not NOT_2087(I9675,g4807);
  not NOT_2088(I13512,g7138);
  not NOT_2089(g3881,g2969);
  not NOT_2090(I5383,g647);
  not NOT_2091(I10280,g5488);
  not NOT_2092(g8971,I15417);
  not NOT_2093(g7738,I14085);
  not NOT_2094(g4585,g2925);
  not NOT_2095(I8264,g3653);
  not NOT_2096(g6621,I11855);
  not NOT_2097(g1944,I5817);
  not NOT_2098(g3897,g3131);
  not NOT_2099(g4041,g2605);
  not NOT_2100(I12915,g7000);
  not NOT_2101(g9092,I15666);
  not NOT_2102(I8360,g1186);
  not NOT_2103(g6313,I11266);
  not NOT_2104(g7078,g6683);
  not NOT_2105(g7340,I13438);
  not NOT_2106(I7377,g3189);
  not NOT_2107(I10157,g5109);
  not NOT_2108(I13831,g7322);
  not NOT_2109(I6036,g130);
  not NOT_2110(I14157,g7547);
  not NOT_2111(I12277,g6681);
  not NOT_2112(I6178,g1220);
  not NOT_2113(g4673,I8928);
  not NOT_2114(g6202,I10949);
  not NOT_2115(g8670,I14804);
  not NOT_2116(I9684,g4813);
  not NOT_2117(g7035,g6543);
  not NOT_2118(I13499,g7134);
  not NOT_2119(I15803,g9148);
  not NOT_2120(I9639,g4685);
  not NOT_2121(g7517,I13731);
  not NOT_2122(I7287,g2561);
  not NOT_2123(g6094,I10716);
  not NOT_2124(I14231,g7566);
  not NOT_2125(I9791,g4779);
  not NOT_2126(I6831,g2185);
  not NOT_2127(g5028,I9372);
  not NOT_2128(g4669,I8922);
  not NOT_2129(g1565,g649);
  not NOT_2130(I8724,g3927);
  not NOT_2131(g5671,I10160);
  not NOT_2132(I11722,g5772);
  not NOT_2133(I12782,g6463);
  not NOT_2134(I13722,g7442);
  not NOT_2135(I16090,g9336);
  not NOT_2136(I6805,g1603);
  not NOT_2137(g3635,g1949);
  not NOT_2138(I13924,g7365);
  not NOT_2139(I5633,g891);
  not NOT_2140(g1681,g929);
  not NOT_2141(g6776,I12199);
  not NOT_2142(I7781,g2605);
  not NOT_2143(I6422,g1805);
  not NOT_2144(g6593,I11793);
  not NOT_2145(g4890,g4075);
  not NOT_2146(I12352,g6752);
  not NOT_2147(I13432,g7280);
  not NOT_2148(g2525,I6354);
  not NOT_2149(g3801,I7262);
  not NOT_2150(I14763,g7834);
  not NOT_2151(I13271,g7067);
  not NOT_2152(g2645,I6419);
  not NOT_2153(I8835,g3954);
  not NOT_2154(g5826,I10503);
  not NOT_2155(I12418,g6572);
  not NOT_2156(I7797,g3019);
  not NOT_2157(g8606,I14683);
  not NOT_2158(I12170,g5956);
  not NOT_2159(g4011,I7762);
  not NOT_2160(I11461,g6094);
  not NOT_2161(g9076,I15622);
  not NOT_2162(g5741,I10280);
  not NOT_2163(g7110,I12918);
  not NOT_2164(I5732,g859);
  not NOT_2165(g6264,g5403);
  not NOT_2166(g7310,I13362);
  not NOT_2167(I11031,g5335);
  not NOT_2168(I13031,g6984);
  not NOT_2169(g5638,g4748);
  not NOT_2170(g6360,I11407);
  not NOT_2171(g2879,I6597);
  not NOT_2172(I13199,g7025);
  not NOT_2173(I11736,g6076);
  not NOT_2174(I11887,g5918);
  not NOT_2175(g9375,I16151);
  not NOT_2176(I7344,g2964);
  not NOT_2177(g2962,g2382);
  not NOT_2178(g5609,g4748);
  not NOT_2179(I15003,g8633);
  not NOT_2180(I8799,g3951);
  not NOT_2181(g2659,g1655);
  not NOT_2182(g6050,g5246);
  not NOT_2183(I12167,g5939);
  not NOT_2184(g2506,I6341);
  not NOT_2185(g1820,g621);
  not NOT_2186(I6437,g1784);
  not NOT_2187(I11696,g5971);
  not NOT_2188(g7236,g6944);
  not NOT_2189(I6302,g1313);
  not NOT_2190(g3091,g1603);
  not NOT_2191(I13843,g7326);
  not NOT_2192(I16026,g9267);
  not NOT_2193(g7762,I14157);
  not NOT_2194(g3491,g1800);
  not NOT_2195(g4080,I7867);
  not NOT_2196(I14076,g7577);
  not NOT_2197(I14085,g7583);
  not NOT_2198(g4573,g2911);
  not NOT_2199(I11764,g6056);
  not NOT_2200(g5758,I10347);
  not NOT_2201(I13764,g7479);
  not NOT_2202(g6724,I12088);
  not NOT_2203(I11365,g5826);
  not NOT_2204(g2275,g990);
  not NOT_2205(g2311,I6090);
  not NOT_2206(I9539,g4018);
  not NOT_2207(g6179,I10896);
  not NOT_2208(I13365,g7267);
  not NOT_2209(g5466,g4890);
  not NOT_2210(g4713,I9014);
  not NOT_2211(I10243,g5026);
  not NOT_2212(g6379,I11464);
  not NOT_2213(I11132,g5624);
  not NOT_2214(g7590,I13915);
  not NOT_2215(g9184,I15830);
  not NOT_2216(I13869,g7338);
  not NOT_2217(I5565,g1296);
  not NOT_2218(g2615,g1563);
  not NOT_2219(g6878,I12505);
  not NOT_2220(g5165,I9621);
  not NOT_2221(g4569,g2906);
  not NOT_2222(g5571,I10032);
  not NOT_2223(g3920,g3097);
  not NOT_2224(I12022,g5874);
  not NOT_2225(g3578,I7053);
  not NOT_2226(g3868,g2948);
  not NOT_2227(g2174,g1319);
  not NOT_2228(g6289,I11194);
  not NOT_2229(g6777,I12202);
  not NOT_2230(I8802,g3963);
  not NOT_2231(g6658,g6224);
  not NOT_2232(g2374,I6220);
  not NOT_2233(g5448,g5137);
  not NOT_2234(g1922,g1251);
  not NOT_2235(I9162,g4272);
  not NOT_2236(g7556,I13846);
  not NOT_2237(I13161,g7080);
  not NOT_2238(I10773,g5708);
  not NOT_2239(g5055,g4477);
  not NOT_2240(I12313,g6730);
  not NOT_2241(g6835,I12376);
  not NOT_2242(g2985,I6733);
  not NOT_2243(I9419,g3916);
  not NOT_2244(I10268,g5471);
  not NOT_2245(g1581,g710);
  not NOT_2246(g5827,I10506);
  not NOT_2247(I12748,g6585);
  not NOT_2248(g6882,I12517);
  not NOT_2249(I6042,g237);
  not NOT_2250(I15651,g9056);
  not NOT_2251(I15672,g9047);
  not NOT_2252(g3582,g2407);
  not NOT_2253(g2284,I6036);
  not NOT_2254(I5914,g1097);
  not NOT_2255(I13225,g7095);
  not NOT_2256(g7064,I12829);
  not NOT_2257(g2239,I5978);
  not NOT_2258(I7314,g2916);
  not NOT_2259(I10180,g4721);
  not NOT_2260(I16148,g9368);
  not NOT_2261(g1597,g973);
  not NOT_2262(g9077,I15625);
  not NOT_2263(g2180,g1318);
  not NOT_2264(g5846,g5367);
  not NOT_2265(g2380,I6242);
  not NOT_2266(I13258,g6907);
  not NOT_2267(I12900,g6947);
  not NOT_2268(I7870,g2827);
  not NOT_2269(I8901,g4122);
  not NOT_2270(g2832,g2184);
  not NOT_2271(I12466,g6687);
  not NOT_2272(g5396,g4692);
  not NOT_2273(I5413,g1016);
  not NOT_2274(g1784,I5636);
  not NOT_2275(g6799,I12268);
  not NOT_2276(I6054,g465);
  not NOT_2277(g2020,I5855);
  not NOT_2278(I10930,g5600);
  not NOT_2279(I15513,g8970);
  not NOT_2280(I11043,g5648);
  not NOT_2281(I6454,g1868);
  not NOT_2282(I12101,g5971);
  not NOT_2283(I6770,g1590);
  not NOT_2284(g6674,I11978);
  not NOT_2285(I13244,g7033);
  not NOT_2286(g7563,I13861);
  not NOT_2287(g8111,I14374);
  not NOT_2288(g5780,I10387);
  not NOT_2289(g4000,g3131);
  not NOT_2290(I10694,g5445);
  not NOT_2291(g4126,I7981);
  not NOT_2292(I10965,g5719);
  not NOT_2293(g6997,I12737);
  not NOT_2294(g7295,I13317);
  not NOT_2295(g2794,g2185);
  not NOT_2296(I11069,g5671);
  not NOT_2297(g9104,I15702);
  not NOT_2298(I5936,g222);
  not NOT_2299(g9099,I15687);
  not NOT_2300(I6532,g1694);
  not NOT_2301(g9304,g9298);
  not NOT_2302(g2931,I6669);
  not NOT_2303(g3721,I7211);
  not NOT_2304(g6238,I11043);
  not NOT_2305(I6553,g2246);
  not NOT_2306(g5662,g5027);
  not NOT_2307(I13810,g7312);
  not NOT_2308(g8174,I14403);
  not NOT_2309(g6332,I11323);
  not NOT_2310(I15717,g9051);
  not NOT_2311(I11955,g5988);
  not NOT_2312(g5418,g5100);
  not NOT_2313(g5467,g4891);
  not NOT_2314(I9025,g4462);
  not NOT_2315(g6353,I11386);
  not NOT_2316(g7194,I13118);
  not NOT_2317(I13879,g7332);
  not NOT_2318(I9425,g3917);
  not NOT_2319(g655,I5383);
  not NOT_2320(g2905,I6629);
  not NOT_2321(I6012,g384);
  not NOT_2322(g6744,I12124);
  not NOT_2323(g7731,I14064);
  not NOT_2324(g6802,I12277);
  not NOT_2325(g8284,I14531);
  not NOT_2326(g2628,g1573);
  not NOT_2327(g3502,g1616);
  not NOT_2328(g8545,g7905);
  not NOT_2329(I6189,g249);
  not NOT_2330(g2630,g1575);
  not NOT_2331(g5493,g4920);
  not NOT_2332(g8180,g7719);
  not NOT_2333(I14279,g7700);
  not NOT_2334(g4608,I8739);
  not NOT_2335(g4924,g4113);
  not NOT_2336(I5775,g1240);
  not NOT_2337(g7966,I14291);
  not NOT_2338(g2100,g1227);
  not NOT_2339(g3940,I7623);
  not NOT_2340(I10469,g5222);
  not NOT_2341(I11967,g5971);
  not NOT_2342(I11994,g6195);
  not NOT_2343(g7471,g7233);
  not NOT_2344(I15723,g9065);
  not NOT_2345(g9044,I15536);
  not NOT_2346(g1942,g828);
  not NOT_2347(I6029,g1207);
  not NOT_2348(g4023,I7788);
  not NOT_2349(I8736,g4008);
  not NOT_2350(I10286,g5519);
  not NOT_2351(I6371,g33);
  not NOT_2352(g1704,I5548);
  not NOT_2353(g5181,I9669);
  not NOT_2354(I12008,g5897);
  not NOT_2355(I9678,g4808);
  not NOT_2356(I15433,g8911);
  not NOT_2357(g5847,I10552);
  not NOT_2358(I6956,g1907);
  not NOT_2359(g6901,g6525);
  not NOT_2360(I14039,g7449);
  not NOT_2361(g4588,g2929);
  not NOT_2362(I11425,g5872);
  not NOT_2363(g5685,I10186);
  not NOT_2364(g5197,g4938);
  not NOT_2365(I13425,g7166);
  not NOT_2366(g5397,g5076);
  not NOT_2367(I8889,g4311);
  not NOT_2368(g6511,I11693);
  not NOT_2369(g703,I5398);
  not NOT_2370(I11458,g6063);
  not NOT_2371(I15811,g9151);
  not NOT_2372(I10815,g5418);
  not NOT_2373(I12454,g6581);
  not NOT_2374(g2973,g1854);
  not NOT_2375(g1810,I5676);
  not NOT_2376(g3430,I6956);
  not NOT_2377(g4665,I8910);
  not NOT_2378(I12712,g6543);
  not NOT_2379(g4051,g3093);
  not NOT_2380(g6092,g5317);
  not NOT_2381(I13918,g7361);
  not NOT_2382(I15971,g9233);
  not NOT_2383(I8871,g3869);
  not NOT_2384(I14187,g7728);
  not NOT_2385(g7150,g6952);
  not NOT_2386(I14677,g7791);
  not NOT_2387(g7350,I13466);
  not NOT_2388(g6864,I12463);
  not NOT_2389(I7195,g1795);
  not NOT_2390(g2969,g2393);
  not NOT_2391(I13444,g7282);
  not NOT_2392(g6714,I12068);
  not NOT_2393(g7773,I14190);
  not NOT_2394(g4146,I8011);
  not NOT_2395(g7009,I12753);
  not NOT_2396(g4633,I8814);
  not NOT_2397(g2323,I6112);
  not NOT_2398(I10937,g5560);
  not NOT_2399(I6963,g1558);
  not NOT_2400(g1568,g658);
  not NOT_2401(I6109,g1214);
  not NOT_2402(I6791,g1967);
  not NOT_2403(g4103,I7922);
  not NOT_2404(I12567,g6721);
  not NOT_2405(I6309,g1336);
  not NOT_2406(g4303,I8268);
  not NOT_2407(I11086,g5397);
  not NOT_2408(I7807,g2595);
  not NOT_2409(g3910,I7523);
  not NOT_2410(I12238,g6637);
  not NOT_2411(g7769,I14178);
  not NOT_2412(I10169,g4873);
  not NOT_2413(I7859,g2804);
  not NOT_2414(g4696,I8983);
  not NOT_2415(g1912,g1524);
  not NOT_2416(g5631,g4938);
  not NOT_2417(g7836,I14260);
  not NOT_2418(I14169,g7715);
  not NOT_2419(g5723,g4938);
  not NOT_2420(g4732,I9034);
  not NOT_2421(g5101,g4259);
  not NOT_2422(I12382,g6772);
  not NOT_2423(I5356,g3837);
  not NOT_2424(g2528,g1260);
  not NOT_2425(I14410,g7697);
  not NOT_2426(g2351,g792);
  not NOT_2427(g2648,I6428);
  not NOT_2428(I8838,g3967);
  not NOT_2429(I12176,g5939);
  not NOT_2430(I8024,g3076);
  not NOT_2431(I12675,g6510);
  not NOT_2432(g6736,I12108);
  not NOT_2433(g8750,g8524);
  not NOT_2434(I10479,g5227);
  not NOT_2435(g6968,I12699);
  not NOT_2436(g2655,g1611);
  not NOT_2437(g8973,I15423);
  not NOT_2438(g1929,g1224);
  not NOT_2439(I12154,g5874);
  not NOT_2440(I5942,g300);
  not NOT_2441(I9369,g3901);
  not NOT_2442(g7229,g6938);
  not NOT_2443(g6623,I11861);
  not NOT_2444(g7993,I14298);
  not NOT_2445(I7255,g1955);
  not NOT_2446(g6076,g5287);
  not NOT_2447(I14015,g7440);
  not NOT_2448(I9407,g4232);
  not NOT_2449(g6889,I12538);
  not NOT_2450(I11656,g5772);
  not NOT_2451(I13656,g7228);
  not NOT_2452(g3589,I7061);
  not NOT_2453(g8040,g7699);
  not NOT_2454(I11353,g5788);
  not NOT_2455(g9036,I15522);
  not NOT_2456(g4443,I8449);
  not NOT_2457(I13353,g7231);
  not NOT_2458(I11680,g5939);
  not NOT_2459(g8969,I15411);
  not NOT_2460(I8477,g3014);
  not NOT_2461(g9178,I15814);
  not NOT_2462(g9378,I16158);
  not NOT_2463(I13144,g7031);
  not NOT_2464(g4116,I7959);
  not NOT_2465(g6375,I11452);
  not NOT_2466(g6871,I12484);
  not NOT_2467(g4316,I8291);
  not NOT_2468(I5954,g89);
  not NOT_2469(g2884,g2238);
  not NOT_2470(g3861,I7386);
  not NOT_2471(g5041,I9393);
  not NOT_2472(g3048,I6784);
  not NOT_2473(g4034,I7811);
  not NOT_2474(I9582,g4694);
  not NOT_2475(I8205,g2655);
  not NOT_2476(g6651,I11933);
  not NOT_2477(g9182,g9178);
  not NOT_2478(I5432,g1176);
  not NOT_2479(g4565,g2901);
  not NOT_2480(g8666,I14792);
  not NOT_2481(g9382,I16168);
  not NOT_2482(I15959,g9217);
  not NOT_2483(I15379,g8882);
  not NOT_2484(I8742,g3919);
  not NOT_2485(g2372,I6214);
  not NOT_2486(g3774,g1770);
  not NOT_2487(I13631,g7248);
  not NOT_2488(I5568,g1409);
  not NOT_2489(g8875,I15211);
  not NOT_2490(g3846,I7341);
  not NOT_2491(g2618,g1566);
  not NOT_2492(g1683,g795);
  not NOT_2493(I16129,g9355);
  not NOT_2494(g6384,I11479);
  not NOT_2495(g2235,I5966);
  not NOT_2496(g2343,g1392);
  not NOT_2497(g6139,I10780);
  not NOT_2498(g5168,I9630);
  not NOT_2499(I12439,g6566);
  not NOT_2500(g5669,I10154);
  not NOT_2501(g4697,I8986);
  not NOT_2502(g6339,I11344);
  not NOT_2503(g4914,g4093);
  not NOT_2504(I14531,g8178);
  not NOT_2505(g2282,g1400);
  not NOT_2506(I7112,g2546);
  not NOT_2507(g1778,g613);
  not NOT_2508(g1894,I5772);
  not NOT_2509(g5058,I9416);
  not NOT_2510(g6838,I12385);
  not NOT_2511(g4596,g3466);
  not NOT_2512(I8754,g3911);
  not NOT_2513(g6024,g5494);
  not NOT_2514(I14178,g7562);
  not NOT_2515(g4013,g3131);
  not NOT_2516(g2134,g1317);
  not NOT_2517(g6795,I12256);
  not NOT_2518(g3780,g1847);
  not NOT_2519(I10186,g5129);
  not NOT_2520(g6737,I12111);
  not NOT_2521(g2334,I6143);
  not NOT_2522(I15681,g9063);
  not NOT_2523(g6809,I12298);
  not NOT_2524(I8273,g2976);
  not NOT_2525(I12349,g6742);
  not NOT_2526(g5743,I10286);
  not NOT_2527(I6419,g1799);
  not NOT_2528(I10373,g5722);
  not NOT_2529(g1782,g624);
  not NOT_2530(I7676,g2584);
  not NOT_2531(g2548,g1351);
  not NOT_2532(I7293,g2955);
  not NOT_2533(I12906,g6918);
  not NOT_2534(I15429,g8899);
  not NOT_2535(I7129,g2495);
  not NOT_2536(I13023,g7040);
  not NOT_2537(g1661,g1405);
  not NOT_2538(I7329,g2920);
  not NOT_2539(I11224,g6255);
  not NOT_2540(g6672,I11974);
  not NOT_2541(g2555,g936);
  not NOT_2542(g6231,I11028);
  not NOT_2543(g3018,I6770);
  not NOT_2544(I11308,g5759);
  not NOT_2545(g2804,g1796);
  not NOT_2546(I12304,g6711);
  not NOT_2547(g9095,I15675);
  not NOT_2548(I13308,g7169);
  not NOT_2549(g5734,I10259);
  not NOT_2550(g1949,g1292);
  not NOT_2551(g6523,I11707);
  not NOT_2552(I9502,g3972);
  not NOT_2553(g3994,g3192);
  not NOT_2554(I8983,g4536);
  not NOT_2555(g9102,I15696);
  not NOT_2556(g9208,g9198);
  not NOT_2557(I15765,g9039);
  not NOT_2558(g9302,g9281);
  not NOT_2559(I8862,g3981);
  not NOT_2560(g6205,g5628);
  not NOT_2561(I14334,g7578);
  not NOT_2562(g8172,I14397);
  not NOT_2563(I15690,g9074);
  not NOT_2564(g2621,g1567);
  not NOT_2565(I8712,g4007);
  not NOT_2566(I7592,g2712);
  not NOT_2567(g5074,I9440);
  not NOT_2568(g3093,g1686);
  not NOT_2569(I6728,g1959);
  not NOT_2570(I8543,g2810);
  not NOT_2571(g5474,g4904);
  not NOT_2572(g1646,g1214);
  not NOT_2573(g7298,I13326);
  not NOT_2574(g4601,I8718);
  not NOT_2575(I7746,g3591);
  not NOT_2576(g6634,I11894);
  not NOT_2577(g8667,I14795);
  not NOT_2578(I13816,g7455);
  not NOT_2579(g8235,I14492);
  not NOT_2580(g2313,I6096);
  not NOT_2581(g6742,I12120);
  not NOT_2582(g1603,I5471);
  not NOT_2583(g6104,g5345);
  not NOT_2584(I14964,g8406);
  not NOT_2585(g6304,I11239);
  not NOT_2586(I15504,g8967);
  not NOT_2587(g2202,g1321);
  not NOT_2588(I12138,g5874);
  not NOT_2589(g4922,g4111);
  not NOT_2590(I10587,g5439);
  not NOT_2591(I13752,g7315);
  not NOT_2592(I11374,g5844);
  not NOT_2593(g3847,I7344);
  not NOT_2594(g2908,g2290);
  not NOT_2595(g5480,g4913);
  not NOT_2596(I6425,g1811);
  not NOT_2597(g5713,g4841);
  not NOT_2598(g4581,g2921);
  not NOT_2599(I12415,g6410);
  not NOT_2600(g3700,g2514);
  not NOT_2601(g9042,I15530);
  not NOT_2602(g2494,g9);
  not NOT_2603(I7953,g3542);
  not NOT_2604(g6754,I12135);
  not NOT_2605(g1583,g718);
  not NOT_2606(g5569,I10028);
  not NOT_2607(g4597,I8706);
  not NOT_2608(I9564,g4703);
  not NOT_2609(I5894,g86);
  not NOT_2610(I11669,g5918);
  not NOT_2611(g7708,I14005);
  not NOT_2612(I13669,g7240);
  not NOT_2613(g9233,I15953);
  not NOT_2614(g7520,I13740);
  not NOT_2615(g8792,I14996);
  not NOT_2616(I11260,g5779);
  not NOT_2617(g6613,I11835);
  not NOT_2618(g3950,g3131);
  not NOT_2619(g4784,I9095);
  not NOT_2620(I10569,g5417);
  not NOT_2621(g4739,I9053);
  not NOT_2622(I11392,g5800);
  not NOT_2623(g1952,g1333);
  not NOT_2624(I9910,g4681);
  not NOT_2625(g6269,I11090);
  not NOT_2626(g5688,I10193);
  not NOT_2627(I6006,g306);
  not NOT_2628(I15533,g9002);
  not NOT_2629(g2965,g2384);
  not NOT_2630(g6983,I12722);
  not NOT_2631(g1616,I5478);
  not NOT_2632(I14747,g8175);
  not NOT_2633(g7176,I13084);
  not NOT_2634(I5475,g1084);
  not NOT_2635(I7716,g3038);
  not NOT_2636(g6572,I11764);
  not NOT_2637(g6862,I12457);
  not NOT_2638(I11559,g6065);
  not NOT_2639(g4079,I7864);
  not NOT_2640(I11525,g5874);
  not NOT_2641(I11488,g6034);
  not NOT_2642(I13559,g7177);
  not NOT_2643(g3562,I7044);
  not NOT_2644(I12484,g6621);
  not NOT_2645(I9609,g4780);
  not NOT_2646(g2264,I5997);
  not NOT_2647(g6712,I12062);
  not NOT_2648(g7405,I13518);
  not NOT_2649(g4668,I8919);
  not NOT_2650(I6087,g318);
  not NOT_2651(I6305,g1333);
  not NOT_2652(g3631,I7098);
  not NOT_2653(g7829,I14251);
  not NOT_2654(g2360,g1435);
  not NOT_2655(g2933,I6673);
  not NOT_2656(g3723,g2096);
  not NOT_2657(I12609,g6571);
  not NOT_2658(g7286,I13290);
  not NOT_2659(g7765,I14166);
  not NOT_2660(I7198,g2509);
  not NOT_2661(I10807,g5294);
  not NOT_2662(g5000,I9325);
  not NOT_2663(I5646,g883);
  not NOT_2664(g8094,g7705);
  not NOT_2665(I14807,g8603);
  not NOT_2666(g2641,g1587);
  not NOT_2667(I14974,g8442);
  not NOT_2668(I9217,g4443);
  not NOT_2669(I10639,g5224);
  not NOT_2670(g4501,g2801);
  not NOT_2671(g6729,g6263);
  not NOT_2672(g6961,I12684);
  not NOT_2673(I13544,g1167);
  not NOT_2674(g3605,g1938);
  not NOT_2675(I13865,g7333);
  not NOT_2676(g2996,g1828);
  not NOT_2677(I9466,g3943);
  not NOT_2678(g5760,I10353);
  not NOT_2679(g9189,I15845);
  not NOT_2680(g7733,I14070);
  not NOT_2681(I12921,g6993);
  not NOT_2682(I13713,g7341);
  not NOT_2683(g9389,I16183);
  not NOT_2684(g1970,I5831);
  not NOT_2685(I6226,g408);
  not NOT_2686(g7270,I13250);
  not NOT_2687(I8805,g3976);
  not NOT_2688(I10265,g5468);
  not NOT_2689(I8916,g4195);
  not NOT_2690(g1925,g825);
  not NOT_2691(g8776,g8585);
  not NOT_2692(g2724,g1814);
  not NOT_2693(g7225,g6936);
  not NOT_2694(g7610,g7450);
  not NOT_2695(g9029,I15501);
  not NOT_2696(g6014,I10614);
  not NOT_2697(I14416,g7727);
  not NOT_2698(g2379,I6239);
  not NOT_2699(I13610,g7227);
  not NOT_2700(I12813,g6607);
  not NOT_2701(I16145,g9367);
  not NOT_2702(g6885,I12526);
  not NOT_2703(I6045,g309);
  not NOT_2704(g4704,I9001);
  not NOT_2705(I13042,g6963);
  not NOT_2706(g6660,I11958);
  not NOT_2707(g6946,I12649);
  not NOT_2708(I13255,g7057);
  not NOT_2709(g2878,g2233);
  not NOT_2710(I13189,g7002);
  not NOT_2711(I7644,g2584);
  not NOT_2712(g5183,I9675);
  not NOT_2713(I13679,g7259);
  not NOT_2714(g7124,g6896);
  not NOT_2715(I12973,g6927);
  not NOT_2716(g5608,g4969);
  not NOT_2717(I9333,g4245);
  not NOT_2718(g2289,I6051);
  not NOT_2719(g6903,I12582);
  not NOT_2720(g2777,g1797);
  not NOT_2721(g9281,I16009);
  not NOT_2722(g5779,I10384);
  not NOT_2723(I10579,g5433);
  not NOT_2724(I9774,g4678);
  not NOT_2725(g4250,I8177);
  not NOT_2726(g2882,g2236);
  not NOT_2727(I11686,g6076);
  not NOT_2728(I11939,g6015);
  not NOT_2729(I7867,g2818);
  not NOT_2730(g9297,I16017);
  not NOT_2731(I13460,g7263);
  not NOT_2732(g4032,I7807);
  not NOT_2733(I11383,g5827);
  not NOT_2734(g2271,I6018);
  not NOT_2735(I9396,g3908);
  not NOT_2736(I13383,g7275);
  not NOT_2737(g1789,g1034);
  not NOT_2738(g7206,I13134);
  not NOT_2739(I6578,g1603);
  not NOT_2740(I6868,g530);
  not NOT_2741(I5616,g979);
  not NOT_2742(g6036,I10643);
  not NOT_2743(I13267,g6913);
  not NOT_2744(g6378,I11461);
  not NOT_2745(I6767,g1933);
  not NOT_2746(g5161,I9609);
  not NOT_2747(I16132,g9356);
  not NOT_2748(I10442,g5215);
  not NOT_2749(I15498,g8974);
  not NOT_2750(g1987,I5842);
  not NOT_2751(g1771,g609);
  not NOT_2752(I7211,g1742);
  not NOT_2753(g7287,I13293);
  not NOT_2754(I14442,g8065);
  not NOT_2755(g6135,I10770);
  not NOT_2756(I5404,g722);
  not NOT_2757(g4568,g2904);
  not NOT_2758(I7386,g3013);
  not NOT_2759(g5665,g4748);
  not NOT_2760(g9109,I15717);
  not NOT_2761(g5051,I9407);
  not NOT_2762(g6335,I11332);
  not NOT_2763(g6831,I12364);
  not NOT_2764(g9309,I16043);
  not NOT_2765(g3531,g1616);
  not NOT_2766(g5127,I9525);
  not NOT_2767(g2674,g1675);
  not NOT_2768(g6288,I11191);
  not NOT_2769(g6382,I11473);
  not NOT_2770(I16161,g9363);
  not NOT_2771(g8179,I14416);
  not NOT_2772(I9018,g3872);
  not NOT_2773(g3743,g1776);
  not NOT_2774(I7599,g2734);
  not NOT_2775(I15924,g9207);
  not NOT_2776(I6015,g437);
  not NOT_2777(I12400,g6767);
  not NOT_2778(g4357,g3679);
  not NOT_2779(g5146,I9564);
  not NOT_2780(g6805,I12286);
  not NOT_2781(g5633,g4895);
  not NOT_2782(I11218,g6161);
  not NOT_2783(I12214,g6507);
  not NOT_2784(g7781,I14214);
  not NOT_2785(g2238,I5975);
  not NOT_2786(g2332,g926);
  not NOT_2787(I10430,g5211);
  not NOT_2788(I13837,g7324);
  not NOT_2789(g3856,I7371);
  not NOT_2790(g2680,g1665);
  not NOT_2791(I14430,g7836);
  not NOT_2792(g2209,I5926);
  not NOT_2793(g2353,g871);
  not NOT_2794(I9493,g4426);
  not NOT_2795(g4929,g4120);
  not NOT_2796(g9201,g9183);
  not NOT_2797(I12328,g6760);
  not NOT_2798(I15753,g9080);
  not NOT_2799(g5696,I10207);
  not NOT_2800(g8882,I15222);
  not NOT_2801(g1945,g1081);
  not NOT_2802(g6947,I12652);
  not NOT_2803(g7510,I13710);
  not NOT_2804(g7245,I13193);
  not NOT_2805(g6798,I12265);
  not NOT_2806(I12538,g6606);
  not NOT_2807(g1738,g741);
  not NOT_2808(g3074,I6800);
  not NOT_2809(I16043,g9285);
  not NOT_2810(g5732,I10253);
  not NOT_2811(g7291,I13305);
  not NOT_2812(g3992,I7723);
  not NOT_2813(I14035,g7310);
  not NOT_2814(I15199,g8792);
  not NOT_2815(I10684,g5258);
  not NOT_2816(I11455,g6087);
  not NOT_2817(g4626,I8793);
  not NOT_2818(I8233,g3588);
  not NOT_2819(I11470,g6095);
  not NOT_2820(g5240,I9752);
  not NOT_2821(g7344,g7150);
  not NOT_2822(I13617,g7276);
  not NOT_2823(g5072,g4457);
  not NOT_2824(g9098,I15684);
  not NOT_2825(I13915,g7360);
  not NOT_2826(g8799,I15007);
  not NOT_2827(I12241,g6640);
  not NOT_2828(I14142,g7551);
  not NOT_2829(g1907,g52);
  not NOT_2830(g5472,I9892);
  not NOT_2831(I9021,g4489);
  not NOT_2832(g6873,I12490);
  not NOT_2833(g7207,I13137);
  not NOT_2834(g6632,I11890);
  not NOT_2835(g6095,I10719);
  not NOT_2836(g3080,g1679);
  not NOT_2837(g8674,I14816);
  not NOT_2838(g6037,I10646);
  not NOT_2839(g3573,g2424);
  not NOT_2840(I15696,g9050);
  not NOT_2841(g3863,I7392);
  not NOT_2842(I5789,g1524);
  not NOT_2843(g1959,g1252);
  not NOT_2844(g2901,g2284);
  not NOT_2845(g7259,g7060);
  not NOT_2846(g6653,I11939);
  not NOT_2847(I13277,g7078);
  not NOT_2848(g6102,g5345);
  not NOT_2849(g6208,I10965);
  not NOT_2850(g6302,I11233);
  not NOT_2851(g8541,g8094);
  not NOT_2852(I13075,g6958);
  not NOT_2853(g2511,g1328);
  not NOT_2854(I7061,g2457);
  not NOT_2855(g6869,I12478);
  not NOT_2856(g1876,g77);
  not NOT_2857(I12771,g6735);
  not NOT_2858(I11467,g6064);
  not NOT_2859(I11494,g6037);
  not NOT_2860(I13595,g7216);
  not NOT_2861(g7488,g7225);
  not NOT_2862(I12235,g6634);
  not NOT_2863(g2092,g1225);
  not NOT_2864(g5434,g5112);
  not NOT_2865(I10193,g4670);
  not NOT_2866(I11037,g5299);
  not NOT_2867(I14130,g7592);
  not NOT_2868(I14193,g7532);
  not NOT_2869(g6752,I12131);
  not NOT_2870(g5147,I9567);
  not NOT_2871(I13782,g7498);
  not NOT_2872(I11984,g6246);
  not NOT_2873(g8802,I15014);
  not NOT_2874(I11419,g5835);
  not NOT_2875(I6428,g1818);
  not NOT_2876(g9019,I15481);
  not NOT_2877(g9362,I16122);
  not NOT_2878(I13419,g7277);
  not NOT_2879(g3857,I7374);
  not NOT_2880(g7951,I14288);
  not NOT_2881(I8706,g3828);
  not NOT_2882(g3976,I7697);
  not NOT_2883(I15225,g8689);
  not NOT_2884(I15708,g9072);
  not NOT_2885(I13822,g7459);
  not NOT_2886(I10475,g5529);
  not NOT_2887(I9301,g4295);
  not NOT_2888(g7114,I12930);
  not NOT_2889(I11266,g5794);
  not NOT_2890(g4661,I8898);
  not NOT_2891(g6786,I12229);
  not NOT_2892(I7145,g2501);
  not NOT_2893(I6564,g2073);
  not NOT_2894(g4075,I7856);
  not NOT_2895(I5945,g333);
  not NOT_2896(I8787,g4012);
  not NOT_2897(g4475,g3818);
  not NOT_2898(g5596,g4841);
  not NOT_2899(g1663,g1416);
  not NOT_2900(I6826,g2185);
  not NOT_2901(g6364,I11419);
  not NOT_2902(g7870,I14270);
  not NOT_2903(g5013,I9341);
  not NOT_2904(g4627,I8796);
  not NOT_2905(I5709,g901);
  not NOT_2906(g8511,I14646);
  not NOT_2907(g9086,I15648);
  not NOT_2908(g1824,I5706);
  not NOT_2909(I5478,g1148);
  not NOT_2910(g6296,I11215);
  not NOT_2911(I11194,g6243);
  not NOT_2912(g4646,I8853);
  not NOT_2913(I7107,g2480);
  not NOT_2914(g2623,g1585);
  not NOT_2915(g6725,I12091);
  not NOT_2916(I9585,g4697);
  not NOT_2917(I10347,g5706);
  not NOT_2918(I10253,g5240);
  not NOT_2919(g5820,I10485);
  not NOT_2920(I7359,g2871);
  not NOT_2921(g9185,I15833);
  not NOT_2922(g4084,I7875);
  not NOT_2923(g4603,I8724);
  not NOT_2924(I5435,g1461);
  not NOT_2925(g7336,I13428);
  not NOT_2926(I13524,g7151);
  not NOT_2927(I15657,g9059);
  not NOT_2928(g9385,I16173);
  not NOT_2929(g8864,I15178);
  not NOT_2930(I15068,g8638);
  not NOT_2931(g7768,I14175);
  not NOT_2932(g1590,I5466);
  not NOT_2933(g1877,g595);
  not NOT_2934(I11401,g5828);
  not NOT_2935(g6553,I11725);
  not NOT_2936(g9070,I15604);
  not NOT_2937(g7594,I13927);
  not NOT_2938(I8745,g3929);
  not NOT_2939(I10236,g5014);
  not NOT_2940(g2375,I6223);
  not NOT_2941(g2871,I6587);
  not NOT_2942(I12725,g6565);
  not NOT_2943(g3220,g1889);
  not NOT_2944(I15337,g8802);
  not NOT_2945(g2651,I6437);
  not NOT_2946(I6217,g105);
  not NOT_2947(g6012,g5367);
  not NOT_2948(g1556,g65);
  not NOT_2949(I13118,g7068);
  not NOT_2950(g3779,g2511);
  not NOT_2951(g4583,g2924);
  not NOT_2952(I11864,g5753);
  not NOT_2953(I14175,g7718);
  not NOT_2954(g2285,I6039);
  not NOT_2955(I7115,g2547);
  not NOT_2956(g6189,I10930);
  not NOT_2957(I8808,g4014);
  not NOT_2958(g6389,I11494);
  not NOT_2959(I7811,g3019);
  not NOT_2960(I16158,g9363);
  not NOT_2961(I9669,g4909);
  not NOT_2962(I13749,g7313);
  not NOT_2963(g7887,I14273);
  not NOT_2964(g7122,I12958);
  not NOT_2965(g4919,g4104);
  not NOT_2966(g3977,g3160);
  not NOT_2967(I6571,g1711);
  not NOT_2968(g6888,I12535);
  not NOT_2969(I6048,g387);
  not NOT_2970(I10516,g5241);
  not NOT_2971(g5581,g4969);
  not NOT_2972(I14264,g7698);
  not NOT_2973(g3588,g2379);
  not NOT_2974(I9531,g4463);
  not NOT_2975(g2184,I5911);
  not NOT_2976(I6711,g1726);
  not NOT_2977(g6371,I11440);
  not NOT_2978(g1785,g615);
  not NOT_2979(g6787,I12232);
  not NOT_2980(g8968,I15408);
  not NOT_2981(g2384,I6254);
  not NOT_2982(I11704,g6076);
  not NOT_2983(g5060,I9422);
  not NOT_2984(I13704,g7352);
  not NOT_2985(I11305,g5807);
  not NOT_2986(g9331,g9321);
  not NOT_2987(g6956,I12669);
  not NOT_2988(I13305,g7168);
  not NOT_2989(g5460,g4684);
  not NOT_2990(g5597,g4969);
  not NOT_2991(I11254,g5793);
  not NOT_2992(g7433,I13562);
  not NOT_2993(g6675,I11981);
  not NOT_2994(g4616,I8763);
  not NOT_2995(I11809,g6285);
  not NOT_2996(I11900,g5847);
  not NOT_2997(g4561,g2900);
  not NOT_2998(g3051,I6791);
  not NOT_2999(I13900,g7356);
  not NOT_3000(I6333,g1345);
  not NOT_3001(I13466,g7122);
  not NOT_3002(I9505,g4300);
  not NOT_3003(g1563,g639);
  not NOT_3004(g2424,g1329);
  not NOT_3005(I12141,g5897);
  not NOT_3006(g2795,g1801);
  not NOT_3007(I8449,g3630);
  not NOT_3008(I12652,g6664);
  not NOT_3009(g9087,I15651);
  not NOT_3010(g9105,I15705);
  not NOT_3011(g5784,I10397);
  not NOT_3012(g4004,g2845);
  not NOT_3013(I15010,g8584);
  not NOT_3014(I15918,g9211);
  not NOT_3015(g9305,I16033);
  not NOT_3016(g5739,I10274);
  not NOT_3017(I8865,g4032);
  not NOT_3018(g7496,I13666);
  not NOT_3019(g4527,g3466);
  not NOT_3020(g7550,I13834);
  not NOT_3021(g6297,I11218);
  not NOT_3022(g3999,I7738);
  not NOT_3023(g4647,I8856);
  not NOT_3024(g8175,I14406);
  not NOT_3025(I8715,g3903);
  not NOT_3026(I7595,g2573);
  not NOT_3027(g8871,I15199);
  not NOT_3028(g3633,I7104);
  not NOT_3029(g2672,I6471);
  not NOT_3030(g2231,I5954);
  not NOT_3031(g7137,I12993);
  not NOT_3032(I14208,g7711);
  not NOT_3033(g8651,I14747);
  not NOT_3034(g2477,g25);
  not NOT_3035(I16017,g9264);
  not NOT_3036(g2643,g1589);
  not NOT_3037(g6684,I11998);
  not NOT_3038(I12135,g5988);
  not NOT_3039(g6639,g6198);
  not NOT_3040(g5668,I10151);
  not NOT_3041(g6338,I11341);
  not NOT_3042(I15598,g8991);
  not NOT_3043(I6509,g1684);
  not NOT_3044(g5294,g5087);
  not NOT_3045(g4503,I8565);
  not NOT_3046(g5840,I10535);
  not NOT_3047(g6963,I12690);
  not NOT_3048(I7978,g3574);
  not NOT_3049(g6791,I12244);
  not NOT_3050(g2205,g13);
  not NOT_3051(I12406,g6773);
  not NOT_3052(g6309,I11254);
  not NOT_3053(g5190,g4938);
  not NOT_3054(g4925,g4114);
  not NOT_3055(I5657,g921);
  not NOT_3056(I12361,g6765);
  not NOT_3057(I7417,g3659);
  not NOT_3058(g3732,g2533);
  not NOT_3059(I6018,g462);
  not NOT_3060(g1557,I5432);
  not NOT_3061(g2634,g1578);
  not NOT_3062(g3753,g2540);
  not NOT_3063(I10614,g5302);
  not NOT_3064(g6808,I12295);
  not NOT_3065(I9573,g4701);
  not NOT_3066(g9045,I15539);
  not NOT_3067(I10436,g5213);
  not NOT_3068(g724,I5401);
  not NOT_3069(I14614,g7832);
  not NOT_3070(g7266,I13238);
  not NOT_3071(g2551,g1360);
  not NOT_3072(I14436,g7904);
  not NOT_3073(g2104,I5879);
  not NOT_3074(g3944,I7635);
  not NOT_3075(I11693,g6076);
  not NOT_3076(g5156,I9594);
  not NOT_3077(g9373,I16145);
  not NOT_3078(g9091,I15663);
  not NOT_3079(g4120,I7967);
  not NOT_3080(I16023,g9267);
  not NOT_3081(I7629,g3633);
  not NOT_3082(g6759,I12148);
  not NOT_3083(I10274,g5524);
  not NOT_3084(I14073,g7627);
  not NOT_3085(I6093,g468);
  not NOT_3086(I8268,g2801);
  not NOT_3087(I13009,g6935);
  not NOT_3088(g1948,g1250);
  not NOT_3089(g8809,I15065);
  not NOT_3090(g7142,I13012);
  not NOT_3091(g6201,I10946);
  not NOT_3092(g2926,g2325);
  not NOT_3093(g7342,I13444);
  not NOT_3094(I11008,g5693);
  not NOT_3095(g9369,I16135);
  not NOT_3096(I10565,g5402);
  not NOT_3097(g6957,I12672);
  not NOT_3098(g7255,I13209);
  not NOT_3099(g4617,I8766);
  not NOT_3100(I8452,g2816);
  not NOT_3101(g649,I5380);
  not NOT_3102(g8672,I14810);
  not NOT_3103(g3316,I6930);
  not NOT_3104(g9059,I15571);
  not NOT_3105(I11476,g6194);
  not NOT_3106(I11485,g6137);
  not NOT_3107(I7800,g2605);
  not NOT_3108(g6449,I11596);
  not NOT_3109(g2273,I6024);
  not NOT_3110(g1814,g630);
  not NOT_3111(g6865,I12466);
  not NOT_3112(I7554,g2573);
  not NOT_3113(g7097,I12881);
  not NOT_3114(g7726,I14049);
  not NOT_3115(I13454,g7147);
  not NOT_3116(g7497,I13669);
  not NOT_3117(I10292,g5577);
  not NOT_3118(g2044,I5861);
  not NOT_3119(g7354,I13478);
  not NOT_3120(g5163,I9615);
  not NOT_3121(g6604,I11818);
  not NOT_3122(g5810,I10463);
  not NOT_3123(I13570,g7198);
  not NOT_3124(I6021,g495);
  not NOT_3125(g6498,I11666);
  not NOT_3126(g2269,I6012);
  not NOT_3127(g1773,g610);
  not NOT_3128(I8486,g2824);
  not NOT_3129(I10409,g5204);
  not NOT_3130(g4547,g3466);
  not NOT_3131(g5053,g4438);
  not NOT_3132(g6833,I12370);
  not NOT_3133(I8730,g3987);
  not NOT_3134(g3533,g2397);
  not NOT_3135(g5453,g4680);
  not NOT_3136(g2862,I6578);
  not NOT_3137(I15631,g9003);
  not NOT_3138(I12463,g6682);
  not NOT_3139(g4892,I9250);
  not NOT_3140(I11239,g6173);
  not NOT_3141(g2712,g2039);
  not NOT_3142(I14136,g7633);
  not NOT_3143(g9227,I15947);
  not NOT_3144(g1769,I5609);
  not NOT_3145(I9126,g3870);
  not NOT_3146(I7902,g2709);
  not NOT_3147(g2543,g1348);
  not NOT_3148(g6896,I12561);
  not NOT_3149(I13238,g6900);
  not NOT_3150(I9760,g4838);
  not NOT_3151(g3013,I6764);
  not NOT_3152(g1918,g822);
  not NOT_3153(g1967,g1432);
  not NOT_3154(g7112,I12924);
  not NOT_3155(g7267,I13241);
  not NOT_3156(I5966,g278);
  not NOT_3157(g5157,I9597);
  not NOT_3158(g2961,I6711);
  not NOT_3159(g4738,I9050);
  not NOT_3160(g8754,g8524);
  not NOT_3161(I5471,g1029);
  not NOT_3162(g6019,g5367);
  not NOT_3163(g6362,I11413);
  not NOT_3164(I13185,g7020);
  not NOT_3165(I6723,g2052);
  not NOT_3166(I13092,g7047);
  not NOT_3167(g7293,I13311);
  not NOT_3168(g2927,I6663);
  not NOT_3169(I12514,g6605);
  not NOT_3170(I5948,g378);
  not NOT_3171(g3936,I7605);
  not NOT_3172(I13518,g7141);
  not NOT_3173(g7129,I12973);
  not NOT_3174(I15571,g8982);
  not NOT_3175(I15308,g8799);
  not NOT_3176(g1822,g761);
  not NOT_3177(g7329,I13407);
  not NOT_3178(g7761,I14154);
  not NOT_3179(g4907,g4087);
  not NOT_3180(g2885,g2239);
  not NOT_3181(g4035,I7814);
  not NOT_3182(g2660,I6451);
  not NOT_3183(g2946,g2365);
  not NOT_3184(I12421,g6486);
  not NOT_3185(I14109,g7590);
  not NOT_3186(g7727,I14052);
  not NOT_3187(I15495,g8973);
  not NOT_3188(g4482,I8520);
  not NOT_3189(I7964,g3488);
  not NOT_3190(g2903,g2286);
  not NOT_3191(g5626,g4748);
  not NOT_3192(g7592,I13921);
  not NOT_3193(I8766,g3960);
  not NOT_3194(I9588,g4704);
  not NOT_3195(g6486,I11648);
  not NOT_3196(I8105,g3339);
  not NOT_3197(I10283,g5643);
  not NOT_3198(g4656,I8883);
  not NOT_3199(g7746,I14109);
  not NOT_3200(g6730,I12098);
  not NOT_3201(g9188,I15842);
  not NOT_3202(g7221,I13157);
  not NOT_3203(I15687,g9071);
  not NOT_3204(g9388,I16180);
  not NOT_3205(g3922,I7561);
  not NOT_3206(I15985,g9237);
  not NOT_3207(I14492,g7829);
  not NOT_3208(g9216,I15924);
  not NOT_3209(g6385,I11482);
  not NOT_3210(g6881,I12514);
  not NOT_3211(I12541,g6614);
  not NOT_3212(I8748,g3997);
  not NOT_3213(g4915,g4094);
  not NOT_3214(I11215,g6156);
  not NOT_3215(g9028,I15498);
  not NOT_3216(g6070,g5317);
  not NOT_3217(I11729,g5772);
  not NOT_3218(g1895,I5775);
  not NOT_3219(g6897,I12564);
  not NOT_3220(g1837,g1007);
  not NOT_3221(I13577,g7186);
  not NOT_3222(g9030,I15504);
  not NOT_3223(g6025,g5367);
  not NOT_3224(I6673,g2246);
  not NOT_3225(g6425,I11556);
  not NOT_3226(I14381,g7596);
  not NOT_3227(I13728,g7439);
  not NOT_3228(g5683,I10180);
  not NOT_3229(I12325,g6755);
  not NOT_3230(I9633,g4800);
  not NOT_3231(g2288,I6048);
  not NOT_3232(I7118,g2484);
  not NOT_3233(I7167,g2505);
  not NOT_3234(I14091,g7589);
  not NOT_3235(g2382,I6248);
  not NOT_3236(g7068,g6556);
  not NOT_3237(I12829,g6441);
  not NOT_3238(I12535,g6599);
  not NOT_3239(I15669,g9045);
  not NOT_3240(g3784,g1768);
  not NOT_3241(I10796,g5397);
  not NOT_3242(g8014,g7564);
  not NOT_3243(I9103,g4374);
  not NOT_3244(I12358,g6761);
  not NOT_3245(I13438,g7143);
  not NOT_3246(g3739,g2536);
  not NOT_3247(I6669,g1698);
  not NOT_3248(g4663,I8904);
  not NOT_3249(I6368,g20);
  not NOT_3250(g2916,I6646);
  not NOT_3251(I15842,g9171);
  not NOT_3252(I8373,g3783);
  not NOT_3253(g5735,I10262);
  not NOT_3254(g1788,g984);
  not NOT_3255(g3995,I7728);
  not NOT_3256(g3937,g2845);
  not NOT_3257(g8903,I15315);
  not NOT_3258(g3079,g1603);
  not NOT_3259(g5782,I10393);
  not NOT_3260(g4002,g3192);
  not NOT_3261(I10390,g5195);
  not NOT_3262(I13906,g7358);
  not NOT_3263(I11284,g5795);
  not NOT_3264(I13284,g7156);
  not NOT_3265(g6131,g5529);
  not NOT_3266(g7576,I13873);
  not NOT_3267(g6331,I11320);
  not NOT_3268(g5075,I9443);
  not NOT_3269(g3840,I7323);
  not NOT_3270(g2947,I6695);
  not NOT_3271(g7716,I14025);
  not NOT_3272(g7149,I13031);
  not NOT_3273(g2798,g1787);
  not NOT_3274(I11622,g5847);
  not NOT_3275(g1842,g764);
  not NOT_3276(g7349,I13463);
  not NOT_3277(g6635,I11897);
  not NOT_3278(I13622,g7279);
  not NOT_3279(g9108,I15714);
  not NOT_3280(g3390,I6949);
  not NOT_3281(g9308,I16040);
  not NOT_3282(I8868,g4035);
  not NOT_3283(g5627,g4673);
  not NOT_3284(g6682,I11994);
  not NOT_3285(g6766,I12167);
  not NOT_3286(g6087,I10705);
  not NOT_3287(I12173,g5918);
  not NOT_3288(g8178,I14413);
  not NOT_3289(g6305,I11242);
  not NOT_3290(g6801,I12274);
  not NOT_3291(I6856,g449);
  not NOT_3292(g4590,g2932);
  not NOT_3293(I10522,g5243);
  not NOT_3294(I15830,g9180);
  not NOT_3295(I8718,g3909);
  not NOT_3296(g3501,g2185);
  not NOT_3297(I9443,g4564);
  not NOT_3298(g5526,g5086);
  not NOT_3299(g7198,I13126);
  not NOT_3300(g4657,I8886);
  not NOT_3301(g7747,I14112);
  not NOT_3302(g7855,I14267);
  not NOT_3303(g9217,I15927);
  not NOT_3304(g2873,g1779);
  not NOT_3305(g1854,g773);
  not NOT_3306(g2632,g1576);
  not NOT_3307(I9116,g4297);
  not NOT_3308(I8261,g3643);
  not NOT_3309(g4556,g2895);
  not NOT_3310(g9066,I15592);
  not NOT_3311(I13653,g7246);
  not NOT_3312(g5084,g4477);
  not NOT_3313(g5603,g4938);
  not NOT_3314(g1941,I5812);
  not NOT_3315(I6474,g1941);
  not NOT_3316(g2495,g26);
  not NOT_3317(I8793,g3923);
  not NOT_3318(I9034,g4317);
  not NOT_3319(g2653,I6443);
  not NOT_3320(g7241,I13185);
  not NOT_3321(g6755,I12138);
  not NOT_3322(g2208,I5923);
  not NOT_3323(g3942,I7629);
  not NOT_3324(I12760,g6685);
  not NOT_3325(g5439,g5058);
  not NOT_3326(g4928,g4119);
  not NOT_3327(I10862,g5364);
  not NOT_3328(g6226,g5658);
  not NOT_3329(g4930,g4121);
  not NOT_3330(g8916,I15334);
  not NOT_3331(g2869,g2224);
  not NOT_3332(I15610,g8995);
  not NOT_3333(I15705,g9068);
  not NOT_3334(I10949,g5513);
  not NOT_3335(g9048,I15546);
  not NOT_3336(g4899,g4080);
  not NOT_3337(g4464,I8486);
  not NOT_3338(I9347,g3896);
  not NOT_3339(g1708,I5552);
  not NOT_3340(I9681,g4811);
  not NOT_3341(g7524,I13752);
  not NOT_3342(g6173,I10882);
  not NOT_3343(g2752,g2389);
  not NOT_3344(g3954,I7655);
  not NOT_3345(g6373,I11446);
  not NOT_3346(I10702,g5529);
  not NOT_3347(I15678,g9060);
  not NOT_3348(g9133,I15773);
  not NOT_3349(g2917,g2309);
  not NOT_3350(g9333,g9323);
  not NOT_3351(g7119,I12945);
  not NOT_3352(g1812,I5682);
  not NOT_3353(g7319,g7124);
  not NOT_3354(I14904,g8629);
  not NOT_3355(I8721,g3918);
  not NOT_3356(g1958,g786);
  not NOT_3357(g2265,I6000);
  not NOT_3358(g6369,I11434);
  not NOT_3359(g7352,I13472);
  not NOT_3360(g7577,I13876);
  not NOT_3361(g6007,g5494);
  not NOT_3362(I12927,g7014);
  not NOT_3363(g9196,g9185);
  not NOT_3364(g7717,I14028);
  not NOT_3365(g6059,g5317);
  not NOT_3366(g6868,I12475);
  not NOT_3367(g5616,g4938);
  not NOT_3368(g3568,g1935);
  not NOT_3369(g8873,I15205);
  not NOT_3370(I13484,g7128);
  not NOT_3371(g1829,I5715);
  not NOT_3372(g8632,I14712);
  not NOT_3373(I5842,g68);
  not NOT_3374(I15065,g8636);
  not NOT_3375(g6767,I12170);
  not NOT_3376(g2364,I6192);
  not NOT_3377(I12649,g6457);
  not NOT_3378(g2233,I5960);
  not NOT_3379(I10183,g5129);
  not NOT_3380(g1911,I5789);
  not NOT_3381(I10397,g5200);
  not NOT_3382(g7211,I13147);
  not NOT_3383(I5392,g694);
  not NOT_3384(g3912,g3192);
  not NOT_3385(I14397,g7686);
  not NOT_3386(g4089,I7888);
  not NOT_3387(I12903,g6905);
  not NOT_3388(g2454,I6294);
  not NOT_3389(I11200,g6251);
  not NOT_3390(g8869,I15193);
  not NOT_3391(g4489,g2826);
  not NOT_3392(g2770,g2210);
  not NOT_3393(g6793,I12250);
  not NOT_3394(I10509,g5237);
  not NOT_3395(g9018,I15478);
  not NOT_3396(g4557,g2896);
  not NOT_3397(g5764,I10369);
  not NOT_3398(g7599,g7450);
  not NOT_3399(g9067,I15595);
  not NOT_3400(g1974,g803);
  not NOT_3401(I10933,g5668);
  not NOT_3402(g7274,I13258);
  not NOT_3403(I15218,g8801);
  not NOT_3404(g6015,I10617);
  not NOT_3405(g4071,I7850);
  not NOT_3406(I6000,g202);
  not NOT_3407(I7341,g2931);
  not NOT_3408(g2532,I6358);
  not NOT_3409(g8752,g8564);
  not NOT_3410(g6227,I11018);
  not NOT_3411(g3929,I7588);
  not NOT_3412(I13921,g7362);
  not NOT_3413(I6326,g1443);
  not NOT_3414(I14851,g8630);
  not NOT_3415(g8917,I15337);
  not NOT_3416(g1796,g617);
  not NOT_3417(g4242,I8161);
  not NOT_3418(g7125,I12965);
  not NOT_3419(g9093,I15669);
  not NOT_3420(I8428,g3611);
  not NOT_3421(g6246,I11055);
  not NOT_3422(I7691,g3651);
  not NOT_3423(I15160,g8631);
  not NOT_3424(I13813,g7314);
  not NOT_3425(g8042,I14325);
  not NOT_3426(g5224,g5114);
  not NOT_3427(g7280,I13274);
  not NOT_3428(g8442,I14623);
  not NOT_3429(g6721,g6257);
  not NOT_3430(g8786,g8545);
  not NOT_3431(g5120,I9512);
  not NOT_3432(I12262,g6656);
  not NOT_3433(g2389,g1230);
  not NOT_3434(g9181,g9177);
  not NOT_3435(g2706,g1821);
  not NOT_3436(g7544,I13816);
  not NOT_3437(I8826,g4023);
  not NOT_3438(g9381,I16165);
  not NOT_3439(I5812,g1243);
  not NOT_3440(g7483,g7226);
  not NOT_3441(I15915,g9194);
  not NOT_3442(I9460,g3941);
  not NOT_3443(I9597,g4738);
  not NOT_3444(I6183,g6);
  not NOT_3445(g4350,I8315);
  not NOT_3446(g2888,I6608);
  not NOT_3447(I6608,g1612);
  not NOT_3448(g9197,g9186);
  not NOT_3449(I6220,g126);
  not NOT_3450(I10574,g5426);
  not NOT_3451(g2371,g944);
  not NOT_3452(I8910,g4200);
  not NOT_3453(g2787,g1807);
  not NOT_3454(g4438,I8446);
  not NOT_3455(g7106,I12906);
  not NOT_3456(I11732,g6076);
  not NOT_3457(g5617,g4969);
  not NOT_3458(g8770,g8545);
  not NOT_3459(g6502,I11672);
  not NOT_3460(I14205,g7710);
  not NOT_3461(g7306,I13350);
  not NOT_3462(g5789,I10412);
  not NOT_3463(g4009,I7758);
  not NOT_3464(g2956,g2375);
  not NOT_3465(I16119,g9351);
  not NOT_3466(I14311,g7566);
  not NOT_3467(g7790,I14227);
  not NOT_3468(g5516,g4924);
  not NOT_3469(I15595,g8990);
  not NOT_3470(g6940,I12639);
  not NOT_3471(I5911,g216);
  not NOT_3472(I8308,g3674);
  not NOT_3473(g7061,g6650);
  not NOT_3474(g7187,I13103);
  not NOT_3475(I7311,g2879);
  not NOT_3476(g5987,g5294);
  not NOT_3477(g1849,I5732);
  not NOT_3478(g3778,g2145);
  not NOT_3479(I13692,g7343);
  not NOT_3480(I13761,g7418);
  not NOT_3481(g642,I5377);
  not NOT_3482(I8883,g4198);
  not NOT_3483(g7756,I14139);
  not NOT_3484(g6388,I11491);
  not NOT_3485(I10592,g5444);
  not NOT_3486(g5299,I9804);
  not NOT_3487(I9840,g4702);
  not NOT_3488(g3735,g1961);
  not NOT_3489(g4918,g4103);
  not NOT_3490(g6216,I10987);
  not NOT_3491(g1781,g622);
  not NOT_3492(I6051,g440);
  not NOT_3493(I7374,g3084);
  not NOT_3494(I10780,g5445);
  not NOT_3495(g8012,I14305);
  not NOT_3496(I6127,g471);
  not NOT_3497(I6451,g1895);
  not NOT_3498(g6028,g5529);
  not NOT_3499(I14780,g8284);
  not NOT_3500(I12247,g6646);
  not NOT_3501(g6671,I11971);
  not NOT_3502(g7904,I14276);
  not NOT_3503(g1797,g627);
  not NOT_3504(g2639,g1583);
  not NOT_3505(g7046,I12806);
  not NOT_3506(I11329,g5825);
  not NOT_3507(g3075,g2216);
  not NOT_3508(g2963,g2383);
  not NOT_3509(g4229,I8140);
  not NOT_3510(I10350,g5707);
  not NOT_3511(I13329,g7247);
  not NOT_3512(g7446,I13595);
  not NOT_3513(g7514,I13722);
  not NOT_3514(g3949,I7644);
  not NOT_3515(g2309,I6084);
  not NOT_3516(g9101,I15693);
  not NOT_3517(I7545,g3589);
  not NOT_3518(I12388,g6403);
  not NOT_3519(g9301,g9260);
  not NOT_3520(g4822,I9177);
  not NOT_3521(g7145,I13023);
  not NOT_3522(g8029,I14318);
  not NOT_3523(I7380,g3461);
  not NOT_3524(g7345,I13451);
  not NOT_3525(I12098,g5956);
  not NOT_3526(g8787,g8564);
  not NOT_3527(I16036,g9282);
  not NOT_3528(I7832,g2768);
  not NOT_3529(g5738,I10271);
  not NOT_3530(g6826,I12349);
  not NOT_3531(g7763,I14160);
  not NOT_3532(g3526,g2185);
  not NOT_3533(g8956,I15382);
  not NOT_3534(g3998,g3097);
  not NOT_3535(g8675,I14819);
  not NOT_3536(g5709,g4841);
  not NOT_3537(I8333,g3721);
  not NOT_3538(g6741,I12117);
  not NOT_3539(I15589,g8988);
  not NOT_3540(g3084,I6820);
  not NOT_3541(g3603,g2092);
  not NOT_3542(I5377,g635);
  not NOT_3543(g785,I5407);
  not NOT_3544(g5478,g5025);
  not NOT_3545(I13241,g7030);
  not NOT_3546(I14413,g7723);
  not NOT_3547(g1694,g21);
  not NOT_3548(g7107,I12909);
  not NOT_3549(g4921,g4202);
  not NOT_3550(g7307,I13353);
  not NOT_3551(g3850,I7353);
  not NOT_3552(I15836,g9165);
  not NOT_3553(g2957,g2376);
  not NOT_3554(I8196,g3654);
  not NOT_3555(g7159,I13051);
  not NOT_3556(I7931,g2780);
  not NOT_3557(g1852,g887);
  not NOT_3558(g1923,I5801);
  not NOT_3559(I6072,g1211);
  not NOT_3560(g6108,g5345);
  not NOT_3561(g7359,I13493);
  not NOT_3562(I9250,g4134);
  not NOT_3563(g5435,g5121);
  not NOT_3564(g6308,I11251);
  not NOT_3565(g5517,g4925);
  not NOT_3566(g5690,g4748);
  not NOT_3567(I9363,g4258);
  not NOT_3568(g7223,I13161);
  not NOT_3569(g5482,g4915);
  not NOT_3570(g1701,I5545);
  not NOT_3571(g6883,I12520);
  not NOT_3572(I9053,g4327);
  not NOT_3573(g8684,I14848);
  not NOT_3574(g3583,g2128);
  not NOT_3575(g4895,g4078);
  not NOT_3576(g8639,I14725);
  not NOT_3577(I6443,g1774);
  not NOT_3578(g7757,I14142);
  not NOT_3579(I7905,g2863);
  not NOT_3580(I11683,g5988);
  not NOT_3581(g4620,I8775);
  not NOT_3582(g8791,g8585);
  not NOT_3583(g4462,I8480);
  not NOT_3584(g2498,I6333);
  not NOT_3585(g6217,g5649);
  not NOT_3586(g3919,I7554);
  not NOT_3587(g6758,I12145);
  not NOT_3588(g6589,g6083);
  not NOT_3589(g1886,I5766);
  not NOT_3590(I7204,g2520);
  not NOT_3591(I16009,g9261);
  not NOT_3592(I15616,g8997);
  not NOT_3593(I5781,g979);
  not NOT_3594(g2833,I6561);
  not NOT_3595(g7522,I13746);
  not NOT_3596(g7115,I12933);
  not NOT_3597(g7251,I13203);
  not NOT_3598(g8808,I15062);
  not NOT_3599(I6434,g1830);
  not NOT_3600(g3952,I7651);
  not NOT_3601(g7315,I13373);
  not NOT_3602(g7811,I14238);
  not NOT_3603(g7047,g6498);
  not NOT_3604(g9368,I16132);
  not NOT_3605(I8994,g4565);
  not NOT_3606(I10046,g4840);
  not NOT_3607(g6861,I12454);
  not NOT_3608(g6365,I11422);
  not NOT_3609(g2584,g1646);
  not NOT_3610(I14046,g7492);
  not NOT_3611(g4788,I9103);
  not NOT_3612(g6048,g5246);
  not NOT_3613(I11515,g5897);
  not NOT_3614(I11991,g5939);
  not NOT_3615(g2539,I6363);
  not NOT_3616(g2896,g2269);
  not NOT_3617(g3561,I7041);
  not NOT_3618(g9058,I15568);
  not NOT_3619(I13515,g7152);
  not NOT_3620(g8759,g8524);
  not NOT_3621(I13882,g7350);
  not NOT_3622(g6711,I12059);
  not NOT_3623(g1870,I5751);
  not NOT_3624(I11407,g5841);
  not NOT_3625(I13407,g7271);
  not NOT_3626(g1825,I5709);
  not NOT_3627(g6827,I12352);
  not NOT_3628(g3527,g1616);
  not NOT_3629(g8957,I15385);
  not NOT_3630(g6133,I10766);
  not NOT_3631(g6333,I11326);
  not NOT_3632(I14282,g7709);
  not NOT_3633(g3647,g2424);
  not NOT_3634(I9929,g5052);
  not NOT_3635(g2162,I5901);
  not NOT_3636(I7973,g3071);
  not NOT_3637(g2268,I6009);
  not NOT_3638(g6774,I12193);
  not NOT_3639(g2362,I6186);
  not NOT_3640(I12629,g6523);
  not NOT_3641(g3764,g2039);
  not NOT_3642(g4085,I7878);
  not NOT_3643(I12451,g6524);
  not NOT_3644(g6846,I12409);
  not NOT_3645(I12472,g6591);
  not NOT_3646(I12220,g6645);
  not NOT_3647(g8865,I15181);
  not NOT_3648(g3546,I7029);
  not NOT_3649(g5002,g4335);
  not NOT_3650(I14743,g8174);
  not NOT_3651(I8847,g4025);
  not NOT_3652(g2052,I5865);
  not NOT_3653(g5402,g5000);
  not NOT_3654(g5824,I10497);
  not NOT_3655(g7595,I13930);
  not NOT_3656(g6803,I12280);
  not NOT_3657(g2452,g23);
  not NOT_3658(g8604,I14677);
  not NOT_3659(g3503,g2407);
  not NOT_3660(g3970,g2845);
  not NOT_3661(g1768,g605);
  not NOT_3662(g9074,I15616);
  not NOT_3663(g6538,I11714);
  not NOT_3664(I13441,g7146);
  not NOT_3665(I5852,g1202);
  not NOT_3666(I5923,g252);
  not NOT_3667(I11206,g6133);
  not NOT_3668(I7323,g2905);
  not NOT_3669(g6780,I12211);
  not NOT_3670(g6509,I11689);
  not NOT_3671(g1806,I5670);
  not NOT_3672(g1943,g1025);
  not NOT_3673(I6820,g1707);
  not NOT_3674(g7243,I13189);
  not NOT_3675(I6936,g1878);
  not NOT_3676(I11725,g6036);
  not NOT_3677(I12776,g6739);
  not NOT_3678(I13725,g7437);
  not NOT_3679(g2728,g2256);
  not NOT_3680(g2486,g959);
  not NOT_3681(g6662,I11964);
  not NOT_3682(g6018,g5494);
  not NOT_3683(I6317,g1339);
  not NOT_3684(g1887,g83);
  not NOT_3685(I16176,g9385);
  not NOT_3686(I13758,g7414);
  not NOT_3687(I15693,g9048);
  not NOT_3688(I12355,g6756);
  not NOT_3689(I13435,g7170);
  not NOT_3690(g1934,g154);
  not NOT_3691(g2185,I5914);
  not NOT_3692(g6290,I11197);
  not NOT_3693(g4640,I8835);
  not NOT_3694(g2881,g2235);
  not NOT_3695(I7648,g2712);
  not NOT_3696(I16154,g9370);
  not NOT_3697(I7875,g3819);
  not NOT_3698(I12370,g6758);
  not NOT_3699(g4031,I7804);
  not NOT_3700(g7130,I12976);
  not NOT_3701(I7655,g2734);
  not NOT_3702(g3617,g1655);
  not NOT_3703(g6093,g5345);
  not NOT_3704(I11744,g6120);
  not NOT_3705(g7542,I13810);
  not NOT_3706(g2470,g42);
  not NOT_3707(g7330,I13410);
  not NOT_3708(g2897,g2270);
  not NOT_3709(g6493,I11659);
  not NOT_3710(g6256,I11069);
  not NOT_3711(I12151,g5847);
  not NOT_3712(g6816,I12319);
  not NOT_3713(g5785,I10400);
  not NOT_3714(I12996,g6934);
  not NOT_3715(g4005,I7746);
  not NOT_3716(I13940,g7355);
  not NOT_3717(I8101,g3259);
  not NOT_3718(I8817,g3935);
  not NOT_3719(I14662,g7783);
  not NOT_3720(g3987,I7716);
  not NOT_3721(g3771,g1853);
  not NOT_3722(I11848,g6159);
  not NOT_3723(I9782,g4720);
  not NOT_3724(I11398,g5823);
  not NOT_3725(I12367,g6754);
  not NOT_3726(I12394,g6759);
  not NOT_3727(I6060,g580);
  not NOT_3728(g6381,I11470);
  not NOT_3729(g4286,g3790);
  not NOT_3730(I11652,g5939);
  not NOT_3731(g6847,I12412);
  not NOT_3732(I6460,g2104);
  not NOT_3733(I6597,g1970);
  not NOT_3734(I10482,g5228);
  not NOT_3735(g3547,g2345);
  not NOT_3736(g6700,g6244);
  not NOT_3737(g6397,I11512);
  not NOT_3738(I10552,g5396);
  not NOT_3739(I8751,g4009);
  not NOT_3740(g3892,g3131);
  not NOT_3741(I11263,g5784);
  not NOT_3742(I10204,g5060);
  not NOT_3743(I9627,g4777);
  not NOT_3744(g2131,g1300);
  not NOT_3745(I6784,g2052);
  not NOT_3746(g2006,g806);
  not NOT_3747(g2331,g933);
  not NOT_3748(I12319,g6741);
  not NOT_3749(g4733,g4202);
  not NOT_3750(I11332,g5832);
  not NOT_3751(g5844,I10545);
  not NOT_3752(I13332,g7241);
  not NOT_3753(g6263,g5688);
  not NOT_3754(g4270,g2573);
  not NOT_3755(I5972,g356);
  not NOT_3756(g2635,g1579);
  not NOT_3757(g1807,g619);
  not NOT_3758(g6950,I12659);
  not NOT_3759(g8881,g8683);
  not NOT_3760(g9126,I15756);
  not NOT_3761(g4610,I8745);
  not NOT_3762(g2105,g1444);
  not NOT_3763(I7667,g3052);
  not NOT_3764(g3945,g3097);
  not NOT_3765(I12059,g5874);
  not NOT_3766(I10786,g5452);
  not NOT_3767(I12025,g5918);
  not NOT_3768(g2487,I6323);
  not NOT_3769(I9084,g4358);
  not NOT_3770(g5731,I10250);
  not NOT_3771(I9603,g4719);
  not NOT_3772(I13962,g7413);
  not NOT_3773(I14786,g8606);
  not NOT_3774(g7512,I13716);
  not NOT_3775(I9484,g3957);
  not NOT_3776(g3991,g3160);
  not NOT_3777(g7090,g6525);
  not NOT_3778(I6294,g1330);
  not NOT_3779(I9850,g4798);
  not NOT_3780(g594,I5368);
  not NOT_3781(I10356,g5711);
  not NOT_3782(I15382,g8883);
  not NOT_3783(I11500,g6219);
  not NOT_3784(g6562,I11736);
  not NOT_3785(g7366,I13512);
  not NOT_3786(g4069,I7844);
  not NOT_3787(I15519,g9019);
  not NOT_3788(g5071,g4438);
  not NOT_3789(g3078,g1603);
  not NOT_3790(g3340,g2474);
  not NOT_3791(I10826,g5434);
  not NOT_3792(I15675,g9058);
  not NOT_3793(I10380,g5448);
  not NOT_3794(g5705,g4841);
  not NOT_3795(g5471,I9889);
  not NOT_3796(g7056,g6520);
  not NOT_3797(g6631,I11887);
  not NOT_3798(g4540,g2882);
  not NOT_3799(g2226,g1320);
  not NOT_3800(I7548,g3590);
  not NOT_3801(I10998,g5672);
  not NOT_3802(I12044,g5847);
  not NOT_3803(g6723,I12085);
  not NOT_3804(g7456,g7174);
  not NOT_3805(I13048,g6956);
  not NOT_3806(g7529,I13767);
  not NOT_3807(g6257,g5685);
  not NOT_3808(g3959,g3097);
  not NOT_3809(g1815,g760);
  not NOT_3810(g6101,g5317);
  not NOT_3811(g7148,I13028);
  not NOT_3812(g6817,I12322);
  not NOT_3813(g9183,g9161);
  not NOT_3814(g6301,I11230);
  not NOT_3815(g7348,I13460);
  not NOT_3816(g3517,g2283);
  not NOT_3817(I11004,g5613);
  not NOT_3818(g3082,g1680);
  not NOT_3819(g9383,g9380);
  not NOT_3820(I8772,g4011);
  not NOT_3821(I7804,g3029);
  not NOT_3822(g9220,g9205);
  not NOT_3823(I11221,g6167);
  not NOT_3824(g7155,I13039);
  not NOT_3825(g7355,I13481);
  not NOT_3826(g6605,I11821);
  not NOT_3827(I7792,g3038);
  not NOT_3828(I12301,g6703);
  not NOT_3829(g8678,I14828);
  not NOT_3830(g1726,g158);
  not NOT_3831(g3876,g3466);
  not NOT_3832(g8131,I14378);
  not NOT_3833(I12120,g5939);
  not NOT_3834(g2373,I6217);
  not NOT_3835(g2091,g819);
  not NOT_3836(g8406,I14614);
  not NOT_3837(I13613,g7273);
  not NOT_3838(g1960,g1268);
  not NOT_3839(g5814,I10475);
  not NOT_3840(g7260,g7064);
  not NOT_3841(g6751,I12128);
  not NOT_3842(g5150,I9576);
  not NOT_3843(I8011,g3225);
  not NOT_3844(I9561,g4695);
  not NOT_3845(g8682,I14844);
  not NOT_3846(g8766,g8545);
  not NOT_3847(g5038,g4457);
  not NOT_3848(I5395,g698);
  not NOT_3849(I8856,g3955);
  not NOT_3850(g2283,I6033);
  not NOT_3851(g7063,I12826);
  not NOT_3852(I12699,g6504);
  not NOT_3853(g9161,I15803);
  not NOT_3854(I16138,g9358);
  not NOT_3855(I13106,g7056);
  not NOT_3856(g9361,I16119);
  not NOT_3857(g2007,g1223);
  not NOT_3858(I13605,g7197);
  not NOT_3859(I10448,g5335);
  not NOT_3860(g7463,g7239);
  not NOT_3861(g5009,g4344);
  not NOT_3862(g2407,I6286);
  not NOT_3863(I6163,g402);
  not NOT_3864(I14448,g7792);
  not NOT_3865(g2920,I6652);
  not NOT_3866(g2868,g2223);
  not NOT_3867(I6363,g16);
  not NOT_3868(I15501,g8975);
  not NOT_3869(g9051,I15553);
  not NOT_3870(I15729,g9073);
  not NOT_3871(g2459,I6299);
  not NOT_3872(I15577,g8984);
  not NOT_3873(g4898,g4079);
  not NOT_3874(g6441,I11586);
  not NOT_3875(I13463,g7264);
  not NOT_3876(g9127,I15759);
  not NOT_3877(g2767,I6509);
  not NOT_3878(g4900,I9258);
  not NOT_3879(g1783,I5633);
  not NOT_3880(I7908,g3516);
  not NOT_3881(g5769,I10380);
  not NOT_3882(I11951,g5847);
  not NOT_3883(I11371,g5840);
  not NOT_3884(g8755,g8545);
  not NOT_3885(g636,I5371);
  not NOT_3886(g7279,I13271);
  not NOT_3887(g8226,I14457);
  not NOT_3888(g5836,g5529);
  not NOT_3889(g4510,g2840);
  not NOT_3890(I13234,g6898);
  not NOT_3891(g4245,I8172);
  not NOT_3892(I12427,g6553);
  not NOT_3893(g7720,I14035);
  not NOT_3894(g7118,I12942);
  not NOT_3895(g5918,I10574);
  not NOT_3896(g2793,I6532);
  not NOT_3897(g7367,I13515);
  not NOT_3898(I12632,g6514);
  not NOT_3899(g9103,I15699);
  not NOT_3900(g9303,g9301);
  not NOT_3901(g1676,g727);
  not NOT_3902(g2015,g33);
  not NOT_3903(I8480,g3640);
  not NOT_3904(g6368,I11431);
  not NOT_3905(g7057,g6644);
  not NOT_3906(g8173,I14400);
  not NOT_3907(g4344,g3124);
  not NOT_3908(g6772,I12187);
  not NOT_3909(I6157,g246);
  not NOT_3910(I12403,g6769);
  not NOT_3911(I12547,g6708);
  not NOT_3912(g1828,g769);
  not NOT_3913(g2664,I6463);
  not NOT_3914(g2246,I5989);
  not NOT_3915(g4259,I8196);
  not NOT_3916(g5822,I10491);
  not NOT_3917(g6890,I12541);
  not NOT_3918(g7549,I13831);
  not NOT_3919(g1830,I5718);
  not NOT_3920(g4694,I8977);
  not NOT_3921(I15622,g8999);
  not NOT_3922(g1727,g596);
  not NOT_3923(g3590,I7064);
  not NOT_3924(g3877,g2960);
  not NOT_3925(I10433,g5212);
  not NOT_3926(I5692,g906);
  not NOT_3927(g8602,g8094);
  not NOT_3928(I10387,g5194);
  not NOT_3929(I12226,g6636);
  not NOT_3930(I14433,g8061);
  not NOT_3931(g7686,I13979);
  not NOT_3932(g8407,g8013);
  not NOT_3933(g4088,I7885);
  not NOT_3934(I12481,g6616);
  not NOT_3935(g9072,I15610);
  not NOT_3936(g3657,I7145);
  not NOT_3937(g4923,g4112);
  not NOT_3938(g2721,g1803);
  not NOT_3939(g6505,I11677);
  not NOT_3940(g8868,I15190);
  not NOT_3941(I14148,g7543);
  not NOT_3942(g6011,g5494);
  not NOT_3943(I5960,g187);
  not NOT_3944(g1746,g290);
  not NOT_3945(I14097,g7595);
  not NOT_3946(g6856,I12439);
  not NOT_3947(g4701,I8994);
  not NOT_3948(I10646,g5364);
  not NOT_3949(g8767,g8564);
  not NOT_3950(g9043,I15533);
  not NOT_3951(g3556,I7036);
  not NOT_3952(I13012,g7071);
  not NOT_3953(I10343,g5704);
  not NOT_3954(I14646,g7790);
  not NOT_3955(g3928,g3097);
  not NOT_3956(I16052,g9291);
  not NOT_3957(g8582,g8094);
  not NOT_3958(g9116,I15738);
  not NOT_3959(g6074,g5317);
  not NOT_3960(g3930,g3097);
  not NOT_3961(g2502,I6337);
  not NOT_3962(g9316,g9302);
  not NOT_3963(I11473,g6069);
  not NOT_3964(I13541,g7209);
  not NOT_3965(g4886,g4071);
  not NOT_3966(I10369,g5716);
  not NOT_3967(g9034,I15516);
  not NOT_3968(I12490,g6625);
  not NOT_3969(g8015,g7689);
  not NOT_3970(g2940,I6686);
  not NOT_3971(g8227,I14460);
  not NOT_3972(g4114,I7953);
  not NOT_3973(g7253,g7049);
  not NOT_3974(I11359,g5810);
  not NOT_3975(I12376,g6766);
  not NOT_3976(I12385,g6397);
  not NOT_3977(I13359,g7255);
  not NOT_3978(I9892,g4879);
  not NOT_3979(g5462,g4886);
  not NOT_3980(g2689,g1670);
  not NOT_3981(g6573,g5868);
  not NOT_3982(g6863,I12460);
  not NOT_3983(I11920,g5874);
  not NOT_3984(I12980,g6929);
  not NOT_3985(I7878,g2829);
  not NOT_3986(g8664,I14786);
  not NOT_3987(I8760,g3931);
  not NOT_3988(I11434,g5789);
  not NOT_3989(g3563,g2007);
  not NOT_3990(I10412,g5205);
  not NOT_3991(g2216,I5933);
  not NOT_3992(g6713,I12065);
  not NOT_3993(g1677,g1532);
  not NOT_3994(g7519,I13737);
  not NOT_3995(g7740,I14091);
  not NOT_3996(g4650,I8865);
  not NOT_3997(I7658,g2562);
  not NOT_3998(I5401,g723);
  not NOT_3999(I12888,g6948);
  not NOT_4000(I13828,g7321);
  not NOT_4001(I5676,g911);
  not NOT_4002(I14133,g7574);
  not NOT_4003(g2671,I6468);
  not NOT_4004(g9210,g9200);
  not NOT_4005(g1576,g691);
  not NOT_4006(g6569,I11747);
  not NOT_4007(g1866,g71);
  not NOT_4008(I7882,g2700);
  not NOT_4009(g5788,I10409);
  not NOT_4010(g4008,I7755);
  not NOT_4011(I10896,g5475);
  not NOT_4012(I6894,g1863);
  not NOT_4013(I11344,g5820);
  not NOT_4014(g3844,I7335);
  not NOT_4015(I13344,g7210);
  not NOT_4016(I15484,g8918);
  not NOT_4017(g1848,g772);
  not NOT_4018(I10716,g5537);
  not NOT_4019(I13682,g7251);
  not NOT_4020(g4594,g2941);
  not NOT_4021(g5842,I10541);
  not NOT_4022(g2826,g2183);
  not NOT_4023(g1747,g599);
  not NOT_4024(g1855,g866);
  not NOT_4025(I6075,g2);
  not NOT_4026(g6857,I12442);
  not NOT_4027(g7586,I13903);
  not NOT_4028(I9907,g4837);
  not NOT_4029(I13173,g7089);
  not NOT_4030(g5192,g4841);
  not NOT_4031(I10582,g5437);
  not NOT_4032(g3557,g1773);
  not NOT_4033(g5085,I9457);
  not NOT_4034(g4806,I9139);
  not NOT_4035(I7981,g3555);
  not NOT_4036(I6949,g2148);
  not NOT_4037(I12190,g5918);
  not NOT_4038(g3966,g3160);
  not NOT_4039(I8977,g3877);
  not NOT_4040(g2910,I6636);
  not NOT_4041(g3071,g1948);
  not NOT_4042(g3705,I7204);
  not NOT_4043(g9117,I15741);
  not NOT_4044(I12520,g6622);
  not NOT_4045(g2638,g1582);
  not NOT_4046(g4065,I7838);
  not NOT_4047(g9317,g9306);
  not NOT_4048(I8161,g3517);
  not NOT_4049(g8689,I14857);
  not NOT_4050(g4122,I7973);
  not NOT_4051(I15921,g9206);
  not NOT_4052(g4465,g3677);
  not NOT_4053(g7141,I13009);
  not NOT_4054(I14925,g8381);
  not NOT_4055(g3948,g3131);
  not NOT_4056(g4934,g4125);
  not NOT_4057(g7341,I13441);
  not NOT_4058(g8216,I14427);
  not NOT_4059(I6646,g2246);
  not NOT_4060(g2308,I6081);
  not NOT_4061(I7132,g2554);
  not NOT_4062(I13134,g7017);
  not NOT_4063(I7332,g2947);
  not NOT_4064(I8665,g3051);
  not NOT_4065(I12211,g6502);
  not NOT_4066(I14112,g7560);
  not NOT_4067(g6326,I11305);
  not NOT_4068(g7525,I13755);
  not NOT_4069(g7710,I14009);
  not NOT_4070(g3955,I7658);
  not NOT_4071(I7680,g2712);
  not NOT_4072(I11506,g6189);
  not NOT_4073(I14378,g7691);
  not NOT_4074(g2883,g2237);
  not NOT_4075(I6084,g240);
  not NOT_4076(I7353,g2833);
  not NOT_4077(g8671,I14807);
  not NOT_4078(I11028,g5642);
  not NOT_4079(I13506,g7148);
  not NOT_4080(I12088,g5874);
  not NOT_4081(I6039,g207);
  not NOT_4082(g4033,g3192);
  not NOT_4083(I13028,g7087);
  not NOT_4084(g6760,I12151);
  not NOT_4085(I14603,g7827);
  not NOT_4086(g5520,g4928);
  not NOT_4087(I15184,g8684);
  not NOT_4088(g4096,I7911);
  not NOT_4089(g8564,g7951);
  not NOT_4090(g3038,g2092);
  not NOT_4091(g1818,I5692);
  not NOT_4092(g1577,g695);
  not NOT_4093(g1867,g878);
  not NOT_4094(g9060,I15574);
  not NOT_4095(I9310,g4268);
  not NOT_4096(I7558,g2734);
  not NOT_4097(I10681,g5686);
  not NOT_4098(g5812,I10469);
  not NOT_4099(g6183,I10914);
  not NOT_4100(g7158,I13048);
  not NOT_4101(g2365,I6195);
  not NOT_4102(I12659,g6459);
  not NOT_4103(g6383,I11476);
  not NOT_4104(g7358,I13490);
  not NOT_4105(g5176,I9654);
  not NOT_4106(g4195,I8094);
  not NOT_4107(I9663,g4809);
  not NOT_4108(g6220,I11001);
  not NOT_4109(g7506,I13698);
  not NOT_4110(I15732,g9076);
  not NOT_4111(g4891,g4076);
  not NOT_4112(I13927,g7366);
  not NOT_4113(g4913,g4092);
  not NOT_4114(I12250,g6651);
  not NOT_4115(g658,I5386);
  not NOT_4116(g8910,I15324);
  not NOT_4117(I16100,g9338);
  not NOT_4118(g6779,I12208);
  not NOT_4119(I14857,g8657);
  not NOT_4120(g3769,g2548);
  not NOT_4121(I6952,g1896);
  not NOT_4122(g8638,I14722);
  not NOT_4123(g3836,I7311);
  not NOT_4124(g5829,I10512);
  not NOT_4125(g7587,I13906);
  not NOT_4126(I13649,g7281);
  not NOT_4127(g5286,g4714);
  not NOT_4128(g1975,g1253);
  not NOT_4129(I5747,g1260);
  not NOT_4130(g4807,I9142);
  not NOT_4131(g6977,g6664);
  not NOT_4132(g7111,I12921);
  not NOT_4133(I5855,g71);
  not NOT_4134(I5398,g702);
  not NOT_4135(g3918,I7551);
  not NOT_4136(g2774,g1813);
  not NOT_4137(g7275,I13261);
  not NOT_4138(g7311,I13365);
  not NOT_4139(g3967,I7680);
  not NOT_4140(I6561,g1715);
  not NOT_4141(I11648,g6028);
  not NOT_4142(I10690,g5538);
  not NOT_4143(g6588,g5836);
  not NOT_4144(I11491,g6010);
  not NOT_4145(I11903,g5939);
  not NOT_4146(g9079,I15631);
  not NOT_4147(I13903,g7357);
  not NOT_4148(g8883,I15225);
  not NOT_4149(g6161,I10842);
  not NOT_4150(I7492,g3561);
  not NOT_4151(g6361,I11410);
  not NOT_4152(g4266,I8202);
  not NOT_4153(g2396,g1033);
  not NOT_4154(I7864,g3812);
  not NOT_4155(I10548,g5260);
  not NOT_4156(I13755,g7317);
  not NOT_4157(g5733,I10256);
  not NOT_4158(g7174,g7097);
  not NOT_4159(g6051,g5246);
  not NOT_4160(g3993,g3192);
  not NOT_4161(g8217,I14430);
  not NOT_4162(I13770,g7491);
  not NOT_4163(I11981,g6246);
  not NOT_4164(I9657,g4784);
  not NOT_4165(I12968,g6925);
  not NOT_4166(g1821,g631);
  not NOT_4167(I15329,g8793);
  not NOT_4168(g6327,I11308);
  not NOT_4169(g2780,I6517);
  not NOT_4170(I6764,g1955);
  not NOT_4171(g3822,g1815);
  not NOT_4172(g5610,g4938);
  not NOT_4173(g2509,g37);
  not NOT_4174(I15539,g9005);
  not NOT_4175(g5073,g4477);
  not NOT_4176(g5796,I10427);
  not NOT_4177(I8565,g3071);
  not NOT_4178(g5473,g4903);
  not NOT_4179(g7284,I13284);
  not NOT_4180(g6146,I10801);
  not NOT_4181(g4081,I7870);
  not NOT_4182(g7239,g6945);
  not NOT_4183(g6346,I11365);
  not NOT_4184(g7545,I13819);
  not NOT_4185(I6970,g1872);
  not NOT_4186(g2662,I6457);
  not NOT_4187(g5124,I9520);
  not NOT_4188(g7180,I13092);
  not NOT_4189(g6103,g5317);
  not NOT_4190(g4692,I8971);
  not NOT_4191(g7591,I13918);
  not NOT_4192(g6303,I11236);
  not NOT_4193(g2467,I6305);
  not NOT_4194(I9064,g4302);
  not NOT_4195(I13767,g7486);
  not NOT_4196(I13794,g7346);
  not NOT_4197(I11395,g5812);
  not NOT_4198(g5469,g4898);
  not NOT_4199(g2290,I6054);
  not NOT_4200(I7262,g2514);
  not NOT_4201(I10128,g4688);
  not NOT_4202(g6696,I12022);
  not NOT_4203(g3921,I7558);
  not NOT_4204(I9785,g4747);
  not NOT_4205(I5577,g172);
  not NOT_4206(g4960,g4259);
  not NOT_4207(g7420,I13537);
  not NOT_4208(I11633,g5897);
  not NOT_4209(g5177,I9657);
  not NOT_4210(I12894,g7009);
  not NOT_4211(g7507,I13701);
  not NOT_4212(g8774,I14964);
  not NOT_4213(g5206,g4938);
  not NOT_4214(I7623,g3631);
  not NOT_4215(g2256,g1324);
  not NOT_4216(I11191,g6155);
  not NOT_4217(g2816,g1685);
  not NOT_4218(I13719,g7334);
  not NOT_4219(g6508,I11686);
  not NOT_4220(g6944,I12643);
  not NOT_4221(g3837,I7314);
  not NOT_4222(g6072,g5345);
  not NOT_4223(I11718,g6115);
  not NOT_4224(g3062,g2100);
  not NOT_4225(I14298,g7678);
  not NOT_4226(g9032,I15510);
  not NOT_4227(I5386,g648);
  not NOT_4228(g3462,g1743);
  not NOT_4229(g1756,g533);
  not NOT_4230(g2381,I6245);
  not NOT_4231(I5975,g381);
  not NOT_4232(I11832,g6274);
  not NOT_4233(g8780,g8524);
  not NOT_4234(g9053,I15557);
  not NOT_4235(I12202,g6481);
  not NOT_4236(g4112,I7947);
  not NOT_4237(g7905,I14279);
  not NOT_4238(g4267,I8205);
  not NOT_4239(g2700,g1744);
  not NOT_4240(I7651,g2573);
  not NOT_4241(I16107,g9337);
  not NOT_4242(I8820,g3952);
  not NOT_4243(I11440,g6009);
  not NOT_4244(g2397,g1272);
  not NOT_4245(I12496,g6592);
  not NOT_4246(g5199,g4841);
  not NOT_4247(g1904,g1021);
  not NOT_4248(I12111,g5956);
  not NOT_4249(g6316,I11275);
  not NOT_4250(g7515,I13725);
  not NOT_4251(I11861,g5747);
  not NOT_4252(g8662,I14780);
  not NOT_4253(g5781,I10390);
  not NOT_4254(g4001,g3160);
  not NOT_4255(g6034,I10639);
  not NOT_4256(g8018,I14315);
  not NOT_4257(I13861,g7330);
  not NOT_4258(I9089,g4566);
  not NOT_4259(g8067,I14342);
  not NOT_4260(g2263,g1394);
  not NOT_4261(g7100,I12888);
  not NOT_4262(I13247,g6906);
  not NOT_4263(I6299,g47);
  not NOT_4264(g7300,I13332);
  not NOT_4265(I11389,g5766);
  not NOT_4266(I11926,g6190);
  not NOT_4267(I12986,g6931);
  not NOT_4268(g5797,I10430);
  not NOT_4269(I15414,g8900);
  not NOT_4270(I13045,g6955);
  not NOT_4271(g6147,I10804);
  not NOT_4272(I5984,g540);
  not NOT_4273(g9157,g9141);
  not NOT_4274(g6347,I11368);
  not NOT_4275(I5939,g275);
  not NOT_4276(I13099,g7054);
  not NOT_4277(g3842,I7329);
  not NOT_4278(I13388,g7149);
  not NOT_4279(g8093,I14370);
  not NOT_4280(g6681,I11991);
  not NOT_4281(I11701,g5772);
  not NOT_4282(g8493,g8041);
  not NOT_4283(I13701,g7349);
  not NOT_4284(I10512,g5238);
  not NOT_4285(g3085,g1945);
  not NOT_4286(I8775,g4019);
  not NOT_4287(I7838,g2781);
  not NOT_4288(I8922,g4229);
  not NOT_4289(I11251,g6152);
  not NOT_4290(I11272,g5758);
  not NOT_4291(g7750,I14121);
  not NOT_4292(g3485,g1737);
  not NOT_4293(g2562,g1652);
  not NOT_4294(g1695,g778);
  not NOT_4295(g6697,I12025);
  not NOT_4296(g1637,g1087);
  not NOT_4297(g5144,I9558);
  not NOT_4298(g4592,g2938);
  not NOT_4299(g5344,I9819);
  not NOT_4300(g6210,I10969);
  not NOT_4301(I5636,g891);
  not NOT_4302(g2631,g1586);
  not NOT_4303(g4746,I9076);
  not NOT_4304(I12877,g6700);
  not NOT_4305(g8181,I14420);
  not NOT_4306(g6596,I11800);
  not NOT_4307(g5207,g4673);
  not NOT_4308(g8381,I14603);
  not NOT_4309(g3854,I7365);
  not NOT_4310(g2817,g1849);
  not NOT_4311(g3941,I7626);
  not NOT_4312(I7672,g3062);
  not NOT_4313(I16135,g9357);
  not NOT_4314(g4703,I8998);
  not NOT_4315(g5819,I10482);
  not NOT_4316(g8685,I14851);
  not NOT_4317(g7440,I13577);
  not NOT_4318(I10445,g5418);
  not NOT_4319(I7523,g2562);
  not NOT_4320(I14445,g8067);
  not NOT_4321(I12196,g6471);
  not NOT_4322(I6078,g95);
  not NOT_4323(g2605,g1639);
  not NOT_4324(I13140,g6954);
  not NOT_4325(I9350,g4503);
  not NOT_4326(g7123,I12961);
  not NOT_4327(g8421,g8017);
  not NOT_4328(g5088,I9466);
  not NOT_4329(I8784,g3949);
  not NOT_4330(I13997,g7432);
  not NOT_4331(I8739,g3910);
  not NOT_4332(g1757,g604);
  not NOT_4333(g5488,I9910);
  not NOT_4334(g4932,g4202);
  not NOT_4335(I12526,g6626);
  not NOT_4336(I15759,g9082);
  not NOT_4337(g5701,g5120);
  not NOT_4338(g6820,I12331);
  not NOT_4339(g4624,I8787);
  not NOT_4340(I9009,g4591);
  not NOT_4341(I6959,g1558);
  not NOT_4342(g3520,g1616);
  not NOT_4343(g6936,I12629);
  not NOT_4344(g3219,I6872);
  not NOT_4345(I6517,g1687);
  not NOT_4346(g3640,I7112);
  not NOT_4347(I16049,g9288);
  not NOT_4348(g6117,I10739);
  not NOT_4349(g1811,I5679);
  not NOT_4350(g6317,I11278);
  not NOT_4351(I7551,g2712);
  not NOT_4352(I7104,g2479);
  not NOT_4353(g3812,g1750);
  not NOT_4354(I12457,g6671);
  not NOT_4355(g7528,I13764);
  not NOT_4356(I14722,g8076);
  not NOT_4357(g7151,I13035);
  not NOT_4358(g3958,g3097);
  not NOT_4359(g7351,I13469);
  not NOT_4360(g4677,I8932);
  not NOT_4361(g6601,g6083);
  not NOT_4362(g7530,I13770);
  not NOT_4363(I12866,g6483);
  not NOT_4364(I8190,g3545);
  not NOT_4365(g8562,g8094);
  not NOT_4366(I9918,g4968);
  not NOT_4367(I10271,g5487);
  not NOT_4368(g5114,I9502);
  not NOT_4369(g4576,g2913);
  not NOT_4370(I15940,g9213);
  not NOT_4371(I13447,g7261);
  not NOT_4372(g8631,I14709);
  not NOT_4373(g2673,I6474);
  not NOT_4374(g6775,I12196);
  not NOT_4375(g3829,I7290);
  not NOT_4376(g6922,g6525);
  not NOT_4377(I5763,g1207);
  not NOT_4378(g3911,I7526);
  not NOT_4379(I6214,g7);
  not NOT_4380(g6581,I11773);
  not NOT_4381(g5825,I10500);
  not NOT_4382(I14342,g7582);
  not NOT_4383(g8605,I14680);
  not NOT_4384(I14145,g7542);
  not NOT_4385(I12256,g6647);
  not NOT_4386(I14031,g7448);
  not NOT_4387(g4198,I8101);
  not NOT_4388(I7044,g2402);
  not NOT_4389(g6597,I11803);
  not NOT_4390(g9075,I15619);
  not NOT_4391(I13451,g7262);
  not NOT_4392(I13472,g7266);
  not NOT_4393(I14199,g7704);
  not NOT_4394(I12280,g6684);
  not NOT_4395(g3974,g3131);
  not NOT_4396(I6663,g2246);
  not NOT_4397(I13628,g7248);
  not NOT_4398(g8751,g8545);
  not NOT_4399(g2458,g30);
  not NOT_4400(I5359,g3839);
  not NOT_4401(g6784,I12223);
  not NOT_4402(g2743,g1808);
  not NOT_4403(g3610,g2424);
  not NOT_4404(g2890,g2264);
  not NOT_4405(g5768,I10377);
  not NOT_4406(I10528,g5245);
  not NOT_4407(I16033,g9282);
  not NOT_4408(g8585,g7993);
  not NOT_4409(g1612,I5475);
  not NOT_4410(I10393,g5196);
  not NOT_4411(g7172,g7092);
  not NOT_4412(g1017,I5419);
  not NOT_4413(I7712,g3657);
  not NOT_4414(I14330,g7538);
  not NOT_4415(g2505,g28);
  not NOT_4416(g8041,g7701);
  not NOT_4417(I15962,g9218);
  not NOT_4418(g2011,I5847);
  not NOT_4419(g3124,g1857);
  not NOT_4420(g5806,I10451);
  not NOT_4421(I5416,g8868);
  not NOT_4422(g1935,g1280);
  not NOT_4423(g3980,g3192);
  not NOT_4424(g6937,I12632);
  not NOT_4425(g7143,g6996);
  not NOT_4426(I11591,g5814);
  not NOT_4427(g2734,g2170);
  not NOT_4428(g7343,I13447);
  not NOT_4429(I13776,g7497);
  not NOT_4430(g9039,I15527);
  not NOT_4431(g4524,g2869);
  not NOT_4432(g6294,I11209);
  not NOT_4433(g6840,I12391);
  not NOT_4434(g4644,I8847);
  not NOT_4435(I6590,g2467);
  not NOT_4436(I13147,g7024);
  not NOT_4437(g8673,I14813);
  not NOT_4438(g3540,g2424);
  not NOT_4439(I15833,g9162);
  not NOT_4440(g4119,I7964);
  not NOT_4441(I9837,g4781);
  not NOT_4442(g6190,I10933);
  not NOT_4443(g2074,I5872);
  not NOT_4444(I6657,g1701);
  not NOT_4445(g6390,I11497);
  not NOT_4446(g7134,I12986);
  not NOT_4447(I12885,g6946);
  not NOT_4448(g7334,I13422);
  not NOT_4449(I13825,g7318);
  not NOT_4450(g2992,g1833);
  not NOT_4451(g4258,I8193);
  not NOT_4452(I11858,g6165);
  not NOT_4453(g4577,g2914);
  not NOT_4454(g6501,I11669);
  not NOT_4455(g7548,I13828);
  not NOT_4456(g8669,I14801);
  not NOT_4457(g4867,I9209);
  not NOT_4458(I13858,g7329);
  not NOT_4459(I14709,g8198);
  not NOT_4460(I10259,g5362);
  not NOT_4461(g6156,I10829);
  not NOT_4462(I12511,g6598);
  not NOT_4463(g6356,I11395);
  not NOT_4464(g5433,g5024);
  not NOT_4465(I10708,g5545);
  not NOT_4466(g7555,I13843);
  not NOT_4467(g1800,g1477);
  not NOT_4468(I12763,g6686);
  not NOT_4469(g3287,I6911);
  not NOT_4470(g8772,g8585);
  not NOT_4471(I7885,g2837);
  not NOT_4472(I5654,g921);
  not NOT_4473(I8357,g1182);
  not NOT_4474(I6930,g1876);
  not NOT_4475(g2573,g1649);
  not NOT_4476(g2863,g1778);
  not NOT_4477(g7792,I14231);
  not NOT_4478(g2480,g44);
  not NOT_4479(I15613,g8996);
  not NOT_4480(I9788,g4711);
  not NOT_4481(g8743,g8524);
  not NOT_4482(g3849,I7350);
  not NOT_4483(g6704,I12044);
  not NOT_4484(I15947,g9221);
  not NOT_4485(g5845,I10548);
  not NOT_4486(g4599,I8712);
  not NOT_4487(g5137,I9539);
  not NOT_4488(g5395,I9840);
  not NOT_4489(g8856,I15160);
  not NOT_4490(g7113,I12927);
  not NOT_4491(g3898,g3160);
  not NOT_4492(g8734,I14904);
  not NOT_4493(g4026,g3192);
  not NOT_4494(g7313,I13369);
  not NOT_4495(g4274,I8218);
  not NOT_4496(g4426,I8428);
  not NOT_4497(I7036,g2454);
  not NOT_4498(g6250,g5679);
  not NOT_4499(g6810,I12301);
  not NOT_4500(g4614,I8757);
  not NOT_4501(g6363,I11416);
  not NOT_4502(g4370,I8351);
  not NOT_4503(I5978,g414);
  not NOT_4504(g3510,g2185);
  not NOT_4505(I10810,g5403);
  not NOT_4506(g6032,g5494);
  not NOT_4507(I11446,g6062);
  not NOT_4508(g4125,I7978);
  not NOT_4509(I14810,g8481);
  not NOT_4510(I11227,g6130);
  not NOT_4511(g6432,I11569);
  not NOT_4512(g5807,I10454);
  not NOT_4513(I14657,g7782);
  not NOT_4514(g7094,g6525);
  not NOT_4515(I12307,g6712);
  not NOT_4516(I11025,g5638);
  not NOT_4517(I12085,g5971);
  not NOT_4518(g2976,I6728);
  not NOT_4519(I7335,g2910);
  not NOT_4520(g1823,g768);
  not NOT_4521(g7494,g7260);
  not NOT_4522(g7518,I13734);
  not NOT_4523(g5266,I9782);
  not NOT_4524(g6568,I11744);
  not NOT_4525(g4544,g2886);
  not NOT_4526(I11203,g6129);
  not NOT_4527(I5542,g1272);
  not NOT_4528(I13203,g7088);
  not NOT_4529(g7776,I14199);
  not NOT_4530(g1649,g1217);
  not NOT_4531(I7749,g3692);
  not NOT_4532(g7593,I13924);
  not NOT_4533(g3819,g1748);
  not NOT_4534(g4636,I8823);
  not NOT_4535(g3694,g2174);
  not NOT_4536(g2326,I6121);
  not NOT_4537(I14792,g8583);
  not NOT_4538(I9520,g3995);
  not NOT_4539(g6357,I11398);
  not NOT_4540(g4106,I7931);
  not NOT_4541(I15507,g8968);
  not NOT_4542(I12942,g7023);
  not NOT_4543(g3852,I7359);
  not NOT_4544(I6471,g1923);
  not NOT_4545(g3923,I7564);
  not NOT_4546(g4306,I8273);
  not NOT_4547(I8778,g3922);
  not NOT_4548(I11281,g5785);
  not NOT_4549(I12268,g6661);
  not NOT_4550(g9320,g9307);
  not NOT_4551(g5481,g4914);
  not NOT_4552(g3488,g1727);
  not NOT_4553(I7947,g3485);
  not NOT_4554(I13281,g7155);
  not NOT_4555(g1698,I5542);
  not NOT_4556(I6242,g1554);
  not NOT_4557(I16173,g9382);
  not NOT_4558(I12655,g6458);
  not NOT_4559(I11377,g5811);
  not NOT_4560(g7264,I13234);
  not NOT_4561(g5726,I10243);
  not NOT_4562(g5154,I9588);
  not NOT_4563(I10919,g5479);
  not NOT_4564(I9005,g4585);
  not NOT_4565(g7160,I13054);
  not NOT_4566(g7360,I13496);
  not NOT_4567(I11562,g5939);
  not NOT_4568(I11645,g5874);
  not NOT_4569(I13562,g7179);
  not NOT_4570(g7521,I13743);
  not NOT_4571(g4622,I8781);
  not NOT_4572(g4027,g2845);
  not NOT_4573(g2183,I5908);
  not NOT_4574(g3951,I7648);
  not NOT_4575(g7050,g6618);
  not NOT_4576(I6254,g536);
  not NOT_4577(g2383,I6251);
  not NOT_4578(g2924,g2314);
  not NOT_4579(I12839,g6630);
  not NOT_4580(I12930,g7019);
  not NOT_4581(I8949,g4116);
  not NOT_4582(I7632,g3634);
  not NOT_4583(I7095,g2539);
  not NOT_4584(I12993,g6933);
  not NOT_4585(I10545,g5259);
  not NOT_4586(g6626,I11870);
  not NOT_4587(I11290,g5818);
  not NOT_4588(I13290,g7158);
  not NOT_4589(I7495,g3562);
  not NOT_4590(I14079,g7579);
  not NOT_4591(g4904,g4085);
  not NOT_4592(g4200,I8105);
  not NOT_4593(I13698,g7348);
  not NOT_4594(I7302,g2825);
  not NOT_4595(I12965,g6924);
  not NOT_4596(I12131,g5918);
  not NOT_4597(g9299,I16023);
  not NOT_4598(I6009,g359);
  not NOT_4599(g3870,g3466);
  not NOT_4600(I8998,g4576);
  not NOT_4601(I5512,g557);
  not NOT_4602(g4003,g3192);
  not NOT_4603(I9974,g4676);
  not NOT_4604(g5112,I9496);
  not NOT_4605(g3825,g1826);
  not NOT_4606(g3650,I7126);
  not NOT_4607(g5267,I9785);
  not NOT_4608(I12487,g6623);
  not NOT_4609(g4841,g4250);
  not NOT_4610(g2161,g1454);
  not NOT_4611(I8084,g3706);
  not NOT_4612(g1652,g1220);
  not NOT_4613(g2361,I6183);
  not NOT_4614(I7752,g3591);
  not NOT_4615(I12502,g6604);
  not NOT_4616(g4191,I8084);
  not NOT_4617(g1843,g771);
  not NOT_4618(g8760,g8545);
  not NOT_4619(g3008,g1816);
  not NOT_4620(I8850,g4031);
  not NOT_4621(g2665,g1661);
  not NOT_4622(g7289,I13299);
  not NOT_4623(g7777,I14202);
  not NOT_4624(g6683,g6237);
  not NOT_4625(g5401,I9845);
  not NOT_4626(I10125,g5127);
  not NOT_4627(g4695,I8980);
  not NOT_4628(I10532,g5253);
  not NOT_4629(g4637,I8826);
  not NOT_4630(I5649,g1389);
  not NOT_4631(g7835,I14257);
  not NOT_4632(g2327,I6124);
  not NOT_4633(g5129,I9531);
  not NOT_4634(g6778,I12205);
  not NOT_4635(g5761,I10356);
  not NOT_4636(g3768,g2253);
  not NOT_4637(I10783,g5542);
  not NOT_4638(g6894,g6525);
  not NOT_4639(I13403,g7269);
  not NOT_4640(I13547,g1170);
  not NOT_4641(g4307,g3700);
  not NOT_4642(g4536,g2877);
  not NOT_4643(g2999,g1823);
  not NOT_4644(I14783,g8324);
  not NOT_4645(g3972,I7691);
  not NOT_4646(g1686,I5531);
  not NOT_4647(g5828,I10509);
  not NOT_4648(g2346,I6154);
  not NOT_4649(g2633,g1577);
  not NOT_4650(I12469,g6586);
  not NOT_4651(g9244,I15974);
  not NOT_4652(I10561,g5265);
  not NOT_4653(I6229,g486);
  not NOT_4654(g8608,I14687);
  not NOT_4655(g8220,I14439);
  not NOT_4656(I10353,g5710);
  not NOT_4657(I12286,g6696);
  not NOT_4658(g6782,I12217);
  not NOT_4659(I7164,g2157);
  not NOT_4660(I10295,g5523);
  not NOT_4661(I8919,g4196);
  not NOT_4662(g3943,I7632);
  not NOT_4663(g9140,I15784);
  not NOT_4664(I9177,g4299);
  not NOT_4665(g9078,I15628);
  not NOT_4666(g9340,I16090);
  not NOT_4667(I13481,g7254);
  not NOT_4668(g5592,g4969);
  not NOT_4669(I14680,g7810);
  not NOT_4670(g6661,I11961);
  not NOT_4671(g6075,g5345);
  not NOT_4672(g4016,g3192);
  not NOT_4673(I8952,g4197);
  not NOT_4674(g699,I5395);
  not NOT_4675(I12038,g5847);
  not NOT_4676(g5746,I10295);
  not NOT_4677(g6475,I11633);
  not NOT_4678(g9035,I15519);
  not NOT_4679(g1670,g1489);
  not NOT_4680(g3465,I6963);
  not NOT_4681(g8977,I15433);
  not NOT_4682(I7296,g2915);
  not NOT_4683(g3934,I7599);
  not NOT_4684(g9082,I15638);
  not NOT_4685(g3230,I6887);
  not NOT_4686(g4522,g2867);
  not NOT_4687(g4115,I7956);
  not NOT_4688(g4251,I8180);
  not NOT_4689(g6292,I11203);
  not NOT_4690(I12187,g5897);
  not NOT_4691(g4811,I9158);
  not NOT_4692(g4642,I8841);
  not NOT_4693(g7541,I13807);
  not NOT_4694(g2944,g2363);
  not NOT_4695(g2240,I5981);
  not NOT_4696(g1938,g1288);
  not NOT_4697(g1813,g620);
  not NOT_4698(g6646,I11920);
  not NOT_4699(g7132,I12980);
  not NOT_4700(I8986,g4552);
  not NOT_4701(g8665,I14789);
  not NOT_4702(g7332,I13416);
  not NOT_4703(I13490,g7130);
  not NOT_4704(g1909,g998);
  not NOT_4705(g7353,I13475);
  not NOT_4706(g6603,I11815);
  not NOT_4707(g3096,I6834);
  not NOT_4708(I5872,g77);
  not NOT_4709(I13956,g7499);
  not NOT_4710(g5468,I9884);
  not NOT_4711(g6850,I12421);
  not NOT_4712(g3496,I6974);
  not NOT_4713(g7744,I14103);
  not NOT_4714(g4654,I8877);
  not NOT_4715(I13103,g7055);
  not NOT_4716(g3845,I7338);
  not NOT_4717(g2316,I6109);
  not NOT_4718(g9214,I15918);
  not NOT_4719(I5989,g1460);
  not NOT_4720(I7389,g3496);
  not NOT_4721(I11824,g6283);
  not NOT_4722(g5677,I10166);
  not NOT_4723(I7706,g2584);
  not NOT_4724(I13888,g7335);
  not NOT_4725(g3891,g3097);
  not NOT_4726(I8925,g4482);
  not NOT_4727(g3913,g2834);
  not NOT_4728(I10289,g5569);
  not NOT_4729(g9110,I15720);
  not NOT_4730(g9310,I16046);
  not NOT_4731(g6702,I12038);
  not NOT_4732(g7558,I13850);
  not NOT_4733(I7888,g3505);
  not NOT_4734(g4595,g2942);
  not NOT_4735(g4537,g2878);
  not NOT_4736(I15927,g9208);
  not NOT_4737(I7029,g2392);
  not NOT_4738(g1687,g10);
  not NOT_4739(I7371,g3050);
  not NOT_4740(g2347,I6157);
  not NOT_4741(I12666,g6476);
  not NOT_4742(g5149,I9573);
  not NOT_4743(I14288,g7705);
  not NOT_4744(I14224,g7722);
  not NOT_4745(I9344,g4341);
  not NOT_4746(I12217,g6631);
  not NOT_4747(I7956,g2810);
  not NOT_4748(g1586,g730);
  not NOT_4749(I6788,g1681);
  not NOT_4750(I12478,g6603);
  not NOT_4751(g2533,g1336);
  not NOT_4752(g8753,I14925);
  not NOT_4753(g3859,I7380);
  not NOT_4754(g4612,I8751);
  not NOT_4755(g7511,I13713);
  not NOT_4756(g4017,g2845);
  not NOT_4757(I15648,g9044);
  not NOT_4758(g2914,g2308);
  not NOT_4759(I8277,g3504);
  not NOT_4760(g5198,g4969);
  not NOT_4761(I9819,g4691);
  not NOT_4762(g8072,I14349);
  not NOT_4763(g9236,I15962);
  not NOT_4764(g2210,g1326);
  not NOT_4765(g6616,I11848);
  not NOT_4766(g4935,g4202);
  not NOT_4767(g7092,I12866);
  not NOT_4768(I5670,g941);
  not NOT_4769(I15604,g8993);
  not NOT_4770(g7492,I13656);
  not NOT_4771(I14816,g8642);
  not NOT_4772(g1570,g665);
  not NOT_4773(g1860,g162);
  not NOT_4774(g8443,g8015);
  not NOT_4775(I6192,g327);
  not NOT_4776(g7574,I13869);
  not NOT_4777(g6004,g5494);
  not NOT_4778(I15770,g9121);
  not NOT_4779(I10687,g5674);
  not NOT_4780(g4629,I8802);
  not NOT_4781(I10976,g5726);
  not NOT_4782(g6404,I11525);
  not NOT_4783(I12223,g6655);
  not NOT_4784(g4328,g3086);
  not NOT_4785(I14687,g7826);
  not NOT_4786(g7714,I14019);
  not NOT_4787(g6647,I11923);
  not NOT_4788(g4130,I7987);
  not NOT_4789(g4542,g2884);
  not NOT_4790(I10752,g5618);
  not NOT_4791(g3815,g1822);
  not NOT_4792(I7338,g2923);
  not NOT_4793(g6764,I12161);
  not NOT_4794(I14374,g7693);
  not NOT_4795(I10643,g5267);
  not NOT_4796(g3692,I7198);
  not NOT_4797(I13088,g7045);
  not NOT_4798(g9222,I15940);
  not NOT_4799(I14643,g7837);
  not NOT_4800(g2936,I6680);
  not NOT_4801(g3497,g2185);
  not NOT_4802(g5524,I9938);
  not NOT_4803(g7580,I13885);
  not NOT_4804(g4800,I9123);
  not NOT_4805(g5644,g4748);
  not NOT_4806(I15845,g9174);
  not NOT_4807(g3960,I7667);
  not NOT_4808(I8892,g4115);
  not NOT_4809(g1879,I5763);
  not NOT_4810(g4554,g2892);
  not NOT_4811(I11497,g6014);
  not NOT_4812(g9064,I15586);
  not NOT_4813(I15990,g9239);
  not NOT_4814(I5552,g1284);
  not NOT_4815(g7262,I13228);
  not NOT_4816(g5152,I9582);
  not NOT_4817(g5258,I9774);
  not NOT_4818(I14260,g7717);
  not NOT_4819(g7736,I14079);
  not NOT_4820(g5818,I10479);
  not NOT_4821(I10842,g5701);
  not NOT_4822(g6224,I11011);
  not NOT_4823(g5577,I10046);
  not NOT_4824(I14668,g7787);
  not NOT_4825(I11659,g5897);
  not NOT_4826(g5717,g4969);
  not NOT_4827(I13126,g6949);
  not NOT_4828(I13659,g7232);
  not NOT_4829(I8945,g4106);
  not NOT_4830(I11987,g6278);
  not NOT_4831(g6320,I11287);
  not NOT_4832(I12373,g6763);
  not NOT_4833(I6431,g1825);
  not NOT_4834(I13250,g7036);
  not NOT_4835(I14489,g7829);
  not NOT_4836(g2922,g2313);
  not NOT_4837(g1587,g734);
  not NOT_4838(g3783,I7255);
  not NOT_4839(g8013,g7561);
  not NOT_4840(I10525,g5244);
  not NOT_4841(I10488,g5230);
  not NOT_4842(I16061,g9294);
  not NOT_4843(I10424,g5209);
  not NOT_4844(g7476,g7229);
  not NOT_4845(I8709,g4191);
  not NOT_4846(g3979,I7702);
  not NOT_4847(I14424,g7652);
  not NOT_4848(I6376,g38);
  not NOT_4849(g5186,I9684);
  not NOT_4850(I10558,g5264);
  not NOT_4851(I8140,g3429);
  not NOT_4852(I12936,g7015);
  not NOT_4853(g9237,I15965);
  not NOT_4854(I9136,g4280);
  not NOT_4855(I11296,g5831);
  not NOT_4856(I9336,g4493);
  not NOT_4857(g6617,I11851);
  not NOT_4858(g6789,I12238);
  not NOT_4859(I13296,g7161);
  not NOT_4860(g4512,g2842);
  not NOT_4861(g2460,I6302);
  not NOT_4862(I7098,g2477);
  not NOT_4863(I8907,g4095);
  not NOT_4864(I11338,g5798);
  not NOT_4865(g7722,I14039);
  not NOT_4866(I12334,g6713);
  not NOT_4867(I13338,g7190);
  not NOT_4868(I9594,g4718);
  not NOT_4869(I7498,g2752);
  not NOT_4870(g5026,I9366);
  not NOT_4871(I6286,g1307);
  not NOT_4872(g3676,g2380);
  not NOT_4873(g9194,g9182);
  not NOT_4874(g5426,g5013);
  not NOT_4875(I6911,g1869);
  not NOT_4876(I8517,g3014);
  not NOT_4877(g7285,I13287);
  not NOT_4878(g2784,g2340);
  not NOT_4879(g5170,I9636);
  not NOT_4880(g3761,g1772);
  not NOT_4881(g4056,g3082);
  not NOT_4882(g7500,I13676);
  not NOT_4883(I11060,g5453);
  not NOT_4884(g9089,I15657);
  not NOT_4885(I13060,g6959);
  not NOT_4886(g6299,I11224);
  not NOT_4887(g5821,I10488);
  not NOT_4888(I11197,g6122);
  not NOT_4889(g3828,I7287);
  not NOT_4890(g4649,I8862);
  not NOT_4891(I7584,g3062);
  not NOT_4892(I11855,g5751);
  not NOT_4893(I6733,g1718);
  not NOT_4894(g3830,I7293);
  not NOT_4895(I6974,g2528);
  not NOT_4896(I15388,g8898);
  not NOT_4897(I15324,g8779);
  not NOT_4898(I6270,g492);
  not NOT_4899(g2937,g2346);
  not NOT_4900(I11870,g5752);
  not NOT_4901(g7139,I12999);
  not NOT_4902(g9071,I15607);
  not NOT_4903(g5939,I10579);
  not NOT_4904(I10705,g5463);
  not NOT_4905(g6892,I12547);
  not NOT_4906(g1832,g763);
  not NOT_4907(g2479,g32);
  not NOT_4908(g7339,I13435);
  not NOT_4909(I13527,g7217);
  not NOT_4910(g2668,g1662);
  not NOT_4911(I14042,g7470);
  not NOT_4912(g1853,g766);
  not NOT_4913(g2840,g2207);
  not NOT_4914(g4698,I8989);
  not NOT_4915(g8775,g8564);
  not NOT_4916(g3746,g2100);
  not NOT_4917(g5083,g4457);
  not NOT_4918(g7838,I14264);
  not NOT_4919(I5879,g1267);
  not NOT_4920(g7024,I12782);
  not NOT_4921(g7424,I13547);
  not NOT_4922(I7362,g2933);
  not NOT_4923(I12909,g7046);
  not NOT_4924(I14270,g7703);
  not NOT_4925(g7737,I14082);
  not NOT_4926(I10678,g5566);
  not NOT_4927(I6124,g399);
  not NOT_4928(g8581,g8094);
  not NOT_4929(I14124,g7591);
  not NOT_4930(g6945,I12646);
  not NOT_4931(I12117,g5918);
  not NOT_4932(g1794,I5646);
  not NOT_4933(I11503,g6220);
  not NOT_4934(g2501,g27);
  not NOT_4935(I11867,g6286);
  not NOT_4936(I11894,g5956);
  not NOT_4937(I10460,g5219);
  not NOT_4938(I13894,g7353);
  not NOT_4939(g4463,I8483);
  not NOT_4940(I14460,g7789);
  not NOT_4941(g6244,g5670);
  not NOT_4942(g7077,g6676);
  not NOT_4943(I9496,g3971);
  not NOT_4944(g7231,I13173);
  not NOT_4945(g3932,I7595);
  not NOT_4946(g5790,I10415);
  not NOT_4947(g7523,I13749);
  not NOT_4948(I9845,g4728);
  not NOT_4949(g6140,I10783);
  not NOT_4950(g3953,g3160);
  not NOT_4951(g6340,I11347);
  not NOT_4952(I11714,g5772);
  not NOT_4953(g9350,I16100);
  not NOT_4954(g5187,I9687);
  not NOT_4955(g5061,I9425);
  not NOT_4956(I14267,g7695);
  not NOT_4957(I14294,g7553);
  not NOT_4958(g6478,I11638);
  not NOT_4959(g8784,g8545);
  not NOT_4960(g2942,g2350);
  not NOT_4961(g5461,g4885);
  not NOT_4962(g4279,g3340);
  not NOT_4963(I11707,g5988);
  not NOT_4964(g7205,I13131);
  not NOT_4965(I13707,g7420);
  not NOT_4966(I13819,g7426);
  not NOT_4967(g5756,I10343);
  not NOT_4968(g6035,g5494);
  not NOT_4969(g6959,I12678);
  not NOT_4970(I7728,g3675);
  not NOT_4971(I11257,g5805);
  not NOT_4972(g5622,g4938);
  not NOT_4973(g4619,I8772);
  not NOT_4974(g5027,I9369);
  not NOT_4975(g6517,I11701);
  not NOT_4976(I11818,g6276);
  not NOT_4977(g3677,g2485);
  not NOT_4978(g5427,g5115);
  not NOT_4979(I15871,g9184);
  not NOT_4980(I11055,g5696);
  not NOT_4981(I13979,g7415);
  not NOT_4982(I5374,g634);
  not NOT_4983(I13496,g7133);
  not NOT_4984(g7742,I14097);
  not NOT_4985(g4652,I8871);
  not NOT_4986(g7551,I13837);
  not NOT_4987(g7104,I12900);
  not NOT_4988(g6876,I12499);
  not NOT_4989(g7099,I12885);
  not NOT_4990(g4057,I7832);
  not NOT_4991(g7304,I13344);
  not NOT_4992(g8668,I14798);
  not NOT_4993(I11978,g6186);
  not NOT_4994(I6849,g368);
  not NOT_4995(g3866,g2945);
  not NOT_4996(g2954,g2374);
  not NOT_4997(g4457,I8477);
  not NOT_4998(g7499,g7258);
  not NOT_4999(I8877,g4274);
  not NOT_5000(g2810,g1922);
  not NOT_5001(g2363,I6189);
  not NOT_5002(g6656,I11948);
  not NOT_5003(g9212,I15912);
  not NOT_5004(I12639,g6506);
  not NOT_5005(I16151,g9369);
  not NOT_5006(g3716,g2522);
  not NOT_5007(g5514,g4922);
  not NOT_5008(I5545,g1276);
  not NOT_5009(g5403,g5088);
  not NOT_5010(g5145,I9561);
  not NOT_5011(g2453,I6291);
  not NOT_5012(I5380,g645);
  not NOT_5013(g5841,I10538);
  not NOT_5014(g3848,I7347);
  not NOT_5015(g1750,g602);
  not NOT_5016(I6900,g1866);
  not NOT_5017(I12265,g6660);
  not NOT_5018(g7754,I14133);
  not NOT_5019(I10160,g5139);
  not NOT_5020(g5763,I10366);
  not NOT_5021(I9142,g4236);
  not NOT_5022(g5191,g4969);
  not NOT_5023(g8156,I14394);
  not NOT_5024(g3855,I7368);
  not NOT_5025(I14160,g7549);
  not NOT_5026(g3398,I6952);
  not NOT_5027(I8928,g4153);
  not NOT_5028(g7273,I13255);
  not NOT_5029(I6245,g142);
  not NOT_5030(I9081,g4357);
  not NOT_5031(I12391,g6744);
  not NOT_5032(g4598,I8709);
  not NOT_5033(g6110,g5335);
  not NOT_5034(g6310,I11257);
  not NOT_5035(I6291,g46);
  not NOT_5036(g7044,g6543);
  not NOT_5037(I10617,g5677);
  not NOT_5038(I15628,g9001);
  not NOT_5039(g4121,I7970);
  not NOT_5040(I5559,g1292);
  not NOT_5041(g2157,I5897);
  not NOT_5042(g7269,I13247);
  not NOT_5043(g6663,I11967);
  not NOT_5044(g4670,I8925);
  not NOT_5045(g5159,I9603);
  not NOT_5046(g4625,I8790);
  not NOT_5047(g7983,I14294);
  not NOT_5048(I10277,g5472);
  not NOT_5049(I11018,g5626);
  not NOT_5050(I13196,g7008);
  not NOT_5051(I7635,g3052);
  not NOT_5052(I13695,g7345);
  not NOT_5053(g6824,I12343);
  not NOT_5054(g7712,I14015);
  not NOT_5055(g1666,g1472);
  not NOT_5056(g3524,g2306);
  not NOT_5057(g4253,g2734);
  not NOT_5058(g2929,g2327);
  not NOT_5059(g4938,I9310);
  not NOT_5060(g6236,I11037);
  not NOT_5061(g4813,I9162);
  not NOT_5062(I12586,g6643);
  not NOT_5063(g7543,I13813);
  not NOT_5064(g5016,I9350);
  not NOT_5065(g5757,g5261);
  not NOT_5066(g8810,I15068);
  not NOT_5067(g3644,g2131);
  not NOT_5068(I7305,g3048);
  not NOT_5069(g8363,g7992);
  not NOT_5070(I15776,g9127);
  not NOT_5071(I16058,g9294);
  not NOT_5072(I10494,g5232);
  not NOT_5073(g4909,I9271);
  not NOT_5074(I12442,g6542);
  not NOT_5075(I5515,g567);
  not NOT_5076(I14623,g7833);
  not NOT_5077(I8844,g3992);
  not NOT_5078(g5522,g4930);
  not NOT_5079(g5115,I9505);
  not NOT_5080(g6877,I12502);
  not NOT_5081(g5811,I10466);
  not NOT_5082(g5642,I10125);
  not NOT_5083(g2626,g1571);
  not NOT_5084(g3577,g2372);
  not NOT_5085(g7534,I13782);
  not NOT_5086(g7729,I14058);
  not NOT_5087(g3867,g2946);
  not NOT_5088(I15950,g9222);
  not NOT_5089(I13457,g7120);
  not NOT_5090(g1655,g1231);
  not NOT_5091(g6657,I11951);
  not NOT_5092(I7755,g3019);
  not NOT_5093(g4552,g2890);
  not NOT_5094(g9062,I15580);
  not NOT_5095(I11917,g5897);
  not NOT_5096(g4606,I8733);
  not NOT_5097(g6556,I11732);
  not NOT_5098(I10418,g5453);
  not NOT_5099(g6222,g5654);
  not NOT_5100(I12041,g5897);
  not NOT_5101(g5874,I10565);
  not NOT_5102(I9001,g4577);
  not NOT_5103(I14822,g8649);
  not NOT_5104(g7014,I12760);
  not NOT_5105(g4687,I8962);
  not NOT_5106(I8966,g4444);
  not NOT_5107(I12430,g6432);
  not NOT_5108(I11001,g5698);
  not NOT_5109(g5654,g4748);
  not NOT_5110(I12493,g6587);
  not NOT_5111(g7414,I13527);
  not NOT_5112(I9129,g4475);
  not NOT_5113(I15394,g8916);
  not NOT_5114(g3975,g3131);
  not NOT_5115(g6064,I10681);
  not NOT_5116(g4586,g2926);
  not NOT_5117(g6899,g6525);
  not NOT_5118(g2683,g1666);
  not NOT_5119(g6785,I12226);
  not NOT_5120(I11689,g5956);
  not NOT_5121(I11923,g5939);
  not NOT_5122(I12340,g6725);
  not NOT_5123(I12983,g6930);
  not NOT_5124(g7513,I13719);
  not NOT_5125(I5969,g303);
  not NOT_5126(I12806,g6602);
  not NOT_5127(I12684,g6472);
  not NOT_5128(I7602,g2562);
  not NOT_5129(g2894,g2267);
  not NOT_5130(I15420,g8881);
  not NOT_5131(g4570,g2907);
  not NOT_5132(g4341,I8308);
  not NOT_5133(g9298,I16020);
  not NOT_5134(g9085,I15645);
  not NOT_5135(I8814,g4028);
  not NOT_5136(g1667,g1481);
  not NOT_5137(g4525,g2870);
  not NOT_5138(g4710,I9009);
  not NOT_5139(g7178,I13088);
  not NOT_5140(g2782,g1616);
  not NOT_5141(g6295,I11212);
  not NOT_5142(g1235,I5422);
  not NOT_5143(g5612,g4814);
  not NOT_5144(I12517,g6613);
  not NOT_5145(g6237,I11040);
  not NOT_5146(g4645,I8850);
  not NOT_5147(I13157,g6997);
  not NOT_5148(g2661,I6454);
  not NOT_5149(g5417,g5006);
  not NOT_5150(g1566,g652);
  not NOT_5151(g7135,I12989);
  not NOT_5152(g6844,I12403);
  not NOT_5153(g7335,I13425);
  not NOT_5154(I11066,g5460);
  not NOT_5155(I13066,g6957);
  not NOT_5156(I13231,g6897);
  not NOT_5157(g7288,I13296);
  not NOT_5158(g6194,I10937);
  not NOT_5159(I5528,g43);
  not NOT_5160(g2627,g1572);
  not NOT_5161(I14118,g7565);
  not NOT_5162(g5128,I9528);
  not NOT_5163(I9624,g4746);
  not NOT_5164(g2292,I6060);
  not NOT_5165(I14022,g7443);
  not NOT_5166(g6089,g5317);
  not NOT_5167(I12193,g6468);
  not NOT_5168(g6731,I12101);
  not NOT_5169(g4607,I8736);
  not NOT_5170(I8769,g3999);
  not NOT_5171(I13876,g7347);
  not NOT_5172(I13885,g7351);
  not NOT_5173(g5542,g5061);
  not NOT_5174(g7022,I12776);
  not NOT_5175(g2646,I6422);
  not NOT_5176(g7422,I13541);
  not NOT_5177(g4659,I8892);
  not NOT_5178(g7749,I14118);
  not NOT_5179(g1555,I5428);
  not NOT_5180(I12523,g6624);
  not NOT_5181(g4358,g3680);
  not NOT_5182(g1804,I5664);
  not NOT_5183(I6887,g2528);
  not NOT_5184(g8683,g8235);
  not NOT_5185(I13854,g7327);
  not NOT_5186(g6071,I10694);
  not NOT_5187(g9219,I15933);
  not NOT_5188(g1792,g616);
  not NOT_5189(g2039,g1228);
  not NOT_5190(g3061,I6795);
  not NOT_5191(g3187,I6860);
  not NOT_5192(g6471,I11627);
  not NOT_5193(g8778,I14974);
  not NOT_5194(I14276,g7720);
  not NOT_5195(I14285,g7625);
  not NOT_5196(g2484,g45);
  not NOT_5197(g9031,I15507);
  not NOT_5198(g5800,I10439);
  not NOT_5199(I5410,g8866);
  not NOT_5200(g3461,I6959);
  not NOT_5201(g6242,I11047);
  not NOT_5202(I14305,g7537);
  not NOT_5203(g9252,I15982);
  not NOT_5204(g4587,g2928);
  not NOT_5205(I12475,g6596);
  not NOT_5206(I6033,g3);
  not NOT_5207(I9576,g4706);
  not NOT_5208(I10466,g5221);
  not NOT_5209(g6948,I12655);
  not NOT_5210(g4111,I7944);
  not NOT_5211(I5839,g1198);
  not NOT_5212(g7560,I13854);
  not NOT_5213(g4275,g3790);
  not NOT_5214(g4311,I8282);
  not NOT_5215(g9376,I16154);
  not NOT_5216(I15738,g9079);
  not NOT_5217(I15562,g8979);
  not NOT_5218(I15645,g9043);
  not NOT_5219(g6955,I12666);
  not NOT_5220(g4615,I8760);
  not NOT_5221(g3904,g3160);
  not NOT_5222(g8661,I14777);
  not NOT_5223(I10177,g4721);
  not NOT_5224(I15699,g9061);
  not NOT_5225(I6096,g521);
  not NOT_5226(g6254,g5683);
  not NOT_5227(g6814,I12313);
  not NOT_5228(g7095,I12877);
  not NOT_5229(g3514,g2424);
  not NOT_5230(g2919,g2311);
  not NOT_5231(g7037,g6525);
  not NOT_5232(g6150,g5287);
  not NOT_5233(g7495,I13663);
  not NOT_5234(g1908,g812);
  not NOT_5235(g7437,I13570);
  not NOT_5236(g6350,I11377);
  not NOT_5237(g7102,I12894);
  not NOT_5238(g7208,I13140);
  not NOT_5239(I6195,g405);
  not NOT_5240(g7302,I13338);
  not NOT_5241(I13550,g1173);
  not NOT_5242(g6038,I10649);
  not NOT_5243(I5667,g916);
  not NOT_5244(I11314,g5781);
  not NOT_5245(I6337,g1348);
  not NOT_5246(g3841,I7326);
  not NOT_5247(I13314,g7160);
  not NOT_5248(I11287,g5806);
  not NOT_5249(g2276,I6029);
  not NOT_5250(I12253,g6427);
  not NOT_5251(g6773,I12190);
  not NOT_5252(I13287,g7157);
  not NOT_5253(g1567,g655);
  not NOT_5254(I16103,g9339);
  not NOT_5255(g7579,I13882);
  not NOT_5256(I14064,g7556);
  not NOT_5257(g6009,I10605);
  not NOT_5258(g3191,I6868);
  not NOT_5259(g4545,g2887);
  not NOT_5260(g2616,g1564);
  not NOT_5261(g7719,g7475);
  not NOT_5262(g2561,g1555);
  not NOT_5263(g5490,g4917);
  not NOT_5264(g691,I5389);
  not NOT_5265(g5823,I10494);
  not NOT_5266(g534,I5365);
  not NOT_5267(g5166,I9624);
  not NOT_5268(I11596,g6228);
  not NOT_5269(g4591,g2937);
  not NOT_5270(g8603,I14674);
  not NOT_5271(I13054,g6960);
  not NOT_5272(g8039,g7696);
  not NOT_5273(g1776,g608);
  not NOT_5274(g6769,I12176);
  not NOT_5275(g7752,I14127);
  not NOT_5276(I11431,g5782);
  not NOT_5277(g9073,I15613);
  not NOT_5278(g6836,I12379);
  not NOT_5279(g4020,I7781);
  not NOT_5280(g6212,I10973);
  not NOT_5281(g2404,g1276);
  not NOT_5282(I5548,g1280);
  not NOT_5283(I8895,g4130);
  not NOT_5284(g2647,I6425);
  not NOT_5285(g5529,g4689);
  not NOT_5286(g3159,I6856);
  not NOT_5287(I10166,g5016);
  not NOT_5288(g5148,I9570);
  not NOT_5289(g3359,I6946);
  not NOT_5290(g5649,g4748);
  not NOT_5291(g6918,I12609);
  not NOT_5292(g6967,I12696);
  not NOT_5293(I5555,g1288);
  not NOT_5294(I11269,g5756);
  not NOT_5295(I14166,g7702);
  not NOT_5296(I14009,g7436);
  not NOT_5297(g2764,g1802);
  not NOT_5298(g7265,g7077);
  not NOT_5299(g9324,I16072);
  not NOT_5300(g7042,g6543);
  not NOT_5301(g2546,I6368);
  not NOT_5302(I11773,g6262);
  not NOT_5303(g5155,I9591);
  not NOT_5304(g4559,g2898);
  not NOT_5305(g9069,I15601);
  not NOT_5306(I11942,g6015);
  not NOT_5307(I11341,g5809);
  not NOT_5308(I13773,g7496);
  not NOT_5309(g3858,I7377);
  not NOT_5310(g7442,I13583);
  not NOT_5311(g8583,I14668);
  not NOT_5312(I13341,g7207);
  not NOT_5313(g4931,I9301);
  not NOT_5314(I6248,g411);
  not NOT_5315(I7564,g2752);
  not NOT_5316(I9258,g4249);
  not NOT_5317(g3757,g1977);
  not NOT_5318(g2970,g2394);
  not NOT_5319(g6229,g5665);
  not NOT_5320(I15481,g8913);
  not NOT_5321(I10485,g5229);
  not NOT_5322(g6993,I12731);
  not NOT_5323(g1933,g1247);
  not NOT_5324(g7164,I13066);
  not NOT_5325(g7364,I13506);
  not NOT_5326(I6081,g118);
  not NOT_5327(g2925,g2324);
  not NOT_5328(g9177,I15811);
  not NOT_5329(g7233,g6940);
  not NOT_5330(g9206,g9196);
  not NOT_5331(I10555,g5529);
  not NOT_5332(I10454,g5217);
  not NOT_5333(g6822,I12337);
  not NOT_5334(g3522,g2407);
  not NOT_5335(I14454,g8177);
  not NOT_5336(g7054,g6511);
  not NOT_5337(g2224,I5945);
  not NOT_5338(g3642,I7118);
  not NOT_5339(I13734,g7422);
  not NOT_5340(g3047,g1736);
  not NOT_5341(I10914,g5448);
  not NOT_5342(I11335,g5839);
  not NOT_5343(g7454,I13610);
  not NOT_5344(g4628,I8799);
  not NOT_5345(I14712,g8059);
  not NOT_5346(I13335,g7206);
  not NOT_5347(g7770,I14181);
  not NOT_5348(g5463,g5085);
  not NOT_5349(I6154,g122);
  not NOT_5350(g7296,I13320);
  not NOT_5351(I6354,g1357);
  not NOT_5352(g4630,I8805);
  not NOT_5353(I13930,g7405);
  not NOT_5354(g7725,I14046);
  not NOT_5355(I11838,g6281);
  not NOT_5356(I5908,g196);
  not NOT_5357(g4300,I8261);
  not NOT_5358(g7532,I13776);
  not NOT_5359(g1724,I5568);
  not NOT_5360(I7308,g3074);
  not NOT_5361(g3874,g2957);
  not NOT_5362(I12208,g6496);
  not NOT_5363(I13131,g6951);
  not NOT_5364(g3654,g2521);
  not NOT_5365(g9199,g9188);
  not NOT_5366(I15784,g9125);
  not NOT_5367(g8647,I14739);
  not NOT_5368(I15956,g9216);
  not NOT_5369(g2617,g1565);
  not NOT_5370(g2906,g2288);
  not NOT_5371(I15385,g8880);
  not NOT_5372(g1878,g80);
  not NOT_5373(g5167,I9627);
  not NOT_5374(I14238,g7608);
  not NOT_5375(g5367,I9834);
  not NOT_5376(g5872,I10561);
  not NOT_5377(I13487,g7129);
  and AND2_0(g7412,g7121,g4841);
  and AND2_1(g6462,g6215,g2424);
  and AND2_2(g8925,g4592,g8754);
  and AND2_3(g4969,g4362,g2216);
  and AND2_4(g7429,g1057,g7212);
  and AND2_5(g9144,g9123,g6096);
  and AND2_6(g9344,g9329,g6211);
  and AND2_7(g4123,g2627,g2617);
  and AND2_8(g8320,g4557,g7951);
  and AND4_0(I8431,g3430,g3398,g3359,g3341);
  and AND2_9(g9259,g9230,g5639);
  and AND2_10(g8277,g162,g8042);
  and AND4_1(I8005,g3430,g3398,g3359,g2106);
  and AND2_11(g4351,g309,g3131);
  and AND2_12(g8299,g591,g8181);
  and AND2_13(g6941,g1126,g6582);
  and AND2_14(g4410,g408,g3160);
  and AND2_15(g8892,g8681,g4969);
  and AND4_2(I7994,g3430,g3398,g3359,g3341);
  and AND2_16(g5552,g1114,g4832);
  and AND2_17(g8945,g4541,g8784);
  and AND2_18(g8738,g8619,g3338);
  and AND2_19(g6431,g5847,g5494);
  and AND2_20(g4172,I8057,I8058);
  and AND2_21(g7449,g7272,g6901);
  and AND2_22(g8709,g2818,g8386);
  and AND2_23(g6176,g1149,g5198);
  and AND2_24(g6005,g5557,g2407);
  and AND2_25(g4343,g306,g3131);
  and AND2_26(g8078,g7463,g7634);
  and AND2_27(g8340,g423,g7920);
  and AND2_28(g6405,g5956,g5494);
  and AND2_29(g4282,g3549,g3568);
  and AND2_30(g7604,g7456,g3466);
  and AND2_31(g1714,g1454,g1450);
  and AND2_32(g5570,g1759,g4841);
  and AND2_33(g8690,g3485,g8363);
  and AND2_34(g7833,g6461,g7601);
  and AND2_35(g4334,g225,g3097);
  and AND2_36(g8876,g8769,g6102);
  and AND2_37(g6733,g685,g5873);
  and AND2_38(g6974,g3613,g6505);
  and AND2_39(g4804,g952,g3876);
  and AND2_40(g8915,g8794,g8239);
  and AND2_41(g7419,g7230,g3530);
  and AND2_42(g8310,g573,g8181);
  and AND2_43(g4494,I8546,I8547);
  and AND2_44(g8824,g264,g8524);
  and AND2_45(g8877,g8773,g6104);
  and AND2_46(g6399,g5971,g5494);
  and AND3_0(I9330,g2784,g2770,g2746);
  and AND2_47(g9142,g9124,g6059);
  and AND2_48(g8928,g4595,g8757);
  and AND2_49(g5020,g579,g3937);
  and AND4_3(g4933,g2746,g2728,g4320,g2770);
  and AND2_50(g8930,g3866,g8760);
  and AND4_4(I8114,g2162,g2149,g2137,g2106);
  and AND2_51(g8064,g7483,g7634);
  and AND2_52(g7678,g7367,g4158);
  and AND2_53(g4724,g828,g4038);
  and AND2_54(g7087,g6440,g5311);
  and AND2_55(g4379,g399,g3160);
  and AND2_56(g8295,g4512,g7905);
  and AND2_57(g8237,g89,g8131);
  and AND2_58(g6923,g6570,g5612);
  and AND3_1(g4878,g2573,g2562,I9222);
  and AND2_59(g8844,g4056,g8602);
  and AND4_5(I8594,g3316,g2057,g2020,g1987);
  and AND3_2(I9166,g4041,g2595,g2584);
  and AND2_60(g8089,g840,g7658);
  and AND2_61(g8731,g2743,g8421);
  and AND2_62(g4271,g3666,g3684);
  and AND2_63(g6951,g5511,g6595);
  and AND2_64(g8071,g7540,g4969);
  and AND2_65(g8705,g2798,g8421);
  and AND2_66(g4799,g951,g4596);
  and AND4_6(I8033,g3430,g3398,g3359,g2106);
  and AND2_67(g8948,g4570,g8789);
  and AND2_68(g5969,g5564,g2424);
  and AND2_69(g7602,g7476,g3466);
  and AND2_70(g7007,g6627,g5072);
  and AND2_71(g5123,g516,g4033);
  and AND2_72(g4132,g2637,g2633);
  and AND4_7(I8496,g3316,g3287,g2020,g1987);
  and AND3_3(g4238,g2695,g2698,I8157);
  and AND2_73(g8814,g3880,g8463);
  and AND2_74(g6408,g669,g6019);
  and AND2_75(g8150,g846,g7658);
  and AND2_76(g4744,g3525,g4296);
  and AND2_77(g8438,g649,g7793);
  and AND2_78(g6972,g5661,g6498);
  and AND2_79(g7415,g7222,g5603);
  and AND2_80(g8836,g348,g8545);
  and AND3_4(g4901,g3723,g4288,I9261);
  and AND2_81(g6433,g778,g6134);
  and AND2_82(g8229,g8180,g5680);
  and AND2_83(g9349,g9340,g5690);
  and AND2_84(g8822,g417,g8564);
  and AND2_85(g6395,g2157,g6007);
  and AND2_86(g8921,g4579,g8747);
  and AND2_87(g7689,g7367,g4417);
  and AND2_88(g5334,g4887,g2424);
  and AND2_89(g5548,g1549,g4826);
  and AND2_90(g4968,g4403,g1760);
  and AND2_91(g6266,g1481,g5285);
  and AND2_92(g8837,g426,g8564);
  and AND2_93(g7030,g6705,g5723);
  and AND2_94(g8062,g7476,g7634);
  and AND2_95(g8620,g751,g8199);
  and AND2_96(g8462,g49,g8199);
  and AND2_97(g9119,g9049,g5345);
  and AND4_8(I8001,g2074,g3287,g2020,g1987);
  and AND2_98(g7564,g7367,g4172);
  and AND2_99(g9258,g9227,g5628);
  and AND4_9(I8401,g3316,g3287,g3264,g3238);
  and AND2_100(g4175,g1110,g3502);
  and AND2_101(g4375,g219,g3097);
  and AND2_102(g5313,g4820,g2407);
  and AND2_103(g6726,g5897,g5367);
  and AND2_104(g6154,g1499,g5713);
  and AND2_105(g8842,g429,g8564);
  and AND2_106(g7609,g7467,g3466);
  and AND2_107(g8298,g553,g8181);
  and AND2_108(g5094,g535,g4004);
  and AND2_109(g9274,g4748,g9255);
  and AND2_110(g4139,I8000,I8001);
  and AND2_111(g4384,g246,g3097);
  and AND2_112(g4838,g4517,g1760);
  and AND2_113(g8854,g443,g8564);
  and AND2_114(g7217,g1142,g6941);
  and AND2_115(g8941,g3882,g8776);
  and AND2_116(g4424,g489,g3192);
  and AND2_117(g6979,g5095,g6511);
  and AND2_118(g5593,g4110,g4969);
  and AND3_5(g6112,g5673,g4841,g5541);
  and AND2_119(g4077,g1284,g3582);
  and AND2_120(g6001,g5540,g2407);
  and AND2_121(g6401,g5971,g5367);
  and AND2_122(g8708,g3557,g8407);
  and AND2_123(g7827,g7575,g7173);
  and AND2_124(g5050,g587,g3970);
  and AND2_125(g1725,g1409,g1416);
  and AND2_126(g6727,g681,g5846);
  and AND2_127(g8405,g741,g8018);
  and AND2_128(g4099,g117,g3647);
  and AND2_129(g4304,g2784,g3779);
  and AND2_130(g8829,g267,g8524);
  and AND2_131(g8286,g180,g8156);
  and AND2_132(g8911,g8798,g7688);
  and AND2_133(g8733,g2996,g8493);
  and AND2_134(g8270,g110,g8131);
  and AND2_135(g8610,g665,g7887);
  and AND2_136(g9345,g9330,g6217);
  and AND3_6(g4269,g2354,g3563,I8209);
  and AND4_10(I8524,g3316,g2057,g3264,g1987);
  and AND2_137(g2781,g1600,g976);
  and AND2_138(g8069,g7456,g7634);
  and AND2_139(g4712,g1179,g4276);
  and AND2_140(g7181,g6124,g7039);
  and AND2_141(g9159,g9138,g6074);
  and AND2_142(g9359,g4748,g9340);
  and AND2_143(g8377,g507,g7966);
  and AND2_144(g7197,g7093,g5055);
  and AND2_145(g7700,g7367,g4494);
  and AND2_146(g7021,g3390,g6673);
  and AND2_147(g4729,g1504,g4059);
  and AND2_148(g4961,g377,g3904);
  and AND2_149(g9016,g8904,g8239);
  and AND2_150(g8287,g4500,g7855);
  and AND4_11(I8186,g3778,g3549,g3568,g3583);
  and AND2_151(g5132,I9534,I9535);
  and AND2_152(g8849,g513,g8585);
  and AND4_12(I7995,g2074,g3287,g2020,g3238);
  and AND2_153(g9251,g4748,g9230);
  and AND2_154(g4414,I8412,I8413);
  and AND3_7(g3313,g2334,g2316,g2298);
  and AND2_155(g7631,g7367,g4187);
  and AND2_156(g8291,g122,g8111);
  and AND2_157(g3094,g945,g1898);
  and AND2_158(g4436,g492,g3192);
  and AND2_159(g6577,g6142,g4160);
  and AND2_160(g7605,g7435,g5607);
  and AND2_161(g4378,g321,g3131);
  and AND2_162(g4135,I7994,I7995);
  and AND2_163(g5092,g456,g4002);
  and AND2_164(g4182,I8071,I8072);
  and AND4_13(g4288,g3563,g3579,g3603,I8240);
  and AND2_165(g9272,g4748,g9248);
  and AND2_166(g8259,g4538,g7855);
  and AND2_167(g5714,g1532,g4733);
  and AND2_168(g8088,g837,g7658);
  and AND2_169(g8852,g362,g8545);
  and AND2_170(g8923,g4587,g8751);
  and AND4_14(I8461,g3316,g3287,g2020,g3238);
  and AND2_171(g7041,g6734,g5206);
  and AND2_172(g4422,g411,g3160);
  and AND2_173(g8701,g2700,g8363);
  and AND2_174(g2768,g1597,g973);
  and AND2_175(g9328,g9324,g6465);
  and AND2_176(g4798,g4216,g1760);
  and AND2_177(g9130,g9054,g5345);
  and AND2_178(g6125,g5548,g4202);
  and AND2_179(g2972,g2397,g2407);
  and AND4_15(I8046,g2074,g2057,g3264,g1987);
  and AND2_180(g8951,g8785,g6072);
  and AND2_181(g8314,g443,g7920);
  and AND2_182(g4437,g540,g2845);
  and AND2_183(g8825,g342,g8545);
  and AND2_184(g8650,g591,g8094);
  and AND3_8(g4302,g3086,g3659,g3124);
  and AND2_185(g1728,g1432,g1439);
  and AND2_186(g8336,g420,g7920);
  and AND2_187(g6061,g5257,g1616);
  and AND2_188(g8943,g4560,g8781);
  and AND2_189(g6046,g1073,g5592);
  and AND4_16(I8115,g2074,g3287,g3264,g1987);
  and AND4_17(I8642,g3430,g3398,g3359,g2106);
  and AND2_190(g8322,g4559,g7993);
  and AND3_9(g6003,g3716,g5633,I10597);
  and AND2_191(g8934,g3873,g8766);
  and AND2_192(g9348,g9333,g6229);
  and AND2_193(g7713,g4403,g7367);
  and AND2_194(g6145,g1489,g5705);
  and AND2_195(g4054,g3767,g2424);
  and AND2_196(g4454,g544,g2845);
  and AND2_197(g5077,g236,g3988);
  and AND2_198(g4532,I8617,I8618);
  and AND2_199(g6107,g5478,g1849);
  and AND2_200(g8845,g432,g8564);
  and AND3_10(I9202,g2605,g4044,g2584);
  and AND2_201(g8337,g498,g7966);
  and AND2_202(g4412,g486,g3192);
  and AND2_203(g5104,g274,g4010);
  and AND2_204(g6757,g5874,g5412);
  and AND2_205(g9279,g9255,g5665);
  and AND2_206(g4389,g480,g3192);
  and AND4_18(I8612,g3430,g3398,g3359,g3341);
  and AND2_207(g6416,g710,g6026);
  and AND4_19(I8417,g3430,g3398,g3359,g2106);
  and AND2_208(g9118,g9046,g5345);
  and AND2_209(g4787,g953,g4547);
  and AND2_210(g6047,g1477,g5596);
  and AND2_211(g8266,g2157,g8042);
  and AND2_212(g6447,g734,g6073);
  and AND2_213(g4956,g295,g3892);
  and AND2_214(g2979,g1494,g1733);
  and AND2_215(g5044,g234,g3959);
  and AND2_216(g8081,g834,g7658);
  and AND2_217(g8815,g258,g8524);
  and AND2_218(g7183,g6132,g7042);
  and AND2_219(g7608,g7367,g4169);
  and AND2_220(g8692,g3462,g8363);
  and AND2_221(g8726,g2795,g8386);
  and AND2_222(g4138,g2638,g2634);
  and AND2_223(g4109,g990,g3790);
  and AND2_224(g4791,g949,g4562);
  and AND2_225(g4707,g812,g4062);
  and AND2_226(g6417,g718,g6027);
  and AND4_20(I8090,g3316,g2057,g2020,g3238);
  and AND4_21(I8490,g3430,g3398,g3359,g3341);
  and AND2_227(g4201,I8108,I8109);
  and AND2_228(g8267,g154,g8042);
  and AND2_229(g8312,g365,g7870);
  and AND2_230(g6629,g6023,g4841);
  and AND3_11(g4957,g2746,g2728,g4320);
  and AND2_231(g4049,g141,g3514);
  and AND4_22(I8456,g3316,g3287,g2020,g1987);
  and AND4_23(I8529,g3316,g2057,g3264,g3238);
  and AND2_232(g8293,g4510,g7855);
  and AND2_233(g8329,g527,g7966);
  and AND2_234(g7696,g7367,g4469);
  and AND2_235(g5513,g4889,g5071);
  and AND2_236(g4098,g985,g3790);
  and AND2_237(g6554,g5762,g1616);
  and AND2_238(g8828,g4573,g8541);
  and AND2_239(g8830,g345,g8545);
  and AND2_240(g8727,g2724,g8421);
  and AND2_241(g5436,g1541,g4926);
  and AND2_242(g7240,g6719,g6894);
  and AND4_24(I8063,g2162,g2149,g2137,g2106);
  and AND2_243(g8703,g3574,g8407);
  and AND2_244(g4268,g2216,g2655);
  and AND2_245(g8932,g3868,g8762);
  and AND2_246(g6166,g1509,g5725);
  and AND2_247(g8624,g754,g8199);
  and AND2_248(g8953,g8758,g6093);
  and AND2_249(g4052,g1276,g3522);
  and AND2_250(g8068,g7687,g5610);
  and AND2_251(g4452,g437,g3160);
  and AND3_12(g6056,g3760,g5286,g1695);
  and AND2_252(g6456,g6116,g2407);
  and AND4_25(I8057,g3430,g3398,g3359,g3341);
  and AND2_253(g7681,g7444,g5099);
  and AND2_254(g9158,g9137,g6070);
  and AND2_255(g5560,g3390,g5036);
  and AND2_256(g4086,g103,g3629);
  and AND2_257(g4728,g190,g4179);
  and AND2_258(g4486,I8528,I8529);
  and AND2_259(g8716,g3506,g8443);
  and AND2_260(g7596,g7428,g7028);
  and AND2_261(g4504,I8568,I8569);
  and AND2_262(g4185,g2636,g2632);
  and AND2_263(g9275,g9241,g5645);
  and AND2_264(g4385,g300,g3131);
  and AND2_265(g8848,g281,g8524);
  and AND2_266(g5579,g4090,g4841);
  and AND2_267(g4425,g536,g2845);
  and AND2_268(g2386,g1130,g1092);
  and AND2_269(g5442,g4679,g4202);
  and AND2_270(g6057,g1061,g5617);
  and AND2_271(g4131,g2630,g2622);
  and AND2_272(g8319,g255,g7838);
  and AND4_26(I8552,g3316,g2057,g3264,g1987);
  and AND2_273(g8258,g142,g8111);
  and AND2_274(g6971,g6424,g4969);
  and AND2_275(g8717,g2764,g8421);
  and AND2_276(g7597,g7316,g4841);
  and AND2_277(g7079,g4259,g6677);
  and AND2_278(g8274,g4580,g7951);
  and AND2_279(g4445,I8455,I8456);
  and AND2_280(g4091,g129,g3639);
  and AND2_281(g4491,g557,g2845);
  and AND2_282(g8325,g184,g8156);
  and AND2_283(g8821,g339,g8545);
  and AND2_284(g4169,I8052,I8053);
  and AND2_285(g5029,g212,g3945);
  and AND2_286(g4369,g580,g2845);
  and AND2_287(g8280,g114,g8111);
  and AND2_288(g8939,g3879,g8772);
  and AND2_289(g4407,g252,g3097);
  and AND2_290(g4059,g1499,g2979);
  and AND2_291(g4868,g4227,g4160);
  and AND2_292(g8306,g4525,g7951);
  and AND2_293(g4793,g3887,g4202);
  and AND2_294(g8461,g658,g7793);
  and AND2_295(g8622,g738,g7811);
  and AND2_296(g4246,g1106,g3226);
  and AND2_297(g8403,g639,g7793);
  and AND2_298(g8841,g351,g8545);
  and AND2_299(g5049,g474,g3969);
  and AND4_27(I8020,g2074,g3287,g2020,g1987);
  and AND2_300(g8695,g2709,g8363);
  and AND2_301(g8307,g432,g7920);
  and AND2_302(g9278,g9252,g5658);
  and AND2_303(g4388,g402,g3160);
  and AND2_304(g8359,g642,g7793);
  and AND2_305(g4216,I8114,I8115);
  and AND2_306(g9143,g9122,g6089);
  and AND2_307(g9343,g9328,g1738);
  and AND2_308(g7626,g7463,g3466);
  and AND2_309(g8858,g524,g8585);
  and AND2_310(g4430,I8436,I8437);
  and AND4_28(I9534,g3019,g3029,g3038,g3052);
  and AND2_311(g9334,g9318,g6205);
  and AND2_312(g8315,g4544,g7993);
  and AND2_313(g4826,g1545,g4239);
  and AND2_314(g6239,g1514,g5314);
  and AND2_315(g5019,g312,g3933);
  and AND2_316(g2935,g1612,g1077);
  and AND2_317(g7683,g1061,g7429);
  and AND2_318(g5452,g4876,g3499);
  and AND2_319(g8654,g570,g8094);
  and AND2_320(g6420,g5918,g5367);
  and AND2_321(g4108,g782,g3655);
  and AND3_13(g4883,g3746,g3723,g4288);
  and AND4_29(I8040,g3430,g3398,g3359,g3341);
  and AND2_322(g4066,g1280,g3532);
  and AND2_323(g8272,g158,g8042);
  and AND2_324(g4466,I8490,I8491);
  and AND2_325(g8978,g8909,g5587);
  and AND2_326(g8612,g673,g7887);
  and AND3_14(g3429,g1454,g1838,g1444);
  and AND2_327(g6204,g5542,g5294);
  and AND2_328(g4365,g237,g3097);
  and AND2_329(g4048,g1288,g3513);
  and AND2_330(g8935,g3874,g8767);
  and AND2_331(g5425,g1528,g4916);
  and AND2_332(g4448,I8460,I8461);
  and AND2_333(g4711,g190,g4072);
  and AND4_30(I8528,g3430,g3398,g3359,g2106);
  and AND2_334(g8328,g4571,g7993);
  and AND2_335(g4133,g2631,g2623);
  and AND2_336(g4333,g1087,g2782);
  and AND2_337(g8542,g661,g7887);
  and AND2_338(g8330,g261,g7838);
  and AND2_339(g4396,g459,g3192);
  and AND2_340(g9160,g9139,g6092);
  and AND2_341(g6040,g1462,g5578);
  and AND2_342(g5105,g354,g4013);
  and AND2_343(g7616,g7367,g4517);
  and AND2_344(g7561,g7367,g4163);
  and AND2_345(g4067,g133,g3539);
  and AND4_31(I8618,g2074,g3287,g3264,g3238);
  and AND3_15(I8143,g2674,g2677,g2680);
  and AND2_346(g3049,g2274,g1844);
  and AND2_347(g8090,g843,g7658);
  and AND2_348(g6151,g1494,g5709);
  and AND2_349(g8823,g4561,g8512);
  and AND2_350(g5045,g293,g3961);
  and AND2_351(g5091,g397,g4001);
  and AND2_352(g4181,g1142,g3512);
  and AND2_353(g8456,g703,g7811);
  and AND2_354(g9271,g4748,g9244);
  and AND2_355(g4397,g483,g3192);
  and AND2_356(g8851,g284,g8524);
  and AND2_357(g4421,g333,g3131);
  and AND2_358(g8698,g3774,g8342);
  and AND2_359(g8260,g138,g8111);
  and AND2_360(g5767,g5344,g3079);
  and AND2_361(g6172,g1514,g5192);
  and AND2_362(g9238,g4748,g9223);
  and AND2_363(g8720,g3825,g8421);
  and AND2_364(g4101,g108,g3649);
  and AND2_365(g8318,g183,g8156);
  and AND2_366(g8652,g563,g8094);
  and AND2_367(g8843,g507,g8585);
  and AND4_32(I8593,g3430,g3398,g3359,g2106);
  and AND2_368(g8457,g724,g7811);
  and AND3_16(I10597,g3769,g3754,g3735);
  and AND2_369(g1753,g819,g815);
  and AND2_370(g8686,g3819,g8342);
  and AND2_371(g7709,g7367,g4529);
  and AND2_372(g8321,g446,g7920);
  and AND2_373(g6908,g6478,g5246);
  and AND2_374(g4168,g1106,g3500);
  and AND2_375(g6567,g6265,g2424);
  and AND2_376(g4368,g318,g3131);
  and AND2_377(g8938,g3878,g8771);
  and AND2_378(g5428,g775,g4707);
  and AND2_379(g8813,g255,g8524);
  and AND2_380(g5030,g233,g3946);
  and AND2_381(g4058,g3656,g2407);
  and AND2_382(g4743,g3518,g4286);
  and AND2_383(g8740,g2966,g8493);
  and AND2_384(g6965,g55,g6489);
  and AND2_385(g4411,g462,g3192);
  and AND2_386(g8687,g3488,g8363);
  and AND2_387(g6160,g1504,g5718);
  and AND2_388(g3226,g1102,g1919);
  and AND2_389(g4074,g137,g3573);
  and AND2_390(g5108,g539,g4017);
  and AND2_391(g6641,g5939,g5494);
  and AND2_392(g7002,g6770,g5054);
  and AND2_393(g6996,g3678,g6552);
  and AND2_394(g5066,g395,g3978);
  and AND2_395(g8860,g527,g8585);
  and AND2_396(g8341,g501,g7966);
  and AND2_397(g8710,g2790,g8421);
  and AND2_398(g9384,g9383,g6245);
  and AND2_399(g8645,g550,g8094);
  and AND3_17(I8209,g2298,g2316,g2334);
  and AND2_400(g7657,g7367,g4201);
  and AND2_401(g8691,g3805,g8342);
  and AND2_402(g5048,g394,g3966);
  and AND2_403(g9024,g8884,g5317);
  and AND2_404(g8879,g8782,g6108);
  and AND2_405(g8607,g8154,g5616);
  and AND2_406(g8962,g8890,g5317);
  and AND2_407(g6611,g3390,g6249);
  and AND2_408(g1739,g803,g799);
  and AND2_409(g8275,g4581,g7993);
  and AND2_410(g8311,g4540,g7905);
  and AND2_411(g4400,g1138,g3614);
  and AND2_412(g6541,g6144,g3510);
  and AND4_33(I8574,g3316,g2057,g2020,g3238);
  and AND2_413(g5018,g232,g3930);
  and AND2_414(g5067,g454,g3980);
  and AND2_415(g5093,g477,g4003);
  and AND2_416(g9273,g4748,g9252);
  and AND2_417(g7557,g7367,g4147);
  and AND2_418(g4383,g222,g3097);
  and AND4_34(g4220,g3533,g3549,g3568,g3583);
  and AND2_419(g8380,g681,g7887);
  and AND2_420(g8832,g501,g8585);
  and AND2_421(g7071,g6639,g1872);
  and AND2_422(g4779,g4176,g1760);
  and AND2_423(g7705,g7367,g4514);
  and AND2_424(g8853,g365,g8545);
  and AND2_425(g7242,g7081,g6899);
  and AND2_426(g4423,g465,g3192);
  and AND2_427(g3188,g2298,g2316);
  and AND2_428(g5700,g1638,g4969);
  and AND2_429(g4361,g471,g3192);
  and AND2_430(g8931,g3867,g8761);
  and AND2_431(g4127,g2628,g2618);
  and AND2_432(g4451,g359,g3131);
  and AND2_433(g4327,g2959,g1867);
  and AND2_434(g6574,g1045,g5984);
  and AND2_435(g7038,g6466,g4841);
  and AND2_436(g8628,g753,g8199);
  and AND2_437(g8300,g126,g8111);
  and AND2_438(g9014,g8906,g8239);
  and AND2_439(g7212,g1053,g7010);
  and AND2_440(g5817,g5395,g3091);
  and AND2_441(g4472,g440,g3160);
  and AND2_442(g3466,g936,g2557);
  and AND2_443(g8440,g714,g7937);
  and AND4_35(I8523,g3430,g3398,g3359,g3341);
  and AND2_444(g5585,g4741,g4841);
  and AND4_36(I8643,g2074,g3287,g3264,g1987);
  and AND4_37(I9535,g3062,g2712,g4253,g2752);
  and AND2_445(g6175,g4332,g5614);
  and AND2_446(g8323,g524,g7966);
  and AND2_447(g9335,g9320,g6206);
  and AND2_448(g5441,g4870,g3497);
  and AND2_449(g4434,g356,g3131);
  and AND3_18(I9261,g3777,g3764,g3746);
  and AND2_450(g4147,I8014,I8015);
  and AND4_38(I8551,g3430,g3398,g3359,g2106);
  and AND2_451(g9022,g8887,g5317);
  and AND2_452(g4681,g4255,g3533);
  and AND2_453(g8151,g849,g7658);
  and AND2_454(g8648,g588,g8094);
  and AND2_455(g7837,g6470,g7610);
  and AND2_456(g5458,g4686,g1616);
  and AND2_457(g3509,g1637,g1616);
  and AND4_39(I8613,g2074,g3287,g3264,g1987);
  and AND2_458(g8839,g4050,g8581);
  and AND2_459(g9037,g8965,g5345);
  and AND2_460(g6643,g1860,g5868);
  and AND2_461(g4936,g214,g3888);
  and AND2_462(g4117,g2626,g2616);
  and AND4_40(g4317,g878,g3086,g1857,g3659);
  and AND2_463(g8278,g4589,g7993);
  and AND2_464(g7192,g7026,g3526);
  and AND2_465(g8282,g179,g8156);
  and AND2_466(g5080,g396,g3991);
  and AND2_467(g5573,g3011,g4841);
  and AND2_468(g8693,g3798,g8342);
  and AND2_469(g8334,g264,g7838);
  and AND4_41(I8014,g3430,g3398,g3359,g3341);
  and AND2_470(g1919,g1098,g1087);
  and AND2_471(g6044,g1467,g5584);
  and AND2_472(g7031,g3390,g6717);
  and AND2_473(g6444,g1676,g6125);
  and AND2_474(g7252,g3591,g6977);
  and AND2_475(g8621,g734,g7937);
  and AND2_476(g4937,g3086,g4309);
  and AND2_477(g8313,g4542,g7951);
  and AND2_478(g4840,g4235,g1980);
  and AND4_42(I8436,g3430,g3398,g3359,g2106);
  and AND2_479(g4190,g1122,g3527);
  and AND2_480(g4390,g560,g2845);
  and AND2_481(g5126,g556,g4037);
  and AND2_482(g9012,g8908,g8239);
  and AND3_19(I8288,g3666,g3684,g3694);
  and AND2_483(g4356,g468,g3192);
  and AND2_484(g9371,g9352,g5917);
  and AND2_485(g6414,g673,g6025);
  and AND2_486(g8264,g105,g8131);
  and AND2_487(g4163,I8040,I8041);
  and AND2_488(g8933,g4511,g8765);
  and AND2_489(g7177,g7016,g5586);
  and AND2_490(g4053,g1292,g3523);
  and AND2_491(g5588,g3028,g4969);
  and AND2_492(g4453,g495,g3192);
  and AND4_43(I8495,g3430,g3398,g3359,g2106);
  and AND4_44(I8437,g3316,g3287,g3264,g1987);
  and AND2_493(g6182,g1519,g5199);
  and AND2_494(g8724,g3822,g8464);
  and AND2_495(g8379,g691,g7793);
  and AND2_496(g7199,g1467,g7003);
  and AND2_497(g6916,g727,g6515);
  and AND2_498(g6022,g5595,g2424);
  and AND2_499(g8878,g8777,g6106);
  and AND2_500(g6422,g714,g6033);
  and AND2_501(g8289,g348,g7870);
  and AND2_502(g8835,g270,g8524);
  and AND2_503(g8271,g130,g8111);
  and AND2_504(g8611,g669,g7887);
  and AND2_505(g5043,g213,g3958);
  and AND3_20(I8296,g3666,g3684,g3707);
  and AND2_506(g6437,g859,g6050);
  and AND2_507(g5443,g1549,g4935);
  and AND2_508(g7694,g7367,g4448);
  and AND2_509(g5116,g355,g4021);
  and AND2_510(g8238,g100,g8131);
  and AND2_511(g5034,g583,g3956);
  and AND2_512(g8332,g417,g7920);
  and AND2_513(g7701,g7367,g4497);
  and AND2_514(g8153,g852,g7658);
  and AND2_515(g4778,g4169,g1760);
  and AND2_516(g8744,g3802,g8464);
  and AND2_517(g7215,g6111,g6984);
  and AND4_45(I8412,g3430,g3398,g3359,g3341);
  and AND2_518(g4782,g4187,g1760);
  and AND2_519(g6042,g1041,g5581);
  and AND4_46(I8029,g2074,g2057,g3264,g1987);
  and AND2_520(g8901,g8804,g5631);
  and AND2_521(g6054,g1057,g5611);
  and AND2_522(g4526,g2642,g741);
  and AND2_523(g7008,g6615,g5083);
  and AND2_524(g2889,g1612,g1077);
  and AND2_525(g7136,g4057,g6953);
  and AND2_526(g5117,g435,g4024);
  and AND2_527(g8714,g2873,g8407);
  and AND2_528(g9025,g8889,g5317);
  and AND4_47(I8109,g2074,g3287,g3264,g3238);
  and AND2_529(g4702,g4243,g1690);
  and AND2_530(g6412,g158,g6024);
  and AND2_531(g7228,g6688,g7090);
  and AND2_532(g6990,g799,g6517);
  and AND2_533(g8262,g4554,g7855);
  and AND2_534(g6171,g5363,g4841);
  and AND2_535(g8736,g3771,g8464);
  and AND2_536(g4276,g2216,g2618);
  and AND2_537(g6429,g168,g6035);
  and AND2_538(g7033,g6716,g5190);
  and AND2_539(g9131,g9055,g5345);
  and AND2_540(g8623,g755,g8199);
  and AND2_541(g8076,g7690,g3521);
  and AND2_542(g7096,g6677,g5101);
  and AND2_543(g8722,g2787,g8386);
  and AND2_544(g7195,g6984,g4226);
  and AND2_545(g1844,g792,g795);
  and AND2_546(g5937,g5562,g2407);
  and AND2_547(g5079,g375,g3990);
  and AND2_548(g4546,g2643,g746);
  and AND2_549(g5479,g5141,g5037);
  and AND2_550(g6745,g1872,g6198);
  and AND2_551(g8285,g118,g8111);
  and AND2_552(g9226,g9220,g5403);
  and AND2_553(g6109,g5453,g5335);
  and AND3_21(g4224,g2680,g2683,I8127);
  and AND2_554(g8384,g636,g7793);
  and AND2_555(g8339,g345,g7870);
  and AND4_48(g4320,g3728,g3750,g3768,I8299);
  and AND2_556(g8838,g504,g8585);
  and AND4_49(I8019,g3430,g3398,g3359,g2106);
  and AND2_557(g8737,g2992,g8493);
  and AND4_50(I8052,g2162,g2149,g2137,g2106);
  and AND2_558(g4906,g4320,g2728);
  and AND2_559(g4789,g2751,g4202);
  and AND2_560(g6049,g1045,g5597);
  and AND2_561(g8077,g859,g7616);
  and AND2_562(g7692,g7367,g4430);
  and AND2_563(g8643,g547,g8094);
  and AND2_564(g6715,g677,g5843);
  and AND2_565(g6098,g5681,g1247);
  and AND2_566(g5032,g313,g3950);
  and AND2_567(g5432,g1537,g4921);
  and AND2_568(g4299,g3233,g3358);
  and AND2_569(g9015,g8905,g8239);
  and AND2_570(g8742,g2973,g8493);
  and AND2_571(g8304,g4523,g7905);
  and AND2_572(g8926,g4593,g8755);
  and AND2_573(g6162,g1134,g5724);
  and AND2_574(g6268,g1092,g5309);
  and AND2_575(g7001,g3722,g6562);
  and AND2_576(g8273,g185,g8156);
  and AND2_577(g6419,g162,g6032);
  and AND2_578(g7676,g7367,g4216);
  and AND2_579(g6052,g1049,g5604);
  and AND4_51(g4078,g3753,g3732,g3712,g3700);
  and AND2_580(g8269,g4569,g7951);
  and AND2_581(g4959,g376,g3898);
  and AND4_52(I8006,g2074,g3287,g2020,g3238);
  and AND2_582(g4435,g414,g3160);
  and AND2_583(g4517,I8593,I8594);
  and AND2_584(g4690,g4081,g3078);
  and AND2_585(g4082,g1296,g3604);
  and AND2_586(g8712,g2804,g8386);
  and AND2_587(g8543,g706,g7887);
  and AND2_588(g7703,g7367,g4504);
  and AND2_589(g8729,g2999,g8493);
  and AND2_590(g8961,g8885,g5317);
  and AND2_591(g9247,g4748,g9227);
  and AND2_592(g8927,g4594,g8756);
  and AND4_53(I8045,g3430,g3398,g3359,g2106);
  and AND2_593(g5894,g1118,g5552);
  and AND2_594(g8660,g1069,g8147);
  and AND2_595(g8946,g4556,g8786);
  and AND2_596(g7677,g7503,g5073);
  and AND4_54(I8491,g3316,g2057,g3264,g3238);
  and AND2_597(g6006,g5575,g2424);
  and AND2_598(g4236,g3260,g3221);
  and AND2_599(g8513,g718,g7937);
  and AND2_600(g6406,g154,g6018);
  and AND2_601(g5475,g3801,g5022);
  and AND2_602(g3190,g1658,g2424);
  and AND2_603(g6105,g5618,g2817);
  and AND4_55(g4877,g3746,g3723,g4288,g3764);
  and AND2_604(g8378,g677,g7887);
  and AND2_605(g6487,g5750,g4969);
  and AND2_606(g7699,g7367,g4486);
  and AND2_607(g8335,g342,g7870);
  and AND2_608(g8831,g423,g8564);
  and AND2_609(g8288,g270,g7838);
  and AND2_610(g8382,g685,g7887);
  and AND2_611(g5484,g1037,g5096);
  and AND4_56(I8015,g2074,g2057,g3264,g3238);
  and AND2_612(g8749,g2989,g8493);
  and AND2_613(g4785,g1678,g4202);
  and AND2_614(g6045,g1472,g5591);
  and AND2_615(g5583,g1775,g4969);
  and AND2_616(g6091,g5712,g5038);
  and AND2_617(g8947,g4558,g8787);
  and AND2_618(g6407,g5956,g5367);
  and AND2_619(g6578,g6218,g3913);
  and AND2_620(g4194,I8089,I8090);
  and AND2_621(g8653,g573,g8094);
  and AND2_622(g4394,g381,g3160);
  and AND2_623(g8302,g4521,g7855);
  and AND2_624(g7186,g6600,g7044);
  and AND2_625(g6582,g1122,g5894);
  and AND2_626(g1733,g1489,g1481);
  and AND2_627(g8719,g2821,g8443);
  and AND2_628(g4705,g190,g3986);
  and AND2_629(g6415,g5988,g5367);
  and AND2_630(g7614,g7367,g4176);
  and AND2_631(g5970,g5605,g2424);
  and AND4_57(I8028,g3430,g3398,g3359,g3341);
  and AND2_632(g8265,g134,g8111);
  and AND2_633(g4955,g215,g3891);
  and AND3_22(g4254,g3583,g3568,g3549);
  and AND2_634(g4814,g150,g4265);
  and AND2_635(g4150,I8019,I8020);
  and AND2_636(g4038,g825,g2949);
  and AND2_637(g9021,g8886,g5317);
  and AND2_638(g8296,g351,g7870);
  and AND2_639(g4409,g384,g3160);
  and AND2_640(g8725,g3008,g8493);
  and AND4_58(I8108,g2162,g2149,g2137,g2106);
  and AND2_641(g6689,g1519,g6239);
  and AND2_642(g7027,g3390,g6698);
  and AND2_643(g5547,g4814,g1819);
  and AND2_644(g7427,g1472,g7199);
  and AND2_645(g1898,g959,g955);
  and AND4_59(I8589,g2074,g3287,g3264,g3238);
  and AND2_646(g6428,g5874,g5494);
  and AND2_647(g6430,g5874,g5384);
  and AND2_648(g7003,g1462,g6689);
  and AND4_60(I8455,g3430,g3398,g3359,g3341);
  and AND2_649(g7695,g7367,g4466);
  and AND2_650(g8281,g168,g8042);
  and AND2_651(g5078,g316,g3989);
  and AND2_652(g6638,g174,g5755);
  and AND2_653(g7536,g4414,g7367);
  and AND2_654(g8297,g429,g7920);
  and AND2_655(g5082,g476,g3994);
  and AND2_656(g8745,g2982,g8493);
  and AND3_23(g4837,g2573,g2562,I9202);
  and AND2_657(g8338,g570,g8181);
  and AND2_658(g8963,g8891,g5317);
  and AND2_659(g4062,g809,g2986);
  and AND2_660(g7416,g7140,g4969);
  and AND2_661(g8309,g550,g8181);
  and AND4_61(I8418,g3316,g3287,g3264,g3238);
  and AND2_662(g6448,g5918,g5384);
  and AND2_663(g6055,g5239,g4202);
  and AND2_664(g7654,g7367,g4142);
  and AND2_665(g4192,g1126,g3531);
  and AND2_666(g4392,g303,g3131);
  and AND2_667(g6196,g4927,g5615);
  and AND2_668(g6396,g661,g6008);
  and AND2_669(g8715,g2761,g8386);
  and AND2_670(g7537,g7363,g7411);
  and AND2_671(g8833,g4583,g8562);
  and AND2_672(g7017,g3390,g6706);
  and AND2_673(g7417,g7144,g1616);
  and AND2_674(g8584,g8146,g7034);
  and AND2_675(g9080,g9011,g5598);
  and AND2_676(g6418,g5897,g5494);
  and AND2_677(g6994,g3658,g6538);
  and AND2_678(g7128,g6926,g3047);
  and AND2_679(g8268,g4568,g7905);
  and AND2_680(g5064,g315,g3975);
  and AND2_681(g8362,g504,g7966);
  and AND2_682(g4958,g296,g3897);
  and AND2_683(g4176,I8063,I8064);
  and AND2_684(g4376,g243,g3097);
  and AND2_685(g7554,g7367,g4139);
  and AND2_686(g5563,g3390,g5070);
  and AND2_687(g1913,g1528,g1532);
  and AND2_688(g6021,g5594,g2424);
  and AND2_689(g6421,g5847,g5384);
  and AND2_690(g8728,g3815,g8464);
  and AND2_691(g8730,g2863,g8407);
  and AND4_62(g4225,g2686,g2689,g2692,g2695);
  and AND2_692(g8385,g695,g7811);
  and AND4_63(I8041,g2074,g2057,g2020,g3238);
  and AND2_693(g4073,g1300,g3567);
  and AND2_694(g4796,g950,g4584);
  and AND2_695(g8070,g863,g7616);
  and AND2_696(g5089,g273,g3998);
  and AND2_697(g4473,g518,g3192);
  and AND2_698(g5489,g4912,g5053);
  and AND2_699(g4124,g2641,g2640);
  and AND2_700(g4469,I8495,I8496);
  and AND2_701(g4377,g297,g3131);
  and AND4_64(I8058,g2074,g2057,g2020,g1987);
  and AND2_702(g8331,g339,g7870);
  and AND2_703(g9023,g8888,g5317);
  and AND4_65(g4287,g3563,g2334,g3579,I8237);
  and AND2_704(g7698,g7367,g4483);
  and AND2_705(g8087,g7471,g7634);
  and AND2_706(g8305,g362,g7870);
  and AND2_707(g4199,g93,g2769);
  and AND2_708(g5438,g1545,g4932);
  and AND2_709(g4781,g4182,g1760);
  and AND2_710(g6041,g5189,g4969);
  and AND2_711(g8748,g2721,g8483);
  and AND2_712(g9327,g9316,g5757);
  and AND2_713(g4797,g3893,g1616);
  and AND2_714(g9146,g9135,g6101);
  and AND2_715(g9346,g9331,g6222);
  and AND2_716(g3002,g871,g1834);
  and AND4_66(I8573,g3430,g3398,g3359,g2106);
  and AND2_717(g6168,g1138,g5191);
  and AND2_718(g7652,g7367,g4194);
  and AND2_719(g6058,g5561,g3501);
  and AND2_720(g7193,g6911,g1616);
  and AND4_67(I8569,g3316,g2057,g2020,g1987);
  and AND2_721(g6743,g730,g5916);
  and AND3_24(g4819,g2573,g2562,I9166);
  and AND2_722(g8283,g267,g7838);
  and AND2_723(g9240,g9223,g5261);
  and AND2_724(g8059,g7682,g7032);
  and AND2_725(g8920,g4578,g8746);
  and AND2_726(g8459,g655,g7793);
  and AND2_727(g6411,g5918,g5494);
  and AND2_728(g8718,g2774,g8386);
  and AND2_729(g7598,g7483,g3466);
  and AND2_730(g3222,g1537,g1913);
  and AND2_731(g8261,g174,g8042);
  and AND2_732(g6474,g6203,g2424);
  and AND2_733(g7625,g7367,g4182);
  and AND2_734(g8793,g8637,g5622);
  and AND2_735(g6992,g6610,g3519);
  and AND2_736(g7232,g6694,g7091);
  and AND4_68(I8000,g3430,g3398,g3359,g3341);
  and AND3_25(g4314,g3694,g3684,g3666);
  and AND4_69(I8400,g3430,g3398,g3359,g3341);
  and AND2_737(g9147,g9136,g6103);
  and AND2_738(g5062,g235,g3973);
  and AND2_739(g9347,g9332,g6226);
  and AND2_740(g4825,g4228,g1964);
  and AND2_741(g8721,g2703,g8464);
  and AND2_742(g7552,g7319,g5749);
  and AND2_743(g7606,g7471,g3466);
  and AND2_744(g4408,g330,g3131);
  and AND2_745(g9013,g8907,g8239);
  and AND2_746(g5298,g1912,g4814);
  and AND2_747(g6976,g4399,g6508);
  and AND2_748(g8940,g4543,g8775);
  and AND4_70(I8588,g3430,g3398,g3359,g3341);
  and AND3_26(g4230,g2683,g3491,I8143);
  and AND2_749(g6400,g150,g6011);
  and AND3_27(I8127,g2699,g2674,g2677);
  and AND2_750(g4433,g278,g3097);
  and AND2_751(g7691,g7367,g4427);
  and AND2_752(g5031,g292,g3948);
  and AND2_753(g7607,g7325,g4969);
  and AND2_754(g8826,g420,g8564);
  and AND2_755(g4395,g405,g3160);
  and AND2_756(g8741,g3787,g8464);
  and AND3_28(g5005,g2728,g4320,I9330);
  and AND2_757(g2827,g1889,g1690);
  and AND2_758(g6423,g5897,g5384);
  and AND2_759(g5765,g1695,g5428);
  and AND4_71(I8240,g2298,g2316,g2334,g2354);
  and AND4_72(I8072,g3316,g3287,g2020,g3238);
  and AND2_760(g8609,g7828,g4969);
  and AND2_761(g8308,g510,g7966);
  and AND2_762(g7615,g7488,g3466);
  and AND2_763(g3229,g1728,g2015);
  and AND2_764(g8066,g7488,g7634);
  and AND4_73(I8034,g2074,g2057,g3264,g3238);
  and AND2_765(g4142,I8005,I8006);
  and AND2_766(g4342,g228,g3097);
  and AND3_29(I9222,g4041,g4044,g2584);
  and AND2_767(g6999,g815,g6556);
  and AND4_74(g4255,g3605,g3644,g3635,I8186);
  and AND2_768(g6633,g5526,g5987);
  and AND2_769(g8711,g3542,g8407);
  and AND2_770(g5069,g566,g3983);
  and AND2_771(g4097,g2624,g2614);
  and AND2_772(g7832,g5343,g7599);
  and AND2_773(g4497,I8551,I8552);
  and AND2_774(g8455,g652,g7793);
  and AND2_775(g4154,g1098,g3495);
  and AND2_776(g8827,g498,g8585);
  and AND2_777(g8333,g563,g8181);
  and AND2_778(g6732,g5874,g5367);
  and AND2_779(g8846,g510,g8585);
  and AND2_780(g6753,g5939,g5384);
  and AND2_781(g7559,g7367,g4155);
  and AND4_75(I8413,g3316,g3287,g3264,g1987);
  and AND2_782(g5287,g786,g4724);
  and AND2_783(g4783,g948,g4527);
  and AND2_784(g6043,g1069,g5582);
  and AND4_76(g4312,g3666,g3684,g3694,g3707);
  and AND2_785(g7628,g7367,g4532);
  and AND2_786(g6434,g855,g6048);
  and AND2_787(g8290,g588,g8181);
  and AND2_788(g4129,g2629,g2621);
  and AND2_789(g8256,g95,g8131);
  and AND2_790(g4830,g4288,g3723);
  and AND2_791(g8816,g336,g8545);
  and AND2_792(g6914,g6483,g5246);
  and AND4_77(I8460,g3430,g3398,g3359,g2106);
  and AND2_793(g6013,g5589,g2424);
  and AND2_794(g6413,g5939,g5367);
  and AND2_795(g8700,g3784,g8342);
  and AND2_796(g7323,g4065,g7171);
  and AND2_797(g8263,g4555,g7905);
  and AND2_798(g8950,g4582,g8791);
  and AND2_799(g4068,g121,g3540);
  and AND4_78(I8079,g3316,g3287,g2020,g1987);
  and AND2_800(g5314,g1509,g4729);
  and AND2_801(g8723,g2706,g8421);
  and AND2_802(g8257,g146,g8042);
  and AND2_803(g8817,g4545,g8482);
  and AND2_804(g8301,g182,g8156);
  and AND2_805(g7010,g1049,g6574);
  and AND2_806(g6060,g1065,g5623);
  and AND2_807(g4699,g1557,g4276);
  and AND2_808(g6460,g6178,g2424);
  and AND2_809(g4398,g567,g2845);
  and AND2_810(g5008,g231,g3920);
  and AND2_811(g7278,g6965,g1745);
  and AND2_812(g6995,g6435,g1616);
  and AND2_813(g8441,g746,g8018);
  and AND2_814(g7235,g6699,g7094);
  and AND4_79(I8432,g3316,g3287,g2020,g3238);
  and AND2_815(g9084,g8964,g5345);
  and AND4_80(I8053,g3316,g3287,g3264,g3238);
  and AND2_816(g7282,g5830,g6939);
  and AND2_817(g5065,g374,g3977);
  and AND2_818(g5122,g436,g4030);
  and AND4_81(g4319,g3728,g3694,g3750,I8296);
  and AND2_819(g7693,g7367,g4445);
  and AND4_82(I8568,g3430,g3398,g3359,g3341);
  and AND2_820(g4352,g387,g3160);
  and AND2_821(g5033,g393,g3953);
  and AND3_30(I8157,g2686,g2689,g2692);
  and AND2_822(g8458,g756,g8199);
  and AND2_823(g5096,g1149,g4400);
  and AND2_824(g4186,g1118,g3520);
  and AND2_825(g9276,g9244,g5649);
  and AND2_826(g4386,g324,g3131);
  and AND2_827(g6954,g5518,g6601);
  and AND2_828(g8074,g855,g7616);
  and AND2_829(g6053,g1053,g5608);
  and AND2_830(g4083,g125,g3610);
  and AND2_831(g8080,g7467,g7634);
  and AND2_832(g4483,I8523,I8524);
  and AND2_833(g3259,g1976,g1960);
  and AND2_834(g8713,g2777,g8421);
  and AND2_835(g5142,g1677,g4202);
  and AND2_836(g6157,g1130,g5717);
  and AND2_837(g5081,g455,g3993);
  and AND2_838(g9120,g9052,g5345);
  and AND2_839(g4187,I8078,I8079);
  and AND2_840(g9277,g9248,g5654);
  and AND2_841(g4387,g378,g3160);
  and AND2_842(g8688,g3812,g8342);
  and AND2_843(g8857,g446,g8564);
  and AND2_844(g8976,g8903,g6588);
  and AND2_845(g4427,I8431,I8432);
  and AND2_846(g4514,I8588,I8589);
  and AND2_847(g5783,g1897,g5287);
  and AND2_848(g7724,g7337,g5938);
  and AND2_849(g7179,g6121,g7035);
  and AND2_850(g4403,I8400,I8401);
  and AND2_851(g8326,g258,g7838);
  and AND2_852(g4145,g2639,g2635);
  and AND2_853(g4391,g249,g3097);
  and AND2_854(g5001,g458,g3912);
  and AND2_855(g7658,g7367,g4150);
  and AND2_856(g4107,g2625,g2615);
  and AND2_857(g1834,g933,g929);
  and AND2_858(g7271,g6436,g6922);
  and AND2_859(g4159,g1102,g3498);
  and AND2_860(g8383,g730,g7937);
  and AND2_861(g8924,g4588,g8752);
  and AND2_862(g7611,g7367,g4507);
  and AND2_863(g8779,g8634,g7037);
  and AND2_864(g6949,g5483,g6589);
  and AND3_31(g4315,g3707,g3728,I8288);
  and AND2_865(g4047,g1272,g3503);
  and AND2_866(g8361,g426,g7920);
  and AND2_867(g6998,g4474,g6555);
  and AND2_868(g7238,g6707,g7098);
  and AND2_869(g5624,g5140,g2794);
  and AND2_870(g7680,g7367,g4166);
  and AND2_871(g8327,g336,g7870);
  and AND2_872(g6039,g1037,g5574);
  and AND2_873(g5068,g475,g3982);
  and AND2_874(g6439,g789,g6150);
  and AND4_83(I8546,g3430,g3398,g3359,g3341);
  and AND2_875(g8303,g284,g7838);
  and AND2_876(g8696,g3743,g8342);
  and AND2_877(g8732,g3808,g8464);
  and AND2_878(g4272,g3233,g3286);
  and AND2_879(g8944,g4539,g8783);
  and AND2_880(g5699,g1667,g4841);
  and AND2_881(g4417,I8417,I8418);
  and AND4_84(I8617,g3430,g3398,g3359,g2106);
  and AND2_882(g7600,g7460,g3466);
  and AND2_883(g4128,g98,g3693);
  and AND2_884(g3081,g1682,g1616);
  and AND2_885(g8316,g513,g7966);
  and AND4_85(I8299,g3666,g3684,g3694,g3707);
  and AND4_86(I8547,g3316,g2057,g2020,g3238);
  and AND2_886(g6970,g5035,g6490);
  and AND2_887(g8147,g1065,g7683);
  and AND2_888(g5119,g543,g4027);
  and AND2_889(g8697,g3761,g8342);
  and AND2_890(g8914,g8795,g8239);
  and AND4_87(g4902,g4304,g2770,g2746,g2728);
  and AND4_88(I8078,g2162,g2149,g2137,g2106);
  and AND2_891(g7175,g6893,g4841);
  and AND2_892(g5599,g4745,g4969);
  and AND2_893(g4490,g521,g3192);
  and AND3_32(g4823,g4238,g4230,g174);
  and AND2_894(g4166,I8045,I8046);
  and AND2_895(g8820,g261,g8524);
  and AND2_896(g4366,g216,g3097);
  and AND2_897(g8936,g3875,g8768);
  and AND2_898(g6771,g146,g6004);
  and AND2_899(g8317,g547,g8181);
  and AND2_900(g4529,I8612,I8613);
  and AND2_901(g5125,g517,g4036);
  and AND2_902(g7184,g6138,g7043);
  and AND2_903(g4155,I8028,I8029);
  and AND2_904(g5984,g1041,g5484);
  and AND2_905(g4355,g390,g3160);
  and AND2_906(g8922,g4586,g8750);
  and AND2_907(g6738,g5847,g5367);
  and AND2_908(g8060,g7535,g4841);
  and AND2_909(g5106,g398,g4015);
  and AND2_910(g6991,g5689,g6520);
  and AND2_911(g8460,g757,g8199);
  and AND2_912(g9038,g8966,g5345);
  and AND2_913(g8739,g3780,g8464);
  and AND2_914(g4720,g190,g4055);
  and AND2_915(g4118,g995,g3790);
  and AND2_916(g4167,g2783,g1616);
  and AND2_917(g4367,g240,g3097);
  and AND3_33(g4872,g1924,g4225,g4224);
  and AND2_918(g7634,g7367,g4549);
  and AND2_919(g8937,g4524,g8770);
  and AND2_920(g8079,g831,g7658);
  and AND2_921(g8294,g281,g7838);
  and AND2_922(g5046,g314,g3962);
  and AND2_923(g8840,g4590,g8582);
  and AND2_924(g4193,g145,g2727);
  and AND2_925(g4393,g327,g3131);
  and AND2_926(g4549,I8642,I8643);
  and AND2_927(g6915,g6493,g5246);
  and AND4_89(I8064,g3316,g3287,g3264,g1987);
  and AND2_928(g8942,g4522,g8780);
  and AND2_929(g2912,g1080,g1945);
  and AND2_930(g5107,g478,g4016);
  and AND2_931(g8704,g2829,g8386);
  and AND2_932(g6002,g5539,g2407);
  and AND2_933(g6402,g665,g6012);
  and AND2_934(g8954,g8763,g6097);
  and AND3_34(I8237,g2298,g2316,g2354);
  and AND2_935(g6762,g5847,g5412);
  and AND2_936(g4740,g2242,g4275);
  and AND4_90(g3258,g2298,g2316,g2334,g2354);
  and AND2_937(g5047,g373,g3964);
  and AND4_91(I8089,g2162,g2149,g2137,g2106);
  and AND2_938(g8912,g8796,g8239);
  and AND4_92(I8071,g2162,g2149,g2137,g2106);
  and AND2_939(g6464,g6177,g2424);
  and AND2_940(g8929,g3865,g8759);
  and AND2_941(g3614,g1134,g2386);
  and AND2_942(g7036,g6728,g5197);
  and AND2_943(g7679,g7447,g5084);
  and AND2_944(g8626,g752,g8199);
  and AND2_945(g3984,g2403,g3085);
  and AND2_946(g5017,g211,g3928);
  and AND2_947(g4691,g4219,g1690);
  and AND2_948(g2949,g822,g1753);
  and AND2_949(g7182,g6902,g4969);
  and AND2_950(g6394,g5988,g5494);
  and AND2_951(g4962,g457,g3905);
  and AND2_952(g4158,I8033,I8034);
  and AND2_953(g6966,g6580,g5580);
  and AND2_954(g8735,g2807,g8443);
  and AND2_955(g8075,g7460,g7634);
  and AND2_956(g8949,g4572,g8790);
  and AND2_957(g7632,g7445,g3548);
  and AND2_958(g7653,g7480,g5754);
  and AND2_959(g8292,g181,g8156);
  and AND2_960(g2952,g2474,g2215);
  and AND2_961(g6438,g4829,g6051);
  and AND2_962(g4284,g3260,g3314);
  and AND2_963(g4239,g1541,g3222);
  and AND2_964(g5090,g317,g4000);
  and AND2_965(g8646,g553,g8094);
  and AND2_966(g6409,g706,g6020);
  and AND2_967(g4180,g1114,g3511);
  and AND2_968(g9270,g4748,g9241);
  and AND2_969(g4380,g584,g2845);
  and AND2_970(g4832,g1110,g4246);
  and AND2_971(g8439,g699,g7811);
  and AND2_972(g2986,g806,g1739);
  and AND2_973(g4420,g275,g3097);
  and AND2_974(g4507,I8573,I8574);
  and AND2_975(g4794,g954,g4574);
  and AND2_976(g8702,g2837,g8386);
  and AND2_977(g8919,g4567,g8743);
  and AND2_978(g8952,g8788,g6075);
  and AND2_979(g8276,g150,g8042);
  and AND2_980(g5063,g294,g3974);
  and AND2_981(g4100,g113,g3648);
  and AND2_982(g7553,g7367,g4135);
  and AND2_983(g8404,g710,g7937);
  and AND2_984(g5118,g479,g4026);
  and AND2_985(g8764,g8231,g4969);
  or OR4_0(g5057,g3939,g3925,g3915,g3907);
  or OR4_1(I14941,g8275,g8323,g8459,g8380);
  or OR2_0(g5193,g5017,g4366);
  or OR2_1(g9291,g9273,g6216);
  or OR2_2(g5549,g2935,g4712);
  or OR2_3(g7029,g6433,g5765);
  or OR2_4(g7787,g4791,g7602);
  or OR2_5(g6249,g4066,g5313);
  or OR3_0(g8906,g8088,g8062,g8699);
  or OR2_6(g5232,g5082,g4412);
  or OR2_7(g8987,g8927,g8826);
  or OR2_8(g5253,g5116,g4451);
  or OR2_9(g7791,g4796,g7606);
  or OR4_2(I8225,g3062,g2712,g2734,g2752);
  or OR4_3(I15250,g8238,g8265,g8272,g8292);
  or OR2_10(g8991,g8931,g8831);
  or OR4_4(I9107,g4133,g4145,g4138,g4132);
  or OR2_11(g9008,g8948,g8857);
  or OR4_5(g2214,g1376,g1377,g1378,g1379);
  or OR2_12(g7575,g7323,g7142);
  or OR2_13(g9136,g8952,g9131);
  or OR3_1(g8907,g8081,g8064,g8707);
  or OR3_2(g8082,g7654,g7628,g7611);
  or OR2_14(g5710,g4958,g4351);
  or OR3_3(I9047,g4155,g4147,g4139);
  or OR2_15(g9122,g8953,g9084);
  or OR3_4(g6270,g1000,g5335,g1909);
  or OR2_16(g6610,g4180,g6061);
  or OR2_17(g6124,g5432,g4789);
  or OR2_18(g6980,g6745,g6028);
  or OR4_6(I14484,g7993,g7966,g7793,g7811);
  or OR2_19(g9137,g8877,g9118);
  or OR2_20(g9337,g9240,g9327);
  or OR2_21(g7086,g4101,g6464);
  or OR4_7(I15055,I15051,I15052,I15053,I15054);
  or OR4_8(I15111,g7951,g7920,g7983,g8181);
  or OR2_22(g5545,g3617,g4824);
  or OR2_23(g7025,g6541,g3095);
  or OR2_24(g4264,g2490,g3315);
  or OR2_25(g8899,g8839,g8652);
  or OR3_5(g8785,g8623,g8656,I14985);
  or OR4_9(I15019,g7951,g7920,g7983,g8181);
  or OR2_26(g6144,g4175,g5458);
  or OR2_27(g9154,g9142,g9021);
  or OR2_28(g9354,g9275,g9344);
  or OR4_10(I15018,g7855,g7838,g7905,g7870);
  or OR2_29(g4179,g207,g3083);
  or OR2_30(g7682,g6044,g7412);
  or OR2_31(g6694,g6151,g5573);
  or OR2_32(g5204,g5033,g4379);
  or OR2_33(g9267,g9251,g6225);
  or OR2_34(g9001,g8941,g8846);
  or OR4_11(g8966,g8741,g8745,g8912,g8850);
  or OR2_35(g7445,g4192,g7193);
  or OR4_12(g5040,g3900,g3895,g3890,g4363);
  or OR2_36(g5440,g4790,g4786);
  or OR4_13(I15102,I15098,I15099,I15100,I15101);
  or OR4_14(g2229,g1371,g1372,g1373,g1374);
  or OR4_15(I14771,g7993,g7966,g7793,g7811);
  or OR4_16(I15231,g8701,g8715,g8730,g8720);
  or OR2_37(g8773,I14959,I14960);
  or OR4_17(g8009,g3591,g7406,g7566,I14302);
  or OR2_38(g8769,I14951,I14952);
  or OR2_39(g7227,g6992,g3128);
  or OR2_40(g6934,g6422,g6430);
  or OR2_41(g8993,g8933,g8835);
  or OR2_42(g6913,g6733,g6738);
  or OR2_43(g5235,g5091,g4422);
  or OR2_44(g5343,g4690,g2862);
  or OR4_18(I15085,g8363,g8342,g8407,g8386);
  or OR2_45(g5566,g3617,g4810);
  or OR4_19(I14759,g7937,g7887,g8029,g8018);
  or OR4_20(I15054,g8363,g8342,g8407,g8386);
  or OR4_21(I15243,I15239,I15240,I15241,I15242);
  or OR4_22(I14758,g7993,g7966,g7793,g7811);
  or OR3_6(g4736,g4532,g4517,I9044);
  or OR2_46(g8895,g8823,g8646);
  or OR2_47(g7428,g6040,g7175);
  or OR2_48(g9352,g9343,g4526);
  or OR2_49(g7826,g4804,g7626);
  or OR3_7(g8788,g8620,g8658,I14990);
  or OR2_50(g5202,g5031,g4377);
  or OR2_51(g5518,g4744,g4118);
  or OR4_23(g4737,g4135,g4529,g4514,I9047);
  or OR2_52(g7165,g6434,g6908);
  or OR2_53(g5264,g5125,g4490);
  or OR4_24(g8176,g7566,g1030,g6664,g6452);
  or OR2_54(g9387,g9349,g9384);
  or OR4_25(g2206,g1363,g1364,g1365,g1366);
  or OR4_26(I14951,g8328,g8316,g8455,g8378);
  or OR4_27(g9046,g8744,g8749,g9016,g8862);
  or OR2_55(g6932,g6417,g6423);
  or OR3_8(I15169,g8483,g8464,g8514);
  or OR2_56(g9003,g8943,g8849);
  or OR4_28(g8796,g8150,g8078,g8070,g8360);
  or OR2_57(g8980,g8920,g8815);
  or OR2_58(g6716,g6162,g5588);
  or OR2_59(g7421,g6745,g7202);
  or OR2_60(g6699,g6154,g5579);
  or OR2_61(g5238,g5094,g4425);
  or OR2_62(g4927,g4318,g1590);
  or OR2_63(g5209,g5044,g4384);
  or OR4_29(I15084,g7951,g7920,g7983,g8181);
  or OR4_30(I15110,g7855,g7838,g7905,g7870);
  or OR2_64(g8900,g8840,g8653);
  or OR2_65(g5511,g4743,g4109);
  or OR2_66(g6717,g4082,g6005);
  or OR2_67(g3160,g1751,g449);
  or OR3_9(g8886,g8727,g8812,I15254);
  or OR4_31(g2230,g1380,g1381,g1382,g1383);
  or OR4_32(I15242,g8697,g8714,g8718,g8719);
  or OR2_68(g5722,g5001,g4361);
  or OR2_69(g2845,g1877,g576);
  or OR4_33(I15230,g8274,g8321,g8298,g8696);
  or OR4_34(I15265,I15261,I15262,I15263,I15264);
  or OR4_35(g4786,g4107,g4097,g4124,I9099);
  or OR3_10(I13553,g1166,g1167,g1170);
  or OR2_70(g8887,I15265,g8819);
  or OR2_71(g7080,g4086,g6462);
  or OR2_72(g4364,g2952,g1725);
  or OR2_73(g9148,g9143,g9024);
  or OR4_36(I14767,g7937,g7887,g8029,g8018);
  or OR2_74(g9355,g9276,g9345);
  or OR2_75(g3541,g1663,g1421);
  or OR3_11(I14990,g8337,g8379,g8543);
  or OR2_76(g5231,g5081,g4411);
  or OR2_77(g5205,g5034,g4380);
  or OR4_37(g8891,g8705,g8811,I15297,I15298);
  or OR4_38(I15041,g7855,g7838,g7905,g7870);
  or OR2_78(g6115,g3617,g5558);
  or OR4_39(I15275,g8693,g8703,g8712,g8717);
  or OR2_79(g4297,g3617,g3602);
  or OR2_80(g7220,g1304,g7062);
  or OR2_81(g5572,g5051,g1236);
  or OR2_82(g8154,g6054,g7607);
  or OR4_40(I14766,g7993,g7966,g7793,g7811);
  or OR2_83(g6935,g6429,g6431);
  or OR3_12(I15165,g8483,g8464,g8514);
  or OR2_84(g8979,g8919,g8813);
  or OR2_85(g5036,g4047,g2972);
  or OR2_86(g3339,g1424,g2014);
  or OR4_41(I15253,g8698,g8711,g8722,g8716);
  or OR2_87(g7443,g7192,g3158);
  or OR4_42(I14754,g7937,g7887,g8029,g8018);
  or OR3_13(I15175,g8483,g8464,g8514);
  or OR4_43(I15264,g8700,g8708,g8726,g8731);
  or OR2_88(g9358,g9279,g9348);
  or OR2_89(g7697,g7419,g3187);
  or OR2_90(g6698,g4073,g6001);
  or OR2_91(g6964,g6447,g6448);
  or OR2_92(g5208,g5043,g4383);
  or OR2_93(g9174,g9147,g8963);
  or OR4_44(I15021,I15017,I15018,I15019,I15020);
  or OR2_94(g9239,g7653,g9226);
  or OR2_95(g5265,g5126,g4491);
  or OR4_45(I15073,g7951,g7920,g7983,g8181);
  or OR4_46(I15274,g8306,g8361,g8299,g8687);
  or OR3_14(g6457,g6196,g6209,g4937);
  or OR2_96(g5233,g5089,g4420);
  or OR2_97(g6686,g4068,g5970);
  or OR3_15(I15292,g8704,g8710,g8805);
  or OR2_98(g8893,g8814,g8643);
  or OR4_47(g7784,g7406,g6664,g3492,I14219);
  or OR2_99(g6121,g5425,g4785);
  or OR3_16(I14366,g7566,g1030,g6664);
  or OR2_100(g5706,g4955,g4342);
  or OR2_101(g6740,g4100,g6022);
  or OR2_102(g4283,g3587,g2665);
  or OR2_103(g8984,g8924,g8822);
  or OR4_48(I15109,g8131,g8111,g8042,g8156);
  or OR2_104(g9123,g8954,g9037);
  or OR4_49(I15283,g8291,g8276,g8325,g8330);
  or OR2_105(g5138,g4108,g3049);
  or OR2_106(g7810,g4799,g7609);
  or OR2_107(g7363,g7136,g6903);
  or OR3_17(I9099,g4127,g4123,g4117);
  or OR2_108(g9151,g9144,g8961);
  or OR2_109(g6525,g6112,g5547);
  or OR2_110(g6710,g55,g6264);
  or OR4_50(I6209,g911,g916,g921,g883);
  or OR3_18(g8904,g8090,g8080,g8706);
  or OR2_111(g5707,g4956,g4343);
  or OR3_19(I14980,g8362,g8403,g8610);
  or OR2_112(g9010,g8950,g8860);
  or OR2_113(g5201,g5030,g4376);
  or OR3_20(g8763,g8232,I14941,I14942);
  or OR3_21(I9044,g4150,g4142,g4549);
  or OR2_114(g8637,g6057,g8071);
  or OR2_115(g5715,g4961,g4355);
  or OR2_116(g9282,g9270,g6238);
  or OR4_51(I15040,g8131,g8111,g8042,g8156);
  or OR2_117(g5052,g4049,g4054);
  or OR4_52(I15252,g8320,g8307,g8317,g8692);
  or OR2_118(g7782,g4783,g7598);
  or OR2_119(g6931,g6416,g6421);
  or OR4_53(I14969,g8315,g8377,g8359,g8611);
  or OR2_120(g5070,g4052,g4058);
  or OR4_54(g2213,g1367,g1368,g1369,g1370);
  or OR2_121(g8982,g8922,g8820);
  or OR2_122(g4055,g187,g3012);
  or OR3_22(g8128,g7566,g6910,g6452);
  or OR3_23(I11603,g6193,g6197,g6175);
  or OR2_123(g9264,g9247,g6242);
  or OR2_124(g6440,g6268,g5700);
  or OR2_125(g6123,g3617,g5556);
  or OR4_55(I15051,g8131,g8111,g8042,g8156);
  or OR4_56(I15072,g7855,g7838,g7905,g7870);
  or OR4_57(I14496,g7937,g7887,g8029,g8018);
  or OR2_126(g8902,g8844,g8654);
  or OR3_24(I15152,g8483,g8464,g8514);
  or OR2_127(g8155,g7632,g3219);
  or OR3_25(g8964,g8915,g8863,I15400);
  or OR2_128(g5227,g5077,g4407);
  or OR4_58(I15020,g8363,g8342,g8407,g8386);
  or OR2_129(g5203,g5032,g4378);
  or OR3_26(I9029,g4504,g4494,g4430);
  or OR2_130(g8989,g8929,g8829);
  or OR4_59(I15113,I15109,I15110,I15111,I15112);
  or OR2_131(g8834,g7096,g8229);
  or OR2_132(g5188,g5008,g4365);
  or OR2_133(g7435,g6052,g7182);
  or OR2_134(g7690,g4181,g7417);
  or OR2_135(g5216,g5062,g4391);
  or OR2_136(g3131,g1749,g368);
  or OR2_137(g8909,g6043,g8764);
  or OR3_27(g4734,g4469,g4448,I9038);
  or OR2_138(g6933,g6419,g6428);
  or OR4_60(I14480,g7937,g7887,g8029,g8018);
  or OR2_139(g9285,g9271,g6221);
  or OR4_61(I6208,g891,g896,g901,g906);
  or OR2_140(g5217,g5063,g4392);
  or OR2_141(g9139,g8879,g9120);
  or OR2_142(g9339,g9259,g9335);
  or OR2_143(g5711,g4959,g4352);
  or OR2_144(g7222,g6049,g6971);
  or OR4_62(I14942,g8439,g8440,g8405,g8460);
  or OR2_145(g4688,g4193,g3190);
  or OR2_146(g5196,g5020,g4369);
  or OR2_147(g6132,g5436,g4793);
  or OR2_148(g8985,g8925,g8824);
  or OR2_149(g7089,g4128,g6474);
  or OR2_150(g5256,g5119,g4454);
  or OR4_63(I14468,g7937,g7887,g8029,g8018);
  or OR4_64(g8794,g8153,g8074,g8069,g8523);
  or OR2_151(g5021,g943,g4501);
  or OR2_152(g7254,g6923,g5298);
  or OR2_153(g6600,g5443,g6055);
  or OR3_28(g8905,g8089,g8087,g8694);
  or OR2_154(g7438,g7184,g6978);
  or OR2_155(g6580,g6039,g6041);
  or OR2_156(g6262,g4074,g5334);
  or OR4_65(I15229,g8262,g8303,g8268,g8312);
  or OR4_66(I14479,g7993,g7966,g7793,g7811);
  or OR4_67(I15228,g8270,g8258,g8281,g8273);
  or OR2_157(g4072,g196,g2995);
  or OR2_158(g9135,g8951,g9130);
  or OR2_159(g9288,g9272,g6235);
  or OR4_68(I15112,g8363,g8342,g8407,g8386);
  or OR2_160(g5673,g4823,g4872);
  or OR2_161(g7062,g4048,g6456);
  or OR2_162(g4413,g2371,g3285);
  or OR3_29(g8884,g8735,g8818,I15232);
  or OR2_163(g7788,g4794,g7604);
  or OR2_164(g8988,g8928,g8827);
  or OR2_165(g6926,g6406,g6411);
  or OR2_166(g8804,g6060,g8609);
  or OR4_69(g9054,g8724,g8729,g9013,g8680);
  or OR4_70(I15298,g8332,g8333,g8686,g8702);
  or OR2_167(g6543,g6125,g1553);
  or OR3_30(g8908,g8079,g8066,g8855);
  or OR4_71(I14772,g7937,g7887,g8029,g8018);
  or OR4_72(I15232,I15228,I15229,I15230,I15231);
  or OR4_73(I15261,g8256,g8271,g8267,g8286);
  or OR2_168(g6927,g6408,g6413);
  or OR2_169(g9171,g9146,g8962);
  or OR4_74(g8965,g8739,g8742,g8914,g8847);
  or OR2_170(g5220,g5066,g4395);
  or OR2_171(g6436,g6266,g5699);
  or OR2_172(g8996,g8936,g8838);
  or OR2_173(g9138,g8878,g9119);
  or OR2_174(g9338,g9258,g9334);
  or OR2_175(g8777,I14969,I14970);
  or OR4_75(g9049,g8732,g8737,g9015,g8861);
  or OR4_76(I15031,g7951,g7920,g7983,g8181);
  or OR2_176(g8981,g8921,g8816);
  or OR3_31(g1690,g1021,g1025,g1018);
  or OR2_177(g8997,g8937,g8841);
  or OR2_178(g6579,g6098,g1975);
  or OR2_179(g7088,g6638,g6641);
  or OR2_180(g6719,g6166,g6171);
  or OR2_181(g6917,g6743,g6753);
  or OR2_182(g9162,g9158,g9022);
  or OR4_77(g4735,g4427,g4414,g4403,I9041);
  or OR4_78(g9052,g8728,g8733,g9014,g8679);
  or OR2_183(g5210,g5045,g4385);
  or OR4_79(g2262,g1384,g1385,g1386,g1387);
  or OR4_80(I15043,g8363,g8342,g8407,g8386);
  or OR2_184(g7825,g4801,g7615);
  or OR2_185(g3760,I7232,I7233);
  or OR3_32(I9041,g4483,g4466,g4445);
  or OR3_33(g5317,g4727,g4737,g4735);
  or OR4_81(I14952,g8456,g8513,g8458,g8236);
  or OR2_186(g6706,g4077,g6002);
  or OR2_187(g7230,g4190,g6995);
  or OR2_188(g9006,g8946,g8853);
  or OR3_34(g8889,I15283,I15284,I15285);
  or OR3_35(I14834,g8483,g8464,g8514);
  or OR2_189(g7337,g7278,g4546);
  or OR2_190(g6138,g5438,g5442);
  or OR4_82(I15086,I15082,I15083,I15084,I15085);
  or OR2_191(g6707,g6160,g5585);
  or OR4_83(g8795,g8151,g8077,g8075,g8279);
  or OR2_192(g7248,g7079,g5652);
  or OR2_193(g1955,g1189,g16);
  or OR2_194(g5704,g4936,g4334);
  or OR2_195(g9007,g8947,g8854);
  or OR2_196(g7081,g6172,g6629);
  or OR2_197(g9261,g9238,g6227);
  or OR2_198(g8634,g6047,g8060);
  or OR4_84(I15017,g8131,g8111,g8042,g8156);
  or OR2_199(g7783,g4787,g7600);
  or OR2_200(g8613,g8082,g7616);
  or OR2_201(g8983,g8923,g8821);
  or OR2_202(g4876,g4159,g4167);
  or OR2_203(g6728,g6168,g5593);
  or OR2_204(g6470,g5817,g2934);
  or OR3_36(g8885,g8723,g8806,I15243);
  or OR4_85(I7232,g2367,g2352,g2378,g2330);
  or OR2_205(g9165,g9159,g9023);
  or OR4_86(I15042,g7951,g7920,g7983,g8181);
  or OR4_87(g9055,g8721,g8725,g9012,g8859);
  or OR2_206(g6445,g6105,g6107);
  or OR3_37(g7258,g7083,g5403,I13220);
  or OR2_207(g6602,g6058,g3092);
  or OR2_208(g4295,g2828,g2668);
  or OR4_88(I15030,g7855,g7838,g7905,g7870);
  or OR2_209(g6920,g6395,g6399);
  or OR2_210(g5561,g4168,g4797);
  or OR3_38(g6459,g6259,g6185,I11603);
  or OR2_211(g6718,g4083,g6006);
  or OR2_212(g7026,g4186,g6554);
  or OR4_89(I14933,g8385,g8404,g8441,g8462);
  or OR3_39(g7426,g1173,g7217,I13553);
  or OR2_213(g7170,g6916,g6444);
  or OR3_40(g7083,g5448,g6267,g6710);
  or OR4_90(I15075,I15071,I15072,I15073,I15074);
  or OR2_214(g8990,g8930,g8830);
  or OR2_215(g8888,I15276,g8807);
  or OR2_216(g7191,g7071,g6980);
  or OR2_217(g5244,g5107,g4436);
  or OR2_218(g5140,g4333,g3509);
  or OR2_219(g7016,g6042,g6487);
  or OR2_220(g9168,g9160,g9025);
  or OR4_91(I15276,I15272,I15273,I15274,I15275);
  or OR3_41(I15285,g8709,g8713,g8803);
  or OR2_221(g5214,g5049,g4389);
  or OR4_92(I15053,g7951,g7920,g7983,g8181);
  or OR4_93(I15254,I15250,I15251,I15252,I15253);
  or OR2_222(g4249,g3617,g1639);
  or OR2_223(g3986,g202,g3129);
  or OR3_42(I14302,g6664,g3492,g979);
  or OR2_224(g9011,g6046,g8892);
  or OR4_94(I15101,g8363,g8342,g8407,g8386);
  or OR2_225(g5236,g5092,g4423);
  or OR2_226(g7272,g6182,g7038);
  or OR2_227(g8896,g8828,g8648);
  or OR2_228(g5222,g5068,g4397);
  or OR2_229(g4812,g2490,g4237);
  or OR2_230(g4829,g863,g4051);
  or OR2_231(g6685,g4067,g5969);
  or OR2_232(g5237,g5093,g4424);
  or OR4_95(I15074,g8363,g8342,g8407,g8386);
  or OR4_96(I15239,g8264,g8260,g8277,g8301);
  or OR2_233(g5194,g5018,g4367);
  or OR2_234(g9000,g8940,g8845);
  or OR2_235(g8897,g8833,g8650);
  or OR2_236(g7166,g6437,g6914);
  or OR2_237(g5242,g5105,g4434);
  or OR2_238(g5254,g5117,g4452);
  or OR4_97(I14932,g8278,g8329,g8461,g8382);
  or OR2_239(g6585,g3617,g6119);
  or OR2_240(g6673,g4053,g5937);
  or OR2_241(g5212,g5047,g4387);
  or OR2_242(g7167,g6438,g6915);
  or OR3_43(g8091,g7215,g6452,I14366);
  or OR4_98(I15083,g7855,g7838,g7905,g7870);
  or OR2_243(g5229,g5079,g4409);
  or OR4_99(I15284,g8335,g8340,g8290,g8691);
  or OR4_100(g6458,g6184,g6259,g6174,g6214);
  or OR2_244(g7834,g7724,g6762);
  or OR2_245(g6734,g6176,g5599);
  or OR2_246(g4870,g4154,g3081);
  or OR2_247(g7687,g6053,g7416);
  or OR2_248(g6688,g6145,g5570);
  or OR4_101(I15052,g7855,g7838,g7905,g7870);
  or OR4_102(I14959,g8322,g8308,g8438,g8612);
  or OR2_249(g5708,g2889,g4699);
  or OR2_250(g5219,g5065,g4394);
  or OR2_251(g6924,g6400,g6405);
  or OR3_44(I15400,g8736,g8748,g8740);
  or OR2_252(g9294,g9274,g6230);
  or OR3_45(g8758,g8655,I14932,I14933);
  or OR2_253(g9356,g9277,g9346);
  or OR2_254(g7020,g3617,g6578);
  or OR4_103(I15241,g8269,g8314,g8309,g8695);
  or OR4_104(I15100,g7951,g7920,g7983,g8181);
  or OR2_255(g9363,g9359,g6210);
  or OR2_256(g6116,g5546,g4681);
  or OR3_46(g6565,g2396,g6131,g1603);
  or OR2_257(g8994,g8934,g8836);
  or OR2_258(g5245,g5108,g4437);
  or OR2_259(g9357,g9278,g9347);
  or OR2_260(g3192,g1756,g530);
  or OR4_105(g4727,g4417,g4172,g4163,I9029);
  or OR2_261(g7040,g6439,g5783);
  or OR2_262(g5259,g5122,g4472);
  or OR3_47(I14831,g8483,g8464,g8514);
  or OR3_48(I9038,g4507,g4497,g4486);
  or OR4_106(I15082,g8131,g8111,g8042,g8156);
  or OR2_263(g5215,g5050,g4390);
  or OR4_107(I14753,g7993,g7966,g7793,g7811);
  or OR2_264(g2368,I6208,I6209);
  or OR2_265(g4747,g3984,g2912);
  or OR3_49(I13220,g58,g6258,g5418);
  or OR4_108(I15263,g8313,g8297,g8310,g8690);
  or OR2_266(g6739,g4099,g6021);
  or OR4_109(I5757,g969,g970,g966,g963);
  or OR3_50(I8363,g2655,g1163,g1160);
  or OR4_110(I14960,g8621,g8622,g8628,g8230);
  or OR2_267(g5228,g5078,g4408);
  or OR2_268(g5230,g5080,g4410);
  or OR3_51(g8890,I15290,I15291,I15292);
  or OR4_111(I15273,g8287,g8334,g8295,g8339);
  or OR2_269(g5195,g5019,g4368);
  or OR2_270(g9004,g8944,g8851);
  or OR2_271(g7202,g6028,g7071);
  or OR4_112(I15033,I15029,I15030,I15031,I15032);
  or OR2_272(g8992,g8932,g8832);
  or OR4_113(I14970,g8457,g8383,g8626,g8233);
  or OR2_273(g4280,I8224,I8225);
  or OR2_274(g6912,g4199,g6567);
  or OR2_275(g5255,g5118,g4453);
  or OR4_114(g4790,g4185,g4131,g4129,I9107);
  or OR2_276(g6929,g6412,g6418);
  or OR2_277(g7450,g6090,g7195);
  or OR4_115(g1872,g971,g962,g972,I5757);
  or OR2_278(g5218,g5064,g4393);
  or OR2_279(g6735,g4091,g6013);
  or OR2_280(g5830,g5714,g5142);
  or OR4_116(I15291,g8331,g8336,g8338,g8688);
  or OR4_117(I7233,g2315,g2385,g2294,g2395);
  or OR2_281(g5221,g5067,g4396);
  or OR4_118(I15029,g8131,g8111,g8042,g8156);
  or OR2_282(g2043,g1263,g1257);
  or OR2_283(g8999,g8939,g8843);
  or OR2_284(g8146,g6045,g7597);
  or OR4_119(I8224,g3019,g3029,g3038,g3052);
  or OR2_285(g5716,g4962,g4356);
  or OR2_286(g6919,g6771,g6394);
  or OR2_287(g9002,g8942,g8848);
  or OR2_288(g6952,g6633,g6204);
  or OR4_120(I15240,g8259,g8294,g8263,g8305);
  or OR4_121(I14495,g7993,g7966,g7793,g7811);
  or OR2_289(g5241,g5104,g4433);
  or OR3_52(I14985,g8341,g8384,g8542);
  or OR2_290(g3097,g1746,g287);
  or OR4_122(I15262,g8293,g8283,g8304,g8289);
  or OR2_291(g6925,g6402,g6407);
  or OR2_292(g6120,g3617,g5555);
  or OR2_293(g5211,g5046,g4386);
  or OR2_294(g6906,g6715,g6726);
  or OR4_123(I15099,g7855,g7838,g7905,g7870);
  or OR4_124(I15098,g8131,g8111,g8042,g8156);
  or OR4_125(I15251,g8302,g8288,g8311,g8296);
  or OR4_126(I15272,g8237,g8300,g8261,g8282);
  or OR2_295(g5483,g4740,g4098);
  or OR4_127(I15032,g8363,g8342,g8407,g8386);
  or OR2_296(g6907,g6727,g6732);
  or OR2_297(g9009,g8949,g8858);
  or OR2_298(g8995,g8935,g8837);
  or OR3_53(I14219,g979,g7566,g1865);
  or OR2_299(g5200,g5029,g4375);
  or OR2_300(g5345,g4736,g4734);
  or OR2_301(g5223,g5069,g4398);
  or OR4_128(I15071,g8131,g8111,g8042,g8156);
  or OR4_129(I14467,g7993,g7966,g7793,g7811);
  or OR3_54(I15147,g8483,g8464,g8514);
  or OR2_302(g6590,g3617,g6153);
  or OR3_55(I15172,g8483,g8464,g8514);
  or OR2_303(g6928,g6409,g6415);
  or OR2_304(g6930,g6414,g6420);
  or OR2_305(g5537,g3617,g4835);
  or OR2_306(g7436,g7183,g6975);
  or OR2_307(g5243,g5106,g4435);
  or OR2_308(g5234,g5090,g4421);
  or OR4_130(I15044,I15040,I15041,I15042,I15043);
  or OR2_309(g6705,g6157,g5583);
  or OR2_310(g8894,g8817,g8645);
  or OR3_56(g8782,g8624,g8659,I14980);
  or OR2_311(g9005,g8945,g8852);
  or OR2_312(g5213,g5048,g4388);
  or OR4_131(I15290,g8285,g8266,g8318,g8326);
  or OR4_132(g4374,g1182,g1186,g1179,I8363);
  or OR2_313(g8998,g8938,g8842);
  or OR2_314(g9124,g8876,g9038);
  or OR2_315(g5698,g5057,g5040);
  or OR4_133(I14485,g7937,g7887,g8029,g8018);
  or OR2_316(g5260,g5123,g4473);
  or OR2_317(g9377,g9371,g6757);
  or OR2_318(g6921,g6396,g6401);
  or OR2_319(g8986,g8926,g8825);
  or OR4_134(I15297,g8280,g8257,g8319,g8327);
  nand NAND2_0(I15888,g9192,I15887);
  nand NAND2_1(I7466,g2982,g1704);
  nand NAND2_2(I10092,g4881,g2177);
  nand NAND2_3(g5686,g5132,g1263);
  nand NAND2_4(I5521,g1098,I5519);
  nand NAND2_5(g4528,I8606,I8607);
  nand NAND2_6(g5625,g2044,g4957);
  nand NAND2_7(I7538,g2996,g1715);
  nand NAND2_8(I11143,g5493,I11142);
  nand NAND2_9(I7467,g2982,I7466);
  nand NAND2_10(g4839,g1879,g4269);
  nand NAND2_11(I10906,g5492,g2605);
  nand NAND2_12(I12575,g6574,g1049);
  nand NAND2_13(I7181,g795,I7179);
  nand NAND2_14(g4235,g1415,g2668);
  nand NAND2_15(g6286,I11178,I11179);
  nand NAND2_16(I7421,g2525,g2703);
  nand NAND2_17(g5141,I9548,I9549);
  nand NAND2_18(g6911,I12597,I12598);
  nand NAND2_19(g4548,I8636,I8637);
  nand NAND2_20(I15855,g9168,g9165);
  nand NAND2_21(I11110,g2734,I11108);
  nand NAND2_22(I11179,g3019,I11177);
  nand NAND2_23(g6473,g5269,g5988);
  nand NAND2_24(I6524,g1102,I6522);
  nand NAND2_25(I11178,g5466,I11177);
  nand NAND2_26(I8510,g2517,g2807);
  nand NAND2_27(I8245,g3506,I8243);
  nand NAND2_28(g4313,g3712,g3700);
  nand NAND2_29(I11186,g3029,I11184);
  nand NAND2_30(g6469,g5918,g5278);
  nand NAND2_31(I13685,g1977,g7237);
  nand NAND2_32(I6258,g837,I6257);
  nand NAND2_33(g6177,I10889,I10890);
  nand NAND2_34(I13800,g7429,g1061);
  nand NAND2_35(I15819,g9148,I15817);
  nand NAND2_36(I15818,g9151,I15817);
  nand NAND2_37(I5600,g1489,I5598);
  nand NAND2_38(g6287,I11185,I11186);
  nand NAND2_39(I9978,g4880,g2092);
  nand NAND2_40(I9243,g4305,I9241);
  nand NAND2_41(I6274,g840,I6273);
  nand NAND3_0(g5284,g4344,g4335,g4963);
  nand NAND2_42(I10745,g2100,I10743);
  nand NAND2_43(g5239,I9746,I9747);
  nand NAND2_44(I9234,g4310,I9233);
  nand NAND2_45(I6170,g843,g911);
  nand NAND2_46(I13587,g2556,g7234);
  nand NAND2_47(g6510,g5278,g5874);
  nand NAND2_48(I6939,g2161,g2051);
  nand NAND2_49(I11117,g3062,I11115);
  nand NAND2_50(g5559,g5132,g1257);
  nand NAND2_51(g3232,g2298,g2276);
  nand NAND2_52(I7531,g2487,g3787);
  nand NAND2_53(g3938,I7610,I7611);
  nand NAND2_54(I7505,g3802,I7503);
  nand NAND2_55(I7011,g2333,I7009);
  nand NAND2_56(I11123,g5517,I11122);
  nand NAND2_57(I11751,g6112,I11750);
  nand NAND2_58(g6701,I12032,I12033);
  nand NAND2_59(g4835,I9195,I9196);
  nand NAND2_60(I13639,g7257,I13638);
  nand NAND2_61(I10329,g2562,I10327);
  nand NAND2_62(g6215,I10981,I10982);
  nand NAND2_63(I6904,g2105,g1838);
  nand NAND2_64(I13638,g7257,g7069);
  nand NAND2_65(I10328,g5467,I10327);
  nand NAND2_66(g5750,I10314,I10315);
  nand NAND2_67(I7480,g3808,I7478);
  nand NAND2_68(I11841,g2548,g6158);
  nand NAND2_69(I7569,g3780,I7567);
  nand NAND2_70(I9964,g1938,I9963);
  nand NAND2_71(g3525,I7010,I7011);
  nand NAND2_72(g4332,g3681,g2368);
  nand NAND2_73(g7535,I13786,I13787);
  nand NAND2_74(I6757,g186,g1983);
  nand NAND2_75(I12051,g5956,g5939);
  nand NAND2_76(g3358,I6940,I6941);
  nand NAND2_77(I11116,g5481,I11115);
  nand NAND2_78(I11615,g6239,I11614);
  nand NAND2_79(I6522,g1919,g1102);
  nand NAND2_80(I9057,g4059,g1504);
  nand NAND2_81(I10991,g5632,g2389);
  nand NAND2_82(I9549,g4307,I9547);
  nand NAND2_83(I8255,g3825,I8253);
  nand NAND2_84(g4492,I8537,I8538);
  nand NAND3_1(g4714,g4344,g4335,g4328);
  nand NAND2_85(I11142,g5493,g3062);
  nand NAND2_86(I7423,g2703,I7421);
  nand NAND2_87(I11165,g3029,I11163);
  nand NAND2_88(I6234,g896,I6232);
  nand NAND2_89(I10744,g5550,I10743);
  nand NAND2_90(g5555,I9979,I9980);
  nand NAND2_91(I10849,g2595,I10847);
  nand NAND2_92(g4889,I9242,I9243);
  nand NAND2_93(g4476,I8511,I8512);
  nand NAND2_94(g6142,I10790,I10791);
  nand NAND2_95(I10848,g5490,I10847);
  nand NAND4_0(g4871,g3635,g3605,g4220,g3644);
  nand NAND2_96(g6497,g5278,g5847);
  nand NAND2_97(I7240,g1658,I7239);
  nand NAND2_98(g5567,g1879,g4883);
  nand NAND2_99(I10361,g1118,I10359);
  nand NAND2_100(I7443,g2973,g1701);
  nand NAND2_101(I13600,g7244,I13598);
  nand NAND2_102(I9691,g5096,g1037);
  nand NAND2_103(g6218,I10992,I10993);
  nand NAND2_104(g4231,g2276,g3258);
  nand NAND2_105(I11137,g3052,I11135);
  nand NAND2_106(I7533,g3787,I7531);
  nand NAND2_107(I11873,g2543,g6187);
  nand NAND2_108(I12552,g1462,I12550);
  nand NAND2_109(I9985,g4836,g2096);
  nand NAND2_110(I11614,g6239,g1519);
  nand NAND2_111(g7093,I12870,I12871);
  nand NAND2_112(g9191,I15856,I15857);
  nand NAND2_113(I6843,g205,I6842);
  nand NAND2_114(I8119,g1904,g3220);
  nand NAND2_115(I11122,g5517,g2712);
  nand NAND2_116(I8152,g38,I8150);
  nand NAND2_117(I7460,g2506,I7459);
  nand NAND2_118(I14473,g8147,I14472);
  nand NAND2_119(I10789,g5512,g2170);
  nand NAND2_120(I7937,g3614,g1138);
  nand NAND2_121(I11136,g5476,I11135);
  nand NAND2_122(I6232,g834,g896);
  nand NAND2_123(I7479,g2502,I7478);
  nand NAND2_124(I10359,g5552,g1118);
  nand NAND2_125(I6813,g210,g2052);
  nand NAND2_126(g1759,I5599,I5600);
  nand NAND2_127(g5558,I10000,I10001);
  nand NAND2_128(I6740,g195,I6739);
  nand NAND2_129(g4513,I8582,I8583);
  nand NAND2_130(I11164,g5469,I11163);
  nand NAND2_131(I8939,g4239,I8938);
  nand NAND2_132(g6119,I10744,I10745);
  nand NAND2_133(g7257,I13214,I13215);
  nand NAND2_134(I7156,g2331,g929);
  nand NAND2_135(g4679,I8939,I8940);
  nand NAND2_136(I11575,g5894,I11574);
  nand NAND2_137(g3518,I6997,I6998);
  nand NAND2_138(I8636,g2481,I8635);
  nand NAND3_2(g4831,g3635,g3605,g4220);
  nand NAND2_139(I11109,g5522,I11108);
  nand NAND2_140(g6893,I12551,I12552);
  nand NAND2_141(I11108,g5522,g2734);
  nand NAND2_142(g6274,I11102,I11103);
  nand NAND2_143(I9151,g3883,g1649);
  nand NAND2_144(I7453,g3226,I7452);
  nand NAND2_145(g6170,I10874,I10875);
  nand NAND2_146(I11750,g6112,g1486);
  nand NAND2_147(I7568,g2481,I7567);
  nand NAND2_148(g6280,I11136,I11137);
  nand NAND2_149(I7157,g2331,I7156);
  nand NAND2_150(I8637,g2743,I8635);
  nand NAND2_151(g4869,g4254,g3533);
  nand NAND2_152(I8536,g2506,g2798);
  nand NAND2_153(I9278,g4313,I9276);
  nand NAND2_154(g3658,I7149,I7150);
  nand NAND3_3(g6187,g5633,g3735,g3716);
  nand NAND2_155(I6275,g906,I6273);
  nand NAND2_156(I9235,g2180,I9233);
  nand NAND2_157(I10981,g5625,I10980);
  nand NAND2_158(g2395,I6274,I6275);
  nand NAND2_159(I9693,g1037,I9691);
  nand NAND2_160(I9548,g1952,I9547);
  nand NAND2_161(g7480,I13639,I13640);
  nand NAND2_162(I10899,g5520,g2752);
  nand NAND2_163(g1678,I5506,I5507);
  nand NAND2_164(I11757,g1758,g6118);
  nand NAND3_4(g5672,g5056,g5039,g5023);
  nand NAND2_165(g6695,I12016,I12017);
  nand NAND2_166(g3680,I7187,I7188);
  nand NAND2_167(g1682,I5520,I5521);
  nand NAND2_168(g6159,I10835,I10836);
  nand NAND2_169(I8537,g2506,I8536);
  nand NAND2_170(I13397,g1057,I13395);
  nand NAND2_171(I6905,g2105,I6904);
  nand NAND2_172(I8243,g2011,g3506);
  nand NAND2_173(I8328,g2721,I8326);
  nand NAND2_174(g2783,I6523,I6524);
  nand NAND2_175(I9965,g4869,I9963);
  nand NAND2_176(I6750,g1733,g1494);
  nand NAND2_177(I13213,g7065,g7082);
  nand NAND2_178(g5712,I10224,I10225);
  nand NAND2_179(g4745,I9070,I9071);
  nand NAND2_180(I11574,g5894,g1122);
  nand NAND3_5(g4309,g3002,g3124,g3659);
  nand NAND2_181(I10061,g4910,I10060);
  nand NAND2_182(I7616,g3008,g1721);
  nand NAND2_183(I8512,g2807,I8510);
  nand NAND2_184(g3889,I7437,I7438);
  nand NAND2_185(I10360,g5552,I10359);
  nand NAND2_186(I8166,g3231,I8164);
  nand NAND2_187(I7503,g2498,g3802);
  nand NAND2_188(g3722,I7215,I7216);
  nand NAND2_189(g4575,I8679,I8680);
  nand NAND2_190(I15863,g9174,I15862);
  nand NAND2_191(I13396,g7212,I13395);
  nand NAND2_192(I14472,g8147,g1069);
  nand NAND2_193(I14246,g1065,I14244);
  nand NAND2_194(I7277,g2497,g1898);
  nand NAND2_195(I10071,g4954,g2253);
  nand NAND2_196(I6172,g911,I6170);
  nand NAND2_197(I7617,g3008,I7616);
  nand NAND2_198(g6902,I12576,I12577);
  nand NAND2_199(I9153,g1649,I9151);
  nand NAND2_200(g7316,I13377,I13378);
  nand NAND2_201(g3231,g1889,g1904);
  nand NAND2_202(I6134,g846,I6133);
  nand NAND2_203(I12080,g5971,I12078);
  nand NAND2_204(I7892,g2979,I7891);
  nand NAND2_205(I8393,g2949,I8392);
  nand NAND2_206(g1910,g1435,g1439);
  nand NAND2_207(I13787,g1477,I13785);
  nand NAND2_208(I12031,g5918,g5897);
  nand NAND2_209(g5632,g2276,g4901);
  nand NAND2_210(g5095,I9476,I9477);
  nand NAND2_211(g4881,g2460,g4315);
  nand NAND2_212(g2352,I6171,I6172);
  nand NAND2_213(I7140,g2397,I7138);
  nand NAND2_214(g6463,g5918,g5278);
  nand NAND2_215(I7478,g2502,g3808);
  nand NAND2_216(I8121,g3220,I8119);
  nand NAND2_217(I6202,g831,I6201);
  nand NAND2_218(I13640,g7069,I13638);
  nand NAND2_219(g3613,I7086,I7087);
  nand NAND2_220(g5752,I10328,I10329);
  nand NAND2_221(I12869,g2536,g6618);
  nand NAND2_222(I8253,g2454,g3825);
  nand NAND2_223(I8938,g4239,g1545);
  nand NAND2_224(I6776,g1134,I6774);
  nand NAND2_225(I8606,g2487,I8605);
  nand NAND2_226(I7214,g815,g2091);
  nand NAND3_6(g4305,g3712,g3700,g3732);
  nand NAND2_227(I9476,g4038,I9475);
  nand NAND2_228(I13003,g7010,I13002);
  nand NAND2_229(I6996,g2275,g2242);
  nand NAND2_230(g5189,I9692,I9693);
  nand NAND2_231(I13786,g7427,I13785);
  nand NAND2_232(I6878,g1910,I6876);
  nand NAND2_233(g3679,I7180,I7181);
  nand NAND2_234(I8607,g2764,I8605);
  nand NAND2_235(I8659,g2471,I8658);
  nand NAND2_236(I9477,g1942,I9475);
  nand NAND2_237(g4227,I8133,I8134);
  nand NAND2_238(I6997,g2275,I6996);
  nand NAND2_239(I12079,g5988,I12078);
  nand NAND2_240(g6570,I11751,I11752);
  nand NAND2_241(I12078,g5988,g5971);
  nand NAND2_242(I12598,g1126,I12596);
  nand NAND2_243(I10889,g5590,I10888);
  nand NAND2_244(I10980,g5625,g2210);
  nand NAND2_245(I10888,g5590,g2259);
  nand NAND2_246(g2315,I6103,I6104);
  nand NAND2_247(g4502,I8559,I8560);
  nand NAND4_1(g6158,g3735,g3716,g5633,g3754);
  nand NAND2_248(g5575,I10039,I10040);
  nand NAND2_249(I11149,g5473,g3038);
  nand NAND2_250(I8559,g2502,I8558);
  nand NAND2_251(g6275,I11109,I11110);
  nand NAND2_252(g6615,I11842,I11843);
  nand NAND2_253(I7150,g1974,I7148);
  nand NAND2_254(g5539,I9947,I9948);
  nand NAND2_255(I7438,g3822,I7436);
  nand NAND2_256(I7009,g2295,g2333);
  nand NAND2_257(I15862,g9174,g9171);
  nand NAND2_258(I12017,g5847,I12015);
  nand NAND2_259(g6284,I11164,I11165);
  nand NAND2_260(g6180,I10900,I10901);
  nand NAND2_261(g4741,I9058,I9059);
  nand NAND2_262(I9946,g2128,g4905);
  nand NAND2_263(g4910,g2460,g4314);
  nand NAND2_264(I10625,g5314,g1514);
  nand NAND2_265(g2330,I6134,I6135);
  nand NAND2_266(g6559,g5814,g6109);
  nand NAND2_267(g3012,I6758,I6759);
  nand NAND2_268(g9202,I15881,I15882);
  nand NAND2_269(g3706,g1556,g2510);
  nand NAND2_270(I9182,g4231,I9181);
  nand NAND2_271(I9382,g4062,I9381);
  nand NAND2_272(I10060,g4910,g2226);
  nand NAND2_273(I10197,g4724,I10196);
  nand NAND2_274(I6500,g1913,I6499);
  nand NAND2_275(I10855,g5521,I10854);
  nand NAND2_276(I8151,g3229,I8150);
  nand NAND2_277(I13378,g1472,I13376);
  nand NAND2_278(I9947,g2128,I9946);
  nand NAND2_279(I11096,g2734,I11094);
  nand NAND2_280(I10867,g5480,I10866);
  nand NAND2_281(I5505,g1532,g1528);
  nand NAND2_282(I13802,g1061,I13800);
  nand NAND2_283(I10315,g1041,I10313);
  nand NAND3_7(g5305,g5009,g4335,g4328);
  nand NAND2_284(I6523,g1919,I6522);
  nand NAND2_285(I10819,g5567,I10818);
  nand NAND2_286(I12016,g5874,I12015);
  nand NAND2_287(I10818,g5567,g2039);
  nand NAND2_288(g5748,I10306,I10307);
  nand NAND2_289(I11549,g5984,g1045);
  nand NAND2_290(g9179,I15818,I15819);
  nand NAND2_291(I7085,g1753,g1918);
  nand NAND2_292(I7485,g2989,g1708);
  nand NAND2_293(I6104,g921,I6102);
  nand NAND2_294(I6499,g1913,g1537);
  nand NAND2_295(g4256,g3233,g1444);
  nand NAND2_296(I8134,g1646,I8132);
  nand NAND2_297(g7503,I13686,I13687);
  nand NAND2_298(I10094,g2177,I10092);
  nand NAND2_299(I6273,g840,g906);
  nand NAND2_300(g2367,I6202,I6203);
  nand NAND2_301(g4700,g2460,g4271);
  nand NAND2_302(I13002,g7010,g1053);
  nand NAND2_303(I9233,g4310,g2180);
  nand NAND2_304(I10019,g2174,I10017);
  nand NAND2_305(g4263,g3260,g1435);
  nand NAND2_306(I10196,g4724,g1958);
  nand NAND2_307(I10018,g4700,I10017);
  nand NAND2_308(g6282,I11150,I11151);
  nand NAND2_309(I10866,g5480,g2605);
  nand NAND2_310(I7270,g955,I7268);
  nand NAND2_311(I10001,g1929,I9999);
  nand NAND2_312(I7610,g2471,I7609);
  nand NAND2_313(I9171,g4244,I9169);
  nand NAND2_314(I10923,g5525,g2752);
  nand NAND2_315(I7069,g1639,I7068);
  nand NAND2_316(I10300,g2562,I10298);
  nand NAND3_8(g7244,g7050,g3757,g3739);
  nand NAND2_317(I7540,g1715,I7538);
  nand NAND2_318(g7140,I13003,I13004);
  nand NAND2_319(g5689,I10197,I10198);
  nand NAND2_320(I9745,g4826,g1549);
  nand NAND2_321(I9963,g1938,g4869);
  nand NAND2_322(g7082,I12853,I12854);
  nand NAND2_323(I6135,g916,I6133);
  nand NAND2_324(g3678,I7173,I7174);
  nand NAND2_325(I15881,g9190,I15880);
  nand NAND2_326(I11080,g2511,I11078);
  nand NAND2_327(I10854,g5521,g2584);
  nand NAND2_328(I6916,g2360,g1732);
  nand NAND2_329(g5564,I10018,I10019);
  nand NAND2_330(I8658,g2471,g2724);
  nand NAND2_331(I5696,g1513,I5695);
  nand NAND2_332(I7510,g2992,g1711);
  nand NAND2_333(I12853,g6701,I12852);
  nand NAND2_334(g4474,I8503,I8504);
  nand NAND2_335(I10314,g5484,I10313);
  nand NAND2_336(I6102,g849,g921);
  nand NAND2_337(I11843,g6158,I11841);
  nand NAND2_338(I10307,g3019,I10305);
  nand NAND2_339(g5589,I10061,I10062);
  nand NAND2_340(I8132,g3232,g1646);
  nand NAND2_341(I8680,g2706,I8678);
  nand NAND2_342(g3602,I7069,I7070);
  nand NAND2_343(I6752,g1494,I6750);
  nand NAND2_344(I6917,g2360,I6916);
  nand NAND2_345(g1775,I5620,I5621);
  nand NAND2_346(I7215,g815,I7214);
  nand NAND2_347(g3767,I7240,I7241);
  nand NAND2_348(I5697,g1524,I5695);
  nand NAND2_349(I8558,g2502,g2790);
  nand NAND2_350(I12053,g5939,I12051);
  nand NAND2_351(I6233,g834,I6232);
  nand NAND2_352(I10335,g5462,I10334);
  nand NAND2_353(g9205,I15898,I15899);
  nand NAND2_354(I8511,g2517,I8510);
  nand NAND2_355(I10993,g2389,I10991);
  nand NAND2_356(I14839,g1073,I14837);
  nand NAND2_357(g5538,g5132,g1266);
  nand NAND2_358(I15897,g9202,g9203);
  nand NAND2_359(I14838,g8660,I14837);
  nand NAND2_360(g7237,g7050,g3739);
  nand NAND2_361(I9070,g4400,I9069);
  nand NAND2_362(g6153,I10819,I10820);
  nand NAND2_363(g6680,g5403,g6252);
  nand NAND2_364(g8239,g8073,g8092);
  nand NAND2_365(I11171,g5477,I11170);
  nand NAND2_366(I6171,g843,I6170);
  nand NAND2_367(I10039,g4893,I10038);
  nand NAND2_368(I10306,g5470,I10305);
  nand NAND2_369(I10038,g4893,g2202);
  nand NAND2_370(g3028,I6775,I6776);
  nand NAND2_371(I11079,g5697,I11078);
  nand NAND2_372(I7891,g2979,g1499);
  nand NAND2_373(I10143,g4707,I10142);
  nand NAND2_374(I13599,g2551,I13598);
  nand NAND2_375(I11078,g5697,g2511);
  nand NAND2_376(I13598,g2551,g7244);
  nand NAND2_377(g5562,I10010,I10011);
  nand NAND2_378(I10791,g2170,I10789);
  nand NAND2_379(I15850,g9154,I15848);
  nand NAND2_380(I8339,g2966,I8338);
  nand NAND2_381(g5257,I9768,I9769);
  nand NAND2_382(I6759,g1983,I6757);
  nand NAND2_383(g5605,I10093,I10094);
  nand NAND2_384(g3883,g2276,g3188);
  nand NAND2_385(I11158,g3052,I11156);
  nand NAND2_386(I6201,g831,g891);
  nand NAND2_387(I9169,g1935,g4244);
  nand NAND2_388(g5751,I10321,I10322);
  nand NAND2_389(I9059,g1504,I9057);
  nand NAND2_390(g6476,g5939,g5269);
  nand NAND2_391(I11144,g3062,I11142);
  nand NAND2_392(I9767,g4832,g1114);
  nand NAND2_393(g6722,I12079,I12080);
  nand NAND2_394(I10223,g2522,g4895);
  nand NAND2_395(g6285,I11171,I11172);
  nand NAND2_396(I12577,g1049,I12575);
  nand NAND2_397(I6539,g2555,I6538);
  nand NAND2_398(I10321,g5459,I10320);
  nand NAND2_399(I13017,g6941,I13016);
  nand NAND2_400(g6424,I11550,I11551);
  nand NAND2_401(I10953,g5565,I10952);
  nand NAND2_402(I15857,g9165,I15855);
  nand NAND2_403(g6477,g5269,g5918);
  nand NAND2_404(g4820,I9170,I9171);
  nand NAND2_405(I10334,g5462,g2573);
  nand NAND2_406(I13687,g7237,I13685);
  nand NAND2_407(I11752,g1486,I11750);
  nand NAND2_408(I7068,g1639,g1643);
  nand NAND2_409(I12852,g6701,g6695);
  nand NAND2_410(I7468,g1704,I7466);
  nand NAND2_411(g6273,I11095,I11096);
  nand NAND2_412(I9826,g4729,g1509);
  nand NAND2_413(I8660,g2724,I8658);
  nand NAND2_414(I10000,g4839,I9999);
  nand NAND2_415(I10908,g2605,I10906);
  nand NAND2_416(I11842,g2548,I11841);
  nand NAND2_417(I7576,g1718,I7574);
  nand NAND2_418(I7149,g799,I7148);
  nand NAND2_419(I12576,g6574,I12575);
  nand NAND2_420(I13016,g6941,g1142);
  nand NAND2_421(g4294,I8244,I8245);
  nand NAND2_422(I8679,g2467,I8678);
  nand NAND2_423(I7241,g2134,I7239);
  nand NAND2_424(I12052,g5956,I12051);
  nand NAND2_425(I15856,g9168,I15855);
  nand NAND2_426(I15880,g9190,g9179);
  nand NAND2_427(I10992,g5632,I10991);
  nand NAND2_428(I9827,g4729,I9826);
  nand NAND2_429(g7069,g5435,g6680);
  nand NAND2_430(I11124,g2712,I11122);
  nand NAND2_431(I8560,g2790,I8558);
  nand NAND2_432(g4954,g4319,g2460);
  nand NAND2_433(g4810,I9152,I9153);
  nand NAND2_434(g7540,I13801,I13802);
  nand NAND2_435(g4363,I8339,I8340);
  nand NAND2_436(I13686,g1977,I13685);
  nand NAND2_437(I9196,g1652,I9194);
  nand NAND2_438(I10835,g5514,I10834);
  nand NAND2_439(g6178,g2205,g5568);
  nand NAND2_440(I7893,g1499,I7891);
  nand NAND2_441(I7186,g2353,g1834);
  nand NAND2_442(I11875,g6187,I11873);
  nand NAND2_443(g4912,I9277,I9278);
  nand NAND2_444(g3890,I7444,I7445);
  nand NAND2_445(I9994,g4871,I9992);
  nand NAND2_446(g3011,I6751,I6752);
  nand NAND2_447(I7939,g1138,I7937);
  nand NAND2_448(I6203,g891,I6201);
  nand NAND2_449(I9181,g4231,g2007);
  nand NAND2_450(g5753,I10335,I10336);
  nand NAND2_451(I8164,g1943,g3231);
  nand NAND2_452(I9381,g4062,g1908);
  nand NAND2_453(I15887,g9192,g9191);
  nand NAND2_454(g7144,I13017,I13018);
  nand NAND2_455(I10142,g4707,g1916);
  nand NAND2_456(I6940,g2161,I6939);
  nand NAND2_457(I7187,g2353,I7186);
  nand NAND2_458(I7461,g3815,I7459);
  nand NAND2_459(g5565,g2044,g4933);
  nand NAND2_460(g5681,g5132,g2043);
  nand NAND2_461(g6265,I11079,I11080);
  nand NAND2_462(g5697,g2044,g5005);
  nand NAND2_463(I11170,g5477,g3038);
  nand NAND2_464(g6164,I10848,I10849);
  nand NAND2_465(I8956,g4246,I8955);
  nand NAND2_466(I6741,g1970,I6739);
  nand NAND2_467(g6770,I12180,I12181);
  nand NAND2_468(I13589,g7234,I13587);
  nand NAND2_469(I13588,g2556,I13587);
  nand NAND2_470(I8338,g2966,g1698);
  nand NAND2_471(g3924,I7568,I7569);
  nand NAND2_472(I10952,g5565,g2340);
  nand NAND2_473(I6758,g186,I6757);
  nand NAND2_474(I6066,g883,I6064);
  nand NAND2_475(g7065,I12833,I12834);
  nand NAND2_476(I11616,g1519,I11614);
  nand NAND2_477(I10790,g5512,I10789);
  nand NAND2_478(I9058,g4059,I9057);
  nand NAND2_479(I10873,g5516,g2595);
  nand NAND2_480(I8957,g1110,I8955);
  nand NAND2_481(g3665,I7157,I7158);
  nand NAND2_482(I6133,g846,g916);
  nand NAND2_483(g6281,I11143,I11144);
  nand NAND2_484(I6774,g2386,g1134);
  nand NAND2_485(I11101,g5491,g2712);
  nand NAND2_486(I11177,g5466,g3019);
  nand NAND2_487(I10834,g5514,g2584);
  nand NAND2_488(I6538,g2555,g2557);
  nand NAND2_489(I9992,g2145,g4871);
  nand NAND2_490(I11874,g2543,I11873);
  nand NAND2_491(I15817,g9151,g9148);
  nand NAND2_492(I12833,g6722,I12832);
  nand NAND2_493(I10320,g5459,g2573);
  nand NAND2_494(I10073,g2253,I10071);
  nand NAND2_495(g8231,I14473,I14474);
  nand NAND2_496(g5363,I9827,I9828);
  nand NAND2_497(g3681,g866,g2368);
  nand NAND2_498(I8504,g2038,I8502);
  nand NAND2_499(g3914,I7532,I7533);
  nand NAND2_500(I12951,g7003,g1467);
  nand NAND3_9(g5568,g2044,g4902,g4320);
  nand NAND2_501(I12033,g5897,I12031);
  nand NAND2_502(I8470,g2525,g2821);
  nand NAND2_503(I7512,g1711,I7510);
  nand NAND2_504(g9203,I15888,I15889);
  nand NAND2_505(I11185,g5474,I11184);
  nand NAND2_506(g4244,g3549,g3533);
  nand NAND2_507(I6257,g837,g901);
  nand NAND2_508(I7148,g799,g1974);
  nand NAND2_509(I9183,g2007,I9181);
  nand NAND2_510(I9383,g1908,I9381);
  nand NAND2_511(I14474,g1069,I14472);
  nand NAND2_512(I8678,g2467,g2706);
  nand NAND2_513(I10327,g5467,g2562);
  nand NAND2_514(g7828,I14245,I14246);
  nand NAND2_515(I8635,g2481,g2743);
  nand NAND2_516(I6751,g1733,I6750);
  nand NAND2_517(g6504,g5269,g5874);
  nand NAND2_518(I13215,g7082,I13213);
  nand NAND2_519(g2378,I6233,I6234);
  nand NAND2_520(I10982,g2210,I10980);
  nand NAND2_521(I7279,g1898,I7277);
  nand NAND2_522(I9999,g4839,g1929);
  nand NAND2_523(g4110,I7938,I7939);
  nand NAND2_524(g4310,g3666,g2460);
  nand NAND2_525(g4824,I9182,I9183);
  nand NAND2_526(g5661,I10143,I10144);
  nand NAND2_527(I8582,g2498,I8581);
  nand NAND2_528(I7938,g3614,I7937);
  nand NAND2_529(I5620,g1092,I5619);
  nand NAND2_530(I10040,g2202,I10038);
  nand NAND2_531(g8798,g6984,g8644);
  nand NAND2_532(g4563,I8659,I8660);
  nand NAND2_533(g6169,I10867,I10868);
  nand NAND2_534(g6283,I11157,I11158);
  nand NAND2_535(g4237,I8151,I8152);
  nand NAND2_536(I11576,g1122,I11574);
  nand NAND2_537(I8502,g2986,g2038);
  nand NAND2_538(I10847,g5490,g2595);
  nand NAND2_539(I8940,g1545,I8938);
  nand NAND2_540(I10062,g2226,I10060);
  nand NAND2_541(I11115,g5481,g3062);
  nand NAND2_542(g5546,I9964,I9965);
  nand NAND2_543(g7325,I13396,I13397);
  nand NAND2_544(I5520,g1087,I5519);
  nand NAND2_545(g6203,I10953,I10954);
  nand NAND2_546(I11184,g5474,g3029);
  nand NAND2_547(I7158,g929,I7156);
  nand NAND2_548(I6924,g1728,I6923);
  nand NAND2_549(I12832,g6722,g6709);
  nand NAND2_550(I10072,g4954,I10071);
  nand NAND2_551(g4836,g4288,g1879);
  nand NAND2_552(g3894,I7460,I7461);
  nand NAND2_553(g6188,I10924,I10925);
  nand NAND2_554(I7174,g2006,I7172);
  nand NAND2_555(I13214,g7065,I13213);
  nand NAND2_556(I10820,g2039,I10818);
  nand NAND2_557(I7239,g1658,g2134);
  nand NAND2_558(I8165,g1943,I8164);
  nand NAND2_559(I7180,g2351,I7179);
  nand NAND2_560(I6103,g849,I6102);
  nand NAND2_561(I8133,g3232,I8132);
  nand NAND2_562(g1819,I5696,I5697);
  nand NAND2_563(I12032,g5918,I12031);
  nand NAND2_564(g5035,I9382,I9383);
  nand NAND2_565(I9954,g2131,I9953);
  nand NAND2_566(I8538,g2798,I8536);
  nand NAND2_567(I15864,g9171,I15862);
  nand NAND2_568(I12871,g6618,I12869);
  nand NAND2_569(g6466,I11615,I11616);
  nand NAND2_570(g7447,I13599,I13600);
  nand NAND2_571(g6165,I10855,I10856);
  nand NAND2_572(g6571,I11758,I11759);
  nand NAND3_10(g5310,g5009,g4335,g4963);
  nand NAND2_573(g4298,I8254,I8255);
  nand NAND2_574(I10743,g5550,g2100);
  nand NAND2_575(g5762,I10360,I10361);
  nand NAND2_576(g3925,I7575,I7576);
  nand NAND2_577(g5590,g2044,g4906);
  nand NAND2_578(I11759,g6118,I11757);
  nand NAND2_579(g5657,g5021,g4381);
  nand NAND2_580(I11758,g1758,I11757);
  nand NAND2_581(g6467,g5956,g5269);
  nand NAND2_582(g5556,I9986,I9987);
  nand NAND2_583(g4219,I8120,I8121);
  nand NAND2_584(g2385,I6258,I6259);
  nand NAND4_2(g7234,g3757,g3739,g7050,g3770);
  nand NAND2_585(g4252,g2276,g3313);
  nand NAND2_586(g3906,I7504,I7505);
  nand NAND2_587(I6775,g2386,I6774);
  nand NAND2_588(I7010,g2295,I7009);
  nand NAND2_589(I10890,g2259,I10888);
  nand NAND2_590(I8605,g2487,g2764);
  nand NAND2_591(g6181,I10907,I10908);
  nand NAND2_592(g4911,g4320,g2044);
  nand NAND2_593(I9475,g4038,g1942);
  nand NAND2_594(I6739,g195,g1970);
  nand NAND2_595(I7172,g1739,g2006);
  nand NAND2_596(I7278,g2497,I7277);
  nand NAND2_597(I11135,g5476,g3052);
  nand NAND2_598(I7618,g1721,I7616);
  nand NAND2_599(g2801,I6539,I6540);
  nand NAND2_600(g5557,I9993,I9994);
  nand NAND2_601(g3907,I7511,I7512);
  nand NAND2_602(I6501,g1537,I6499);
  nand NAND2_603(I13004,g1053,I13002);
  nand NAND2_604(I9276,g2533,g4313);
  nand NAND2_605(g3656,I7139,I7140);
  nand NAND2_606(g3915,I7539,I7540);
  nand NAND2_607(g4399,I8393,I8394);
  nand NAND2_608(I9986,g4836,I9985);
  nand NAND2_609(I7567,g2481,g3780);
  nand NAND2_610(I9277,g2533,I9276);
  nand NAND2_611(I11163,g5469,g3029);
  nand NAND2_612(I12551,g6689,I12550);
  nand NAND2_613(g7121,I12952,I12953);
  nand NAND2_614(I9987,g2096,I9985);
  nand NAND2_615(g3899,I7479,I7480);
  nand NAND2_616(I9547,g1952,g4307);
  nand NAND2_617(I7179,g2351,g795);
  nand NAND2_618(I8326,g2011,g2721);
  nand NAND2_619(I12181,g6163,I12179);
  nand NAND2_620(I10011,g4821,I10009);
  nand NAND2_621(I7611,g3771,I7609);
  nand NAND2_622(I10627,g1514,I10625);
  nand NAND2_623(g4887,I9234,I9235);
  nand NAND2_624(g4228,g1408,g2665);
  nand NAND2_625(I10925,g2752,I10923);
  nand NAND2_626(I6998,g2242,I6996);
  nand NAND2_627(I8327,g2011,I8326);
  nand NAND2_628(g6023,I10626,I10627);
  nand NAND2_629(I7511,g2992,I7510);
  nand NAND2_630(g2333,g985,g990);
  nand NAND2_631(I8472,g2821,I8470);
  nand NAND2_632(I7574,g2999,g1718);
  nand NAND2_633(g9190,I15849,I15850);
  nand NAND2_634(I12870,g2536,I12869);
  nand NAND2_635(I6925,g33,I6923);
  nand NAND2_636(I13395,g7212,g1057);
  nand NAND2_637(g5540,I9954,I9955);
  nand NAND2_638(I10626,g5314,I10625);
  nand NAND2_639(I14245,g7683,I14244);
  nand NAND2_640(I10299,g5461,I10298);
  nand NAND2_641(g3895,I7467,I7468);
  nand NAND2_642(I10298,g5461,g2562);
  nand NAND2_643(g6472,g5971,g5269);
  nand NAND2_644(I6906,g1838,I6904);
  nand NAND2_645(I5599,g1481,I5598);
  nand NAND2_646(I9194,g4252,g1652);
  nand NAND2_647(I10856,g2584,I10854);
  nand NAND2_648(I15882,g9179,I15880);
  nand NAND2_649(I7139,g2404,I7138);
  nand NAND2_650(I9071,g1149,I9069);
  nand NAND2_651(I9242,g2540,I9241);
  nand NAND3_11(g5291,g4344,g5002,g4963);
  nand NAND2_652(I9948,g4905,I9946);
  nand NAND2_653(I8581,g2498,g2777);
  nand NAND2_654(I9955,g4831,I9953);
  nand NAND2_655(g2751,I6500,I6501);
  nand NAND2_656(I6876,g1967,g1910);
  nand NAND2_657(I9769,g1114,I9767);
  nand NAND2_658(I10080,g2256,I10078);
  nand NAND2_659(I10924,g5525,I10923);
  nand NAND2_660(I15849,g9162,I15848);
  nand NAND2_661(g3286,I6905,I6906);
  nand NAND2_662(I15848,g9162,g9154);
  nand NAND2_663(I9993,g2145,I9992);
  nand NAND2_664(I12597,g6582,I12596);
  nand NAND2_665(I5695,g1513,g1524);
  nand NAND2_666(I7444,g2973,I7443);
  nand NAND2_667(I7269,g2486,I7268);
  nand NAND2_668(I10198,g1958,I10196);
  nand NAND2_669(g5594,I10072,I10073);
  nand NAND2_670(I13785,g7427,g1477);
  nand NAND2_671(I6877,g1967,I6876);
  nand NAND2_672(I10868,g2605,I10866);
  nand NAND2_673(g2474,g1405,g1412);
  nand NAND2_674(I12854,g6695,I12852);
  nand NAND2_675(I10225,g4895,I10223);
  nand NAND2_676(I11151,g3038,I11149);
  nand NAND2_677(I11172,g3038,I11170);
  nand NAND2_678(I6064,g852,g883);
  nand NAND2_679(g4893,g2460,g4312);
  nand NAND2_680(g5550,g1879,g4830);
  nand NAND2_681(I14244,g7683,g1065);
  nand NAND2_682(g3900,I7486,I7487);
  nand NAND2_683(g6163,g5633,g3716);
  nand NAND2_684(I7436,g2517,g3822);
  nand NAND2_685(I12550,g6689,g1462);
  nand NAND2_686(g4821,g4220,g3605);
  nand NAND2_687(I6844,g2016,I6842);
  nand NAND2_688(I12596,g6582,g1126);
  nand NAND2_689(I7422,g2525,I7421);
  nand NAND2_690(I13377,g7199,I13376);
  nand NAND2_691(I12180,g1961,I12179);
  nand NAND2_692(I10010,g1949,I10009);
  nand NAND2_693(g3886,I7422,I7423);
  nand NAND2_694(I6814,g210,I6813);
  nand NAND2_695(I10079,g4911,I10078);
  nand NAND2_696(I7437,g2517,I7436);
  nand NAND2_697(g3314,I6917,I6918);
  nand NAND2_698(I10078,g4911,g2256);
  nand NAND3_12(g5312,g5009,g5002,g4963);
  nand NAND2_699(I10322,g2573,I10320);
  nand NAND2_700(g2051,g1444,g1450);
  nand NAND2_701(I10901,g2752,I10899);
  nand NAND2_702(I6918,g1732,I6916);
  nand NAND2_703(I9980,g2092,I9978);
  nand NAND2_704(I9069,g4400,g1149);
  nand NAND2_705(I8583,g2777,I8581);
  nand NAND2_706(g4359,I8327,I8328);
  nand NAND2_707(I10144,g1916,I10142);
  nand NAND2_708(I11551,g1045,I11549);
  nand NAND2_709(g3887,I7429,I7430);
  nand NAND2_710(I7454,g1106,I7452);
  nand NAND2_711(I10336,g2573,I10334);
  nand NAND2_712(g6627,I11874,I11875);
  nand NAND2_713(I7532,g2487,I7531);
  nand NAND2_714(I10017,g4700,g2174);
  nand NAND2_715(I5619,g1092,g1130);
  nand NAND2_716(I13376,g7199,g1472);
  nand NAND2_717(I11103,g2712,I11101);
  nand NAND2_718(I11095,g5515,I11094);
  nand NAND2_719(g8633,g8176,g6232);
  nand NAND2_720(I8503,g2986,I8502);
  nand NAND2_721(g4880,g4287,g1879);
  nand NAND3_13(g5576,g4894,g4888,g4884);
  nand NAND2_722(I10224,g2522,I10223);
  nand NAND2_723(I7429,g3222,I7428);
  nand NAND2_724(I8120,g1904,I8119);
  nand NAND2_725(I12015,g5874,g5847);
  nand NAND2_726(I5598,g1481,g1489);
  nand NAND2_727(g6276,I11116,I11117);
  nand NAND2_728(g4243,I8165,I8166);
  nand NAND2_729(g5747,I10299,I10300);
  nand NAND2_730(I6842,g205,g2016);
  nand NAND2_731(I7138,g2404,g2397);
  nand NAND2_732(I10954,g2340,I10952);
  nand NAND2_733(I6941,g2051,I6939);
  nand NAND2_734(g6503,g5269,g5897);
  nand NAND2_735(I5519,g1087,g1098);
  nand NAND2_736(I12179,g1961,g6163);
  nand NAND2_737(g8681,I14838,I14839);
  nand NAND2_738(I15899,g9203,I15897);
  nand NAND2_739(I15898,g9202,I15897);
  nand NAND2_740(I12953,g1467,I12951);
  nand NAND2_741(I8244,g2011,I8243);
  nand NAND2_742(g6277,I11123,I11124);
  nand NAND2_743(I7575,g2999,I7574);
  nand NAND2_744(I8340,g1698,I8338);
  nand NAND2_745(g4090,I7892,I7893);
  nand NAND2_746(I9768,g4832,I9767);
  nand NAND2_747(g6516,g5897,g5278);
  nand NAND2_748(g3129,I6843,I6844);
  nand NAND2_749(g4456,I8471,I8472);
  nand NAND2_750(I7539,g2996,I7538);
  nand NAND2_751(g2995,I6740,I6741);
  nand NAND2_752(g2294,I6065,I6066);
  nand NAND2_753(g3221,I6877,I6878);
  nand NAND2_754(I7268,g2486,g955);
  nand NAND2_755(I5506,g1532,I5505);
  nand NAND2_756(I7452,g3226,g1106);
  nand NAND2_757(g6709,I12052,I12053);
  nand NAND2_758(I6540,g2557,I6538);
  nand NAND2_759(I10093,g4881,I10092);
  nand NAND2_760(I9195,g4252,I9194);
  nand NAND2_761(I7086,g1753,I7085);
  nand NAND2_762(I7486,g2989,I7485);
  nand NAND2_763(g6435,I11575,I11576);
  nand NAND2_764(g6482,g5269,g5847);
  nand NAND2_765(I7504,g2498,I7503);
  nand NAND2_766(I10875,g2595,I10873);
  nand NAND2_767(I7070,g1643,I7068);
  nand NAND2_768(I14837,g8660,g1073);
  nand NAND2_769(g4686,I8956,I8957);
  nand NAND2_770(I11094,g5515,g2734);
  nand NAND2_771(I5507,g1528,I5505);
  nand NAND2_772(I11150,g5473,I11149);
  nand NAND2_773(I13801,g7429,I13800);
  nand NAND2_774(I9692,g5096,I9691);
  nand NAND2_775(g7444,I13588,I13589);
  nand NAND2_776(I13018,g1142,I13016);
  nand NAND2_777(I6259,g901,I6257);
  nand NAND2_778(I7087,g1918,I7085);
  nand NAND2_779(I7487,g1708,I7485);
  nand NAND2_780(I6923,g1728,g33);
  nand NAND2_781(g3818,I7278,I7279);
  nand NAND2_782(I8394,g1925,I8392);
  nand NAND2_783(I9979,g4880,I9978);
  nand NAND2_784(g3893,I7453,I7454);
  nand NAND2_785(I7445,g1701,I7443);
  nand NAND2_786(I7173,g1739,I7172);
  nand NAND2_787(I8471,g2525,I8470);
  nand NAND2_788(I9828,g1509,I9826);
  nand NAND2_789(g5595,I10079,I10080);
  nand NAND2_790(I8955,g4246,g1110);
  nand NAND2_791(g9192,I15863,I15864);
  nand NAND2_792(I8254,g2454,I8253);
  nand NAND2_793(I10836,g2584,I10834);
  nand NAND2_794(I9746,g4826,I9745);
  nand NAND2_795(I7459,g2506,g3815);
  nand NAND2_796(I11102,g5491,I11101);
  nand NAND2_797(I11157,g5482,I11156);
  nand NAND2_798(g3939,I7617,I7618);
  nand NAND2_799(I8150,g3229,g38);
  nand NAND2_800(g3083,I6814,I6815);
  nand NAND2_801(I9953,g2131,g4831);
  nand NAND4_3(g4879,g2595,g2584,g4270,g4281);
  nand NAND2_802(I10313,g5484,g1041);
  nand NAND2_803(I6065,g852,I6064);
  nand NAND2_804(I10305,g5470,g3019);
  nand NAND2_805(I10900,g5520,I10899);
  nand NAND2_806(I9747,g1549,I9745);
  nand NAND2_807(g8627,g6232,g8091);
  nand NAND2_808(I11550,g5984,I11549);
  nand NAND2_809(I9241,g2540,g4305);
  nand NAND2_810(g5512,g1879,g4877);
  nand NAND2_811(I7188,g1834,I7186);
  nand NAND2_812(I10874,g5516,I10873);
  nand NAND2_813(I7216,g2091,I7214);
  nand NAND2_814(I12952,g7003,I12951);
  nand NAND2_815(I7428,g3222,g1541);
  nand NAND2_816(I10009,g1949,g4821);
  nand NAND2_817(I7430,g1541,I7428);
  nand NAND2_818(I11156,g5482,g3052);
  nand NAND2_819(I9152,g3883,I9151);
  nand NAND2_820(I5621,g1130,I5619);
  nand NAND2_821(I6815,g2052,I6813);
  nand NAND2_822(g4905,g4282,g3533);
  nand NAND2_823(g3811,I7269,I7270);
  nand NAND2_824(g3315,I6924,I6925);
  nand NAND2_825(I10907,g5492,I10906);
  nand NAND2_826(I7609,g2471,g3771);
  nand NAND2_827(I12834,g6709,I12832);
  nand NAND2_828(I8392,g2949,g1925);
  nand NAND2_829(I9170,g1935,I9169);
  nand NAND2_830(I15889,g9191,I15887);
  nor NOR4_0(g4884,g4492,g4476,g4456,g4294);
  nor NOR3_0(g8656,g8199,I14758,I14759);
  nor NOR2_0(g3260,g1728,g2490);
  nor NOR2_1(g5615,g4714,g3002);
  nor NOR3_1(g8236,g8199,I14495,I14496);
  nor NOR2_2(g4160,g1231,g2834);
  nor NOR2_3(g7406,g7191,g1600);
  nor NOR2_4(g6259,g3002,g5312);
  nor NOR4_1(g6465,g5403,g5802,g5769,g5790);
  nor NOR4_2(g3515,g1388,g2262,g2230,g2214);
  nor NOR3_2(g8812,g8443,g8421,I15086);
  nor NOR2_5(g3528,g2343,g1391);
  nor NOR2_6(g8073,g7658,g7654);
  nor NOR2_7(g3555,g2359,g1398);
  nor NOR3_3(g8819,g8443,g8421,I15113);
  nor NOR3_4(g8694,g7658,g8613,g7634);
  nor NOR3_5(g8806,g8443,g8421,I15044);
  nor NOR3_6(g8230,g8199,I14467,I14468);
  nor NOR3_7(g8807,g8443,g8421,I15055);
  nor NOR4_3(g4888,g4548,g4528,g4513,g4502);
  nor NOR3_8(g8859,g8493,g8239,I15165);
  nor NOR2_8(g7326,g7194,g6999);
  nor NOR3_9(g8699,g7658,g8613,g7634);
  nor NOR3_10(g8855,g7658,g8613,g7634);
  nor NOR2_9(g8644,g4146,g8128);
  nor NOR2_10(g6193,g1926,g5310);
  nor NOR3_11(g8818,g8443,g8421,I15102);
  nor NOR2_11(g3885,g3310,g3466);
  nor NOR2_12(g6174,g1855,g5305);
  nor NOR2_13(g3233,g1714,g1459);
  nor NOR3_12(g8811,g8443,g8421,I15075);
  nor NOR2_14(g8629,g6270,g8009);
  nor NOR4_4(g8279,g7658,g7616,g8082,g7634);
  nor NOR4_5(g3504,g1375,g2229,g2213,g2206);
  nor NOR4_6(g8625,g1000,g6573,g1860,g8009);
  nor NOR3_13(g8232,g8199,I14479,I14480);
  nor NOR3_14(g8659,g8199,I14771,I14772);
  nor NOR2_15(g6209,g2332,g5305);
  nor NOR4_7(g8630,g6110,g7784,g3591,g1864);
  nor NOR2_16(g6184,g875,g5291);
  nor NOR3_15(g8655,g8199,I14753,I14754);
  nor NOR2_17(g5772,g5428,g1888);
  nor NOR2_18(g2521,g65,g62);
  nor NOR2_19(g7324,g7189,g6994);
  nor NOR4_8(g5023,g3894,g3889,g3886,g4359);
  nor NOR4_9(g8360,g7658,g7616,g8082,g7634);
  nor NOR4_10(g8641,g6559,g162,g7784,g3591);
  nor NOR2_20(g3505,g2263,g1395);
  nor NOR3_16(g8658,g8199,I14766,I14767);
  nor NOR3_17(g8680,g8493,g8239,I14834);
  nor NOR3_18(g4894,g4298,g4575,g4563);
  nor NOR2_21(g7314,g7180,g6972);
  nor NOR4_11(g8092,g7634,g7628,g7616,g7611);
  nor NOR2_22(g7322,g7188,g6991);
  nor NOR4_12(g8523,g7658,g7616,g8082,g7634);
  nor NOR2_23(g7312,g7178,g6970);
  nor NOR2_24(g6452,g6270,g2245);
  nor NOR2_25(g2014,g1421,g1416);
  nor NOR3_19(g8862,g8493,g8239,I15172);
  nor NOR2_26(g6185,g5305,g1590);
  nor NOR3_20(g8679,g8493,g8239,I14831);
  nor NOR4_13(g5039,g3924,g3914,g3906,g3899);
  nor NOR3_21(g8805,g8443,g8421,I15033);
  nor NOR3_22(g7152,g6253,g7083,g5418);
  nor NOR3_23(g6664,g5836,g1901,g1788);
  nor NOR2_27(g1980,g1430,g1431);
  nor NOR3_24(g8233,g8199,I14484,I14485);
  nor NOR3_25(g8706,g7658,g8613,g7634);
  nor NOR4_14(g6910,g1011,g1837,g6559,g1008);
  nor NOR3_26(g8707,g7658,g8613,g7634);
  nor NOR2_28(g7328,g7196,g7001);
  nor NOR2_29(g3516,g2282,g1401);
  nor NOR4_15(g6197,g875,g866,g1590,g5291);
  nor NOR2_30(g8635,g1034,g8128);
  nor NOR2_31(g8801,g8635,g3790);
  nor NOR2_32(g3310,g936,g2557);
  nor NOR2_33(g7318,g7185,g6979);
  nor NOR2_34(g7321,g7187,g6990);
  nor NOR3_27(g3237,g1444,g1838,g1454);
  nor NOR3_28(g8861,g8493,g8239,I15169);
  nor NOR2_35(g4354,g1424,g3541);
  nor NOR3_29(g8803,g8443,g8421,I15021);
  nor NOR2_36(g4676,g3885,g3094);
  nor NOR3_30(g8847,g8493,g8239,I15147);
  nor NOR2_37(g4349,g2496,g3310);
  nor NOR3_31(g3225,g1021,g1025,g1889);
  nor NOR2_38(g7566,g7421,g1597);
  nor NOR3_32(g8863,g8493,g8239,I15175);
  nor NOR2_39(g1964,g1428,g1429);
  nor NOR3_33(g7209,g1789,g146,g6984);
  nor NOR3_34(g5614,g3002,g1590,g4714);
  nor NOR2_40(g4318,g3681,g1590);
  nor NOR2_41(g6214,g878,g5284);
  nor NOR2_42(g4232,g1934,g3591);
  nor NOR3_35(g6489,g5802,g5769,g5790);
  nor NOR3_36(g3790,g985,g990,g2295);
  nor NOR3_37(g5056,g3556,g2872,g3938);
  nor NOR3_38(g8850,g8493,g8239,I15152);

endmodule

