
module c1908(N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34,
     N37, N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76,
     N79, N82, N85, N88, N91, N94, N99, N104, N2753, N2754, N2755,
     N2756, N2762, N2767, N2768, N2779, N2780, N2781, N2782, N2783,
     N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888, N2889,
     N2890, N2891, N2892, N2899);
//   input N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37,
       N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79,
       N82, N85, N88, N91, N94, N99, N104;
//   output N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780,
       N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886,
       N2887, N2888, N2889, N2890, N2891, N2892, N2899;
  wire N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37,
       N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79,
       N82, N85, N88, N91, N94, N99, N104;
  wire N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780,
       N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886,
       N2887, N2888, N2889, N2890, N2891, N2892, N2899;
  wire N190, N194, N197, N201, N206, N209, N212, N216;
  wire N220, N225, N229, N232, N235, N239, N243, N247;
  wire N251, N252, N253, N263, N266, N269, N272, N275;
  wire N277, N280, N290, N306, N550, N574, N586, N592;
  wire N601, N602, N603, N608, N612, N643, N655, N682;
  wire N685, N724, N886, N887, N893, N896, N899, N903;
  wire N907, N910, N921, N922, N923, N926, N991, N1054;
  wire N1055, N1063, N1064, N1067, N1068, N1119, N1120, N1121;
  wire N1122, N1128, N1129, N1130, N1131, N1132, N1133, N1150;
  wire N1155, N1157, N1158, N1159, N1160, N1162, N1163, N1167;
  wire N1171, N1188, N1206, N1210, N1214, N1221, N1226, N1232;
  wire N1235, N1243, N1246, N1249, N1264, N1267, N1309, N1311;
  wire N1313, N1315, N1317, N1319, N1334, N1344, N1345, N1346;
  wire N1348, N1350, N1352, N1358, N1364, N1370, N1376, N1386;
  wire N1387, N1388, N1389, N1396, N1397, N1398, N1399, N1412;
  wire N1433, N1434, N1438, N1439, N1440, N1443, N1444, N1447;
  wire N1448, N1453, N1454, N1457, N1458, N1459, N1460, N1462;
  wire N1464, N1472, N1478, N1481, N1484, N1487, N1489, N1493;
  wire N1495, N1496, N1498, N1510, N1513, N1517, N1521, N1526;
  wire N1527, N1528, N1529, N1530, N1531, N1532, N1546, N1554;
  wire N1557, N1561, N1567, N1568, N1571, N1576, N1594, N1596;
  wire N1636, N1638, N1671, N1672, N1678, N1685, N1688, N1706;
  wire N1708, N1712, N1720, N1723, N1740, N1741, N1742, N1746;
  wire N1748, N1759, N1769, N1772, N1773, N1774, N1784, N1788;
  wire N1795, N1796, N1798, N1801, N1802, N1809, N1821, N1822;
  wire N1825, N1826, N1827, N1830, N1838, N1848, N1850, N1852;
  wire N1855, N1857, N1858, N1878, N1882, N1883, N1884, N1885;
  wire N1889, N1898, N1910, N1911, N1912, N1913, N1915, N1919;
  wire N1920, N1936, N1938, N1941, N1947, N1965, N1968, N1975;
  wire N1976, N1979, N1987, N2000, N2003, N2004, N2005, N2008;
  wire N2012, N2014, N2016, N2018, N2019, N2020, N2022, N2023;
  wire N2024, N2026, N2036, N2038, N2040, N2041, N2047, N2052;
  wire N2055, N2060, N2062, N2067, N2076, N2077, N2078, N2081;
  wire N2104, N2119, N2129, N2143, N2214, N2215, N2222, N2223;
  wire N2226, N2227, N2230, N2232, N2234, N2236, N2240, N2244;
  wire N2250, N2253, N2256, N2266, N2272, N2279, N2340, N2353;
  wire N2361, N2375, N2384, N2385, N2386, N2426, N2427, N2537;
  wire N2540, N2543, N2546, N2549, N2552, N2555, N2558, N2561;
  wire N2564, N2567, N2570, N2573, N2576, N2594, N2597, N2600;
  wire N2603, N2606, N2611, N2614, N2617, N2620, N2627, N2628;
  wire N2629, N2630, N2631, N2632, N2633, N2634, N2639, N2642;
  wire N2645, N2648, N2651, N2655, N2658, N2661, N2664, N2669;
  wire N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2682;
  wire N2683, N2688, N2689, N2690, N2691, N2720, N2721, N2722;
  wire N2723, N2724, N2725, N2726, N2727, N2728, N2729, N2730;
  wire N2731, N2732, N2733, N2734, N2735, N2736, N2737, N2738;
  wire N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746;
  wire N2747, N2750, N2757, N2758, N2759, N2760, N2761, N2763;
  wire N2764, N2765, N2766, N2773, N2776, N2789, N2800, N2807;
  wire N2808, N2809, N2810, N2812, N2815, N2818, N2821, N2824;
  wire N2827, N2828, N2829, N2843, N2846, N2850, N2851, N2852;
  wire N2853, N2854, N2857, N2858, N2859, N2860, N2861, N2862;
  wire N2863, N2866, N2867, N2868, N2869, N2870, N2871, N2872;
  wire N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880;
  wire N2881, N2882, N2883, N2895, N2896, N2897, N2898, n_59;
  wire n_66, n_71, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86;
  and AND2_87 (N574, N63, N275);
  and AND2_91 (N586, N66, N275);
  and AND2_123 (N682, N251, N104);
  and AND2_124 (N685, N252, N104);
  and AND2_594 (N1965, N1910, N601);
  and AND2_595 (N1968, N602, N1912);
  and AND2_653 (N2104, N2012, N2047);
  and AND2_654 (N2119, N1979, N2047);
  and AND2_655 (N2129, N2012, N2026);
  and AND2_656 (N2143, N1979, N2026);
  and AND2_693 (N2266, N899, N2240);
  and AND2_695 (N2272, N903, N2244);
  and AND2_701 (N2340, N2067, N2250);
  and AND2_702 (N2353, N2041, N2250);
  and AND2_703 (N2361, N2067, N2236);
  and AND2_704 (N2375, N2041, N2236);
  and AND2_706 (N2385, N1163, N2253);
  and AND2_707 (N2386, N899, N2253);
  and AND2_708 (N2426, N1167, N2256);
  and AND2_709 (N2427, N903, N2256);
  and AND2_810 (N2773, N2745, N275);
  and AND2_811 (N2776, N2746, N275);
  and AND2_869 (N2886, N2876, N550);
  and AND2_870 (N2887, N550, N2877);
  and AND2_871 (N2888, N550, N2878);
  and AND2_872 (N2889, N2879, N550);
  and AND2_873 (N2890, N550, N2880);
  and AND2_880 (N2899, N2898, N550);
  and AND3_93 (N592, N49, N253, N275);
  and AND3_110 (N643, N56, N69, N275);
  and AND3_114 (N655, N60, N69, N275);
  and AND3_137 (N724, N53, N253, N275);
  and AND3_175 (N926, N99, N275, N603);
  and AND3_830 (N2815, N76, N94, N2789);
  and AND3_831 (N2818, N82, N94, N2789);
  and AND3_832 (N2821, N85, N94, N2789);
  and AND3_836 (N2829, N79, N94, N2789);
  nand NAND2_17 (N251, N63, N88);
  nand NAND2_18 (N252, N66, N91);
  nand NAND2_75 (N550, N306, N104);
  nand NAND2_96 (N601, N104, N277);
  nand NAND2_97 (N602, N104, N280);
  nand NAND2_98 (N603, N69, N72);
  nand NAND2_99 (N608, N69, N290);
  nand NAND2_100 (N612, N253, N290);
  nand NAND2_160 (N899, N53, N612);
  nand NAND2_161 (N903, N60, N608);
  nand NAND2_162 (N907, N49, N612);
  nand NAND2_163 (N910, N56, N608);
  nand NAND2_233 (N1054, N216, N10);
  nand NAND2_234 (N1055, N201, N22);
  nand NAND2_235 (N1063, N239, N25);
  nand NAND2_236 (N1064, N220, N40);
  nand NAND2_237 (N1067, N655, N37);
  nand NAND2_238 (N1068, N235, N896);
  nand NAND2_239 (N1119, N216, N13);
  nand NAND2_240 (N1120, N206, N22);
  nand NAND2_241 (N1121, N243, N991);
  nand NAND2_242 (N1122, N724, N43);
  nand NAND2_243 (N1128, N216, N16);
  nand NAND2_244 (N1129, N209, N22);
  nand NAND2_245 (N1130, N243, N28);
  nand NAND2_246 (N1131, N225, N43);
  nand NAND2_247 (N1132, N225, N19);
  nand NAND2_248 (N1133, N212, N28);
  nand NAND2_251 (N1150, N1054, N1055);
  nand NAND2_259 (N1158, N1063, N1064);
  nand NAND2_261 (N1160, N592, N1);
  nand NAND2_263 (N1162, N1067, N1068);
  nand NAND2_268 (N1171, N921, N923);
  nand NAND2_269 (N1188, N922, N923);
  nand NAND2_271 (N1206, N194, N7);
  nand NAND2_275 (N1210, N209, N19);
  nand NAND2_279 (N1214, N243, N46);
  nand NAND2_286 (N1221, N232, N37);
  nand NAND2_291 (N1226, N239, N10);
  nand NAND2_297 (N1232, N1119, N1120);
  nand NAND2_298 (N1235, N1121, N1122);
  nand NAND2_304 (N1243, N1128, N1129);
  nand NAND2_305 (N1246, N1130, N1131);
  nand NAND2_306 (N1249, N1132, N1133);
  nand NAND2_312 (N1267, N190, N1159);
  nand NAND2_313 (N1309, N197, N4);
  nand NAND2_315 (N1311, N212, N16);
  nand NAND2_317 (N1313, N247, N43);
  nand NAND2_319 (N1315, N235, N34);
  nand NAND2_321 (N1317, N201, N40);
  nand NAND2_328 (N1344, N1267, N1160);
  nand NAND2_329 (N1345, N1249, N10);
  nand NAND2_335 (N1352, N1309, N1206);
  nand NAND2_337 (N1358, N1311, N1210);
  nand NAND2_339 (N1364, N1313, N1214);
  nand NAND2_341 (N1370, N1315, N1221);
  nand NAND2_343 (N1376, N1317, N1226);
  nand NAND2_347 (N1387, N1232, N4);
  nand NAND2_349 (N1389, N1235, N31);
  nand NAND2_353 (N1397, N1243, N7);
  nand NAND2_355 (N1399, N1246, N34);
  nand NAND2_357 (N1412, N201, N1346);
  nand NAND2_361 (N1433, N194, N1386);
  nand NAND2_362 (N1434, N229, N1388);
  nand NAND2_363 (N1438, N197, N1396);
  nand NAND2_364 (N1439, N232, N1398);
  nand NAND2_366 (N1443, N1352, N1);
  nand NAND2_370 (N1447, N1358, N13);
  nand NAND2_374 (N1453, N1364, N28);
  nand NAND2_378 (N1457, N1370, N31);
  nand NAND2_380 (N1459, N1376, N1157);
  nand NAND2_383 (N1462, N1158, N46);
  nand NAND2_385 (N1464, N1345, N1412);
  nand NAND2_390 (N1472, N1387, N1433);
  nand NAND2_393 (N1478, N1389, N1434);
  nand NAND2_394 (N1481, N1399, N1439);
  nand NAND2_395 (N1484, N1397, N1438);
  nand NAND2_396 (N1487, N190, N1444);
  nand NAND2_398 (N1489, N206, N1448);
  nand NAND2_402 (N1493, N225, N1454);
  nand NAND2_404 (N1495, N229, N1458);
  nand NAND2_405 (N1496, N586, N1460);
  nand NAND2_406 (N1498, N247, N1319);
  nand NAND2_412 (N1513, N1443, N1487);
  nand NAND2_414 (N1517, N1447, N1489);
  nand NAND2_416 (N1521, N1453, N1493);
  nand NAND2_418 (N1526, N1457, N1495);
  nand NAND2_419 (N1527, N1459, N1496);
  nand NAND2_421 (N1529, N1462, N1498);
  nand NAND2_432 (N1567, N1484, N1531);
  nand NAND2_433 (N1568, N1481, N1532);
  nand NAND2_440 (N1594, N1529, N1530);
  nand NAND2_442 (N1596, N1567, N1568);
  nand NAND2_452 (N1636, N1478, N1576);
  nand NAND2_453 (N1638, N1576, N1464);
  nand NAND2_462 (N1671, N1596, N893);
  nand NAND2_466 (N1678, N1521, N25);
  nand NAND2_472 (N1685, N1594, N1636);
  nand NAND2_473 (N1688, N1510, N1529);
  nand NAND2_476 (N1706, N643, N1672);
  nand NAND2_478 (N1708, N1546, N1561);
  nand NAND2_482 (N1712, N220, N1554);
  nand NAND2_486 (N1720, N1554, N1557);
  nand NAND2_488 (N1723, N1638, N1688);
  nand NAND2_494 (N1740, N1685, N1528);
  nand NAND2_496 (N1742, N1671, N1706);
  nand NAND2_497 (N1746, N1517, N1513);
  nand NAND2_499 (N1748, N1678, N1712);
  nand NAND2_501 (N1759, N1526, N1521);
  nand NAND2_507 (N1769, N1472, N1741);
  nand NAND2_508 (N1772, N1723, N1162);
  nand NAND2_510 (N1774, N1708, N1746);
  nand NAND2_513 (N1784, N1554, N1546);
  nand NAND2_517 (N1788, N1720, N1759);
  nand NAND2_520 (N1795, N1748, N1155);
  nand NAND2_522 (N1798, N1740, N1769);
  nand NAND2_523 (N1801, N1334, N1773);
  nand NAND2_524 (N1802, N1742, N290);
  nand NAND2_527 (N1809, N1513, N1521);
  nand NAND2_532 (N1821, N1774, N1150);
  nand NAND2_536 (N1825, N574, N1796);
  nand NAND2_537 (N1826, N1788, N1158);
  nand NAND2_539 (N1830, N1772, N1801);
  nand NAND2_541 (N1838, N1809, N1784);
  nand NAND2_543 (N1848, N1264, N1822);
  nand NAND2_545 (N1850, N1795, N1825);
  nand NAND2_546 (N1852, N1319, N1827);
  nand NAND2_547 (N1855, N1788, N1517);
  nand NAND2_550 (N1858, N1798, N290);
  nand NAND2_557 (N1878, N1821, N1848);
  nand NAND2_559 (N1882, N1838, N1526);
  nand NAND2_561 (N1884, N1826, N1852);
  nand NAND2_562 (N1885, N1561, N1827);
  nand NAND2_563 (N1889, N1830, N290);
  nand NAND2_570 (N1911, N1557, N1883);
  nand NAND2_572 (N1913, N1855, N1885);
  nand NAND2_574 (N1919, N1802, N85);
  nand NAND2_583 (N1936, N1882, N1911);
  nand NAND2_586 (N1941, N272, N1920);
  nand NAND2_596 (N1975, N1858, N82);
  nand NAND2_600 (N1979, N1919, N1941);
  nand NAND2_605 (N2000, N1878, N1850);
  nand NAND2_607 (N2003, N1947, N1344);
  nand NAND2_608 (N2004, N1889, N1350);
  nand NAND2_612 (N2008, N269, N1976);
  nand NAND2_616 (N2014, N1878, N1898);
  nand NAND2_618 (N2016, N1936, N1527);
  nand NAND2_621 (N2020, N1898, N1910);
  nand NAND2_623 (N2022, N1987, N1571);
  nand NAND2_624 (N2023, N1440, N1913);
  nand NAND2_625 (N2024, N910, N2005);
  nand NAND2_627 (N2026, N1975, N2008);
  nand NAND2_631 (N2036, N1850, N1910);
  nand NAND2_633 (N2038, N2020, N2000);
  nand NAND2_635 (N2040, N2023, N2003);
  nand NAND2_636 (N2041, N2004, N2024);
  nand NAND2_639 (N2052, N2036, N2014);
  nand NAND2_640 (N2055, N2022, N2016);
  nand NAND2_643 (N2062, N2040, N290);
  nand NAND2_649 (N2078, N2060, N290);
  nand NAND2_650 (N2081, N2055, N290);
  nand NAND2_663 (N2214, N2062, N79);
  nand NAND2_667 (N2222, N2078, N1348);
  nand NAND2_671 (N2226, N2081, N76);
  nand NAND2_675 (N2230, N266, N2215);
  nand NAND2_677 (N2232, N907, N2223);
  nand NAND2_679 (N2234, N263, N2227);
  nand NAND2_681 (N2236, N2214, N2230);
  nand NAND2_683 (N2240, N2222, N2232);
  nand NAND2_685 (N2244, N2226, N2234);
  nand NAND2_750 (N2669, N2558, N190);
  nand NAND2_752 (N2671, N2561, N194);
  nand NAND2_754 (N2673, N2564, N197);
  nand NAND2_756 (N2675, N2567, N201);
  nand NAND2_758 (N2682, N2570, N225);
  nand NAND2_760 (N2688, N2573, N243);
  nand NAND2_762 (N2690, N2576, N247);
  nand NAND2_765 (N2720, N1, N2670);
  nand NAND2_766 (N2721, N4, N2672);
  nand NAND2_767 (N2722, N7, N2674);
  nand NAND2_768 (N2723, N10, N2676);
  nand NAND2_769 (N2724, N2639, N206);
  nand NAND2_771 (N2726, N2642, N209);
  nand NAND2_773 (N2728, N2645, N212);
  nand NAND2_775 (N2730, N2648, N216);
  nand NAND2_777 (N2732, N2651, N220);
  nand NAND2_779 (N2734, N28, N2683);
  nand NAND2_780 (N2735, N2655, N229);
  nand NAND2_782 (N2737, N2658, N232);
  nand NAND2_784 (N2739, N2661, N235);
  nand NAND2_786 (N2741, N2664, N239);
  nand NAND2_788 (N2743, N43, N2689);
  nand NAND2_789 (N2744, N46, N2691);
  nand NAND2_794 (N2753, N2669, N2720);
  nand NAND2_795 (N2754, N2671, N2721);
  nand NAND2_796 (N2755, N2673, N2722);
  nand NAND2_797 (N2756, N2675, N2723);
  nand NAND2_798 (N2757, N13, N2725);
  nand NAND2_799 (N2758, N16, N2727);
  nand NAND2_800 (N2759, N19, N2729);
  nand NAND2_801 (N2760, N22, N2731);
  nand NAND2_802 (N2761, N25, N2733);
  nand NAND2_803 (N2762, N2682, N2734);
  nand NAND2_804 (N2763, N31, N2736);
  nand NAND2_805 (N2764, N34, N2738);
  nand NAND2_806 (N2765, N37, N2740);
  nand NAND2_807 (N2766, N40, N2742);
  nand NAND2_808 (N2767, N2688, N2743);
  nand NAND2_809 (N2768, N2690, N2744);
  nand NAND2_812 (N2779, N2724, N2757);
  nand NAND2_813 (N2780, N2726, N2758);
  nand NAND2_814 (N2781, N2728, N2759);
  nand NAND2_815 (N2782, N2730, N2760);
  nand NAND2_816 (N2783, N2732, N2761);
  nand NAND2_817 (N2784, N2735, N2763);
  nand NAND2_818 (N2785, N2737, N2764);
  nand NAND2_819 (N2786, N2739, N2765);
  nand NAND2_820 (N2787, N2741, N2766);
  nand NAND2_822 (N2789, N2747, N2750);
  nand NAND2_824 (N2807, N2773, N2018);
  nand NAND2_826 (N2809, N2776, N2019);
  nand NAND2_834 (N2827, N1965, N2808);
  nand NAND2_835 (N2828, N1968, N2810);
  nand NAND2_837 (N2843, N2807, N2827);
  nand NAND2_838 (N2846, N2809, N2828);
  nand NAND2_839 (N2850, N2812, N2076);
  nand NAND2_840 (N2851, N2815, N2077);
  nand NAND2_841 (N2852, N2818, N1915);
  nand NAND2_842 (N2853, N2821, N1857);
  nand NAND2_843 (N2854, N2824, N1938);
  nand NAND2_850 (N2863, N2829, N1947);
  nand NAND2_851 (N2866, N2052, N2857);
  nand NAND2_852 (N2867, N2055, N2858);
  nand NAND2_853 (N2868, N1798, N2859);
  nand NAND2_854 (N2869, N1742, N2860);
  nand NAND2_855 (N2870, N1830, N2861);
  nand NAND2_856 (N2871, N2843, N886);
  nand NAND2_858 (N2873, N2846, N887);
  nand NAND2_860 (N2875, N1913, N2862);
  nand NAND2_861 (N2876, N2866, N2850);
  nand NAND2_862 (N2877, N2867, N2851);
  nand NAND2_863 (N2878, N2868, N2852);
  nand NAND2_864 (N2879, N2869, N2853);
  nand NAND2_865 (N2880, N2870, N2854);
  nand NAND2_866 (N2881, N682, N2872);
  nand NAND2_867 (N2882, N685, N2874);
  nand NAND2_868 (N2883, N2875, N2863);
  nand NAND2_874 (N2891, N2871, N2881);
  nand NAND2_875 (N2892, N2873, N2882);
  nand NAND2_876 (N2895, N2883, N1440);
  nand NAND2_878 (N2897, N1344, N2896);
  nand NAND2_879 (N2898, N2895, N2897);
  nand NAND4_172 (N921, N277, N94, N104, N603);
  nand NAND4_173 (N922, N280, N94, N104, N603);
  nand NAND5_710 (N2537, N2266, N2272, N2361, N2104, N1171);
  nand NAND5_711 (N2540, N2266, N2272, N2340, N2129, N1171);
  nand NAND5_712 (N2543, N2266, N2272, N2340, N2119, N1171);
  nand NAND5_713 (N2546, N2266, N2272, N2353, N2104, N1171);
  nand NAND5_714 (N2549, N2266, N2272, N2375, N2119, N1188);
  nand NAND5_715 (N2552, N2266, N2272, N2361, N2143, N1188);
  nand NAND5_716 (N2555, N2266, N2272, N2375, N2129, N1188);
  nand NAND5_724 (N2594, N2266, N2427, N2361, N2129, N1171);
  nand NAND5_725 (N2597, N2266, N2427, N2361, N2119, N1171);
  nand NAND5_726 (N2600, N2266, N2427, N2375, N2104, N1171);
  nand NAND5_727 (N2603, N2266, N2427, N2340, N2143, N1171);
  nand NAND5_728 (N2606, N2266, N2427, N2353, N2129, N1188);
  nand NAND5_729 (N2611, N2386, N2272, N2361, N2129, N1188);
  nand NAND5_730 (N2614, N2386, N2272, N2361, N2119, N1188);
  nand NAND5_731 (N2617, N2386, N2272, N2375, N2104, N1188);
  nand NAND5_732 (N2620, N2386, N2272, N2353, N2129, N1188);
  nand NAND5_733 (N2627, N2266, N2427, N2340, N2104, N926);
  nand NAND5_734 (N2628, N2386, N2272, N2340, N2104, N926);
  nand NAND5_735 (N2629, N2386, N2427, N2361, N2104, N926);
  nand NAND5_736 (N2630, N2386, N2427, N2340, N2129, N926);
  nand NAND5_737 (N2631, N2386, N2427, N2340, N2119, N926);
  nand NAND5_738 (N2632, N2386, N2427, N2353, N2104, N926);
  nand NAND5_739 (N2633, N2386, N2426, N2340, N2104, N926);
  nand NAND5_740 (N2634, N2385, N2427, N2340, N2104, N926);
  nand NAND8_696 (N2279, N2067, N2012, N2047, N2250, N899, N2256,
       N2253, N903);
  nand NAND8_790 (N2745, N2537, N2540, N2543, N2546, N2594, N2597,
       N2600, N2603);
  nand NAND8_791 (N2746, N2606, N2549, N2611, N2614, N2617, N2620,
       N2552, N2555);
  nor NOR2_828 (N2811, N2384, N2800);
  not NOT1_1 (N190, N1);
  not NOT1_2 (N194, N4);
  not NOT1_3 (N197, N7);
  not NOT1_4 (N201, N10);
  not NOT1_5 (N206, N13);
  not NOT1_6 (N209, N16);
  not NOT1_7 (N212, N19);
  not NOT1_8 (N216, N22);
  not NOT1_9 (N220, N25);
  not NOT1_10 (N225, N28);
  not NOT1_11 (N229, N31);
  not NOT1_12 (N232, N34);
  not NOT1_13 (N235, N37);
  not NOT1_14 (N239, N40);
  not NOT1_15 (N243, N43);
  not NOT1_16 (N247, N46);
  not NOT1_19 (N253, N72);
  not NOT1_23 (N263, N76);
  not NOT1_24 (N266, N79);
  not NOT1_25 (N269, N82);
  not NOT1_26 (N272, N85);
  not NOT1_27 (N275, N104);
  not NOT1_29 (N277, N88);
  not NOT1_30 (N280, N91);
  not NOT1_32 (N290, N94);
  not NOT1_36 (N306, N99);
  not NOT1_147 (N886, N682);
  not NOT1_148 (N887, N685);
  not NOT1_154 (N893, N643);
  not NOT1_157 (N896, N655);
  not NOT1_204 (N991, N724);
  not NOT1_256 (N1155, N574);
  not NOT1_258 (N1157, N586);
  not NOT1_260 (N1159, N592);
  not NOT1_264 (N1163, N899);
  not NOT1_266 (N1167, N903);
  not NOT1_311 (N1264, N1150);
  not NOT1_323 (N1319, N1158);
  not NOT1_327 (N1334, N1162);
  not NOT1_330 (N1346, N1249);
  not NOT1_331 (N1348, N907);
  not NOT1_333 (N1350, N910);
  not NOT1_346 (N1386, N1232);
  not NOT1_348 (N1388, N1235);
  not NOT1_352 (N1396, N1243);
  not NOT1_354 (N1398, N1246);
  not NOT1_365 (N1440, N1344);
  not NOT1_367 (N1444, N1352);
  not NOT1_371 (N1448, N1358);
  not NOT1_375 (N1454, N1364);
  not NOT1_379 (N1458, N1370);
  not NOT1_381 (N1460, N1376);
  not NOT1_411 (N1510, N1464);
  not NOT1_420 (N1528, N1472);
  not NOT1_422 (N1530, N1478);
  not NOT1_423 (N1531, N1481);
  not NOT1_424 (N1532, N1484);
  not NOT1_428 (N1546, N1513);
  not NOT1_429 (N1554, N1521);
  not NOT1_430 (N1557, N1526);
  not NOT1_431 (N1561, N1517);
  not NOT1_435 (N1571, N1527);
  not NOT1_436 (N1576, N1529);
  not NOT1_463 (N1672, N1596);
  not NOT1_495 (N1741, N1685);
  not NOT1_509 (N1773, N1723);
  not NOT1_521 (N1796, N1748);
  not NOT1_533 (N1822, N1774);
  not NOT1_538 (N1827, N1788);
  not NOT1_549 (N1857, N1742);
  not NOT1_560 (N1883, N1838);
  not NOT1_567 (N1898, N1850);
  not NOT1_569 (N1910, N1878);
  not NOT1_571 (N1912, N1884);
  not NOT1_573 (N1915, N1798);
  not NOT1_575 (N1920, N1802);
  not NOT1_585 (N1938, N1830);
  not NOT1_589 (N1947, N1913);
  not NOT1_597 (N1976, N1858);
  not NOT1_603 (N1987, N1936);
  not NOT1_609 (N2005, N1889);
  not NOT1_614 (N2012, N1979);
  not NOT1_619 (N2018, N1965);
  not NOT1_620 (N2019, N1968);
  not NOT1_638 (N2047, N2026);
  not NOT1_641 (N2060, N2038);
  not NOT1_644 (N2067, N2041);
  not NOT1_647 (N2076, N2052);
  not NOT1_648 (N2077, N2055);
  not NOT1_664 (N2215, N2062);
  not NOT1_668 (N2223, N2078);
  not NOT1_672 (N2227, N2081);
  not NOT1_687 (N2250, N2236);
  not NOT1_688 (N2253, N2240);
  not NOT1_689 (N2256, N2244);
  not NOT1_751 (N2670, N2558);
  not NOT1_753 (N2672, N2561);
  not NOT1_755 (N2674, N2564);
  not NOT1_757 (N2676, N2567);
  not NOT1_759 (N2683, N2570);
  not NOT1_761 (N2689, N2573);
  not NOT1_763 (N2691, N2576);
  not NOT1_770 (N2725, N2639);
  not NOT1_772 (N2727, N2642);
  not NOT1_774 (N2729, N2645);
  not NOT1_776 (N2731, N2648);
  not NOT1_778 (N2733, N2651);
  not NOT1_781 (N2736, N2655);
  not NOT1_783 (N2738, N2658);
  not NOT1_785 (N2740, N2661);
  not NOT1_787 (N2742, N2664);
  not NOT1_825 (N2808, N2773);
  not NOT1_827 (N2810, N2776);
  not NOT1_844 (N2857, N2812);
  not NOT1_845 (N2858, N2815);
  not NOT1_846 (N2859, N2818);
  not NOT1_847 (N2860, N2821);
  not NOT1_848 (N2861, N2824);
  not NOT1_849 (N2862, N2829);
  not NOT1_857 (N2872, N2843);
  not NOT1_859 (N2874, N2846);
  not NOT1_877 (N2896, N2883);
  and g1 (N2384, N275, N2279, N306);
  and g2 (n_59, N2266, N2272);
  and g3 (N2558, N2361, N2104, N1171, n_59);
  and g5 (N2561, N2340, N2129, N1171, n_59);
  and g7 (N2564, N2340, N2119, N1171, n_59);
  and g9 (N2567, N2353, N2104, N1171, n_59);
  and g11 (N2570, N2375, N2119, N1188, n_59);
  and g13 (N2573, N2361, N2143, N1188, n_59);
  and g15 (N2576, N2375, N2129, N1188, n_59);
  and g16 (n_66, N2266, N2427);
  and g17 (N2639, N2361, N2129, N1171, n_66);
  and g19 (N2642, N2361, N2119, N1171, n_66);
  and g21 (N2645, N2375, N2104, N1171, n_66);
  and g23 (N2648, N2340, N2143, N1171, n_66);
  and g25 (N2651, N2353, N2129, N1188, n_66);
  and g26 (n_71, N2386, N2272);
  and g27 (N2655, N2361, N2129, N1188, n_71);
  and g29 (N2658, N2361, N2119, N1188, n_71);
  and g31 (N2661, N2375, N2104, N1188, n_71);
  and g33 (N2664, N2353, N2129, N1188, n_71);
  and g34 (n_75, N275, N2279, N99, N2747);
  and g35 (n_76, N2750, N2627, N2628);
  and g36 (n_77, N2629, N2630, N2631);
  and g37 (n_78, N2632, N2633, N2634);
  and g38 (N2800, n_75, n_76, n_77, n_78);
  and g39 (n_79, N2537, N2540);
  and g40 (n_80, N2543, N2546);
  and g41 (n_81, N2594, N2597);
  and g42 (n_82, N2600, N2603);
  and g43 (N2747, n_79, n_80, n_81, n_82);
  and g44 (n_83, N2606, N2549);
  and g45 (n_84, N2611, N2614);
  and g46 (n_85, N2617, N2620);
  and g47 (n_86, N2552, N2555);
  and g48 (N2750, n_83, n_84, n_85, n_86);
  and g49 (N2812, N49, N612, N94, N2789);
  and g50 (N2824, N56, N608, N94, N2789);
  not g51 (N923, N926);
endmodule

