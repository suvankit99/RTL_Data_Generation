
module ctrl(\opcode[0] , \opcode[1] , \opcode[2] , \opcode[3] ,
     \opcode[4] , \op_ext[0] , \op_ext[1] , \sel_reg_dst[0] ,
     \sel_reg_dst[1] , \sel_alu_opB[0] , \sel_alu_opB[1] , \alu_op[0] ,
     \alu_op[1] , \alu_op[2] , \alu_op_ext[0] , \alu_op_ext[1] ,
     \alu_op_ext[2] , \alu_op_ext[3] , halt, reg_write, sel_pc_opA,
     sel_pc_opB, beqz, bnez, bgez, bltz, jump, Cin, invA, invB, sign,
     mem_write, sel_wb);
  input \opcode[0] , \opcode[1] , \opcode[2] , \opcode[3] , \opcode[4]
       , \op_ext[0] , \op_ext[1] ;
  output \sel_reg_dst[0] , \sel_reg_dst[1] , \sel_alu_opB[0] ,
       \sel_alu_opB[1] , \alu_op[0] , \alu_op[1] , \alu_op[2] ,
       \alu_op_ext[0] , \alu_op_ext[1] , \alu_op_ext[2] ,
       \alu_op_ext[3] , halt, reg_write, sel_pc_opA, sel_pc_opB, beqz,
       bnez, bgez, bltz, jump, Cin, invA, invB, sign, mem_write, sel_wb;
  wire \opcode[0] , \opcode[1] , \opcode[2] , \opcode[3] , \opcode[4] ,
       \op_ext[0] , \op_ext[1] ;
  wire \sel_reg_dst[0] , \sel_reg_dst[1] , \sel_alu_opB[0] ,
       \sel_alu_opB[1] , \alu_op[0] , \alu_op[1] , \alu_op[2] ,
       \alu_op_ext[0] , \alu_op_ext[1] , \alu_op_ext[2] ,
       \alu_op_ext[3] , halt, reg_write, sel_pc_opA, sel_pc_opB, beqz,
       bnez, bgez, bltz, jump, Cin, invA, invB, sign, mem_write, sel_wb;
  wire n35, n36, n37, n38, n39, n40, n41, n42;
  wire n43, n44, n45, n46, n47, n48, n50, n51;
  wire n52, n53, n54, n55, n56, n57, n58, n59;
  wire n60, n61, n63, n64, n65, n66, n67, n68;
  wire n69, n71, n72, n73, n74, n75, n76, n77;
  wire n78, n80, n81, n82, n83, n84, n85, n86;
  wire n87, n88, n89, n90, n91, n92, n93, n94;
  wire n95, n96, n97, n99, n100, n101, n102, n103;
  wire n104, n106, n107, n108, n109, n110, n111, n112;
  wire n113, n114, n115, n117, n118, n119, n120, n121;
  wire n123, n124, n125, n126, n127, n128, n129, n131;
  wire n132, n134, n135, n136, n137, n139, n140, n141;
  wire n142, n143, n145, n146, n147, n148, n149, n150;
  wire n151, n153, n154, n156, n158, n159, n160, n161;
  wire n162, n164, n165, n166, n167, n169, n170, n171;
  wire n173, n174, n175, n177, n179, n180, n181, n182;
  wire n183, n184, n185, n186, n188, n189, n190, n191;
  wire n192, n193, n194, n195, n197, n198, n200, n201;
  wire n202, n203, n205, n206, n207, n_4, n_7, n_8;
  wire n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17;
  wire n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25;
  wire n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41;
  wire n_42, n_43, n_44, n_45, n_46, n_49, n_50, n_51;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140;
//   assign sign = 1'b1;
  not g1 (n_4, \opcode[1] );
  and g2 (n35, \opcode[0] , n_4);
  and g3 (n36, \opcode[3] , \opcode[4] );
  and g4 (n37, n35, n36);
  and g5 (n38, \opcode[1] , \opcode[3] );
  and g6 (n39, \opcode[4] , n38);
  not g7 (n_7, n37);
  not g8 (n_8, n39);
  and g9 (n40, n_7, n_8);
  not g10 (n_10, \opcode[2] );
  not g11 (n_11, n40);
  and g12 (n41, n_10, n_11);
  and g13 (n42, n_4, \opcode[3] );
  and g14 (n43, \opcode[4] , n42);
  not g15 (n_12, \opcode[3] );
  not g16 (n_13, \opcode[4] );
  and g17 (n44, n_12, n_13);
  not g18 (n_14, n36);
  not g19 (n_15, n44);
  and g20 (n45, n_14, n_15);
  not g21 (n_16, n45);
  and g22 (n46, \opcode[1] , n_16);
  not g23 (n_17, n43);
  not g24 (n_18, n46);
  and g25 (n47, n_17, n_18);
  not g26 (n_19, n47);
  and g27 (n48, \opcode[2] , n_19);
  or g28 (\sel_reg_dst[0] , n41, n48);
  not g29 (n_20, \opcode[0] );
  and g30 (n50, n_20, n_14);
  not g31 (n_21, n50);
  and g32 (n51, n_20, n_21);
  not g33 (n_22, n51);
  and g34 (n52, n_4, n_22);
  and g35 (n53, n_12, n_15);
  not g36 (n_23, n53);
  and g37 (n54, \opcode[1] , n_23);
  not g38 (n_24, n52);
  not g39 (n_25, n54);
  and g40 (n55, n_24, n_25);
  not g41 (n_26, n55);
  and g42 (n56, n_10, n_26);
  and g43 (n57, n_12, \opcode[4] );
  not g44 (n_27, n57);
  and g45 (n58, n_12, n_27);
  not g46 (n_28, n58);
  and g47 (n59, \opcode[1] , n_28);
  not g48 (n_29, n59);
  and g49 (n60, \opcode[1] , n_29);
  not g50 (n_30, n60);
  and g51 (n61, \opcode[2] , n_30);
  not g52 (n_31, n56);
  not g53 (n_32, n61);
  and g54 (\sel_reg_dst[1] , n_31, n_32);
  and g55 (n63, n_20, n_16);
  and g56 (n64, \opcode[3] , n_14);
  not g57 (n_33, n64);
  and g58 (n65, \opcode[0] , n_33);
  not g59 (n_34, n63);
  not g60 (n_35, n65);
  and g61 (n66, n_34, n_35);
  not g62 (n_36, n66);
  and g63 (n67, \opcode[1] , n_36);
  not g64 (n_37, n67);
  and g65 (n68, n_24, n_37);
  not g66 (n_38, n68);
  and g67 (n69, n_10, n_38);
  not g68 (n_39, n69);
  and g69 (\sel_alu_opB[0] , n_10, n_39);
  and g70 (n71, n_20, n_12);
  and g71 (n72, n_27, n71);
  and g72 (n73, \opcode[0] , n_16);
  not g73 (n_40, n72);
  not g74 (n_41, n73);
  and g75 (n74, n_40, n_41);
  not g76 (n_42, n74);
  and g77 (n75, n_4, n_42);
  not g78 (n_43, n75);
  and g79 (n76, n_25, n_43);
  not g80 (n_44, n76);
  and g81 (n77, n_10, n_44);
  and g82 (n78, \opcode[2] , n_23);
  not g83 (n_45, n77);
  not g84 (n_46, n78);
  and g85 (\sel_alu_opB[1] , n_45, n_46);
  and g86 (n80, n_20, \opcode[3] );
  and g87 (n81, \opcode[4] , \op_ext[0] );
  and g88 (n82, n80, n81);
  not g89 (n_49, \op_ext[1] );
  and g90 (n83, \opcode[3] , n_49);
  and g91 (n84, n_14, n83);
  not g92 (n_50, \op_ext[0] );
  and g93 (n85, \opcode[3] , n_50);
  and g94 (n86, n_14, n85);
  and g95 (n87, \opcode[3] , \op_ext[0] );
  not g96 (n_51, n86);
  not g97 (n_52, n87);
  and g98 (n88, n_51, n_52);
  not g99 (n_53, n88);
  and g100 (n89, \op_ext[1] , n_53);
  not g101 (n_54, n84);
  not g102 (n_55, n89);
  and g103 (n90, n_54, n_55);
  not g104 (n_56, n90);
  and g105 (n91, \opcode[0] , n_56);
  not g106 (n_57, n82);
  not g107 (n_58, n91);
  and g108 (n92, n_57, n_58);
  not g109 (n_59, n92);
  and g110 (n93, \opcode[1] , n_59);
  not g111 (n_60, n93);
  and g112 (n94, n_10, n_60);
  and g113 (n95, \opcode[0] , n_23);
  not g114 (n_61, n95);
  and g115 (n96, \opcode[0] , n_61);
  not g116 (n_62, n96);
  and g117 (n97, \opcode[2] , n_62);
  not g118 (n_63, n94);
  not g119 (n_64, n97);
  and g120 (\alu_op[0] , n_63, n_64);
  and g121 (n99, \opcode[3] , \op_ext[1] );
  not g122 (n_65, n99);
  and g123 (n100, n_54, n_65);
  not g124 (n_66, n100);
  and g125 (n101, \opcode[1] , n_66);
  not g126 (n_67, n101);
  and g127 (n102, n_10, n_67);
  and g128 (n103, \opcode[1] , n_25);
  not g129 (n_68, n103);
  and g130 (n104, \opcode[2] , n_68);
  not g131 (n_69, n102);
  not g132 (n_70, n104);
  and g133 (\alu_op[1] , n_69, n_70);
  and g134 (n106, n_4, n_14);
  and g135 (n107, n_15, n106);
  and g136 (n108, n_15, n50);
  and g137 (n109, \opcode[0] , n_28);
  not g138 (n_71, n108);
  not g139 (n_72, n109);
  and g140 (n110, n_71, n_72);
  not g141 (n_73, n110);
  and g142 (n111, \opcode[1] , n_73);
  not g143 (n_74, n107);
  not g144 (n_75, n111);
  and g145 (n112, n_74, n_75);
  not g146 (n_76, n112);
  and g147 (n113, n_10, n_76);
  and g148 (n114, \opcode[2] , \opcode[3] );
  and g149 (n115, \opcode[4] , n114);
  or g150 (\alu_op[2] , n113, n115);
  and g151 (n117, n_4, n_10);
  and g152 (n118, n_24, n117);
  and g153 (n119, \opcode[1] , n_42);
  not g154 (n_77, n119);
  and g155 (n120, n_7, n_77);
  not g156 (n_78, n120);
  and g157 (n121, \opcode[2] , n_78);
  or g158 (\alu_op_ext[0] , n118, n121);
  and g159 (n123, n_20, n_23);
  not g160 (n_79, n123);
  and g161 (n124, n_20, n_79);
  not g162 (n_80, n124);
  and g163 (n125, \opcode[1] , n_80);
  and g164 (n126, \opcode[1] , n_10);
  not g165 (n_81, n125);
  and g166 (n127, n_81, n126);
  and g167 (n128, \opcode[1] , \opcode[2] );
  and g168 (n129, n_16, n128);
  or g169 (\alu_op_ext[1] , n127, n129);
  not g170 (n_82, n106);
  and g171 (n131, n_82, n_81);
  not g172 (n_83, n131);
  and g173 (n132, n_10, n_83);
  not g174 (n_84, n132);
  and g175 (\alu_op_ext[2] , n_32, n_84);
  not g176 (n_85, n80);
  and g177 (n134, n_85, n_72);
  not g178 (n_86, n134);
  and g179 (n135, \opcode[1] , n_86);
  and g180 (n136, n_10, n_74);
  not g181 (n_87, n135);
  and g182 (n137, n_87, n136);
  not g183 (n_88, n137);
  and g184 (\alu_op_ext[3] , n_46, n_88);
  and g185 (n139, n_20, n_28);
  not g186 (n_89, n139);
  and g187 (n140, n_20, n_89);
  not g188 (n_90, n140);
  and g189 (n141, n_4, n_90);
  not g190 (n_91, n141);
  and g191 (n142, n_4, n_91);
  not g192 (n_92, n142);
  and g193 (n143, n_10, n_92);
  not g194 (n_93, n143);
  and g195 (halt, n_10, n_93);
  and g196 (n145, n_4, n_86);
  not g197 (n_94, n145);
  and g198 (n146, n_29, n_94);
  not g199 (n_95, n146);
  and g200 (n147, n_10, n_95);
  and g201 (n148, n_4, \opcode[4] );
  and g202 (n149, \opcode[1] , n_33);
  not g203 (n_96, n148);
  not g204 (n_97, n149);
  and g205 (n150, n_96, n_97);
  not g206 (n_98, n150);
  and g207 (n151, \opcode[2] , n_98);
  or g208 (reg_write, n147, n151);
  and g209 (n153, \opcode[0] , n_72);
  not g210 (n_99, n153);
  and g211 (n154, \opcode[2] , n_99);
  not g212 (n_100, n154);
  and g213 (sel_pc_opA, \opcode[2] , n_100);
  and g214 (n156, \opcode[2] , n_90);
  not g215 (n_101, n156);
  and g216 (sel_pc_opB, \opcode[2] , n_101);
  and g217 (n158, n_20, n_33);
  not g218 (n_102, n158);
  and g219 (n159, n_20, n_102);
  not g220 (n_103, n159);
  and g221 (n160, n_4, n_103);
  not g222 (n_104, n160);
  and g223 (n161, n_4, n_104);
  not g224 (n_105, n161);
  and g225 (n162, \opcode[2] , n_105);
  not g226 (n_106, n162);
  and g227 (beqz, \opcode[2] , n_106);
  and g228 (n164, \opcode[0] , n_35);
  not g229 (n_107, n164);
  and g230 (n165, n_4, n_107);
  not g231 (n_108, n165);
  and g232 (n166, n_4, n_108);
  not g233 (n_109, n166);
  and g234 (n167, \opcode[2] , n_109);
  not g235 (n_110, n167);
  and g236 (bnez, \opcode[2] , n_110);
  and g237 (n169, \opcode[1] , n_107);
  not g238 (n_111, n169);
  and g239 (n170, \opcode[1] , n_111);
  not g240 (n_112, n170);
  and g241 (n171, \opcode[2] , n_112);
  not g242 (n_113, n171);
  and g243 (bgez, \opcode[2] , n_113);
  and g244 (n173, \opcode[1] , n_103);
  not g245 (n_114, n173);
  and g246 (n174, \opcode[1] , n_114);
  not g247 (n_115, n174);
  and g248 (n175, \opcode[2] , n_115);
  not g249 (n_116, n175);
  and g250 (bltz, \opcode[2] , n_116);
  and g251 (n177, \opcode[2] , n_28);
  not g252 (n_117, n177);
  and g253 (jump, \opcode[2] , n_117);
  and g254 (n179, \opcode[0] , \opcode[1] );
  and g255 (n180, n_53, n179);
  and g256 (n181, n35, n_35);
  not g257 (n_118, n181);
  and g258 (n182, n_10, n_118);
  not g259 (n_119, n180);
  and g260 (n183, n_119, n182);
  and g261 (n184, \opcode[1] , n_22);
  not g262 (n_120, n184);
  and g263 (n185, n_82, n_120);
  not g264 (n_121, n185);
  and g265 (n186, \opcode[2] , n_121);
  not g266 (n_122, n183);
  not g267 (n_123, n186);
  and g268 (Cin, n_122, n_123);
  and g269 (n188, \op_ext[0] , n36);
  not g270 (n_124, n188);
  and g271 (n189, n_49, n_124);
  not g272 (n_125, n189);
  and g273 (n190, n_49, n_125);
  not g274 (n_126, n190);
  and g275 (n191, \opcode[0] , n_126);
  not g276 (n_127, n191);
  and g277 (n192, \opcode[0] , n_127);
  not g278 (n_128, n192);
  and g279 (n193, \opcode[1] , n_128);
  not g280 (n_129, n193);
  and g281 (n194, n_108, n_129);
  not g282 (n_130, n194);
  and g283 (n195, n_10, n_130);
  not g284 (n_131, n195);
  and g285 (invA, n_10, n_131);
  and g286 (n197, n_56, n179);
  not g287 (n_132, n197);
  and g288 (n198, n_10, n_132);
  not g289 (n_133, n198);
  and g290 (invB, n_123, n_133);
  and g291 (n200, n_4, n_80);
  and g292 (n201, \opcode[1] , n_62);
  not g293 (n_134, n200);
  not g294 (n_135, n201);
  and g295 (n202, n_134, n_135);
  not g296 (n_136, n202);
  and g297 (n203, n_10, n_136);
  not g298 (n_137, n203);
  and g299 (mem_write, n_10, n_137);
  and g300 (n205, n_4, n_62);
  not g301 (n_138, n205);
  and g302 (n206, n_4, n_138);
  not g303 (n_139, n206);
  and g304 (n207, n_10, n_139);
  not g305 (n_140, n207);
  and g306 (sel_wb, n_10, n_140);
endmodule

