
module i2c(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007,
     pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016,
     pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025,
     pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034,
     pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043,
     pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052,
     pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061,
     pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070,
     pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
     pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
     pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097,
     pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
     pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
     pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
     pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
     pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
     pi143, pi144, pi145, pi146, po000, po001, po002, po003, po004,
     po005, po006, po007, po008, po009, po010, po011, po012, po013,
     po014, po015, po016, po017, po018, po019, po020, po021, po022,
     po023, po024, po025, po026, po027, po028, po029, po030, po031,
     po032, po033, po034, po035, po036, po037, po038, po039, po040,
     po041, po042, po043, po044, po045, po046, po047, po048, po049,
     po050, po051, po052, po053, po054, po055, po056, po057, po058,
     po059, po060, po061, po062, po063, po064, po065, po066, po067,
     po068, po069, po070, po071, po072, po073, po074, po075, po076,
     po077, po078, po079, po080, po081, po082, po083, po084, po085,
     po086, po087, po088, po089, po090, po091, po092, po093, po094,
     po095, po096, po097, po098, po099, po100, po101, po102, po103,
     po104, po105, po106, po107, po108, po109, po110, po111, po112,
     po113, po114, po115, po116, po117, po118, po119, po120, po121,
     po122, po123, po124, po125, po126, po127, po128, po129, po130,
     po131, po132, po133, po134, po135, po136, po137, po138, po139,
     po140, po141);
  input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
       pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017,
       pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026,
       pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035,
       pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044,
       pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053,
       pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062,
       pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071,
       pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080,
       pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
       pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
       pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
       pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
       pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
       pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
       pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
       pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008,
       po009, po010, po011, po012, po013, po014, po015, po016, po017,
       po018, po019, po020, po021, po022, po023, po024, po025, po026,
       po027, po028, po029, po030, po031, po032, po033, po034, po035,
       po036, po037, po038, po039, po040, po041, po042, po043, po044,
       po045, po046, po047, po048, po049, po050, po051, po052, po053,
       po054, po055, po056, po057, po058, po059, po060, po061, po062,
       po063, po064, po065, po066, po067, po068, po069, po070, po071,
       po072, po073, po074, po075, po076, po077, po078, po079, po080,
       po081, po082, po083, po084, po085, po086, po087, po088, po089,
       po090, po091, po092, po093, po094, po095, po096, po097, po098,
       po099, po100, po101, po102, po103, po104, po105, po106, po107,
       po108, po109, po110, po111, po112, po113, po114, po115, po116,
       po117, po118, po119, po120, po121, po122, po123, po124, po125,
       po126, po127, po128, po129, po130, po131, po132, po133, po134,
       po135, po136, po137, po138, po139, po140, po141;
  wire pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
       pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017,
       pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026,
       pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035,
       pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044,
       pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053,
       pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062,
       pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071,
       pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080,
       pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
       pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
       pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
       pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
       pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
       pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
       pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
       pi144, pi145, pi146;
  wire po000, po001, po002, po003, po004, po005, po006, po007, po008,
       po009, po010, po011, po012, po013, po014, po015, po016, po017,
       po018, po019, po020, po021, po022, po023, po024, po025, po026,
       po027, po028, po029, po030, po031, po032, po033, po034, po035,
       po036, po037, po038, po039, po040, po041, po042, po043, po044,
       po045, po046, po047, po048, po049, po050, po051, po052, po053,
       po054, po055, po056, po057, po058, po059, po060, po061, po062,
       po063, po064, po065, po066, po067, po068, po069, po070, po071,
       po072, po073, po074, po075, po076, po077, po078, po079, po080,
       po081, po082, po083, po084, po085, po086, po087, po088, po089,
       po090, po091, po092, po093, po094, po095, po096, po097, po098,
       po099, po100, po101, po102, po103, po104, po105, po106, po107,
       po108, po109, po110, po111, po112, po113, po114, po115, po116,
       po117, po118, po119, po120, po121, po122, po123, po124, po125,
       po126, po127, po128, po129, po130, po131, po132, po133, po134,
       po135, po136, po137, po138, po139, po140, po141;
  wire n291, n294, n295, n298, n299, n300, n301, n302;
  wire n305, n306, n307, n308, n309, n310, n311, n312;
  wire n313, n314, n315, n317, n319, n320, n321, n322;
  wire n323, n324, n325, n326, n327, n328, n332, n333;
  wire n334, n335, n336, n337, n338, n339, n341, n344;
  wire n345, n346, n347, n350, n351, n352, n353, n354;
  wire n355, n356, n357, n358, n360, n362, n363, n364;
  wire n365, n366, n367, n368, n369, n370, n371, n375;
  wire n376, n377, n379, n380, n381, n383, n384, n385;
  wire n387, n388, n389, n390, n391, n394, n395, n396;
  wire n397, n398, n399, n401, n403, n404, n405, n406;
  wire n407, n408, n409, n410, n411, n412, n413, n414;
  wire n416, n417, n418, n419, n423, n424, n425, n426;
  wire n427, n428, n433, n434, n435, n436, n437, n438;
  wire n440, n445, n447, n448, n449, n450, n454, n455;
  wire n456, n458, n459, n468, n469, n470, n472, n473;
  wire n479, n482, n483, n484, n486, n487, n488, n494;
  wire n495, n496, n498, n503, n507, n508, n509, n511;
  wire n515, n519, n520, n521, n523, n530, n531, n532;
  wire n534, n540, n541, n542, n544, n548, n549, n553;
  wire n554, n555, n557, n564, n565, n566, n568, n570;
  wire n572, n573, n575, n576, n577, n578, n579, n580;
  wire n581, n582, n583, n584, n588, n589, n590, n591;
  wire n592, n593, n595, n600, n601, n602, n604, n612;
  wire n616, n617, n618, n620, n624, n625, n626, n628;
  wire n634, n635, n636, n638, n639, n640, n641, n642;
  wire n645, n646, n647, n648, n649, n650, n653, n654;
  wire n655, n656, n657, n658, n659, n660, n662, n668;
  wire n669, n670, n672, n681, n682, n683, n685, n686;
  wire n688, n689, n690, n691, n692, n693, n694, n695;
  wire n696, n697, n698, n699, n700, n701, n702, n703;
  wire n704, n705, n709, n713, n714, n715, n716, n717;
  wire n718, n719, n720, n721, n722, n723, n724, n725;
  wire n726, n727, n728, n729, n730, n731, n732, n733;
  wire n734, n735, n736, n737, n738, n739, n740, n741;
  wire n742, n743, n744, n745, n746, n747, n748, n749;
  wire n750, n751, n752, n753, n754, n755, n756, n757;
  wire n758, n759, n761, n762, n763, n764, n765, n766;
  wire n767, n768, n769, n770, n773, n774, n776, n777;
  wire n778, n779, n780, n781, n782, n783, n784, n787;
  wire n788, n790, n791, n792, n793, n794, n795, n796;
  wire n797, n798, n799, n802, n803, n804, n805, n806;
  wire n807, n808, n809, n810, n811, n812, n813, n814;
  wire n815, n816, n817, n818, n819, n820, n821, n822;
  wire n823, n824, n825, n826, n827, n829, n830, n831;
  wire n832, n833, n834, n835, n836, n837, n838, n839;
  wire n840, n841, n842, n843, n844, n845, n846, n847;
  wire n848, n849, n850, n851, n852, n853, n854, n855;
  wire n856, n857, n858, n859, n861, n862, n863, n864;
  wire n865, n866, n868, n869, n870, n871, n872, n873;
  wire n875, n876, n877, n878, n879, n880, n882, n883;
  wire n884, n885, n886, n887, n889, n890, n891, n892;
  wire n893, n894, n896, n897, n898, n899, n900, n901;
  wire n903, n904, n905, n906, n907, n908, n910, n911;
  wire n912, n913, n914, n915, n917, n918, n919, n920;
  wire n921, n922, n923, n924, n927, n930, n931, n932;
  wire n933, n934, n935, n936, n940, n941, n942, n943;
  wire n944, n945, n947, n948, n949, n950, n951, n952;
  wire n953, n956, n957, n958, n959, n960, n961, n965;
  wire n966, n967, n968, n969, n972, n973, n974, n975;
  wire n976, n979, n983, n984, n985, n986, n987, n988;
  wire n989, n990, n991, n992, n993, n994, n995, n996;
  wire n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007;
  wire n1008, n1009, n1010, n1013, n1017, n1018, n1019, n1020;
  wire n1021, n1022, n1023, n1024, n1026, n1027, n1028, n1029;
  wire n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  wire n1038, n1039, n1040, n1041, n1044, n1048, n1049, n1050;
  wire n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058;
  wire n1059, n1060, n1064, n1065, n1066, n1067, n1068, n1069;
  wire n1070, n1071, n1072, n1076, n1080, n1081, n1082, n1083;
  wire n1084, n1085, n1087, n1089, n1090, n1091, n1092, n1096;
  wire n1100, n1101, n1102, n1103, n1104, n1107, n1108, n1109;
  wire n1112, n1113, n1114, n1115, n1116, n1117, n1119, n1120;
  wire n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128;
  wire n1129, n1130, n1131, n1132, n1136, n1137, n1138, n1140;
  wire n1141, n1142, n1144, n1147, n1148, n1149, n1150, n1151;
  wire n1152, n1157, n1158, n1159, n1162, n1164, n1165, n1166;
  wire n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174;
  wire n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182;
  wire n1183, n1184, n1185, n1187, n1188, n1189, n1190, n1191;
  wire n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199;
  wire n1200, n1201, n1202, n1203, n1205, n1208, n1209, n1214;
  wire n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;
  wire n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230;
  wire n1231, n1232, n1233, n1234, n1236, n1237, n1238, n1245;
  wire n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253;
  wire n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263;
  wire n1265, n1266, n1267, n1268, n1270, n1271, n1272, n1273;
  wire n1274, n1276, n1277, n1278, n1280, n1281, n1282, n1283;
  wire n1285, n1286, n1287, n1288, n1290, n1291, n1292, n1293;
  wire n1295, n1296, n1297, n1298, n1300, n1301, n1302, n1304;
  wire n1305, n1306, n1308, n1309, n1310, n1312, n1313, n1314;
  wire n1316, n1317, n1318, n1320, n1321, n1322, n1324, n1325;
  wire n1326, n1327, n1328, n1330, n1331, n1332, n1334, n1335;
  wire n1336, n1338, n1339, n1340, n1342, n1343, n1344, n1346;
  wire n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354;
  wire n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362;
  wire n1363, n1365, n1366, n1367, n1369, n1370, n1371, n1372;
  wire n1377, n1378, n1379, n1381, n1382, n1383, n1385, n1386;
  wire n1387, n1388, n1389, n1391, n1392, n1393, n1395, n1396;
  wire n1397, n1399, n1400, n1401, n1403, n1404, n1405, n1407;
  wire n1408, n1409, n1411, n1412, n1413, n1414, n1415, n1416;
  wire n1417, n1419, n1420, n1421, n1422, n1423, n1424, n1425;
  wire n1426, n1428, n1429, n1430, n1432, n1433, n1434, n1436;
  wire n1437, n1438, n1440, n1441, n1442, n1444, n1445, n1446;
  wire n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455;
  wire n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463;
  wire n1464, n1466, n1467, n1468, n1469, n1470, n1471, n1472;
  wire n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1481;
  wire n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489;
  wire n1490, n1491, n1492, n1493, n1494, n1496, n1497, n1498;
  wire n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506;
  wire n1507, n1508, n1509, n1511, n1512, n1513, n1514, n1515;
  wire n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523;
  wire n1524, n1525, n1526, n1527, n1529, n1530, n1531, n1532;
  wire n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541;
  wire n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549;
  wire n1550, n1552, n1553, n1554, n1555, n1556, n1557, n1558;
  wire n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566;
  wire n1567, n1568, n1570, n1571, n1575, n1576, n1580, n1581;
  wire n1582, n1583, n1584, n1585, n1586, n1588, n1589, n1590;
  wire n1591, n1592, n1594, n1595, n1596, n1597, n1598, n1600;
  wire n1601, n1602, n1603, n1604, n1608, n1613, n1614, n1615;
  wire n1616, n1619, n1620, n1621, n1623, n1628, n1629, n1631;
  wire n_4, n_5, n_8, n_9, n_12, n_13, n_15, n_17;
  wire n_20, n_21, n_24, n_25, n_28, n_29, n_32, n_33;
  wire n_35, n_37, n_38, n_39, n_41, n_42, n_43, n_47;
  wire n_48, n_49, n_50, n_51, n_53, n_54, n_55, n_56;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_67, n_68, n_70, n_71, n_73, n_74, n_75, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_88;
  wire n_89, n_90, n_91, n_96, n_97, n_100, n_101, n_104;
  wire n_105, n_108, n_109, n_112, n_113, n_116, n_117, n_120;
  wire n_121, n_123, n_125, n_127, n_128, n_129, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_142;
  wire n_143, n_144, n_146, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_159, n_160, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_198, n_199, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_239, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_257, n_258, n_260, n_261, n_262, n_264, n_265, n_266;
  wire n_267, n_269, n_270, n_273, n_274, n_276, n_278, n_279;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_305, n_306;
  wire n_307, n_308, n_310, n_311, n_312, n_313, n_314, n_315;
  wire n_316, n_317, n_318, n_319, n_320, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_383;
  wire n_385, n_386, n_388, n_389, n_391, n_392, n_393, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_420, n_421, n_422, n_423, n_424, n_425, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_472, n_473, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_490, n_491, n_492;
  wire n_493, n_494, n_495, n_496, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_513, n_515, n_516, n_517;
  wire n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_568, n_569, n_571, n_572, n_574, n_575;
  wire n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_587, n_588, n_593, n_594, n_595;
  wire n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_604;
  wire n_605, n_607, n_609, n_610, n_611, n_613, n_614, n_615;
  wire n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623;
  wire n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631;
  wire n_632, n_633, n_634, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_665, n_666;
  wire n_670, n_671, n_676, n_678, n_679, n_680, n_682, n_683;
  wire n_684, n_686, n_687, n_688, n_690, n_691, n_692, n_693;
  wire n_694, n_696, n_697, n_698, n_699, n_700, n_702, n_703;
  wire n_704, n_705, n_706, n_708, n_709, n_710, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_728, n_729, n_730;
  wire n_731, n_733, n_734, n_735, n_737, n_738, n_739, n_741;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
  wire n_760, n_762, n_763, n_764, n_765, n_766, n_767, n_769;
  wire n_770, n_771, n_772, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787;
  wire n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811;
  wire n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819;
  wire n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_872, n_873, n_874, n_875, n_876, n_877;
  wire n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885;
  wire n_886, n_887, n_888, n_889, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902;
  wire n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_927;
  wire n_928, n_929, n_930, n_931, n_932, n_933, n_935, n_936;
  wire n_937, n_938, n_939, n_940, n_941, n_942, n_944, n_946;
  wire n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954;
  wire n_955, n_956, n_957, n_958, n_960, n_961, n_962, n_963;
  wire n_964, n_965, n_966, n_969, n_970, n_972, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1150, n_1151, n_1152, n_1154;
  wire n_1156, n_1157, n_1158, n_1159, n_1161, n_1162, n_1163, n_1164;
  wire n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172;
  wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1181;
  wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189;
  wire n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197;
  wire n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213;
  wire n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
//   assign po014 = pi128;
  assign po013 = pi130;
//   assign po012 = 1'b1;
  assign po011 = pi000;
  assign po010 = pi001;
  assign po009 = pi121;
  assign po008 = pi126;
  assign po007 = pi101;
  assign po006 = pi107;
  assign po005 = pi105;
  assign po004 = pi102;
//   assign po003 = pi103;
//   assign po002 = pi104;
  assign po001 = pi083;
//   assign po000 = pi108;
  not g1 (n_4, pi013);
  not g2 (n_5, pi014);
  and g3 (n291, n_4, n_5);
  not g4 (n_8, pi006);
  not g5 (n_9, pi007);
  not g8 (n_12, pi017);
  not g9 (n_13, pi021);
  and g10 (n294, n_12, n_13);
  not g11 (n_15, pi008);
  and g12 (n295, n_15, n294);
  not g13 (n_17, pi012);
  not g16 (n_20, pi018);
  not g17 (n_21, pi019);
  and g18 (n298, n_20, n_21);
  not g19 (n_24, pi004);
  not g20 (n_25, pi016);
  and g21 (n299, n_24, n_25);
  and g22 (n300, n298, n299);
  not g23 (n_28, pi005);
  not g24 (n_29, pi022);
  and g25 (n301, n_28, n_29);
  not g26 (n_32, pi009);
  not g27 (n_33, pi011);
  and g28 (n302, n_32, n_33);
  not g32 (n_35, n305);
  and g33 (n306, pi054, n_35);
  not g34 (n_37, pi000);
  not g35 (n_38, n306);
  and g36 (n307, n_37, n_38);
  not g37 (n_39, n302);
  and g38 (n308, n301, n_39);
  not g39 (n_41, pi056);
  and g40 (n309, n_41, n308);
  not g41 (n_42, n301);
  and g42 (n310, n_41, n_42);
  and g43 (n311, n_15, n_13);
  and g44 (n312, n_9, pi013);
  and g45 (n313, n311, n312);
  and g46 (n314, n_9, n311);
  not g47 (n_43, n311);
  and g48 (n315, pi007, n_43);
  and g52 (n317, pi008, pi021);
  not g56 (n_47, n313);
  not g57 (n_48, n319);
  and g58 (n320, n_47, n_48);
  not g59 (n_49, n320);
  and g60 (n321, n_5, n_49);
  and g61 (n322, n_4, pi014);
  and g62 (n323, n314, n322);
  not g63 (n_50, n321);
  not g64 (n_51, n323);
  and g65 (n324, n_50, n_51);
  not g66 (n_53, pi010);
  not g67 (n_54, n324);
  and g68 (n325, n_53, n_54);
  and g69 (n326, pi010, n291);
  and g70 (n327, n314, n326);
  not g71 (n_55, n325);
  not g72 (n_56, n327);
  and g73 (n328, n_55, n_56);
  and g78 (n332, n_8, n_17);
  not g80 (n_58, n310);
  not g81 (n_59, n333);
  and g82 (n334, n_58, n_59);
  not g83 (n_60, n334);
  and g84 (n335, n302, n_60);
  not g85 (n_61, n309);
  not g86 (n_62, n335);
  and g87 (n336, n_61, n_62);
  not g88 (n_63, n336);
  and g89 (n337, pi054, n_63);
  not g90 (n_64, n307);
  not g91 (n_65, n337);
  and g92 (n338, n_64, n_65);
  not g93 (n_67, pi129);
  not g94 (n_68, n338);
  and g95 (n339, n_67, n_68);
  not g96 (n_70, n339);
  or g97 (po015, pi003, n_70);
  and g98 (n341, n_33, n_17);
  and g101 (n344, n_53, n_29);
  and g102 (n345, n_9, n_4);
  and g103 (n346, n_28, n_8);
  and g104 (n347, n345, n346);
  and g108 (n351, n_12, pi054);
  not g109 (n_71, n350);
  and g110 (n352, n_71, n351);
  not g111 (n_73, pi001);
  not g112 (n_74, n352);
  and g113 (n353, n_73, n_74);
  and g114 (n354, n_5, pi054);
  and g115 (n355, n_15, n_33);
  and g116 (n356, n294, n355);
  and g117 (n357, n_28, n332);
  not g118 (n_75, n332);
  and g119 (n358, pi005, n_75);
  and g123 (n360, pi006, pi012);
  and g127 (n363, pi007, n357);
  not g128 (n_79, n362);
  not g129 (n_80, n363);
  and g130 (n364, n_79, n_80);
  not g131 (n_81, n364);
  and g132 (n365, n_4, n_81);
  and g133 (n366, n312, n357);
  not g134 (n_82, n365);
  not g135 (n_83, n366);
  and g136 (n367, n_82, n_83);
  not g137 (n_84, n367);
  and g138 (n368, n_32, n_84);
  and g139 (n369, n345, n357);
  and g140 (n370, pi009, n369);
  not g141 (n_85, n368);
  not g142 (n_86, n370);
  and g143 (n371, n_85, n_86);
  not g149 (n_88, n353);
  not g150 (n_89, n375);
  and g151 (n376, n_88, n_89);
  not g152 (n_90, n376);
  and g153 (n377, n_67, n_90);
  not g154 (n_91, n377);
  or g155 (po016, pi003, n_91);
  and g156 (n379, pi122, pi127);
  not g157 (n_96, pi045);
  not g158 (n_97, pi048);
  and g159 (n380, n_96, n_97);
  not g160 (n_100, pi043);
  not g161 (n_101, pi047);
  and g162 (n381, n_100, n_101);
  not g164 (n_104, pi015);
  not g165 (n_105, pi020);
  and g166 (n383, n_104, n_105);
  not g167 (n_108, pi024);
  not g168 (n_109, pi049);
  and g169 (n384, n_108, n_109);
  and g170 (n385, n383, n384);
  not g172 (n_112, pi041);
  not g173 (n_113, pi046);
  and g174 (n387, n_112, n_113);
  not g175 (n_116, pi038);
  not g176 (n_117, pi050);
  and g177 (n388, n_116, n_117);
  and g178 (n389, n387, n388);
  not g179 (n_120, pi042);
  not g180 (n_121, pi044);
  and g181 (n390, n_120, n_121);
  not g182 (n_123, pi040);
  and g183 (n391, n_123, n390);
  not g184 (n_125, pi002);
  not g188 (n_127, n394);
  and g189 (n395, pi082, n_127);
  not g190 (n_128, n379);
  not g191 (n_129, n395);
  and g192 (n396, n_128, n_129);
  not g193 (n_131, pi065);
  and g194 (n397, n_131, n396);
  and g195 (n398, n_108, n_96);
  and g196 (n399, n_101, n_97);
  and g198 (n401, n_109, n383);
  and g200 (n403, n_116, n_123);
  and g201 (n404, n390, n403);
  and g202 (n405, n_113, n_117);
  and g203 (n406, n_112, n405);
  and g204 (n407, n404, n406);
  and g205 (n408, n_100, n407);
  not g207 (n_132, n409);
  and g208 (n410, pi082, n_132);
  not g209 (n_133, pi082);
  and g210 (n411, n_133, n379);
  not g211 (n_134, n410);
  not g212 (n_135, n411);
  and g213 (n412, n_134, n_135);
  not g214 (n_136, n412);
  and g215 (n413, pi002, n_136);
  not g216 (n_137, n397);
  not g217 (n_138, n413);
  and g218 (n414, n_137, n_138);
  not g219 (n_139, n414);
  and g220 (po017, n_67, n_139);
  and g221 (n416, n_32, n_5);
  and g222 (n417, n344, n416);
  and g223 (n418, n347, n417);
  and g224 (n419, n_15, n_12);
  not g229 (n_142, pi061);
  not g230 (n_143, pi118);
  and g231 (n424, n_142, n_143);
  not g232 (n_144, n423);
  and g233 (n425, n_144, n424);
  not g234 (n_146, pi123);
  and g235 (n426, pi000, n_146);
  not g236 (n_148, pi113);
  and g237 (n427, n_148, n426);
  not g238 (n_149, n425);
  not g239 (n_150, n427);
  and g240 (n428, n_149, n_150);
  not g241 (n_151, n428);
  and g242 (po018, n_67, n_151);
  and g246 (n433, pi054, n300);
  and g247 (n434, n356, n433);
  not g249 (n_152, pi054);
  and g250 (n436, pi004, n_152);
  not g251 (n_153, n435);
  not g252 (n_154, n436);
  and g253 (n437, n_153, n_154);
  not g254 (n_155, n437);
  and g255 (n438, n_67, n_155);
  not g256 (n_156, pi003);
  and g257 (po019, n_156, n438);
  and g258 (n440, pi005, n_152);
  not g260 (n_159, pi025);
  not g261 (n_160, pi029);
  and g265 (n445, n_4, n417);
  not g267 (n_163, pi059);
  and g268 (n447, n_163, n356);
  and g269 (n448, n_25, pi054);
  and g270 (n449, n_24, n_21);
  and g271 (n450, n_20, n449);
  not g276 (n_164, n440);
  not g277 (n_165, n454);
  and g278 (n455, n_164, n_165);
  not g279 (n_166, n455);
  and g280 (n456, n_67, n_166);
  and g281 (po020, n_156, n456);
  and g282 (n458, pi006, n_152);
  and g283 (n459, n_28, n_9);
  not g285 (n_167, pi028);
  not g294 (n_168, n458);
  not g295 (n_169, n468);
  and g296 (n469, n_168, n_169);
  not g297 (n_170, n469);
  and g298 (n470, n_67, n_170);
  and g299 (po021, n_156, n470);
  and g300 (n472, pi007, n_152);
  and g301 (n473, n_20, n_13);
  and g307 (n479, n_8, n341);
  not g311 (n_171, n472);
  not g312 (n_172, n482);
  and g313 (n483, n_171, n_172);
  not g314 (n_173, n483);
  and g315 (n484, n_67, n_173);
  and g316 (po022, n_156, n484);
  and g317 (n486, pi008, n_152);
  and g318 (n487, n369, n417);
  and g319 (n488, n_12, n_20);
  not g326 (n_174, n486);
  not g327 (n_175, n494);
  and g328 (n495, n_174, n_175);
  not g329 (n_176, n495);
  and g330 (n496, n_67, n_176);
  and g331 (po023, n_156, n496);
  and g332 (n498, pi009, n_152);
  and g337 (n503, n419, n473);
  not g342 (n_177, n498);
  not g343 (n_178, n507);
  and g344 (n508, n_177, n_178);
  not g345 (n_179, n508);
  and g346 (n509, n_67, n_179);
  and g347 (po024, n_156, n509);
  and g348 (n511, pi010, n_152);
  and g352 (n515, n459, n479);
  not g357 (n_180, n511);
  not g358 (n_181, n519);
  and g359 (n520, n_180, n_181);
  not g360 (n_182, n520);
  and g361 (n521, n_67, n_182);
  and g362 (po025, n_156, n521);
  and g363 (n523, pi011, n_152);
  not g371 (n_183, n523);
  not g372 (n_184, n530);
  and g373 (n531, n_183, n_184);
  not g374 (n_185, n531);
  and g375 (n532, n_67, n_185);
  and g376 (po026, n_156, n532);
  and g377 (n534, pi012, n_152);
  not g384 (n_186, n534);
  not g385 (n_187, n540);
  and g386 (n541, n_186, n_187);
  not g387 (n_188, n541);
  and g388 (n542, n_67, n_188);
  and g389 (po027, n_156, n542);
  and g390 (n544, pi013, n_152);
  and g394 (n548, n_159, pi029);
  and g395 (n549, n_167, n548);
  not g400 (n_189, n544);
  not g401 (n_190, n553);
  and g402 (n554, n_189, n_190);
  not g403 (n_191, n554);
  and g404 (n555, n_67, n_191);
  and g405 (po028, n_156, n555);
  and g406 (n557, pi014, n_152);
  not g414 (n_192, n557);
  not g415 (n_193, n564);
  and g416 (n565, n_192, n_193);
  not g417 (n_194, n565);
  and g418 (n566, n_67, n_194);
  and g419 (po029, n_156, n566);
  and g420 (n568, n_112, n_100);
  and g422 (n570, n_96, n384);
  and g424 (n572, n_113, n388);
  and g425 (n573, n391, n572);
  not g428 (n_195, n575);
  and g429 (n576, pi082, n_195);
  not g430 (n_196, n576);
  and g431 (n577, n_128, n_196);
  not g432 (n_198, pi070);
  and g433 (n578, n_198, n577);
  and g434 (n579, n_97, n381);
  and g435 (n580, n570, n579);
  and g436 (n581, n407, n580);
  not g437 (n_199, n581);
  and g438 (n582, pi015, n_199);
  and g439 (n583, n_96, n399);
  and g440 (n584, n_125, n_105);
  not g446 (n_201, n582);
  not g447 (n_202, n588);
  and g448 (n589, n_201, n_202);
  not g449 (n_203, n589);
  and g450 (n590, pi082, n_203);
  and g451 (n591, pi015, n411);
  not g452 (n_204, n590);
  not g453 (n_205, n591);
  and g454 (n592, n_204, n_205);
  not g455 (n_206, n578);
  and g456 (n593, n_206, n592);
  not g457 (n_207, n593);
  and g458 (po030, n_67, n_207);
  and g459 (n595, pi016, n_152);
  not g465 (n_208, n595);
  not g466 (n_209, n600);
  and g467 (n601, n_208, n_209);
  not g468 (n_210, n601);
  and g469 (n602, n_67, n_210);
  and g470 (po031, n_156, n602);
  and g471 (n604, pi017, n_152);
  and g479 (n612, n_33, n311);
  not g484 (n_211, n604);
  not g485 (n_212, n616);
  and g486 (n617, n_211, n_212);
  not g487 (n_213, n617);
  and g488 (n618, n_67, n_213);
  and g489 (po032, n_156, n618);
  and g490 (n620, pi018, n_152);
  not g495 (n_214, n620);
  not g496 (n_215, n624);
  and g497 (n625, n_214, n_215);
  not g498 (n_216, n625);
  and g499 (n626, n_67, n_216);
  and g500 (po033, n_156, n626);
  and g501 (n628, pi019, n_152);
  not g508 (n_217, n628);
  not g509 (n_218, n634);
  and g510 (n635, n_217, n_218);
  not g511 (n_219, n635);
  and g512 (n636, n_67, n_219);
  and g513 (po034, n_156, n636);
  and g514 (n638, n381, n387);
  and g515 (n639, n_108, n380);
  and g516 (n640, n638, n639);
  and g517 (n641, n_123, n_120);
  and g518 (n642, n388, n641);
  not g522 (n_220, n645);
  and g523 (n646, pi082, n_220);
  not g524 (n_221, n646);
  and g525 (n647, n_128, n_221);
  not g526 (n_223, pi071);
  and g527 (n648, n_223, n647);
  and g528 (n649, n_117, n403);
  and g529 (n650, n_104, n_109);
  not g533 (n_224, n653);
  and g534 (n654, pi020, n_224);
  and g535 (n655, pi002, n645);
  not g536 (n_225, n654);
  not g537 (n_226, n655);
  and g538 (n656, n_225, n_226);
  not g539 (n_227, n656);
  and g540 (n657, pi082, n_227);
  and g541 (n658, pi020, n411);
  not g542 (n_228, n657);
  not g543 (n_229, n658);
  and g544 (n659, n_228, n_229);
  not g545 (n_230, n648);
  and g546 (n660, n_230, n659);
  not g547 (n_231, n660);
  and g548 (po035, n_67, n_231);
  and g549 (n662, pi021, n_152);
  not g556 (n_232, n662);
  not g557 (n_233, n668);
  and g558 (n669, n_232, n_233);
  not g559 (n_234, n669);
  and g560 (n670, n_67, n_234);
  and g561 (po036, n_156, n670);
  and g562 (n672, pi022, n_152);
  not g572 (n_235, n672);
  not g573 (n_236, n681);
  and g574 (n682, n_235, n_236);
  not g575 (n_237, n682);
  and g576 (n683, n_67, n_237);
  and g577 (po037, n_156, n683);
  not g578 (n_239, pi023);
  and g579 (n685, n_239, pi055);
  not g580 (n_241, n685);
  and g581 (n686, n_67, n_241);
  and g582 (po038, pi061, n686);
  and g583 (n688, n_101, n568);
  and g584 (n689, n380, n688);
  and g585 (n690, n573, n689);
  not g586 (n_242, n690);
  and g587 (n691, pi082, n_242);
  and g588 (n692, n584, n650);
  not g589 (n_243, n692);
  and g590 (n693, pi082, n_243);
  not g591 (n_244, n693);
  and g592 (n694, n379, n_244);
  not g593 (n_245, n691);
  not g594 (n_246, n694);
  and g595 (n695, n_245, n_246);
  not g596 (n_247, n695);
  and g597 (n696, n_108, n_247);
  and g598 (n697, n_125, n_96);
  and g599 (n698, n399, n697);
  and g600 (n699, n401, n698);
  and g601 (n700, n408, n699);
  not g602 (n_248, n700);
  and g603 (n701, pi082, n_248);
  not g604 (n_249, n701);
  and g605 (n702, n_128, n_249);
  and g606 (n703, pi063, n702);
  and g607 (n704, n_100, n387);
  and g608 (n705, n583, n704);
  and g619 (n713, pi085, pi116);
  not g620 (n_257, pi085);
  not g621 (n_258, pi110);
  and g622 (n714, n_257, n_258);
  not g623 (n_260, pi096);
  and g624 (n715, n_260, n714);
  not g625 (n_261, n713);
  not g626 (n_262, n715);
  and g627 (n716, n_261, n_262);
  not g628 (n_264, n716);
  and g629 (n717, pi100, n_264);
  not g630 (n_265, pi116);
  and g631 (n718, pi025, n_265);
  and g632 (n719, pi085, n718);
  not g633 (n_266, n717);
  not g634 (n_267, n719);
  and g635 (n720, n_266, n_267);
  not g636 (n_269, pi026);
  not g637 (n_270, n720);
  and g638 (n721, n_269, n_270);
  not g639 (n_273, pi051);
  not g640 (n_274, pi052);
  and g641 (n722, n_273, n_274);
  not g642 (n_276, pi039);
  and g643 (n723, n_276, n722);
  not g644 (n_278, pi095);
  not g645 (n_279, pi100);
  and g646 (n724, n_278, n_279);
  not g647 (n_281, pi097);
  and g648 (n725, n_281, n724);
  not g649 (n_282, n725);
  and g650 (n726, n_258, n_282);
  not g651 (n_283, n726);
  and g652 (n727, pi025, n_283);
  and g653 (n728, pi026, pi116);
  not g654 (n_284, n727);
  not g655 (n_285, n728);
  and g656 (n729, n_284, n_285);
  not g657 (n_286, n723);
  not g658 (n_287, n729);
  and g659 (n730, n_286, n_287);
  and g660 (n731, pi026, n718);
  not g661 (n_288, n730);
  not g662 (n_289, n731);
  and g663 (n732, n_288, n_289);
  not g664 (n_290, n732);
  and g665 (n733, n_257, n_290);
  not g666 (n_291, n721);
  not g667 (n_292, n733);
  and g668 (n734, n_291, n_292);
  not g669 (n_294, pi027);
  not g670 (n_295, n734);
  and g671 (n735, n_294, n_295);
  and g672 (n736, n_276, n_274);
  and g673 (n737, n_273, n736);
  and g674 (n738, pi116, n737);
  not g675 (n_296, n718);
  not g676 (n_297, n738);
  and g677 (n739, n_296, n_297);
  not g678 (n_298, n739);
  and g679 (n740, pi027, n_298);
  and g680 (n741, n723, n727);
  not g681 (n_299, n740);
  not g682 (n_300, n741);
  and g683 (n742, n_299, n_300);
  and g684 (n743, n_269, n_257);
  not g685 (n_301, n742);
  and g686 (n744, n_301, n743);
  not g687 (n_302, n735);
  not g688 (n_303, n744);
  and g689 (n745, n_302, n_303);
  not g690 (n_305, pi053);
  not g691 (n_306, n745);
  and g692 (n746, n_305, n_306);
  and g693 (n747, pi025, n_269);
  and g694 (n748, n_265, n747);
  and g695 (n749, pi053, n_257);
  and g696 (n750, n_294, n749);
  and g697 (n751, n748, n750);
  not g698 (n_307, n746);
  not g699 (n_308, n751);
  and g700 (n752, n_307, n_308);
  not g701 (n_310, pi058);
  not g702 (n_311, n752);
  and g703 (n753, n_310, n_311);
  and g704 (n754, n_294, n_257);
  and g705 (n755, n_305, pi058);
  and g706 (n756, n754, n755);
  and g707 (n757, n748, n756);
  not g708 (n_312, n753);
  not g709 (n_313, n757);
  and g710 (n758, n_312, n_313);
  not g711 (n_314, n758);
  and g712 (n759, n_67, n_314);
  and g713 (po040, n_156, n759);
  and g714 (n761, pi085, n_265);
  not g715 (n_315, n761);
  and g716 (n762, n_258, n_315);
  and g717 (n763, n_285, n762);
  and g718 (n764, n_260, n763);
  and g719 (n765, n_269, n713);
  not g720 (n_316, n764);
  not g721 (n_317, n765);
  and g722 (n766, n_316, n_317);
  not g723 (n_318, n766);
  and g724 (n767, pi100, n_318);
  and g725 (n768, n_257, n_297);
  and g726 (n769, pi026, n768);
  not g727 (n_319, n767);
  not g728 (n_320, n769);
  and g729 (n770, n_319, n_320);
  and g733 (n773, n_294, n_305);
  and g734 (n774, n_310, n773);
  and g736 (n776, pi095, n_260);
  and g737 (n777, pi027, pi116);
  not g738 (n_322, n777);
  and g739 (n778, n762, n_322);
  and g740 (n779, n776, n778);
  and g741 (n780, n_294, n713);
  not g742 (n_323, n779);
  not g743 (n_324, n780);
  and g744 (n781, n_323, n_324);
  not g745 (n_325, n781);
  and g746 (n782, n_279, n_325);
  and g747 (n783, pi027, n768);
  not g748 (n_326, n782);
  not g749 (n_327, n783);
  and g750 (n784, n_326, n_327);
  and g754 (n787, n_305, n_310);
  and g755 (n788, n_269, n787);
  and g757 (n790, n_269, n_286);
  and g758 (n791, n_294, n737);
  not g759 (n_329, n790);
  not g760 (n_330, n791);
  and g761 (n792, n_329, n_330);
  not g762 (n_331, n792);
  and g763 (n793, n_283, n_331);
  and g764 (n794, pi026, n_294);
  and g765 (n795, n_269, pi027);
  not g766 (n_332, n794);
  not g767 (n_333, n795);
  and g768 (n796, n_332, n_333);
  not g769 (n_334, n796);
  and g770 (n797, n_265, n_334);
  not g771 (n_335, n793);
  not g772 (n_336, n797);
  and g773 (n798, n_335, n_336);
  not g774 (n_337, n798);
  and g775 (n799, pi028, n_337);
  and g779 (n803, n728, n737);
  not g780 (n_338, n802);
  not g781 (n_339, n803);
  and g782 (n804, n_338, n_339);
  not g783 (n_340, n804);
  and g784 (n805, n_294, n_340);
  and g785 (n806, n777, n790);
  not g786 (n_341, n805);
  not g787 (n_342, n806);
  and g788 (n807, n_341, n_342);
  not g789 (n_343, n799);
  and g790 (n808, n_343, n807);
  not g791 (n_344, n808);
  and g792 (n809, n_257, n_344);
  and g793 (n810, pi028, n_265);
  and g794 (n811, n_279, pi116);
  not g795 (n_345, n810);
  not g796 (n_346, n811);
  and g797 (n812, n_345, n_346);
  not g798 (n_347, n812);
  and g799 (n813, pi085, n_347);
  and g800 (n814, n_269, n_294);
  and g801 (n815, n813, n814);
  not g802 (n_348, n809);
  not g803 (n_349, n815);
  and g804 (n816, n_348, n_349);
  not g805 (n_350, n816);
  and g806 (n817, n_305, n_350);
  and g807 (n818, n_294, pi028);
  and g808 (n819, n_265, n818);
  and g809 (n820, n_269, n749);
  and g810 (n821, n819, n820);
  not g811 (n_351, n817);
  not g812 (n_352, n821);
  and g813 (n822, n_351, n_352);
  not g814 (n_353, n822);
  and g815 (n823, n_310, n_353);
  and g816 (n824, n743, n755);
  and g817 (n825, n819, n824);
  not g818 (n_354, n823);
  not g819 (n_355, n825);
  and g820 (n826, n_354, n_355);
  not g821 (n_356, n826);
  and g822 (n827, n_67, n_356);
  and g823 (po043, n_156, n827);
  and g824 (n829, pi029, pi110);
  and g825 (n830, pi097, n_258);
  and g826 (n831, n_260, n830);
  and g827 (n832, pi029, n_281);
  not g828 (n_357, n831);
  not g829 (n_358, n832);
  and g830 (n833, n_357, n_358);
  not g831 (n_359, n833);
  and g832 (n834, n724, n_359);
  not g833 (n_360, n829);
  not g834 (n_361, n834);
  and g835 (n835, n_360, n_361);
  not g836 (n_362, n835);
  and g837 (n836, n_310, n_362);
  and g838 (n837, pi097, pi116);
  and g839 (n838, pi029, n_265);
  not g840 (n_363, n837);
  not g841 (n_364, n838);
  and g842 (n839, n_363, n_364);
  not g843 (n_365, n839);
  and g844 (n840, pi058, n_365);
  not g845 (n_366, n836);
  not g846 (n_367, n840);
  and g847 (n841, n_366, n_367);
  not g848 (n_368, n841);
  and g849 (n842, n_305, n_368);
  and g850 (n843, pi053, n_310);
  and g851 (n844, n838, n843);
  not g852 (n_369, n842);
  not g853 (n_370, n844);
  and g854 (n845, n_369, n_370);
  not g855 (n_371, n845);
  and g856 (n846, n_294, n_371);
  and g857 (n847, pi027, n838);
  and g858 (n848, n787, n847);
  not g859 (n_372, n846);
  not g860 (n_373, n848);
  and g861 (n849, n_372, n_373);
  not g862 (n_374, n849);
  and g863 (n850, n_257, n_374);
  and g864 (n851, pi085, n774);
  and g865 (n852, n838, n851);
  not g866 (n_375, n850);
  not g867 (n_376, n852);
  and g868 (n853, n_375, n_376);
  not g869 (n_377, n853);
  and g870 (n854, n_269, n_377);
  and g871 (n855, n754, n787);
  and g872 (n856, pi026, n855);
  and g873 (n857, n838, n856);
  not g874 (n_378, n854);
  not g875 (n_379, n857);
  and g876 (n858, n_378, n_379);
  not g877 (n_380, n858);
  and g878 (n859, n_67, n_380);
  and g879 (po044, n_156, n859);
  not g880 (n_383, pi109);
  and g881 (n861, pi030, n_383);
  and g882 (n862, pi060, pi109);
  not g883 (n_385, n861);
  not g884 (n_386, n862);
  and g885 (n863, n_385, n_386);
  not g886 (n_388, pi106);
  not g887 (n_389, n863);
  and g888 (n864, n_388, n_389);
  and g889 (n865, pi088, pi106);
  not g890 (n_391, n864);
  not g891 (n_392, n865);
  and g892 (n866, n_391, n_392);
  not g893 (n_393, n866);
  and g894 (po045, n_67, n_393);
  and g895 (n868, pi089, pi106);
  and g896 (n869, pi030, pi109);
  and g897 (n870, pi031, n_383);
  not g898 (n_396, n869);
  not g899 (n_397, n870);
  and g900 (n871, n_396, n_397);
  not g901 (n_398, n871);
  and g902 (n872, n_388, n_398);
  not g903 (n_399, n868);
  not g904 (n_400, n872);
  and g905 (n873, n_399, n_400);
  not g906 (n_401, n873);
  and g907 (po046, n_67, n_401);
  and g908 (n875, pi099, pi106);
  and g909 (n876, pi031, pi109);
  and g910 (n877, pi032, n_383);
  not g911 (n_404, n876);
  not g912 (n_405, n877);
  and g913 (n878, n_404, n_405);
  not g914 (n_406, n878);
  and g915 (n879, n_388, n_406);
  not g916 (n_407, n875);
  not g917 (n_408, n879);
  and g918 (n880, n_407, n_408);
  not g919 (n_409, n880);
  and g920 (po047, n_67, n_409);
  and g921 (n882, pi090, pi106);
  and g922 (n883, pi032, pi109);
  and g923 (n884, pi033, n_383);
  not g924 (n_412, n883);
  not g925 (n_413, n884);
  and g926 (n885, n_412, n_413);
  not g927 (n_414, n885);
  and g928 (n886, n_388, n_414);
  not g929 (n_415, n882);
  not g930 (n_416, n886);
  and g931 (n887, n_415, n_416);
  not g932 (n_417, n887);
  and g933 (po048, n_67, n_417);
  and g934 (n889, pi091, pi106);
  and g935 (n890, pi033, pi109);
  and g936 (n891, pi034, n_383);
  not g937 (n_420, n890);
  not g938 (n_421, n891);
  and g939 (n892, n_420, n_421);
  not g940 (n_422, n892);
  and g941 (n893, n_388, n_422);
  not g942 (n_423, n889);
  not g943 (n_424, n893);
  and g944 (n894, n_423, n_424);
  not g945 (n_425, n894);
  and g946 (po049, n_67, n_425);
  and g947 (n896, pi092, pi106);
  and g948 (n897, pi034, pi109);
  and g949 (n898, pi035, n_383);
  not g950 (n_428, n897);
  not g951 (n_429, n898);
  and g952 (n899, n_428, n_429);
  not g953 (n_430, n899);
  and g954 (n900, n_388, n_430);
  not g955 (n_431, n896);
  not g956 (n_432, n900);
  and g957 (n901, n_431, n_432);
  not g958 (n_433, n901);
  and g959 (po050, n_67, n_433);
  and g960 (n903, pi098, pi106);
  and g961 (n904, pi035, pi109);
  and g962 (n905, pi036, n_383);
  not g963 (n_436, n904);
  not g964 (n_437, n905);
  and g965 (n906, n_436, n_437);
  not g966 (n_438, n906);
  and g967 (n907, n_388, n_438);
  not g968 (n_439, n903);
  not g969 (n_440, n907);
  and g970 (n908, n_439, n_440);
  not g971 (n_441, n908);
  and g972 (po051, n_67, n_441);
  and g973 (n910, pi093, pi106);
  and g974 (n911, pi036, pi109);
  and g975 (n912, pi037, n_383);
  not g976 (n_444, n911);
  not g977 (n_445, n912);
  and g978 (n913, n_444, n_445);
  not g979 (n_446, n913);
  and g980 (n914, n_388, n_446);
  not g981 (n_447, n910);
  not g982 (n_448, n914);
  and g983 (n915, n_447, n_448);
  not g984 (n_449, n915);
  and g985 (po052, n_67, n_449);
  not g986 (n_450, n391);
  and g987 (n917, pi082, n_450);
  and g988 (n918, n406, n579);
  and g989 (n919, n385, n697);
  and g990 (n920, n918, n919);
  not g991 (n_451, n920);
  and g992 (n921, pi082, n_451);
  not g993 (n_452, n921);
  and g994 (n922, n379, n_452);
  not g995 (n_453, n917);
  not g996 (n_454, n922);
  and g997 (n923, n_453, n_454);
  not g998 (n_455, n923);
  and g999 (n924, n_116, n_455);
  not g1006 (n_456, n930);
  and g1007 (n931, pi082, n_456);
  not g1008 (n_457, n931);
  and g1009 (n932, n_128, n_457);
  and g1010 (n933, pi074, n932);
  and g1011 (n934, n_121, pi082);
  and g1012 (n935, pi038, n641);
  and g1013 (n936, n934, n935);
  and g1020 (n940, n_273, pi109);
  and g1021 (n941, n736, n940);
  not g1022 (n_462, n941);
  and g1023 (n942, n_388, n_462);
  and g1024 (n943, pi109, n722);
  not g1025 (n_463, n943);
  and g1026 (n944, pi039, n_463);
  not g1027 (n_464, n944);
  and g1028 (n945, n942, n_464);
  not g1029 (n_465, n945);
  and g1030 (po054, n_67, n_465);
  not g1031 (n_466, n390);
  and g1032 (n947, pi082, n_466);
  and g1033 (n948, n579, n919);
  and g1034 (n949, n389, n948);
  not g1035 (n_467, n949);
  and g1036 (n950, pi082, n_467);
  not g1037 (n_468, n950);
  and g1038 (n951, n379, n_468);
  not g1039 (n_469, n947);
  not g1040 (n_470, n951);
  and g1041 (n952, n_469, n_470);
  not g1042 (n_471, n952);
  and g1043 (n953, n_123, n_471);
  not g1047 (n_472, n956);
  and g1048 (n957, pi082, n_472);
  not g1049 (n_473, n957);
  and g1050 (n958, n_128, n_473);
  and g1051 (n959, pi073, n958);
  and g1052 (n960, pi040, pi082);
  and g1053 (n961, n390, n960);
  not g1060 (n_478, n573);
  and g1061 (n965, pi082, n_478);
  not g1062 (n_479, n948);
  and g1063 (n966, pi082, n_479);
  not g1064 (n_480, n966);
  and g1065 (n967, n379, n_480);
  not g1066 (n_481, n965);
  not g1067 (n_482, n967);
  and g1068 (n968, n_481, n_482);
  not g1069 (n_483, n968);
  and g1070 (n969, n_112, n_483);
  not g1074 (n_484, n972);
  and g1075 (n973, pi082, n_484);
  not g1076 (n_485, n973);
  and g1077 (n974, n_128, n_485);
  and g1078 (n975, pi076, n974);
  and g1079 (n976, n403, n405);
  and g1089 (n983, pi044, pi082);
  and g1090 (n984, n688, n976);
  and g1091 (n985, n927, n984);
  not g1092 (n_490, n985);
  and g1093 (n986, pi082, n_490);
  not g1094 (n_491, n986);
  and g1095 (n987, n379, n_491);
  not g1096 (n_492, n983);
  not g1097 (n_493, n987);
  and g1098 (n988, n_492, n_493);
  not g1099 (n_494, n988);
  and g1100 (n989, n_120, n_494);
  and g1101 (n990, n_121, n649);
  and g1102 (n991, n638, n990);
  and g1103 (n992, n927, n991);
  not g1104 (n_495, n992);
  and g1105 (n993, pi082, n_495);
  not g1106 (n_496, n993);
  and g1107 (n994, n_128, n_496);
  and g1108 (n995, pi072, n994);
  and g1109 (n996, pi042, n934);
  not g1116 (n_501, n407);
  and g1117 (n1000, pi082, n_501);
  and g1118 (n1001, n385, n698);
  not g1119 (n_502, n1001);
  and g1120 (n1002, pi082, n_502);
  not g1121 (n_503, n1002);
  and g1122 (n1003, n379, n_503);
  not g1123 (n_504, n1000);
  not g1124 (n_505, n1003);
  and g1125 (n1004, n_504, n_505);
  not g1126 (n_506, n1004);
  and g1127 (n1005, n_100, n_506);
  and g1128 (n1006, n_101, n407);
  and g1129 (n1007, n927, n1006);
  not g1130 (n_507, n1007);
  and g1131 (n1008, pi082, n_507);
  not g1132 (n_508, n1008);
  and g1133 (n1009, n_128, n_508);
  and g1134 (n1010, pi077, n1009);
  and g1144 (n1017, n638, n642);
  and g1145 (n1018, n927, n1017);
  not g1146 (n_513, n1018);
  and g1147 (n1019, pi082, n_513);
  and g1148 (n1020, pi067, n_128);
  and g1149 (n1021, n_121, n379);
  not g1150 (n_515, n1020);
  not g1151 (n_516, n1021);
  and g1152 (n1022, n_515, n_516);
  not g1153 (n_517, n1019);
  not g1154 (n_518, n1022);
  and g1155 (n1023, n_517, n_518);
  and g1156 (n1024, n_67, n_492);
  not g1157 (n_519, n1023);
  and g1158 (po059, n_519, n1024);
  and g1159 (n1026, n399, n704);
  and g1160 (n1027, n388, n391);
  and g1161 (n1028, n1026, n1027);
  not g1162 (n_520, n1028);
  and g1163 (n1029, pi082, n_520);
  and g1164 (n1030, n_108, n692);
  not g1165 (n_521, n1030);
  and g1166 (n1031, pi082, n_521);
  not g1167 (n_522, n1031);
  and g1168 (n1032, n379, n_522);
  not g1169 (n_523, n1029);
  not g1170 (n_524, n1032);
  and g1171 (n1033, n_523, n_524);
  not g1172 (n_525, n1033);
  and g1173 (n1034, n_96, n_525);
  and g1174 (n1035, n_125, n399);
  and g1175 (n1036, n385, n1035);
  and g1176 (n1037, n408, n1036);
  not g1177 (n_526, n1037);
  and g1178 (n1038, pi082, n_526);
  not g1179 (n_527, n1038);
  and g1180 (n1039, n_128, n_527);
  and g1181 (n1040, pi068, n1039);
  and g1182 (n1041, n_116, n641);
  not g1192 (n_532, n1027);
  and g1193 (n1048, pi082, n_532);
  and g1194 (n1049, n688, n927);
  not g1195 (n_533, n1049);
  and g1196 (n1050, pi082, n_533);
  not g1197 (n_534, n1050);
  and g1198 (n1051, n379, n_534);
  not g1199 (n_535, n1048);
  not g1200 (n_536, n1051);
  and g1201 (n1052, n_535, n_536);
  not g1202 (n_537, n1052);
  and g1203 (n1053, n_113, n_537);
  and g1204 (n1054, n_117, n404);
  and g1205 (n1055, n1049, n1054);
  not g1206 (n_538, n1055);
  and g1207 (n1056, pi082, n_538);
  not g1208 (n_539, n1056);
  and g1209 (n1057, n_128, n_539);
  and g1210 (n1058, pi075, n1057);
  and g1211 (n1059, pi046, pi082);
  and g1212 (n1060, n1054, n1059);
  not g1219 (n_544, n408);
  and g1220 (n1064, pi082, n_544);
  not g1221 (n_545, n927);
  and g1222 (n1065, pi082, n_545);
  not g1223 (n_546, n1065);
  and g1224 (n1066, n379, n_546);
  not g1225 (n_547, n1064);
  not g1226 (n_548, n1066);
  and g1227 (n1067, n_547, n_548);
  not g1228 (n_549, n1067);
  and g1229 (n1068, n_101, n_549);
  and g1230 (n1069, n408, n927);
  not g1231 (n_550, n1069);
  and g1232 (n1070, pi082, n_550);
  not g1233 (n_551, n1070);
  and g1234 (n1071, n_128, n_551);
  and g1235 (n1072, pi064, n1071);
  and g1246 (n1080, n638, n1027);
  not g1247 (n_556, n1080);
  and g1248 (n1081, pi082, n_556);
  not g1249 (n_557, n919);
  and g1250 (n1082, pi082, n_557);
  not g1251 (n_558, n1082);
  and g1252 (n1083, n379, n_558);
  not g1253 (n_559, n1081);
  not g1254 (n_560, n1083);
  and g1255 (n1084, n_559, n_560);
  not g1256 (n_561, n1084);
  and g1257 (n1085, n_97, n_561);
  and g1259 (n1087, n398, n401);
  not g1262 (n_562, n1089);
  and g1263 (n1090, pi082, n_562);
  not g1264 (n_563, n1090);
  and g1265 (n1091, n_128, n_563);
  and g1266 (n1092, pi062, n1091);
  and g1277 (n1100, n384, n1054);
  and g1278 (n1101, n705, n1100);
  not g1279 (n_568, n1101);
  and g1280 (n1102, pi082, n_568);
  not g1281 (n_569, n1102);
  and g1282 (n1103, n_128, n_569);
  not g1283 (n_571, pi069);
  and g1284 (n1104, n_571, n1103);
  not g1288 (n_572, n1107);
  and g1289 (n1108, pi049, n_572);
  and g1290 (n1109, n_125, n383);
  not g1295 (n_574, n1108);
  not g1296 (n_575, n1112);
  and g1297 (n1113, n_574, n_575);
  not g1298 (n_576, n1113);
  and g1299 (n1114, pi082, n_576);
  and g1300 (n1115, pi049, n411);
  not g1301 (n_577, n1114);
  not g1302 (n_578, n1115);
  and g1303 (n1116, n_577, n_578);
  not g1304 (n_579, n1104);
  and g1305 (n1117, n_579, n1116);
  not g1306 (n_580, n1117);
  and g1307 (po064, n_67, n_580);
  not g1308 (n_581, n404);
  and g1309 (n1119, pi082, n_581);
  and g1310 (n1120, n704, n1035);
  and g1311 (n1121, n1087, n1120);
  not g1312 (n_582, n1121);
  and g1313 (n1122, pi082, n_582);
  not g1314 (n_583, n1122);
  and g1315 (n1123, n379, n_583);
  not g1316 (n_584, n1119);
  not g1317 (n_585, n1123);
  and g1318 (n1124, n_584, n_585);
  not g1319 (n_586, n1124);
  and g1320 (n1125, n_117, n_586);
  and g1321 (n1126, n404, n638);
  and g1322 (n1127, n927, n1126);
  not g1323 (n_587, n1127);
  and g1324 (n1128, pi082, n_587);
  not g1325 (n_588, n1128);
  and g1326 (n1129, n_128, n_588);
  and g1327 (n1130, pi066, n1129);
  and g1328 (n1131, pi050, n1041);
  and g1329 (n1132, n934, n1131);
  and g1336 (n1136, pi051, n_383);
  not g1337 (n_593, n940);
  not g1338 (n_594, n1136);
  and g1339 (n1137, n_593, n_594);
  and g1340 (n1138, n_388, n1137);
  not g1341 (n_595, n1138);
  and g1342 (po066, n_67, n_595);
  and g1343 (n1140, pi052, n_593);
  and g1344 (n1141, n_388, n_463);
  not g1345 (n_596, n1140);
  and g1346 (n1142, n_596, n1141);
  not g1347 (n_597, n1142);
  and g1348 (po067, n_67, n_597);
  and g1349 (n1144, pi058, pi116);
  not g1353 (n_598, n1144);
  not g1354 (n_599, n1147);
  and g1355 (n1148, n_598, n_599);
  not g1356 (n_600, n1148);
  and g1357 (n1149, n_305, n_600);
  and g1358 (n1150, pi097, n1149);
  and g1359 (n1151, n_265, n843);
  not g1360 (n_601, n1150);
  not g1361 (n_602, n1151);
  and g1362 (n1152, n_601, n_602);
  and g1368 (n1157, n408, n1001);
  not g1369 (n_604, n1157);
  and g1370 (n1158, pi082, n_604);
  not g1371 (n_605, n1158);
  and g1372 (n1159, n_128, n_605);
  or g1373 (po069, pi129, n1159);
  or g1374 (po129, pi123, pi129);
  not g1375 (n_607, pi122);
  and g1376 (n1162, pi114, n_607);
  not g1377 (n_609, po129);
  and g1378 (po070, n_609, n1162);
  and g1379 (n1164, n_269, pi058);
  and g1380 (n1165, pi026, n_310);
  and g1381 (n1166, pi116, n1165);
  not g1382 (n_610, n1164);
  not g1383 (n_611, n1166);
  and g1384 (n1167, n_610, n_611);
  not g1385 (n_613, n1167);
  and g1386 (n1168, pi094, n_613);
  and g1387 (n1169, pi058, n_265);
  and g1388 (n1170, pi037, n_265);
  not g1389 (n_614, n1170);
  and g1390 (n1171, n_610, n_614);
  not g1391 (n_615, n1169);
  not g1392 (n_616, n1171);
  and g1393 (n1172, n_615, n_616);
  not g1394 (n_617, n1168);
  not g1395 (n_618, n1172);
  and g1396 (n1173, n_617, n_618);
  not g1397 (n_619, n1173);
  and g1398 (n1174, n_305, n_619);
  and g1399 (n1175, n_269, pi037);
  and g1400 (n1176, n_310, n1175);
  not g1401 (n_620, n1174);
  not g1402 (n_621, n1176);
  and g1403 (n1177, n_620, n_621);
  not g1404 (n_622, n1177);
  and g1405 (n1178, n_257, n_622);
  and g1406 (n1179, n787, n1175);
  not g1407 (n_623, n1178);
  not g1408 (n_624, n1179);
  and g1409 (n1180, n_623, n_624);
  not g1410 (n_625, n1180);
  and g1411 (n1181, n_294, n_625);
  and g1412 (n1182, n_257, n787);
  and g1413 (n1183, n1175, n1182);
  not g1414 (n_626, n1181);
  not g1415 (n_627, n1183);
  and g1416 (n1184, n_626, n_627);
  not g1417 (n_628, n1184);
  and g1418 (n1185, n_67, n_628);
  and g1419 (po071, n_156, n1185);
  and g1420 (n1187, n_269, n_305);
  and g1421 (n1188, pi026, pi053);
  not g1422 (n_629, n1188);
  and g1423 (n1189, n_257, n_629);
  not g1424 (n_630, n1187);
  not g1425 (n_631, n1189);
  and g1426 (n1190, n_630, n_631);
  not g1427 (n_632, n1190);
  and g1428 (n1191, n_310, n_632);
  and g1429 (n1192, n_257, n1187);
  and g1430 (n1193, n_265, n1192);
  not g1431 (n_633, n1191);
  not g1432 (n_634, n1193);
  and g1433 (n1194, n_633, n_634);
  not g1434 (n_636, n1194);
  and g1435 (n1195, pi057, n_636);
  and g1436 (n1196, pi060, n1144);
  and g1437 (n1197, n1192, n1196);
  not g1438 (n_637, n1195);
  not g1439 (n_638, n1197);
  and g1440 (n1198, n_637, n_638);
  not g1441 (n_639, n1198);
  and g1442 (n1199, n_294, n_639);
  and g1443 (n1200, pi057, n_310);
  and g1444 (n1201, n1192, n1200);
  not g1445 (n_640, n1199);
  not g1446 (n_641, n1201);
  and g1447 (n1202, n_640, n_641);
  not g1448 (n_642, n1202);
  and g1449 (n1203, n_67, n_642);
  and g1450 (po072, n_156, n1203);
  and g1451 (n1205, n814, n1169);
  not g1455 (n_643, n1205);
  not g1456 (n_644, n1208);
  and g1457 (n1209, n_643, n_644);
  not g1463 (n_646, n755);
  not g1464 (n_647, n843);
  and g1465 (n1214, n_646, n_647);
  not g1466 (n_648, n1214);
  and g1467 (n1215, n_265, n_648);
  and g1468 (n1216, n_283, n787);
  not g1469 (n_649, n1215);
  not g1470 (n_650, n1216);
  and g1471 (n1217, n_649, n_650);
  not g1472 (n_651, n1217);
  and g1473 (n1218, pi059, n_651);
  and g1474 (n1219, n726, n787);
  and g1475 (n1220, pi096, n1219);
  not g1476 (n_652, n1218);
  not g1477 (n_653, n1220);
  and g1478 (n1221, n_652, n_653);
  not g1479 (n_654, n1221);
  and g1480 (n1222, n_257, n_654);
  and g1481 (n1223, pi059, n_265);
  and g1482 (n1224, pi085, n787);
  and g1483 (n1225, n1223, n1224);
  not g1484 (n_655, n1222);
  not g1485 (n_656, n1225);
  and g1486 (n1226, n_655, n_656);
  not g1487 (n_657, n1226);
  and g1488 (n1227, n_294, n_657);
  and g1489 (n1228, pi027, n1182);
  and g1490 (n1229, n1223, n1228);
  not g1491 (n_658, n1227);
  not g1492 (n_659, n1229);
  and g1493 (n1230, n_658, n_659);
  not g1494 (n_660, n1230);
  and g1495 (n1231, n_269, n_660);
  and g1496 (n1232, n856, n1223);
  not g1497 (n_661, n1231);
  not g1498 (n_662, n1232);
  and g1499 (n1233, n_661, n_662);
  not g1500 (n_663, n1233);
  and g1501 (n1234, n_67, n_663);
  and g1502 (po074, n_156, n1234);
  not g1503 (n_665, pi117);
  and g1504 (n1236, n_665, n_607);
  not g1505 (n_666, n1236);
  and g1506 (n1237, pi060, n_666);
  and g1507 (n1238, pi123, n1236);
  or g1508 (po075, n1237, n1238);
  not g1513 (n_670, pi137);
  not g1514 (n_671, pi138);
  and g1517 (n1245, pi132, pi133);
  and g1518 (n1246, pi131, n1245);
  not g1520 (n_676, n1247);
  and g1521 (n1248, pi062, n_676);
  and g1522 (n1249, pi136, n_670);
  not g1523 (n_678, pi140);
  and g1524 (n1250, n_678, n1249);
  and g1525 (n1251, n_671, n1246);
  and g1526 (n1252, n1250, n1251);
  not g1527 (n_679, n1248);
  not g1528 (n_680, n1252);
  and g1529 (n1253, n_679, n_680);
  or g1530 (po077, pi129, n1253);
  and g1531 (n1255, pi063, n_676);
  not g1532 (n_682, pi142);
  and g1533 (n1256, n_682, n1249);
  and g1534 (n1257, n1251, n1256);
  not g1535 (n_683, n1255);
  not g1536 (n_684, n1257);
  and g1537 (n1258, n_683, n_684);
  or g1538 (po078, pi129, n1258);
  and g1539 (n1260, pi064, n_676);
  not g1540 (n_686, pi139);
  and g1541 (n1261, n_686, n1249);
  and g1542 (n1262, n1251, n1261);
  not g1543 (n_687, n1260);
  not g1544 (n_688, n1262);
  and g1545 (n1263, n_687, n_688);
  or g1546 (po079, pi129, n1263);
  and g1547 (n1265, pi065, n_676);
  not g1548 (n_690, pi146);
  and g1549 (n1266, n_690, n1249);
  and g1550 (n1267, n1251, n1266);
  not g1551 (n_691, n1265);
  not g1552 (n_692, n1267);
  and g1553 (n1268, n_691, n_692);
  or g1554 (po080, pi129, n1268);
  not g1555 (n_693, pi136);
  and g1556 (n1270, n_693, n_670);
  and g1557 (n1271, n1251, n1270);
  not g1558 (n_694, n1271);
  and g1559 (n1272, pi066, n_694);
  not g1560 (n_696, pi143);
  and g1561 (n1273, n_696, n1271);
  not g1562 (n_697, n1272);
  not g1563 (n_698, n1273);
  and g1564 (n1274, n_697, n_698);
  or g1565 (po081, pi129, n1274);
  and g1566 (n1276, pi067, n_694);
  and g1567 (n1277, n_686, n1271);
  not g1568 (n_699, n1276);
  not g1569 (n_700, n1277);
  and g1570 (n1278, n_699, n_700);
  or g1571 (po082, pi129, n1278);
  and g1572 (n1280, pi068, n_676);
  not g1573 (n_702, pi141);
  and g1574 (n1281, n_702, n1249);
  and g1575 (n1282, n1251, n1281);
  not g1576 (n_703, n1280);
  not g1577 (n_704, n1282);
  and g1578 (n1283, n_703, n_704);
  or g1579 (po083, pi129, n1283);
  and g1580 (n1285, pi069, n_676);
  and g1581 (n1286, n_696, n1249);
  and g1582 (n1287, n1251, n1286);
  not g1583 (n_705, n1285);
  not g1584 (n_706, n1287);
  and g1585 (n1288, n_705, n_706);
  or g1586 (po084, pi129, n1288);
  and g1587 (n1290, pi070, n_676);
  not g1588 (n_708, pi144);
  and g1589 (n1291, n_708, n1249);
  and g1590 (n1292, n1251, n1291);
  not g1591 (n_709, n1290);
  not g1592 (n_710, n1292);
  and g1593 (n1293, n_709, n_710);
  or g1594 (po085, pi129, n1293);
  and g1595 (n1295, pi071, n_676);
  not g1596 (n_712, pi145);
  and g1597 (n1296, n_712, n1249);
  and g1598 (n1297, n1251, n1296);
  not g1599 (n_713, n1295);
  not g1600 (n_714, n1297);
  and g1601 (n1298, n_713, n_714);
  or g1602 (po086, pi129, n1298);
  and g1603 (n1300, pi072, n_694);
  and g1604 (n1301, n_678, n1271);
  not g1605 (n_715, n1300);
  not g1606 (n_716, n1301);
  and g1607 (n1302, n_715, n_716);
  or g1608 (po087, pi129, n1302);
  and g1609 (n1304, pi073, n_694);
  and g1610 (n1305, n_702, n1271);
  not g1611 (n_717, n1304);
  not g1612 (n_718, n1305);
  and g1613 (n1306, n_717, n_718);
  or g1614 (po088, pi129, n1306);
  and g1615 (n1308, pi074, n_694);
  and g1616 (n1309, n_682, n1271);
  not g1617 (n_719, n1308);
  not g1618 (n_720, n1309);
  and g1619 (n1310, n_719, n_720);
  or g1620 (po089, pi129, n1310);
  and g1621 (n1312, pi075, n_694);
  and g1622 (n1313, n_708, n1271);
  not g1623 (n_721, n1312);
  not g1624 (n_722, n1313);
  and g1625 (n1314, n_721, n_722);
  or g1626 (po090, pi129, n1314);
  and g1627 (n1316, pi076, n_694);
  and g1628 (n1317, n_712, n1271);
  not g1629 (n_723, n1316);
  not g1630 (n_724, n1317);
  and g1631 (n1318, n_723, n_724);
  or g1632 (po091, pi129, n1318);
  and g1633 (n1320, pi077, n_694);
  and g1634 (n1321, n_690, n1271);
  not g1635 (n_725, n1320);
  not g1636 (n_726, n1321);
  and g1637 (n1322, n_725, n_726);
  or g1638 (po092, pi129, n1322);
  and g1639 (n1324, n_693, pi137);
  and g1640 (n1325, n1251, n1324);
  not g1641 (n_728, n1325);
  and g1642 (n1326, pi078, n_728);
  and g1643 (n1327, pi142, n1325);
  not g1644 (n_729, n1326);
  not g1645 (n_730, n1327);
  and g1646 (n1328, n_729, n_730);
  not g1647 (n_731, n1328);
  and g1648 (po093, n_67, n_731);
  and g1649 (n1330, pi079, n_728);
  and g1650 (n1331, pi143, n1325);
  not g1651 (n_733, n1330);
  not g1652 (n_734, n1331);
  and g1653 (n1332, n_733, n_734);
  not g1654 (n_735, n1332);
  and g1655 (po094, n_67, n_735);
  and g1656 (n1334, pi080, n_728);
  and g1657 (n1335, pi144, n1325);
  not g1658 (n_737, n1334);
  not g1659 (n_738, n1335);
  and g1660 (n1336, n_737, n_738);
  not g1661 (n_739, n1336);
  and g1662 (po095, n_67, n_739);
  and g1663 (n1338, pi081, n_728);
  and g1664 (n1339, pi145, n1325);
  not g1665 (n_741, n1338);
  not g1666 (n_742, n1339);
  and g1667 (n1340, n_741, n_742);
  not g1668 (n_743, n1340);
  and g1669 (po096, n_67, n_743);
  and g1670 (n1342, pi082, n_728);
  and g1671 (n1343, pi146, n1325);
  not g1672 (n_744, n1342);
  not g1673 (n_745, n1343);
  and g1674 (n1344, n_744, n_745);
  not g1675 (n_746, n1344);
  and g1676 (po097, n_67, n_746);
  and g1677 (n1346, pi089, pi138);
  not g1678 (n_747, pi062);
  and g1679 (n1347, n_747, n_671);
  not g1680 (n_748, n1346);
  not g1681 (n_749, n1347);
  and g1682 (n1348, n_748, n_749);
  not g1683 (n_750, n1348);
  and g1684 (n1349, pi136, n_750);
  and g1685 (n1350, pi119, pi138);
  not g1686 (n_752, pi072);
  and g1687 (n1351, n_752, n_671);
  not g1688 (n_753, n1350);
  not g1689 (n_754, n1351);
  and g1690 (n1352, n_753, n_754);
  not g1691 (n_755, n1352);
  and g1692 (n1353, n_693, n_755);
  not g1693 (n_756, n1349);
  not g1694 (n_757, n1353);
  and g1695 (n1354, n_756, n_757);
  not g1696 (n_758, n1354);
  and g1697 (n1355, n_670, n_758);
  not g1698 (n_760, pi115);
  and g1699 (n1356, n_760, pi138);
  and g1700 (n1357, pi087, n_671);
  not g1701 (n_762, n1356);
  not g1702 (n_763, n1357);
  and g1703 (n1358, n_762, n_763);
  not g1704 (n_764, n1358);
  and g1705 (n1359, n_693, n_764);
  and g1706 (n1360, pi136, n_671);
  and g1707 (n1361, pi031, n1360);
  not g1708 (n_765, n1359);
  not g1709 (n_766, n1361);
  and g1710 (n1362, n_765, n_766);
  not g1711 (n_767, n1362);
  and g1712 (n1363, pi137, n_767);
  or g1713 (po098, n1355, n1363);
  and g1714 (n1365, pi084, n_728);
  and g1715 (n1366, pi141, n1325);
  not g1716 (n_769, n1365);
  not g1717 (n_770, n1366);
  and g1718 (n1367, n_769, n_770);
  not g1719 (n_771, n1367);
  and g1720 (po099, n_67, n_771);
  and g1721 (n1369, n_257, n_282);
  and g1722 (n1370, n_258, n1369);
  and g1723 (n1371, pi096, n1370);
  not g1724 (n_772, n1371);
  and g1725 (n1372, n_315, n_772);
  and g1731 (n1377, pi086, n_728);
  and g1732 (n1378, pi139, n1325);
  not g1733 (n_775, n1377);
  not g1734 (n_776, n1378);
  and g1735 (n1379, n_775, n_776);
  not g1736 (n_777, n1379);
  and g1737 (po101, n_67, n_777);
  and g1738 (n1381, pi087, n_728);
  and g1739 (n1382, pi140, n1325);
  not g1740 (n_778, n1381);
  not g1741 (n_779, n1382);
  and g1742 (n1383, n_778, n_779);
  not g1743 (n_780, n1383);
  and g1744 (po102, n_67, n_780);
  and g1745 (n1385, pi136, pi137);
  and g1746 (n1386, n1251, n1385);
  not g1747 (n_781, n1386);
  and g1748 (n1387, pi088, n_781);
  and g1749 (n1388, pi139, n1386);
  not g1750 (n_782, n1387);
  not g1751 (n_783, n1388);
  and g1752 (n1389, n_782, n_783);
  not g1753 (n_784, n1389);
  and g1754 (po103, n_67, n_784);
  and g1755 (n1391, pi089, n_781);
  and g1756 (n1392, pi140, n1386);
  not g1757 (n_785, n1391);
  not g1758 (n_786, n1392);
  and g1759 (n1393, n_785, n_786);
  not g1760 (n_787, n1393);
  and g1761 (po104, n_67, n_787);
  and g1762 (n1395, pi090, n_781);
  and g1763 (n1396, pi142, n1386);
  not g1764 (n_788, n1395);
  not g1765 (n_789, n1396);
  and g1766 (n1397, n_788, n_789);
  not g1767 (n_790, n1397);
  and g1768 (po105, n_67, n_790);
  and g1769 (n1399, pi091, n_781);
  and g1770 (n1400, pi143, n1386);
  not g1771 (n_791, n1399);
  not g1772 (n_792, n1400);
  and g1773 (n1401, n_791, n_792);
  not g1774 (n_793, n1401);
  and g1775 (po106, n_67, n_793);
  and g1776 (n1403, pi092, n_781);
  and g1777 (n1404, pi144, n1386);
  not g1778 (n_794, n1403);
  not g1779 (n_795, n1404);
  and g1780 (n1405, n_794, n_795);
  not g1781 (n_796, n1405);
  and g1782 (po107, n_67, n_796);
  and g1783 (n1407, pi093, n_781);
  and g1784 (n1408, pi146, n1386);
  not g1785 (n_797, n1407);
  not g1786 (n_798, n1408);
  and g1787 (n1409, n_797, n_798);
  not g1788 (n_799, n1409);
  and g1789 (po108, n_67, n_799);
  and g1790 (n1411, pi082, n_670);
  and g1791 (n1412, n_693, n1411);
  and g1792 (n1413, pi138, n1246);
  and g1793 (n1414, n1412, n1413);
  not g1794 (n_800, n1414);
  and g1795 (n1415, pi094, n_800);
  and g1796 (n1416, pi142, n1414);
  not g1797 (n_801, n1415);
  not g1798 (n_802, n1416);
  and g1799 (n1417, n_801, n_802);
  not g1800 (n_803, n1417);
  and g1801 (po109, n_67, n_803);
  not g1802 (n_804, n1246);
  and g1803 (n1419, n_156, n_804);
  and g1804 (n1420, n_258, n1419);
  and g1805 (n1421, pi138, n1412);
  not g1806 (n_805, n1421);
  and g1807 (n1422, n1246, n_805);
  not g1808 (n_806, n1420);
  not g1809 (n_807, n1422);
  and g1810 (n1423, n_806, n_807);
  not g1811 (n_808, n1423);
  and g1812 (n1424, pi095, n_808);
  and g1813 (n1425, pi143, n1414);
  not g1814 (n_809, n1424);
  not g1815 (n_810, n1425);
  and g1816 (n1426, n_809, n_810);
  not g1817 (n_811, n1426);
  and g1818 (po110, n_67, n_811);
  and g1819 (n1428, pi096, n_808);
  and g1820 (n1429, pi146, n1414);
  not g1821 (n_812, n1428);
  not g1822 (n_813, n1429);
  and g1823 (n1430, n_812, n_813);
  not g1824 (n_814, n1430);
  and g1825 (po111, n_67, n_814);
  and g1826 (n1432, pi097, n_808);
  and g1827 (n1433, pi145, n1414);
  not g1828 (n_815, n1432);
  not g1829 (n_816, n1433);
  and g1830 (n1434, n_815, n_816);
  not g1831 (n_817, n1434);
  and g1832 (po112, n_67, n_817);
  and g1833 (n1436, pi098, n_781);
  and g1834 (n1437, pi145, n1386);
  not g1835 (n_818, n1436);
  not g1836 (n_819, n1437);
  and g1837 (n1438, n_818, n_819);
  not g1838 (n_820, n1438);
  and g1839 (po113, n_67, n_820);
  and g1840 (n1440, pi099, n_781);
  and g1841 (n1441, pi141, n1386);
  not g1842 (n_821, n1440);
  not g1843 (n_822, n1441);
  and g1844 (n1442, n_821, n_822);
  not g1845 (n_823, n1442);
  and g1846 (po114, n_67, n_823);
  and g1847 (n1444, pi100, n_808);
  and g1848 (n1445, pi144, n1414);
  not g1849 (n_824, n1444);
  not g1850 (n_825, n1445);
  and g1851 (n1446, n_824, n_825);
  not g1852 (n_826, n1446);
  and g1853 (po115, n_67, n_826);
  and g1854 (n1448, pi124, pi138);
  not g1855 (n_828, pi077);
  and g1856 (n1449, n_828, n_671);
  not g1857 (n_829, n1448);
  not g1858 (n_830, n1449);
  and g1859 (n1450, n_829, n_830);
  not g1860 (n_831, n1450);
  and g1861 (n1451, n_693, n_831);
  and g1862 (n1452, n_131, n_671);
  and g1863 (n1453, pi093, pi138);
  not g1864 (n_832, n1452);
  not g1865 (n_833, n1453);
  and g1866 (n1454, n_832, n_833);
  not g1867 (n_834, n1454);
  and g1868 (n1455, pi136, n_834);
  not g1869 (n_835, n1451);
  not g1870 (n_836, n1455);
  and g1871 (n1456, n_835, n_836);
  not g1872 (n_837, n1456);
  and g1873 (n1457, n_670, n_837);
  and g1874 (n1458, pi037, n1360);
  and g1875 (n1459, pi096, pi138);
  and g1876 (n1460, pi082, n_671);
  not g1877 (n_838, n1459);
  not g1878 (n_839, n1460);
  and g1879 (n1461, n_838, n_839);
  not g1880 (n_840, n1461);
  and g1881 (n1462, n_693, n_840);
  not g1882 (n_841, n1458);
  not g1883 (n_842, n1462);
  and g1884 (n1463, n_841, n_842);
  not g1885 (n_843, n1463);
  and g1886 (n1464, pi137, n_843);
  or g1887 (po116, n1457, n1464);
  and g1888 (n1466, pi091, n1249);
  and g1889 (n1467, pi095, n1324);
  not g1890 (n_844, n1466);
  not g1891 (n_845, n1467);
  and g1892 (n1468, n_844, n_845);
  not g1893 (n_846, n1468);
  and g1894 (n1469, pi138, n_846);
  and g1895 (n1470, pi079, n_693);
  and g1896 (n1471, pi034, pi136);
  not g1897 (n_847, n1470);
  not g1898 (n_848, n1471);
  and g1899 (n1472, n_847, n_848);
  not g1900 (n_849, n1472);
  and g1901 (n1473, pi137, n_849);
  and g1902 (n1474, n_571, pi136);
  not g1903 (n_850, pi066);
  and g1904 (n1475, n_850, n_693);
  not g1905 (n_851, n1474);
  not g1906 (n_852, n1475);
  and g1907 (n1476, n_851, n_852);
  not g1908 (n_853, n1476);
  and g1909 (n1477, n_670, n_853);
  not g1910 (n_854, n1473);
  not g1911 (n_855, n1477);
  and g1912 (n1478, n_854, n_855);
  not g1913 (n_856, n1478);
  and g1914 (n1479, n_671, n_856);
  or g1915 (po117, n1469, n1479);
  and g1916 (n1481, pi090, n1249);
  and g1917 (n1482, pi094, n1324);
  not g1918 (n_857, n1481);
  not g1919 (n_858, n1482);
  and g1920 (n1483, n_857, n_858);
  not g1921 (n_859, n1483);
  and g1922 (n1484, pi138, n_859);
  and g1923 (n1485, pi078, n_693);
  and g1924 (n1486, pi033, pi136);
  not g1925 (n_860, n1485);
  not g1926 (n_861, n1486);
  and g1927 (n1487, n_860, n_861);
  not g1928 (n_862, n1487);
  and g1929 (n1488, pi137, n_862);
  not g1930 (n_863, pi063);
  and g1931 (n1489, n_863, pi136);
  not g1932 (n_864, pi074);
  and g1933 (n1490, n_864, n_693);
  not g1934 (n_865, n1489);
  not g1935 (n_866, n1490);
  and g1936 (n1491, n_865, n_866);
  not g1937 (n_867, n1491);
  and g1938 (n1492, n_670, n_867);
  not g1939 (n_868, n1488);
  not g1940 (n_869, n1492);
  and g1941 (n1493, n_868, n_869);
  not g1942 (n_870, n1493);
  and g1943 (n1494, n_671, n_870);
  or g1944 (po118, n1484, n1494);
  and g1945 (n1496, pi099, n1249);
  not g1946 (n_872, pi112);
  and g1947 (n1497, n_872, n1324);
  not g1948 (n_873, n1496);
  not g1949 (n_874, n1497);
  and g1950 (n1498, n_873, n_874);
  not g1951 (n_875, n1498);
  and g1952 (n1499, pi138, n_875);
  not g1953 (n_876, pi068);
  and g1954 (n1500, n_876, pi136);
  not g1955 (n_877, pi073);
  and g1956 (n1501, n_877, n_693);
  not g1957 (n_878, n1500);
  not g1958 (n_879, n1501);
  and g1959 (n1502, n_878, n_879);
  not g1960 (n_880, n1502);
  and g1961 (n1503, n_670, n_880);
  and g1962 (n1504, pi084, n_693);
  and g1963 (n1505, pi032, pi136);
  not g1964 (n_881, n1504);
  not g1965 (n_882, n1505);
  and g1966 (n1506, n_881, n_882);
  not g1967 (n_883, n1506);
  and g1968 (n1507, pi137, n_883);
  not g1969 (n_884, n1503);
  not g1970 (n_885, n1507);
  and g1971 (n1508, n_884, n_885);
  not g1972 (n_886, n1508);
  and g1973 (n1509, n_671, n_886);
  or g1974 (po119, n1499, n1509);
  and g1975 (n1511, pi092, pi138);
  and g1976 (n1512, n_198, n_671);
  not g1977 (n_887, n1511);
  not g1978 (n_888, n1512);
  and g1979 (n1513, n_887, n_888);
  not g1980 (n_889, n1513);
  and g1981 (n1514, pi136, n_889);
  and g1982 (n1515, pi125, pi138);
  not g1983 (n_891, pi075);
  and g1984 (n1516, n_891, n_671);
  not g1985 (n_892, n1515);
  not g1986 (n_893, n1516);
  and g1987 (n1517, n_892, n_893);
  not g1988 (n_894, n1517);
  and g1989 (n1518, n_693, n_894);
  not g1990 (n_895, n1514);
  not g1991 (n_896, n1518);
  and g1992 (n1519, n_895, n_896);
  not g1993 (n_897, n1519);
  and g1994 (n1520, n_670, n_897);
  and g1995 (n1521, pi080, n_671);
  and g1996 (n1522, pi100, pi138);
  not g1997 (n_898, n1521);
  not g1998 (n_899, n1522);
  and g1999 (n1523, n_898, n_899);
  not g2000 (n_900, n1523);
  and g2001 (n1524, n_693, n_900);
  and g2002 (n1525, pi035, n1360);
  not g2003 (n_901, n1524);
  not g2004 (n_902, n1525);
  and g2005 (n1526, n_901, n_902);
  not g2006 (n_903, n1526);
  and g2007 (n1527, pi137, n_903);
  or g2008 (po120, n1520, n1527);
  and g2009 (n1529, n788, n1370);
  and g2010 (n1530, n_294, n1529);
  not g2011 (n_904, n1530);
  and g2012 (n1531, n_261, n_904);
  not g2013 (n_905, n1531);
  and g2014 (n1532, n_67, n_905);
  and g2015 (po121, n_156, n1532);
  and g2016 (n1534, pi098, pi138);
  and g2017 (n1535, n_223, n_671);
  not g2018 (n_906, n1534);
  not g2019 (n_907, n1535);
  and g2020 (n1536, n_906, n_907);
  not g2021 (n_908, n1536);
  and g2022 (n1537, pi136, n_908);
  not g2023 (n_909, pi076);
  and g2024 (n1538, n_909, n_671);
  and g2025 (n1539, pi023, pi138);
  not g2026 (n_910, n1538);
  not g2027 (n_911, n1539);
  and g2028 (n1540, n_910, n_911);
  not g2029 (n_912, n1540);
  and g2030 (n1541, n_693, n_912);
  not g2031 (n_913, n1537);
  not g2032 (n_914, n1541);
  and g2033 (n1542, n_913, n_914);
  not g2034 (n_915, n1542);
  and g2035 (n1543, n_670, n_915);
  and g2036 (n1544, pi036, n1360);
  and g2037 (n1545, pi081, n_671);
  and g2038 (n1546, pi097, pi138);
  not g2039 (n_916, n1545);
  not g2040 (n_917, n1546);
  and g2041 (n1547, n_916, n_917);
  not g2042 (n_918, n1547);
  and g2043 (n1548, n_693, n_918);
  not g2044 (n_919, n1544);
  not g2045 (n_920, n1548);
  and g2046 (n1549, n_919, n_920);
  not g2047 (n_921, n1549);
  and g2048 (n1550, pi137, n_921);
  or g2049 (po122, n1543, n1550);
  and g2050 (n1552, pi088, pi138);
  not g2051 (n_922, pi064);
  and g2052 (n1553, n_922, n_671);
  not g2053 (n_923, n1552);
  not g2054 (n_924, n1553);
  and g2055 (n1554, n_923, n_924);
  not g2056 (n_925, n1554);
  and g2057 (n1555, pi136, n_925);
  and g2058 (n1556, pi120, pi138);
  not g2059 (n_927, pi067);
  and g2060 (n1557, n_927, n_671);
  not g2061 (n_928, n1556);
  not g2062 (n_929, n1557);
  and g2063 (n1558, n_928, n_929);
  not g2064 (n_930, n1558);
  and g2065 (n1559, n_693, n_930);
  not g2066 (n_931, n1555);
  not g2067 (n_932, n1559);
  and g2068 (n1560, n_931, n_932);
  not g2069 (n_933, n1560);
  and g2070 (n1561, n_670, n_933);
  and g2071 (n1562, pi086, n_671);
  and g2072 (n1563, pi111, pi138);
  not g2073 (n_935, n1562);
  not g2074 (n_936, n1563);
  and g2075 (n1564, n_935, n_936);
  not g2076 (n_937, n1564);
  and g2077 (n1565, n_693, n_937);
  and g2078 (n1566, pi030, n1360);
  not g2079 (n_938, n1565);
  not g2080 (n_939, n1566);
  and g2081 (n1567, n_938, n_939);
  not g2082 (n_940, n1567);
  and g2083 (n1568, pi137, n_940);
  or g2084 (po123, n1561, n1568);
  not g2085 (n_941, n737);
  and g2086 (n1570, n_941, n795);
  not g2087 (n_942, n1570);
  and g2088 (n1571, n_332, n_942);
  and g2093 (n1575, n_281, n755);
  not g2094 (n_944, n1575);
  and g2095 (n1576, n_647, n_944);
  and g2100 (n1580, pi111, n_805);
  and g2101 (n1581, n_693, pi139);
  and g2102 (n1582, n_670, pi138);
  and g2103 (n1583, pi082, n1582);
  and g2104 (n1584, n1581, n1583);
  not g2105 (n_946, n1580);
  not g2106 (n_947, n1584);
  and g2107 (n1585, n_946, n_947);
  not g2108 (n_948, n1585);
  and g2109 (n1586, n1246, n_948);
  and g2110 (po126, n_67, n1586);
  and g2111 (n1588, n_693, pi141);
  and g2112 (n1589, n1583, n1588);
  and g2113 (n1590, n_872, n_805);
  not g2114 (n_949, n1589);
  not g2115 (n_950, n1590);
  and g2116 (n1591, n_949, n_950);
  not g2117 (n_951, n1591);
  and g2118 (n1592, n1246, n_951);
  and g2119 (po127, n_67, n1592);
  and g2120 (n1594, n_152, n_148);
  and g2121 (n1595, n_33, n_29);
  not g2122 (n_952, n1595);
  and g2123 (n1596, pi054, n_952);
  not g2124 (n_953, n1594);
  not g2125 (n_954, n1596);
  and g2126 (n1597, n_953, n_954);
  not g2127 (n_955, n1597);
  and g2128 (n1598, n_67, n_955);
  and g2129 (po128, n_156, n1598);
  and g2130 (n1600, n_693, pi140);
  and g2131 (n1601, n1583, n1600);
  and g2132 (n1602, n_760, n_805);
  not g2133 (n_956, n1601);
  not g2134 (n_957, n1602);
  and g2135 (n1603, n_956, n_957);
  not g2136 (n_958, n1603);
  and g2137 (n1604, n1246, n_958);
  and g2138 (po130, n_67, n1604);
  or g2146 (po132, n_607, pi129);
  and g2147 (n1613, n_152, pi118);
  and g2148 (n1614, pi054, n_163);
  and g2149 (n1615, n549, n1614);
  not g2150 (n_960, n1613);
  not g2151 (n_961, n1615);
  and g2152 (n1616, n_960, n_961);
  not g2153 (n_962, n1616);
  and g2154 (po133, n_67, n_962);
  not g2155 (n_963, n724);
  and g2156 (po134, n_67, n_963);
  not g2157 (n_964, pi120);
  and g2158 (n1619, n_258, n_964);
  and g2159 (n1620, n_156, n1619);
  not g2160 (n_965, n1620);
  and g2161 (n1621, n_67, n_965);
  not g2162 (n_966, pi111);
  and g2163 (po135, n_966, n1621);
  and g2164 (n1623, pi081, pi120);
  and g2165 (po136, n_67, n1623);
  or g2166 (po137, pi129, pi134);
  or g2167 (po138, pi129, pi135);
  and g2168 (po139, pi057, n_67);
  and g2169 (n1628, n_260, pi125);
  not g2170 (n_969, n1628);
  and g2171 (n1629, n_156, n_969);
  not g2172 (n_970, n1629);
  and g2173 (po140, n_67, n_970);
  not g2174 (n_972, pi126);
  and g2175 (n1631, n_972, pi132);
  and g2176 (po141, pi133, n1631);
  and g2177 (n_1110, n291, n_8);
  and g2178 (n_1111, n_9, n_17);
  and g2179 (n_1112, n295, n300);
  and g2180 (n_1113, n301, n302);
  and g2181 (n305, n_1110, n_1111, n_1112, n_1113);
  and g2182 (n_1115, n_1114, n_12);
  not g2183 (n_1114, n328);
  and g2184 (n333, n300, n301, n332, n_1115);
  and g2185 (n319, n_1116, n_1117, n_1118, n_4);
  not g2186 (n_1116, n314);
  not g2187 (n_1117, n315);
  not g2188 (n_1118, n317);
  and g2189 (n_1120, n_1119, n344);
  not g2190 (n_1119, n371);
  and g2191 (n375, n354, n356, n300, n_1120);
  and g2192 (n_1121, n300, n311);
  and g2193 (n_1122, n341, n344);
  and g2194 (n350, n_5, n347, n_1121, n_1122);
  and g2195 (n362, n_1123, n_1124, n_1125, n_9);
  not g2196 (n_1123, n357);
  not g2197 (n_1124, n358);
  not g2198 (n_1125, n360);
  and g2199 (n_1126, n380, n381);
  and g2200 (n_1127, n385, n389);
  and g2201 (n394, n_125, n391, n_1126, n_1127);
  and g2202 (n409, n398, n399, n401, n408);
  and g2203 (n_1128, n418, n341);
  and g2204 (n423, n419, n_13, n300, n_1128);
  and g2205 (n_1129, n369, n416);
  and g2206 (n435, pi010, n_29, n434, n_1129);
  and g2207 (n_1130, n_9, n332, pi028);
  and g2208 (n_1131, n_159, n_160, n445);
  and g2209 (n_1132, n447, n448);
  and g2210 (n_1133, n_28, n450);
  and g2211 (n454, n_1130, n_1131, n_1132, n_1133);
  and g2212 (n_1134, n445, n459, n_17);
  and g2213 (n_1135, n_167, pi025, n_160);
  and g2215 (n_1137, n_8, n450);
  and g2216 (n468, n_1134, n_1135, n_1132, n_1137);
  and g2217 (n_1138, n473, pi008, n_12);
  and g2218 (n_1139, n448, n_9);
  and g2219 (n_1140, n449, n445);
  and g2220 (n_1141, n_28, n479);
  and g2221 (n482, n_1138, n_1139, n_1140, n_1141);
  and g2222 (n_1142, n487, n488);
  and g2223 (n_1143, n_33, pi021);
  and g2224 (n_1144, n448, n_15);
  and g2225 (n494, n449, n_1142, n_1143, n_1144);
  and g2226 (n_1145, n291, n344, n332);
  and g2227 (n_1146, pi011, n459);
  and g2228 (n_1147, n503, n448);
  and g2229 (n_1148, n_32, n449);
  and g2230 (n507, n_1145, n_1146, n_1147, n_1148);
  and g2232 (n_1150, n_53, n449);
  and g2233 (n_1151, n515, n322);
  and g2234 (n_1152, n_32, n_29);
  and g2235 (n519, n_1147, n_1150, n_1151, n_1152);
  and g2237 (n_1154, n_33, n449);
  and g2239 (n_1156, n_53, pi022);
  and g2240 (n530, n_1147, n_1154, n_1129, n_1156);
  and g2241 (n_1157, n448, n_17);
  and g2242 (n_1158, n449, pi018);
  and g2243 (n_1159, n295, n_33);
  and g2244 (n540, n418, n_1157, n_1158, n_1159);
  and g2246 (n_1161, n_4, n450);
  and g2247 (n_1162, n357, n549);
  and g2248 (n_1163, n_9, n417);
  and g2249 (n553, n_1132, n_1161, n_1162, n_1163);
  and g2250 (n_1164, n503, n449);
  and g2251 (n_1165, n_25, n354);
  and g2252 (n_1166, n515, n344);
  and g2253 (n_1167, n_32, pi013);
  and g2254 (n564, n_1164, n_1165, n_1166, n_1167);
  and g2255 (n_1168, n399, n568);
  and g2256 (n575, n570, n_104, n573, n_1168);
  and g2257 (n_1170, n_1169, n583);
  not g2258 (n_1169, n584);
  and g2259 (n588, n384, n408, n_104, n_1170);
  and g2260 (n_1171, n434, n417);
  and g2261 (n_1172, n345, n_28);
  and g2262 (n600, pi006, n_17, n_1171, n_1172);
  and g2263 (n_1173, n445, n_9, n346);
  and g2264 (n_1174, n_17, n_159, n_167);
  and g2265 (n_1175, n450, n_25, n351);
  and g2266 (n_1176, n612, n_160, pi059);
  and g2267 (n616, n_1173, n_1174, n_1175, n_1176);
  and g2268 (n_1177, n487, n356);
  and g2269 (n624, n450, pi016, pi054, n_1177);
  and g2270 (n_1178, n487, pi017);
  and g2271 (n_1179, n612, n448);
  and g2273 (n634, n_20, n_1178, n_1179, n449);
  and g2274 (n645, n640, n642, n_121, n401);
  and g2275 (n653, n640, n649, n390, n650);
  and g2276 (n_1181, n487, n355);
  and g2277 (n_1182, n488, n299);
  and g2278 (n_1183, pi019, n_13);
  and g2279 (n668, pi054, n_1181, n_1182, n_1183);
  and g2280 (n_1184, n503, n448, n_29);
  and g2281 (n_1185, n449, n291, n_32);
  and g2282 (n_1186, n_53, n479);
  and g2283 (n_1187, pi005, n_9);
  and g2284 (n681, n_1184, n_1185, n_1186, n_1187);
  and g2285 (po039, n_1188, n_1189, n_1190, n_67);
  not g2286 (n_1188, n696);
  not g2287 (n_1189, n703);
  not g2288 (n_1190, n709);
  and g2289 (n_1191, n705, n649);
  and g2290 (n709, n390, pi024, pi082, n_1191);
  and g2291 (po041, n_1192, n_156, n_67, n774);
  not g2292 (n_1192, n770);
  and g2293 (po042, n_1193, n_156, n_67, n788);
  not g2294 (n_1193, n784);
  and g2295 (n802, n776, n_258, n_269, n_279);
  and g2296 (po053, n_1194, n_1195, n_1196, n_67);
  not g2297 (n_1194, n924);
  not g2298 (n_1195, n933);
  not g2299 (n_1196, n936);
  and g2300 (n930, n927, n638, n_117, n391);
  and g2301 (n927, n401, n398, n_125, n_97);
  and g2302 (po055, n_1197, n_1198, n_1199, n_67);
  not g2303 (n_1197, n953);
  not g2304 (n_1198, n959);
  not g2305 (n_1199, n961);
  and g2306 (n956, n927, n638, n388, n390);
  and g2307 (po056, n_1200, n_1201, n_1202, n_67);
  not g2308 (n_1200, n969);
  not g2309 (n_1201, n975);
  not g2310 (n_1202, n979);
  and g2311 (n979, n976, n390, pi041, pi082);
  and g2312 (n972, n927, n404, n381, n405);
  and g2313 (po057, n_1203, n_1204, n_1205, n_67);
  not g2314 (n_1203, n989);
  not g2315 (n_1204, n995);
  not g2316 (n_1205, n996);
  and g2317 (po058, n_1206, n_1207, n_1208, n_67);
  not g2318 (n_1206, n1005);
  not g2319 (n_1207, n1010);
  not g2320 (n_1208, n1013);
  and g2321 (n1013, n389, n934, pi043, n641);
  and g2322 (po060, n_1209, n_1210, n_1211, n_67);
  not g2323 (n_1209, n1034);
  not g2324 (n_1210, n1040);
  not g2325 (n_1211, n1044);
  and g2326 (n1044, n918, n934, pi045, n1041);
  and g2327 (po061, n_1212, n_1213, n_1214, n_67);
  not g2328 (n_1212, n1053);
  not g2329 (n_1213, n1058);
  not g2330 (n_1214, n1060);
  and g2331 (po062, n_1215, n_1216, n_1217, n_67);
  not g2332 (n_1215, n1068);
  not g2333 (n_1216, n1072);
  not g2334 (n_1217, n1076);
  and g2335 (n_1218, n568, n572);
  and g2336 (n1076, n934, pi047, n641, n_1218);
  and g2337 (po063, n_1219, n_1220, n_1221, n_67);
  not g2338 (n_1219, n1085);
  not g2339 (n_1220, n1092);
  not g2340 (n_1221, n1096);
  and g2341 (n_1222, n381, n406);
  and g2342 (n1096, n934, pi048, n1041, n_1222);
  and g2343 (n1089, n408, n_125, n_101, n1087);
  and g2344 (n1112, n_1223, n380, n638, n1100);
  not g2345 (n_1223, n1109);
  and g2346 (n1107, n705, n990, n_108, n_120);
  and g2347 (po065, n_1224, n_1225, n_1226, n_67);
  not g2348 (n_1224, n1125);
  not g2349 (n_1225, n1130);
  not g2350 (n_1226, n1132);
  and g2351 (n_1228, n_1227, n_269);
  not g2352 (n_1227, n1152);
  and g2353 (po068, n754, n_156, n_67, n_1228);
  and g2354 (n1147, n724, n_260, n_310, n_258);
  and g2355 (n_1230, n_1229, n_257);
  not g2356 (n_1229, n1209);
  and g2357 (po073, n_305, n_156, n_67, n_1230);
  and g2358 (n1208, n737, n_310, pi116, n_334);
  and g2359 (po076, n_1231, n_67, n_607, pi123);
  not g2360 (n_1231, pi114);
  and g2361 (n1247, pi136, n_670, n_671, n1246);
  and g2362 (n_1233, n_1232, n_269);
  not g2363 (n_1232, n1372);
  and g2364 (po100, n774, n_156, n_67, n_1233);
  and g2365 (po124, n_1234, pi116, n_156, n_67);
  not g2366 (n_1234, n1571);
  and g2367 (po125, n_1235, pi116, n_156, n_67);
  not g2368 (n_1235, n1576);
  and g2369 (po131, n_1236, pi054, n_156, n_67);
  not g2370 (n_1236, n1608);
  and g2371 (n1608, n_24, n_17, n_9, n_32);
endmodule

