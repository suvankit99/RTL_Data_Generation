
module max(\in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
     \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
     \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
     \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
     \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
     \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
     \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
     \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
     \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
     \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
     \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
     \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
     \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
     \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
     \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
     \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
     \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101]
     , \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] ,
     \in0[107] , \in0[108] , \in0[109] , \in0[110] , \in0[111] ,
     \in0[112] , \in0[113] , \in0[114] , \in0[115] , \in0[116] ,
     \in0[117] , \in0[118] , \in0[119] , \in0[120] , \in0[121] ,
     \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
     \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] ,
     \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
     \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
     \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
     \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
     \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
     \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
     \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
     \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
     \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
     \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
     \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
     \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
     \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
     \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
     \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
     \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
     \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] ,
     \in1[106] , \in1[107] , \in1[108] , \in1[109] , \in1[110] ,
     \in1[111] , \in1[112] , \in1[113] , \in1[114] , \in1[115] ,
     \in1[116] , \in1[117] , \in1[118] , \in1[119] , \in1[120] ,
     \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
     \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
     \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
     \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
     \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
     \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
     \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
     \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
     \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
     \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
     \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
     \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
     \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
     \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
     \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
     \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
     \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
     \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
     \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] ,
     \in2[105] , \in2[106] , \in2[107] , \in2[108] , \in2[109] ,
     \in2[110] , \in2[111] , \in2[112] , \in2[113] , \in2[114] ,
     \in2[115] , \in2[116] , \in2[117] , \in2[118] , \in2[119] ,
     \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
     \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
     \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
     \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
     \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
     \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
     \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
     \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
     \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
     \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
     \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
     \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
     \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
     \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
     \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
     \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
     \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
     \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
     \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] ,
     \in3[104] , \in3[105] , \in3[106] , \in3[107] , \in3[108] ,
     \in3[109] , \in3[110] , \in3[111] , \in3[112] , \in3[113] ,
     \in3[114] , \in3[115] , \in3[116] , \in3[117] , \in3[118] ,
     \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
     \in3[124] , \in3[125] , \in3[126] , \in3[127] , \result[0] ,
     \result[1] , \result[2] , \result[3] , \result[4] , \result[5] ,
     \result[6] , \result[7] , \result[8] , \result[9] , \result[10] ,
     \result[11] , \result[12] , \result[13] , \result[14] ,
     \result[15] , \result[16] , \result[17] , \result[18] ,
     \result[19] , \result[20] , \result[21] , \result[22] ,
     \result[23] , \result[24] , \result[25] , \result[26] ,
     \result[27] , \result[28] , \result[29] , \result[30] ,
     \result[31] , \result[32] , \result[33] , \result[34] ,
     \result[35] , \result[36] , \result[37] , \result[38] ,
     \result[39] , \result[40] , \result[41] , \result[42] ,
     \result[43] , \result[44] , \result[45] , \result[46] ,
     \result[47] , \result[48] , \result[49] , \result[50] ,
     \result[51] , \result[52] , \result[53] , \result[54] ,
     \result[55] , \result[56] , \result[57] , \result[58] ,
     \result[59] , \result[60] , \result[61] , \result[62] ,
     \result[63] , \result[64] , \result[65] , \result[66] ,
     \result[67] , \result[68] , \result[69] , \result[70] ,
     \result[71] , \result[72] , \result[73] , \result[74] ,
     \result[75] , \result[76] , \result[77] , \result[78] ,
     \result[79] , \result[80] , \result[81] , \result[82] ,
     \result[83] , \result[84] , \result[85] , \result[86] ,
     \result[87] , \result[88] , \result[89] , \result[90] ,
     \result[91] , \result[92] , \result[93] , \result[94] ,
     \result[95] , \result[96] , \result[97] , \result[98] ,
     \result[99] , \result[100] , \result[101] , \result[102] ,
     \result[103] , \result[104] , \result[105] , \result[106] ,
     \result[107] , \result[108] , \result[109] , \result[110] ,
     \result[111] , \result[112] , \result[113] , \result[114] ,
     \result[115] , \result[116] , \result[117] , \result[118] ,
     \result[119] , \result[120] , \result[121] , \result[122] ,
     \result[123] , \result[124] , \result[125] , \result[126] ,
     \result[127] , \address[0] , \address[1] );
//   input \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
       \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
       \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17]
       , \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] ,
       \in0[23] , \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28]
       , \in0[29] , \in0[30] , \in0[31] , \in0[32] , \in0[33] ,
       \in0[34] , \in0[35] , \in0[36] , \in0[37] , \in0[38] , \in0[39]
       , \in0[40] , \in0[41] , \in0[42] , \in0[43] , \in0[44] ,
       \in0[45] , \in0[46] , \in0[47] , \in0[48] , \in0[49] , \in0[50]
       , \in0[51] , \in0[52] , \in0[53] , \in0[54] , \in0[55] ,
       \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] , \in0[61]
       , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
       \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72]
       , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
       \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83]
       , \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] ,
       \in0[89] , \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94]
       , \in0[95] , \in0[96] , \in0[97] , \in0[98] , \in0[99] ,
       \in0[100] , \in0[101] , \in0[102] , \in0[103] , \in0[104] ,
       \in0[105] , \in0[106] , \in0[107] , \in0[108] , \in0[109] ,
       \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
       \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
       \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] ,
       \in0[125] , \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2]
       , \in1[3] , \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] ,
       \in1[9] , \in1[10] , \in1[11] , \in1[12] , \in1[13] , \in1[14] ,
       \in1[15] , \in1[16] , \in1[17] , \in1[18] , \in1[19] , \in1[20]
       , \in1[21] , \in1[22] , \in1[23] , \in1[24] , \in1[25] ,
       \in1[26] , \in1[27] , \in1[28] , \in1[29] , \in1[30] , \in1[31]
       , \in1[32] , \in1[33] , \in1[34] , \in1[35] , \in1[36] ,
       \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] , \in1[42]
       , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
       \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53]
       , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
       \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64]
       , \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] ,
       \in1[70] , \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75]
       , \in1[76] , \in1[77] , \in1[78] , \in1[79] , \in1[80] ,
       \in1[81] , \in1[82] , \in1[83] , \in1[84] , \in1[85] , \in1[86]
       , \in1[87] , \in1[88] , \in1[89] , \in1[90] , \in1[91] ,
       \in1[92] , \in1[93] , \in1[94] , \in1[95] , \in1[96] , \in1[97]
       , \in1[98] , \in1[99] , \in1[100] , \in1[101] , \in1[102] ,
       \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
       \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
       \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] ,
       \in1[118] , \in1[119] , \in1[120] , \in1[121] , \in1[122] ,
       \in1[123] , \in1[124] , \in1[125] , \in1[126] , \in1[127] ,
       \in2[0] , \in2[1] , \in2[2] , \in2[3] , \in2[4] , \in2[5] ,
       \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] , \in2[11] ,
       \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] , \in2[17]
       , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
       \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28]
       , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
       \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39]
       , \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] ,
       \in2[45] , \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50]
       , \in2[51] , \in2[52] , \in2[53] , \in2[54] , \in2[55] ,
       \in2[56] , \in2[57] , \in2[58] , \in2[59] , \in2[60] , \in2[61]
       , \in2[62] , \in2[63] , \in2[64] , \in2[65] , \in2[66] ,
       \in2[67] , \in2[68] , \in2[69] , \in2[70] , \in2[71] , \in2[72]
       , \in2[73] , \in2[74] , \in2[75] , \in2[76] , \in2[77] ,
       \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] , \in2[83]
       , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
       \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94]
       , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
       \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] ,
       \in2[105] , \in2[106] , \in2[107] , \in2[108] , \in2[109] ,
       \in2[110] , \in2[111] , \in2[112] , \in2[113] , \in2[114] ,
       \in2[115] , \in2[116] , \in2[117] , \in2[118] , \in2[119] ,
       \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
       \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2]
       , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
       \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
       \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20]
       , \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] ,
       \in3[26] , \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31]
       , \in3[32] , \in3[33] , \in3[34] , \in3[35] , \in3[36] ,
       \in3[37] , \in3[38] , \in3[39] , \in3[40] , \in3[41] , \in3[42]
       , \in3[43] , \in3[44] , \in3[45] , \in3[46] , \in3[47] ,
       \in3[48] , \in3[49] , \in3[50] , \in3[51] , \in3[52] , \in3[53]
       , \in3[54] , \in3[55] , \in3[56] , \in3[57] , \in3[58] ,
       \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] , \in3[64]
       , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
       \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75]
       , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
       \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86]
       , \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] ,
       \in3[92] , \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97]
       , \in3[98] , \in3[99] , \in3[100] , \in3[101] , \in3[102] ,
       \in3[103] , \in3[104] , \in3[105] , \in3[106] , \in3[107] ,
       \in3[108] , \in3[109] , \in3[110] , \in3[111] , \in3[112] ,
       \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
       \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
       \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
//   output \result[0] , \result[1] , \result[2] , \result[3] , \result[4]
       , \result[5] , \result[6] , \result[7] , \result[8] , \result[9]
       , \result[10] , \result[11] , \result[12] , \result[13] ,
       \result[14] , \result[15] , \result[16] , \result[17] ,
       \result[18] , \result[19] , \result[20] , \result[21] ,
       \result[22] , \result[23] , \result[24] , \result[25] ,
       \result[26] , \result[27] , \result[28] , \result[29] ,
       \result[30] , \result[31] , \result[32] , \result[33] ,
       \result[34] , \result[35] , \result[36] , \result[37] ,
       \result[38] , \result[39] , \result[40] , \result[41] ,
       \result[42] , \result[43] , \result[44] , \result[45] ,
       \result[46] , \result[47] , \result[48] , \result[49] ,
       \result[50] , \result[51] , \result[52] , \result[53] ,
       \result[54] , \result[55] , \result[56] , \result[57] ,
       \result[58] , \result[59] , \result[60] , \result[61] ,
       \result[62] , \result[63] , \result[64] , \result[65] ,
       \result[66] , \result[67] , \result[68] , \result[69] ,
       \result[70] , \result[71] , \result[72] , \result[73] ,
       \result[74] , \result[75] , \result[76] , \result[77] ,
       \result[78] , \result[79] , \result[80] , \result[81] ,
       \result[82] , \result[83] , \result[84] , \result[85] ,
       \result[86] , \result[87] , \result[88] , \result[89] ,
       \result[90] , \result[91] , \result[92] , \result[93] ,
       \result[94] , \result[95] , \result[96] , \result[97] ,
       \result[98] , \result[99] , \result[100] , \result[101] ,
       \result[102] , \result[103] , \result[104] , \result[105] ,
       \result[106] , \result[107] , \result[108] , \result[109] ,
       \result[110] , \result[111] , \result[112] , \result[113] ,
       \result[114] , \result[115] , \result[116] , \result[117] ,
       \result[118] , \result[119] , \result[120] , \result[121] ,
       \result[122] , \result[123] , \result[124] , \result[125] ,
       \result[126] , \result[127] , \address[0] , \address[1] ;
  wire \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
       \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
       \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17]
       , \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] ,
       \in0[23] , \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28]
       , \in0[29] , \in0[30] , \in0[31] , \in0[32] , \in0[33] ,
       \in0[34] , \in0[35] , \in0[36] , \in0[37] , \in0[38] , \in0[39]
       , \in0[40] , \in0[41] , \in0[42] , \in0[43] , \in0[44] ,
       \in0[45] , \in0[46] , \in0[47] , \in0[48] , \in0[49] , \in0[50]
       , \in0[51] , \in0[52] , \in0[53] , \in0[54] , \in0[55] ,
       \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] , \in0[61]
       , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
       \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72]
       , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
       \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83]
       , \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] ,
       \in0[89] , \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94]
       , \in0[95] , \in0[96] , \in0[97] , \in0[98] , \in0[99] ,
       \in0[100] , \in0[101] , \in0[102] , \in0[103] , \in0[104] ,
       \in0[105] , \in0[106] , \in0[107] , \in0[108] , \in0[109] ,
       \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
       \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
       \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] ,
       \in0[125] , \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2]
       , \in1[3] , \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] ,
       \in1[9] , \in1[10] , \in1[11] , \in1[12] , \in1[13] , \in1[14] ,
       \in1[15] , \in1[16] , \in1[17] , \in1[18] , \in1[19] , \in1[20]
       , \in1[21] , \in1[22] , \in1[23] , \in1[24] , \in1[25] ,
       \in1[26] , \in1[27] , \in1[28] , \in1[29] , \in1[30] , \in1[31]
       , \in1[32] , \in1[33] , \in1[34] , \in1[35] , \in1[36] ,
       \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] , \in1[42]
       , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
       \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53]
       , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
       \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64]
       , \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] ,
       \in1[70] , \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75]
       , \in1[76] , \in1[77] , \in1[78] , \in1[79] , \in1[80] ,
       \in1[81] , \in1[82] , \in1[83] , \in1[84] , \in1[85] , \in1[86]
       , \in1[87] , \in1[88] , \in1[89] , \in1[90] , \in1[91] ,
       \in1[92] , \in1[93] , \in1[94] , \in1[95] , \in1[96] , \in1[97]
       , \in1[98] , \in1[99] , \in1[100] , \in1[101] , \in1[102] ,
       \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
       \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
       \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] ,
       \in1[118] , \in1[119] , \in1[120] , \in1[121] , \in1[122] ,
       \in1[123] , \in1[124] , \in1[125] , \in1[126] , \in1[127] ,
       \in2[0] , \in2[1] , \in2[2] , \in2[3] , \in2[4] , \in2[5] ,
       \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] , \in2[11] ,
       \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] , \in2[17]
       , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
       \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28]
       , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
       \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39]
       , \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] ,
       \in2[45] , \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50]
       , \in2[51] , \in2[52] , \in2[53] , \in2[54] , \in2[55] ,
       \in2[56] , \in2[57] , \in2[58] , \in2[59] , \in2[60] , \in2[61]
       , \in2[62] , \in2[63] , \in2[64] , \in2[65] , \in2[66] ,
       \in2[67] , \in2[68] , \in2[69] , \in2[70] , \in2[71] , \in2[72]
       , \in2[73] , \in2[74] , \in2[75] , \in2[76] , \in2[77] ,
       \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] , \in2[83]
       , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
       \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94]
       , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
       \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] ,
       \in2[105] , \in2[106] , \in2[107] , \in2[108] , \in2[109] ,
       \in2[110] , \in2[111] , \in2[112] , \in2[113] , \in2[114] ,
       \in2[115] , \in2[116] , \in2[117] , \in2[118] , \in2[119] ,
       \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
       \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2]
       , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
       \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
       \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20]
       , \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] ,
       \in3[26] , \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31]
       , \in3[32] , \in3[33] , \in3[34] , \in3[35] , \in3[36] ,
       \in3[37] , \in3[38] , \in3[39] , \in3[40] , \in3[41] , \in3[42]
       , \in3[43] , \in3[44] , \in3[45] , \in3[46] , \in3[47] ,
       \in3[48] , \in3[49] , \in3[50] , \in3[51] , \in3[52] , \in3[53]
       , \in3[54] , \in3[55] , \in3[56] , \in3[57] , \in3[58] ,
       \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] , \in3[64]
       , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
       \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75]
       , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
       \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86]
       , \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] ,
       \in3[92] , \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97]
       , \in3[98] , \in3[99] , \in3[100] , \in3[101] , \in3[102] ,
       \in3[103] , \in3[104] , \in3[105] , \in3[106] , \in3[107] ,
       \in3[108] , \in3[109] , \in3[110] , \in3[111] , \in3[112] ,
       \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
       \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
       \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  wire \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
       \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
       \result[10] , \result[11] , \result[12] , \result[13] ,
       \result[14] , \result[15] , \result[16] , \result[17] ,
       \result[18] , \result[19] , \result[20] , \result[21] ,
       \result[22] , \result[23] , \result[24] , \result[25] ,
       \result[26] , \result[27] , \result[28] , \result[29] ,
       \result[30] , \result[31] , \result[32] , \result[33] ,
       \result[34] , \result[35] , \result[36] , \result[37] ,
       \result[38] , \result[39] , \result[40] , \result[41] ,
       \result[42] , \result[43] , \result[44] , \result[45] ,
       \result[46] , \result[47] , \result[48] , \result[49] ,
       \result[50] , \result[51] , \result[52] , \result[53] ,
       \result[54] , \result[55] , \result[56] , \result[57] ,
       \result[58] , \result[59] , \result[60] , \result[61] ,
       \result[62] , \result[63] , \result[64] , \result[65] ,
       \result[66] , \result[67] , \result[68] , \result[69] ,
       \result[70] , \result[71] , \result[72] , \result[73] ,
       \result[74] , \result[75] , \result[76] , \result[77] ,
       \result[78] , \result[79] , \result[80] , \result[81] ,
       \result[82] , \result[83] , \result[84] , \result[85] ,
       \result[86] , \result[87] , \result[88] , \result[89] ,
       \result[90] , \result[91] , \result[92] , \result[93] ,
       \result[94] , \result[95] , \result[96] , \result[97] ,
       \result[98] , \result[99] , \result[100] , \result[101] ,
       \result[102] , \result[103] , \result[104] , \result[105] ,
       \result[106] , \result[107] , \result[108] , \result[109] ,
       \result[110] , \result[111] , \result[112] , \result[113] ,
       \result[114] , \result[115] , \result[116] , \result[117] ,
       \result[118] , \result[119] , \result[120] , \result[121] ,
       \result[122] , \result[123] , \result[124] , \result[125] ,
       \result[126] , \result[127] , \address[0] , \address[1] ;
  wire n643, n644, n645, n646, n647, n648, n649, n650;
  wire n651, n652, n653, n654, n655, n656, n657, n658;
  wire n659, n660, n661, n662, n663, n664, n665, n666;
  wire n667, n668, n669, n670, n671, n672, n673, n674;
  wire n675, n676, n677, n678, n679, n680, n681, n682;
  wire n683, n684, n685, n686, n687, n688, n689, n690;
  wire n691, n692, n693, n694, n695, n696, n697, n698;
  wire n699, n700, n701, n702, n703, n704, n705, n706;
  wire n707, n708, n709, n710, n711, n712, n713, n714;
  wire n715, n716, n717, n718, n719, n720, n721, n722;
  wire n723, n724, n725, n726, n727, n728, n729, n730;
  wire n731, n732, n733, n734, n735, n736, n737, n738;
  wire n739, n740, n741, n742, n743, n744, n745, n746;
  wire n747, n748, n749, n750, n751, n752, n753, n754;
  wire n755, n756, n757, n758, n759, n760, n761, n762;
  wire n763, n764, n765, n766, n767, n768, n769, n770;
  wire n771, n772, n773, n774, n775, n776, n777, n778;
  wire n779, n780, n781, n782, n783, n784, n785, n786;
  wire n787, n788, n789, n790, n791, n792, n793, n794;
  wire n795, n796, n797, n798, n799, n800, n801, n802;
  wire n803, n804, n805, n806, n807, n808, n809, n810;
  wire n811, n812, n813, n814, n815, n816, n817, n818;
  wire n819, n820, n821, n822, n823, n824, n825, n826;
  wire n827, n828, n829, n830, n831, n832, n833, n834;
  wire n835, n836, n837, n838, n839, n840, n841, n842;
  wire n843, n844, n845, n846, n847, n848, n849, n850;
  wire n851, n852, n853, n854, n855, n856, n857, n858;
  wire n859, n860, n861, n862, n863, n864, n865, n866;
  wire n867, n868, n869, n870, n871, n872, n873, n874;
  wire n875, n876, n877, n878, n879, n880, n881, n882;
  wire n883, n884, n885, n886, n887, n888, n889, n890;
  wire n891, n892, n893, n894, n895, n896, n897, n898;
  wire n899, n900, n901, n902, n903, n904, n905, n906;
  wire n907, n908, n909, n910, n911, n912, n913, n914;
  wire n915, n916, n917, n918, n919, n920, n921, n922;
  wire n923, n924, n925, n926, n927, n928, n929, n930;
  wire n931, n932, n933, n934, n935, n936, n937, n938;
  wire n939, n940, n944, n945, n946, n947, n948, n949;
  wire n950, n951, n952, n953, n954, n955, n956, n957;
  wire n958, n959, n960, n961, n962, n966, n967, n971;
  wire n975, n976, n977, n978, n979, n980, n981, n982;
  wire n983, n984, n985, n986, n987, n991, n992, n993;
  wire n994, n995, n996, n997, n998, n999, n1000, n1001;
  wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009;
  wire n1012, n1013, n1017, n1021, n1022, n1025, n1026, n1027;
  wire n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  wire n1036, n1039, n1042, n1043, n1044, n1045, n1046, n1047;
  wire n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057;
  wire n1058, n1059, n1060, n1061, n1064, n1067, n1070, n1071;
  wire n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079;
  wire n1080, n1081, n1084, n1087, n1088, n1089, n1090, n1091;
  wire n1092, n1095, n1096, n1097, n1098, n1099, n1100, n1101;
  wire n1102, n1103, n1104, n1105, n1106, n1109, n1112, n1115;
  wire n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123;
  wire n1124, n1125, n1126, n1129, n1132, n1133, n1134, n1135;
  wire n1136, n1137, n1140, n1141, n1142, n1143, n1144, n1145;
  wire n1146, n1147, n1148, n1149, n1150, n1151, n1154, n1157;
  wire n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167;
  wire n1168, n1169, n1170, n1171, n1174, n1177, n1178, n1179;
  wire n1180, n1181, n1182, n1185, n1186, n1187, n1188, n1189;
  wire n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197;
  wire n1198, n1199, n1200, n1203, n1204, n1205, n1206, n1207;
  wire n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215;
  wire n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223;
  wire n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231;
  wire n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239;
  wire n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247;
  wire n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255;
  wire n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263;
  wire n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271;
  wire n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279;
  wire n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287;
  wire n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295;
  wire n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303;
  wire n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311;
  wire n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319;
  wire n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327;
  wire n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335;
  wire n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343;
  wire n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351;
  wire n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359;
  wire n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367;
  wire n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;
  wire n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383;
  wire n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391;
  wire n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399;
  wire n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407;
  wire n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415;
  wire n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423;
  wire n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431;
  wire n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439;
  wire n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447;
  wire n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455;
  wire n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463;
  wire n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471;
  wire n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479;
  wire n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487;
  wire n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495;
  wire n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503;
  wire n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511;
  wire n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522;
  wire n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530;
  wire n1531, n1532, n1533, n1537, n1538, n1542, n1546, n1547;
  wire n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555;
  wire n1556, n1557, n1558, n1562, n1563, n1564, n1565, n1566;
  wire n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574;
  wire n1575, n1576, n1577, n1578, n1579, n1580, n1583, n1584;
  wire n1588, n1592, n1593, n1596, n1597, n1598, n1599, n1600;
  wire n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1610;
  wire n1613, n1614, n1615, n1616, n1617, n1618, n1621, n1622;
  wire n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630;
  wire n1631, n1632, n1635, n1638, n1641, n1642, n1643, n1644;
  wire n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652;
  wire n1655, n1658, n1659, n1660, n1661, n1662, n1663, n1666;
  wire n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674;
  wire n1675, n1676, n1677, n1680, n1683, n1686, n1687, n1688;
  wire n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696;
  wire n1697, n1700, n1703, n1704, n1705, n1706, n1707, n1708;
  wire n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718;
  wire n1719, n1720, n1721, n1722, n1725, n1728, n1731, n1732;
  wire n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740;
  wire n1741, n1742, n1745, n1748, n1749, n1750, n1751, n1752;
  wire n1753, n1756, n1757, n1758, n1759, n1760, n1761, n1762;
  wire n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770;
  wire n1771, n1774, n1775, n1776, n1777, n1778, n1779, n1780;
  wire n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788;
  wire n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796;
  wire n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804;
  wire n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812;
  wire n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820;
  wire n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828;
  wire n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836;
  wire n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844;
  wire n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852;
  wire n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860;
  wire n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868;
  wire n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876;
  wire n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884;
  wire n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892;
  wire n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900;
  wire n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908;
  wire n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916;
  wire n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924;
  wire n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932;
  wire n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940;
  wire n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948;
  wire n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956;
  wire n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964;
  wire n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972;
  wire n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980;
  wire n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988;
  wire n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996;
  wire n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004;
  wire n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012;
  wire n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020;
  wire n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;
  wire n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036;
  wire n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044;
  wire n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052;
  wire n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060;
  wire n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068;
  wire n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076;
  wire n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084;
  wire n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092;
  wire n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100;
  wire n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108;
  wire n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116;
  wire n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124;
  wire n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132;
  wire n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140;
  wire n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148;
  wire n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156;
  wire n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164;
  wire n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172;
  wire n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180;
  wire n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188;
  wire n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196;
  wire n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204;
  wire n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212;
  wire n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220;
  wire n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228;
  wire n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236;
  wire n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244;
  wire n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252;
  wire n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260;
  wire n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268;
  wire n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276;
  wire n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284;
  wire n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292;
  wire n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300;
  wire n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308;
  wire n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316;
  wire n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324;
  wire n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332;
  wire n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340;
  wire n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348;
  wire n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356;
  wire n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364;
  wire n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372;
  wire n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380;
  wire n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388;
  wire n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396;
  wire n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404;
  wire n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412;
  wire n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420;
  wire n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428;
  wire n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436;
  wire n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444;
  wire n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452;
  wire n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460;
  wire n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468;
  wire n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476;
  wire n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484;
  wire n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492;
  wire n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500;
  wire n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508;
  wire n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516;
  wire n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524;
  wire n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532;
  wire n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540;
  wire n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548;
  wire n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556;
  wire n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564;
  wire n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572;
  wire n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580;
  wire n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588;
  wire n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596;
  wire n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604;
  wire n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612;
  wire n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620;
  wire n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628;
  wire n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636;
  wire n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644;
  wire n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652;
  wire n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660;
  wire n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668;
  wire n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676;
  wire n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684;
  wire n2685, n2686, n2687, n2688, n2689, n2692, n2693, n2694;
  wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702;
  wire n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710;
  wire n2714, n2715, n2719, n2723, n2724, n2725, n2726, n2727;
  wire n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735;
  wire n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743;
  wire n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751;
  wire n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759;
  wire n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767;
  wire n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775;
  wire n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783;
  wire n2784, n2787, n2788, n2789, n2790, n2791, n2792, n2793;
  wire n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801;
  wire n2802, n2803, n2804, n2805, n2808, n2809, n2813, n2817;
  wire n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827;
  wire n2828, n2829, n2830, n2831, n2834, n2837, n2838, n2839;
  wire n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847;
  wire n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855;
  wire n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863;
  wire n2864, n2865, n2866, n2869, n2870, n2871, n2872, n2873;
  wire n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2883;
  wire n2886, n2889, n2890, n2891, n2892, n2893, n2894, n2895;
  wire n2896, n2897, n2898, n2899, n2900, n2903, n2906, n2907;
  wire n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915;
  wire n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923;
  wire n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931;
  wire n2932, n2933, n2934, n2935, n2938, n2939, n2940, n2941;
  wire n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949;
  wire n2952, n2955, n2958, n2959, n2960, n2961, n2962, n2963;
  wire n2964, n2965, n2966, n2967, n2968, n2969, n2972, n2975;
  wire n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983;
  wire n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991;
  wire n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999;
  wire n3000, n3001, n3002, n3003, n3004, n3007, n3008, n3009;
  wire n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017;
  wire n3018, n3021, n3024, n3027, n3028, n3029, n3030, n3031;
  wire n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3041;
  wire n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051;
  wire n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059;
  wire n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067;
  wire n3068, n3069, n3070, n3071, n3072, n3073, n3076, n3077;
  wire n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085;
  wire n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093;
  wire n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101;
  wire n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109;
  wire n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119;
  wire n3120, n3122, n3123, n3125, n3126, n3128, n3129, n3131;
  wire n3132, n3134, n3135, n3137, n3138, n3140, n3141, n3143;
  wire n3144, n3146, n3147, n3149, n3150, n3152, n3153, n3155;
  wire n3156, n3158, n3159, n3161, n3162, n3164, n3165, n3167;
  wire n3168, n3170, n3171, n3173, n3174, n3176, n3177, n3179;
  wire n3180, n3182, n3183, n3185, n3186, n3188, n3189, n3191;
  wire n3192, n3194, n3195, n3197, n3198, n3200, n3201, n3203;
  wire n3204, n3206, n3207, n3209, n3210, n3212, n3213, n3215;
  wire n3216, n3218, n3219, n3221, n3222, n3224, n3225, n3227;
  wire n3228, n3230, n3231, n3233, n3234, n3236, n3237, n3239;
  wire n3240, n3242, n3243, n3245, n3246, n3248, n3249, n3251;
  wire n3252, n3254, n3255, n3257, n3258, n3260, n3261, n3263;
  wire n3264, n3266, n3267, n3269, n3270, n3272, n3273, n3275;
  wire n3276, n3278, n3279, n3281, n3282, n3284, n3285, n3287;
  wire n3288, n3290, n3291, n3293, n3294, n3296, n3297, n3299;
  wire n3300, n3302, n3303, n3305, n3306, n3308, n3309, n3311;
  wire n3312, n3314, n3315, n3317, n3318, n3320, n3321, n3323;
  wire n3324, n3326, n3327, n3329, n3330, n3332, n3333, n3335;
  wire n3336, n3338, n3339, n3341, n3342, n3344, n3345, n3347;
  wire n3348, n3350, n3351, n3353, n3354, n3356, n3357, n3359;
  wire n3360, n3362, n3363, n3365, n3366, n3368, n3369, n3371;
  wire n3372, n3374, n3375, n3377, n3378, n3380, n3381, n3383;
  wire n3384, n3386, n3387, n3389, n3390, n3392, n3393, n3395;
  wire n3396, n3398, n3399, n3401, n3402, n3404, n3405, n3407;
  wire n3408, n3410, n3411, n3413, n3414, n3416, n3417, n3419;
  wire n3420, n3422, n3423, n3425, n3426, n3428, n3429, n3431;
  wire n3432, n3434, n3435, n3437, n3438, n3440, n3441, n3443;
  wire n3444, n3446, n3447, n3449, n3450, n3452, n3453, n3455;
  wire n3456, n3458, n3459, n3461, n3462, n3464, n3465, n3467;
  wire n3468, n3470, n3471, n3473, n3474, n3476, n3477, n3479;
  wire n3480, n3482, n3483, n3485, n3486, n3488, n3489, n3491;
  wire n3492, n3494, n3495, n3497, n3498, n3500, n3501, n3503;
  wire n3505, n3506, n_3, n_4, n_6, n_8, n_9, n_11;
  wire n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_23;
  wire n_26, n_29, n_31, n_32, n_34, n_38, n_39, n_41;
  wire n_43, n_44, n_46, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_59, n_60, n_62, n_64, n_65, n_67;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_79;
  wire n_82, n_85, n_87, n_88, n_90, n_94, n_95, n_97;
  wire n_99, n_100, n_102, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_115, n_116, n_118, n_120, n_121, n_123;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_135;
  wire n_138, n_141, n_143, n_144, n_146, n_150, n_151, n_153;
  wire n_155, n_156, n_158, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_171, n_172, n_174, n_176, n_177, n_179;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_191;
  wire n_194, n_196, n_197, n_199, n_203, n_204, n_206, n_208;
  wire n_209, n_211, n_214, n_216, n_217, n_220, n_221, n_223;
  wire n_225, n_226, n_228, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_251, n_252, n_254, n_256;
  wire n_257, n_259, n_262, n_264, n_265, n_268, n_269, n_271;
  wire n_273, n_274, n_276, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_298, n_301, n_304, n_307;
  wire n_310, n_313, n_316, n_319, n_322, n_325, n_328, n_331;
  wire n_334, n_337, n_340, n_343, n_346, n_349, n_352, n_355;
  wire n_358, n_361, n_365, n_368, n_370, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_386, n_388, n_389, n_390, n_391, n_392;
  wire n_394, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_412, n_414, n_415, n_416, n_417, n_418, n_420, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_458, n_460, n_461, n_462, n_463, n_464;
  wire n_466, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_504, n_506, n_507, n_508;
  wire n_509, n_510, n_512, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_550, n_553;
  wire n_555, n_556, n_558, n_561, n_563, n_564, n_566, n_569;
  wire n_572, n_574, n_575, n_576, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_602, n_611;
  wire n_614, n_617, n_619, n_620, n_622, n_625, n_627, n_628;
  wire n_630, n_633, n_636, n_638, n_639, n_640, n_643, n_644;
  wire n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
  wire n_661, n_666, n_675, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_699, n_702, n_704, n_705, n_707, n_710, n_712, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_733, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_755, n_758, n_760, n_761, n_763, n_766, n_768, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_789, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_811, n_814, n_816, n_817, n_819, n_822, n_824, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835;
  wire n_836, n_837, n_838, n_845, n_848, n_849, n_850, n_851;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_867, n_870, n_872, n_873, n_875, n_878, n_880, n_883;
  wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
  wire n_892, n_893, n_895, n_899, n_901, n_904, n_906, n_907;
  wire n_908, n_911, n_912, n_913, n_914, n_915, n_916, n_917;
  wire n_918, n_919, n_920, n_921, n_922, n_925, n_926, n_928;
  wire n_930, n_931, n_933, n_937, n_938, n_939, n_940, n_941;
  wire n_942, n_943, n_945, n_948, n_951, n_953, n_954, n_956;
  wire n_960, n_961, n_963, n_965, n_966, n_968, n_972, n_973;
  wire n_974, n_975, n_976, n_977, n_978, n_981, n_982, n_984;
  wire n_986, n_987, n_989, n_993, n_994, n_995, n_996, n_997;
  wire n_998, n_999, n_1001, n_1004, n_1007, n_1009, n_1010, n_1012;
  wire n_1016, n_1017, n_1019, n_1021, n_1022, n_1024, n_1028, n_1029;
  wire n_1030, n_1031, n_1032, n_1033, n_1034, n_1037, n_1038, n_1040;
  wire n_1042, n_1043, n_1045, n_1049, n_1050, n_1051, n_1052, n_1053;
  wire n_1054, n_1055, n_1057, n_1060, n_1063, n_1065, n_1066, n_1068;
  wire n_1072, n_1073, n_1075, n_1077, n_1078, n_1080, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1093, n_1094, n_1096;
  wire n_1098, n_1099, n_1101, n_1105, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1113, n_1116, n_1118, n_1119, n_1121, n_1125;
  wire n_1126, n_1128, n_1130, n_1131, n_1133, n_1136, n_1138, n_1139;
  wire n_1142, n_1143, n_1145, n_1147, n_1148, n_1150, n_1154, n_1155;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1173;
  wire n_1174, n_1176, n_1178, n_1179, n_1181, n_1184, n_1186, n_1187;
  wire n_1190, n_1191, n_1193, n_1195, n_1196, n_1198, n_1202, n_1203;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1220;
  wire n_1223, n_1226, n_1229, n_1232, n_1235, n_1238, n_1241, n_1244;
  wire n_1247, n_1250, n_1253, n_1256, n_1259, n_1262, n_1265, n_1268;
  wire n_1271, n_1274, n_1277, n_1280, n_1283, n_1287, n_1290, n_1291;
  wire n_1292, n_1294, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1309, n_1311;
  wire n_1312, n_1313, n_1314, n_1315, n_1317, n_1319, n_1320, n_1321;
  wire n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329;
  wire n_1330, n_1331, n_1332, n_1333, n_1335, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1343, n_1345, n_1346, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1381, n_1383;
  wire n_1384, n_1385, n_1386, n_1387, n_1389, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409;
  wire n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425;
  wire n_1427, n_1429, n_1430, n_1431, n_1432, n_1433, n_1435, n_1437;
  wire n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469;
  wire n_1470, n_1471, n_1473, n_1476, n_1478, n_1479, n_1481, n_1484;
  wire n_1486, n_1487, n_1489, n_1492, n_1495, n_1497, n_1498, n_1499;
  wire n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509;
  wire n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1525, n_1534, n_1537, n_1540, n_1542, n_1543;
  wire n_1545, n_1548, n_1550, n_1551, n_1553, n_1556, n_1559, n_1561;
  wire n_1562, n_1563, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571;
  wire n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579;
  wire n_1580, n_1581, n_1582, n_1583, n_1584, n_1589, n_1598, n_1602;
  wire n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610;
  wire n_1611, n_1612, n_1613, n_1614, n_1622, n_1625, n_1627, n_1628;
  wire n_1630, n_1633, n_1635, n_1638, n_1639, n_1640, n_1641, n_1642;
  wire n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1656;
  wire n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666;
  wire n_1667, n_1668, n_1669, n_1670, n_1678, n_1681, n_1683, n_1684;
  wire n_1686, n_1689, n_1691, n_1694, n_1695, n_1696, n_1697, n_1698;
  wire n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1712;
  wire n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722;
  wire n_1723, n_1724, n_1725, n_1726, n_1734, n_1737, n_1739, n_1740;
  wire n_1742, n_1745, n_1747, n_1750, n_1751, n_1752, n_1753, n_1754;
  wire n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1768;
  wire n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778;
  wire n_1779, n_1780, n_1781, n_1782, n_1790, n_1793, n_1795, n_1796;
  wire n_1798, n_1801, n_1803, n_1806, n_1807, n_1808, n_1809, n_1810;
  wire n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1818, n_1822;
  wire n_1824, n_1827, n_1829, n_1830, n_1831, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844;
  wire n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852;
  wire n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860;
  wire n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868;
  wire n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884;
  wire n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892;
  wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
  wire n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916;
  wire n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924;
  wire n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932;
  wire n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940;
  wire n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948;
  wire n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956;
  wire n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964;
  wire n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972;
  wire n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980;
  wire n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988;
  wire n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996;
  wire n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004;
  wire n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012;
  wire n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020;
  wire n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028;
  wire n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036;
  wire n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
  wire n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052;
  wire n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060;
  wire n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068;
  wire n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076;
  wire n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092;
  wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100;
  wire n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108;
  wire n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116;
  wire n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124;
  wire n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132;
  wire n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140;
  wire n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148;
  wire n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156;
  wire n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164;
  wire n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172;
  wire n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180;
  wire n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188;
  wire n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196;
  wire n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204;
  wire n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212;
  wire n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220;
  wire n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228;
  wire n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236;
  wire n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244;
  wire n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252;
  wire n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260;
  wire n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268;
  wire n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276;
  wire n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284;
  wire n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292;
  wire n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300;
  wire n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308;
  wire n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316;
  wire n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324;
  wire n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332;
  wire n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356;
  wire n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364;
  wire n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372;
  wire n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380;
  wire n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388;
  wire n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396;
  wire n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404;
  wire n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412;
  wire n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420;
  wire n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428;
  wire n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436;
  wire n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468;
  wire n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476;
  wire n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484;
  wire n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492;
  wire n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500;
  wire n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508;
  wire n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516;
  wire n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524;
  wire n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532;
  wire n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540;
  wire n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548;
  wire n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556;
  wire n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564;
  wire n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572;
  wire n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580;
  wire n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, n_2588;
  wire n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596;
  wire n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604;
  wire n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612;
  wire n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620;
  wire n_2621, n_2622, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630;
  wire n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638;
  wire n_2639, n_2640, n_2641, n_2642, n_2648, n_2656, n_2657, n_2658;
  wire n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666;
  wire n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674;
  wire n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682;
  wire n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690;
  wire n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698;
  wire n_2699, n_2700, n_2701, n_2702, n_2705, n_2706, n_2707, n_2708;
  wire n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716;
  wire n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2728;
  wire n_2736, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745;
  wire n_2746, n_2747, n_2748, n_2749, n_2750, n_2757, n_2758, n_2759;
  wire n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767;
  wire n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775;
  wire n_2776, n_2777, n_2778, n_2779, n_2782, n_2783, n_2784, n_2785;
  wire n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793;
  wire n_2800, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809;
  wire n_2810, n_2811, n_2812, n_2813, n_2814, n_2821, n_2822, n_2823;
  wire n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831;
  wire n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839;
  wire n_2840, n_2841, n_2842, n_2843, n_2846, n_2847, n_2848, n_2849;
  wire n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857;
  wire n_2864, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873;
  wire n_2874, n_2875, n_2876, n_2877, n_2878, n_2885, n_2886, n_2887;
  wire n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895;
  wire n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903;
  wire n_2904, n_2905, n_2906, n_2907, n_2910, n_2911, n_2912, n_2913;
  wire n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, n_2921;
  wire n_2928, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937;
  wire n_2938, n_2939, n_2940, n_2941, n_2942, n_2949, n_2950, n_2951;
  wire n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959;
  wire n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967;
  wire n_2968, n_2969, n_2970, n_2971, n_2974, n_2975, n_2976, n_2977;
  wire n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985;
  wire n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993;
  wire n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001;
  wire n_3002, n_3003, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011;
  wire n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3020;
  wire n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028;
  wire n_3029, n_3030, n_3031, n_3161, n_3162, n_3163, n_3164, n_3165;
  wire n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173;
  wire n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181;
  wire n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189;
  wire n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197;
  wire n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205;
  wire n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213;
  wire n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221;
  wire n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229;
  wire n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237;
  wire n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, n_3245;
  wire n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253;
  wire n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261;
  wire n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269;
  wire n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276, n_3277;
  wire n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, n_3285;
  wire n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293;
  wire n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301;
  wire n_3302, n_3303, n_3304, n_3305, n_3306;
  not g1 (n_3, \in3[119] );
  and g2 (n643, \in2[119] , n_3);
  not g3 (n_4, \in2[119] );
  and g4 (n644, n_4, \in3[119] );
  not g5 (n_6, \in2[118] );
  and g6 (n645, n_6, \in3[118] );
  not g7 (n_8, n644);
  not g8 (n_9, n645);
  and g9 (n646, n_8, n_9);
  not g10 (n_11, \in2[117] );
  and g11 (n647, n_11, \in3[117] );
  not g12 (n_15, \in3[116] );
  and g13 (n648, \in2[116] , n_15);
  not g14 (n_16, n647);
  and g15 (n649, n_16, n648);
  not g16 (n_17, \in3[117] );
  and g17 (n650, \in2[117] , n_17);
  not g18 (n_18, n649);
  not g19 (n_19, n650);
  and g20 (n651, n_18, n_19);
  not g21 (n_20, n651);
  and g22 (n652, n646, n_20);
  not g23 (n_21, \in3[118] );
  and g24 (n653, n_21, n_8);
  and g25 (n654, \in2[118] , n653);
  not g26 (n_23, \in2[112] );
  and g27 (n655, n_23, \in3[112] );
  not g28 (n_26, \in2[115] );
  and g29 (n656, n_26, \in3[115] );
  not g30 (n_29, \in2[114] );
  and g31 (n657, n_29, \in3[114] );
  not g32 (n_31, n656);
  not g33 (n_32, n657);
  and g34 (n658, n_31, n_32);
  not g35 (n_34, \in2[113] );
  and g36 (n659, n_34, \in3[113] );
  not g37 (n_38, \in3[111] );
  and g38 (n660, \in2[111] , n_38);
  not g39 (n_39, \in2[111] );
  and g40 (n661, n_39, \in3[111] );
  not g41 (n_41, \in2[110] );
  and g42 (n662, n_41, \in3[110] );
  not g43 (n_43, n661);
  not g44 (n_44, n662);
  and g45 (n663, n_43, n_44);
  not g46 (n_46, \in2[109] );
  and g47 (n664, n_46, \in3[109] );
  not g48 (n_50, \in3[108] );
  and g49 (n665, \in2[108] , n_50);
  not g50 (n_51, n664);
  and g51 (n666, n_51, n665);
  not g52 (n_52, \in3[109] );
  and g53 (n667, \in2[109] , n_52);
  not g54 (n_53, n666);
  not g55 (n_54, n667);
  and g56 (n668, n_53, n_54);
  not g57 (n_55, n668);
  and g58 (n669, n663, n_55);
  not g59 (n_56, \in3[110] );
  and g60 (n670, n_56, n_43);
  and g61 (n671, \in2[110] , n670);
  not g62 (n_59, \in3[103] );
  and g63 (n672, \in2[103] , n_59);
  not g64 (n_60, \in2[103] );
  and g65 (n673, n_60, \in3[103] );
  not g66 (n_62, \in2[102] );
  and g67 (n674, n_62, \in3[102] );
  not g68 (n_64, n673);
  not g69 (n_65, n674);
  and g70 (n675, n_64, n_65);
  not g71 (n_67, \in2[101] );
  and g72 (n676, n_67, \in3[101] );
  not g73 (n_71, \in3[100] );
  and g74 (n677, \in2[100] , n_71);
  not g75 (n_72, n676);
  and g76 (n678, n_72, n677);
  not g77 (n_73, \in3[101] );
  and g78 (n679, \in2[101] , n_73);
  not g79 (n_74, n678);
  not g80 (n_75, n679);
  and g81 (n680, n_74, n_75);
  not g82 (n_76, n680);
  and g83 (n681, n675, n_76);
  not g84 (n_77, \in3[102] );
  and g85 (n682, n_77, n_64);
  and g86 (n683, \in2[102] , n682);
  not g87 (n_79, \in2[96] );
  and g88 (n684, n_79, \in3[96] );
  not g89 (n_82, \in2[99] );
  and g90 (n685, n_82, \in3[99] );
  not g91 (n_85, \in2[98] );
  and g92 (n686, n_85, \in3[98] );
  not g93 (n_87, n685);
  not g94 (n_88, n686);
  and g95 (n687, n_87, n_88);
  not g96 (n_90, \in2[97] );
  and g97 (n688, n_90, \in3[97] );
  not g98 (n_94, \in3[95] );
  and g99 (n689, \in2[95] , n_94);
  not g100 (n_95, \in2[95] );
  and g101 (n690, n_95, \in3[95] );
  not g102 (n_97, \in2[94] );
  and g103 (n691, n_97, \in3[94] );
  not g104 (n_99, n690);
  not g105 (n_100, n691);
  and g106 (n692, n_99, n_100);
  not g107 (n_102, \in2[93] );
  and g108 (n693, n_102, \in3[93] );
  not g109 (n_106, \in3[92] );
  and g110 (n694, \in2[92] , n_106);
  not g111 (n_107, n693);
  and g112 (n695, n_107, n694);
  not g113 (n_108, \in3[93] );
  and g114 (n696, \in2[93] , n_108);
  not g115 (n_109, n695);
  not g116 (n_110, n696);
  and g117 (n697, n_109, n_110);
  not g118 (n_111, n697);
  and g119 (n698, n692, n_111);
  not g120 (n_112, \in3[94] );
  and g121 (n699, n_112, n_99);
  and g122 (n700, \in2[94] , n699);
  not g123 (n_115, \in3[87] );
  and g124 (n701, \in2[87] , n_115);
  not g125 (n_116, \in2[87] );
  and g126 (n702, n_116, \in3[87] );
  not g127 (n_118, \in2[86] );
  and g128 (n703, n_118, \in3[86] );
  not g129 (n_120, n702);
  not g130 (n_121, n703);
  and g131 (n704, n_120, n_121);
  not g132 (n_123, \in2[85] );
  and g133 (n705, n_123, \in3[85] );
  not g134 (n_127, \in3[84] );
  and g135 (n706, \in2[84] , n_127);
  not g136 (n_128, n705);
  and g137 (n707, n_128, n706);
  not g138 (n_129, \in3[85] );
  and g139 (n708, \in2[85] , n_129);
  not g140 (n_130, n707);
  not g141 (n_131, n708);
  and g142 (n709, n_130, n_131);
  not g143 (n_132, n709);
  and g144 (n710, n704, n_132);
  not g145 (n_133, \in3[86] );
  and g146 (n711, n_133, n_120);
  and g147 (n712, \in2[86] , n711);
  not g148 (n_135, \in2[80] );
  and g149 (n713, n_135, \in3[80] );
  not g150 (n_138, \in2[83] );
  and g151 (n714, n_138, \in3[83] );
  not g152 (n_141, \in2[82] );
  and g153 (n715, n_141, \in3[82] );
  not g154 (n_143, n714);
  not g155 (n_144, n715);
  and g156 (n716, n_143, n_144);
  not g157 (n_146, \in2[81] );
  and g158 (n717, n_146, \in3[81] );
  not g159 (n_150, \in3[79] );
  and g160 (n718, \in2[79] , n_150);
  not g161 (n_151, \in2[79] );
  and g162 (n719, n_151, \in3[79] );
  not g163 (n_153, \in2[78] );
  and g164 (n720, n_153, \in3[78] );
  not g165 (n_155, n719);
  not g166 (n_156, n720);
  and g167 (n721, n_155, n_156);
  not g168 (n_158, \in2[77] );
  and g169 (n722, n_158, \in3[77] );
  not g170 (n_162, \in3[76] );
  and g171 (n723, \in2[76] , n_162);
  not g172 (n_163, n722);
  and g173 (n724, n_163, n723);
  not g174 (n_164, \in3[77] );
  and g175 (n725, \in2[77] , n_164);
  not g176 (n_165, n724);
  not g177 (n_166, n725);
  and g178 (n726, n_165, n_166);
  not g179 (n_167, n726);
  and g180 (n727, n721, n_167);
  not g181 (n_168, \in3[78] );
  and g182 (n728, n_168, n_155);
  and g183 (n729, \in2[78] , n728);
  not g184 (n_171, \in3[71] );
  and g185 (n730, \in2[71] , n_171);
  not g186 (n_172, \in2[71] );
  and g187 (n731, n_172, \in3[71] );
  not g188 (n_174, \in2[70] );
  and g189 (n732, n_174, \in3[70] );
  not g190 (n_176, n731);
  not g191 (n_177, n732);
  and g192 (n733, n_176, n_177);
  not g193 (n_179, \in2[69] );
  and g194 (n734, n_179, \in3[69] );
  not g195 (n_183, \in3[68] );
  and g196 (n735, \in2[68] , n_183);
  not g197 (n_184, n734);
  and g198 (n736, n_184, n735);
  not g199 (n_185, \in3[69] );
  and g200 (n737, \in2[69] , n_185);
  not g201 (n_186, n736);
  not g202 (n_187, n737);
  and g203 (n738, n_186, n_187);
  not g204 (n_188, n738);
  and g205 (n739, n733, n_188);
  not g206 (n_189, \in3[70] );
  and g207 (n740, n_189, n_176);
  and g208 (n741, \in2[70] , n740);
  not g209 (n_191, \in2[67] );
  and g210 (n742, n_191, \in3[67] );
  not g211 (n_194, \in2[66] );
  and g212 (n743, n_194, \in3[66] );
  not g213 (n_196, n742);
  not g214 (n_197, n743);
  and g215 (n744, n_196, n_197);
  not g216 (n_199, \in2[65] );
  and g217 (n745, n_199, \in3[65] );
  not g218 (n_203, \in3[63] );
  and g219 (n746, \in2[63] , n_203);
  not g220 (n_204, \in2[63] );
  and g221 (n747, n_204, \in3[63] );
  not g222 (n_206, \in2[62] );
  and g223 (n748, n_206, \in3[62] );
  not g224 (n_208, n747);
  not g225 (n_209, n748);
  and g226 (n749, n_208, n_209);
  not g227 (n_211, \in2[60] );
  and g228 (n750, n_211, \in3[60] );
  not g229 (n_214, \in2[61] );
  and g230 (n751, n_214, \in3[61] );
  not g231 (n_216, n750);
  not g232 (n_217, n751);
  and g233 (n752, n_216, n_217);
  and g234 (n753, n749, n752);
  not g235 (n_220, \in3[59] );
  and g236 (n754, \in2[59] , n_220);
  not g237 (n_221, \in2[59] );
  and g238 (n755, n_221, \in3[59] );
  not g239 (n_223, \in2[58] );
  and g240 (n756, n_223, \in3[58] );
  not g241 (n_225, n755);
  not g242 (n_226, n756);
  and g243 (n757, n_225, n_226);
  not g244 (n_228, \in2[57] );
  and g245 (n758, n_228, \in3[57] );
  not g246 (n_232, \in3[56] );
  and g247 (n759, \in2[56] , n_232);
  not g248 (n_233, n758);
  and g249 (n760, n_233, n759);
  not g250 (n_234, \in3[57] );
  and g251 (n761, \in2[57] , n_234);
  not g252 (n_235, n760);
  not g253 (n_236, n761);
  and g254 (n762, n_235, n_236);
  not g255 (n_237, \in3[58] );
  and g256 (n763, \in2[58] , n_237);
  not g257 (n_238, n763);
  and g258 (n764, n762, n_238);
  not g259 (n_239, n764);
  and g260 (n765, n757, n_239);
  not g261 (n_240, n754);
  not g262 (n_241, n765);
  and g263 (n766, n_240, n_241);
  not g264 (n_242, n766);
  and g265 (n767, n753, n_242);
  not g266 (n_243, \in3[60] );
  and g267 (n768, \in2[60] , n_243);
  and g268 (n769, n_217, n768);
  not g269 (n_244, \in3[61] );
  and g270 (n770, \in2[61] , n_244);
  not g271 (n_245, n769);
  not g272 (n_246, n770);
  and g273 (n771, n_245, n_246);
  not g274 (n_247, n771);
  and g275 (n772, n749, n_247);
  not g276 (n_248, \in3[62] );
  and g277 (n773, n_248, n_208);
  and g278 (n774, \in2[62] , n773);
  not g279 (n_251, \in3[47] );
  and g280 (n775, \in2[47] , n_251);
  not g281 (n_252, \in2[47] );
  and g282 (n776, n_252, \in3[47] );
  not g283 (n_254, \in2[46] );
  and g284 (n777, n_254, \in3[46] );
  not g285 (n_256, n776);
  not g286 (n_257, n777);
  and g287 (n778, n_256, n_257);
  not g288 (n_259, \in2[44] );
  and g289 (n779, n_259, \in3[44] );
  not g290 (n_262, \in2[45] );
  and g291 (n780, n_262, \in3[45] );
  not g292 (n_264, n779);
  not g293 (n_265, n780);
  and g294 (n781, n_264, n_265);
  and g295 (n782, n778, n781);
  not g296 (n_268, \in3[43] );
  and g297 (n783, \in2[43] , n_268);
  not g298 (n_269, \in2[43] );
  and g299 (n784, n_269, \in3[43] );
  not g300 (n_271, \in2[42] );
  and g301 (n785, n_271, \in3[42] );
  not g302 (n_273, n784);
  not g303 (n_274, n785);
  and g304 (n786, n_273, n_274);
  not g305 (n_276, \in2[41] );
  and g306 (n787, n_276, \in3[41] );
  not g307 (n_280, \in3[40] );
  and g308 (n788, \in2[40] , n_280);
  not g309 (n_281, n787);
  and g310 (n789, n_281, n788);
  not g311 (n_282, \in3[41] );
  and g312 (n790, \in2[41] , n_282);
  not g313 (n_283, n789);
  not g314 (n_284, n790);
  and g315 (n791, n_283, n_284);
  not g316 (n_285, \in3[42] );
  and g317 (n792, \in2[42] , n_285);
  not g318 (n_286, n792);
  and g319 (n793, n791, n_286);
  not g320 (n_287, n793);
  and g321 (n794, n786, n_287);
  not g322 (n_288, n783);
  not g323 (n_289, n794);
  and g324 (n795, n_288, n_289);
  not g325 (n_290, n795);
  and g326 (n796, n782, n_290);
  not g327 (n_291, \in3[44] );
  and g328 (n797, \in2[44] , n_291);
  and g329 (n798, n_265, n797);
  not g330 (n_292, \in3[45] );
  and g331 (n799, \in2[45] , n_292);
  not g332 (n_293, n798);
  not g333 (n_294, n799);
  and g334 (n800, n_293, n_294);
  not g335 (n_295, n800);
  and g336 (n801, n778, n_295);
  not g337 (n_296, \in3[46] );
  and g338 (n802, n_296, n_256);
  and g339 (n803, \in2[46] , n802);
  not g340 (n_298, \in2[32] );
  and g341 (n804, n_298, \in3[32] );
  not g342 (n_301, \in2[31] );
  and g343 (n805, n_301, \in3[31] );
  not g344 (n_304, \in2[30] );
  and g345 (n806, n_304, \in3[30] );
  not g346 (n_307, \in2[29] );
  and g347 (n807, n_307, \in3[29] );
  not g348 (n_310, \in2[28] );
  and g349 (n808, n_310, \in3[28] );
  not g350 (n_313, \in2[27] );
  and g351 (n809, n_313, \in3[27] );
  not g352 (n_316, \in2[26] );
  and g353 (n810, n_316, \in3[26] );
  not g354 (n_319, \in2[23] );
  and g355 (n811, n_319, \in3[23] );
  not g356 (n_322, \in2[22] );
  and g357 (n812, n_322, \in3[22] );
  not g358 (n_325, \in2[21] );
  and g359 (n813, n_325, \in3[21] );
  not g360 (n_328, \in2[20] );
  and g361 (n814, n_328, \in3[20] );
  not g362 (n_331, \in2[19] );
  and g363 (n815, n_331, \in3[19] );
  not g364 (n_334, \in2[18] );
  and g365 (n816, n_334, \in3[18] );
  not g366 (n_337, \in2[15] );
  and g367 (n817, n_337, \in3[15] );
  not g368 (n_340, \in2[14] );
  and g369 (n818, n_340, \in3[14] );
  not g370 (n_343, \in2[13] );
  and g371 (n819, n_343, \in3[13] );
  not g372 (n_346, \in2[12] );
  and g373 (n820, n_346, \in3[12] );
  not g374 (n_349, \in2[11] );
  and g375 (n821, n_349, \in3[11] );
  not g376 (n_352, \in2[10] );
  and g377 (n822, n_352, \in3[10] );
  not g378 (n_355, \in2[7] );
  and g379 (n823, n_355, \in3[7] );
  not g380 (n_358, \in2[6] );
  and g381 (n824, n_358, \in3[6] );
  not g382 (n_361, \in2[3] );
  and g383 (n825, n_361, \in3[3] );
  not g384 (n_365, \in3[0] );
  and g385 (n826, \in2[0] , n_365);
  and g386 (n827, \in2[1] , n826);
  not g387 (n_368, n827);
  and g388 (n828, \in3[1] , n_368);
  not g389 (n_370, \in2[2] );
  and g390 (n829, n_370, \in3[2] );
  not g391 (n_372, \in2[1] );
  not g392 (n_373, n826);
  and g393 (n830, n_372, n_373);
  not g394 (n_374, n829);
  not g395 (n_375, n830);
  and g396 (n831, n_374, n_375);
  not g397 (n_376, n828);
  and g398 (n832, n_376, n831);
  not g399 (n_377, \in3[2] );
  and g400 (n833, \in2[2] , n_377);
  not g401 (n_378, n832);
  not g402 (n_379, n833);
  and g403 (n834, n_378, n_379);
  not g404 (n_380, n825);
  not g405 (n_381, n834);
  and g406 (n835, n_380, n_381);
  not g407 (n_382, \in3[3] );
  and g408 (n836, \in2[3] , n_382);
  not g409 (n_383, n835);
  not g410 (n_384, n836);
  and g411 (n837, n_383, n_384);
  not g412 (n_386, \in2[4] );
  and g413 (n838, n_386, n837);
  not g414 (n_388, \in3[4] );
  not g415 (n_389, n838);
  and g416 (n839, n_388, n_389);
  not g417 (n_390, n837);
  and g418 (n840, \in2[4] , n_390);
  not g419 (n_391, n839);
  not g420 (n_392, n840);
  and g421 (n841, n_391, n_392);
  not g422 (n_394, \in2[5] );
  and g423 (n842, n_394, n841);
  not g424 (n_396, \in3[5] );
  not g425 (n_397, n842);
  and g426 (n843, n_396, n_397);
  not g427 (n_398, n841);
  and g428 (n844, \in2[5] , n_398);
  not g429 (n_399, n843);
  not g430 (n_400, n844);
  and g431 (n845, n_399, n_400);
  not g432 (n_401, n824);
  not g433 (n_402, n845);
  and g434 (n846, n_401, n_402);
  not g435 (n_403, \in3[6] );
  and g436 (n847, \in2[6] , n_403);
  not g437 (n_404, n846);
  not g438 (n_405, n847);
  and g439 (n848, n_404, n_405);
  not g440 (n_406, n823);
  not g441 (n_407, n848);
  and g442 (n849, n_406, n_407);
  not g443 (n_408, \in3[7] );
  and g444 (n850, \in2[7] , n_408);
  not g445 (n_409, n849);
  not g446 (n_410, n850);
  and g447 (n851, n_409, n_410);
  not g448 (n_412, \in2[8] );
  and g449 (n852, n_412, n851);
  not g450 (n_414, \in3[8] );
  not g451 (n_415, n852);
  and g452 (n853, n_414, n_415);
  not g453 (n_416, n851);
  and g454 (n854, \in2[8] , n_416);
  not g455 (n_417, n853);
  not g456 (n_418, n854);
  and g457 (n855, n_417, n_418);
  not g458 (n_420, \in2[9] );
  and g459 (n856, n_420, n855);
  not g460 (n_422, \in3[9] );
  not g461 (n_423, n856);
  and g462 (n857, n_422, n_423);
  not g463 (n_424, n855);
  and g464 (n858, \in2[9] , n_424);
  not g465 (n_425, n857);
  not g466 (n_426, n858);
  and g467 (n859, n_425, n_426);
  not g468 (n_427, n822);
  not g469 (n_428, n859);
  and g470 (n860, n_427, n_428);
  not g471 (n_429, \in3[10] );
  and g472 (n861, \in2[10] , n_429);
  not g473 (n_430, n860);
  not g474 (n_431, n861);
  and g475 (n862, n_430, n_431);
  not g476 (n_432, n821);
  not g477 (n_433, n862);
  and g478 (n863, n_432, n_433);
  not g479 (n_434, \in3[11] );
  and g480 (n864, \in2[11] , n_434);
  not g481 (n_435, n863);
  not g482 (n_436, n864);
  and g483 (n865, n_435, n_436);
  not g484 (n_437, n820);
  not g485 (n_438, n865);
  and g486 (n866, n_437, n_438);
  not g487 (n_439, \in3[12] );
  and g488 (n867, \in2[12] , n_439);
  not g489 (n_440, n866);
  not g490 (n_441, n867);
  and g491 (n868, n_440, n_441);
  not g492 (n_442, n819);
  not g493 (n_443, n868);
  and g494 (n869, n_442, n_443);
  not g495 (n_444, \in3[13] );
  and g496 (n870, \in2[13] , n_444);
  not g497 (n_445, n869);
  not g498 (n_446, n870);
  and g499 (n871, n_445, n_446);
  not g500 (n_447, n818);
  not g501 (n_448, n871);
  and g502 (n872, n_447, n_448);
  not g503 (n_449, \in3[14] );
  and g504 (n873, \in2[14] , n_449);
  not g505 (n_450, n872);
  not g506 (n_451, n873);
  and g507 (n874, n_450, n_451);
  not g508 (n_452, n817);
  not g509 (n_453, n874);
  and g510 (n875, n_452, n_453);
  not g511 (n_454, \in3[15] );
  and g512 (n876, \in2[15] , n_454);
  not g513 (n_455, n875);
  not g514 (n_456, n876);
  and g515 (n877, n_455, n_456);
  not g516 (n_458, \in2[16] );
  and g517 (n878, n_458, n877);
  not g518 (n_460, \in3[16] );
  not g519 (n_461, n878);
  and g520 (n879, n_460, n_461);
  not g521 (n_462, n877);
  and g522 (n880, \in2[16] , n_462);
  not g523 (n_463, n879);
  not g524 (n_464, n880);
  and g525 (n881, n_463, n_464);
  not g526 (n_466, \in2[17] );
  and g527 (n882, n_466, n881);
  not g528 (n_468, \in3[17] );
  not g529 (n_469, n882);
  and g530 (n883, n_468, n_469);
  not g531 (n_470, n881);
  and g532 (n884, \in2[17] , n_470);
  not g533 (n_471, n883);
  not g534 (n_472, n884);
  and g535 (n885, n_471, n_472);
  not g536 (n_473, n816);
  not g537 (n_474, n885);
  and g538 (n886, n_473, n_474);
  not g539 (n_475, \in3[18] );
  and g540 (n887, \in2[18] , n_475);
  not g541 (n_476, n886);
  not g542 (n_477, n887);
  and g543 (n888, n_476, n_477);
  not g544 (n_478, n815);
  not g545 (n_479, n888);
  and g546 (n889, n_478, n_479);
  not g547 (n_480, \in3[19] );
  and g548 (n890, \in2[19] , n_480);
  not g549 (n_481, n889);
  not g550 (n_482, n890);
  and g551 (n891, n_481, n_482);
  not g552 (n_483, n814);
  not g553 (n_484, n891);
  and g554 (n892, n_483, n_484);
  not g555 (n_485, \in3[20] );
  and g556 (n893, \in2[20] , n_485);
  not g557 (n_486, n892);
  not g558 (n_487, n893);
  and g559 (n894, n_486, n_487);
  not g560 (n_488, n813);
  not g561 (n_489, n894);
  and g562 (n895, n_488, n_489);
  not g563 (n_490, \in3[21] );
  and g564 (n896, \in2[21] , n_490);
  not g565 (n_491, n895);
  not g566 (n_492, n896);
  and g567 (n897, n_491, n_492);
  not g568 (n_493, n812);
  not g569 (n_494, n897);
  and g570 (n898, n_493, n_494);
  not g571 (n_495, \in3[22] );
  and g572 (n899, \in2[22] , n_495);
  not g573 (n_496, n898);
  not g574 (n_497, n899);
  and g575 (n900, n_496, n_497);
  not g576 (n_498, n811);
  not g577 (n_499, n900);
  and g578 (n901, n_498, n_499);
  not g579 (n_500, \in3[23] );
  and g580 (n902, \in2[23] , n_500);
  not g581 (n_501, n901);
  not g582 (n_502, n902);
  and g583 (n903, n_501, n_502);
  not g584 (n_504, \in2[24] );
  and g585 (n904, n_504, n903);
  not g586 (n_506, \in3[24] );
  not g587 (n_507, n904);
  and g588 (n905, n_506, n_507);
  not g589 (n_508, n903);
  and g590 (n906, \in2[24] , n_508);
  not g591 (n_509, n905);
  not g592 (n_510, n906);
  and g593 (n907, n_509, n_510);
  not g594 (n_512, \in2[25] );
  and g595 (n908, n_512, n907);
  not g596 (n_514, \in3[25] );
  not g597 (n_515, n908);
  and g598 (n909, n_514, n_515);
  not g599 (n_516, n907);
  and g600 (n910, \in2[25] , n_516);
  not g601 (n_517, n909);
  not g602 (n_518, n910);
  and g603 (n911, n_517, n_518);
  not g604 (n_519, n810);
  not g605 (n_520, n911);
  and g606 (n912, n_519, n_520);
  not g607 (n_521, \in3[26] );
  and g608 (n913, \in2[26] , n_521);
  not g609 (n_522, n912);
  not g610 (n_523, n913);
  and g611 (n914, n_522, n_523);
  not g612 (n_524, n809);
  not g613 (n_525, n914);
  and g614 (n915, n_524, n_525);
  not g615 (n_526, \in3[27] );
  and g616 (n916, \in2[27] , n_526);
  not g617 (n_527, n915);
  not g618 (n_528, n916);
  and g619 (n917, n_527, n_528);
  not g620 (n_529, n808);
  not g621 (n_530, n917);
  and g622 (n918, n_529, n_530);
  not g623 (n_531, \in3[28] );
  and g624 (n919, \in2[28] , n_531);
  not g625 (n_532, n918);
  not g626 (n_533, n919);
  and g627 (n920, n_532, n_533);
  not g628 (n_534, n807);
  not g629 (n_535, n920);
  and g630 (n921, n_534, n_535);
  not g631 (n_536, \in3[29] );
  and g632 (n922, \in2[29] , n_536);
  not g633 (n_537, n921);
  not g634 (n_538, n922);
  and g635 (n923, n_537, n_538);
  not g636 (n_539, n806);
  not g637 (n_540, n923);
  and g638 (n924, n_539, n_540);
  not g639 (n_541, \in3[30] );
  and g640 (n925, \in2[30] , n_541);
  not g641 (n_542, n924);
  not g642 (n_543, n925);
  and g643 (n926, n_542, n_543);
  not g644 (n_544, n805);
  not g645 (n_545, n926);
  and g646 (n927, n_544, n_545);
  not g647 (n_546, \in3[31] );
  and g648 (n928, \in2[31] , n_546);
  not g649 (n_547, n927);
  not g650 (n_548, n928);
  and g651 (n929, n_547, n_548);
  not g652 (n_550, \in2[39] );
  and g653 (n930, n_550, \in3[39] );
  not g654 (n_553, \in2[38] );
  and g655 (n931, n_553, \in3[38] );
  not g656 (n_555, n930);
  not g657 (n_556, n931);
  and g658 (n932, n_555, n_556);
  not g659 (n_558, \in2[36] );
  and g660 (n933, n_558, \in3[36] );
  not g661 (n_561, \in2[37] );
  and g662 (n934, n_561, \in3[37] );
  not g663 (n_563, n933);
  not g664 (n_564, n934);
  and g665 (n935, n_563, n_564);
  and g666 (n936, n932, n935);
  not g667 (n_566, \in2[33] );
  and g668 (n937, n_566, \in3[33] );
  not g669 (n_569, \in2[35] );
  and g670 (n938, n_569, \in3[35] );
  not g671 (n_572, \in2[34] );
  and g672 (n939, n_572, \in3[34] );
  not g673 (n_574, n938);
  not g674 (n_575, n939);
  and g675 (n940, n_574, n_575);
  not g676 (n_576, n937);
  not g683 (n_579, \in3[39] );
  and g684 (n945, \in2[39] , n_579);
  not g685 (n_580, \in3[36] );
  and g686 (n946, \in2[36] , n_580);
  and g687 (n947, n_564, n946);
  not g688 (n_581, \in3[37] );
  and g689 (n948, \in2[37] , n_581);
  not g690 (n_582, n947);
  not g691 (n_583, n948);
  and g692 (n949, n_582, n_583);
  not g693 (n_584, n949);
  and g694 (n950, n932, n_584);
  not g695 (n_585, \in3[38] );
  and g696 (n951, n_585, n_555);
  and g697 (n952, \in2[38] , n951);
  not g698 (n_586, \in3[35] );
  and g699 (n953, \in2[35] , n_586);
  not g700 (n_587, \in3[32] );
  and g701 (n954, n_587, n_576);
  and g702 (n955, \in2[32] , n954);
  not g703 (n_588, \in3[33] );
  and g704 (n956, \in2[33] , n_588);
  not g705 (n_589, n955);
  not g706 (n_590, n956);
  and g707 (n957, n_589, n_590);
  not g708 (n_591, \in3[34] );
  and g709 (n958, \in2[34] , n_591);
  not g710 (n_592, n958);
  and g711 (n959, n957, n_592);
  not g712 (n_593, n959);
  and g713 (n960, n940, n_593);
  not g714 (n_594, n953);
  not g715 (n_595, n960);
  and g716 (n961, n_594, n_595);
  not g717 (n_596, n961);
  and g718 (n962, n936, n_596);
  not g728 (n_602, \in2[40] );
  and g729 (n967, n_602, \in3[40] );
  not g745 (n_611, \in2[48] );
  and g746 (n976, n_611, \in3[48] );
  not g747 (n_614, \in2[55] );
  and g748 (n977, n_614, \in3[55] );
  not g749 (n_617, \in2[54] );
  and g750 (n978, n_617, \in3[54] );
  not g751 (n_619, n977);
  not g752 (n_620, n978);
  and g753 (n979, n_619, n_620);
  not g754 (n_622, \in2[53] );
  and g755 (n980, n_622, \in3[53] );
  not g756 (n_625, \in2[52] );
  and g757 (n981, n_625, \in3[52] );
  not g758 (n_627, n980);
  not g759 (n_628, n981);
  and g760 (n982, n_627, n_628);
  and g761 (n983, n979, n982);
  not g762 (n_630, \in2[49] );
  and g763 (n984, n_630, \in3[49] );
  not g764 (n_633, \in2[51] );
  and g765 (n985, n_633, \in3[51] );
  not g766 (n_636, \in2[50] );
  and g767 (n986, n_636, \in3[50] );
  not g768 (n_638, n985);
  not g769 (n_639, n986);
  and g770 (n987, n_638, n_639);
  not g771 (n_640, n984);
  not g778 (n_643, \in3[55] );
  and g779 (n992, \in2[55] , n_643);
  not g780 (n_644, \in3[51] );
  and g781 (n993, \in2[51] , n_644);
  not g782 (n_645, \in3[48] );
  and g783 (n994, n_645, n_640);
  and g784 (n995, \in2[48] , n994);
  not g785 (n_646, \in3[49] );
  and g786 (n996, \in2[49] , n_646);
  not g787 (n_647, n995);
  not g788 (n_648, n996);
  and g789 (n997, n_647, n_648);
  not g790 (n_649, \in3[50] );
  and g791 (n998, \in2[50] , n_649);
  not g792 (n_650, n998);
  and g793 (n999, n997, n_650);
  not g794 (n_651, n999);
  and g795 (n1000, n987, n_651);
  not g796 (n_652, n993);
  not g797 (n_653, n1000);
  and g798 (n1001, n_652, n_653);
  not g799 (n_654, n1001);
  and g800 (n1002, n983, n_654);
  not g801 (n_655, \in3[52] );
  and g802 (n1003, \in2[52] , n_655);
  and g803 (n1004, n_627, n1003);
  not g804 (n_656, \in3[53] );
  and g805 (n1005, \in2[53] , n_656);
  not g806 (n_657, n1004);
  not g807 (n_658, n1005);
  and g808 (n1006, n_657, n_658);
  not g809 (n_659, \in3[54] );
  and g810 (n1007, \in2[54] , n_659);
  not g811 (n_660, n1007);
  and g812 (n1008, n1006, n_660);
  not g813 (n_661, n1008);
  and g814 (n1009, n979, n_661);
  not g822 (n_666, \in2[56] );
  and g823 (n1013, n_666, \in3[56] );
  not g839 (n_675, \in2[64] );
  and g840 (n1022, n_675, \in3[64] );
  not g844 (n_679, n745);
  not g847 (n_680, \in3[67] );
  and g848 (n1026, \in2[67] , n_680);
  not g849 (n_681, \in3[64] );
  and g850 (n1027, \in2[64] , n_681);
  and g851 (n1028, n_679, n1027);
  not g852 (n_682, \in3[65] );
  and g853 (n1029, \in2[65] , n_682);
  not g854 (n_683, n1028);
  not g855 (n_684, n1029);
  and g856 (n1030, n_683, n_684);
  not g857 (n_685, \in3[66] );
  and g858 (n1031, \in2[66] , n_685);
  not g859 (n_686, n1031);
  and g860 (n1032, n1030, n_686);
  not g861 (n_687, n1032);
  and g862 (n1033, n744, n_687);
  not g863 (n_688, n1026);
  not g864 (n_689, n1033);
  and g865 (n1034, n_688, n_689);
  not g866 (n_690, n1025);
  and g867 (n1035, n_690, n1034);
  not g868 (n_691, \in2[68] );
  and g869 (n1036, n_691, \in3[68] );
  not g882 (n_699, \in2[75] );
  and g883 (n1043, n_699, \in3[75] );
  not g884 (n_702, \in2[74] );
  and g885 (n1044, n_702, \in3[74] );
  not g886 (n_704, n1043);
  not g887 (n_705, n1044);
  and g888 (n1045, n_704, n_705);
  not g889 (n_707, \in2[73] );
  and g890 (n1046, n_707, \in3[73] );
  not g891 (n_710, \in2[72] );
  and g892 (n1047, n_710, \in3[72] );
  not g893 (n_712, n1046);
  not g899 (n_715, \in3[75] );
  and g900 (n1051, \in2[75] , n_715);
  not g901 (n_716, \in3[72] );
  and g902 (n1052, \in2[72] , n_716);
  and g903 (n1053, n_712, n1052);
  not g904 (n_717, \in3[73] );
  and g905 (n1054, \in2[73] , n_717);
  not g906 (n_718, n1053);
  not g907 (n_719, n1054);
  and g908 (n1055, n_718, n_719);
  not g909 (n_720, \in3[74] );
  and g910 (n1056, \in2[74] , n_720);
  not g911 (n_721, n1056);
  and g912 (n1057, n1055, n_721);
  not g913 (n_722, n1057);
  and g914 (n1058, n1045, n_722);
  not g915 (n_723, n1051);
  not g916 (n_724, n1058);
  and g917 (n1059, n_723, n_724);
  not g918 (n_725, n1050);
  and g919 (n1060, n_725, n1059);
  not g920 (n_726, \in2[76] );
  and g921 (n1061, n_726, \in3[76] );
  not g934 (n_733, n717);
  not g940 (n_736, \in3[83] );
  and g941 (n1071, \in2[83] , n_736);
  not g942 (n_737, \in3[80] );
  and g943 (n1072, n_737, n_733);
  and g944 (n1073, \in2[80] , n1072);
  not g945 (n_738, \in3[81] );
  and g946 (n1074, \in2[81] , n_738);
  not g947 (n_739, n1073);
  not g948 (n_740, n1074);
  and g949 (n1075, n_739, n_740);
  not g950 (n_741, \in3[82] );
  and g951 (n1076, \in2[82] , n_741);
  not g952 (n_742, n1076);
  and g953 (n1077, n1075, n_742);
  not g954 (n_743, n1077);
  and g955 (n1078, n716, n_743);
  not g956 (n_744, n1071);
  not g957 (n_745, n1078);
  and g958 (n1079, n_744, n_745);
  not g959 (n_746, n1070);
  and g960 (n1080, n_746, n1079);
  not g961 (n_747, \in2[84] );
  and g962 (n1081, n_747, \in3[84] );
  not g975 (n_755, \in2[91] );
  and g976 (n1088, n_755, \in3[91] );
  not g977 (n_758, \in2[90] );
  and g978 (n1089, n_758, \in3[90] );
  not g979 (n_760, n1088);
  not g980 (n_761, n1089);
  and g981 (n1090, n_760, n_761);
  not g982 (n_763, \in2[89] );
  and g983 (n1091, n_763, \in3[89] );
  not g984 (n_766, \in2[88] );
  and g985 (n1092, n_766, \in3[88] );
  not g986 (n_768, n1091);
  not g992 (n_771, \in3[91] );
  and g993 (n1096, \in2[91] , n_771);
  not g994 (n_772, \in3[88] );
  and g995 (n1097, \in2[88] , n_772);
  and g996 (n1098, n_768, n1097);
  not g997 (n_773, \in3[89] );
  and g998 (n1099, \in2[89] , n_773);
  not g999 (n_774, n1098);
  not g1000 (n_775, n1099);
  and g1001 (n1100, n_774, n_775);
  not g1002 (n_776, \in3[90] );
  and g1003 (n1101, \in2[90] , n_776);
  not g1004 (n_777, n1101);
  and g1005 (n1102, n1100, n_777);
  not g1006 (n_778, n1102);
  and g1007 (n1103, n1090, n_778);
  not g1008 (n_779, n1096);
  not g1009 (n_780, n1103);
  and g1010 (n1104, n_779, n_780);
  not g1011 (n_781, n1095);
  and g1012 (n1105, n_781, n1104);
  not g1013 (n_782, \in2[92] );
  and g1014 (n1106, n_782, \in3[92] );
  not g1027 (n_789, n688);
  not g1033 (n_792, \in3[99] );
  and g1034 (n1116, \in2[99] , n_792);
  not g1035 (n_793, \in3[96] );
  and g1036 (n1117, n_793, n_789);
  and g1037 (n1118, \in2[96] , n1117);
  not g1038 (n_794, \in3[97] );
  and g1039 (n1119, \in2[97] , n_794);
  not g1040 (n_795, n1118);
  not g1041 (n_796, n1119);
  and g1042 (n1120, n_795, n_796);
  not g1043 (n_797, \in3[98] );
  and g1044 (n1121, \in2[98] , n_797);
  not g1045 (n_798, n1121);
  and g1046 (n1122, n1120, n_798);
  not g1047 (n_799, n1122);
  and g1048 (n1123, n687, n_799);
  not g1049 (n_800, n1116);
  not g1050 (n_801, n1123);
  and g1051 (n1124, n_800, n_801);
  not g1052 (n_802, n1115);
  and g1053 (n1125, n_802, n1124);
  not g1054 (n_803, \in2[100] );
  and g1055 (n1126, n_803, \in3[100] );
  not g1068 (n_811, \in2[107] );
  and g1069 (n1133, n_811, \in3[107] );
  not g1070 (n_814, \in2[106] );
  and g1071 (n1134, n_814, \in3[106] );
  not g1072 (n_816, n1133);
  not g1073 (n_817, n1134);
  and g1074 (n1135, n_816, n_817);
  not g1075 (n_819, \in2[105] );
  and g1076 (n1136, n_819, \in3[105] );
  not g1077 (n_822, \in2[104] );
  and g1078 (n1137, n_822, \in3[104] );
  not g1079 (n_824, n1136);
  not g1085 (n_827, \in3[107] );
  and g1086 (n1141, \in2[107] , n_827);
  not g1087 (n_828, \in3[104] );
  and g1088 (n1142, \in2[104] , n_828);
  and g1089 (n1143, n_824, n1142);
  not g1090 (n_829, \in3[105] );
  and g1091 (n1144, \in2[105] , n_829);
  not g1092 (n_830, n1143);
  not g1093 (n_831, n1144);
  and g1094 (n1145, n_830, n_831);
  not g1095 (n_832, \in3[106] );
  and g1096 (n1146, \in2[106] , n_832);
  not g1097 (n_833, n1146);
  and g1098 (n1147, n1145, n_833);
  not g1099 (n_834, n1147);
  and g1100 (n1148, n1135, n_834);
  not g1101 (n_835, n1141);
  not g1102 (n_836, n1148);
  and g1103 (n1149, n_835, n_836);
  not g1104 (n_837, n1140);
  and g1105 (n1150, n_837, n1149);
  not g1106 (n_838, \in2[108] );
  and g1107 (n1151, n_838, \in3[108] );
  not g1120 (n_845, n659);
  not g1126 (n_848, \in3[115] );
  and g1127 (n1161, \in2[115] , n_848);
  not g1128 (n_849, \in3[112] );
  and g1129 (n1162, n_849, n_845);
  and g1130 (n1163, \in2[112] , n1162);
  not g1131 (n_850, \in3[113] );
  and g1132 (n1164, \in2[113] , n_850);
  not g1133 (n_851, n1163);
  not g1134 (n_852, n1164);
  and g1135 (n1165, n_851, n_852);
  not g1136 (n_853, \in3[114] );
  and g1137 (n1166, \in2[114] , n_853);
  not g1138 (n_854, n1166);
  and g1139 (n1167, n1165, n_854);
  not g1140 (n_855, n1167);
  and g1141 (n1168, n658, n_855);
  not g1142 (n_856, n1161);
  not g1143 (n_857, n1168);
  and g1144 (n1169, n_856, n_857);
  not g1145 (n_858, n1160);
  and g1146 (n1170, n_858, n1169);
  not g1147 (n_859, \in2[116] );
  and g1148 (n1171, n_859, \in3[116] );
  not g1161 (n_867, \in2[123] );
  and g1162 (n1178, n_867, \in3[123] );
  not g1163 (n_870, \in2[122] );
  and g1164 (n1179, n_870, \in3[122] );
  not g1165 (n_872, n1178);
  not g1166 (n_873, n1179);
  and g1167 (n1180, n_872, n_873);
  not g1168 (n_875, \in2[121] );
  and g1169 (n1181, n_875, \in3[121] );
  not g1170 (n_878, \in2[120] );
  and g1171 (n1182, n_878, \in3[120] );
  not g1172 (n_880, n1181);
  not g1178 (n_883, \in3[123] );
  and g1179 (n1186, \in2[123] , n_883);
  not g1180 (n_884, \in3[120] );
  and g1181 (n1187, \in2[120] , n_884);
  and g1182 (n1188, n_880, n1187);
  not g1183 (n_885, \in3[121] );
  and g1184 (n1189, \in2[121] , n_885);
  not g1185 (n_886, n1188);
  not g1186 (n_887, n1189);
  and g1187 (n1190, n_886, n_887);
  not g1188 (n_888, \in3[122] );
  and g1189 (n1191, \in2[122] , n_888);
  not g1190 (n_889, n1191);
  and g1191 (n1192, n1190, n_889);
  not g1192 (n_890, n1192);
  and g1193 (n1193, n1180, n_890);
  not g1194 (n_891, n1186);
  not g1195 (n_892, n1193);
  and g1196 (n1194, n_891, n_892);
  not g1197 (n_893, n1185);
  and g1198 (n1195, n_893, n1194);
  not g1199 (n_895, \in2[124] );
  and g1200 (n1196, n_895, \in3[124] );
  not g1201 (n_899, \in3[127] );
  and g1202 (n1197, \in2[127] , n_899);
  not g1203 (n_901, \in2[126] );
  and g1204 (n1198, n_901, \in3[126] );
  not g1205 (n_904, \in2[125] );
  and g1206 (n1199, n_904, \in3[125] );
  not g1207 (n_906, n1198);
  not g1208 (n_907, n1199);
  and g1209 (n1200, n_906, n_907);
  not g1210 (n_908, n1197);
  not g1216 (n_911, \in3[124] );
  and g1217 (n1204, \in2[124] , n_911);
  not g1218 (n_912, \in3[125] );
  and g1219 (n1205, \in2[125] , n_912);
  not g1220 (n_913, n1204);
  not g1221 (n_914, n1205);
  and g1222 (n1206, n_913, n_914);
  not g1223 (n_915, n1206);
  and g1224 (n1207, n1200, n_915);
  not g1225 (n_916, \in3[126] );
  and g1226 (n1208, \in2[126] , n_916);
  not g1227 (n_917, n1207);
  not g1228 (n_918, n1208);
  and g1229 (n1209, n_917, n_918);
  not g1230 (n_919, n1209);
  and g1231 (n1210, n_908, n_919);
  not g1232 (n_920, n1203);
  not g1233 (n_921, n1210);
  and g1234 (n1211, n_920, n_921);
  and g1235 (n1212, n_899, n1211);
  not g1236 (n_922, n1212);
  and g1237 (n1213, \in2[127] , n_922);
  not g1238 (n_925, \in1[119] );
  and g1239 (n1214, \in0[119] , n_925);
  not g1240 (n_926, \in0[119] );
  and g1241 (n1215, n_926, \in1[119] );
  not g1242 (n_928, \in0[118] );
  and g1243 (n1216, n_928, \in1[118] );
  not g1244 (n_930, n1215);
  not g1245 (n_931, n1216);
  and g1246 (n1217, n_930, n_931);
  not g1247 (n_933, \in0[117] );
  and g1248 (n1218, n_933, \in1[117] );
  not g1249 (n_937, \in1[116] );
  and g1250 (n1219, \in0[116] , n_937);
  not g1251 (n_938, n1218);
  and g1252 (n1220, n_938, n1219);
  not g1253 (n_939, \in1[117] );
  and g1254 (n1221, \in0[117] , n_939);
  not g1255 (n_940, n1220);
  not g1256 (n_941, n1221);
  and g1257 (n1222, n_940, n_941);
  not g1258 (n_942, n1222);
  and g1259 (n1223, n1217, n_942);
  not g1260 (n_943, \in1[118] );
  and g1261 (n1224, n_943, n_930);
  and g1262 (n1225, \in0[118] , n1224);
  not g1263 (n_945, \in0[112] );
  and g1264 (n1226, n_945, \in1[112] );
  not g1265 (n_948, \in0[115] );
  and g1266 (n1227, n_948, \in1[115] );
  not g1267 (n_951, \in0[114] );
  and g1268 (n1228, n_951, \in1[114] );
  not g1269 (n_953, n1227);
  not g1270 (n_954, n1228);
  and g1271 (n1229, n_953, n_954);
  not g1272 (n_956, \in0[113] );
  and g1273 (n1230, n_956, \in1[113] );
  not g1274 (n_960, \in1[111] );
  and g1275 (n1231, \in0[111] , n_960);
  not g1276 (n_961, \in0[111] );
  and g1277 (n1232, n_961, \in1[111] );
  not g1278 (n_963, \in0[110] );
  and g1279 (n1233, n_963, \in1[110] );
  not g1280 (n_965, n1232);
  not g1281 (n_966, n1233);
  and g1282 (n1234, n_965, n_966);
  not g1283 (n_968, \in0[109] );
  and g1284 (n1235, n_968, \in1[109] );
  not g1285 (n_972, \in1[108] );
  and g1286 (n1236, \in0[108] , n_972);
  not g1287 (n_973, n1235);
  and g1288 (n1237, n_973, n1236);
  not g1289 (n_974, \in1[109] );
  and g1290 (n1238, \in0[109] , n_974);
  not g1291 (n_975, n1237);
  not g1292 (n_976, n1238);
  and g1293 (n1239, n_975, n_976);
  not g1294 (n_977, n1239);
  and g1295 (n1240, n1234, n_977);
  not g1296 (n_978, \in1[110] );
  and g1297 (n1241, n_978, n_965);
  and g1298 (n1242, \in0[110] , n1241);
  not g1299 (n_981, \in1[103] );
  and g1300 (n1243, \in0[103] , n_981);
  not g1301 (n_982, \in0[103] );
  and g1302 (n1244, n_982, \in1[103] );
  not g1303 (n_984, \in0[102] );
  and g1304 (n1245, n_984, \in1[102] );
  not g1305 (n_986, n1244);
  not g1306 (n_987, n1245);
  and g1307 (n1246, n_986, n_987);
  not g1308 (n_989, \in0[101] );
  and g1309 (n1247, n_989, \in1[101] );
  not g1310 (n_993, \in1[100] );
  and g1311 (n1248, \in0[100] , n_993);
  not g1312 (n_994, n1247);
  and g1313 (n1249, n_994, n1248);
  not g1314 (n_995, \in1[101] );
  and g1315 (n1250, \in0[101] , n_995);
  not g1316 (n_996, n1249);
  not g1317 (n_997, n1250);
  and g1318 (n1251, n_996, n_997);
  not g1319 (n_998, n1251);
  and g1320 (n1252, n1246, n_998);
  not g1321 (n_999, \in1[102] );
  and g1322 (n1253, n_999, n_986);
  and g1323 (n1254, \in0[102] , n1253);
  not g1324 (n_1001, \in0[96] );
  and g1325 (n1255, n_1001, \in1[96] );
  not g1326 (n_1004, \in0[99] );
  and g1327 (n1256, n_1004, \in1[99] );
  not g1328 (n_1007, \in0[98] );
  and g1329 (n1257, n_1007, \in1[98] );
  not g1330 (n_1009, n1256);
  not g1331 (n_1010, n1257);
  and g1332 (n1258, n_1009, n_1010);
  not g1333 (n_1012, \in0[97] );
  and g1334 (n1259, n_1012, \in1[97] );
  not g1335 (n_1016, \in1[95] );
  and g1336 (n1260, \in0[95] , n_1016);
  not g1337 (n_1017, \in0[95] );
  and g1338 (n1261, n_1017, \in1[95] );
  not g1339 (n_1019, \in0[94] );
  and g1340 (n1262, n_1019, \in1[94] );
  not g1341 (n_1021, n1261);
  not g1342 (n_1022, n1262);
  and g1343 (n1263, n_1021, n_1022);
  not g1344 (n_1024, \in0[93] );
  and g1345 (n1264, n_1024, \in1[93] );
  not g1346 (n_1028, \in1[92] );
  and g1347 (n1265, \in0[92] , n_1028);
  not g1348 (n_1029, n1264);
  and g1349 (n1266, n_1029, n1265);
  not g1350 (n_1030, \in1[93] );
  and g1351 (n1267, \in0[93] , n_1030);
  not g1352 (n_1031, n1266);
  not g1353 (n_1032, n1267);
  and g1354 (n1268, n_1031, n_1032);
  not g1355 (n_1033, n1268);
  and g1356 (n1269, n1263, n_1033);
  not g1357 (n_1034, \in1[94] );
  and g1358 (n1270, n_1034, n_1021);
  and g1359 (n1271, \in0[94] , n1270);
  not g1360 (n_1037, \in1[87] );
  and g1361 (n1272, \in0[87] , n_1037);
  not g1362 (n_1038, \in0[87] );
  and g1363 (n1273, n_1038, \in1[87] );
  not g1364 (n_1040, \in0[86] );
  and g1365 (n1274, n_1040, \in1[86] );
  not g1366 (n_1042, n1273);
  not g1367 (n_1043, n1274);
  and g1368 (n1275, n_1042, n_1043);
  not g1369 (n_1045, \in0[85] );
  and g1370 (n1276, n_1045, \in1[85] );
  not g1371 (n_1049, \in1[84] );
  and g1372 (n1277, \in0[84] , n_1049);
  not g1373 (n_1050, n1276);
  and g1374 (n1278, n_1050, n1277);
  not g1375 (n_1051, \in1[85] );
  and g1376 (n1279, \in0[85] , n_1051);
  not g1377 (n_1052, n1278);
  not g1378 (n_1053, n1279);
  and g1379 (n1280, n_1052, n_1053);
  not g1380 (n_1054, n1280);
  and g1381 (n1281, n1275, n_1054);
  not g1382 (n_1055, \in1[86] );
  and g1383 (n1282, n_1055, n_1042);
  and g1384 (n1283, \in0[86] , n1282);
  not g1385 (n_1057, \in0[80] );
  and g1386 (n1284, n_1057, \in1[80] );
  not g1387 (n_1060, \in0[83] );
  and g1388 (n1285, n_1060, \in1[83] );
  not g1389 (n_1063, \in0[82] );
  and g1390 (n1286, n_1063, \in1[82] );
  not g1391 (n_1065, n1285);
  not g1392 (n_1066, n1286);
  and g1393 (n1287, n_1065, n_1066);
  not g1394 (n_1068, \in0[81] );
  and g1395 (n1288, n_1068, \in1[81] );
  not g1396 (n_1072, \in1[79] );
  and g1397 (n1289, \in0[79] , n_1072);
  not g1398 (n_1073, \in0[79] );
  and g1399 (n1290, n_1073, \in1[79] );
  not g1400 (n_1075, \in0[78] );
  and g1401 (n1291, n_1075, \in1[78] );
  not g1402 (n_1077, n1290);
  not g1403 (n_1078, n1291);
  and g1404 (n1292, n_1077, n_1078);
  not g1405 (n_1080, \in0[77] );
  and g1406 (n1293, n_1080, \in1[77] );
  not g1407 (n_1084, \in1[76] );
  and g1408 (n1294, \in0[76] , n_1084);
  not g1409 (n_1085, n1293);
  and g1410 (n1295, n_1085, n1294);
  not g1411 (n_1086, \in1[77] );
  and g1412 (n1296, \in0[77] , n_1086);
  not g1413 (n_1087, n1295);
  not g1414 (n_1088, n1296);
  and g1415 (n1297, n_1087, n_1088);
  not g1416 (n_1089, n1297);
  and g1417 (n1298, n1292, n_1089);
  not g1418 (n_1090, \in1[78] );
  and g1419 (n1299, n_1090, n_1077);
  and g1420 (n1300, \in0[78] , n1299);
  not g1421 (n_1093, \in1[71] );
  and g1422 (n1301, \in0[71] , n_1093);
  not g1423 (n_1094, \in0[71] );
  and g1424 (n1302, n_1094, \in1[71] );
  not g1425 (n_1096, \in0[70] );
  and g1426 (n1303, n_1096, \in1[70] );
  not g1427 (n_1098, n1302);
  not g1428 (n_1099, n1303);
  and g1429 (n1304, n_1098, n_1099);
  not g1430 (n_1101, \in0[69] );
  and g1431 (n1305, n_1101, \in1[69] );
  not g1432 (n_1105, \in1[68] );
  and g1433 (n1306, \in0[68] , n_1105);
  not g1434 (n_1106, n1305);
  and g1435 (n1307, n_1106, n1306);
  not g1436 (n_1107, \in1[69] );
  and g1437 (n1308, \in0[69] , n_1107);
  not g1438 (n_1108, n1307);
  not g1439 (n_1109, n1308);
  and g1440 (n1309, n_1108, n_1109);
  not g1441 (n_1110, n1309);
  and g1442 (n1310, n1304, n_1110);
  not g1443 (n_1111, \in1[70] );
  and g1444 (n1311, n_1111, n_1098);
  and g1445 (n1312, \in0[70] , n1311);
  not g1446 (n_1113, \in0[67] );
  and g1447 (n1313, n_1113, \in1[67] );
  not g1448 (n_1116, \in0[66] );
  and g1449 (n1314, n_1116, \in1[66] );
  not g1450 (n_1118, n1313);
  not g1451 (n_1119, n1314);
  and g1452 (n1315, n_1118, n_1119);
  not g1453 (n_1121, \in0[65] );
  and g1454 (n1316, n_1121, \in1[65] );
  not g1455 (n_1125, \in1[63] );
  and g1456 (n1317, \in0[63] , n_1125);
  not g1457 (n_1126, \in0[63] );
  and g1458 (n1318, n_1126, \in1[63] );
  not g1459 (n_1128, \in0[62] );
  and g1460 (n1319, n_1128, \in1[62] );
  not g1461 (n_1130, n1318);
  not g1462 (n_1131, n1319);
  and g1463 (n1320, n_1130, n_1131);
  not g1464 (n_1133, \in0[60] );
  and g1465 (n1321, n_1133, \in1[60] );
  not g1466 (n_1136, \in0[61] );
  and g1467 (n1322, n_1136, \in1[61] );
  not g1468 (n_1138, n1321);
  not g1469 (n_1139, n1322);
  and g1470 (n1323, n_1138, n_1139);
  and g1471 (n1324, n1320, n1323);
  not g1472 (n_1142, \in1[59] );
  and g1473 (n1325, \in0[59] , n_1142);
  not g1474 (n_1143, \in0[59] );
  and g1475 (n1326, n_1143, \in1[59] );
  not g1476 (n_1145, \in0[58] );
  and g1477 (n1327, n_1145, \in1[58] );
  not g1478 (n_1147, n1326);
  not g1479 (n_1148, n1327);
  and g1480 (n1328, n_1147, n_1148);
  not g1481 (n_1150, \in0[57] );
  and g1482 (n1329, n_1150, \in1[57] );
  not g1483 (n_1154, \in1[56] );
  and g1484 (n1330, \in0[56] , n_1154);
  not g1485 (n_1155, n1329);
  and g1486 (n1331, n_1155, n1330);
  not g1487 (n_1156, \in1[57] );
  and g1488 (n1332, \in0[57] , n_1156);
  not g1489 (n_1157, n1331);
  not g1490 (n_1158, n1332);
  and g1491 (n1333, n_1157, n_1158);
  not g1492 (n_1159, \in1[58] );
  and g1493 (n1334, \in0[58] , n_1159);
  not g1494 (n_1160, n1334);
  and g1495 (n1335, n1333, n_1160);
  not g1496 (n_1161, n1335);
  and g1497 (n1336, n1328, n_1161);
  not g1498 (n_1162, n1325);
  not g1499 (n_1163, n1336);
  and g1500 (n1337, n_1162, n_1163);
  not g1501 (n_1164, n1337);
  and g1502 (n1338, n1324, n_1164);
  not g1503 (n_1165, \in1[60] );
  and g1504 (n1339, \in0[60] , n_1165);
  and g1505 (n1340, n_1139, n1339);
  not g1506 (n_1166, \in1[61] );
  and g1507 (n1341, \in0[61] , n_1166);
  not g1508 (n_1167, n1340);
  not g1509 (n_1168, n1341);
  and g1510 (n1342, n_1167, n_1168);
  not g1511 (n_1169, n1342);
  and g1512 (n1343, n1320, n_1169);
  not g1513 (n_1170, \in1[62] );
  and g1514 (n1344, n_1170, n_1130);
  and g1515 (n1345, \in0[62] , n1344);
  not g1516 (n_1173, \in1[47] );
  and g1517 (n1346, \in0[47] , n_1173);
  not g1518 (n_1174, \in0[47] );
  and g1519 (n1347, n_1174, \in1[47] );
  not g1520 (n_1176, \in0[46] );
  and g1521 (n1348, n_1176, \in1[46] );
  not g1522 (n_1178, n1347);
  not g1523 (n_1179, n1348);
  and g1524 (n1349, n_1178, n_1179);
  not g1525 (n_1181, \in0[44] );
  and g1526 (n1350, n_1181, \in1[44] );
  not g1527 (n_1184, \in0[45] );
  and g1528 (n1351, n_1184, \in1[45] );
  not g1529 (n_1186, n1350);
  not g1530 (n_1187, n1351);
  and g1531 (n1352, n_1186, n_1187);
  and g1532 (n1353, n1349, n1352);
  not g1533 (n_1190, \in1[43] );
  and g1534 (n1354, \in0[43] , n_1190);
  not g1535 (n_1191, \in0[43] );
  and g1536 (n1355, n_1191, \in1[43] );
  not g1537 (n_1193, \in0[42] );
  and g1538 (n1356, n_1193, \in1[42] );
  not g1539 (n_1195, n1355);
  not g1540 (n_1196, n1356);
  and g1541 (n1357, n_1195, n_1196);
  not g1542 (n_1198, \in0[41] );
  and g1543 (n1358, n_1198, \in1[41] );
  not g1544 (n_1202, \in1[40] );
  and g1545 (n1359, \in0[40] , n_1202);
  not g1546 (n_1203, n1358);
  and g1547 (n1360, n_1203, n1359);
  not g1548 (n_1204, \in1[41] );
  and g1549 (n1361, \in0[41] , n_1204);
  not g1550 (n_1205, n1360);
  not g1551 (n_1206, n1361);
  and g1552 (n1362, n_1205, n_1206);
  not g1553 (n_1207, \in1[42] );
  and g1554 (n1363, \in0[42] , n_1207);
  not g1555 (n_1208, n1363);
  and g1556 (n1364, n1362, n_1208);
  not g1557 (n_1209, n1364);
  and g1558 (n1365, n1357, n_1209);
  not g1559 (n_1210, n1354);
  not g1560 (n_1211, n1365);
  and g1561 (n1366, n_1210, n_1211);
  not g1562 (n_1212, n1366);
  and g1563 (n1367, n1353, n_1212);
  not g1564 (n_1213, \in1[44] );
  and g1565 (n1368, \in0[44] , n_1213);
  and g1566 (n1369, n_1187, n1368);
  not g1567 (n_1214, \in1[45] );
  and g1568 (n1370, \in0[45] , n_1214);
  not g1569 (n_1215, n1369);
  not g1570 (n_1216, n1370);
  and g1571 (n1371, n_1215, n_1216);
  not g1572 (n_1217, n1371);
  and g1573 (n1372, n1349, n_1217);
  not g1574 (n_1218, \in1[46] );
  and g1575 (n1373, n_1218, n_1178);
  and g1576 (n1374, \in0[46] , n1373);
  not g1577 (n_1220, \in0[32] );
  and g1578 (n1375, n_1220, \in1[32] );
  not g1579 (n_1223, \in0[31] );
  and g1580 (n1376, n_1223, \in1[31] );
  not g1581 (n_1226, \in0[30] );
  and g1582 (n1377, n_1226, \in1[30] );
  not g1583 (n_1229, \in0[29] );
  and g1584 (n1378, n_1229, \in1[29] );
  not g1585 (n_1232, \in0[28] );
  and g1586 (n1379, n_1232, \in1[28] );
  not g1587 (n_1235, \in0[27] );
  and g1588 (n1380, n_1235, \in1[27] );
  not g1589 (n_1238, \in0[26] );
  and g1590 (n1381, n_1238, \in1[26] );
  not g1591 (n_1241, \in0[23] );
  and g1592 (n1382, n_1241, \in1[23] );
  not g1593 (n_1244, \in0[22] );
  and g1594 (n1383, n_1244, \in1[22] );
  not g1595 (n_1247, \in0[21] );
  and g1596 (n1384, n_1247, \in1[21] );
  not g1597 (n_1250, \in0[20] );
  and g1598 (n1385, n_1250, \in1[20] );
  not g1599 (n_1253, \in0[19] );
  and g1600 (n1386, n_1253, \in1[19] );
  not g1601 (n_1256, \in0[18] );
  and g1602 (n1387, n_1256, \in1[18] );
  not g1603 (n_1259, \in0[15] );
  and g1604 (n1388, n_1259, \in1[15] );
  not g1605 (n_1262, \in0[14] );
  and g1606 (n1389, n_1262, \in1[14] );
  not g1607 (n_1265, \in0[13] );
  and g1608 (n1390, n_1265, \in1[13] );
  not g1609 (n_1268, \in0[12] );
  and g1610 (n1391, n_1268, \in1[12] );
  not g1611 (n_1271, \in0[11] );
  and g1612 (n1392, n_1271, \in1[11] );
  not g1613 (n_1274, \in0[10] );
  and g1614 (n1393, n_1274, \in1[10] );
  not g1615 (n_1277, \in0[7] );
  and g1616 (n1394, n_1277, \in1[7] );
  not g1617 (n_1280, \in0[6] );
  and g1618 (n1395, n_1280, \in1[6] );
  not g1619 (n_1283, \in0[3] );
  and g1620 (n1396, n_1283, \in1[3] );
  not g1621 (n_1287, \in1[0] );
  and g1622 (n1397, \in0[0] , n_1287);
  not g1623 (n_1290, \in1[1] );
  and g1624 (n1398, \in0[1] , n_1290);
  not g1625 (n_1291, n1397);
  not g1626 (n_1292, n1398);
  and g1627 (n1399, n_1291, n_1292);
  not g1628 (n_1294, \in0[2] );
  and g1629 (n1400, n_1294, \in1[2] );
  not g1630 (n_1296, \in0[1] );
  and g1631 (n1401, n_1296, \in1[1] );
  not g1632 (n_1297, n1400);
  not g1633 (n_1298, n1401);
  and g1634 (n1402, n_1297, n_1298);
  not g1635 (n_1299, n1399);
  and g1636 (n1403, n_1299, n1402);
  not g1637 (n_1300, \in1[2] );
  and g1638 (n1404, \in0[2] , n_1300);
  not g1639 (n_1301, n1403);
  not g1640 (n_1302, n1404);
  and g1641 (n1405, n_1301, n_1302);
  not g1642 (n_1303, n1396);
  not g1643 (n_1304, n1405);
  and g1644 (n1406, n_1303, n_1304);
  not g1645 (n_1305, \in1[3] );
  and g1646 (n1407, \in0[3] , n_1305);
  not g1647 (n_1306, n1406);
  not g1648 (n_1307, n1407);
  and g1649 (n1408, n_1306, n_1307);
  not g1650 (n_1309, \in0[4] );
  and g1651 (n1409, n_1309, n1408);
  not g1652 (n_1311, \in1[4] );
  not g1653 (n_1312, n1409);
  and g1654 (n1410, n_1311, n_1312);
  not g1655 (n_1313, n1408);
  and g1656 (n1411, \in0[4] , n_1313);
  not g1657 (n_1314, n1410);
  not g1658 (n_1315, n1411);
  and g1659 (n1412, n_1314, n_1315);
  not g1660 (n_1317, \in0[5] );
  and g1661 (n1413, n_1317, n1412);
  not g1662 (n_1319, \in1[5] );
  not g1663 (n_1320, n1413);
  and g1664 (n1414, n_1319, n_1320);
  not g1665 (n_1321, n1412);
  and g1666 (n1415, \in0[5] , n_1321);
  not g1667 (n_1322, n1414);
  not g1668 (n_1323, n1415);
  and g1669 (n1416, n_1322, n_1323);
  not g1670 (n_1324, n1395);
  not g1671 (n_1325, n1416);
  and g1672 (n1417, n_1324, n_1325);
  not g1673 (n_1326, \in1[6] );
  and g1674 (n1418, \in0[6] , n_1326);
  not g1675 (n_1327, n1417);
  not g1676 (n_1328, n1418);
  and g1677 (n1419, n_1327, n_1328);
  not g1678 (n_1329, n1394);
  not g1679 (n_1330, n1419);
  and g1680 (n1420, n_1329, n_1330);
  not g1681 (n_1331, \in1[7] );
  and g1682 (n1421, \in0[7] , n_1331);
  not g1683 (n_1332, n1420);
  not g1684 (n_1333, n1421);
  and g1685 (n1422, n_1332, n_1333);
  not g1686 (n_1335, \in0[8] );
  and g1687 (n1423, n_1335, n1422);
  not g1688 (n_1337, \in1[8] );
  not g1689 (n_1338, n1423);
  and g1690 (n1424, n_1337, n_1338);
  not g1691 (n_1339, n1422);
  and g1692 (n1425, \in0[8] , n_1339);
  not g1693 (n_1340, n1424);
  not g1694 (n_1341, n1425);
  and g1695 (n1426, n_1340, n_1341);
  not g1696 (n_1343, \in0[9] );
  and g1697 (n1427, n_1343, n1426);
  not g1698 (n_1345, \in1[9] );
  not g1699 (n_1346, n1427);
  and g1700 (n1428, n_1345, n_1346);
  not g1701 (n_1347, n1426);
  and g1702 (n1429, \in0[9] , n_1347);
  not g1703 (n_1348, n1428);
  not g1704 (n_1349, n1429);
  and g1705 (n1430, n_1348, n_1349);
  not g1706 (n_1350, n1393);
  not g1707 (n_1351, n1430);
  and g1708 (n1431, n_1350, n_1351);
  not g1709 (n_1352, \in1[10] );
  and g1710 (n1432, \in0[10] , n_1352);
  not g1711 (n_1353, n1431);
  not g1712 (n_1354, n1432);
  and g1713 (n1433, n_1353, n_1354);
  not g1714 (n_1355, n1392);
  not g1715 (n_1356, n1433);
  and g1716 (n1434, n_1355, n_1356);
  not g1717 (n_1357, \in1[11] );
  and g1718 (n1435, \in0[11] , n_1357);
  not g1719 (n_1358, n1434);
  not g1720 (n_1359, n1435);
  and g1721 (n1436, n_1358, n_1359);
  not g1722 (n_1360, n1391);
  not g1723 (n_1361, n1436);
  and g1724 (n1437, n_1360, n_1361);
  not g1725 (n_1362, \in1[12] );
  and g1726 (n1438, \in0[12] , n_1362);
  not g1727 (n_1363, n1437);
  not g1728 (n_1364, n1438);
  and g1729 (n1439, n_1363, n_1364);
  not g1730 (n_1365, n1390);
  not g1731 (n_1366, n1439);
  and g1732 (n1440, n_1365, n_1366);
  not g1733 (n_1367, \in1[13] );
  and g1734 (n1441, \in0[13] , n_1367);
  not g1735 (n_1368, n1440);
  not g1736 (n_1369, n1441);
  and g1737 (n1442, n_1368, n_1369);
  not g1738 (n_1370, n1389);
  not g1739 (n_1371, n1442);
  and g1740 (n1443, n_1370, n_1371);
  not g1741 (n_1372, \in1[14] );
  and g1742 (n1444, \in0[14] , n_1372);
  not g1743 (n_1373, n1443);
  not g1744 (n_1374, n1444);
  and g1745 (n1445, n_1373, n_1374);
  not g1746 (n_1375, n1388);
  not g1747 (n_1376, n1445);
  and g1748 (n1446, n_1375, n_1376);
  not g1749 (n_1377, \in1[15] );
  and g1750 (n1447, \in0[15] , n_1377);
  not g1751 (n_1378, n1446);
  not g1752 (n_1379, n1447);
  and g1753 (n1448, n_1378, n_1379);
  not g1754 (n_1381, \in0[16] );
  and g1755 (n1449, n_1381, n1448);
  not g1756 (n_1383, \in1[16] );
  not g1757 (n_1384, n1449);
  and g1758 (n1450, n_1383, n_1384);
  not g1759 (n_1385, n1448);
  and g1760 (n1451, \in0[16] , n_1385);
  not g1761 (n_1386, n1450);
  not g1762 (n_1387, n1451);
  and g1763 (n1452, n_1386, n_1387);
  not g1764 (n_1389, \in0[17] );
  and g1765 (n1453, n_1389, n1452);
  not g1766 (n_1391, \in1[17] );
  not g1767 (n_1392, n1453);
  and g1768 (n1454, n_1391, n_1392);
  not g1769 (n_1393, n1452);
  and g1770 (n1455, \in0[17] , n_1393);
  not g1771 (n_1394, n1454);
  not g1772 (n_1395, n1455);
  and g1773 (n1456, n_1394, n_1395);
  not g1774 (n_1396, n1387);
  not g1775 (n_1397, n1456);
  and g1776 (n1457, n_1396, n_1397);
  not g1777 (n_1398, \in1[18] );
  and g1778 (n1458, \in0[18] , n_1398);
  not g1779 (n_1399, n1457);
  not g1780 (n_1400, n1458);
  and g1781 (n1459, n_1399, n_1400);
  not g1782 (n_1401, n1386);
  not g1783 (n_1402, n1459);
  and g1784 (n1460, n_1401, n_1402);
  not g1785 (n_1403, \in1[19] );
  and g1786 (n1461, \in0[19] , n_1403);
  not g1787 (n_1404, n1460);
  not g1788 (n_1405, n1461);
  and g1789 (n1462, n_1404, n_1405);
  not g1790 (n_1406, n1385);
  not g1791 (n_1407, n1462);
  and g1792 (n1463, n_1406, n_1407);
  not g1793 (n_1408, \in1[20] );
  and g1794 (n1464, \in0[20] , n_1408);
  not g1795 (n_1409, n1463);
  not g1796 (n_1410, n1464);
  and g1797 (n1465, n_1409, n_1410);
  not g1798 (n_1411, n1384);
  not g1799 (n_1412, n1465);
  and g1800 (n1466, n_1411, n_1412);
  not g1801 (n_1413, \in1[21] );
  and g1802 (n1467, \in0[21] , n_1413);
  not g1803 (n_1414, n1466);
  not g1804 (n_1415, n1467);
  and g1805 (n1468, n_1414, n_1415);
  not g1806 (n_1416, n1383);
  not g1807 (n_1417, n1468);
  and g1808 (n1469, n_1416, n_1417);
  not g1809 (n_1418, \in1[22] );
  and g1810 (n1470, \in0[22] , n_1418);
  not g1811 (n_1419, n1469);
  not g1812 (n_1420, n1470);
  and g1813 (n1471, n_1419, n_1420);
  not g1814 (n_1421, n1382);
  not g1815 (n_1422, n1471);
  and g1816 (n1472, n_1421, n_1422);
  not g1817 (n_1423, \in1[23] );
  and g1818 (n1473, \in0[23] , n_1423);
  not g1819 (n_1424, n1472);
  not g1820 (n_1425, n1473);
  and g1821 (n1474, n_1424, n_1425);
  not g1822 (n_1427, \in0[24] );
  and g1823 (n1475, n_1427, n1474);
  not g1824 (n_1429, \in1[24] );
  not g1825 (n_1430, n1475);
  and g1826 (n1476, n_1429, n_1430);
  not g1827 (n_1431, n1474);
  and g1828 (n1477, \in0[24] , n_1431);
  not g1829 (n_1432, n1476);
  not g1830 (n_1433, n1477);
  and g1831 (n1478, n_1432, n_1433);
  not g1832 (n_1435, \in0[25] );
  and g1833 (n1479, n_1435, n1478);
  not g1834 (n_1437, \in1[25] );
  not g1835 (n_1438, n1479);
  and g1836 (n1480, n_1437, n_1438);
  not g1837 (n_1439, n1478);
  and g1838 (n1481, \in0[25] , n_1439);
  not g1839 (n_1440, n1480);
  not g1840 (n_1441, n1481);
  and g1841 (n1482, n_1440, n_1441);
  not g1842 (n_1442, n1381);
  not g1843 (n_1443, n1482);
  and g1844 (n1483, n_1442, n_1443);
  not g1845 (n_1444, \in1[26] );
  and g1846 (n1484, \in0[26] , n_1444);
  not g1847 (n_1445, n1483);
  not g1848 (n_1446, n1484);
  and g1849 (n1485, n_1445, n_1446);
  not g1850 (n_1447, n1380);
  not g1851 (n_1448, n1485);
  and g1852 (n1486, n_1447, n_1448);
  not g1853 (n_1449, \in1[27] );
  and g1854 (n1487, \in0[27] , n_1449);
  not g1855 (n_1450, n1486);
  not g1856 (n_1451, n1487);
  and g1857 (n1488, n_1450, n_1451);
  not g1858 (n_1452, n1379);
  not g1859 (n_1453, n1488);
  and g1860 (n1489, n_1452, n_1453);
  not g1861 (n_1454, \in1[28] );
  and g1862 (n1490, \in0[28] , n_1454);
  not g1863 (n_1455, n1489);
  not g1864 (n_1456, n1490);
  and g1865 (n1491, n_1455, n_1456);
  not g1866 (n_1457, n1378);
  not g1867 (n_1458, n1491);
  and g1868 (n1492, n_1457, n_1458);
  not g1869 (n_1459, \in1[29] );
  and g1870 (n1493, \in0[29] , n_1459);
  not g1871 (n_1460, n1492);
  not g1872 (n_1461, n1493);
  and g1873 (n1494, n_1460, n_1461);
  not g1874 (n_1462, n1377);
  not g1875 (n_1463, n1494);
  and g1876 (n1495, n_1462, n_1463);
  not g1877 (n_1464, \in1[30] );
  and g1878 (n1496, \in0[30] , n_1464);
  not g1879 (n_1465, n1495);
  not g1880 (n_1466, n1496);
  and g1881 (n1497, n_1465, n_1466);
  not g1882 (n_1467, n1376);
  not g1883 (n_1468, n1497);
  and g1884 (n1498, n_1467, n_1468);
  not g1885 (n_1469, \in1[31] );
  and g1886 (n1499, \in0[31] , n_1469);
  not g1887 (n_1470, n1498);
  not g1888 (n_1471, n1499);
  and g1889 (n1500, n_1470, n_1471);
  not g1890 (n_1473, \in0[39] );
  and g1891 (n1501, n_1473, \in1[39] );
  not g1892 (n_1476, \in0[38] );
  and g1893 (n1502, n_1476, \in1[38] );
  not g1894 (n_1478, n1501);
  not g1895 (n_1479, n1502);
  and g1896 (n1503, n_1478, n_1479);
  not g1897 (n_1481, \in0[36] );
  and g1898 (n1504, n_1481, \in1[36] );
  not g1899 (n_1484, \in0[37] );
  and g1900 (n1505, n_1484, \in1[37] );
  not g1901 (n_1486, n1504);
  not g1902 (n_1487, n1505);
  and g1903 (n1506, n_1486, n_1487);
  and g1904 (n1507, n1503, n1506);
  not g1905 (n_1489, \in0[33] );
  and g1906 (n1508, n_1489, \in1[33] );
  not g1907 (n_1492, \in0[35] );
  and g1908 (n1509, n_1492, \in1[35] );
  not g1909 (n_1495, \in0[34] );
  and g1910 (n1510, n_1495, \in1[34] );
  not g1911 (n_1497, n1509);
  not g1912 (n_1498, n1510);
  and g1913 (n1511, n_1497, n_1498);
  not g1914 (n_1499, n1508);
  not g1921 (n_1502, \in1[39] );
  and g1922 (n1516, \in0[39] , n_1502);
  not g1923 (n_1503, \in1[36] );
  and g1924 (n1517, \in0[36] , n_1503);
  and g1925 (n1518, n_1487, n1517);
  not g1926 (n_1504, \in1[37] );
  and g1927 (n1519, \in0[37] , n_1504);
  not g1928 (n_1505, n1518);
  not g1929 (n_1506, n1519);
  and g1930 (n1520, n_1505, n_1506);
  not g1931 (n_1507, n1520);
  and g1932 (n1521, n1503, n_1507);
  not g1933 (n_1508, \in1[38] );
  and g1934 (n1522, n_1508, n_1478);
  and g1935 (n1523, \in0[38] , n1522);
  not g1936 (n_1509, \in1[35] );
  and g1937 (n1524, \in0[35] , n_1509);
  not g1938 (n_1510, \in1[32] );
  and g1939 (n1525, n_1510, n_1499);
  and g1940 (n1526, \in0[32] , n1525);
  not g1941 (n_1511, \in1[33] );
  and g1942 (n1527, \in0[33] , n_1511);
  not g1943 (n_1512, n1526);
  not g1944 (n_1513, n1527);
  and g1945 (n1528, n_1512, n_1513);
  not g1946 (n_1514, \in1[34] );
  and g1947 (n1529, \in0[34] , n_1514);
  not g1948 (n_1515, n1529);
  and g1949 (n1530, n1528, n_1515);
  not g1950 (n_1516, n1530);
  and g1951 (n1531, n1511, n_1516);
  not g1952 (n_1517, n1524);
  not g1953 (n_1518, n1531);
  and g1954 (n1532, n_1517, n_1518);
  not g1955 (n_1519, n1532);
  and g1956 (n1533, n1507, n_1519);
  not g1966 (n_1525, \in0[40] );
  and g1967 (n1538, n_1525, \in1[40] );
  not g1983 (n_1534, \in0[48] );
  and g1984 (n1547, n_1534, \in1[48] );
  not g1985 (n_1537, \in0[55] );
  and g1986 (n1548, n_1537, \in1[55] );
  not g1987 (n_1540, \in0[54] );
  and g1988 (n1549, n_1540, \in1[54] );
  not g1989 (n_1542, n1548);
  not g1990 (n_1543, n1549);
  and g1991 (n1550, n_1542, n_1543);
  not g1992 (n_1545, \in0[53] );
  and g1993 (n1551, n_1545, \in1[53] );
  not g1994 (n_1548, \in0[52] );
  and g1995 (n1552, n_1548, \in1[52] );
  not g1996 (n_1550, n1551);
  not g1997 (n_1551, n1552);
  and g1998 (n1553, n_1550, n_1551);
  and g1999 (n1554, n1550, n1553);
  not g2000 (n_1553, \in0[49] );
  and g2001 (n1555, n_1553, \in1[49] );
  not g2002 (n_1556, \in0[51] );
  and g2003 (n1556, n_1556, \in1[51] );
  not g2004 (n_1559, \in0[50] );
  and g2005 (n1557, n_1559, \in1[50] );
  not g2006 (n_1561, n1556);
  not g2007 (n_1562, n1557);
  and g2008 (n1558, n_1561, n_1562);
  not g2009 (n_1563, n1555);
  not g2016 (n_1566, \in1[55] );
  and g2017 (n1563, \in0[55] , n_1566);
  not g2018 (n_1567, \in1[51] );
  and g2019 (n1564, \in0[51] , n_1567);
  not g2020 (n_1568, \in1[48] );
  and g2021 (n1565, n_1568, n_1563);
  and g2022 (n1566, \in0[48] , n1565);
  not g2023 (n_1569, \in1[49] );
  and g2024 (n1567, \in0[49] , n_1569);
  not g2025 (n_1570, n1566);
  not g2026 (n_1571, n1567);
  and g2027 (n1568, n_1570, n_1571);
  not g2028 (n_1572, \in1[50] );
  and g2029 (n1569, \in0[50] , n_1572);
  not g2030 (n_1573, n1569);
  and g2031 (n1570, n1568, n_1573);
  not g2032 (n_1574, n1570);
  and g2033 (n1571, n1558, n_1574);
  not g2034 (n_1575, n1564);
  not g2035 (n_1576, n1571);
  and g2036 (n1572, n_1575, n_1576);
  not g2037 (n_1577, n1572);
  and g2038 (n1573, n1554, n_1577);
  not g2039 (n_1578, \in1[52] );
  and g2040 (n1574, \in0[52] , n_1578);
  and g2041 (n1575, n_1550, n1574);
  not g2042 (n_1579, \in1[53] );
  and g2043 (n1576, \in0[53] , n_1579);
  not g2044 (n_1580, n1575);
  not g2045 (n_1581, n1576);
  and g2046 (n1577, n_1580, n_1581);
  not g2047 (n_1582, \in1[54] );
  and g2048 (n1578, \in0[54] , n_1582);
  not g2049 (n_1583, n1578);
  and g2050 (n1579, n1577, n_1583);
  not g2051 (n_1584, n1579);
  and g2052 (n1580, n1550, n_1584);
  not g2060 (n_1589, \in0[56] );
  and g2061 (n1584, n_1589, \in1[56] );
  not g2077 (n_1598, \in0[64] );
  and g2078 (n1593, n_1598, \in1[64] );
  not g2082 (n_1602, n1316);
  not g2085 (n_1603, \in1[67] );
  and g2086 (n1597, \in0[67] , n_1603);
  not g2087 (n_1604, \in1[64] );
  and g2088 (n1598, \in0[64] , n_1604);
  and g2089 (n1599, n_1602, n1598);
  not g2090 (n_1605, \in1[65] );
  and g2091 (n1600, \in0[65] , n_1605);
  not g2092 (n_1606, n1599);
  not g2093 (n_1607, n1600);
  and g2094 (n1601, n_1606, n_1607);
  not g2095 (n_1608, \in1[66] );
  and g2096 (n1602, \in0[66] , n_1608);
  not g2097 (n_1609, n1602);
  and g2098 (n1603, n1601, n_1609);
  not g2099 (n_1610, n1603);
  and g2100 (n1604, n1315, n_1610);
  not g2101 (n_1611, n1597);
  not g2102 (n_1612, n1604);
  and g2103 (n1605, n_1611, n_1612);
  not g2104 (n_1613, n1596);
  and g2105 (n1606, n_1613, n1605);
  not g2106 (n_1614, \in0[68] );
  and g2107 (n1607, n_1614, \in1[68] );
  not g2120 (n_1622, \in0[75] );
  and g2121 (n1614, n_1622, \in1[75] );
  not g2122 (n_1625, \in0[74] );
  and g2123 (n1615, n_1625, \in1[74] );
  not g2124 (n_1627, n1614);
  not g2125 (n_1628, n1615);
  and g2126 (n1616, n_1627, n_1628);
  not g2127 (n_1630, \in0[73] );
  and g2128 (n1617, n_1630, \in1[73] );
  not g2129 (n_1633, \in0[72] );
  and g2130 (n1618, n_1633, \in1[72] );
  not g2131 (n_1635, n1617);
  not g2137 (n_1638, \in1[75] );
  and g2138 (n1622, \in0[75] , n_1638);
  not g2139 (n_1639, \in1[72] );
  and g2140 (n1623, \in0[72] , n_1639);
  and g2141 (n1624, n_1635, n1623);
  not g2142 (n_1640, \in1[73] );
  and g2143 (n1625, \in0[73] , n_1640);
  not g2144 (n_1641, n1624);
  not g2145 (n_1642, n1625);
  and g2146 (n1626, n_1641, n_1642);
  not g2147 (n_1643, \in1[74] );
  and g2148 (n1627, \in0[74] , n_1643);
  not g2149 (n_1644, n1627);
  and g2150 (n1628, n1626, n_1644);
  not g2151 (n_1645, n1628);
  and g2152 (n1629, n1616, n_1645);
  not g2153 (n_1646, n1622);
  not g2154 (n_1647, n1629);
  and g2155 (n1630, n_1646, n_1647);
  not g2156 (n_1648, n1621);
  and g2157 (n1631, n_1648, n1630);
  not g2158 (n_1649, \in0[76] );
  and g2159 (n1632, n_1649, \in1[76] );
  not g2172 (n_1656, n1288);
  not g2178 (n_1659, \in1[83] );
  and g2179 (n1642, \in0[83] , n_1659);
  not g2180 (n_1660, \in1[80] );
  and g2181 (n1643, n_1660, n_1656);
  and g2182 (n1644, \in0[80] , n1643);
  not g2183 (n_1661, \in1[81] );
  and g2184 (n1645, \in0[81] , n_1661);
  not g2185 (n_1662, n1644);
  not g2186 (n_1663, n1645);
  and g2187 (n1646, n_1662, n_1663);
  not g2188 (n_1664, \in1[82] );
  and g2189 (n1647, \in0[82] , n_1664);
  not g2190 (n_1665, n1647);
  and g2191 (n1648, n1646, n_1665);
  not g2192 (n_1666, n1648);
  and g2193 (n1649, n1287, n_1666);
  not g2194 (n_1667, n1642);
  not g2195 (n_1668, n1649);
  and g2196 (n1650, n_1667, n_1668);
  not g2197 (n_1669, n1641);
  and g2198 (n1651, n_1669, n1650);
  not g2199 (n_1670, \in0[84] );
  and g2200 (n1652, n_1670, \in1[84] );
  not g2213 (n_1678, \in0[91] );
  and g2214 (n1659, n_1678, \in1[91] );
  not g2215 (n_1681, \in0[90] );
  and g2216 (n1660, n_1681, \in1[90] );
  not g2217 (n_1683, n1659);
  not g2218 (n_1684, n1660);
  and g2219 (n1661, n_1683, n_1684);
  not g2220 (n_1686, \in0[89] );
  and g2221 (n1662, n_1686, \in1[89] );
  not g2222 (n_1689, \in0[88] );
  and g2223 (n1663, n_1689, \in1[88] );
  not g2224 (n_1691, n1662);
  not g2230 (n_1694, \in1[91] );
  and g2231 (n1667, \in0[91] , n_1694);
  not g2232 (n_1695, \in1[88] );
  and g2233 (n1668, \in0[88] , n_1695);
  and g2234 (n1669, n_1691, n1668);
  not g2235 (n_1696, \in1[89] );
  and g2236 (n1670, \in0[89] , n_1696);
  not g2237 (n_1697, n1669);
  not g2238 (n_1698, n1670);
  and g2239 (n1671, n_1697, n_1698);
  not g2240 (n_1699, \in1[90] );
  and g2241 (n1672, \in0[90] , n_1699);
  not g2242 (n_1700, n1672);
  and g2243 (n1673, n1671, n_1700);
  not g2244 (n_1701, n1673);
  and g2245 (n1674, n1661, n_1701);
  not g2246 (n_1702, n1667);
  not g2247 (n_1703, n1674);
  and g2248 (n1675, n_1702, n_1703);
  not g2249 (n_1704, n1666);
  and g2250 (n1676, n_1704, n1675);
  not g2251 (n_1705, \in0[92] );
  and g2252 (n1677, n_1705, \in1[92] );
  not g2265 (n_1712, n1259);
  not g2271 (n_1715, \in1[99] );
  and g2272 (n1687, \in0[99] , n_1715);
  not g2273 (n_1716, \in1[96] );
  and g2274 (n1688, n_1716, n_1712);
  and g2275 (n1689, \in0[96] , n1688);
  not g2276 (n_1717, \in1[97] );
  and g2277 (n1690, \in0[97] , n_1717);
  not g2278 (n_1718, n1689);
  not g2279 (n_1719, n1690);
  and g2280 (n1691, n_1718, n_1719);
  not g2281 (n_1720, \in1[98] );
  and g2282 (n1692, \in0[98] , n_1720);
  not g2283 (n_1721, n1692);
  and g2284 (n1693, n1691, n_1721);
  not g2285 (n_1722, n1693);
  and g2286 (n1694, n1258, n_1722);
  not g2287 (n_1723, n1687);
  not g2288 (n_1724, n1694);
  and g2289 (n1695, n_1723, n_1724);
  not g2290 (n_1725, n1686);
  and g2291 (n1696, n_1725, n1695);
  not g2292 (n_1726, \in0[100] );
  and g2293 (n1697, n_1726, \in1[100] );
  not g2306 (n_1734, \in0[107] );
  and g2307 (n1704, n_1734, \in1[107] );
  not g2308 (n_1737, \in0[106] );
  and g2309 (n1705, n_1737, \in1[106] );
  not g2310 (n_1739, n1704);
  not g2311 (n_1740, n1705);
  and g2312 (n1706, n_1739, n_1740);
  not g2313 (n_1742, \in0[105] );
  and g2314 (n1707, n_1742, \in1[105] );
  not g2315 (n_1745, \in0[104] );
  and g2316 (n1708, n_1745, \in1[104] );
  not g2317 (n_1747, n1707);
  not g2323 (n_1750, \in1[107] );
  and g2324 (n1712, \in0[107] , n_1750);
  not g2325 (n_1751, \in1[104] );
  and g2326 (n1713, \in0[104] , n_1751);
  and g2327 (n1714, n_1747, n1713);
  not g2328 (n_1752, \in1[105] );
  and g2329 (n1715, \in0[105] , n_1752);
  not g2330 (n_1753, n1714);
  not g2331 (n_1754, n1715);
  and g2332 (n1716, n_1753, n_1754);
  not g2333 (n_1755, \in1[106] );
  and g2334 (n1717, \in0[106] , n_1755);
  not g2335 (n_1756, n1717);
  and g2336 (n1718, n1716, n_1756);
  not g2337 (n_1757, n1718);
  and g2338 (n1719, n1706, n_1757);
  not g2339 (n_1758, n1712);
  not g2340 (n_1759, n1719);
  and g2341 (n1720, n_1758, n_1759);
  not g2342 (n_1760, n1711);
  and g2343 (n1721, n_1760, n1720);
  not g2344 (n_1761, \in0[108] );
  and g2345 (n1722, n_1761, \in1[108] );
  not g2358 (n_1768, n1230);
  not g2364 (n_1771, \in1[115] );
  and g2365 (n1732, \in0[115] , n_1771);
  not g2366 (n_1772, \in1[112] );
  and g2367 (n1733, n_1772, n_1768);
  and g2368 (n1734, \in0[112] , n1733);
  not g2369 (n_1773, \in1[113] );
  and g2370 (n1735, \in0[113] , n_1773);
  not g2371 (n_1774, n1734);
  not g2372 (n_1775, n1735);
  and g2373 (n1736, n_1774, n_1775);
  not g2374 (n_1776, \in1[114] );
  and g2375 (n1737, \in0[114] , n_1776);
  not g2376 (n_1777, n1737);
  and g2377 (n1738, n1736, n_1777);
  not g2378 (n_1778, n1738);
  and g2379 (n1739, n1229, n_1778);
  not g2380 (n_1779, n1732);
  not g2381 (n_1780, n1739);
  and g2382 (n1740, n_1779, n_1780);
  not g2383 (n_1781, n1731);
  and g2384 (n1741, n_1781, n1740);
  not g2385 (n_1782, \in0[116] );
  and g2386 (n1742, n_1782, \in1[116] );
  not g2399 (n_1790, \in0[123] );
  and g2400 (n1749, n_1790, \in1[123] );
  not g2401 (n_1793, \in0[122] );
  and g2402 (n1750, n_1793, \in1[122] );
  not g2403 (n_1795, n1749);
  not g2404 (n_1796, n1750);
  and g2405 (n1751, n_1795, n_1796);
  not g2406 (n_1798, \in0[121] );
  and g2407 (n1752, n_1798, \in1[121] );
  not g2408 (n_1801, \in0[120] );
  and g2409 (n1753, n_1801, \in1[120] );
  not g2410 (n_1803, n1752);
  not g2416 (n_1806, \in1[123] );
  and g2417 (n1757, \in0[123] , n_1806);
  not g2418 (n_1807, \in1[120] );
  and g2419 (n1758, \in0[120] , n_1807);
  and g2420 (n1759, n_1803, n1758);
  not g2421 (n_1808, \in1[121] );
  and g2422 (n1760, \in0[121] , n_1808);
  not g2423 (n_1809, n1759);
  not g2424 (n_1810, n1760);
  and g2425 (n1761, n_1809, n_1810);
  not g2426 (n_1811, \in1[122] );
  and g2427 (n1762, \in0[122] , n_1811);
  not g2428 (n_1812, n1762);
  and g2429 (n1763, n1761, n_1812);
  not g2430 (n_1813, n1763);
  and g2431 (n1764, n1751, n_1813);
  not g2432 (n_1814, n1757);
  not g2433 (n_1815, n1764);
  and g2434 (n1765, n_1814, n_1815);
  not g2435 (n_1816, n1756);
  and g2436 (n1766, n_1816, n1765);
  not g2437 (n_1818, \in0[124] );
  and g2438 (n1767, n_1818, \in1[124] );
  not g2439 (n_1822, \in1[127] );
  and g2440 (n1768, \in0[127] , n_1822);
  not g2441 (n_1824, \in0[126] );
  and g2442 (n1769, n_1824, \in1[126] );
  not g2443 (n_1827, \in0[125] );
  and g2444 (n1770, n_1827, \in1[125] );
  not g2445 (n_1829, n1769);
  not g2446 (n_1830, n1770);
  and g2447 (n1771, n_1829, n_1830);
  not g2448 (n_1831, n1768);
  not g2454 (n_1834, \in1[124] );
  and g2455 (n1775, \in0[124] , n_1834);
  not g2456 (n_1835, \in1[125] );
  and g2457 (n1776, \in0[125] , n_1835);
  not g2458 (n_1836, n1775);
  not g2459 (n_1837, n1776);
  and g2460 (n1777, n_1836, n_1837);
  not g2461 (n_1838, n1777);
  and g2462 (n1778, n1771, n_1838);
  not g2463 (n_1839, \in1[126] );
  and g2464 (n1779, \in0[126] , n_1839);
  not g2465 (n_1840, n1778);
  not g2466 (n_1841, n1779);
  and g2467 (n1780, n_1840, n_1841);
  not g2468 (n_1842, n1780);
  and g2469 (n1781, n_1831, n_1842);
  not g2470 (n_1843, n1774);
  not g2471 (n_1844, n1781);
  and g2472 (n1782, n_1843, n_1844);
  and g2473 (n1783, n_1822, n1782);
  not g2474 (n_1845, n1783);
  and g2475 (n1784, \in0[127] , n_1845);
  not g2476 (n_1846, n1784);
  and g2477 (n1785, n1213, n_1846);
  not g2478 (n_1847, \in0[127] );
  and g2479 (n1786, n_1847, \in1[127] );
  not g2480 (n_1848, n1786);
  and g2481 (n1787, n1782, n_1848);
  and g2482 (n1788, \in1[119] , n1787);
  not g2483 (n_1849, n1787);
  and g2484 (n1789, \in0[119] , n_1849);
  not g2485 (n_1850, n1788);
  not g2486 (n_1851, n1789);
  and g2487 (n1790, n_1850, n_1851);
  not g2488 (n_1852, \in2[127] );
  and g2489 (n1791, n_1852, \in3[127] );
  not g2490 (n_1853, n1791);
  and g2491 (n1792, n1211, n_1853);
  and g2492 (n1793, \in3[119] , n1792);
  not g2493 (n_1854, n1792);
  and g2494 (n1794, \in2[119] , n_1854);
  not g2495 (n_1855, n1793);
  not g2496 (n_1856, n1794);
  and g2497 (n1795, n_1855, n_1856);
  not g2498 (n_1857, n1790);
  and g2499 (n1796, n_1857, n1795);
  not g2500 (n_1858, n1795);
  and g2501 (n1797, n1790, n_1858);
  and g2502 (n1798, \in3[118] , n1792);
  and g2503 (n1799, \in2[118] , n_1854);
  not g2504 (n_1859, n1798);
  not g2505 (n_1860, n1799);
  and g2506 (n1800, n_1859, n_1860);
  and g2507 (n1801, \in1[118] , n1787);
  and g2508 (n1802, \in0[118] , n_1849);
  not g2509 (n_1861, n1801);
  not g2510 (n_1862, n1802);
  and g2511 (n1803, n_1861, n_1862);
  not g2512 (n_1863, n1800);
  and g2513 (n1804, n_1863, n1803);
  not g2514 (n_1864, n1797);
  not g2515 (n_1865, n1804);
  and g2516 (n1805, n_1864, n_1865);
  and g2517 (n1806, \in1[116] , n1787);
  and g2518 (n1807, \in0[116] , n_1849);
  not g2519 (n_1866, n1806);
  not g2520 (n_1867, n1807);
  and g2521 (n1808, n_1866, n_1867);
  and g2522 (n1809, \in1[117] , n1787);
  and g2523 (n1810, \in0[117] , n_1849);
  not g2524 (n_1868, n1809);
  not g2525 (n_1869, n1810);
  and g2526 (n1811, n_1868, n_1869);
  and g2527 (n1812, \in3[117] , n1792);
  and g2528 (n1813, \in2[117] , n_1854);
  not g2529 (n_1870, n1812);
  not g2530 (n_1871, n1813);
  and g2531 (n1814, n_1870, n_1871);
  not g2532 (n_1872, n1814);
  and g2533 (n1815, n1811, n_1872);
  and g2534 (n1816, \in3[116] , n1792);
  and g2535 (n1817, \in2[116] , n_1854);
  not g2536 (n_1873, n1816);
  not g2537 (n_1874, n1817);
  and g2538 (n1818, n_1873, n_1874);
  not g2539 (n_1875, n1815);
  and g2540 (n1819, n_1875, n1818);
  not g2541 (n_1876, n1808);
  and g2542 (n1820, n_1876, n1819);
  not g2543 (n_1877, n1811);
  and g2544 (n1821, n_1877, n1814);
  not g2545 (n_1878, n1820);
  not g2546 (n_1879, n1821);
  and g2547 (n1822, n_1878, n_1879);
  not g2548 (n_1880, n1822);
  and g2549 (n1823, n1805, n_1880);
  not g2550 (n_1881, n1803);
  and g2551 (n1824, n1800, n_1881);
  and g2552 (n1825, n_1864, n1824);
  and g2553 (n1826, \in3[112] , n1792);
  and g2554 (n1827, \in2[112] , n_1854);
  not g2555 (n_1882, n1826);
  not g2556 (n_1883, n1827);
  and g2557 (n1828, n_1882, n_1883);
  and g2558 (n1829, \in1[112] , n1787);
  and g2559 (n1830, \in0[112] , n_1849);
  not g2560 (n_1884, n1829);
  not g2561 (n_1885, n1830);
  and g2562 (n1831, n_1884, n_1885);
  not g2563 (n_1886, n1828);
  and g2564 (n1832, n_1886, n1831);
  and g2565 (n1833, \in1[115] , n1787);
  and g2566 (n1834, \in0[115] , n_1849);
  not g2567 (n_1887, n1833);
  not g2568 (n_1888, n1834);
  and g2569 (n1835, n_1887, n_1888);
  and g2570 (n1836, \in3[115] , n1792);
  and g2571 (n1837, \in2[115] , n_1854);
  not g2572 (n_1889, n1836);
  not g2573 (n_1890, n1837);
  and g2574 (n1838, n_1889, n_1890);
  not g2575 (n_1891, n1838);
  and g2576 (n1839, n1835, n_1891);
  and g2577 (n1840, \in3[114] , n1792);
  and g2578 (n1841, \in2[114] , n_1854);
  not g2579 (n_1892, n1840);
  not g2580 (n_1893, n1841);
  and g2581 (n1842, n_1892, n_1893);
  and g2582 (n1843, \in1[114] , n1787);
  and g2583 (n1844, \in0[114] , n_1849);
  not g2584 (n_1894, n1843);
  not g2585 (n_1895, n1844);
  and g2586 (n1845, n_1894, n_1895);
  not g2587 (n_1896, n1842);
  and g2588 (n1846, n_1896, n1845);
  not g2589 (n_1897, n1839);
  not g2590 (n_1898, n1846);
  and g2591 (n1847, n_1897, n_1898);
  and g2592 (n1848, \in1[113] , n1787);
  and g2593 (n1849, \in0[113] , n_1849);
  not g2594 (n_1899, n1848);
  not g2595 (n_1900, n1849);
  and g2596 (n1850, n_1899, n_1900);
  and g2597 (n1851, \in3[113] , n1792);
  and g2598 (n1852, \in2[113] , n_1854);
  not g2599 (n_1901, n1851);
  not g2600 (n_1902, n1852);
  and g2601 (n1853, n_1901, n_1902);
  not g2602 (n_1903, n1853);
  and g2603 (n1854, n1850, n_1903);
  and g2604 (n1855, \in1[111] , n1787);
  and g2605 (n1856, \in0[111] , n_1849);
  not g2606 (n_1904, n1855);
  not g2607 (n_1905, n1856);
  and g2608 (n1857, n_1904, n_1905);
  and g2609 (n1858, \in3[111] , n1792);
  and g2610 (n1859, \in2[111] , n_1854);
  not g2611 (n_1906, n1858);
  not g2612 (n_1907, n1859);
  and g2613 (n1860, n_1906, n_1907);
  not g2614 (n_1908, n1857);
  and g2615 (n1861, n_1908, n1860);
  not g2616 (n_1909, n1860);
  and g2617 (n1862, n1857, n_1909);
  and g2618 (n1863, \in3[110] , n1792);
  and g2619 (n1864, \in2[110] , n_1854);
  not g2620 (n_1910, n1863);
  not g2621 (n_1911, n1864);
  and g2622 (n1865, n_1910, n_1911);
  and g2623 (n1866, \in1[110] , n1787);
  and g2624 (n1867, \in0[110] , n_1849);
  not g2625 (n_1912, n1866);
  not g2626 (n_1913, n1867);
  and g2627 (n1868, n_1912, n_1913);
  not g2628 (n_1914, n1865);
  and g2629 (n1869, n_1914, n1868);
  not g2630 (n_1915, n1862);
  not g2631 (n_1916, n1869);
  and g2632 (n1870, n_1915, n_1916);
  and g2633 (n1871, \in1[109] , n1787);
  and g2634 (n1872, \in0[109] , n_1849);
  not g2635 (n_1917, n1871);
  not g2636 (n_1918, n1872);
  and g2637 (n1873, n_1917, n_1918);
  and g2638 (n1874, \in3[109] , n1792);
  and g2639 (n1875, \in2[109] , n_1854);
  not g2640 (n_1919, n1874);
  not g2641 (n_1920, n1875);
  and g2642 (n1876, n_1919, n_1920);
  not g2643 (n_1921, n1876);
  and g2644 (n1877, n1873, n_1921);
  and g2645 (n1878, \in1[108] , n1787);
  and g2646 (n1879, \in0[108] , n_1849);
  not g2647 (n_1922, n1878);
  not g2648 (n_1923, n1879);
  and g2649 (n1880, n_1922, n_1923);
  and g2650 (n1881, \in3[108] , n1792);
  and g2651 (n1882, \in2[108] , n_1854);
  not g2652 (n_1924, n1881);
  not g2653 (n_1925, n1882);
  and g2654 (n1883, n_1924, n_1925);
  not g2655 (n_1926, n1880);
  and g2656 (n1884, n_1926, n1883);
  not g2657 (n_1927, n1877);
  and g2658 (n1885, n_1927, n1884);
  not g2659 (n_1928, n1873);
  and g2660 (n1886, n_1928, n1876);
  not g2661 (n_1929, n1885);
  not g2662 (n_1930, n1886);
  and g2663 (n1887, n_1929, n_1930);
  not g2664 (n_1931, n1887);
  and g2665 (n1888, n1870, n_1931);
  not g2666 (n_1932, n1868);
  and g2667 (n1889, n1865, n_1932);
  and g2668 (n1890, n_1915, n1889);
  and g2669 (n1891, \in1[103] , n1787);
  and g2670 (n1892, \in0[103] , n_1849);
  not g2671 (n_1933, n1891);
  not g2672 (n_1934, n1892);
  and g2673 (n1893, n_1933, n_1934);
  and g2674 (n1894, \in3[103] , n1792);
  and g2675 (n1895, \in2[103] , n_1854);
  not g2676 (n_1935, n1894);
  not g2677 (n_1936, n1895);
  and g2678 (n1896, n_1935, n_1936);
  not g2679 (n_1937, n1893);
  and g2680 (n1897, n_1937, n1896);
  not g2681 (n_1938, n1896);
  and g2682 (n1898, n1893, n_1938);
  and g2683 (n1899, \in3[102] , n1792);
  and g2684 (n1900, \in2[102] , n_1854);
  not g2685 (n_1939, n1899);
  not g2686 (n_1940, n1900);
  and g2687 (n1901, n_1939, n_1940);
  and g2688 (n1902, \in1[102] , n1787);
  and g2689 (n1903, \in0[102] , n_1849);
  not g2690 (n_1941, n1902);
  not g2691 (n_1942, n1903);
  and g2692 (n1904, n_1941, n_1942);
  not g2693 (n_1943, n1901);
  and g2694 (n1905, n_1943, n1904);
  not g2695 (n_1944, n1898);
  not g2696 (n_1945, n1905);
  and g2697 (n1906, n_1944, n_1945);
  and g2698 (n1907, \in1[101] , n1787);
  and g2699 (n1908, \in0[101] , n_1849);
  not g2700 (n_1946, n1907);
  not g2701 (n_1947, n1908);
  and g2702 (n1909, n_1946, n_1947);
  and g2703 (n1910, \in3[101] , n1792);
  and g2704 (n1911, \in2[101] , n_1854);
  not g2705 (n_1948, n1910);
  not g2706 (n_1949, n1911);
  and g2707 (n1912, n_1948, n_1949);
  not g2708 (n_1950, n1912);
  and g2709 (n1913, n1909, n_1950);
  and g2710 (n1914, \in1[100] , n1787);
  and g2711 (n1915, \in0[100] , n_1849);
  not g2712 (n_1951, n1914);
  not g2713 (n_1952, n1915);
  and g2714 (n1916, n_1951, n_1952);
  and g2715 (n1917, \in3[100] , n1792);
  and g2716 (n1918, \in2[100] , n_1854);
  not g2717 (n_1953, n1917);
  not g2718 (n_1954, n1918);
  and g2719 (n1919, n_1953, n_1954);
  not g2720 (n_1955, n1916);
  and g2721 (n1920, n_1955, n1919);
  not g2722 (n_1956, n1913);
  and g2723 (n1921, n_1956, n1920);
  not g2724 (n_1957, n1909);
  and g2725 (n1922, n_1957, n1912);
  not g2726 (n_1958, n1921);
  not g2727 (n_1959, n1922);
  and g2728 (n1923, n_1958, n_1959);
  not g2729 (n_1960, n1923);
  and g2730 (n1924, n1906, n_1960);
  not g2731 (n_1961, n1904);
  and g2732 (n1925, n1901, n_1961);
  and g2733 (n1926, n_1944, n1925);
  and g2734 (n1927, \in3[96] , n1792);
  and g2735 (n1928, \in2[96] , n_1854);
  not g2736 (n_1962, n1927);
  not g2737 (n_1963, n1928);
  and g2738 (n1929, n_1962, n_1963);
  and g2739 (n1930, \in1[96] , n1787);
  and g2740 (n1931, \in0[96] , n_1849);
  not g2741 (n_1964, n1930);
  not g2742 (n_1965, n1931);
  and g2743 (n1932, n_1964, n_1965);
  not g2744 (n_1966, n1929);
  and g2745 (n1933, n_1966, n1932);
  and g2746 (n1934, \in1[99] , n1787);
  and g2747 (n1935, \in0[99] , n_1849);
  not g2748 (n_1967, n1934);
  not g2749 (n_1968, n1935);
  and g2750 (n1936, n_1967, n_1968);
  and g2751 (n1937, \in3[99] , n1792);
  and g2752 (n1938, \in2[99] , n_1854);
  not g2753 (n_1969, n1937);
  not g2754 (n_1970, n1938);
  and g2755 (n1939, n_1969, n_1970);
  not g2756 (n_1971, n1939);
  and g2757 (n1940, n1936, n_1971);
  and g2758 (n1941, \in3[98] , n1792);
  and g2759 (n1942, \in2[98] , n_1854);
  not g2760 (n_1972, n1941);
  not g2761 (n_1973, n1942);
  and g2762 (n1943, n_1972, n_1973);
  and g2763 (n1944, \in1[98] , n1787);
  and g2764 (n1945, \in0[98] , n_1849);
  not g2765 (n_1974, n1944);
  not g2766 (n_1975, n1945);
  and g2767 (n1946, n_1974, n_1975);
  not g2768 (n_1976, n1943);
  and g2769 (n1947, n_1976, n1946);
  not g2770 (n_1977, n1940);
  not g2771 (n_1978, n1947);
  and g2772 (n1948, n_1977, n_1978);
  and g2773 (n1949, \in1[97] , n1787);
  and g2774 (n1950, \in0[97] , n_1849);
  not g2775 (n_1979, n1949);
  not g2776 (n_1980, n1950);
  and g2777 (n1951, n_1979, n_1980);
  and g2778 (n1952, \in3[97] , n1792);
  and g2779 (n1953, \in2[97] , n_1854);
  not g2780 (n_1981, n1952);
  not g2781 (n_1982, n1953);
  and g2782 (n1954, n_1981, n_1982);
  not g2783 (n_1983, n1954);
  and g2784 (n1955, n1951, n_1983);
  and g2785 (n1956, \in1[95] , n1787);
  and g2786 (n1957, \in0[95] , n_1849);
  not g2787 (n_1984, n1956);
  not g2788 (n_1985, n1957);
  and g2789 (n1958, n_1984, n_1985);
  and g2790 (n1959, \in3[95] , n1792);
  and g2791 (n1960, \in2[95] , n_1854);
  not g2792 (n_1986, n1959);
  not g2793 (n_1987, n1960);
  and g2794 (n1961, n_1986, n_1987);
  not g2795 (n_1988, n1958);
  and g2796 (n1962, n_1988, n1961);
  not g2797 (n_1989, n1961);
  and g2798 (n1963, n1958, n_1989);
  and g2799 (n1964, \in3[94] , n1792);
  and g2800 (n1965, \in2[94] , n_1854);
  not g2801 (n_1990, n1964);
  not g2802 (n_1991, n1965);
  and g2803 (n1966, n_1990, n_1991);
  and g2804 (n1967, \in1[94] , n1787);
  and g2805 (n1968, \in0[94] , n_1849);
  not g2806 (n_1992, n1967);
  not g2807 (n_1993, n1968);
  and g2808 (n1969, n_1992, n_1993);
  not g2809 (n_1994, n1966);
  and g2810 (n1970, n_1994, n1969);
  not g2811 (n_1995, n1963);
  not g2812 (n_1996, n1970);
  and g2813 (n1971, n_1995, n_1996);
  and g2814 (n1972, \in1[93] , n1787);
  and g2815 (n1973, \in0[93] , n_1849);
  not g2816 (n_1997, n1972);
  not g2817 (n_1998, n1973);
  and g2818 (n1974, n_1997, n_1998);
  and g2819 (n1975, \in3[93] , n1792);
  and g2820 (n1976, \in2[93] , n_1854);
  not g2821 (n_1999, n1975);
  not g2822 (n_2000, n1976);
  and g2823 (n1977, n_1999, n_2000);
  not g2824 (n_2001, n1977);
  and g2825 (n1978, n1974, n_2001);
  and g2826 (n1979, \in1[92] , n1787);
  and g2827 (n1980, \in0[92] , n_1849);
  not g2828 (n_2002, n1979);
  not g2829 (n_2003, n1980);
  and g2830 (n1981, n_2002, n_2003);
  and g2831 (n1982, \in3[92] , n1792);
  and g2832 (n1983, \in2[92] , n_1854);
  not g2833 (n_2004, n1982);
  not g2834 (n_2005, n1983);
  and g2835 (n1984, n_2004, n_2005);
  not g2836 (n_2006, n1981);
  and g2837 (n1985, n_2006, n1984);
  not g2838 (n_2007, n1978);
  and g2839 (n1986, n_2007, n1985);
  not g2840 (n_2008, n1974);
  and g2841 (n1987, n_2008, n1977);
  not g2842 (n_2009, n1986);
  not g2843 (n_2010, n1987);
  and g2844 (n1988, n_2009, n_2010);
  not g2845 (n_2011, n1988);
  and g2846 (n1989, n1971, n_2011);
  not g2847 (n_2012, n1969);
  and g2848 (n1990, n1966, n_2012);
  and g2849 (n1991, n_1995, n1990);
  and g2850 (n1992, \in1[87] , n1787);
  and g2851 (n1993, \in0[87] , n_1849);
  not g2852 (n_2013, n1992);
  not g2853 (n_2014, n1993);
  and g2854 (n1994, n_2013, n_2014);
  and g2855 (n1995, \in3[87] , n1792);
  and g2856 (n1996, \in2[87] , n_1854);
  not g2857 (n_2015, n1995);
  not g2858 (n_2016, n1996);
  and g2859 (n1997, n_2015, n_2016);
  not g2860 (n_2017, n1994);
  and g2861 (n1998, n_2017, n1997);
  not g2862 (n_2018, n1997);
  and g2863 (n1999, n1994, n_2018);
  and g2864 (n2000, \in3[86] , n1792);
  and g2865 (n2001, \in2[86] , n_1854);
  not g2866 (n_2019, n2000);
  not g2867 (n_2020, n2001);
  and g2868 (n2002, n_2019, n_2020);
  and g2869 (n2003, \in1[86] , n1787);
  and g2870 (n2004, \in0[86] , n_1849);
  not g2871 (n_2021, n2003);
  not g2872 (n_2022, n2004);
  and g2873 (n2005, n_2021, n_2022);
  not g2874 (n_2023, n2002);
  and g2875 (n2006, n_2023, n2005);
  not g2876 (n_2024, n1999);
  not g2877 (n_2025, n2006);
  and g2878 (n2007, n_2024, n_2025);
  and g2879 (n2008, \in1[85] , n1787);
  and g2880 (n2009, \in0[85] , n_1849);
  not g2881 (n_2026, n2008);
  not g2882 (n_2027, n2009);
  and g2883 (n2010, n_2026, n_2027);
  and g2884 (n2011, \in3[85] , n1792);
  and g2885 (n2012, \in2[85] , n_1854);
  not g2886 (n_2028, n2011);
  not g2887 (n_2029, n2012);
  and g2888 (n2013, n_2028, n_2029);
  not g2889 (n_2030, n2013);
  and g2890 (n2014, n2010, n_2030);
  and g2891 (n2015, \in1[84] , n1787);
  and g2892 (n2016, \in0[84] , n_1849);
  not g2893 (n_2031, n2015);
  not g2894 (n_2032, n2016);
  and g2895 (n2017, n_2031, n_2032);
  and g2896 (n2018, \in3[84] , n1792);
  and g2897 (n2019, \in2[84] , n_1854);
  not g2898 (n_2033, n2018);
  not g2899 (n_2034, n2019);
  and g2900 (n2020, n_2033, n_2034);
  not g2901 (n_2035, n2017);
  and g2902 (n2021, n_2035, n2020);
  not g2903 (n_2036, n2014);
  and g2904 (n2022, n_2036, n2021);
  not g2905 (n_2037, n2010);
  and g2906 (n2023, n_2037, n2013);
  not g2907 (n_2038, n2022);
  not g2908 (n_2039, n2023);
  and g2909 (n2024, n_2038, n_2039);
  not g2910 (n_2040, n2024);
  and g2911 (n2025, n2007, n_2040);
  not g2912 (n_2041, n2005);
  and g2913 (n2026, n2002, n_2041);
  and g2914 (n2027, n_2024, n2026);
  and g2915 (n2028, \in3[80] , n1792);
  and g2916 (n2029, \in2[80] , n_1854);
  not g2917 (n_2042, n2028);
  not g2918 (n_2043, n2029);
  and g2919 (n2030, n_2042, n_2043);
  and g2920 (n2031, \in1[80] , n1787);
  and g2921 (n2032, \in0[80] , n_1849);
  not g2922 (n_2044, n2031);
  not g2923 (n_2045, n2032);
  and g2924 (n2033, n_2044, n_2045);
  not g2925 (n_2046, n2030);
  and g2926 (n2034, n_2046, n2033);
  and g2927 (n2035, \in1[83] , n1787);
  and g2928 (n2036, \in0[83] , n_1849);
  not g2929 (n_2047, n2035);
  not g2930 (n_2048, n2036);
  and g2931 (n2037, n_2047, n_2048);
  and g2932 (n2038, \in3[83] , n1792);
  and g2933 (n2039, \in2[83] , n_1854);
  not g2934 (n_2049, n2038);
  not g2935 (n_2050, n2039);
  and g2936 (n2040, n_2049, n_2050);
  not g2937 (n_2051, n2040);
  and g2938 (n2041, n2037, n_2051);
  and g2939 (n2042, \in3[82] , n1792);
  and g2940 (n2043, \in2[82] , n_1854);
  not g2941 (n_2052, n2042);
  not g2942 (n_2053, n2043);
  and g2943 (n2044, n_2052, n_2053);
  and g2944 (n2045, \in1[82] , n1787);
  and g2945 (n2046, \in0[82] , n_1849);
  not g2946 (n_2054, n2045);
  not g2947 (n_2055, n2046);
  and g2948 (n2047, n_2054, n_2055);
  not g2949 (n_2056, n2044);
  and g2950 (n2048, n_2056, n2047);
  not g2951 (n_2057, n2041);
  not g2952 (n_2058, n2048);
  and g2953 (n2049, n_2057, n_2058);
  and g2954 (n2050, \in1[81] , n1787);
  and g2955 (n2051, \in0[81] , n_1849);
  not g2956 (n_2059, n2050);
  not g2957 (n_2060, n2051);
  and g2958 (n2052, n_2059, n_2060);
  and g2959 (n2053, \in3[81] , n1792);
  and g2960 (n2054, \in2[81] , n_1854);
  not g2961 (n_2061, n2053);
  not g2962 (n_2062, n2054);
  and g2963 (n2055, n_2061, n_2062);
  not g2964 (n_2063, n2055);
  and g2965 (n2056, n2052, n_2063);
  and g2966 (n2057, \in1[79] , n1787);
  and g2967 (n2058, \in0[79] , n_1849);
  not g2968 (n_2064, n2057);
  not g2969 (n_2065, n2058);
  and g2970 (n2059, n_2064, n_2065);
  and g2971 (n2060, \in3[79] , n1792);
  and g2972 (n2061, \in2[79] , n_1854);
  not g2973 (n_2066, n2060);
  not g2974 (n_2067, n2061);
  and g2975 (n2062, n_2066, n_2067);
  not g2976 (n_2068, n2059);
  and g2977 (n2063, n_2068, n2062);
  not g2978 (n_2069, n2062);
  and g2979 (n2064, n2059, n_2069);
  and g2980 (n2065, \in3[78] , n1792);
  and g2981 (n2066, \in2[78] , n_1854);
  not g2982 (n_2070, n2065);
  not g2983 (n_2071, n2066);
  and g2984 (n2067, n_2070, n_2071);
  and g2985 (n2068, \in1[78] , n1787);
  and g2986 (n2069, \in0[78] , n_1849);
  not g2987 (n_2072, n2068);
  not g2988 (n_2073, n2069);
  and g2989 (n2070, n_2072, n_2073);
  not g2990 (n_2074, n2067);
  and g2991 (n2071, n_2074, n2070);
  not g2992 (n_2075, n2064);
  not g2993 (n_2076, n2071);
  and g2994 (n2072, n_2075, n_2076);
  and g2995 (n2073, \in1[77] , n1787);
  and g2996 (n2074, \in0[77] , n_1849);
  not g2997 (n_2077, n2073);
  not g2998 (n_2078, n2074);
  and g2999 (n2075, n_2077, n_2078);
  and g3000 (n2076, \in3[77] , n1792);
  and g3001 (n2077, \in2[77] , n_1854);
  not g3002 (n_2079, n2076);
  not g3003 (n_2080, n2077);
  and g3004 (n2078, n_2079, n_2080);
  not g3005 (n_2081, n2078);
  and g3006 (n2079, n2075, n_2081);
  and g3007 (n2080, \in1[76] , n1787);
  and g3008 (n2081, \in0[76] , n_1849);
  not g3009 (n_2082, n2080);
  not g3010 (n_2083, n2081);
  and g3011 (n2082, n_2082, n_2083);
  and g3012 (n2083, \in3[76] , n1792);
  and g3013 (n2084, \in2[76] , n_1854);
  not g3014 (n_2084, n2083);
  not g3015 (n_2085, n2084);
  and g3016 (n2085, n_2084, n_2085);
  not g3017 (n_2086, n2082);
  and g3018 (n2086, n_2086, n2085);
  not g3019 (n_2087, n2079);
  and g3020 (n2087, n_2087, n2086);
  not g3021 (n_2088, n2075);
  and g3022 (n2088, n_2088, n2078);
  not g3023 (n_2089, n2087);
  not g3024 (n_2090, n2088);
  and g3025 (n2089, n_2089, n_2090);
  not g3026 (n_2091, n2089);
  and g3027 (n2090, n2072, n_2091);
  not g3028 (n_2092, n2070);
  and g3029 (n2091, n2067, n_2092);
  and g3030 (n2092, n_2075, n2091);
  and g3031 (n2093, \in1[71] , n1787);
  and g3032 (n2094, \in0[71] , n_1849);
  not g3033 (n_2093, n2093);
  not g3034 (n_2094, n2094);
  and g3035 (n2095, n_2093, n_2094);
  and g3036 (n2096, \in3[71] , n1792);
  and g3037 (n2097, \in2[71] , n_1854);
  not g3038 (n_2095, n2096);
  not g3039 (n_2096, n2097);
  and g3040 (n2098, n_2095, n_2096);
  not g3041 (n_2097, n2095);
  and g3042 (n2099, n_2097, n2098);
  not g3043 (n_2098, n2098);
  and g3044 (n2100, n2095, n_2098);
  and g3045 (n2101, \in3[70] , n1792);
  and g3046 (n2102, \in2[70] , n_1854);
  not g3047 (n_2099, n2101);
  not g3048 (n_2100, n2102);
  and g3049 (n2103, n_2099, n_2100);
  and g3050 (n2104, \in1[70] , n1787);
  and g3051 (n2105, \in0[70] , n_1849);
  not g3052 (n_2101, n2104);
  not g3053 (n_2102, n2105);
  and g3054 (n2106, n_2101, n_2102);
  not g3055 (n_2103, n2103);
  and g3056 (n2107, n_2103, n2106);
  not g3057 (n_2104, n2100);
  not g3058 (n_2105, n2107);
  and g3059 (n2108, n_2104, n_2105);
  and g3060 (n2109, \in1[69] , n1787);
  and g3061 (n2110, \in0[69] , n_1849);
  not g3062 (n_2106, n2109);
  not g3063 (n_2107, n2110);
  and g3064 (n2111, n_2106, n_2107);
  and g3065 (n2112, \in3[69] , n1792);
  and g3066 (n2113, \in2[69] , n_1854);
  not g3067 (n_2108, n2112);
  not g3068 (n_2109, n2113);
  and g3069 (n2114, n_2108, n_2109);
  not g3070 (n_2110, n2114);
  and g3071 (n2115, n2111, n_2110);
  and g3072 (n2116, \in1[68] , n1787);
  and g3073 (n2117, \in0[68] , n_1849);
  not g3074 (n_2111, n2116);
  not g3075 (n_2112, n2117);
  and g3076 (n2118, n_2111, n_2112);
  and g3077 (n2119, \in3[68] , n1792);
  and g3078 (n2120, \in2[68] , n_1854);
  not g3079 (n_2113, n2119);
  not g3080 (n_2114, n2120);
  and g3081 (n2121, n_2113, n_2114);
  not g3082 (n_2115, n2118);
  and g3083 (n2122, n_2115, n2121);
  not g3084 (n_2116, n2115);
  and g3085 (n2123, n_2116, n2122);
  not g3086 (n_2117, n2111);
  and g3087 (n2124, n_2117, n2114);
  not g3088 (n_2118, n2123);
  not g3089 (n_2119, n2124);
  and g3090 (n2125, n_2118, n_2119);
  not g3091 (n_2120, n2125);
  and g3092 (n2126, n2108, n_2120);
  not g3093 (n_2121, n2106);
  and g3094 (n2127, n2103, n_2121);
  and g3095 (n2128, n_2104, n2127);
  and g3096 (n2129, \in1[67] , n1787);
  and g3097 (n2130, \in0[67] , n_1849);
  not g3098 (n_2122, n2129);
  not g3099 (n_2123, n2130);
  and g3100 (n2131, n_2122, n_2123);
  and g3101 (n2132, \in3[67] , n1792);
  and g3102 (n2133, \in2[67] , n_1854);
  not g3103 (n_2124, n2132);
  not g3104 (n_2125, n2133);
  and g3105 (n2134, n_2124, n_2125);
  not g3106 (n_2126, n2134);
  and g3107 (n2135, n2131, n_2126);
  and g3108 (n2136, \in3[66] , n1792);
  and g3109 (n2137, \in2[66] , n_1854);
  not g3110 (n_2127, n2136);
  not g3111 (n_2128, n2137);
  and g3112 (n2138, n_2127, n_2128);
  and g3113 (n2139, \in1[66] , n1787);
  and g3114 (n2140, \in0[66] , n_1849);
  not g3115 (n_2129, n2139);
  not g3116 (n_2130, n2140);
  and g3117 (n2141, n_2129, n_2130);
  not g3118 (n_2131, n2138);
  and g3119 (n2142, n_2131, n2141);
  not g3120 (n_2132, n2135);
  not g3121 (n_2133, n2142);
  and g3122 (n2143, n_2132, n_2133);
  and g3123 (n2144, \in3[64] , n1792);
  and g3124 (n2145, \in2[64] , n_1854);
  not g3125 (n_2134, n2144);
  not g3126 (n_2135, n2145);
  and g3127 (n2146, n_2134, n_2135);
  and g3128 (n2147, \in1[64] , n1787);
  and g3129 (n2148, \in0[64] , n_1849);
  not g3130 (n_2136, n2147);
  not g3131 (n_2137, n2148);
  and g3132 (n2149, n_2136, n_2137);
  not g3133 (n_2138, n2146);
  and g3134 (n2150, n_2138, n2149);
  and g3135 (n2151, \in1[65] , n1787);
  and g3136 (n2152, \in0[65] , n_1849);
  not g3137 (n_2139, n2151);
  not g3138 (n_2140, n2152);
  and g3139 (n2153, n_2139, n_2140);
  and g3140 (n2154, \in3[65] , n1792);
  and g3141 (n2155, \in2[65] , n_1854);
  not g3142 (n_2141, n2154);
  not g3143 (n_2142, n2155);
  and g3144 (n2156, n_2141, n_2142);
  not g3145 (n_2143, n2156);
  and g3146 (n2157, n2153, n_2143);
  and g3147 (n2158, \in1[63] , n1787);
  and g3148 (n2159, \in0[63] , n_1849);
  not g3149 (n_2144, n2158);
  not g3150 (n_2145, n2159);
  and g3151 (n2160, n_2144, n_2145);
  and g3152 (n2161, \in3[63] , n1792);
  and g3153 (n2162, \in2[63] , n_1854);
  not g3154 (n_2146, n2161);
  not g3155 (n_2147, n2162);
  and g3156 (n2163, n_2146, n_2147);
  not g3157 (n_2148, n2160);
  and g3158 (n2164, n_2148, n2163);
  not g3159 (n_2149, n2163);
  and g3160 (n2165, n2160, n_2149);
  and g3161 (n2166, \in3[62] , n1792);
  and g3162 (n2167, \in2[62] , n_1854);
  not g3163 (n_2150, n2166);
  not g3164 (n_2151, n2167);
  and g3165 (n2168, n_2150, n_2151);
  and g3166 (n2169, \in1[62] , n1787);
  and g3167 (n2170, \in0[62] , n_1849);
  not g3168 (n_2152, n2169);
  not g3169 (n_2153, n2170);
  and g3170 (n2171, n_2152, n_2153);
  not g3171 (n_2154, n2168);
  and g3172 (n2172, n_2154, n2171);
  not g3173 (n_2155, n2165);
  not g3174 (n_2156, n2172);
  and g3175 (n2173, n_2155, n_2156);
  and g3176 (n2174, \in1[60] , n1787);
  and g3177 (n2175, \in0[60] , n_1849);
  not g3178 (n_2157, n2174);
  not g3179 (n_2158, n2175);
  and g3180 (n2176, n_2157, n_2158);
  and g3181 (n2177, \in3[60] , n1792);
  and g3182 (n2178, \in2[60] , n_1854);
  not g3183 (n_2159, n2177);
  not g3184 (n_2160, n2178);
  and g3185 (n2179, n_2159, n_2160);
  not g3186 (n_2161, n2179);
  and g3187 (n2180, n2176, n_2161);
  and g3188 (n2181, \in1[61] , n1787);
  and g3189 (n2182, \in0[61] , n_1849);
  not g3190 (n_2162, n2181);
  not g3191 (n_2163, n2182);
  and g3192 (n2183, n_2162, n_2163);
  and g3193 (n2184, \in3[61] , n1792);
  and g3194 (n2185, \in2[61] , n_1854);
  not g3195 (n_2164, n2184);
  not g3196 (n_2165, n2185);
  and g3197 (n2186, n_2164, n_2165);
  not g3198 (n_2166, n2186);
  and g3199 (n2187, n2183, n_2166);
  not g3200 (n_2167, n2180);
  not g3201 (n_2168, n2187);
  and g3202 (n2188, n_2167, n_2168);
  and g3203 (n2189, n2173, n2188);
  and g3204 (n2190, \in1[59] , n1787);
  and g3205 (n2191, \in0[59] , n_1849);
  not g3206 (n_2169, n2190);
  not g3207 (n_2170, n2191);
  and g3208 (n2192, n_2169, n_2170);
  and g3209 (n2193, \in3[59] , n1792);
  and g3210 (n2194, \in2[59] , n_1854);
  not g3211 (n_2171, n2193);
  not g3212 (n_2172, n2194);
  and g3213 (n2195, n_2171, n_2172);
  not g3214 (n_2173, n2192);
  and g3215 (n2196, n_2173, n2195);
  not g3216 (n_2174, n2195);
  and g3217 (n2197, n2192, n_2174);
  and g3218 (n2198, \in1[58] , n1787);
  and g3219 (n2199, \in0[58] , n_1849);
  not g3220 (n_2175, n2198);
  not g3221 (n_2176, n2199);
  and g3222 (n2200, n_2175, n_2176);
  and g3223 (n2201, \in3[58] , n1792);
  and g3224 (n2202, \in2[58] , n_1854);
  not g3225 (n_2177, n2201);
  not g3226 (n_2178, n2202);
  and g3227 (n2203, n_2177, n_2178);
  not g3228 (n_2179, n2203);
  and g3229 (n2204, n2200, n_2179);
  not g3230 (n_2180, n2197);
  not g3231 (n_2181, n2204);
  and g3232 (n2205, n_2180, n_2181);
  and g3233 (n2206, \in1[57] , n1787);
  and g3234 (n2207, \in0[57] , n_1849);
  not g3235 (n_2182, n2206);
  not g3236 (n_2183, n2207);
  and g3237 (n2208, n_2182, n_2183);
  and g3238 (n2209, \in3[57] , n1792);
  and g3239 (n2210, \in2[57] , n_1854);
  not g3240 (n_2184, n2209);
  not g3241 (n_2185, n2210);
  and g3242 (n2211, n_2184, n_2185);
  not g3243 (n_2186, n2211);
  and g3244 (n2212, n2208, n_2186);
  and g3245 (n2213, \in1[56] , n1787);
  and g3246 (n2214, \in0[56] , n_1849);
  not g3247 (n_2187, n2213);
  not g3248 (n_2188, n2214);
  and g3249 (n2215, n_2187, n_2188);
  and g3250 (n2216, \in3[56] , n1792);
  and g3251 (n2217, \in2[56] , n_1854);
  not g3252 (n_2189, n2216);
  not g3253 (n_2190, n2217);
  and g3254 (n2218, n_2189, n_2190);
  not g3255 (n_2191, n2215);
  and g3256 (n2219, n_2191, n2218);
  not g3257 (n_2192, n2212);
  and g3258 (n2220, n_2192, n2219);
  not g3259 (n_2193, n2208);
  and g3260 (n2221, n_2193, n2211);
  not g3261 (n_2194, n2220);
  not g3262 (n_2195, n2221);
  and g3263 (n2222, n_2194, n_2195);
  not g3264 (n_2196, n2200);
  and g3265 (n2223, n_2196, n2203);
  not g3266 (n_2197, n2223);
  and g3267 (n2224, n2222, n_2197);
  not g3268 (n_2198, n2224);
  and g3269 (n2225, n2205, n_2198);
  not g3270 (n_2199, n2196);
  not g3271 (n_2200, n2225);
  and g3272 (n2226, n_2199, n_2200);
  not g3273 (n_2201, n2226);
  and g3274 (n2227, n2189, n_2201);
  not g3275 (n_2202, n2176);
  and g3276 (n2228, n_2202, n2179);
  and g3277 (n2229, n_2168, n2228);
  not g3278 (n_2203, n2183);
  and g3279 (n2230, n_2203, n2186);
  not g3280 (n_2204, n2229);
  not g3281 (n_2205, n2230);
  and g3282 (n2231, n_2204, n_2205);
  not g3283 (n_2206, n2231);
  and g3284 (n2232, n2173, n_2206);
  not g3285 (n_2207, n2171);
  and g3286 (n2233, n2168, n_2207);
  and g3287 (n2234, n_2155, n2233);
  and g3288 (n2235, \in1[47] , n1787);
  and g3289 (n2236, \in0[47] , n_1849);
  not g3290 (n_2208, n2235);
  not g3291 (n_2209, n2236);
  and g3292 (n2237, n_2208, n_2209);
  and g3293 (n2238, \in3[47] , n1792);
  and g3294 (n2239, \in2[47] , n_1854);
  not g3295 (n_2210, n2238);
  not g3296 (n_2211, n2239);
  and g3297 (n2240, n_2210, n_2211);
  not g3298 (n_2212, n2237);
  and g3299 (n2241, n_2212, n2240);
  not g3300 (n_2213, n2240);
  and g3301 (n2242, n2237, n_2213);
  and g3302 (n2243, \in3[46] , n1792);
  and g3303 (n2244, \in2[46] , n_1854);
  not g3304 (n_2214, n2243);
  not g3305 (n_2215, n2244);
  and g3306 (n2245, n_2214, n_2215);
  and g3307 (n2246, \in1[46] , n1787);
  and g3308 (n2247, \in0[46] , n_1849);
  not g3309 (n_2216, n2246);
  not g3310 (n_2217, n2247);
  and g3311 (n2248, n_2216, n_2217);
  not g3312 (n_2218, n2245);
  and g3313 (n2249, n_2218, n2248);
  not g3314 (n_2219, n2242);
  not g3315 (n_2220, n2249);
  and g3316 (n2250, n_2219, n_2220);
  and g3317 (n2251, \in1[44] , n1787);
  and g3318 (n2252, \in0[44] , n_1849);
  not g3319 (n_2221, n2251);
  not g3320 (n_2222, n2252);
  and g3321 (n2253, n_2221, n_2222);
  and g3322 (n2254, \in3[44] , n1792);
  and g3323 (n2255, \in2[44] , n_1854);
  not g3324 (n_2223, n2254);
  not g3325 (n_2224, n2255);
  and g3326 (n2256, n_2223, n_2224);
  not g3327 (n_2225, n2256);
  and g3328 (n2257, n2253, n_2225);
  and g3329 (n2258, \in1[45] , n1787);
  and g3330 (n2259, \in0[45] , n_1849);
  not g3331 (n_2226, n2258);
  not g3332 (n_2227, n2259);
  and g3333 (n2260, n_2226, n_2227);
  and g3334 (n2261, \in3[45] , n1792);
  and g3335 (n2262, \in2[45] , n_1854);
  not g3336 (n_2228, n2261);
  not g3337 (n_2229, n2262);
  and g3338 (n2263, n_2228, n_2229);
  not g3339 (n_2230, n2263);
  and g3340 (n2264, n2260, n_2230);
  not g3341 (n_2231, n2257);
  not g3342 (n_2232, n2264);
  and g3343 (n2265, n_2231, n_2232);
  and g3344 (n2266, n2250, n2265);
  and g3345 (n2267, \in1[43] , n1787);
  and g3346 (n2268, \in0[43] , n_1849);
  not g3347 (n_2233, n2267);
  not g3348 (n_2234, n2268);
  and g3349 (n2269, n_2233, n_2234);
  and g3350 (n2270, \in3[43] , n1792);
  and g3351 (n2271, \in2[43] , n_1854);
  not g3352 (n_2235, n2270);
  not g3353 (n_2236, n2271);
  and g3354 (n2272, n_2235, n_2236);
  not g3355 (n_2237, n2269);
  and g3356 (n2273, n_2237, n2272);
  not g3357 (n_2238, n2272);
  and g3358 (n2274, n2269, n_2238);
  and g3359 (n2275, \in1[42] , n1787);
  and g3360 (n2276, \in0[42] , n_1849);
  not g3361 (n_2239, n2275);
  not g3362 (n_2240, n2276);
  and g3363 (n2277, n_2239, n_2240);
  and g3364 (n2278, \in3[42] , n1792);
  and g3365 (n2279, \in2[42] , n_1854);
  not g3366 (n_2241, n2278);
  not g3367 (n_2242, n2279);
  and g3368 (n2280, n_2241, n_2242);
  not g3369 (n_2243, n2280);
  and g3370 (n2281, n2277, n_2243);
  not g3371 (n_2244, n2274);
  not g3372 (n_2245, n2281);
  and g3373 (n2282, n_2244, n_2245);
  and g3374 (n2283, \in1[41] , n1787);
  and g3375 (n2284, \in0[41] , n_1849);
  not g3376 (n_2246, n2283);
  not g3377 (n_2247, n2284);
  and g3378 (n2285, n_2246, n_2247);
  and g3379 (n2286, \in3[41] , n1792);
  and g3380 (n2287, \in2[41] , n_1854);
  not g3381 (n_2248, n2286);
  not g3382 (n_2249, n2287);
  and g3383 (n2288, n_2248, n_2249);
  not g3384 (n_2250, n2288);
  and g3385 (n2289, n2285, n_2250);
  and g3386 (n2290, \in1[40] , n1787);
  and g3387 (n2291, \in0[40] , n_1849);
  not g3388 (n_2251, n2290);
  not g3389 (n_2252, n2291);
  and g3390 (n2292, n_2251, n_2252);
  and g3391 (n2293, \in3[40] , n1792);
  and g3392 (n2294, \in2[40] , n_1854);
  not g3393 (n_2253, n2293);
  not g3394 (n_2254, n2294);
  and g3395 (n2295, n_2253, n_2254);
  not g3396 (n_2255, n2292);
  and g3397 (n2296, n_2255, n2295);
  not g3398 (n_2256, n2289);
  and g3399 (n2297, n_2256, n2296);
  not g3400 (n_2257, n2285);
  and g3401 (n2298, n_2257, n2288);
  not g3402 (n_2258, n2297);
  not g3403 (n_2259, n2298);
  and g3404 (n2299, n_2258, n_2259);
  not g3405 (n_2260, n2277);
  and g3406 (n2300, n_2260, n2280);
  not g3407 (n_2261, n2300);
  and g3408 (n2301, n2299, n_2261);
  not g3409 (n_2262, n2301);
  and g3410 (n2302, n2282, n_2262);
  not g3411 (n_2263, n2273);
  not g3412 (n_2264, n2302);
  and g3413 (n2303, n_2263, n_2264);
  not g3414 (n_2265, n2303);
  and g3415 (n2304, n2266, n_2265);
  not g3416 (n_2266, n2253);
  and g3417 (n2305, n_2266, n2256);
  and g3418 (n2306, n_2232, n2305);
  not g3419 (n_2267, n2260);
  and g3420 (n2307, n_2267, n2263);
  not g3421 (n_2268, n2306);
  not g3422 (n_2269, n2307);
  and g3423 (n2308, n_2268, n_2269);
  not g3424 (n_2270, n2308);
  and g3425 (n2309, n2250, n_2270);
  not g3426 (n_2271, n2248);
  and g3427 (n2310, n2245, n_2271);
  and g3428 (n2311, n_2219, n2310);
  and g3429 (n2312, \in3[32] , n1792);
  and g3430 (n2313, \in2[32] , n_1854);
  not g3431 (n_2272, n2312);
  not g3432 (n_2273, n2313);
  and g3433 (n2314, n_2272, n_2273);
  and g3434 (n2315, \in1[32] , n1787);
  and g3435 (n2316, \in0[32] , n_1849);
  not g3436 (n_2274, n2315);
  not g3437 (n_2275, n2316);
  and g3438 (n2317, n_2274, n_2275);
  not g3439 (n_2276, n2314);
  and g3440 (n2318, n_2276, n2317);
  and g3441 (n2319, \in1[31] , n1787);
  and g3442 (n2320, \in0[31] , n_1849);
  not g3443 (n_2277, n2319);
  not g3444 (n_2278, n2320);
  and g3445 (n2321, n_2277, n_2278);
  and g3446 (n2322, \in3[31] , n1792);
  and g3447 (n2323, \in2[31] , n_1854);
  not g3448 (n_2279, n2322);
  not g3449 (n_2280, n2323);
  and g3450 (n2324, n_2279, n_2280);
  not g3451 (n_2281, n2324);
  and g3452 (n2325, n2321, n_2281);
  and g3453 (n2326, \in1[30] , n1787);
  and g3454 (n2327, \in0[30] , n_1849);
  not g3455 (n_2282, n2326);
  not g3456 (n_2283, n2327);
  and g3457 (n2328, n_2282, n_2283);
  and g3458 (n2329, \in3[30] , n1792);
  and g3459 (n2330, \in2[30] , n_1854);
  not g3460 (n_2284, n2329);
  not g3461 (n_2285, n2330);
  and g3462 (n2331, n_2284, n_2285);
  not g3463 (n_2286, n2331);
  and g3464 (n2332, n2328, n_2286);
  and g3465 (n2333, \in1[29] , n1787);
  and g3466 (n2334, \in0[29] , n_1849);
  not g3467 (n_2287, n2333);
  not g3468 (n_2288, n2334);
  and g3469 (n2335, n_2287, n_2288);
  and g3470 (n2336, \in3[29] , n1792);
  and g3471 (n2337, \in2[29] , n_1854);
  not g3472 (n_2289, n2336);
  not g3473 (n_2290, n2337);
  and g3474 (n2338, n_2289, n_2290);
  not g3475 (n_2291, n2338);
  and g3476 (n2339, n2335, n_2291);
  and g3477 (n2340, \in1[28] , n1787);
  and g3478 (n2341, \in0[28] , n_1849);
  not g3479 (n_2292, n2340);
  not g3480 (n_2293, n2341);
  and g3481 (n2342, n_2292, n_2293);
  and g3482 (n2343, \in3[28] , n1792);
  and g3483 (n2344, \in2[28] , n_1854);
  not g3484 (n_2294, n2343);
  not g3485 (n_2295, n2344);
  and g3486 (n2345, n_2294, n_2295);
  not g3487 (n_2296, n2345);
  and g3488 (n2346, n2342, n_2296);
  and g3489 (n2347, \in1[27] , n1787);
  and g3490 (n2348, \in0[27] , n_1849);
  not g3491 (n_2297, n2347);
  not g3492 (n_2298, n2348);
  and g3493 (n2349, n_2297, n_2298);
  and g3494 (n2350, \in3[27] , n1792);
  and g3495 (n2351, \in2[27] , n_1854);
  not g3496 (n_2299, n2350);
  not g3497 (n_2300, n2351);
  and g3498 (n2352, n_2299, n_2300);
  not g3499 (n_2301, n2352);
  and g3500 (n2353, n2349, n_2301);
  and g3501 (n2354, \in1[26] , n1787);
  and g3502 (n2355, \in0[26] , n_1849);
  not g3503 (n_2302, n2354);
  not g3504 (n_2303, n2355);
  and g3505 (n2356, n_2302, n_2303);
  and g3506 (n2357, \in3[26] , n1792);
  and g3507 (n2358, \in2[26] , n_1854);
  not g3508 (n_2304, n2357);
  not g3509 (n_2305, n2358);
  and g3510 (n2359, n_2304, n_2305);
  not g3511 (n_2306, n2359);
  and g3512 (n2360, n2356, n_2306);
  and g3513 (n2361, \in3[25] , n1792);
  and g3514 (n2362, \in2[25] , n_1854);
  not g3515 (n_2307, n2361);
  not g3516 (n_2308, n2362);
  and g3517 (n2363, n_2307, n_2308);
  and g3518 (n2364, \in3[24] , n1792);
  and g3519 (n2365, \in2[24] , n_1854);
  not g3520 (n_2309, n2364);
  not g3521 (n_2310, n2365);
  and g3522 (n2366, n_2309, n_2310);
  and g3523 (n2367, \in1[23] , n1787);
  and g3524 (n2368, \in0[23] , n_1849);
  not g3525 (n_2311, n2367);
  not g3526 (n_2312, n2368);
  and g3527 (n2369, n_2311, n_2312);
  and g3528 (n2370, \in3[23] , n1792);
  and g3529 (n2371, \in2[23] , n_1854);
  not g3530 (n_2313, n2370);
  not g3531 (n_2314, n2371);
  and g3532 (n2372, n_2313, n_2314);
  not g3533 (n_2315, n2372);
  and g3534 (n2373, n2369, n_2315);
  and g3535 (n2374, \in1[22] , n1787);
  and g3536 (n2375, \in0[22] , n_1849);
  not g3537 (n_2316, n2374);
  not g3538 (n_2317, n2375);
  and g3539 (n2376, n_2316, n_2317);
  and g3540 (n2377, \in3[22] , n1792);
  and g3541 (n2378, \in2[22] , n_1854);
  not g3542 (n_2318, n2377);
  not g3543 (n_2319, n2378);
  and g3544 (n2379, n_2318, n_2319);
  not g3545 (n_2320, n2379);
  and g3546 (n2380, n2376, n_2320);
  and g3547 (n2381, \in1[21] , n1787);
  and g3548 (n2382, \in0[21] , n_1849);
  not g3549 (n_2321, n2381);
  not g3550 (n_2322, n2382);
  and g3551 (n2383, n_2321, n_2322);
  and g3552 (n2384, \in3[21] , n1792);
  and g3553 (n2385, \in2[21] , n_1854);
  not g3554 (n_2323, n2384);
  not g3555 (n_2324, n2385);
  and g3556 (n2386, n_2323, n_2324);
  not g3557 (n_2325, n2386);
  and g3558 (n2387, n2383, n_2325);
  and g3559 (n2388, \in1[20] , n1787);
  and g3560 (n2389, \in0[20] , n_1849);
  not g3561 (n_2326, n2388);
  not g3562 (n_2327, n2389);
  and g3563 (n2390, n_2326, n_2327);
  and g3564 (n2391, \in3[20] , n1792);
  and g3565 (n2392, \in2[20] , n_1854);
  not g3566 (n_2328, n2391);
  not g3567 (n_2329, n2392);
  and g3568 (n2393, n_2328, n_2329);
  not g3569 (n_2330, n2393);
  and g3570 (n2394, n2390, n_2330);
  and g3571 (n2395, \in1[19] , n1787);
  and g3572 (n2396, \in0[19] , n_1849);
  not g3573 (n_2331, n2395);
  not g3574 (n_2332, n2396);
  and g3575 (n2397, n_2331, n_2332);
  and g3576 (n2398, \in3[19] , n1792);
  and g3577 (n2399, \in2[19] , n_1854);
  not g3578 (n_2333, n2398);
  not g3579 (n_2334, n2399);
  and g3580 (n2400, n_2333, n_2334);
  not g3581 (n_2335, n2400);
  and g3582 (n2401, n2397, n_2335);
  and g3583 (n2402, \in1[18] , n1787);
  and g3584 (n2403, \in0[18] , n_1849);
  not g3585 (n_2336, n2402);
  not g3586 (n_2337, n2403);
  and g3587 (n2404, n_2336, n_2337);
  and g3588 (n2405, \in3[18] , n1792);
  and g3589 (n2406, \in2[18] , n_1854);
  not g3590 (n_2338, n2405);
  not g3591 (n_2339, n2406);
  and g3592 (n2407, n_2338, n_2339);
  not g3593 (n_2340, n2407);
  and g3594 (n2408, n2404, n_2340);
  and g3595 (n2409, \in3[17] , n1792);
  and g3596 (n2410, \in2[17] , n_1854);
  not g3597 (n_2341, n2409);
  not g3598 (n_2342, n2410);
  and g3599 (n2411, n_2341, n_2342);
  and g3600 (n2412, \in3[16] , n1792);
  and g3601 (n2413, \in2[16] , n_1854);
  not g3602 (n_2343, n2412);
  not g3603 (n_2344, n2413);
  and g3604 (n2414, n_2343, n_2344);
  and g3605 (n2415, \in1[15] , n1787);
  and g3606 (n2416, \in0[15] , n_1849);
  not g3607 (n_2345, n2415);
  not g3608 (n_2346, n2416);
  and g3609 (n2417, n_2345, n_2346);
  and g3610 (n2418, \in3[15] , n1792);
  and g3611 (n2419, \in2[15] , n_1854);
  not g3612 (n_2347, n2418);
  not g3613 (n_2348, n2419);
  and g3614 (n2420, n_2347, n_2348);
  not g3615 (n_2349, n2420);
  and g3616 (n2421, n2417, n_2349);
  and g3617 (n2422, \in1[14] , n1787);
  and g3618 (n2423, \in0[14] , n_1849);
  not g3619 (n_2350, n2422);
  not g3620 (n_2351, n2423);
  and g3621 (n2424, n_2350, n_2351);
  and g3622 (n2425, \in3[14] , n1792);
  and g3623 (n2426, \in2[14] , n_1854);
  not g3624 (n_2352, n2425);
  not g3625 (n_2353, n2426);
  and g3626 (n2427, n_2352, n_2353);
  not g3627 (n_2354, n2427);
  and g3628 (n2428, n2424, n_2354);
  and g3629 (n2429, \in1[13] , n1787);
  and g3630 (n2430, \in0[13] , n_1849);
  not g3631 (n_2355, n2429);
  not g3632 (n_2356, n2430);
  and g3633 (n2431, n_2355, n_2356);
  and g3634 (n2432, \in3[13] , n1792);
  and g3635 (n2433, \in2[13] , n_1854);
  not g3636 (n_2357, n2432);
  not g3637 (n_2358, n2433);
  and g3638 (n2434, n_2357, n_2358);
  not g3639 (n_2359, n2434);
  and g3640 (n2435, n2431, n_2359);
  and g3641 (n2436, \in1[12] , n1787);
  and g3642 (n2437, \in0[12] , n_1849);
  not g3643 (n_2360, n2436);
  not g3644 (n_2361, n2437);
  and g3645 (n2438, n_2360, n_2361);
  and g3646 (n2439, \in3[12] , n1792);
  and g3647 (n2440, \in2[12] , n_1854);
  not g3648 (n_2362, n2439);
  not g3649 (n_2363, n2440);
  and g3650 (n2441, n_2362, n_2363);
  not g3651 (n_2364, n2441);
  and g3652 (n2442, n2438, n_2364);
  and g3653 (n2443, \in1[11] , n1787);
  and g3654 (n2444, \in0[11] , n_1849);
  not g3655 (n_2365, n2443);
  not g3656 (n_2366, n2444);
  and g3657 (n2445, n_2365, n_2366);
  and g3658 (n2446, \in3[11] , n1792);
  and g3659 (n2447, \in2[11] , n_1854);
  not g3660 (n_2367, n2446);
  not g3661 (n_2368, n2447);
  and g3662 (n2448, n_2367, n_2368);
  not g3663 (n_2369, n2448);
  and g3664 (n2449, n2445, n_2369);
  and g3665 (n2450, \in1[10] , n1787);
  and g3666 (n2451, \in0[10] , n_1849);
  not g3667 (n_2370, n2450);
  not g3668 (n_2371, n2451);
  and g3669 (n2452, n_2370, n_2371);
  and g3670 (n2453, \in3[10] , n1792);
  and g3671 (n2454, \in2[10] , n_1854);
  not g3672 (n_2372, n2453);
  not g3673 (n_2373, n2454);
  and g3674 (n2455, n_2372, n_2373);
  not g3675 (n_2374, n2455);
  and g3676 (n2456, n2452, n_2374);
  and g3677 (n2457, \in3[9] , n1792);
  and g3678 (n2458, \in2[9] , n_1854);
  not g3679 (n_2375, n2457);
  not g3680 (n_2376, n2458);
  and g3681 (n2459, n_2375, n_2376);
  and g3682 (n2460, \in3[8] , n1792);
  and g3683 (n2461, \in2[8] , n_1854);
  not g3684 (n_2377, n2460);
  not g3685 (n_2378, n2461);
  and g3686 (n2462, n_2377, n_2378);
  and g3687 (n2463, \in1[7] , n1787);
  and g3688 (n2464, \in0[7] , n_1849);
  not g3689 (n_2379, n2463);
  not g3690 (n_2380, n2464);
  and g3691 (n2465, n_2379, n_2380);
  and g3692 (n2466, \in3[7] , n1792);
  and g3693 (n2467, \in2[7] , n_1854);
  not g3694 (n_2381, n2466);
  not g3695 (n_2382, n2467);
  and g3696 (n2468, n_2381, n_2382);
  not g3697 (n_2383, n2468);
  and g3698 (n2469, n2465, n_2383);
  and g3699 (n2470, \in3[6] , n1792);
  and g3700 (n2471, \in2[6] , n_1854);
  not g3701 (n_2384, n2470);
  not g3702 (n_2385, n2471);
  and g3703 (n2472, n_2384, n_2385);
  and g3704 (n2473, \in1[6] , n1787);
  and g3705 (n2474, \in0[6] , n_1849);
  not g3706 (n_2386, n2473);
  not g3707 (n_2387, n2474);
  and g3708 (n2475, n_2386, n_2387);
  and g3709 (n2476, \in3[5] , n1792);
  and g3710 (n2477, \in2[5] , n_1854);
  not g3711 (n_2388, n2476);
  not g3712 (n_2389, n2477);
  and g3713 (n2478, n_2388, n_2389);
  and g3714 (n2479, \in1[5] , n1787);
  and g3715 (n2480, \in0[5] , n_1849);
  not g3716 (n_2390, n2479);
  not g3717 (n_2391, n2480);
  and g3718 (n2481, n_2390, n_2391);
  and g3719 (n2482, \in3[4] , n1792);
  and g3720 (n2483, \in2[4] , n_1854);
  not g3721 (n_2392, n2482);
  not g3722 (n_2393, n2483);
  and g3723 (n2484, n_2392, n_2393);
  and g3724 (n2485, \in1[4] , n1787);
  and g3725 (n2486, \in0[4] , n_1849);
  not g3726 (n_2394, n2485);
  not g3727 (n_2395, n2486);
  and g3728 (n2487, n_2394, n_2395);
  and g3729 (n2488, \in1[3] , n1787);
  and g3730 (n2489, \in0[3] , n_1849);
  not g3731 (n_2396, n2488);
  not g3732 (n_2397, n2489);
  and g3733 (n2490, n_2396, n_2397);
  and g3734 (n2491, \in3[3] , n1792);
  and g3735 (n2492, \in2[3] , n_1854);
  not g3736 (n_2398, n2491);
  not g3737 (n_2399, n2492);
  and g3738 (n2493, n_2398, n_2399);
  not g3739 (n_2400, n2493);
  and g3740 (n2494, n2490, n_2400);
  and g3741 (n2495, \in3[1] , n1792);
  and g3742 (n2496, \in2[1] , n_1854);
  not g3743 (n_2401, n2495);
  not g3744 (n_2402, n2496);
  and g3745 (n2497, n_2401, n_2402);
  and g3746 (n2498, \in1[0] , n1787);
  and g3747 (n2499, \in0[0] , n_1849);
  not g3748 (n_2403, n2498);
  not g3749 (n_2404, n2499);
  and g3750 (n2500, n_2403, n_2404);
  and g3751 (n2501, \in3[0] , n1792);
  and g3752 (n2502, \in2[0] , n_1854);
  not g3753 (n_2405, n2501);
  not g3754 (n_2406, n2502);
  and g3755 (n2503, n_2405, n_2406);
  not g3756 (n_2407, n2500);
  and g3757 (n2504, n_2407, n2503);
  and g3758 (n2505, n2497, n2504);
  and g3759 (n2506, \in1[1] , n1787);
  and g3760 (n2507, \in0[1] , n_1849);
  not g3761 (n_2408, n2506);
  not g3762 (n_2409, n2507);
  and g3763 (n2508, n_2408, n_2409);
  not g3764 (n_2410, n2505);
  and g3765 (n2509, n_2410, n2508);
  and g3766 (n2510, \in1[2] , n1787);
  and g3767 (n2511, \in0[2] , n_1849);
  not g3768 (n_2411, n2510);
  not g3769 (n_2412, n2511);
  and g3770 (n2512, n_2411, n_2412);
  and g3771 (n2513, \in3[2] , n1792);
  and g3772 (n2514, \in2[2] , n_1854);
  not g3773 (n_2413, n2513);
  not g3774 (n_2414, n2514);
  and g3775 (n2515, n_2413, n_2414);
  not g3776 (n_2415, n2515);
  and g3777 (n2516, n2512, n_2415);
  not g3778 (n_2416, n2497);
  not g3779 (n_2417, n2504);
  and g3780 (n2517, n_2416, n_2417);
  not g3781 (n_2418, n2516);
  not g3782 (n_2419, n2517);
  and g3783 (n2518, n_2418, n_2419);
  not g3784 (n_2420, n2509);
  and g3785 (n2519, n_2420, n2518);
  not g3786 (n_2421, n2512);
  and g3787 (n2520, n_2421, n2515);
  not g3788 (n_2422, n2519);
  not g3789 (n_2423, n2520);
  and g3790 (n2521, n_2422, n_2423);
  not g3791 (n_2424, n2494);
  not g3792 (n_2425, n2521);
  and g3793 (n2522, n_2424, n_2425);
  not g3794 (n_2426, n2490);
  and g3795 (n2523, n_2426, n2493);
  not g3796 (n_2427, n2522);
  not g3797 (n_2428, n2523);
  and g3798 (n2524, n_2427, n_2428);
  and g3799 (n2525, n2487, n2524);
  not g3800 (n_2429, n2525);
  and g3801 (n2526, n2484, n_2429);
  not g3802 (n_2430, n2487);
  not g3803 (n_2431, n2524);
  and g3804 (n2527, n_2430, n_2431);
  not g3805 (n_2432, n2526);
  not g3806 (n_2433, n2527);
  and g3807 (n2528, n_2432, n_2433);
  and g3808 (n2529, n2481, n2528);
  not g3809 (n_2434, n2529);
  and g3810 (n2530, n2478, n_2434);
  not g3811 (n_2435, n2481);
  not g3812 (n_2436, n2528);
  and g3813 (n2531, n_2435, n_2436);
  not g3814 (n_2437, n2530);
  not g3815 (n_2438, n2531);
  and g3816 (n2532, n_2437, n_2438);
  and g3817 (n2533, n2475, n2532);
  not g3818 (n_2439, n2533);
  and g3819 (n2534, n2472, n_2439);
  not g3820 (n_2440, n2475);
  not g3821 (n_2441, n2532);
  and g3822 (n2535, n_2440, n_2441);
  not g3823 (n_2442, n2534);
  not g3824 (n_2443, n2535);
  and g3825 (n2536, n_2442, n_2443);
  not g3826 (n_2444, n2469);
  not g3827 (n_2445, n2536);
  and g3828 (n2537, n_2444, n_2445);
  not g3829 (n_2446, n2465);
  and g3830 (n2538, n_2446, n2468);
  not g3831 (n_2447, n2537);
  not g3832 (n_2448, n2538);
  and g3833 (n2539, n_2447, n_2448);
  and g3834 (n2540, \in1[8] , n1787);
  and g3835 (n2541, \in0[8] , n_1849);
  not g3836 (n_2449, n2540);
  not g3837 (n_2450, n2541);
  and g3838 (n2542, n_2449, n_2450);
  and g3839 (n2543, n2539, n2542);
  not g3840 (n_2451, n2543);
  and g3841 (n2544, n2462, n_2451);
  not g3842 (n_2452, n2539);
  not g3843 (n_2453, n2542);
  and g3844 (n2545, n_2452, n_2453);
  not g3845 (n_2454, n2544);
  not g3846 (n_2455, n2545);
  and g3847 (n2546, n_2454, n_2455);
  and g3848 (n2547, \in1[9] , n1787);
  and g3849 (n2548, \in0[9] , n_1849);
  not g3850 (n_2456, n2547);
  not g3851 (n_2457, n2548);
  and g3852 (n2549, n_2456, n_2457);
  and g3853 (n2550, n2546, n2549);
  not g3854 (n_2458, n2550);
  and g3855 (n2551, n2459, n_2458);
  not g3856 (n_2459, n2546);
  not g3857 (n_2460, n2549);
  and g3858 (n2552, n_2459, n_2460);
  not g3859 (n_2461, n2551);
  not g3860 (n_2462, n2552);
  and g3861 (n2553, n_2461, n_2462);
  not g3862 (n_2463, n2456);
  not g3863 (n_2464, n2553);
  and g3864 (n2554, n_2463, n_2464);
  not g3865 (n_2465, n2452);
  and g3866 (n2555, n_2465, n2455);
  not g3867 (n_2466, n2554);
  not g3868 (n_2467, n2555);
  and g3869 (n2556, n_2466, n_2467);
  not g3870 (n_2468, n2449);
  not g3871 (n_2469, n2556);
  and g3872 (n2557, n_2468, n_2469);
  not g3873 (n_2470, n2445);
  and g3874 (n2558, n_2470, n2448);
  not g3875 (n_2471, n2557);
  not g3876 (n_2472, n2558);
  and g3877 (n2559, n_2471, n_2472);
  not g3878 (n_2473, n2442);
  not g3879 (n_2474, n2559);
  and g3880 (n2560, n_2473, n_2474);
  not g3881 (n_2475, n2438);
  and g3882 (n2561, n_2475, n2441);
  not g3883 (n_2476, n2560);
  not g3884 (n_2477, n2561);
  and g3885 (n2562, n_2476, n_2477);
  not g3886 (n_2478, n2435);
  not g3887 (n_2479, n2562);
  and g3888 (n2563, n_2478, n_2479);
  not g3889 (n_2480, n2431);
  and g3890 (n2564, n_2480, n2434);
  not g3891 (n_2481, n2563);
  not g3892 (n_2482, n2564);
  and g3893 (n2565, n_2481, n_2482);
  not g3894 (n_2483, n2428);
  not g3895 (n_2484, n2565);
  and g3896 (n2566, n_2483, n_2484);
  not g3897 (n_2485, n2424);
  and g3898 (n2567, n_2485, n2427);
  not g3899 (n_2486, n2566);
  not g3900 (n_2487, n2567);
  and g3901 (n2568, n_2486, n_2487);
  not g3902 (n_2488, n2421);
  not g3903 (n_2489, n2568);
  and g3904 (n2569, n_2488, n_2489);
  not g3905 (n_2490, n2417);
  and g3906 (n2570, n_2490, n2420);
  not g3907 (n_2491, n2569);
  not g3908 (n_2492, n2570);
  and g3909 (n2571, n_2491, n_2492);
  and g3910 (n2572, \in1[16] , n1787);
  and g3911 (n2573, \in0[16] , n_1849);
  not g3912 (n_2493, n2572);
  not g3913 (n_2494, n2573);
  and g3914 (n2574, n_2493, n_2494);
  and g3915 (n2575, n2571, n2574);
  not g3916 (n_2495, n2575);
  and g3917 (n2576, n2414, n_2495);
  not g3918 (n_2496, n2571);
  not g3919 (n_2497, n2574);
  and g3920 (n2577, n_2496, n_2497);
  not g3921 (n_2498, n2576);
  not g3922 (n_2499, n2577);
  and g3923 (n2578, n_2498, n_2499);
  and g3924 (n2579, \in1[17] , n1787);
  and g3925 (n2580, \in0[17] , n_1849);
  not g3926 (n_2500, n2579);
  not g3927 (n_2501, n2580);
  and g3928 (n2581, n_2500, n_2501);
  and g3929 (n2582, n2578, n2581);
  not g3930 (n_2502, n2582);
  and g3931 (n2583, n2411, n_2502);
  not g3932 (n_2503, n2578);
  not g3933 (n_2504, n2581);
  and g3934 (n2584, n_2503, n_2504);
  not g3935 (n_2505, n2583);
  not g3936 (n_2506, n2584);
  and g3937 (n2585, n_2505, n_2506);
  not g3938 (n_2507, n2408);
  not g3939 (n_2508, n2585);
  and g3940 (n2586, n_2507, n_2508);
  not g3941 (n_2509, n2404);
  and g3942 (n2587, n_2509, n2407);
  not g3943 (n_2510, n2586);
  not g3944 (n_2511, n2587);
  and g3945 (n2588, n_2510, n_2511);
  not g3946 (n_2512, n2401);
  not g3947 (n_2513, n2588);
  and g3948 (n2589, n_2512, n_2513);
  not g3949 (n_2514, n2397);
  and g3950 (n2590, n_2514, n2400);
  not g3951 (n_2515, n2589);
  not g3952 (n_2516, n2590);
  and g3953 (n2591, n_2515, n_2516);
  not g3954 (n_2517, n2394);
  not g3955 (n_2518, n2591);
  and g3956 (n2592, n_2517, n_2518);
  not g3957 (n_2519, n2390);
  and g3958 (n2593, n_2519, n2393);
  not g3959 (n_2520, n2592);
  not g3960 (n_2521, n2593);
  and g3961 (n2594, n_2520, n_2521);
  not g3962 (n_2522, n2387);
  not g3963 (n_2523, n2594);
  and g3964 (n2595, n_2522, n_2523);
  not g3965 (n_2524, n2383);
  and g3966 (n2596, n_2524, n2386);
  not g3967 (n_2525, n2595);
  not g3968 (n_2526, n2596);
  and g3969 (n2597, n_2525, n_2526);
  not g3970 (n_2527, n2380);
  not g3971 (n_2528, n2597);
  and g3972 (n2598, n_2527, n_2528);
  not g3973 (n_2529, n2376);
  and g3974 (n2599, n_2529, n2379);
  not g3975 (n_2530, n2598);
  not g3976 (n_2531, n2599);
  and g3977 (n2600, n_2530, n_2531);
  not g3978 (n_2532, n2373);
  not g3979 (n_2533, n2600);
  and g3980 (n2601, n_2532, n_2533);
  not g3981 (n_2534, n2369);
  and g3982 (n2602, n_2534, n2372);
  not g3983 (n_2535, n2601);
  not g3984 (n_2536, n2602);
  and g3985 (n2603, n_2535, n_2536);
  and g3986 (n2604, \in1[24] , n1787);
  and g3987 (n2605, \in0[24] , n_1849);
  not g3988 (n_2537, n2604);
  not g3989 (n_2538, n2605);
  and g3990 (n2606, n_2537, n_2538);
  and g3991 (n2607, n2603, n2606);
  not g3992 (n_2539, n2607);
  and g3993 (n2608, n2366, n_2539);
  not g3994 (n_2540, n2603);
  not g3995 (n_2541, n2606);
  and g3996 (n2609, n_2540, n_2541);
  not g3997 (n_2542, n2608);
  not g3998 (n_2543, n2609);
  and g3999 (n2610, n_2542, n_2543);
  and g4000 (n2611, \in1[25] , n1787);
  and g4001 (n2612, \in0[25] , n_1849);
  not g4002 (n_2544, n2611);
  not g4003 (n_2545, n2612);
  and g4004 (n2613, n_2544, n_2545);
  and g4005 (n2614, n2610, n2613);
  not g4006 (n_2546, n2614);
  and g4007 (n2615, n2363, n_2546);
  not g4008 (n_2547, n2610);
  not g4009 (n_2548, n2613);
  and g4010 (n2616, n_2547, n_2548);
  not g4011 (n_2549, n2615);
  not g4012 (n_2550, n2616);
  and g4013 (n2617, n_2549, n_2550);
  not g4014 (n_2551, n2360);
  not g4015 (n_2552, n2617);
  and g4016 (n2618, n_2551, n_2552);
  not g4017 (n_2553, n2356);
  and g4018 (n2619, n_2553, n2359);
  not g4019 (n_2554, n2618);
  not g4020 (n_2555, n2619);
  and g4021 (n2620, n_2554, n_2555);
  not g4022 (n_2556, n2353);
  not g4023 (n_2557, n2620);
  and g4024 (n2621, n_2556, n_2557);
  not g4025 (n_2558, n2349);
  and g4026 (n2622, n_2558, n2352);
  not g4027 (n_2559, n2621);
  not g4028 (n_2560, n2622);
  and g4029 (n2623, n_2559, n_2560);
  not g4030 (n_2561, n2346);
  not g4031 (n_2562, n2623);
  and g4032 (n2624, n_2561, n_2562);
  not g4033 (n_2563, n2342);
  and g4034 (n2625, n_2563, n2345);
  not g4035 (n_2564, n2624);
  not g4036 (n_2565, n2625);
  and g4037 (n2626, n_2564, n_2565);
  not g4038 (n_2566, n2339);
  not g4039 (n_2567, n2626);
  and g4040 (n2627, n_2566, n_2567);
  not g4041 (n_2568, n2335);
  and g4042 (n2628, n_2568, n2338);
  not g4043 (n_2569, n2627);
  not g4044 (n_2570, n2628);
  and g4045 (n2629, n_2569, n_2570);
  not g4046 (n_2571, n2332);
  not g4047 (n_2572, n2629);
  and g4048 (n2630, n_2571, n_2572);
  not g4049 (n_2573, n2328);
  and g4050 (n2631, n_2573, n2331);
  not g4051 (n_2574, n2630);
  not g4052 (n_2575, n2631);
  and g4053 (n2632, n_2574, n_2575);
  not g4054 (n_2576, n2325);
  not g4055 (n_2577, n2632);
  and g4056 (n2633, n_2576, n_2577);
  not g4057 (n_2578, n2321);
  and g4058 (n2634, n_2578, n2324);
  not g4059 (n_2579, n2633);
  not g4060 (n_2580, n2634);
  and g4061 (n2635, n_2579, n_2580);
  and g4062 (n2636, \in1[39] , n1787);
  and g4063 (n2637, \in0[39] , n_1849);
  not g4064 (n_2581, n2636);
  not g4065 (n_2582, n2637);
  and g4066 (n2638, n_2581, n_2582);
  and g4067 (n2639, \in3[39] , n1792);
  and g4068 (n2640, \in2[39] , n_1854);
  not g4069 (n_2583, n2639);
  not g4070 (n_2584, n2640);
  and g4071 (n2641, n_2583, n_2584);
  not g4072 (n_2585, n2641);
  and g4073 (n2642, n2638, n_2585);
  and g4074 (n2643, \in3[38] , n1792);
  and g4075 (n2644, \in2[38] , n_1854);
  not g4076 (n_2586, n2643);
  not g4077 (n_2587, n2644);
  and g4078 (n2645, n_2586, n_2587);
  and g4079 (n2646, \in1[38] , n1787);
  and g4080 (n2647, \in0[38] , n_1849);
  not g4081 (n_2588, n2646);
  not g4082 (n_2589, n2647);
  and g4083 (n2648, n_2588, n_2589);
  not g4084 (n_2590, n2645);
  and g4085 (n2649, n_2590, n2648);
  not g4086 (n_2591, n2642);
  not g4087 (n_2592, n2649);
  and g4088 (n2650, n_2591, n_2592);
  and g4089 (n2651, \in1[36] , n1787);
  and g4090 (n2652, \in0[36] , n_1849);
  not g4091 (n_2593, n2651);
  not g4092 (n_2594, n2652);
  and g4093 (n2653, n_2593, n_2594);
  and g4094 (n2654, \in3[36] , n1792);
  and g4095 (n2655, \in2[36] , n_1854);
  not g4096 (n_2595, n2654);
  not g4097 (n_2596, n2655);
  and g4098 (n2656, n_2595, n_2596);
  not g4099 (n_2597, n2656);
  and g4100 (n2657, n2653, n_2597);
  and g4101 (n2658, \in1[37] , n1787);
  and g4102 (n2659, \in0[37] , n_1849);
  not g4103 (n_2598, n2658);
  not g4104 (n_2599, n2659);
  and g4105 (n2660, n_2598, n_2599);
  and g4106 (n2661, \in3[37] , n1792);
  and g4107 (n2662, \in2[37] , n_1854);
  not g4108 (n_2600, n2661);
  not g4109 (n_2601, n2662);
  and g4110 (n2663, n_2600, n_2601);
  not g4111 (n_2602, n2663);
  and g4112 (n2664, n2660, n_2602);
  not g4113 (n_2603, n2657);
  not g4114 (n_2604, n2664);
  and g4115 (n2665, n_2603, n_2604);
  and g4116 (n2666, n2650, n2665);
  and g4117 (n2667, \in1[33] , n1787);
  and g4118 (n2668, \in0[33] , n_1849);
  not g4119 (n_2605, n2667);
  not g4120 (n_2606, n2668);
  and g4121 (n2669, n_2605, n_2606);
  and g4122 (n2670, \in3[33] , n1792);
  and g4123 (n2671, \in2[33] , n_1854);
  not g4124 (n_2607, n2670);
  not g4125 (n_2608, n2671);
  and g4126 (n2672, n_2607, n_2608);
  not g4127 (n_2609, n2672);
  and g4128 (n2673, n2669, n_2609);
  and g4129 (n2674, \in1[35] , n1787);
  and g4130 (n2675, \in0[35] , n_1849);
  not g4131 (n_2610, n2674);
  not g4132 (n_2611, n2675);
  and g4133 (n2676, n_2610, n_2611);
  and g4134 (n2677, \in3[35] , n1792);
  and g4135 (n2678, \in2[35] , n_1854);
  not g4136 (n_2612, n2677);
  not g4137 (n_2613, n2678);
  and g4138 (n2679, n_2612, n_2613);
  not g4139 (n_2614, n2679);
  and g4140 (n2680, n2676, n_2614);
  and g4141 (n2681, \in3[34] , n1792);
  and g4142 (n2682, \in2[34] , n_1854);
  not g4143 (n_2615, n2681);
  not g4144 (n_2616, n2682);
  and g4145 (n2683, n_2615, n_2616);
  and g4146 (n2684, \in1[34] , n1787);
  and g4147 (n2685, \in0[34] , n_1849);
  not g4148 (n_2617, n2684);
  not g4149 (n_2618, n2685);
  and g4150 (n2686, n_2617, n_2618);
  not g4151 (n_2619, n2683);
  and g4152 (n2687, n_2619, n2686);
  not g4153 (n_2620, n2680);
  not g4154 (n_2621, n2687);
  and g4155 (n2688, n_2620, n_2621);
  not g4156 (n_2622, n2673);
  and g4157 (n2689, n_2622, n2688);
  not g4163 (n_2625, n2638);
  and g4164 (n2693, n_2625, n2641);
  not g4165 (n_2626, n2653);
  and g4166 (n2694, n_2626, n2656);
  and g4167 (n2695, n_2604, n2694);
  not g4168 (n_2627, n2660);
  and g4169 (n2696, n_2627, n2663);
  not g4170 (n_2628, n2695);
  not g4171 (n_2629, n2696);
  and g4172 (n2697, n_2628, n_2629);
  not g4173 (n_2630, n2697);
  and g4174 (n2698, n2650, n_2630);
  and g4175 (n2699, n_2591, n2645);
  not g4176 (n_2631, n2648);
  and g4177 (n2700, n_2631, n2699);
  not g4178 (n_2632, n2676);
  and g4179 (n2701, n_2632, n2679);
  and g4180 (n2702, n_2620, n2683);
  not g4181 (n_2633, n2686);
  and g4182 (n2703, n_2633, n2702);
  not g4183 (n_2634, n2317);
  and g4184 (n2704, n2314, n_2634);
  not g4185 (n_2635, n2669);
  and g4186 (n2705, n_2635, n2672);
  not g4187 (n_2636, n2704);
  not g4188 (n_2637, n2705);
  and g4189 (n2706, n_2636, n_2637);
  not g4190 (n_2638, n2706);
  and g4191 (n2707, n2689, n_2638);
  not g4192 (n_2639, n2703);
  not g4193 (n_2640, n2707);
  and g4194 (n2708, n_2639, n_2640);
  not g4195 (n_2641, n2701);
  and g4196 (n2709, n_2641, n2708);
  not g4197 (n_2642, n2709);
  and g4198 (n2710, n2666, n_2642);
  not g4208 (n_2648, n2295);
  and g4209 (n2715, n2292, n_2648);
  and g4225 (n2724, \in3[48] , n1792);
  and g4226 (n2725, \in2[48] , n_1854);
  not g4227 (n_2656, n2724);
  not g4228 (n_2657, n2725);
  and g4229 (n2726, n_2656, n_2657);
  and g4230 (n2727, \in1[48] , n1787);
  and g4231 (n2728, \in0[48] , n_1849);
  not g4232 (n_2658, n2727);
  not g4233 (n_2659, n2728);
  and g4234 (n2729, n_2658, n_2659);
  not g4235 (n_2660, n2726);
  and g4236 (n2730, n_2660, n2729);
  and g4237 (n2731, \in1[55] , n1787);
  and g4238 (n2732, \in0[55] , n_1849);
  not g4239 (n_2661, n2731);
  not g4240 (n_2662, n2732);
  and g4241 (n2733, n_2661, n_2662);
  and g4242 (n2734, \in3[55] , n1792);
  and g4243 (n2735, \in2[55] , n_1854);
  not g4244 (n_2663, n2734);
  not g4245 (n_2664, n2735);
  and g4246 (n2736, n_2663, n_2664);
  not g4247 (n_2665, n2736);
  and g4248 (n2737, n2733, n_2665);
  and g4249 (n2738, \in3[54] , n1792);
  and g4250 (n2739, \in2[54] , n_1854);
  not g4251 (n_2666, n2738);
  not g4252 (n_2667, n2739);
  and g4253 (n2740, n_2666, n_2667);
  and g4254 (n2741, \in1[54] , n1787);
  and g4255 (n2742, \in0[54] , n_1849);
  not g4256 (n_2668, n2741);
  not g4257 (n_2669, n2742);
  and g4258 (n2743, n_2668, n_2669);
  not g4259 (n_2670, n2740);
  and g4260 (n2744, n_2670, n2743);
  not g4261 (n_2671, n2737);
  not g4262 (n_2672, n2744);
  and g4263 (n2745, n_2671, n_2672);
  and g4264 (n2746, \in1[53] , n1787);
  and g4265 (n2747, \in0[53] , n_1849);
  not g4266 (n_2673, n2746);
  not g4267 (n_2674, n2747);
  and g4268 (n2748, n_2673, n_2674);
  and g4269 (n2749, \in3[53] , n1792);
  and g4270 (n2750, \in2[53] , n_1854);
  not g4271 (n_2675, n2749);
  not g4272 (n_2676, n2750);
  and g4273 (n2751, n_2675, n_2676);
  not g4274 (n_2677, n2751);
  and g4275 (n2752, n2748, n_2677);
  and g4276 (n2753, \in3[52] , n1792);
  and g4277 (n2754, \in2[52] , n_1854);
  not g4278 (n_2678, n2753);
  not g4279 (n_2679, n2754);
  and g4280 (n2755, n_2678, n_2679);
  and g4281 (n2756, \in1[52] , n1787);
  and g4282 (n2757, \in0[52] , n_1849);
  not g4283 (n_2680, n2756);
  not g4284 (n_2681, n2757);
  and g4285 (n2758, n_2680, n_2681);
  not g4286 (n_2682, n2755);
  and g4287 (n2759, n_2682, n2758);
  not g4288 (n_2683, n2752);
  not g4289 (n_2684, n2759);
  and g4290 (n2760, n_2683, n_2684);
  and g4291 (n2761, n2745, n2760);
  and g4292 (n2762, \in1[49] , n1787);
  and g4293 (n2763, \in0[49] , n_1849);
  not g4294 (n_2685, n2762);
  not g4295 (n_2686, n2763);
  and g4296 (n2764, n_2685, n_2686);
  and g4297 (n2765, \in3[49] , n1792);
  and g4298 (n2766, \in2[49] , n_1854);
  not g4299 (n_2687, n2765);
  not g4300 (n_2688, n2766);
  and g4301 (n2767, n_2687, n_2688);
  not g4302 (n_2689, n2767);
  and g4303 (n2768, n2764, n_2689);
  and g4304 (n2769, \in1[51] , n1787);
  and g4305 (n2770, \in0[51] , n_1849);
  not g4306 (n_2690, n2769);
  not g4307 (n_2691, n2770);
  and g4308 (n2771, n_2690, n_2691);
  and g4309 (n2772, \in3[51] , n1792);
  and g4310 (n2773, \in2[51] , n_1854);
  not g4311 (n_2692, n2772);
  not g4312 (n_2693, n2773);
  and g4313 (n2774, n_2692, n_2693);
  not g4314 (n_2694, n2774);
  and g4315 (n2775, n2771, n_2694);
  and g4316 (n2776, \in3[50] , n1792);
  and g4317 (n2777, \in2[50] , n_1854);
  not g4318 (n_2695, n2776);
  not g4319 (n_2696, n2777);
  and g4320 (n2778, n_2695, n_2696);
  and g4321 (n2779, \in1[50] , n1787);
  and g4322 (n2780, \in0[50] , n_1849);
  not g4323 (n_2697, n2779);
  not g4324 (n_2698, n2780);
  and g4325 (n2781, n_2697, n_2698);
  not g4326 (n_2699, n2778);
  and g4327 (n2782, n_2699, n2781);
  not g4328 (n_2700, n2775);
  not g4329 (n_2701, n2782);
  and g4330 (n2783, n_2700, n_2701);
  not g4331 (n_2702, n2768);
  and g4332 (n2784, n_2702, n2783);
  not g4338 (n_2705, n2733);
  and g4339 (n2788, n_2705, n2736);
  not g4340 (n_2706, n2771);
  and g4341 (n2789, n_2706, n2774);
  and g4342 (n2790, n_2700, n2778);
  not g4343 (n_2707, n2781);
  and g4344 (n2791, n_2707, n2790);
  not g4345 (n_2708, n2729);
  and g4346 (n2792, n2726, n_2708);
  not g4347 (n_2709, n2764);
  and g4348 (n2793, n_2709, n2767);
  not g4349 (n_2710, n2792);
  not g4350 (n_2711, n2793);
  and g4351 (n2794, n_2710, n_2711);
  not g4352 (n_2712, n2794);
  and g4353 (n2795, n2784, n_2712);
  not g4354 (n_2713, n2791);
  not g4355 (n_2714, n2795);
  and g4356 (n2796, n_2713, n_2714);
  not g4357 (n_2715, n2789);
  and g4358 (n2797, n_2715, n2796);
  not g4359 (n_2716, n2797);
  and g4360 (n2798, n2761, n_2716);
  not g4361 (n_2717, n2758);
  and g4362 (n2799, n2755, n_2717);
  and g4363 (n2800, n_2683, n2799);
  not g4364 (n_2718, n2748);
  and g4365 (n2801, n_2718, n2751);
  not g4366 (n_2719, n2800);
  not g4367 (n_2720, n2801);
  and g4368 (n2802, n_2719, n_2720);
  not g4369 (n_2721, n2743);
  and g4370 (n2803, n2740, n_2721);
  not g4371 (n_2722, n2803);
  and g4372 (n2804, n2802, n_2722);
  not g4373 (n_2723, n2804);
  and g4374 (n2805, n2745, n_2723);
  not g4382 (n_2728, n2218);
  and g4383 (n2809, n2215, n_2728);
  not g4399 (n_2736, n2157);
  not g4405 (n_2739, n2131);
  and g4406 (n2821, n_2739, n2134);
  and g4407 (n2822, n2146, n_2736);
  not g4408 (n_2740, n2149);
  and g4409 (n2823, n_2740, n2822);
  not g4410 (n_2741, n2153);
  and g4411 (n2824, n_2741, n2156);
  not g4412 (n_2742, n2823);
  not g4413 (n_2743, n2824);
  and g4414 (n2825, n_2742, n_2743);
  not g4415 (n_2744, n2141);
  and g4416 (n2826, n2138, n_2744);
  not g4417 (n_2745, n2826);
  and g4418 (n2827, n2825, n_2745);
  not g4419 (n_2746, n2827);
  and g4420 (n2828, n2143, n_2746);
  not g4421 (n_2747, n2821);
  not g4422 (n_2748, n2828);
  and g4423 (n2829, n_2747, n_2748);
  not g4424 (n_2749, n2820);
  and g4425 (n2830, n_2749, n2829);
  not g4426 (n_2750, n2121);
  and g4427 (n2831, n2118, n_2750);
  and g4440 (n2838, \in1[75] , n1787);
  and g4441 (n2839, \in0[75] , n_1849);
  not g4442 (n_2757, n2838);
  not g4443 (n_2758, n2839);
  and g4444 (n2840, n_2757, n_2758);
  and g4445 (n2841, \in3[75] , n1792);
  and g4446 (n2842, \in2[75] , n_1854);
  not g4447 (n_2759, n2841);
  not g4448 (n_2760, n2842);
  and g4449 (n2843, n_2759, n_2760);
  not g4450 (n_2761, n2843);
  and g4451 (n2844, n2840, n_2761);
  and g4452 (n2845, \in3[74] , n1792);
  and g4453 (n2846, \in2[74] , n_1854);
  not g4454 (n_2762, n2845);
  not g4455 (n_2763, n2846);
  and g4456 (n2847, n_2762, n_2763);
  and g4457 (n2848, \in1[74] , n1787);
  and g4458 (n2849, \in0[74] , n_1849);
  not g4459 (n_2764, n2848);
  not g4460 (n_2765, n2849);
  and g4461 (n2850, n_2764, n_2765);
  not g4462 (n_2766, n2847);
  and g4463 (n2851, n_2766, n2850);
  not g4464 (n_2767, n2844);
  not g4465 (n_2768, n2851);
  and g4466 (n2852, n_2767, n_2768);
  and g4467 (n2853, \in1[73] , n1787);
  and g4468 (n2854, \in0[73] , n_1849);
  not g4469 (n_2769, n2853);
  not g4470 (n_2770, n2854);
  and g4471 (n2855, n_2769, n_2770);
  and g4472 (n2856, \in3[73] , n1792);
  and g4473 (n2857, \in2[73] , n_1854);
  not g4474 (n_2771, n2856);
  not g4475 (n_2772, n2857);
  and g4476 (n2858, n_2771, n_2772);
  not g4477 (n_2773, n2858);
  and g4478 (n2859, n2855, n_2773);
  and g4479 (n2860, \in3[72] , n1792);
  and g4480 (n2861, \in2[72] , n_1854);
  not g4481 (n_2774, n2860);
  not g4482 (n_2775, n2861);
  and g4483 (n2862, n_2774, n_2775);
  and g4484 (n2863, \in1[72] , n1787);
  and g4485 (n2864, \in0[72] , n_1849);
  not g4486 (n_2776, n2863);
  not g4487 (n_2777, n2864);
  and g4488 (n2865, n_2776, n_2777);
  not g4489 (n_2778, n2862);
  and g4490 (n2866, n_2778, n2865);
  not g4491 (n_2779, n2859);
  not g4497 (n_2782, n2840);
  and g4498 (n2870, n_2782, n2843);
  not g4499 (n_2783, n2865);
  and g4500 (n2871, n2862, n_2783);
  and g4501 (n2872, n_2779, n2871);
  not g4502 (n_2784, n2855);
  and g4503 (n2873, n_2784, n2858);
  not g4504 (n_2785, n2872);
  not g4505 (n_2786, n2873);
  and g4506 (n2874, n_2785, n_2786);
  not g4507 (n_2787, n2850);
  and g4508 (n2875, n2847, n_2787);
  not g4509 (n_2788, n2875);
  and g4510 (n2876, n2874, n_2788);
  not g4511 (n_2789, n2876);
  and g4512 (n2877, n2852, n_2789);
  not g4513 (n_2790, n2870);
  not g4514 (n_2791, n2877);
  and g4515 (n2878, n_2790, n_2791);
  not g4516 (n_2792, n2869);
  and g4517 (n2879, n_2792, n2878);
  not g4518 (n_2793, n2085);
  and g4519 (n2880, n2082, n_2793);
  not g4532 (n_2800, n2056);
  not g4538 (n_2803, n2037);
  and g4539 (n2890, n_2803, n2040);
  and g4540 (n2891, n2030, n_2800);
  not g4541 (n_2804, n2033);
  and g4542 (n2892, n_2804, n2891);
  not g4543 (n_2805, n2052);
  and g4544 (n2893, n_2805, n2055);
  not g4545 (n_2806, n2892);
  not g4546 (n_2807, n2893);
  and g4547 (n2894, n_2806, n_2807);
  not g4548 (n_2808, n2047);
  and g4549 (n2895, n2044, n_2808);
  not g4550 (n_2809, n2895);
  and g4551 (n2896, n2894, n_2809);
  not g4552 (n_2810, n2896);
  and g4553 (n2897, n2049, n_2810);
  not g4554 (n_2811, n2890);
  not g4555 (n_2812, n2897);
  and g4556 (n2898, n_2811, n_2812);
  not g4557 (n_2813, n2889);
  and g4558 (n2899, n_2813, n2898);
  not g4559 (n_2814, n2020);
  and g4560 (n2900, n2017, n_2814);
  and g4573 (n2907, \in1[91] , n1787);
  and g4574 (n2908, \in0[91] , n_1849);
  not g4575 (n_2821, n2907);
  not g4576 (n_2822, n2908);
  and g4577 (n2909, n_2821, n_2822);
  and g4578 (n2910, \in3[91] , n1792);
  and g4579 (n2911, \in2[91] , n_1854);
  not g4580 (n_2823, n2910);
  not g4581 (n_2824, n2911);
  and g4582 (n2912, n_2823, n_2824);
  not g4583 (n_2825, n2912);
  and g4584 (n2913, n2909, n_2825);
  and g4585 (n2914, \in3[90] , n1792);
  and g4586 (n2915, \in2[90] , n_1854);
  not g4587 (n_2826, n2914);
  not g4588 (n_2827, n2915);
  and g4589 (n2916, n_2826, n_2827);
  and g4590 (n2917, \in1[90] , n1787);
  and g4591 (n2918, \in0[90] , n_1849);
  not g4592 (n_2828, n2917);
  not g4593 (n_2829, n2918);
  and g4594 (n2919, n_2828, n_2829);
  not g4595 (n_2830, n2916);
  and g4596 (n2920, n_2830, n2919);
  not g4597 (n_2831, n2913);
  not g4598 (n_2832, n2920);
  and g4599 (n2921, n_2831, n_2832);
  and g4600 (n2922, \in1[89] , n1787);
  and g4601 (n2923, \in0[89] , n_1849);
  not g4602 (n_2833, n2922);
  not g4603 (n_2834, n2923);
  and g4604 (n2924, n_2833, n_2834);
  and g4605 (n2925, \in3[89] , n1792);
  and g4606 (n2926, \in2[89] , n_1854);
  not g4607 (n_2835, n2925);
  not g4608 (n_2836, n2926);
  and g4609 (n2927, n_2835, n_2836);
  not g4610 (n_2837, n2927);
  and g4611 (n2928, n2924, n_2837);
  and g4612 (n2929, \in3[88] , n1792);
  and g4613 (n2930, \in2[88] , n_1854);
  not g4614 (n_2838, n2929);
  not g4615 (n_2839, n2930);
  and g4616 (n2931, n_2838, n_2839);
  and g4617 (n2932, \in1[88] , n1787);
  and g4618 (n2933, \in0[88] , n_1849);
  not g4619 (n_2840, n2932);
  not g4620 (n_2841, n2933);
  and g4621 (n2934, n_2840, n_2841);
  not g4622 (n_2842, n2931);
  and g4623 (n2935, n_2842, n2934);
  not g4624 (n_2843, n2928);
  not g4630 (n_2846, n2909);
  and g4631 (n2939, n_2846, n2912);
  not g4632 (n_2847, n2934);
  and g4633 (n2940, n2931, n_2847);
  and g4634 (n2941, n_2843, n2940);
  not g4635 (n_2848, n2924);
  and g4636 (n2942, n_2848, n2927);
  not g4637 (n_2849, n2941);
  not g4638 (n_2850, n2942);
  and g4639 (n2943, n_2849, n_2850);
  not g4640 (n_2851, n2919);
  and g4641 (n2944, n2916, n_2851);
  not g4642 (n_2852, n2944);
  and g4643 (n2945, n2943, n_2852);
  not g4644 (n_2853, n2945);
  and g4645 (n2946, n2921, n_2853);
  not g4646 (n_2854, n2939);
  not g4647 (n_2855, n2946);
  and g4648 (n2947, n_2854, n_2855);
  not g4649 (n_2856, n2938);
  and g4650 (n2948, n_2856, n2947);
  not g4651 (n_2857, n1984);
  and g4652 (n2949, n1981, n_2857);
  not g4665 (n_2864, n1955);
  not g4671 (n_2867, n1936);
  and g4672 (n2959, n_2867, n1939);
  and g4673 (n2960, n1929, n_2864);
  not g4674 (n_2868, n1932);
  and g4675 (n2961, n_2868, n2960);
  not g4676 (n_2869, n1951);
  and g4677 (n2962, n_2869, n1954);
  not g4678 (n_2870, n2961);
  not g4679 (n_2871, n2962);
  and g4680 (n2963, n_2870, n_2871);
  not g4681 (n_2872, n1946);
  and g4682 (n2964, n1943, n_2872);
  not g4683 (n_2873, n2964);
  and g4684 (n2965, n2963, n_2873);
  not g4685 (n_2874, n2965);
  and g4686 (n2966, n1948, n_2874);
  not g4687 (n_2875, n2959);
  not g4688 (n_2876, n2966);
  and g4689 (n2967, n_2875, n_2876);
  not g4690 (n_2877, n2958);
  and g4691 (n2968, n_2877, n2967);
  not g4692 (n_2878, n1919);
  and g4693 (n2969, n1916, n_2878);
  and g4706 (n2976, \in1[107] , n1787);
  and g4707 (n2977, \in0[107] , n_1849);
  not g4708 (n_2885, n2976);
  not g4709 (n_2886, n2977);
  and g4710 (n2978, n_2885, n_2886);
  and g4711 (n2979, \in3[107] , n1792);
  and g4712 (n2980, \in2[107] , n_1854);
  not g4713 (n_2887, n2979);
  not g4714 (n_2888, n2980);
  and g4715 (n2981, n_2887, n_2888);
  not g4716 (n_2889, n2981);
  and g4717 (n2982, n2978, n_2889);
  and g4718 (n2983, \in3[106] , n1792);
  and g4719 (n2984, \in2[106] , n_1854);
  not g4720 (n_2890, n2983);
  not g4721 (n_2891, n2984);
  and g4722 (n2985, n_2890, n_2891);
  and g4723 (n2986, \in1[106] , n1787);
  and g4724 (n2987, \in0[106] , n_1849);
  not g4725 (n_2892, n2986);
  not g4726 (n_2893, n2987);
  and g4727 (n2988, n_2892, n_2893);
  not g4728 (n_2894, n2985);
  and g4729 (n2989, n_2894, n2988);
  not g4730 (n_2895, n2982);
  not g4731 (n_2896, n2989);
  and g4732 (n2990, n_2895, n_2896);
  and g4733 (n2991, \in1[105] , n1787);
  and g4734 (n2992, \in0[105] , n_1849);
  not g4735 (n_2897, n2991);
  not g4736 (n_2898, n2992);
  and g4737 (n2993, n_2897, n_2898);
  and g4738 (n2994, \in3[105] , n1792);
  and g4739 (n2995, \in2[105] , n_1854);
  not g4740 (n_2899, n2994);
  not g4741 (n_2900, n2995);
  and g4742 (n2996, n_2899, n_2900);
  not g4743 (n_2901, n2996);
  and g4744 (n2997, n2993, n_2901);
  and g4745 (n2998, \in3[104] , n1792);
  and g4746 (n2999, \in2[104] , n_1854);
  not g4747 (n_2902, n2998);
  not g4748 (n_2903, n2999);
  and g4749 (n3000, n_2902, n_2903);
  and g4750 (n3001, \in1[104] , n1787);
  and g4751 (n3002, \in0[104] , n_1849);
  not g4752 (n_2904, n3001);
  not g4753 (n_2905, n3002);
  and g4754 (n3003, n_2904, n_2905);
  not g4755 (n_2906, n3000);
  and g4756 (n3004, n_2906, n3003);
  not g4757 (n_2907, n2997);
  not g4763 (n_2910, n2978);
  and g4764 (n3008, n_2910, n2981);
  not g4765 (n_2911, n3003);
  and g4766 (n3009, n3000, n_2911);
  and g4767 (n3010, n_2907, n3009);
  not g4768 (n_2912, n2993);
  and g4769 (n3011, n_2912, n2996);
  not g4770 (n_2913, n3010);
  not g4771 (n_2914, n3011);
  and g4772 (n3012, n_2913, n_2914);
  not g4773 (n_2915, n2988);
  and g4774 (n3013, n2985, n_2915);
  not g4775 (n_2916, n3013);
  and g4776 (n3014, n3012, n_2916);
  not g4777 (n_2917, n3014);
  and g4778 (n3015, n2990, n_2917);
  not g4779 (n_2918, n3008);
  not g4780 (n_2919, n3015);
  and g4781 (n3016, n_2918, n_2919);
  not g4782 (n_2920, n3007);
  and g4783 (n3017, n_2920, n3016);
  not g4784 (n_2921, n1883);
  and g4785 (n3018, n1880, n_2921);
  not g4798 (n_2928, n1854);
  not g4804 (n_2931, n1835);
  and g4805 (n3028, n_2931, n1838);
  and g4806 (n3029, n1828, n_2928);
  not g4807 (n_2932, n1831);
  and g4808 (n3030, n_2932, n3029);
  not g4809 (n_2933, n1850);
  and g4810 (n3031, n_2933, n1853);
  not g4811 (n_2934, n3030);
  not g4812 (n_2935, n3031);
  and g4813 (n3032, n_2934, n_2935);
  not g4814 (n_2936, n1845);
  and g4815 (n3033, n1842, n_2936);
  not g4816 (n_2937, n3033);
  and g4817 (n3034, n3032, n_2937);
  not g4818 (n_2938, n3034);
  and g4819 (n3035, n1847, n_2938);
  not g4820 (n_2939, n3028);
  not g4821 (n_2940, n3035);
  and g4822 (n3036, n_2939, n_2940);
  not g4823 (n_2941, n3027);
  and g4824 (n3037, n_2941, n3036);
  not g4825 (n_2942, n1818);
  and g4826 (n3038, n1808, n_2942);
  and g4839 (n3045, \in1[123] , n1787);
  and g4840 (n3046, \in0[123] , n_1849);
  not g4841 (n_2949, n3045);
  not g4842 (n_2950, n3046);
  and g4843 (n3047, n_2949, n_2950);
  and g4844 (n3048, \in3[123] , n1792);
  and g4845 (n3049, \in2[123] , n_1854);
  not g4846 (n_2951, n3048);
  not g4847 (n_2952, n3049);
  and g4848 (n3050, n_2951, n_2952);
  not g4849 (n_2953, n3050);
  and g4850 (n3051, n3047, n_2953);
  and g4851 (n3052, \in3[122] , n1792);
  and g4852 (n3053, \in2[122] , n_1854);
  not g4853 (n_2954, n3052);
  not g4854 (n_2955, n3053);
  and g4855 (n3054, n_2954, n_2955);
  and g4856 (n3055, \in1[122] , n1787);
  and g4857 (n3056, \in0[122] , n_1849);
  not g4858 (n_2956, n3055);
  not g4859 (n_2957, n3056);
  and g4860 (n3057, n_2956, n_2957);
  not g4861 (n_2958, n3054);
  and g4862 (n3058, n_2958, n3057);
  not g4863 (n_2959, n3051);
  not g4864 (n_2960, n3058);
  and g4865 (n3059, n_2959, n_2960);
  and g4866 (n3060, \in1[121] , n1787);
  and g4867 (n3061, \in0[121] , n_1849);
  not g4868 (n_2961, n3060);
  not g4869 (n_2962, n3061);
  and g4870 (n3062, n_2961, n_2962);
  and g4871 (n3063, \in3[121] , n1792);
  and g4872 (n3064, \in2[121] , n_1854);
  not g4873 (n_2963, n3063);
  not g4874 (n_2964, n3064);
  and g4875 (n3065, n_2963, n_2964);
  not g4876 (n_2965, n3065);
  and g4877 (n3066, n3062, n_2965);
  and g4878 (n3067, \in3[120] , n1792);
  and g4879 (n3068, \in2[120] , n_1854);
  not g4880 (n_2966, n3067);
  not g4881 (n_2967, n3068);
  and g4882 (n3069, n_2966, n_2967);
  and g4883 (n3070, \in1[120] , n1787);
  and g4884 (n3071, \in0[120] , n_1849);
  not g4885 (n_2968, n3070);
  not g4886 (n_2969, n3071);
  and g4887 (n3072, n_2968, n_2969);
  not g4888 (n_2970, n3069);
  and g4889 (n3073, n_2970, n3072);
  not g4890 (n_2971, n3066);
  not g4896 (n_2974, n3047);
  and g4897 (n3077, n_2974, n3050);
  and g4898 (n3078, n_2971, n3069);
  not g4899 (n_2975, n3072);
  and g4900 (n3079, n_2975, n3078);
  not g4901 (n_2976, n3062);
  and g4902 (n3080, n_2976, n3065);
  not g4903 (n_2977, n3079);
  not g4904 (n_2978, n3080);
  and g4905 (n3081, n_2977, n_2978);
  not g4906 (n_2979, n3057);
  and g4907 (n3082, n3054, n_2979);
  not g4908 (n_2980, n3082);
  and g4909 (n3083, n3081, n_2980);
  not g4910 (n_2981, n3083);
  and g4911 (n3084, n3059, n_2981);
  not g4912 (n_2982, n3077);
  not g4913 (n_2983, n3084);
  and g4914 (n3085, n_2982, n_2983);
  not g4915 (n_2984, n3076);
  and g4916 (n3086, n_2984, n3085);
  and g4917 (n3087, \in1[124] , n1787);
  and g4918 (n3088, \in0[124] , n_1849);
  not g4919 (n_2985, n3087);
  not g4920 (n_2986, n3088);
  and g4921 (n3089, n_2985, n_2986);
  and g4922 (n3090, \in3[124] , n1792);
  and g4923 (n3091, \in2[124] , n_1854);
  not g4924 (n_2987, n3090);
  not g4925 (n_2988, n3091);
  and g4926 (n3092, n_2987, n_2988);
  not g4927 (n_2989, n3092);
  and g4928 (n3093, n3089, n_2989);
  not g4929 (n_2990, n1213);
  and g4930 (n3094, n_2990, n1784);
  and g4931 (n3095, \in1[126] , n1787);
  and g4932 (n3096, \in0[126] , n_1849);
  not g4933 (n_2991, n3095);
  not g4934 (n_2992, n3096);
  and g4935 (n3097, n_2991, n_2992);
  and g4936 (n3098, \in3[126] , n1792);
  and g4937 (n3099, \in2[126] , n_1854);
  not g4938 (n_2993, n3098);
  not g4939 (n_2994, n3099);
  and g4940 (n3100, n_2993, n_2994);
  not g4941 (n_2995, n3100);
  and g4942 (n3101, n3097, n_2995);
  and g4943 (n3102, \in1[125] , n1787);
  and g4944 (n3103, \in0[125] , n_1849);
  not g4945 (n_2996, n3102);
  not g4946 (n_2997, n3103);
  and g4947 (n3104, n_2996, n_2997);
  and g4948 (n3105, \in3[125] , n1792);
  and g4949 (n3106, \in2[125] , n_1854);
  not g4950 (n_2998, n3105);
  not g4951 (n_2999, n3106);
  and g4952 (n3107, n_2998, n_2999);
  not g4953 (n_3000, n3107);
  and g4954 (n3108, n3104, n_3000);
  not g4955 (n_3001, n3101);
  not g4956 (n_3002, n3108);
  and g4957 (n3109, n_3001, n_3002);
  not g4958 (n_3003, n3094);
  not g4964 (n_3006, n3089);
  and g4965 (n3113, n_3006, n3092);
  not g4966 (n_3007, n3104);
  and g4967 (n3114, n_3007, n3107);
  not g4968 (n_3008, n3113);
  not g4969 (n_3009, n3114);
  and g4970 (n3115, n_3008, n_3009);
  not g4971 (n_3010, n3115);
  and g4972 (n3116, n3109, n_3010);
  not g4973 (n_3011, n3097);
  and g4974 (n3117, n_3011, n3100);
  not g4975 (n_3012, n3116);
  not g4976 (n_3013, n3117);
  and g4977 (n3118, n_3012, n_3013);
  not g4978 (n_3014, n3118);
  and g4979 (n3119, n_3003, n_3014);
  not g4980 (n_3015, n3112);
  not g4981 (n_3016, n3119);
  and g4982 (n3120, n_3015, n_3016);
  not g4983 (n_3017, n1785);
  and g4984 (\address[1] , n_3017, n3120);
  not g4985 (n_3018, n2503);
  and g4986 (n3122, n_3018, \address[1] );
  not g4987 (n_3020, \address[1] );
  and g4988 (n3123, n_2407, n_3020);
  or g4989 (\result[0] , n3122, n3123);
  and g4990 (n3125, n_2416, \address[1] );
  not g4991 (n_3021, n2508);
  and g4992 (n3126, n_3021, n_3020);
  or g4993 (\result[1] , n3125, n3126);
  and g4994 (n3128, n_2415, \address[1] );
  and g4995 (n3129, n_2421, n_3020);
  or g4996 (\result[2] , n3128, n3129);
  and g4997 (n3131, n_2400, \address[1] );
  and g4998 (n3132, n_2426, n_3020);
  or g4999 (\result[3] , n3131, n3132);
  not g5000 (n_3022, n2484);
  and g5001 (n3134, n_3022, \address[1] );
  and g5002 (n3135, n_2430, n_3020);
  or g5003 (\result[4] , n3134, n3135);
  not g5004 (n_3023, n2478);
  and g5005 (n3137, n_3023, \address[1] );
  and g5006 (n3138, n_2435, n_3020);
  or g5007 (\result[5] , n3137, n3138);
  not g5008 (n_3024, n2472);
  and g5009 (n3140, n_3024, \address[1] );
  and g5010 (n3141, n_2440, n_3020);
  or g5011 (\result[6] , n3140, n3141);
  and g5012 (n3143, n_2383, \address[1] );
  and g5013 (n3144, n_2446, n_3020);
  or g5014 (\result[7] , n3143, n3144);
  not g5015 (n_3025, n2462);
  and g5016 (n3146, n_3025, \address[1] );
  and g5017 (n3147, n_2453, n_3020);
  or g5018 (\result[8] , n3146, n3147);
  not g5019 (n_3026, n2459);
  and g5020 (n3149, n_3026, \address[1] );
  and g5021 (n3150, n_2460, n_3020);
  or g5022 (\result[9] , n3149, n3150);
  and g5023 (n3152, n_2374, \address[1] );
  and g5024 (n3153, n_2465, n_3020);
  or g5025 (\result[10] , n3152, n3153);
  and g5026 (n3155, n_2369, \address[1] );
  and g5027 (n3156, n_2470, n_3020);
  or g5028 (\result[11] , n3155, n3156);
  and g5029 (n3158, n_2364, \address[1] );
  and g5030 (n3159, n_2475, n_3020);
  or g5031 (\result[12] , n3158, n3159);
  and g5032 (n3161, n_2359, \address[1] );
  and g5033 (n3162, n_2480, n_3020);
  or g5034 (\result[13] , n3161, n3162);
  and g5035 (n3164, n_2354, \address[1] );
  and g5036 (n3165, n_2485, n_3020);
  or g5037 (\result[14] , n3164, n3165);
  and g5038 (n3167, n_2349, \address[1] );
  and g5039 (n3168, n_2490, n_3020);
  or g5040 (\result[15] , n3167, n3168);
  not g5041 (n_3027, n2414);
  and g5042 (n3170, n_3027, \address[1] );
  and g5043 (n3171, n_2497, n_3020);
  or g5044 (\result[16] , n3170, n3171);
  not g5045 (n_3028, n2411);
  and g5046 (n3173, n_3028, \address[1] );
  and g5047 (n3174, n_2504, n_3020);
  or g5048 (\result[17] , n3173, n3174);
  and g5049 (n3176, n_2340, \address[1] );
  and g5050 (n3177, n_2509, n_3020);
  or g5051 (\result[18] , n3176, n3177);
  and g5052 (n3179, n_2335, \address[1] );
  and g5053 (n3180, n_2514, n_3020);
  or g5054 (\result[19] , n3179, n3180);
  and g5055 (n3182, n_2330, \address[1] );
  and g5056 (n3183, n_2519, n_3020);
  or g5057 (\result[20] , n3182, n3183);
  and g5058 (n3185, n_2325, \address[1] );
  and g5059 (n3186, n_2524, n_3020);
  or g5060 (\result[21] , n3185, n3186);
  and g5061 (n3188, n_2320, \address[1] );
  and g5062 (n3189, n_2529, n_3020);
  or g5063 (\result[22] , n3188, n3189);
  and g5064 (n3191, n_2315, \address[1] );
  and g5065 (n3192, n_2534, n_3020);
  or g5066 (\result[23] , n3191, n3192);
  not g5067 (n_3029, n2366);
  and g5068 (n3194, n_3029, \address[1] );
  and g5069 (n3195, n_2541, n_3020);
  or g5070 (\result[24] , n3194, n3195);
  not g5071 (n_3030, n2363);
  and g5072 (n3197, n_3030, \address[1] );
  and g5073 (n3198, n_2548, n_3020);
  or g5074 (\result[25] , n3197, n3198);
  and g5075 (n3200, n_2306, \address[1] );
  and g5076 (n3201, n_2553, n_3020);
  or g5077 (\result[26] , n3200, n3201);
  and g5078 (n3203, n_2301, \address[1] );
  and g5079 (n3204, n_2558, n_3020);
  or g5080 (\result[27] , n3203, n3204);
  and g5081 (n3206, n_2296, \address[1] );
  and g5082 (n3207, n_2563, n_3020);
  or g5083 (\result[28] , n3206, n3207);
  and g5084 (n3209, n_2291, \address[1] );
  and g5085 (n3210, n_2568, n_3020);
  or g5086 (\result[29] , n3209, n3210);
  and g5087 (n3212, n_2286, \address[1] );
  and g5088 (n3213, n_2573, n_3020);
  or g5089 (\result[30] , n3212, n3213);
  and g5090 (n3215, n_2281, \address[1] );
  and g5091 (n3216, n_2578, n_3020);
  or g5092 (\result[31] , n3215, n3216);
  and g5093 (n3218, n_2276, \address[1] );
  and g5094 (n3219, n_2634, n_3020);
  or g5095 (\result[32] , n3218, n3219);
  and g5096 (n3221, n_2609, \address[1] );
  and g5097 (n3222, n_2635, n_3020);
  or g5098 (\result[33] , n3221, n3222);
  and g5099 (n3224, n_2619, \address[1] );
  and g5100 (n3225, n_2633, n_3020);
  or g5101 (\result[34] , n3224, n3225);
  and g5102 (n3227, n_2614, \address[1] );
  and g5103 (n3228, n_2632, n_3020);
  or g5104 (\result[35] , n3227, n3228);
  and g5105 (n3230, n_2597, \address[1] );
  and g5106 (n3231, n_2626, n_3020);
  or g5107 (\result[36] , n3230, n3231);
  and g5108 (n3233, n_2602, \address[1] );
  and g5109 (n3234, n_2627, n_3020);
  or g5110 (\result[37] , n3233, n3234);
  and g5111 (n3236, n_2590, \address[1] );
  and g5112 (n3237, n_2631, n_3020);
  or g5113 (\result[38] , n3236, n3237);
  and g5114 (n3239, n_2585, \address[1] );
  and g5115 (n3240, n_2625, n_3020);
  or g5116 (\result[39] , n3239, n3240);
  and g5117 (n3242, n_2648, \address[1] );
  and g5118 (n3243, n_2255, n_3020);
  or g5119 (\result[40] , n3242, n3243);
  and g5120 (n3245, n_2250, \address[1] );
  and g5121 (n3246, n_2257, n_3020);
  or g5122 (\result[41] , n3245, n3246);
  and g5123 (n3248, n_2243, \address[1] );
  and g5124 (n3249, n_2260, n_3020);
  or g5125 (\result[42] , n3248, n3249);
  and g5126 (n3251, n_2238, \address[1] );
  and g5127 (n3252, n_2237, n_3020);
  or g5128 (\result[43] , n3251, n3252);
  and g5129 (n3254, n_2225, \address[1] );
  and g5130 (n3255, n_2266, n_3020);
  or g5131 (\result[44] , n3254, n3255);
  and g5132 (n3257, n_2230, \address[1] );
  and g5133 (n3258, n_2267, n_3020);
  or g5134 (\result[45] , n3257, n3258);
  and g5135 (n3260, n_2218, \address[1] );
  and g5136 (n3261, n_2271, n_3020);
  or g5137 (\result[46] , n3260, n3261);
  and g5138 (n3263, n_2213, \address[1] );
  and g5139 (n3264, n_2212, n_3020);
  or g5140 (\result[47] , n3263, n3264);
  and g5141 (n3266, n_2660, \address[1] );
  and g5142 (n3267, n_2708, n_3020);
  or g5143 (\result[48] , n3266, n3267);
  and g5144 (n3269, n_2689, \address[1] );
  and g5145 (n3270, n_2709, n_3020);
  or g5146 (\result[49] , n3269, n3270);
  and g5147 (n3272, n_2699, \address[1] );
  and g5148 (n3273, n_2707, n_3020);
  or g5149 (\result[50] , n3272, n3273);
  and g5150 (n3275, n_2694, \address[1] );
  and g5151 (n3276, n_2706, n_3020);
  or g5152 (\result[51] , n3275, n3276);
  and g5153 (n3278, n_2682, \address[1] );
  and g5154 (n3279, n_2717, n_3020);
  or g5155 (\result[52] , n3278, n3279);
  and g5156 (n3281, n_2677, \address[1] );
  and g5157 (n3282, n_2718, n_3020);
  or g5158 (\result[53] , n3281, n3282);
  and g5159 (n3284, n_2670, \address[1] );
  and g5160 (n3285, n_2721, n_3020);
  or g5161 (\result[54] , n3284, n3285);
  and g5162 (n3287, n_2665, \address[1] );
  and g5163 (n3288, n_2705, n_3020);
  or g5164 (\result[55] , n3287, n3288);
  and g5165 (n3290, n_2728, \address[1] );
  and g5166 (n3291, n_2191, n_3020);
  or g5167 (\result[56] , n3290, n3291);
  and g5168 (n3293, n_2186, \address[1] );
  and g5169 (n3294, n_2193, n_3020);
  or g5170 (\result[57] , n3293, n3294);
  and g5171 (n3296, n_2179, \address[1] );
  and g5172 (n3297, n_2196, n_3020);
  or g5173 (\result[58] , n3296, n3297);
  and g5174 (n3299, n_2174, \address[1] );
  and g5175 (n3300, n_2173, n_3020);
  or g5176 (\result[59] , n3299, n3300);
  and g5177 (n3302, n_2161, \address[1] );
  and g5178 (n3303, n_2202, n_3020);
  or g5179 (\result[60] , n3302, n3303);
  and g5180 (n3305, n_2166, \address[1] );
  and g5181 (n3306, n_2203, n_3020);
  or g5182 (\result[61] , n3305, n3306);
  and g5183 (n3308, n_2154, \address[1] );
  and g5184 (n3309, n_2207, n_3020);
  or g5185 (\result[62] , n3308, n3309);
  and g5186 (n3311, n_2149, \address[1] );
  and g5187 (n3312, n_2148, n_3020);
  or g5188 (\result[63] , n3311, n3312);
  and g5189 (n3314, n_2138, \address[1] );
  and g5190 (n3315, n_2740, n_3020);
  or g5191 (\result[64] , n3314, n3315);
  and g5192 (n3317, n_2143, \address[1] );
  and g5193 (n3318, n_2741, n_3020);
  or g5194 (\result[65] , n3317, n3318);
  and g5195 (n3320, n_2131, \address[1] );
  and g5196 (n3321, n_2744, n_3020);
  or g5197 (\result[66] , n3320, n3321);
  and g5198 (n3323, n_2126, \address[1] );
  and g5199 (n3324, n_2739, n_3020);
  or g5200 (\result[67] , n3323, n3324);
  and g5201 (n3326, n_2750, \address[1] );
  and g5202 (n3327, n_2115, n_3020);
  or g5203 (\result[68] , n3326, n3327);
  and g5204 (n3329, n_2110, \address[1] );
  and g5205 (n3330, n_2117, n_3020);
  or g5206 (\result[69] , n3329, n3330);
  and g5207 (n3332, n_2103, \address[1] );
  and g5208 (n3333, n_2121, n_3020);
  or g5209 (\result[70] , n3332, n3333);
  and g5210 (n3335, n_2098, \address[1] );
  and g5211 (n3336, n_2097, n_3020);
  or g5212 (\result[71] , n3335, n3336);
  and g5213 (n3338, n_2778, \address[1] );
  and g5214 (n3339, n_2783, n_3020);
  or g5215 (\result[72] , n3338, n3339);
  and g5216 (n3341, n_2773, \address[1] );
  and g5217 (n3342, n_2784, n_3020);
  or g5218 (\result[73] , n3341, n3342);
  and g5219 (n3344, n_2766, \address[1] );
  and g5220 (n3345, n_2787, n_3020);
  or g5221 (\result[74] , n3344, n3345);
  and g5222 (n3347, n_2761, \address[1] );
  and g5223 (n3348, n_2782, n_3020);
  or g5224 (\result[75] , n3347, n3348);
  and g5225 (n3350, n_2793, \address[1] );
  and g5226 (n3351, n_2086, n_3020);
  or g5227 (\result[76] , n3350, n3351);
  and g5228 (n3353, n_2081, \address[1] );
  and g5229 (n3354, n_2088, n_3020);
  or g5230 (\result[77] , n3353, n3354);
  and g5231 (n3356, n_2074, \address[1] );
  and g5232 (n3357, n_2092, n_3020);
  or g5233 (\result[78] , n3356, n3357);
  and g5234 (n3359, n_2069, \address[1] );
  and g5235 (n3360, n_2068, n_3020);
  or g5236 (\result[79] , n3359, n3360);
  and g5237 (n3362, n_2046, \address[1] );
  and g5238 (n3363, n_2804, n_3020);
  or g5239 (\result[80] , n3362, n3363);
  and g5240 (n3365, n_2063, \address[1] );
  and g5241 (n3366, n_2805, n_3020);
  or g5242 (\result[81] , n3365, n3366);
  and g5243 (n3368, n_2056, \address[1] );
  and g5244 (n3369, n_2808, n_3020);
  or g5245 (\result[82] , n3368, n3369);
  and g5246 (n3371, n_2051, \address[1] );
  and g5247 (n3372, n_2803, n_3020);
  or g5248 (\result[83] , n3371, n3372);
  and g5249 (n3374, n_2814, \address[1] );
  and g5250 (n3375, n_2035, n_3020);
  or g5251 (\result[84] , n3374, n3375);
  and g5252 (n3377, n_2030, \address[1] );
  and g5253 (n3378, n_2037, n_3020);
  or g5254 (\result[85] , n3377, n3378);
  and g5255 (n3380, n_2023, \address[1] );
  and g5256 (n3381, n_2041, n_3020);
  or g5257 (\result[86] , n3380, n3381);
  and g5258 (n3383, n_2018, \address[1] );
  and g5259 (n3384, n_2017, n_3020);
  or g5260 (\result[87] , n3383, n3384);
  and g5261 (n3386, n_2842, \address[1] );
  and g5262 (n3387, n_2847, n_3020);
  or g5263 (\result[88] , n3386, n3387);
  and g5264 (n3389, n_2837, \address[1] );
  and g5265 (n3390, n_2848, n_3020);
  or g5266 (\result[89] , n3389, n3390);
  and g5267 (n3392, n_2830, \address[1] );
  and g5268 (n3393, n_2851, n_3020);
  or g5269 (\result[90] , n3392, n3393);
  and g5270 (n3395, n_2825, \address[1] );
  and g5271 (n3396, n_2846, n_3020);
  or g5272 (\result[91] , n3395, n3396);
  and g5273 (n3398, n_2857, \address[1] );
  and g5274 (n3399, n_2006, n_3020);
  or g5275 (\result[92] , n3398, n3399);
  and g5276 (n3401, n_2001, \address[1] );
  and g5277 (n3402, n_2008, n_3020);
  or g5278 (\result[93] , n3401, n3402);
  and g5279 (n3404, n_1994, \address[1] );
  and g5280 (n3405, n_2012, n_3020);
  or g5281 (\result[94] , n3404, n3405);
  and g5282 (n3407, n_1989, \address[1] );
  and g5283 (n3408, n_1988, n_3020);
  or g5284 (\result[95] , n3407, n3408);
  and g5285 (n3410, n_1966, \address[1] );
  and g5286 (n3411, n_2868, n_3020);
  or g5287 (\result[96] , n3410, n3411);
  and g5288 (n3413, n_1983, \address[1] );
  and g5289 (n3414, n_2869, n_3020);
  or g5290 (\result[97] , n3413, n3414);
  and g5291 (n3416, n_1976, \address[1] );
  and g5292 (n3417, n_2872, n_3020);
  or g5293 (\result[98] , n3416, n3417);
  and g5294 (n3419, n_1971, \address[1] );
  and g5295 (n3420, n_2867, n_3020);
  or g5296 (\result[99] , n3419, n3420);
  and g5297 (n3422, n_2878, \address[1] );
  and g5298 (n3423, n_1955, n_3020);
  or g5299 (\result[100] , n3422, n3423);
  and g5300 (n3425, n_1950, \address[1] );
  and g5301 (n3426, n_1957, n_3020);
  or g5302 (\result[101] , n3425, n3426);
  and g5303 (n3428, n_1943, \address[1] );
  and g5304 (n3429, n_1961, n_3020);
  or g5305 (\result[102] , n3428, n3429);
  and g5306 (n3431, n_1938, \address[1] );
  and g5307 (n3432, n_1937, n_3020);
  or g5308 (\result[103] , n3431, n3432);
  and g5309 (n3434, n_2906, \address[1] );
  and g5310 (n3435, n_2911, n_3020);
  or g5311 (\result[104] , n3434, n3435);
  and g5312 (n3437, n_2901, \address[1] );
  and g5313 (n3438, n_2912, n_3020);
  or g5314 (\result[105] , n3437, n3438);
  and g5315 (n3440, n_2894, \address[1] );
  and g5316 (n3441, n_2915, n_3020);
  or g5317 (\result[106] , n3440, n3441);
  and g5318 (n3443, n_2889, \address[1] );
  and g5319 (n3444, n_2910, n_3020);
  or g5320 (\result[107] , n3443, n3444);
  and g5321 (n3446, n_2921, \address[1] );
  and g5322 (n3447, n_1926, n_3020);
  or g5323 (\result[108] , n3446, n3447);
  and g5324 (n3449, n_1921, \address[1] );
  and g5325 (n3450, n_1928, n_3020);
  or g5326 (\result[109] , n3449, n3450);
  and g5327 (n3452, n_1914, \address[1] );
  and g5328 (n3453, n_1932, n_3020);
  or g5329 (\result[110] , n3452, n3453);
  and g5330 (n3455, n_1909, \address[1] );
  and g5331 (n3456, n_1908, n_3020);
  or g5332 (\result[111] , n3455, n3456);
  and g5333 (n3458, n_1886, \address[1] );
  and g5334 (n3459, n_2932, n_3020);
  or g5335 (\result[112] , n3458, n3459);
  and g5336 (n3461, n_1903, \address[1] );
  and g5337 (n3462, n_2933, n_3020);
  or g5338 (\result[113] , n3461, n3462);
  and g5339 (n3464, n_1896, \address[1] );
  and g5340 (n3465, n_2936, n_3020);
  or g5341 (\result[114] , n3464, n3465);
  and g5342 (n3467, n_1891, \address[1] );
  and g5343 (n3468, n_2931, n_3020);
  or g5344 (\result[115] , n3467, n3468);
  and g5345 (n3470, n_2942, \address[1] );
  and g5346 (n3471, n_1876, n_3020);
  or g5347 (\result[116] , n3470, n3471);
  and g5348 (n3473, n_1872, \address[1] );
  and g5349 (n3474, n_1877, n_3020);
  or g5350 (\result[117] , n3473, n3474);
  and g5351 (n3476, n_1863, \address[1] );
  and g5352 (n3477, n_1881, n_3020);
  or g5353 (\result[118] , n3476, n3477);
  and g5354 (n3479, n_1858, \address[1] );
  and g5355 (n3480, n_1857, n_3020);
  or g5356 (\result[119] , n3479, n3480);
  and g5357 (n3482, n_2970, \address[1] );
  and g5358 (n3483, n_2975, n_3020);
  or g5359 (\result[120] , n3482, n3483);
  and g5360 (n3485, n_2965, \address[1] );
  and g5361 (n3486, n_2976, n_3020);
  or g5362 (\result[121] , n3485, n3486);
  and g5363 (n3488, n_2958, \address[1] );
  and g5364 (n3489, n_2979, n_3020);
  or g5365 (\result[122] , n3488, n3489);
  and g5366 (n3491, n_2953, \address[1] );
  and g5367 (n3492, n_2974, n_3020);
  or g5368 (\result[123] , n3491, n3492);
  and g5369 (n3494, n_2989, \address[1] );
  and g5370 (n3495, n_3006, n_3020);
  or g5371 (\result[124] , n3494, n3495);
  and g5372 (n3497, n_3000, \address[1] );
  and g5373 (n3498, n_3007, n_3020);
  or g5374 (\result[125] , n3497, n3498);
  and g5375 (n3500, n_2995, \address[1] );
  and g5376 (n3501, n_3011, n_3020);
  or g5377 (\result[126] , n3500, n3501);
  and g5378 (n3503, n_2990, n3120);
  not g5379 (n_3031, n3503);
  and g5380 (\result[127] , n1784, n_3031);
  and g5381 (n3505, n1792, \address[1] );
  and g5382 (n3506, n1787, n_3020);
  or g5383 (\address[0] , n3505, n3506);
  and g5384 (n3112, n_3161, n_3162, n_3003, n3109);
  not g5385 (n_3161, n3086);
  not g5386 (n_3162, n3093);
  and g5387 (n1203, n_3163, n_3164, n_908, n1200);
  not g5388 (n_3163, n1195);
  not g5389 (n_3164, n1196);
  and g5390 (n3076, n_3165, n_3166, n3059, n_2971);
  not g5391 (n_3165, n3044);
  not g5392 (n_3166, n3073);
  and g5393 (n1774, n_3167, n_3168, n_1831, n1771);
  not g5394 (n_3167, n1766);
  not g5395 (n_3168, n1767);
  nor g5396 (n3044, n1796, n1823, n1825, n3041);
  and g5397 (n1185, n_3169, n_3170, n1180, n_880);
  not g5398 (n_3169, n1177);
  not g5399 (n_3170, n1182);
  and g5400 (n3041, n_3171, n_3172, n1805, n_1875);
  not g5401 (n_3171, n3037);
  not g5402 (n_3172, n3038);
  nor g5403 (n1177, n643, n652, n654, n1174);
  and g5404 (n1756, n_3173, n_3174, n1751, n_1803);
  not g5405 (n_3173, n1748);
  not g5406 (n_3174, n1753);
  and g5407 (n1174, n_3175, n_3176, n646, n_16);
  not g5408 (n_3175, n1170);
  not g5409 (n_3176, n1171);
  nor g5410 (n1748, n1214, n1223, n1225, n1745);
  and g5411 (n3027, n_3177, n_3178, n1847, n_2928);
  not g5412 (n_3177, n1832);
  not g5413 (n_3178, n3024);
  and g5414 (n1745, n_3179, n_3180, n1217, n_938);
  not g5415 (n_3179, n1741);
  not g5416 (n_3180, n1742);
  nor g5417 (n3024, n1861, n1888, n1890, n3021);
  and g5418 (n1160, n_3181, n_3182, n658, n_845);
  not g5419 (n_3181, n655);
  not g5420 (n_3182, n1157);
  and g5421 (n3021, n_3183, n_3184, n1870, n_1927);
  not g5422 (n_3183, n3017);
  not g5423 (n_3184, n3018);
  nor g5424 (n1157, n660, n669, n671, n1154);
  and g5425 (n1731, n_3185, n_3186, n1229, n_1768);
  not g5426 (n_3185, n1226);
  not g5427 (n_3186, n1728);
  and g5428 (n1154, n_3187, n_3188, n663, n_51);
  not g5429 (n_3187, n1150);
  not g5430 (n_3188, n1151);
  nor g5431 (n1728, n1231, n1240, n1242, n1725);
  and g5432 (n3007, n_3189, n_3190, n2990, n_2907);
  not g5433 (n_3189, n2975);
  not g5434 (n_3190, n3004);
  and g5435 (n1725, n_3191, n_3192, n1234, n_973);
  not g5436 (n_3191, n1721);
  not g5437 (n_3192, n1722);
  nor g5438 (n2975, n1897, n1924, n1926, n2972);
  and g5439 (n1140, n_3193, n_3194, n1135, n_824);
  not g5440 (n_3193, n1132);
  not g5441 (n_3194, n1137);
  and g5442 (n2972, n_3195, n_3196, n1906, n_1956);
  not g5443 (n_3195, n2968);
  not g5444 (n_3196, n2969);
  nor g5445 (n1132, n672, n681, n683, n1129);
  and g5446 (n1711, n_3197, n_3198, n1706, n_1747);
  not g5447 (n_3197, n1703);
  not g5448 (n_3198, n1708);
  and g5449 (n1129, n_3199, n_3200, n675, n_72);
  not g5450 (n_3199, n1125);
  not g5451 (n_3200, n1126);
  nor g5452 (n1703, n1243, n1252, n1254, n1700);
  and g5453 (n2958, n_3201, n_3202, n1948, n_2864);
  not g5454 (n_3201, n1933);
  not g5455 (n_3202, n2955);
  and g5456 (n1700, n_3203, n_3204, n1246, n_994);
  not g5457 (n_3203, n1696);
  not g5458 (n_3204, n1697);
  nor g5459 (n2955, n1962, n1989, n1991, n2952);
  and g5460 (n1115, n_3205, n_3206, n687, n_789);
  not g5461 (n_3205, n684);
  not g5462 (n_3206, n1112);
  and g5463 (n2952, n_3207, n_3208, n1971, n_2007);
  not g5464 (n_3207, n2948);
  not g5465 (n_3208, n2949);
  nor g5466 (n1112, n689, n698, n700, n1109);
  and g5467 (n1686, n_3209, n_3210, n1258, n_1712);
  not g5468 (n_3209, n1255);
  not g5469 (n_3210, n1683);
  and g5470 (n1109, n_3211, n_3212, n692, n_107);
  not g5471 (n_3211, n1105);
  not g5472 (n_3212, n1106);
  nor g5473 (n1683, n1260, n1269, n1271, n1680);
  and g5474 (n2938, n_3213, n_3214, n2921, n_2843);
  not g5475 (n_3213, n2906);
  not g5476 (n_3214, n2935);
  and g5477 (n1680, n_3215, n_3216, n1263, n_1029);
  not g5478 (n_3215, n1676);
  not g5479 (n_3216, n1677);
  nor g5480 (n2906, n1998, n2025, n2027, n2903);
  and g5481 (n1095, n_3217, n_3218, n1090, n_768);
  not g5482 (n_3217, n1087);
  not g5483 (n_3218, n1092);
  and g5484 (n2903, n_3219, n_3220, n2007, n_2036);
  not g5485 (n_3219, n2899);
  not g5486 (n_3220, n2900);
  nor g5487 (n1087, n701, n710, n712, n1084);
  and g5488 (n1666, n_3221, n_3222, n1661, n_1691);
  not g5489 (n_3221, n1658);
  not g5490 (n_3222, n1663);
  and g5491 (n1084, n_3223, n_3224, n704, n_128);
  not g5492 (n_3223, n1080);
  not g5493 (n_3224, n1081);
  nor g5494 (n1658, n1272, n1281, n1283, n1655);
  and g5495 (n2889, n_3225, n_3226, n2049, n_2800);
  not g5496 (n_3225, n2034);
  not g5497 (n_3226, n2886);
  and g5498 (n1655, n_3227, n_3228, n1275, n_1050);
  not g5499 (n_3227, n1651);
  not g5500 (n_3228, n1652);
  nor g5501 (n2886, n2063, n2090, n2092, n2883);
  and g5502 (n1070, n_3229, n_3230, n716, n_733);
  not g5503 (n_3229, n713);
  not g5504 (n_3230, n1067);
  and g5505 (n2883, n_3231, n_3232, n2072, n_2087);
  not g5506 (n_3231, n2879);
  not g5507 (n_3232, n2880);
  nor g5508 (n1067, n718, n727, n729, n1064);
  and g5509 (n1641, n_3233, n_3234, n1287, n_1656);
  not g5510 (n_3233, n1284);
  not g5511 (n_3234, n1638);
  and g5512 (n1064, n_3235, n_3236, n721, n_163);
  not g5513 (n_3235, n1060);
  not g5514 (n_3236, n1061);
  nor g5515 (n1638, n1289, n1298, n1300, n1635);
  and g5516 (n2869, n_3237, n_3238, n2852, n_2779);
  not g5517 (n_3237, n2837);
  not g5518 (n_3238, n2866);
  and g5519 (n1635, n_3239, n_3240, n1292, n_1085);
  not g5520 (n_3239, n1631);
  not g5521 (n_3240, n1632);
  nor g5522 (n2837, n2099, n2126, n2128, n2834);
  and g5523 (n1050, n_3241, n_3242, n1045, n_712);
  not g5524 (n_3241, n1042);
  not g5525 (n_3242, n1047);
  and g5526 (n2834, n_3243, n_3244, n2108, n_2116);
  not g5527 (n_3243, n2830);
  not g5528 (n_3244, n2831);
  nor g5529 (n1042, n730, n739, n741, n1039);
  and g5530 (n1621, n_3245, n_3246, n1616, n_1635);
  not g5531 (n_3245, n1613);
  not g5532 (n_3246, n1618);
  and g5533 (n1039, n_3247, n_3248, n733, n_184);
  not g5534 (n_3247, n1035);
  not g5535 (n_3248, n1036);
  nor g5536 (n1613, n1301, n1310, n1312, n1610);
  and g5537 (n2820, n_3249, n_3250, n2143, n_2736);
  not g5538 (n_3249, n2150);
  not g5539 (n_3250, n2817);
  and g5540 (n1610, n_3251, n_3252, n1304, n_1106);
  not g5541 (n_3251, n1606);
  not g5542 (n_3252, n1607);
  nor g5543 (n_3256, n2164, n2227);
  and g5544 (n2817, n_3253, n_3254, n_3255, n_3256);
  not g5545 (n_3253, n2232);
  not g5546 (n_3254, n2234);
  not g5547 (n_3255, n2813);
  and g5548 (n1025, n_3257, n_3258, n744, n_679);
  not g5549 (n_3257, n1021);
  not g5550 (n_3258, n1022);
  nor g5551 (n_3259, n2808, n2809);
  and g5552 (n2813, n2205, n2189, n_2192, n_3259);
  nor g5553 (n_3263, n746, n767);
  and g5554 (n1021, n_3260, n_3261, n_3262, n_3263);
  not g5555 (n_3260, n772);
  not g5556 (n_3261, n774);
  not g5557 (n_3262, n1017);
  and g5558 (n1596, n_3264, n_3265, n1315, n_1602);
  not g5559 (n_3264, n1592);
  not g5560 (n_3265, n1593);
  nor g5561 (n2808, n2787, n2788, n2798, n2805);
  nor g5562 (n_3266, n1012, n1013);
  and g5563 (n1017, n757, n753, n_233, n_3266);
  nor g5564 (n_3270, n1317, n1338);
  and g5565 (n1592, n_3267, n_3268, n_3269, n_3270);
  not g5566 (n_3267, n1343);
  not g5567 (n_3268, n1345);
  not g5568 (n_3269, n1588);
  and g5569 (n2787, n_3271, n_3272, n2761, n2784);
  not g5570 (n_3271, n2723);
  not g5571 (n_3272, n2730);
  nor g5572 (n1012, n991, n992, n1002, n1009);
  nor g5573 (n_3273, n1583, n1584);
  and g5574 (n1588, n1328, n1324, n_1155, n_3273);
  nor g5575 (n_3277, n2241, n2304);
  and g5576 (n2723, n_3274, n_3275, n_3276, n_3277);
  not g5577 (n_3274, n2309);
  not g5578 (n_3275, n2311);
  not g5579 (n_3276, n2719);
  nor g5580 (n_3278, n975, n976);
  and g5581 (n991, n983, n_640, n987, n_3278);
  nor g5582 (n1583, n1562, n1563, n1573, n1580);
  nor g5583 (n_3279, n2714, n2715);
  and g5584 (n2719, n2266, n2282, n_2256, n_3279);
  nor g5585 (n_3283, n775, n796);
  and g5586 (n975, n_3280, n_3281, n_3282, n_3283);
  not g5587 (n_3280, n801);
  not g5588 (n_3281, n803);
  not g5589 (n_3282, n971);
  nor g5590 (n_3284, n1546, n1547);
  and g5591 (n1562, n1554, n_1563, n1558, n_3284);
  nor g5592 (n_3288, n2692, n2693);
  and g5593 (n2714, n_3285, n_3286, n_3287, n_3288);
  not g5594 (n_3285, n2698);
  not g5595 (n_3286, n2700);
  not g5596 (n_3287, n2710);
  nor g5597 (n_3289, n966, n967);
  and g5598 (n971, n782, n786, n_281, n_3289);
  nor g5599 (n_3293, n1346, n1367);
  and g5600 (n1546, n_3290, n_3291, n_3292, n_3293);
  not g5601 (n_3290, n1372);
  not g5602 (n_3291, n1374);
  not g5603 (n_3292, n1542);
  and g5604 (n2692, n_3294, n_3295, n2666, n2689);
  not g5605 (n_3294, n2318);
  not g5606 (n_3295, n2635);
  nor g5607 (n_3299, n944, n945);
  and g5608 (n966, n_3296, n_3297, n_3298, n_3299);
  not g5609 (n_3296, n950);
  not g5610 (n_3297, n952);
  not g5611 (n_3298, n962);
  nor g5612 (n_3300, n1537, n1538);
  and g5613 (n1542, n1353, n1357, n_1203, n_3300);
  nor g5614 (n_3301, n804, n929);
  and g5615 (n944, n936, n_576, n940, n_3301);
  nor g5616 (n_3305, n1515, n1516);
  and g5617 (n1537, n_3302, n_3303, n_3304, n_3305);
  not g5618 (n_3302, n1521);
  not g5619 (n_3303, n1523);
  not g5620 (n_3304, n1533);
  nor g5621 (n_3306, n1375, n1500);
  and g5622 (n1515, n1507, n_1499, n1511, n_3306);
endmodule

