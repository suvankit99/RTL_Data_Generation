
module c5315(N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31,
     N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70,
     N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97,
     N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118,
     N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131,
     N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155,
     N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188,
     N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225,
     N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264,
     N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302,
     N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341,
     N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389,
     N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514,
     N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574,
     N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599,
     N603, N607, N610, N613, N616, N619, N625, N631, N709, N816, N1066,
     N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145,
     N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061,
     N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357,
     N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279,
     N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646,
     N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363,
     N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471,
     N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515,
     N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601,
     N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699,
     N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735,
     N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755,
     N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123,
     N8124, N8127, N8128);
  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34,
       N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73,
       N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97,
       N100, N103, N106, N109, N112, N113, N114, N115, N116, N117,
       N118, N119, N120, N121, N122, N123, N126, N127, N128, N129,
       N130, N131, N132, N135, N136, N137, N140, N141, N145, N146,
       N149, N152, N155, N158, N161, N164, N167, N170, N173, N176,
       N179, N182, N185, N188, N191, N194, N197, N200, N203, N206,
       N209, N210, N217, N218, N225, N226, N233, N234, N241, N242,
       N245, N248, N251, N254, N257, N264, N265, N272, N273, N280,
       N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
       N316, N323, N324, N331, N332, N335, N338, N341, N348, N351,
       N358, N361, N366, N369, N372, N373, N374, N386, N389, N400,
       N411, N422, N435, N446, N457, N468, N479, N490, N503, N514,
       N523, N534, N545, N549, N552, N556, N559, N562, N566, N571,
       N574, N577, N580, N583, N588, N591, N592, N595, N596, N597,
       N598, N599, N603, N607, N610, N613, N616, N619, N625, N631;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142,
       N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972,
       N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584,
       N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272,
       N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388,
       N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926,
       N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467,
       N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504,
       N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521,
       N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
       N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705,
       N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741,
       N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761,
       N8075, N8076, N8123, N8124, N8127, N8128;
  wire N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34,
       N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73,
       N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97,
       N100, N103, N106, N109, N112, N113, N114, N115, N116, N117,
       N118, N119, N120, N121, N122, N123, N126, N127, N128, N129,
       N130, N131, N132, N135, N136, N137, N140, N141, N145, N146,
       N149, N152, N155, N158, N161, N164, N167, N170, N173, N176,
       N179, N182, N185, N188, N191, N194, N197, N200, N203, N206,
       N209, N210, N217, N218, N225, N226, N233, N234, N241, N242,
       N245, N248, N251, N254, N257, N264, N265, N272, N273, N280,
       N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
       N316, N323, N324, N331, N332, N335, N338, N341, N348, N351,
       N358, N361, N366, N369, N372, N373, N374, N386, N389, N400,
       N411, N422, N435, N446, N457, N468, N479, N490, N503, N514,
       N523, N534, N545, N549, N552, N556, N559, N562, N566, N571,
       N574, N577, N580, N583, N588, N591, N592, N595, N596, N597,
       N598, N599, N603, N607, N610, N613, N616, N619, N625, N631;
  wire N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142,
       N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972,
       N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584,
       N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272,
       N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388,
       N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926,
       N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467,
       N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504,
       N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521,
       N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
       N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705,
       N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741,
       N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761,
       N8075, N8076, N8123, N8124, N8127, N8128;
  wire N1042, N1043, N1067, N1080, N1092, N1104, N1146, N1148;
  wire N1149, N1150, N1151, N1157, N1219, N1475, N1588, N1660;
  wire N1755, N1758, N2349, N2350, N2585, N2586, N2587, N2588;
  wire N2589, N2591, N2592, N2593, N2594, N2595, N2596, N2597;
  wire N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605;
  wire N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613;
  wire N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621;
  wire N2622, N2624, N2625, N2626, N2628, N2629, N2630, N2631;
  wire N2632, N2633, N2634, N2635, N2636, N2637, N2653, N2664;
  wire N2703, N2709, N2710, N2711, N2712, N2713, N2714, N2715;
  wire N2728, N2739, N2778, N2779, N2790, N2801, N2812, N2823;
  wire N2825, N2827, N2829, N2831, N2832, N2833, N2834, N2835;
  wire N2836, N2837, N2838, N2839, N2841, N2843, N2845, N2847;
  wire N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855;
  wire N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874;
  wire N2875, N2876, N2901, N2902, N2903, N2905, N2907, N2908;
  wire N2909, N2910, N2911, N2912, N2915, N2917, N2919, N2920;
  wire N2921, N2922, N2923, N2924, N2925, N2934, N2935, N2936;
  wire N2937, N2938, N2939, N2940, N2941, N2942, N2954, N2955;
  wire N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963;
  wire N2969, N2970, N2971, N2979, N2980, N2981, N2982, N2983;
  wire N2984, N2985, N2986, N2999, N3013, N3023, N3024, N3025;
  wire N3026, N3027, N3028, N3029, N3030, N3032, N3063, N3068;
  wire N3071, N3072, N3142, N3401, N3402, N3403, N3404, N3405;
  wire N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413;
  wire N3414, N3415, N3416, N3444, N3445, N3446, N3447, N3448;
  wire N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456;
  wire N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466;
  wire N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3502;
  wire N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511;
  wire N3512, N3513, N3514, N3515, N3558, N3559, N3560, N3561;
  wire N3562, N3563, N3605, N3606, N3607, N3608, N3609, N3610;
  wire N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621;
  wire N3622, N3623, N3624, N3627, N3628, N3629, N3630, N3631;
  wire N3632, N3633, N3634, N3635, N3638, N3641, N3642, N3643;
  wire N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651;
  wire N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659;
  wire N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667;
  wire N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675;
  wire N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683;
  wire N3684, N3685, N3686, N3687, N3688, N3689, N3700, N3701;
  wire N3702, N3703, N3704, N3705, N3708, N3709, N3710, N3711;
  wire N3712, N3713, N3715, N3716, N3717, N3718, N3719, N3720;
  wire N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728;
  wire N3729, N3730, N3731, N3732, N3738, N3739, N3740, N3742;
  wire N3743, N3744, N3745, N3746, N3747, N3753, N3757, N3758;
  wire N3761, N3763, N3764, N3765, N3766, N3767, N3768, N3769;
  wire N3770, N3771, N3775, N3781, N3782, N3783, N3784, N3785;
  wire N3786, N3787, N3788, N3789, N3793, N3797, N3800, N3801;
  wire N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809;
  wire N3810, N3813, N3816, N3823, N3824, N3827, N3828, N3829;
  wire N3831, N3834, N3835, N3836, N3837, N3838, N3839, N3840;
  wire N3841, N3842, N3849, N3855, N3861, N3867, N3873, N3881;
  wire N3887, N3893, N3908, N3909, N3911, N3914, N3915, N3916;
  wire N3917, N3918, N3919, N3920, N3921, N3927, N3933, N3942;
  wire N3948, N3956, N3962, N3968, N3975, N3976, N3977, N3980;
  wire N3982, N3987, N3988, N3989, N3990, N3991, N3998, N4008;
  wire N4011, N4024, N4027, N4031, N4032, N4033, N4034, N4035;
  wire N4036, N4037, N4038, N4039, N4040, N4042, N4067, N4088;
  wire N4091, N4094, N4097, N4100, N4103, N4106, N4109, N4144;
  wire N4147, N4153, N4156, N4159, N4183, N4185, N4188, N4191;
  wire N4196, N4197, N4198, N4199, N4200, N4203, N4223, N4224;
  wire N4225, N4228, N4231, N4234, N4237, N4240, N4243, N4246;
  wire N4249, N4252, N4264, N4267, N4268, N4273, N4274, N4276;
  wire N4277, N4280, N4284, N4290, N4297, N4298, N4301, N4305;
  wire N4310, N4357, N4364, N4379, N4385, N4392, N4396, N4400;
  wire N4405, N4515, N4521, N4523, N4524, N4547, N4575, N4608;
  wire N4627, N4701, N4702, N4721, N4724, N4725, N4726, N4727;
  wire N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735;
  wire N4736, N4741, N4855, N4856, N4939, N4953, N4954, N4955;
  wire N4956, N4957, N4958, N4959, N4960, N4961, N4965, N4966;
  wire N4967, N4968, N4972, N4973, N4974, N4975, N4976, N4978;
  wire N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986;
  wire N4987, N5049, N5052, N5053, N5054, N5057, N5058, N5059;
  wire N5060, N5061, N5062, N5063, N5065, N5066, N5069, N5070;
  wire N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078;
  wire N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086;
  wire N5087, N5106, N5107, N5108, N5109, N5110, N5111, N5112;
  wire N5113, N5114, N5115, N5116, N5117, N5119, N5120, N5137;
  wire N5140, N5145, N5147, N5148, N5153, N5154, N5155, N5156;
  wire N5160, N5161, N5162, N5163, N5164, N5165, N5176, N5232;
  wire N5233, N5234, N5235, N5236, N5239, N5241, N5242, N5243;
  wire N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5261;
  wire N5262, N5263, N5264, N5274, N5275, N5303, N5304, N5305;
  wire N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5315;
  wire N5319, N5324, N5328, N5331, N5332, N5346, N5363, N5364;
  wire N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5377;
  wire N5382, N5385, N5389, N5396, N5407, N5418, N5424, N5431;
  wire N5441, N5452, N5462, N5469, N5562, N5573, N5579, N5595;
  wire N5606, N5616, N5622, N5692, N5696, N5700, N5703, N5707;
  wire N5711, N5728, N5736, N5739, N5742, N5745, N5755, N5756;
  wire N5954, N5955, N5956, N6023, N6024, N6025, N6028, N6044;
  wire N6066, N6067, N6068, N6069, N6071, N6072, N6073, N6074;
  wire N6079, N6080, N6083, N6084, N6085, N6088, N6089, N6091;
  wire N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101;
  wire N6102, N6103, N6104, N6105, N6106, N6107, N6117, N6127;
  wire N6133, N6138, N6139, N6140, N6143, N6144, N6146, N6147;
  wire N6149, N6152, N6153, N6154, N6155, N6156, N6157, N6158;
  wire N6159, N6160, N6161, N6162, N6163, N6164, N6175, N6184;
  wire N6189, N6194, N6197, N6200, N6203, N6206, N6221, N6234;
  wire N6235, N6373, N6374, N6375, N6376, N6377, N6378, N6382;
  wire N6386, N6397, N6411, N6419, N6427, N6434, N6437, N6445;
  wire N6469, N6471, N6473, N6474, N6475, N6476, N6477, N6478;
  wire N6482, N6486, N6490, N6494, N6500, N6504, N6508, N6512;
  wire N6536, N6539, N6553, N6556, N6566, N6569, N6572, N6575;
  wire N6580, N6584, N6587, N6606, N6609, N6619, N6622, N6630;
  wire N6631, N6632, N6633, N6634, N6637, N6650, N6651, N6653;
  wire N6657, N6660, N6661, N6662, N6664, N6666, N6668, N6670;
  wire N6672, N6675, N6689, N6690, N6691, N6693, N6695, N6698;
  wire N6699, N6700, N6703, N6708, N6710, N6712, N6713, N6714;
  wire N6715, N6718, N6719, N6720, N6721, N6722, N6792, N6795;
  wire N6801, N6802, N6806, N6807, N6808, N6809, N6810, N6811;
  wire N6812, N6814, N6815, N6816, N6817, N6823, N6824, N6825;
  wire N6826, N6827, N6828, N6829, N6830, N6831, N6834, N6835;
  wire N6836, N6837, N6838, N6839, N6841, N6842, N6843, N6844;
  wire N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857;
  wire N6860, N6861, N6862, N6863, N6866, N6872, N6873, N6874;
  wire N6875, N6876, N6879, N6880, N6881, N6889, N6890, N6891;
  wire N6894, N6895, N6896, N6897, N6900, N6901, N6909, N6912;
  wire N6913, N6914, N6915, N6916, N6919, N6922, N6923, N6932;
  wire N6935, N6936, N6937, N6938, N6939, N6940, N6946, N6947;
  wire N6948, N6949, N6953, N6954, N6955, N6956, N6957, N6958;
  wire N6964, N6965, N6966, N6967, N6973, N6974, N6975, N6976;
  wire N6977, N6978, N6979, N6987, N6990, N6999, N7002, N7003;
  wire N7006, N7011, N7012, N7013, N7016, N7018, N7019, N7020;
  wire N7021, N7022, N7023, N7028, N7031, N7034, N7037, N7040;
  wire N7041, N7044, N7045, N7046, N7047, N7048, N7049, N7054;
  wire N7057, N7060, N7064, N7065, N7072, N7073, N7075, N7076;
  wire N7079, N7080, N7084, N7085, N7087, N7088, N7089, N7090;
  wire N7094, N7097, N7101, N7114, N7115, N7116, N7125, N7126;
  wire N7127, N7130, N7131, N7139, N7140, N7141, N7146, N7147;
  wire N7149, N7150, N7151, N7152, N7153, N7158, N7159, N7160;
  wire N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180;
  wire N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188;
  wire N7189, N7190, N7196, N7197, N7198, N7204, N7205, N7206;
  wire N7207, N7208, N7209, N7212, N7215, N7216, N7217, N7218;
  wire N7219, N7222, N7225, N7228, N7229, N7236, N7239, N7242;
  wire N7245, N7250, N7257, N7260, N7263, N7268, N7269, N7270;
  wire N7276, N7282, N7288, N7294, N7300, N7301, N7304, N7310;
  wire N7320, N7321, N7328, N7338, N7339, N7340, N7341, N7342;
  wire N7349, N7357, N7364, N7402, N7405, N7406, N7407, N7408;
  wire N7409, N7412, N7415, N7416, N7417, N7418, N7419, N7420;
  wire N7421, N7433, N7434, N7435, N7436, N7437, N7438, N7439;
  wire N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447;
  wire N7448, N7450, N7451, N7452, N7453, N7454, N7455, N7456;
  wire N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464;
  wire N7468, N7479, N7481, N7482, N7483, N7484, N7485, N7486;
  wire N7487, N7488, N7489, N7492, N7493, N7498, N7499, N7500;
  wire N7505, N7507, N7508, N7509, N7510, N7512, N7513, N7514;
  wire N7525, N7526, N7529, N7530, N7531, N7537, N7543, N7549;
  wire N7555, N7561, N7567, N7573, N7579, N7582, N7585, N7586;
  wire N7587, N7588, N7589, N7592, N7595, N7598, N7599, N7624;
  wire N7625, N7636, N7657, N7658, N7665, N7666, N7667, N7668;
  wire N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676;
  wire N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684;
  wire N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692;
  wire N7693, N7694, N7695, N7696, N7697, N7708, N7709, N7710;
  wire N7711, N7712, N7715, N7718, N7719, N7720, N7721, N7722;
  wire N7723, N7724, N7727, N7728, N7729, N7730, N7731, N7732;
  wire N7733, N7734, N7743, N7744, N7749, N7750, N7751, N7762;
  wire N7765, N7768, N7769, N7770, N7771, N7772, N7775, N7778;
  wire N7781, N7782, N7787, N7788, N7795, N7796, N7797, N7798;
  wire N7799, N7800, N7803, N7806, N7807, N7808, N7809, N7810;
  wire N7811, N7812, N7815, N7816, N7821, N7822, N7823, N7826;
  wire N7829, N7832, N7833, N7834, N7835, N7836, N7839, N7842;
  wire N7845, N7846, N7851, N7852, N7859, N7860, N7861, N7862;
  wire N7863, N7864, N7867, N7870, N7871, N7872, N7873, N7874;
  wire N7875, N7876, N7879, N7880, N7885, N7886, N7887, N7890;
  wire N7893, N7896, N7897, N7898, N7899, N7900, N7903, N7906;
  wire N7909, N7910, N7917, N7918, N7923, N7924, N7925, N7926;
  wire N7927, N7928, N7929, N7930, N7931, N7932, N7935, N7938;
  wire N7939, N7940, N7943, N7944, N7945, N7946, N7951, N7954;
  wire N7957, N7960, N7963, N7966, N7967, N7968, N7969, N7970;
  wire N7973, N7974, N7984, N7985, N7987, N7988, N7989, N7990;
  wire N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998;
  wire N8001, N8004, N8009, N8013, N8017, N8020, N8021, N8022;
  wire N8023, N8025, N8026, N8027, N8031, N8032, N8033, N8034;
  wire N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042;
  wire N8043, N8044, N8045, N8048, N8055, N8056, N8057, N8058;
  wire N8059, N8060, N8061, N8064, N8071, N8072, N8073, N8074;
  wire N8077, N8078, N8079, N8082, N8089, N8090, N8093, N8096;
  wire N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120;
  wire N8121, N8122, N8125, N8126, n_303, n_305, n_306, n_307;
  wire n_308, n_309, n_314, n_316, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331;
  assign N-6927 = N6925;
  assign N6926 = N6924;
  assign N4278 = N4275;
  assign N3604 = N299;
  assign N3360 = N1;
  assign N3359 = N1;
  assign N3358 = N1;
  assign N3357 = N1;
  assign N2584 = N1141;
  assign N2527 = N299;
  assign N2387 = N549;
  assign N2309 = N1;
  assign N2142 = N141;
  assign N2139 = N137;
  assign N1143 = N1137;
  assign N1142 = N1137;
  assign N1066 = N592;
  assign N816 = N293;
  assign N709 = N141;
  and AND2_3 (N1042, N135, N631);
  and AND2_13 (N1140, N552, N562);
  and AND2_20 (N1147, N141, N145);
  and AND2_23 (N1150, N1043, N27);
  and AND2_24 (N1151, N386, N556);
  and AND2_71 (N1475, N27, N31);
  and AND2_192 (N2054, N136, N1148);
  and AND2_198 (N2349, N1104, N514);
  and AND2_243 (N2625, N619, N625);
  and AND2_309 (N2835, N1067, N210);
  and AND2_310 (N2836, N1067, N218);
  and AND2_311 (N2837, N1067, N226);
  and AND2_312 (N2838, N1067, N234);
  and AND2_325 (N2851, N1067, N257);
  and AND2_326 (N2852, N1067, N265);
  and AND2_327 (N2853, N1067, N273);
  and AND2_328 (N2854, N1067, N281);
  and AND2_331 (N2867, N292, N335);
  and AND2_332 (N2868, N288, N335);
  and AND2_333 (N2869, N280, N335);
  and AND2_334 (N2870, N272, N335);
  and AND2_335 (N2871, N264, N335);
  and AND2_336 (N2872, N241, N335);
  and AND2_337 (N2873, N233, N335);
  and AND2_338 (N2874, N225, N335);
  and AND2_339 (N2875, N217, N335);
  and AND2_340 (N2876, N209, N335);
  and AND2_350 (N2907, N248, N302);
  and AND2_353 (N2910, N242, N293);
  and AND2_354 (N2911, N242, N308);
  and AND2_355 (N2912, N242, N316);
  and AND2_366 (N2923, N1067, N324);
  and AND2_367 (N2924, N1067, N341);
  and AND2_368 (N2925, N1067, N351);
  and AND2_381 (N2938, N242, N257);
  and AND2_382 (N2939, N242, N265);
  and AND2_383 (N2940, N242, N273);
  and AND2_384 (N2941, N242, N281);
  and AND2_387 (N2954, N372, N332);
  and AND2_388 (N2955, N366, N332);
  and AND2_389 (N2956, N358, N332);
  and AND2_390 (N2957, N348, N332);
  and AND2_391 (N2958, N338, N332);
  and AND2_392 (N2959, N331, N332);
  and AND2_393 (N2960, N323, N332);
  and AND2_394 (N2961, N315, N332);
  and AND2_395 (N2962, N307, N332);
  and AND2_396 (N2963, N299, N332);
  and AND2_398 (N2969, N83, N1588);
  and AND2_399 (N2970, N86, N1588);
  and AND2_400 (N2971, N88, N1588);
  and AND2_409 (N2980, N248, N514);
  and AND2_412 (N2983, N242, N324);
  and AND2_414 (N2985, N242, N341);
  and AND2_415 (N2986, N242, N351);
  and AND2_434 (N3013, N248, N361);
  and AND2_448 (N3027, N242, N210);
  and AND2_449 (N3028, N242, N218);
  and AND2_450 (N3029, N242, N226);
  and AND2_451 (N3030, N242, N234);
  and AND2_462 (N3071, N97, N625);
  and AND2_463 (N3072, N94, N625);
  and AND2_499 (N3405, N1080, N2823);
  and AND2_500 (N3406, N1080, N2825);
  and AND2_501 (N3407, N1080, N2827);
  and AND2_502 (N3408, N1080, N2829);
  and AND2_507 (N3413, N1080, N2839);
  and AND2_508 (N3414, N1080, N2841);
  and AND2_509 (N3415, N1080, N2843);
  and AND2_510 (N3416, N1080, N2845);
  and AND2_511 (N3444, N251, N2902);
  and AND2_514 (N3447, N254, N2901);
  and AND2_515 (N3448, N254, N2903);
  and AND2_516 (N3449, N254, N2905);
  and AND2_520 (N3453, N1080, N1660);
  and AND2_521 (N3454, N1080, N2915);
  and AND2_522 (N3455, N1080, N2917);
  and AND2_523 (N3456, N2920, N2350);
  and AND2_528 (N3463, N254, N2839);
  and AND2_529 (N3464, N254, N2841);
  and AND2_530 (N3465, N254, N2843);
  and AND2_531 (N3466, N254, N2845);
  and AND2_536 (N3485, N254, N1660);
  and AND2_537 (N3486, N254, N2915);
  and AND2_538 (N3487, N254, N2917);
  and AND2_545 (N3502, N251, N2999);
  and AND2_551 (N3508, N254, N2823);
  and AND2_552 (N3509, N254, N2825);
  and AND2_553 (N3510, N254, N2827);
  and AND2_554 (N3511, N254, N2829);
  and AND2_573 (N3614, N1588, N2623);
  and AND2_574 (N3615, N588, N2623);
  and AND2_639 (N3680, N289, N2855);
  and AND2_640 (N3681, N281, N2855);
  and AND2_641 (N3682, N273, N2855);
  and AND2_642 (N3683, N265, N2855);
  and AND2_643 (N3684, N257, N2855);
  and AND2_644 (N3685, N234, N2855);
  and AND2_645 (N3686, N226, N2855);
  and AND2_646 (N3687, N218, N2855);
  and AND2_647 (N3688, N210, N2855);
  and AND2_648 (N3689, N206, N2855);
  and AND2_670 (N3723, N369, N2942);
  and AND2_671 (N3724, N361, N2942);
  and AND2_672 (N3725, N351, N2942);
  and AND2_673 (N3726, N341, N2942);
  and AND2_674 (N3727, N324, N2942);
  and AND2_675 (N3728, N316, N2942);
  and AND2_676 (N3729, N308, N2942);
  and AND2_677 (N3730, N302, N2942);
  and AND2_678 (N3731, N293, N2942);
  and AND2_680 (N3738, N83, N588);
  and AND2_681 (N3739, N87, N588);
  and AND2_682 (N3740, N34, N588);
  and AND2_703 (N3761, N242, N206);
  and AND2_740 (N3816, N3482, N2984);
  and AND2_792 (N3982, N254, N3753);
  and AND2_806 (N4031, N3828, N1475);
  and AND2_811 (N4036, N3829, N1475);
  and AND2_817 (N4042, N3831, N1475);
  and AND2_818 (N4067, N3732, N514);
  and AND2_820 (N4088, N3834, N3668);
  and AND2_821 (N4091, N3835, N3669);
  and AND2_822 (N4094, N3836, N3670);
  and AND2_823 (N4097, N3837, N3671);
  and AND2_824 (N4100, N3838, N3676);
  and AND2_825 (N4103, N3839, N3677);
  and AND2_826 (N4106, N3840, N3678);
  and AND2_827 (N4109, N3841, N3679);
  and AND2_828 (N4144, N3908, N3703);
  and AND2_829 (N4147, N3909, N3704);
  and AND2_831 (N4153, N3914, N3711);
  and AND2_832 (N4156, N3915, N3712);
  and AND2_833 (N4159, N3916, N3713);
  and AND2_842 (N4198, N3920, N3722);
  and AND2_853 (N4225, N3918, N3720);
  and AND2_854 (N4228, N3919, N3721);
  and AND2_855 (N4231, N3991, N3770);
  and AND2_856 (N4234, N3917, N3719);
  and AND2_857 (N4237, N3989, N3768);
  and AND2_858 (N4240, N3990, N3769);
  and AND2_859 (N4243, N3988, N3767);
  and AND2_860 (N4246, N3976, N3746);
  and AND2_861 (N4249, N3977, N3747);
  and AND2_862 (N4252, N3975, N3745);
  and AND2_868 (N4268, N446, N3893);
  and AND2_880 (N4280, N3887, N457);
  and AND2_881 (N4284, N3881, N468);
  and AND2_882 (N4290, N422, N3873);
  and AND2_883 (N4297, N3867, N435);
  and AND2_884 (N4298, N3861, N389);
  and AND2_885 (N4301, N3855, N400);
  and AND2_886 (N4305, N3849, N411);
  and AND2_887 (N4310, N3842, N374);
  and AND2_899 (N4379, N3956, N479);
  and AND2_900 (N4385, N490, N3948);
  and AND2_901 (N4392, N3942, N503);
  and AND2_902 (N4396, N3933, N523);
  and AND2_903 (N4400, N3927, N534);
  and AND2_991 (N4737, N4273, N141);
  and AND2_992 (N4738, N4274, N141);
  and AND2_993 (N4739, N4276, N141);
  and AND2_994 (N4740, N4277, N141);
  and AND2_1000 (N4939, N4515, N4185);
  and AND2_1045 (N5065, N4357, N3962);
  and AND2_1097 (N5117, N4364, N4379);
  and AND2_1099 (N5119, N54, N4405);
  and AND2_1297 (N5954, N5264, N4396);
  and AND2_1320 (N6071, N5389, N4280);
  and AND2_1330 (N6083, N5396, N4284);
  and AND2_1335 (N6088, N5407, N4290);
  and AND2_1336 (N6089, N5418, N5407);
  and AND2_1339 (N6094, N5424, N4298);
  and AND2_1343 (N6098, N5431, N4301);
  and AND2_1347 (N6102, N4305, N5441);
  and AND2_1350 (N6105, N5452, N4310);
  and AND2_1352 (N6107, N4, N5462);
  and AND2_1379 (N6138, N5462, N5452);
  and AND2_1385 (N6146, N5562, N4385);
  and AND2_1386 (N6147, N5573, N5562);
  and AND2_1389 (N6152, N5579, N4067);
  and AND2_1396 (N6159, N4400, N5595);
  and AND2_1399 (N6162, N5606, N3921);
  and AND2_1424 (N6194, N4405, N5606);
  and AND2_1546 (N6641, N6080, N6117);
  and AND2_1547 (N6643, N6140, N6149);
  and AND2_1548 (N6646, N6140, N6175);
  and AND2_1549 (N6648, N6080, N6091);
  and AND2_1560 (N6664, N6091, N4);
  and AND2_1574 (N6693, N6149, N54);
  and AND2_1621 (N6801, N6080, N6397);
  and AND2_1622 (N6802, N6427, N6140);
  and AND2_1677 (N6879, N4357, N6478);
  and AND2_1678 (N6880, N6478, N132);
  and AND2_1758 (N7040, N6817, N6079);
  and AND2_1759 (N7041, N6831, N6675);
  and AND2_1769 (N7064, N6844, N6139);
  and AND2_1770 (N7065, N6857, N6703);
  and AND2_1795 (N7125, N6817, N7018);
  and AND2_1796 (N7126, N6817, N7020);
  and AND2_1797 (N7127, N6817, N7022);
  and AND2_1800 (N7139, N6844, N7044);
  and AND2_1801 (N7140, N6844, N7046);
  and AND2_1802 (N7141, N6844, N7048);
  and AND2_1820 (N7173, N7115, N7023);
  and AND2_1821 (N7174, N7116, N7023);
  and AND2_1822 (N7175, N6940, N7023);
  and AND2_1823 (N7176, N5418, N7023);
  and AND2_1825 (N7178, N7130, N7049);
  and AND2_1826 (N7179, N7131, N7049);
  and AND2_1827 (N7180, N6958, N7049);
  and AND2_1828 (N7181, N5573, N7049);
  and AND2_1957 (N7479, N7301, N3068);
  and AND2_1975 (N7506, N7435, N137);
  and AND2_1980 (N7511, N7443, N137);
  and AND2_1997 (N7530, N7402, N3068);
  and AND2_2017 (N7600, N7505, N137);
  and AND2_2018 (N7601, N7507, N137);
  and AND2_2019 (N7602, N7508, N137);
  and AND2_2020 (N7603, N7509, N137);
  and AND2_2021 (N7604, N7510, N137);
  and AND2_2022 (N7605, N7512, N137);
  and AND2_2023 (N7606, N7513, N137);
  and AND2_2024 (N7607, N7514, N137);
  and AND2_2025 (N7624, N6979, N7489);
  and AND2_2026 (N7625, N7489, N7250);
  and AND2_2027 (N7626, N1149, N7525);
  and AND2_2109 (N7754, N7727, N137);
  and AND2_2110 (N7755, N7728, N137);
  and AND2_2111 (N7756, N7729, N137);
  and AND2_2112 (N7757, N7730, N137);
  and AND2_2113 (N7758, N7731, N137);
  and AND2_2114 (N7759, N7732, N137);
  and AND2_2115 (N7760, N7733, N137);
  and AND2_2116 (N7761, N7734, N137);
  and AND2_2254 (N8035, N583, N8025);
  and AND2_2260 (N8041, N566, N8037);
  and AND2_2262 (N8043, N8040, N1157);
  and AND2_2263 (N8044, N8042, N1219);
  and AND2_2280 (N8077, N8073, N619);
  and AND2_2281 (N8078, N8074, N619);
  and AND2_2284 (N8089, N8079, N3063);
  and AND2_2285 (N8090, N8082, N3063);
  and AND2_2304 (N8125, N8121, N137);
  and AND2_2305 (N8126, N8122, N137);
  and AND3_203 (N2585, N170, N571, N574);
  and AND3_204 (N2586, N173, N571, N574);
  and AND3_205 (N2587, N167, N571, N574);
  and AND3_206 (N2588, N164, N571, N574);
  and AND3_207 (N2589, N161, N571, N574);
  and AND3_209 (N2591, N185, N571, N574);
  and AND3_210 (N2592, N158, N571, N574);
  and AND3_211 (N2593, N152, N571, N574);
  and AND3_212 (N2594, N146, N571, N574);
  and AND3_213 (N2595, N170, N577, N580);
  and AND3_214 (N2596, N173, N577, N580);
  and AND3_215 (N2597, N167, N577, N580);
  and AND3_216 (N2598, N164, N577, N580);
  and AND3_217 (N2599, N161, N577, N580);
  and AND3_218 (N2600, N185, N577, N580);
  and AND3_219 (N2601, N158, N577, N580);
  and AND3_220 (N2602, N152, N577, N580);
  and AND3_221 (N2603, N146, N577, N580);
  and AND3_222 (N2604, N106, N613, N616);
  and AND3_223 (N2605, N61, N610, N607);
  and AND3_224 (N2606, N106, N610, N607);
  and AND3_225 (N2607, N49, N610, N607);
  and AND3_226 (N2608, N103, N610, N607);
  and AND3_227 (N2609, N40, N610, N607);
  and AND3_228 (N2610, N37, N610, N607);
  and AND3_229 (N2611, N20, N610, N607);
  and AND3_230 (N2612, N17, N610, N607);
  and AND3_231 (N2613, N70, N610, N607);
  and AND3_232 (N2614, N64, N610, N607);
  and AND3_233 (N2615, N49, N613, N616);
  and AND3_234 (N2616, N103, N613, N616);
  and AND3_235 (N2617, N40, N613, N616);
  and AND3_236 (N2618, N37, N613, N616);
  and AND3_237 (N2619, N20, N613, N616);
  and AND3_238 (N2620, N17, N613, N616);
  and AND3_239 (N2621, N70, N613, N616);
  and AND3_240 (N2622, N64, N613, N616);
  and AND3_242 (N2624, N123, N1758, N599);
  and AND3_244 (N2626, N61, N613, N616);
  and AND3_271 (N2703, N179, N571, N574);
  and AND3_292 (N2778, N179, N577, N580);
  and AND3_305 (N2831, N1104, N457, N210);
  and AND3_306 (N2832, N1104, N468, N218);
  and AND3_307 (N2833, N1104, N422, N226);
  and AND3_308 (N2834, N1104, N435, N234);
  and AND3_321 (N2847, N1104, N389, N257);
  and AND3_322 (N2848, N1104, N400, N265);
  and AND3_323 (N2849, N1104, N411, N273);
  and AND3_324 (N2850, N1104, N374, N281);
  and AND3_351 (N2908, N248, N479, N308);
  and AND3_352 (N2909, N248, N490, N316);
  and AND3_362 (N2919, N1104, N503, N324);
  and AND3_364 (N2921, N1104, N523, N341);
  and AND3_365 (N2922, N1104, N534, N351);
  and AND3_377 (N2934, N248, N389, N257);
  and AND3_378 (N2935, N248, N400, N265);
  and AND3_379 (N2936, N248, N411, N273);
  and AND3_380 (N2937, N248, N374, N281);
  and AND3_408 (N2979, N248, N503, N324);
  and AND3_410 (N2981, N248, N523, N341);
  and AND3_411 (N2982, N248, N534, N351);
  and AND3_444 (N3023, N248, N457, N210);
  and AND3_445 (N3024, N248, N468, N218);
  and AND3_446 (N3025, N248, N422, N226);
  and AND3_447 (N3026, N248, N435, N234);
  and AND3_495 (N3401, N457, N1092, N2823);
  and AND3_496 (N3402, N468, N1092, N2825);
  and AND3_497 (N3403, N422, N1092, N2827);
  and AND3_498 (N3404, N435, N1092, N2829);
  and AND3_503 (N3409, N389, N1092, N2839);
  and AND3_504 (N3410, N400, N1092, N2841);
  and AND3_505 (N3411, N411, N1092, N2843);
  and AND3_506 (N3412, N374, N1092, N2845);
  and AND3_512 (N3445, N479, N251, N2903);
  and AND3_513 (N3446, N490, N251, N2905);
  and AND3_517 (N3450, N503, N1092, N1660);
  and AND3_518 (N3451, N523, N1092, N2915);
  and AND3_519 (N3452, N534, N1092, N2917);
  and AND3_524 (N3459, N389, N251, N2839);
  and AND3_525 (N3460, N400, N251, N2841);
  and AND3_526 (N3461, N411, N251, N2843);
  and AND3_527 (N3462, N374, N251, N2845);
  and AND3_532 (N3481, N503, N251, N1660);
  and AND3_534 (N3483, N523, N251, N2915);
  and AND3_535 (N3484, N534, N251, N2917);
  and AND3_547 (N3504, N457, N251, N2823);
  and AND3_548 (N3505, N468, N251, N2825);
  and AND3_549 (N3506, N422, N251, N2827);
  and AND3_550 (N3507, N435, N251, N2829);
  and AND3_575 (N3616, N200, N2653, N574);
  and AND3_576 (N3617, N203, N2653, N574);
  and AND3_577 (N3618, N197, N2653, N574);
  and AND3_578 (N3619, N194, N2653, N574);
  and AND3_579 (N3620, N191, N2653, N574);
  and AND3_580 (N3621, N182, N2653, N574);
  and AND3_581 (N3622, N188, N2653, N574);
  and AND3_582 (N3623, N155, N2653, N574);
  and AND3_583 (N3624, N149, N2653, N574);
  and AND3_586 (N3627, N200, N2728, N580);
  and AND3_587 (N3628, N203, N2728, N580);
  and AND3_588 (N3629, N197, N2728, N580);
  and AND3_589 (N3630, N194, N2728, N580);
  and AND3_590 (N3631, N191, N2728, N580);
  and AND3_591 (N3632, N182, N2728, N580);
  and AND3_592 (N3633, N188, N2728, N580);
  and AND3_593 (N3634, N155, N2728, N580);
  and AND3_594 (N3635, N149, N2728, N580);
  and AND3_597 (N3638, N109, N2801, N616);
  and AND3_600 (N3641, N11, N2779, N607);
  and AND3_601 (N3642, N109, N2779, N607);
  and AND3_602 (N3643, N46, N2779, N607);
  and AND3_603 (N3644, N100, N2779, N607);
  and AND3_604 (N3645, N91, N2779, N607);
  and AND3_605 (N3646, N43, N2779, N607);
  and AND3_606 (N3647, N76, N2779, N607);
  and AND3_607 (N3648, N73, N2779, N607);
  and AND3_608 (N3649, N67, N2779, N607);
  and AND3_609 (N3650, N14, N2779, N607);
  and AND3_610 (N3651, N46, N2801, N616);
  and AND3_611 (N3652, N100, N2801, N616);
  and AND3_612 (N3653, N91, N2801, N616);
  and AND3_613 (N3654, N43, N2801, N616);
  and AND3_614 (N3655, N76, N2801, N616);
  and AND3_615 (N3656, N73, N2801, N616);
  and AND3_616 (N3657, N67, N2801, N616);
  and AND3_617 (N3658, N14, N2801, N616);
  and AND3_618 (N3659, N120, N3068, N625);
  and AND3_619 (N3660, N11, N2801, N616);
  and AND3_620 (N3661, N118, N3068, N625);
  and AND3_621 (N3662, N176, N2653, N574);
  and AND3_622 (N3663, N176, N2728, N580);
  and AND3_700 (N3758, N248, N446, N206);
  and AND3_717 (N3781, N117, N3068, N625);
  and AND3_718 (N3782, N126, N3068, N625);
  and AND3_719 (N3783, N127, N3068, N625);
  and AND3_720 (N3784, N128, N3068, N625);
  and AND3_721 (N3785, N131, N3068, N625);
  and AND3_722 (N3786, N129, N3068, N625);
  and AND3_723 (N3787, N119, N3068, N625);
  and AND3_724 (N3788, N130, N3068, N625);
  and AND3_728 (N3800, N122, N3068, N625);
  and AND3_729 (N3801, N113, N3068, N625);
  and AND3_730 (N3802, N53, N3068, N625);
  and AND3_731 (N3803, N114, N3068, N625);
  and AND3_732 (N3804, N115, N3068, N625);
  and AND3_733 (N3805, N52, N3068, N625);
  and AND3_734 (N3806, N112, N3068, N625);
  and AND3_735 (N3807, N116, N3068, N625);
  and AND3_736 (N3808, N121, N3068, N625);
  and AND3_737 (N3809, N123, N3068, N625);
  and AND3_790 (N3980, N446, N251, N3753);
  and AND3_800 (N3998, N3456, N3068, N3063);
  and AND3_807 (N4032, N24, N1588, N1475);
  and AND3_808 (N4033, N25, N588, N1475);
  and AND3_809 (N4034, N26, N1588, N1475);
  and AND3_810 (N4035, N81, N588, N1475);
  and AND3_812 (N4037, N79, N1588, N1475);
  and AND3_813 (N4038, N23, N588, N1475);
  and AND3_814 (N4039, N82, N1588, N1475);
  and AND3_815 (N4040, N80, N588, N1475);
  and AND3_840 (N4196, N3775, N3771, N1660);
  and AND3_841 (N4197, N3987, N3068, N3063);
  and AND3_923 (N4547, N3911, N3068, N3063);
  and AND3_995 (N4741, N3705, N1758, N1755);
  and AND3_1003 (N4953, N4188, N3775, N324);
  and AND3_1004 (N4954, N3771, N4191, N324);
  and AND3_1005 (N4955, N4191, N4188, N1660);
  and AND3_1006 (N4956, N4109, N3068, N3063);
  and AND3_1007 (N4957, N4106, N3068, N3063);
  and AND3_1008 (N4958, N4103, N3068, N3063);
  and AND3_1009 (N4959, N4100, N3068, N3063);
  and AND3_1010 (N4960, N4159, N3068, N3063);
  and AND3_1011 (N4961, N4156, N3068, N3063);
  and AND3_1022 (N4978, N3793, N3789, N3797);
  and AND3_1023 (N4979, N4203, N4200, N3797);
  and AND3_1024 (N4980, N4097, N3068, N3063);
  and AND3_1025 (N4981, N4094, N3068, N3063);
  and AND3_1026 (N4982, N4091, N3068, N3063);
  and AND3_1027 (N4983, N4088, N3068, N3063);
  and AND3_1028 (N4984, N4153, N3068, N3063);
  and AND3_1029 (N4985, N4147, N3068, N3063);
  and AND3_1030 (N4986, N4144, N3068, N3063);
  and AND3_1031 (N4987, N3705, N3068, N3063);
  and AND3_1046 (N5066, N4364, N4357, N4379);
  and AND3_1137 (N5163, N4200, N3793, N4976);
  and AND3_1138 (N5164, N3789, N4203, N4976);
  and AND3_1139 (N5165, N4939, N3068, N3063);
  and AND3_1175 (N5240, N5060, N5061, N3757);
  and AND3_1237 (N5388, N5062, N5063, N5241);
  and AND3_1321 (N6072, N5396, N5389, N4284);
  and AND3_1331 (N6084, N5407, N4290, N5396);
  and AND3_1332 (N6085, N5418, N5407, N5396);
  and AND3_1340 (N6095, N5431, N5424, N4301);
  and AND3_1344 (N6099, N5441, N4305, N5431);
  and AND3_1348 (N6103, N5452, N5441, N4310);
  and AND3_1351 (N6106, N4, N5462, N5452);
  and AND3_1374 (N6133, N5462, N5441, N5452);
  and AND3_1382 (N6143, N5562, N4385, N4364);
  and AND3_1383 (N6144, N5573, N5562, N4364);
  and AND3_1390 (N6153, N5264, N5579, N4396);
  and AND3_1393 (N6156, N5595, N4400, N5264);
  and AND3_1397 (N6160, N5606, N5595, N3921);
  and AND3_1400 (N6163, N54, N4405, N5606);
  and AND3_1419 (N6189, N4405, N5595, N5606);
  and AND3_1506 (N6473, N5315, N4524, N5319);
  and AND3_1507 (N6474, N6025, N4198, N5319);
  and AND3_1508 (N6475, N5324, N3757, N5328);
  and AND3_1509 (N6476, N6028, N3987, N5328);
  and AND3_1584 (N6712, N5696, N5692, N5700);
  and AND3_1585 (N6713, N6200, N6197, N5700);
  and AND3_1586 (N6714, N5707, N5703, N5711);
  and AND3_1587 (N6715, N6206, N6203, N5711);
  and AND3_1589 (N6718, N6164, N619, N3063);
  and AND3_1590 (N6719, N4198, N5315, N6469);
  and AND3_1591 (N6720, N4524, N6025, N6469);
  and AND3_1592 (N6721, N3987, N5324, N6471);
  and AND3_1593 (N6722, N3757, N6028, N6471);
  and AND3_1666 (N6860, N6197, N5696, N6708);
  and AND3_1667 (N6861, N5692, N6200, N6708);
  and AND3_1668 (N6862, N6203, N5707, N6710);
  and AND3_1669 (N6863, N5703, N6206, N6710);
  and AND3_1743 (N7011, N6866, N2653, N2664);
  and AND3_1744 (N7012, N6866, N2728, N2739);
  and AND3_1745 (N7013, N6866, N2779, N2790);
  and AND3_1747 (N7016, N6866, N2801, N2812);
  and AND3_1792 (N7114, N6979, N603, N1755);
  and AND3_1803 (N7146, N6932, N619, N3063);
  and AND3_1804 (N7147, N6967, N619, N3063);
  and AND3_1834 (N7187, N7037, N619, N3063);
  and AND3_1835 (N7188, N7034, N619, N3063);
  and AND3_1836 (N7189, N7031, N619, N3063);
  and AND3_1838 (N7196, N7060, N619, N3063);
  and AND3_1839 (N7197, N7057, N619, N3063);
  and AND3_1844 (N7207, N7028, N619, N3063);
  and AND3_1845 (N7208, N7054, N619, N3063);
  and AND3_1879 (N7338, N7190, N571, N2664);
  and AND3_1880 (N7339, N7198, N2653, N2664);
  and AND3_1881 (N7340, N7190, N577, N2739);
  and AND3_1882 (N7341, N7198, N2728, N2739);
  and AND3_1883 (N7342, N7190, N610, N2790);
  and AND3_1884 (N7349, N7198, N2779, N2790);
  and AND3_1885 (N7357, N7198, N2801, N2812);
  and AND3_1887 (N7364, N7190, N613, N2812);
  and AND3_1914 (N7433, N7310, N2653, N2664);
  and AND3_1915 (N7434, N7304, N571, N2664);
  and AND3_1917 (N7436, N7270, N571, N2664);
  and AND3_1918 (N7437, N7288, N2653, N2664);
  and AND3_1919 (N7438, N7276, N571, N2664);
  and AND3_1920 (N7439, N7294, N2653, N2664);
  and AND3_1921 (N7440, N7282, N571, N2664);
  and AND3_1922 (N7441, N7310, N2728, N2739);
  and AND3_1923 (N7442, N7304, N577, N2739);
  and AND3_1925 (N7444, N7270, N577, N2739);
  and AND3_1926 (N7445, N7288, N2728, N2739);
  and AND3_1927 (N7446, N7276, N577, N2739);
  and AND3_1928 (N7447, N7294, N2728, N2739);
  and AND3_1929 (N7448, N7282, N577, N2739);
  and AND3_1931 (N7450, N7310, N2779, N2790);
  and AND3_1932 (N7451, N7304, N610, N2790);
  and AND3_1933 (N7452, N7294, N2779, N2790);
  and AND3_1934 (N7453, N7282, N610, N2790);
  and AND3_1935 (N7454, N7288, N2779, N2790);
  and AND3_1936 (N7455, N7276, N610, N2790);
  and AND3_1937 (N7456, N7270, N610, N2790);
  and AND3_1938 (N7457, N7310, N2801, N2812);
  and AND3_1939 (N7458, N7304, N613, N2812);
  and AND3_1940 (N7459, N7294, N2801, N2812);
  and AND3_1941 (N7460, N7282, N613, N2812);
  and AND3_1942 (N7461, N7288, N2801, N2812);
  and AND3_1943 (N7462, N7276, N613, N2812);
  and AND3_1944 (N7463, N7270, N613, N2812);
  and AND3_1945 (N7464, N7250, N603, N599);
  and AND3_1958 (N7481, N7245, N619, N3063);
  and AND3_1959 (N7482, N7242, N619, N3063);
  and AND3_1960 (N7483, N7239, N619, N3063);
  and AND3_1961 (N7484, N7236, N619, N3063);
  and AND3_1962 (N7485, N7263, N619, N3063);
  and AND3_1963 (N7486, N7260, N619, N3063);
  and AND3_1964 (N7487, N7257, N619, N3063);
  and AND3_1965 (N7488, N7250, N619, N3063);
  and AND3_1993 (N7526, N7468, N3068, N3063);
  and AND3_2029 (N7636, N7529, N3068, N3063);
  and AND3_2033 (N7666, N7555, N2653, N2664);
  and AND3_2034 (N7667, N7531, N571, N2664);
  and AND3_2035 (N7668, N7561, N2653, N2664);
  and AND3_2036 (N7669, N7537, N571, N2664);
  and AND3_2037 (N7670, N7567, N2653, N2664);
  and AND3_2038 (N7671, N7543, N571, N2664);
  and AND3_2039 (N7672, N7573, N2653, N2664);
  and AND3_2040 (N7673, N7549, N571, N2664);
  and AND3_2041 (N7674, N7555, N2728, N2739);
  and AND3_2042 (N7675, N7531, N577, N2739);
  and AND3_2043 (N7676, N7561, N2728, N2739);
  and AND3_2044 (N7677, N7537, N577, N2739);
  and AND3_2045 (N7678, N7567, N2728, N2739);
  and AND3_2046 (N7679, N7543, N577, N2739);
  and AND3_2047 (N7680, N7573, N2728, N2739);
  and AND3_2048 (N7681, N7549, N577, N2739);
  and AND3_2049 (N7682, N7573, N2801, N2812);
  and AND3_2050 (N7683, N7549, N613, N2812);
  and AND3_2051 (N7684, N7573, N2779, N2790);
  and AND3_2052 (N7685, N7549, N610, N2790);
  and AND3_2053 (N7686, N7567, N2779, N2790);
  and AND3_2054 (N7687, N7543, N610, N2790);
  and AND3_2055 (N7688, N7561, N2779, N2790);
  and AND3_2056 (N7689, N7537, N610, N2790);
  and AND3_2057 (N7690, N7555, N2779, N2790);
  and AND3_2058 (N7691, N7531, N610, N2790);
  and AND3_2059 (N7692, N7567, N2801, N2812);
  and AND3_2060 (N7693, N7543, N613, N2812);
  and AND3_2061 (N7694, N7561, N2801, N2812);
  and AND3_2062 (N7695, N7537, N613, N2812);
  and AND3_2063 (N7696, N7555, N2801, N2812);
  and AND3_2064 (N7697, N7531, N613, N2812);
  and AND3_2227 (N7988, N7957, N6831, N1157);
  and AND3_2228 (N7989, N7954, N6397, N1157);
  and AND3_2229 (N7990, N7957, N7041, N566);
  and AND3_2230 (N7991, N7954, N7177, N566);
  and AND3_2233 (N7994, N7963, N6857, N1219);
  and AND3_2234 (N7995, N7960, N6427, N1219);
  and AND3_2235 (N7996, N7963, N7065, N583);
  and AND3_2236 (N7997, N7960, N7182, N583);
  and AND3_2274 (N8071, N8064, N619, N3063);
  and AND3_2275 (N8072, N8061, N619, N3063);
  and AND3_2292 (N8113, N8096, N2779, N2790);
  and AND3_2293 (N8114, N8093, N610, N2790);
  and AND3_2294 (N8115, N8096, N2801, N2812);
  and AND3_2295 (N8116, N8093, N613, N2812);
  and AND3_2296 (N8117, N8096, N2653, N2664);
  and AND3_2297 (N8118, N8093, N571, N2664);
  and AND3_2298 (N8119, N8096, N2728, N2739);
  and AND3_2299 (N8120, N8093, N577, N2739);
  and AND4_1041 (N5060, N4724, N4725, N3700, N4027);
  and AND4_1042 (N5061, N4726, N4727, N3827, N4728);
  and AND4_1043 (N5062, N4729, N4730, N4731, N4732);
  and AND4_1044 (N5063, N4733, N4734, N4735, N4736);
  and AND4_1322 (N6073, N5407, N5389, N4290, N5396);
  and AND4_1323 (N6074, N5562, N4357, N4385, N4364);
  and AND4_1329 (N6080, N5396, N5418, N5407, N5389);
  and AND4_1341 (N6096, N5441, N5424, N4305, N5431);
  and AND4_1345 (N6100, N5452, N5441, N4310, N5431);
  and AND4_1349 (N6104, N4, N5462, N5441, N5452);
  and AND4_1368 (N6127, N5462, N5441, N5431, N5452);
  and AND4_1381 (N6140, N4364, N5573, N5562, N4357);
  and AND4_1391 (N6154, N5595, N5579, N4400, N5264);
  and AND4_1394 (N6157, N5606, N5595, N3921, N5264);
  and AND4_1398 (N6161, N54, N4405, N5595, N5606);
  and AND4_1414 (N6184, N4405, N5595, N5264, N5606);
  nand NAND2_19 (N1146, N373, N1);
  nand NAND2_208 (N2590, N1475, N140);
  nand NAND2_555 (N3512, N369, N2999);
  nand NAND2_556 (N3513, N361, N3032);
  nand NAND2_557 (N3514, N351, N2915);
  nand NAND2_558 (N3515, N341, N2917);
  nand NAND2_559 (N3558, N289, N2845);
  nand NAND2_560 (N3559, N281, N3142);
  nand NAND2_561 (N3560, N273, N2841);
  nand NAND2_562 (N3561, N265, N2843);
  nand NAND2_563 (N3562, N257, N2829);
  nand NAND2_564 (N3563, N234, N2839);
  nand NAND2_566 (N3605, N316, N2903);
  nand NAND2_567 (N3606, N308, N2905);
  nand NAND2_568 (N3607, N302, N2901);
  nand NAND2_569 (N3608, N293, N2902);
  nand NAND2_570 (N3609, N226, N2825);
  nand NAND2_571 (N3610, N218, N2827);
  nand NAND2_713 (N3771, N3512, N3513);
  nand NAND2_714 (N3775, N3514, N3515);
  nand NAND2_725 (N3789, N3558, N3559);
  nand NAND2_726 (N3793, N3560, N3561);
  nand NAND2_727 (N3797, N3562, N3563);
  nand NAND2_738 (N3810, N3607, N3608);
  nand NAND2_739 (N3813, N3605, N3606);
  nand NAND2_743 (N3823, N206, N2823);
  nand NAND2_744 (N3824, N3609, N3610);
  nand NAND2_804 (N4024, N210, N3753);
  nand NAND2_866 (N4264, N4024, N3823);
  nand NAND2_974 (N4701, N3813, N4223);
  nand NAND2_975 (N4702, N3810, N4224);
  nand NAND2_977 (N4721, N3911, N4027);
  nand NAND2_997 (N4856, N3732, N2712);
  nand NAND2_1019 (N4975, N4252, N4199);
  nand NAND2_1032 (N5049, N4701, N4702);
  nand NAND2_1038 (N5057, N3705, N3700);
  nand NAND2_1040 (N5059, N4264, N4267);
  nand NAND2_1050 (N5070, N3893, N2628);
  nand NAND2_1052 (N5072, N3887, N2629);
  nand NAND2_1054 (N5074, N3881, N2630);
  nand NAND2_1056 (N5076, N3873, N2631);
  nand NAND2_1058 (N5078, N3867, N2632);
  nand NAND2_1060 (N5080, N3861, N2633);
  nand NAND2_1062 (N5082, N3855, N2634);
  nand NAND2_1064 (N5084, N3849, N2635);
  nand NAND2_1066 (N5086, N3842, N2636);
  nand NAND2_1087 (N5107, N3956, N2709);
  nand NAND2_1089 (N5109, N3948, N2710);
  nand NAND2_1091 (N5111, N3942, N2711);
  nand NAND2_1092 (N5112, N514, N4855);
  nand NAND2_1094 (N5114, N3933, N2713);
  nand NAND2_1096 (N5116, N3927, N2714);
  nand NAND2_1116 (N5137, N3921, N4521);
  nand NAND2_1119 (N5140, N3942, N4855);
  nand NAND2_1124 (N5145, N3893, N4523);
  nand NAND2_1129 (N5153, N4228, N4965);
  nand NAND2_1130 (N5154, N4225, N4966);
  nand NAND2_1131 (N5155, N4234, N4967);
  nand NAND2_1132 (N5156, N4231, N4968);
  nand NAND2_1134 (N5160, N4249, N4972);
  nand NAND2_1135 (N5161, N4246, N4973);
  nand NAND2_1136 (N5162, N3816, N4974);
  nand NAND2_1169 (N5232, N4240, N5052);
  nand NAND2_1170 (N5233, N4237, N5053);
  nand NAND2_1171 (N5234, N4147, N4725);
  nand NAND2_1172 (N5235, N4144, N4724);
  nand NAND2_1173 (N5236, N4721, N5057);
  nand NAND2_1174 (N5239, N3824, N5058);
  nand NAND2_1177 (N5242, N446, N5069);
  nand NAND2_1178 (N5243, N457, N5071);
  nand NAND2_1179 (N5244, N468, N5073);
  nand NAND2_1180 (N5245, N422, N5075);
  nand NAND2_1181 (N5246, N435, N5077);
  nand NAND2_1182 (N5247, N389, N5079);
  nand NAND2_1183 (N5248, N400, N5081);
  nand NAND2_1184 (N5249, N411, N5083);
  nand NAND2_1185 (N5250, N374, N5085);
  nand NAND2_1195 (N5261, N479, N5106);
  nand NAND2_1196 (N5262, N490, N5108);
  nand NAND2_1197 (N5263, N503, N5110);
  nand NAND2_1198 (N5264, N5112, N4856);
  nand NAND2_1199 (N5274, N523, N5113);
  nand NAND2_1200 (N5275, N534, N5115);
  nand NAND2_1207 (N5303, N3933, N5115);
  nand NAND2_1208 (N5304, N3927, N5113);
  nand NAND2_1209 (N5305, N4008, N4405);
  nand NAND2_1210 (N5306, N3732, N5110);
  nand NAND2_1211 (N5307, N3867, N5075);
  nand NAND2_1212 (N5308, N3873, N5077);
  nand NAND2_1213 (N5309, N3881, N5071);
  nand NAND2_1214 (N5310, N3887, N5073);
  nand NAND2_1215 (N5311, N4011, N5069);
  nand NAND2_1217 (N5315, N5153, N5154);
  nand NAND2_1218 (N5319, N5155, N5156);
  nand NAND2_1219 (N5324, N5160, N5161);
  nand NAND2_1220 (N5328, N5162, N4975);
  nand NAND2_1224 (N5363, N3948, N5106);
  nand NAND2_1225 (N5364, N3956, N5108);
  nand NAND2_1227 (N5366, N3968, N4364);
  nand NAND2_1228 (N5367, N3842, N5083);
  nand NAND2_1229 (N5368, N3849, N5085);
  nand NAND2_1230 (N5369, N3855, N5079);
  nand NAND2_1231 (N5370, N3861, N5081);
  nand NAND2_1232 (N5371, N5148, N5147);
  nand NAND2_1234 (N5377, N5232, N5233);
  nand NAND2_1235 (N5382, N5234, N5235);
  nand NAND2_1236 (N5385, N5239, N5059);
  nand NAND2_1238 (N5389, N5242, N5070);
  nand NAND2_1239 (N5396, N5243, N5072);
  nand NAND2_1240 (N5407, N5244, N5074);
  nand NAND2_1241 (N5418, N5245, N5076);
  nand NAND2_1242 (N5424, N5246, N5078);
  nand NAND2_1243 (N5431, N5247, N5080);
  nand NAND2_1244 (N5441, N5248, N5082);
  nand NAND2_1245 (N5452, N5249, N5084);
  nand NAND2_1246 (N5462, N5250, N5086);
  nand NAND2_1257 (N5562, N5261, N5107);
  nand NAND2_1258 (N5573, N5262, N5109);
  nand NAND2_1259 (N5579, N5263, N5111);
  nand NAND2_1260 (N5595, N5274, N5114);
  nand NAND2_1261 (N5606, N5275, N5116);
  nand NAND2_1262 (N5616, N4405, N2715);
  nand NAND2_1276 (N5692, N5303, N5304);
  nand NAND2_1277 (N5696, N5137, N5305);
  nand NAND2_1278 (N5700, N5306, N5140);
  nand NAND2_1279 (N5703, N5307, N5308);
  nand NAND2_1280 (N5707, N5309, N5310);
  nand NAND2_1281 (N5711, N5145, N5311);
  nand NAND2_1291 (N5736, N5365, N5366);
  nand NAND2_1292 (N5739, N5363, N5364);
  nand NAND2_1293 (N5742, N5369, N5370);
  nand NAND2_1294 (N5745, N5367, N5368);
  nand NAND2_1296 (N5756, N5332, N5331);
  nand NAND2_1298 (N5955, N54, N3921);
  nand NAND2_1303 (N6024, N5371, N5312);
  nand NAND2_1316 (N6066, N4939, N5054);
  nand NAND2_1319 (N6069, N5382, N5755);
  nand NAND2_1401 (N6164, N5616, N5955);
  nand NAND2_1433 (N6221, N5049, N6023);
  nand NAND2_1435 (N6235, N5756, N6044);
  nand NAND2_1484 (N6377, N4243, N5241);
  nand NAND2_1485 (N6378, N5236, N6068);
  nand NAND2_1501 (N6716, N6221, N6024);
  nand NAND2_1510 (N6477, N5385, N6234);
  nand NAND2_1511 (N6478, N4357, N132);
  nand NAND2_1539 (N6630, N5739, N6373);
  nand NAND2_1540 (N6631, N5736, N6374);
  nand NAND2_1541 (N6632, N5745, N6375);
  nand NAND2_1542 (N6633, N5742, N6376);
  nand NAND2_1543 (N6634, N6377, N6066);
  nand NAND2_1544 (N6637, N6069, N6378);
  nand NAND2_1550 (N6650, N5462, N2637);
  nand NAND2_1556 (N6660, N5407, N5087);
  nand NAND2_1558 (N6662, N5407, N5469);
  nand NAND2_1570 (N6689, N5562, N5120);
  nand NAND2_1572 (N6691, N5562, N5622);
  nand NAND2_1577 (N6699, N5606, N5956);
  nand NAND2_1594 (N6877, N6477, N6235);
  nand NAND2_1619 (N6792, N6630, N6631);
  nand NAND2_1620 (N6795, N6632, N6633);
  nand NAND2_1626 (N6806, N4, N6651);
  nand NAND2_1628 (N6808, N6482, N6653);
  nand NAND2_1630 (N6810, N6486, N6653);
  nand NAND2_1632 (N6812, N6490, N6657);
  nand NAND2_1634 (N6814, N6494, N6657);
  nand NAND2_1635 (N6815, N4575, N6661);
  nand NAND2_1636 (N6816, N4290, N6661);
  nand NAND2_1639 (N6824, N6500, N6666);
  nand NAND2_1641 (N6826, N6504, N6668);
  nand NAND2_1643 (N6828, N6508, N6670);
  nand NAND2_1645 (N6830, N6512, N6672);
  nand NAND2_1648 (N6835, N6566, N3968);
  nand NAND2_1650 (N6837, N6569, N3968);
  nand NAND2_1652 (N6839, N6572, N3962);
  nand NAND2_1654 (N6841, N6575, N3962);
  nand NAND2_1655 (N6842, N4627, N6690);
  nand NAND2_1656 (N6843, N4385, N6690);
  nand NAND2_1659 (N6851, N6580, N6695);
  nand NAND2_1661 (N6853, N6584, N6434);
  nand NAND2_1663 (N6855, N6587, N6698);
  nand NAND2_1664 (N6856, N5346, N6700);
  nand NAND2_1684 (N6890, N6536, N5176);
  nand NAND2_1688 (N6896, N6553, N5728);
  nand NAND2_1699 (N6915, N6619, N4405);
  nand NAND2_1703 (N6923, N6634, N6067);
  nand NAND2_1709 (N6932, N6650, N6806);
  nand NAND2_1710 (N6935, N5389, N6807);
  nand NAND2_1711 (N6936, N5389, N6809);
  nand NAND2_1712 (N6937, N5396, N6811);
  nand NAND2_1713 (N6938, N5396, N6411);
  nand NAND2_1714 (N6939, N6660, N6815);
  nand NAND2_1715 (N6940, N6662, N6816);
  nand NAND2_1716 (N6946, N5424, N6823);
  nand NAND2_1717 (N6947, N5431, N6825);
  nand NAND2_1718 (N6948, N5441, N6827);
  nand NAND2_1719 (N6949, N5452, N6829);
  nand NAND2_1720 (N6953, N4357, N6834);
  nand NAND2_1721 (N6954, N4357, N6836);
  nand NAND2_1722 (N6955, N4364, N6838);
  nand NAND2_1723 (N6956, N4364, N6437);
  nand NAND2_1724 (N6957, N6689, N6842);
  nand NAND2_1725 (N6958, N6691, N6843);
  nand NAND2_1726 (N6964, N5579, N6850);
  nand NAND2_1727 (N6965, N5264, N6852);
  nand NAND2_1728 (N6966, N5595, N6854);
  nand NAND2_1729 (N6967, N6699, N6856);
  nand NAND2_1737 (N6987, N4608, N6889);
  nand NAND2_1738 (N6990, N4310, N6895);
  nand NAND2_1739 (N6999, N3921, N6914);
  nand NAND2_1740 (N7002, N5377, N6922);
  nand NAND2_1741 (N7003, N6873, N6872);
  nand NAND2_1742 (N7006, N6875, N6874);
  nand NAND2_1748 (N7018, N6935, N6808);
  nand NAND2_1749 (N7019, N6936, N6810);
  nand NAND2_1750 (N7020, N6937, N6812);
  nand NAND2_1751 (N7021, N6938, N6814);
  nand NAND2_1754 (N7028, N6946, N6824);
  nand NAND2_1755 (N7031, N6947, N6826);
  nand NAND2_1756 (N7034, N6948, N6828);
  nand NAND2_1757 (N7037, N6949, N6830);
  nand NAND2_1760 (N7044, N6953, N6835);
  nand NAND2_1761 (N7045, N6954, N6837);
  nand NAND2_1762 (N7046, N6955, N6839);
  nand NAND2_1763 (N7047, N6956, N6841);
  nand NAND2_1766 (N7054, N6964, N6851);
  nand NAND2_1767 (N7057, N6965, N6853);
  nand NAND2_1768 (N7060, N6966, N6855);
  nand NAND2_1772 (N7073, N6881, N5087);
  nand NAND2_1774 (N7075, N6494, N5469);
  nand NAND2_1775 (N7076, N6890, N6987);
  nand NAND2_1777 (N7080, N6896, N6990);
  nand NAND2_1780 (N7085, N6901, N5120);
  nand NAND2_1782 (N7087, N6575, N5622);
  nand NAND2_1784 (N7089, N6909, N6912);
  nand NAND2_1785 (N7090, N6915, N6999);
  nand NAND2_1787 (N7094, N6974, N6973);
  nand NAND2_1788 (N7097, N6976, N6975);
  nand NAND2_1789 (N7101, N7002, N6923);
  nand NAND2_1807 (N7151, N7006, N6876);
  nand NAND2_1808 (N7152, N4575, N7072);
  nand NAND2_1809 (N7153, N4290, N6411);
  nand NAND2_1810 (N7158, N4627, N7084);
  nand NAND2_1811 (N7159, N4385, N6437);
  nand NAND2_1812 (N7160, N6606, N7088);
  nand NAND2_1831 (N7184, N7094, N6977);
  nand NAND2_1833 (N7186, N7097, N6978);
  nand NAND2_1841 (N7204, N7101, N7149);
  nand NAND2_1843 (N7206, N6637, N7150);
  nand NAND2_1846 (N7209, N7073, N7152);
  nand NAND2_1847 (N7212, N7075, N7153);
  nand NAND2_1849 (N7216, N7076, N7079);
  nand NAND2_1851 (N7218, N7080, N6419);
  nand NAND2_1852 (N7219, N7085, N7158);
  nand NAND2_1853 (N7222, N7087, N7159);
  nand NAND2_1854 (N7225, N7089, N7160);
  nand NAND2_1856 (N7229, N7090, N6445);
  nand NAND2_1865 (N7268, N6792, N7183);
  nand NAND2_1866 (N7269, N6795, N7185);
  nand NAND2_1872 (N7300, N7003, N7205);
  nand NAND2_1873 (N7301, N7206, N7151);
  nand NAND2_1876 (N7320, N6891, N7215);
  nand NAND2_1877 (N7321, N6897, N7217);
  nand NAND2_1878 (N7328, N6916, N7228);
  nand NAND2_1889 (N7474, N7268, N7184);
  nand NAND2_1890 (N7476, N7269, N7186);
  nand NAND2_1891 (N7402, N7204, N7300);
  nand NAND2_1893 (N7406, N7209, N6807);
  nand NAND2_1895 (N7408, N7212, N6809);
  nand NAND2_1896 (N7409, N7320, N7216);
  nand NAND2_1897 (N7412, N7321, N7218);
  nand NAND2_1899 (N7416, N7219, N6834);
  nand NAND2_1901 (N7418, N7222, N6836);
  nand NAND2_1903 (N7420, N7225, N6913);
  nand NAND2_1904 (N7421, N7328, N7229);
  nand NAND2_1966 (N7489, N6979, N7250);
  nand NAND2_1967 (N7492, N6482, N7405);
  nand NAND2_1968 (N7493, N6486, N7407);
  nand NAND2_1969 (N7498, N6566, N7415);
  nand NAND2_1970 (N7499, N6569, N7417);
  nand NAND2_1971 (N7500, N6609, N7419);
  nand NAND2_2006 (N7579, N7492, N7406);
  nand NAND2_2007 (N7582, N7493, N7408);
  nand NAND2_2009 (N7586, N7409, N6894);
  nand NAND2_2011 (N7588, N7412, N6900);
  nand NAND2_2012 (N7589, N7498, N7416);
  nand NAND2_2013 (N7592, N7499, N7418);
  nand NAND2_2014 (N7595, N7500, N7420);
  nand NAND2_2016 (N7599, N7421, N6919);
  nand NAND2_2030 (N7657, N6539, N7585);
  nand NAND2_2031 (N7658, N6556, N7587);
  nand NAND2_2032 (N7665, N6622, N7598);
  nand NAND2_2076 (N7709, N7579, N6079);
  nand NAND2_2078 (N7711, N7582, N6079);
  nand NAND2_2079 (N7712, N7657, N7586);
  nand NAND2_2080 (N7715, N7658, N7588);
  nand NAND2_2082 (N7719, N7589, N6139);
  nand NAND2_2084 (N7721, N7592, N6139);
  nand NAND2_2086 (N7723, N7595, N3921);
  nand NAND2_2087 (N7724, N7665, N7599);
  nand NAND2_2104 (N7743, N5418, N7708);
  nand NAND2_2105 (N7744, N5418, N7710);
  nand NAND2_2106 (N7749, N5573, N7718);
  nand NAND2_2107 (N7750, N5573, N7720);
  nand NAND2_2108 (N7751, N4405, N7722);
  nand NAND2_2117 (N7762, N7743, N7709);
  nand NAND2_2118 (N7765, N7744, N7711);
  nand NAND2_2120 (N7769, N7712, N6651);
  nand NAND2_2122 (N7771, N7715, N6651);
  nand NAND2_2123 (N7772, N7749, N7719);
  nand NAND2_2124 (N7775, N7750, N7721);
  nand NAND2_2125 (N7778, N7751, N7723);
  nand NAND2_2127 (N7782, N7724, N3921);
  nand NAND2_2128 (N7787, N5462, N7768);
  nand NAND2_2129 (N7788, N5462, N7770);
  nand NAND2_2130 (N7795, N4405, N7781);
  nand NAND2_2132 (N7797, N7762, N6661);
  nand NAND2_2134 (N7799, N7765, N6661);
  nand NAND2_2135 (N7800, N7787, N7769);
  nand NAND2_2136 (N7803, N7788, N7771);
  nand NAND2_2138 (N7807, N7772, N6690);
  nand NAND2_2140 (N7809, N7775, N6690);
  nand NAND2_2142 (N7811, N7778, N6700);
  nand NAND2_2143 (N7812, N7795, N7782);
  nand NAND2_2144 (N7815, N5407, N7796);
  nand NAND2_2145 (N7816, N5407, N7798);
  nand NAND2_2146 (N7821, N5562, N7806);
  nand NAND2_2147 (N7822, N5562, N7808);
  nand NAND2_2148 (N7823, N5606, N7810);
  nand NAND2_2149 (N7826, N7815, N7797);
  nand NAND2_2150 (N7829, N7816, N7799);
  nand NAND2_2152 (N7833, N7800, N6672);
  nand NAND2_2154 (N7835, N7803, N6672);
  nand NAND2_2155 (N7836, N7821, N7807);
  nand NAND2_2156 (N7839, N7822, N7809);
  nand NAND2_2157 (N7842, N7823, N7811);
  nand NAND2_2159 (N7846, N7812, N6700);
  nand NAND2_2160 (N7851, N5452, N7832);
  nand NAND2_2161 (N7852, N5452, N7834);
  nand NAND2_2162 (N7859, N5606, N7845);
  nand NAND2_2164 (N7861, N7826, N6653);
  nand NAND2_2166 (N7863, N7829, N6653);
  nand NAND2_2167 (N7864, N7851, N7833);
  nand NAND2_2168 (N7867, N7852, N7835);
  nand NAND2_2170 (N7871, N7836, N3968);
  nand NAND2_2172 (N7873, N7839, N3968);
  nand NAND2_2174 (N7875, N7842, N6695);
  nand NAND2_2175 (N7876, N7859, N7846);
  nand NAND2_2176 (N7879, N5389, N7860);
  nand NAND2_2177 (N7880, N5389, N7862);
  nand NAND2_2178 (N7885, N4357, N7870);
  nand NAND2_2179 (N7886, N4357, N7872);
  nand NAND2_2180 (N7887, N5579, N7874);
  nand NAND2_2181 (N7890, N7879, N7861);
  nand NAND2_2182 (N7893, N7880, N7863);
  nand NAND2_2184 (N7897, N7864, N6666);
  nand NAND2_2186 (N7899, N7867, N6666);
  nand NAND2_2187 (N7900, N7885, N7871);
  nand NAND2_2188 (N7903, N7886, N7873);
  nand NAND2_2189 (N7906, N7887, N7875);
  nand NAND2_2191 (N7910, N7876, N6695);
  nand NAND2_2192 (N7917, N5424, N7896);
  nand NAND2_2193 (N7918, N5424, N7898);
  nand NAND2_2194 (N7923, N5579, N7909);
  nand NAND2_2196 (N7925, N7890, N6657);
  nand NAND2_2198 (N7927, N7893, N6657);
  nand NAND2_2200 (N7929, N7900, N3962);
  nand NAND2_2202 (N7931, N7903, N3962);
  nand NAND2_2203 (N7932, N7917, N7897);
  nand NAND2_2204 (N7935, N7918, N7899);
  nand NAND2_2206 (N7939, N7906, N6698);
  nand NAND2_2207 (N7940, N7923, N7910);
  nand NAND2_2208 (N7943, N5396, N7924);
  nand NAND2_2209 (N7944, N5396, N7926);
  nand NAND2_2210 (N7945, N4364, N7928);
  nand NAND2_2211 (N7946, N4364, N7930);
  nand NAND2_2212 (N7951, N5595, N7938);
  nand NAND2_2213 (N7954, N7943, N7925);
  nand NAND2_2214 (N7957, N7944, N7927);
  nand NAND2_2215 (N7960, N7945, N7929);
  nand NAND2_2216 (N7963, N7946, N7931);
  nand NAND2_2218 (N7967, N7932, N6670);
  nand NAND2_2220 (N7969, N7935, N6670);
  nand NAND2_2221 (N7970, N7951, N7939);
  nand NAND2_2223 (N7974, N7940, N6698);
  nand NAND2_2224 (N7984, N5441, N7966);
  nand NAND2_2225 (N7985, N5441, N7968);
  nand NAND2_2226 (N7987, N5595, N7973);
  nand NAND2_2232 (N7993, N7970, N6434);
  nand NAND2_2237 (N7998, N7984, N7967);
  nand NAND2_2238 (N8001, N7985, N7969);
  nand NAND2_2239 (N8004, N7987, N7974);
  nand NAND2_2240 (N8009, N5264, N7992);
  nand NAND2_2244 (N8021, N7998, N6668);
  nand NAND2_2246 (N8023, N8001, N6668);
  nand NAND2_2247 (N8025, N8009, N7993);
  nand NAND2_2249 (N8027, N8004, N6434);
  nand NAND2_2250 (N8031, N5431, N8020);
  nand NAND2_2251 (N8032, N5431, N8022);
  nand NAND2_2253 (N8034, N5264, N8026);
  nand NAND2_2256 (N8037, N8031, N8021);
  nand NAND2_2257 (N8038, N8032, N8023);
  nand NAND2_2258 (N8039, N8034, N8027);
  nand NAND2_2266 (N8055, N8045, N8033);
  nand NAND2_2268 (N8057, N8048, N8036);
  nand NAND2_2270 (N8059, N8013, N8056);
  nand NAND2_2271 (N8060, N8017, N8058);
  nand NAND2_2272 (N8061, N8055, N8059);
  nand NAND2_2273 (N8064, N8057, N8060);
  nor NOR2_933 (N4575, N422, N3873);
  nor NOR2_944 (N4608, N374, N3842);
  nor NOR2_950 (N4627, N490, N3948);
  nor NOR2_1126 (N5147, N4953, N4196);
  nor NOR2_1127 (N5148, N4954, N4955);
  nor NOR2_1221 (N5331, N5163, N4978);
  nor NOR2_1222 (N5332, N5164, N4979);
  nor NOR2_1515 (N6494, N4284, N6088);
  nor NOR2_1529 (N6575, N4379, N6146);
  nor NOR2_1671 (N6872, N6719, N6473);
  nor NOR2_1672 (N6873, N6720, N6474);
  nor NOR2_1673 (N6874, N6721, N6475);
  nor NOR2_1674 (N6875, N6722, N6476);
  nor NOR2_1730 (N6973, N6860, N6712);
  nor NOR2_1731 (N6974, N6861, N6713);
  nor NOR2_1732 (N6975, N6862, N6714);
  nor NOR2_1733 (N6976, N6863, N6715);
  nor NOR3_1513 (N6486, N4280, N6083, N6084);
  nor NOR3_1524 (N6553, N4301, N6102, N6103);
  nor NOR3_1527 (N6569, N3962, N5117, N6143);
  nor NOR3_1537 (N6619, N4396, N6159, N6160);
  nor NOR4_1525 (N6556, N4298, N6098, N6099, N6100);
  nor NOR4_1538 (N6622, N4067, N5954, N6156, N6157);
  not NOT1_4 (N1043, N591);
  not NOT1_6 (N1067, N595);
  not NOT1_7 (N1080, N596);
  not NOT1_8 (N1092, N597);
  not NOT1_9 (N1104, N598);
  not NOT1_10 (N1137, N545);
  not NOT1_11 (N1138, N348);
  not NOT1_12 (N1139, N366);
  not NOT1_14 (N1141, N549);
  not NOT1_17 (N1144, N338);
  not NOT1_18 (N1145, N358);
  not NOT1_21 (N1148, N592);
  not NOT1_22 (N1149, N1042);
  not NOT1_25 (N1152, N245);
  not NOT1_26 (N1153, N552);
  not NOT1_27 (N1154, N562);
  not NOT1_28 (N1155, N559);
  not NOT1_30 (N1157, N566);
  not NOT1_38 (N1219, N583);
  not NOT1_98 (N1588, N588);
  not NOT1_121 (N1660, N324);
  not NOT1_131 (N1755, N599);
  not NOT1_132 (N1758, N603);
  not NOT1_191 (N1972, N1146);
  not NOT1_193 (N2060, N1150);
  not NOT1_194 (N2061, N1151);
  not NOT1_241 (N2623, N1475);
  not NOT1_246 (N2628, N446);
  not NOT1_247 (N2629, N457);
  not NOT1_248 (N2630, N468);
  not NOT1_249 (N2631, N422);
  not NOT1_250 (N2632, N435);
  not NOT1_251 (N2633, N389);
  not NOT1_252 (N2634, N400);
  not NOT1_253 (N2635, N411);
  not NOT1_254 (N2636, N374);
  not NOT1_255 (N2637, N4);
  not NOT1_266 (N2653, N571);
  not NOT1_267 (N2664, N574);
  not NOT1_273 (N2709, N479);
  not NOT1_274 (N2710, N490);
  not NOT1_275 (N2711, N503);
  not NOT1_276 (N2712, N514);
  not NOT1_277 (N2713, N523);
  not NOT1_278 (N2714, N534);
  not NOT1_279 (N2715, N54);
  not NOT1_287 (N2728, N577);
  not NOT1_288 (N2739, N580);
  not NOT1_293 (N2779, N610);
  not NOT1_294 (N2790, N607);
  not NOT1_295 (N2801, N613);
  not NOT1_296 (N2812, N616);
  not NOT1_297 (N2823, N210);
  not NOT1_299 (N2825, N218);
  not NOT1_301 (N2827, N226);
  not NOT1_303 (N2829, N234);
  not NOT1_313 (N2839, N257);
  not NOT1_315 (N2841, N265);
  not NOT1_317 (N2843, N273);
  not NOT1_319 (N2845, N281);
  not NOT1_329 (N2855, N335);
  not NOT1_344 (N2901, N293);
  not NOT1_345 (N2902, N302);
  not NOT1_346 (N2903, N308);
  not NOT1_348 (N2905, N316);
  not NOT1_358 (N2915, N341);
  not NOT1_360 (N2917, N351);
  not NOT1_363 (N2920, N2349);
  not NOT1_385 (N2942, N332);
  not NOT1_428 (N2999, N361);
  not NOT1_453 (N3032, N369);
  not NOT1_460 (N3063, N625);
  not NOT1_461 (N3068, N619);
  not NOT1_473 (N3142, N289);
  not NOT1_533 (N3482, N2980);
  not NOT1_572 (N3613, N299);
  not NOT1_695 (N3753, N206);
  not NOT1_745 (N3827, N3456);
  not NOT1_750 (N3834, N3664);
  not NOT1_751 (N3835, N3665);
  not NOT1_752 (N3836, N3666);
  not NOT1_753 (N3837, N3667);
  not NOT1_754 (N3838, N3672);
  not NOT1_755 (N3839, N3673);
  not NOT1_756 (N3840, N3674);
  not NOT1_757 (N3841, N3675);
  not NOT1_767 (N3908, N3701);
  not NOT1_768 (N3909, N3702);
  not NOT1_769 (N3911, N3700);
  not NOT1_770 (N3914, N3708);
  not NOT1_771 (N3915, N3709);
  not NOT1_772 (N3916, N3710);
  not NOT1_773 (N3917, N3715);
  not NOT1_774 (N3918, N3716);
  not NOT1_775 (N3919, N3717);
  not NOT1_776 (N3920, N3718);
  not NOT1_785 (N3975, N3742);
  not NOT1_786 (N3976, N3743);
  not NOT1_787 (N3977, N3744);
  not NOT1_795 (N3987, N3757);
  not NOT1_796 (N3988, N3763);
  not NOT1_797 (N3989, N3764);
  not NOT1_798 (N3990, N3765);
  not NOT1_799 (N3991, N3766);
  not NOT1_805 (N4027, N3705);
  not NOT1_838 (N4188, N3771);
  not NOT1_839 (N4191, N3775);
  not NOT1_843 (N4199, N3816);
  not NOT1_844 (N4200, N3789);
  not NOT1_845 (N4203, N3793);
  not NOT1_851 (N4223, N3810);
  not NOT1_852 (N4224, N3813);
  not NOT1_867 (N4267, N3824);
  not NOT1_872 (N4272, N4031);
  not NOT1_875 (N4275, N4036);
  not NOT1_879 (N4279, N4042);
  not NOT1_896 (N4357, N3968);
  not NOT1_897 (N4364, N3962);
  not NOT1_904 (N4405, N3921);
  not NOT1_917 (N4515, N4183);
  not NOT1_919 (N4521, N4008);
  not NOT1_920 (N4523, N4011);
  not NOT1_921 (N4524, N4198);
  not NOT1_978 (N4724, N4147);
  not NOT1_979 (N4725, N4144);
  not NOT1_980 (N4726, N4159);
  not NOT1_981 (N4727, N4156);
  not NOT1_982 (N4728, N4153);
  not NOT1_983 (N4729, N4097);
  not NOT1_984 (N4730, N4094);
  not NOT1_985 (N4731, N4091);
  not NOT1_986 (N4732, N4088);
  not NOT1_987 (N4733, N4109);
  not NOT1_988 (N4734, N4106);
  not NOT1_989 (N4735, N4103);
  not NOT1_990 (N4736, N4100);
  not NOT1_996 (N4855, N3732);
  not NOT1_1012 (N4965, N4225);
  not NOT1_1013 (N4966, N4228);
  not NOT1_1014 (N4967, N4231);
  not NOT1_1015 (N4968, N4234);
  not NOT1_1016 (N4972, N4246);
  not NOT1_1017 (N4973, N4249);
  not NOT1_1018 (N4974, N4252);
  not NOT1_1020 (N4976, N3797);
  not NOT1_1033 (N5052, N4237);
  not NOT1_1034 (N5053, N4240);
  not NOT1_1035 (N5054, N4243);
  not NOT1_1039 (N5058, N4264);
  not NOT1_1049 (N5069, N3893);
  not NOT1_1051 (N5071, N3887);
  not NOT1_1053 (N5073, N3881);
  not NOT1_1055 (N5075, N3873);
  not NOT1_1057 (N5077, N3867);
  not NOT1_1059 (N5079, N3861);
  not NOT1_1061 (N5081, N3855);
  not NOT1_1063 (N5083, N3849);
  not NOT1_1065 (N5085, N3842);
  not NOT1_1067 (N5087, N4575);
  not NOT1_1086 (N5106, N3956);
  not NOT1_1088 (N5108, N3948);
  not NOT1_1090 (N5110, N3942);
  not NOT1_1093 (N5113, N3933);
  not NOT1_1095 (N5115, N3927);
  not NOT1_1100 (N5120, N4627);
  not NOT1_1144 (N5176, N4608);
  not NOT1_1176 (N5241, N4939);
  not NOT1_1216 (N5312, N5049);
  not NOT1_1247 (N5469, N4290);
  not NOT1_1268 (N5622, N4385);
  not NOT1_1284 (N5728, N4310);
  not NOT1_1295 (N5755, N5236);
  not NOT1_1299 (N5956, N5346);
  not NOT1_1302 (N6023, N5371);
  not NOT1_1304 (N6025, N5315);
  not NOT1_1305 (N6028, N5324);
  not NOT1_1310 (N6044, N5385);
  not NOT1_1317 (N6067, N5377);
  not NOT1_1318 (N6068, N5382);
  not NOT1_1328 (N6079, N5418);
  not NOT1_1380 (N6139, N5573);
  not NOT1_1425 (N6197, N5692);
  not NOT1_1426 (N6200, N5696);
  not NOT1_1427 (N6203, N5703);
  not NOT1_1428 (N6206, N5707);
  not NOT1_1434 (N6234, N5756);
  not NOT1_1480 (N6373, N5736);
  not NOT1_1481 (N6374, N5739);
  not NOT1_1482 (N6375, N5742);
  not NOT1_1483 (N6376, N5745);
  not NOT1_1495 (N6434, N5264);
  not NOT1_1502 (N6469, N5319);
  not NOT1_1504 (N6471, N5328);
  not NOT1_1551 (N6651, N5462);
  not NOT1_1552 (N6653, N5389);
  not NOT1_1554 (N6657, N5396);
  not NOT1_1557 (N6661, N5407);
  not NOT1_1561 (N6666, N5424);
  not NOT1_1562 (N6668, N5431);
  not NOT1_1563 (N6670, N5441);
  not NOT1_1564 (N6672, N5452);
  not NOT1_1565 (N6675, N6117);
  not NOT1_1571 (N6690, N5562);
  not NOT1_1575 (N6695, N5579);
  not NOT1_1576 (N6698, N5595);
  not NOT1_1578 (N6700, N5606);
  not NOT1_1579 (N6703, N6175);
  not NOT1_1580 (N6708, N5700);
  not NOT1_1582 (N6710, N5711);
  not NOT1_1627 (N6807, N6482);
  not NOT1_1629 (N6809, N6486);
  not NOT1_1631 (N6811, N6490);
  not NOT1_1633 (N6411, N6494);
  not NOT1_1638 (N6823, N6500);
  not NOT1_1640 (N6825, N6504);
  not NOT1_1642 (N6827, N6508);
  not NOT1_1644 (N6829, N6512);
  not NOT1_1646 (N6831, N6397);
  not NOT1_1647 (N6834, N6566);
  not NOT1_1649 (N6836, N6569);
  not NOT1_1651 (N6838, N6572);
  not NOT1_1653 (N6437, N6575);
  not NOT1_1658 (N6850, N6580);
  not NOT1_1660 (N6852, N6584);
  not NOT1_1662 (N6854, N6587);
  not NOT1_1665 (N6857, N6427);
  not NOT1_1675 (N6876, N6637);
  not NOT1_1683 (N6889, N6536);
  not NOT1_1686 (N6894, N6539);
  not NOT1_1687 (N6895, N6553);
  not NOT1_1689 (N6897, N6419);
  not NOT1_1690 (N6900, N6556);
  not NOT1_1696 (N6912, N6606);
  not NOT1_1697 (N6913, N6609);
  not NOT1_1698 (N6914, N6619);
  not NOT1_1700 (N6916, N6445);
  not NOT1_1701 (N6919, N6622);
  not NOT1_1702 (N6922, N6634);
  not NOT1_1734 (N6977, N6792);
  not NOT1_1735 (N6978, N6795);
  not NOT1_1746 (N7015, N6866);
  not NOT1_1752 (N7022, N6939);
  not NOT1_1753 (N7023, N6817);
  not NOT1_1764 (N7048, N6957);
  not NOT1_1765 (N7049, N6844);
  not NOT1_1771 (N7072, N6881);
  not NOT1_1776 (N7079, N6891);
  not NOT1_1779 (N7084, N6901);
  not NOT1_1783 (N7088, N6909);
  not NOT1_1793 (N7115, N7019);
  not NOT1_1794 (N7116, N7021);
  not NOT1_1798 (N7130, N7045);
  not NOT1_1799 (N7131, N7047);
  not NOT1_1805 (N7149, N7003);
  not NOT1_1806 (N7150, N7006);
  not NOT1_1824 (N7177, N7041);
  not NOT1_1829 (N7182, N7065);
  not NOT1_1830 (N7183, N7094);
  not NOT1_1832 (N7185, N7097);
  not NOT1_1842 (N7205, N7101);
  not NOT1_1848 (N7215, N7076);
  not NOT1_1850 (N7217, N7080);
  not NOT1_1855 (N7228, N7090);
  not NOT1_1886 (N7363, N7198);
  not NOT1_1888 (N7365, N7190);
  not NOT1_1892 (N7405, N7209);
  not NOT1_1894 (N7407, N7212);
  not NOT1_1898 (N7415, N7219);
  not NOT1_1900 (N7417, N7222);
  not NOT1_1902 (N7419, N7225);
  not NOT1_1912 (N7432, N7250);
  not NOT1_1946 (N7465, N7310);
  not NOT1_1947 (N7466, N7294);
  not NOT1_1948 (N7467, N7288);
  not NOT1_1949 (N7468, N7301);
  not NOT1_1951 (N7470, N7304);
  not NOT1_1952 (N7471, N7282);
  not NOT1_1953 (N7472, N7276);
  not NOT1_1954 (N7473, N7270);
  not NOT1_1996 (N7529, N7402);
  not NOT1_2008 (N7585, N7409);
  not NOT1_2010 (N7587, N7412);
  not NOT1_2015 (N7598, N7421);
  not NOT1_2066 (N7699, N7573);
  not NOT1_2067 (N7700, N7567);
  not NOT1_2068 (N7701, N7561);
  not NOT1_2069 (N7702, N7555);
  not NOT1_2071 (N7704, N7549);
  not NOT1_2072 (N7705, N7543);
  not NOT1_2073 (N7706, N7537);
  not NOT1_2074 (N7707, N7531);
  not NOT1_2075 (N7708, N7579);
  not NOT1_2077 (N7710, N7582);
  not NOT1_2081 (N7718, N7589);
  not NOT1_2083 (N7720, N7592);
  not NOT1_2085 (N7722, N7595);
  not NOT1_2119 (N7768, N7712);
  not NOT1_2121 (N7770, N7715);
  not NOT1_2126 (N7781, N7724);
  not NOT1_2131 (N7796, N7762);
  not NOT1_2133 (N7798, N7765);
  not NOT1_2137 (N7806, N7772);
  not NOT1_2139 (N7808, N7775);
  not NOT1_2141 (N7810, N7778);
  not NOT1_2151 (N7832, N7800);
  not NOT1_2153 (N7834, N7803);
  not NOT1_2158 (N7845, N7812);
  not NOT1_2163 (N7860, N7826);
  not NOT1_2165 (N7862, N7829);
  not NOT1_2169 (N7870, N7836);
  not NOT1_2171 (N7872, N7839);
  not NOT1_2173 (N7874, N7842);
  not NOT1_2183 (N7896, N7864);
  not NOT1_2185 (N7898, N7867);
  not NOT1_2190 (N7909, N7876);
  not NOT1_2195 (N7924, N7890);
  not NOT1_2197 (N7926, N7893);
  not NOT1_2199 (N7928, N7900);
  not NOT1_2201 (N7930, N7903);
  not NOT1_2205 (N7938, N7906);
  not NOT1_2217 (N7966, N7932);
  not NOT1_2219 (N7968, N7935);
  not NOT1_2222 (N7973, N7940);
  not NOT1_2231 (N7992, N7970);
  not NOT1_2243 (N8020, N7998);
  not NOT1_2245 (N8022, N8001);
  not NOT1_2248 (N8026, N8004);
  not NOT1_2252 (N8033, N8013);
  not NOT1_2255 (N8036, N8017);
  not NOT1_2259 (N8040, N8038);
  not NOT1_2261 (N8042, N8039);
  not NOT1_2267 (N8056, N8045);
  not NOT1_2269 (N8058, N8048);
  not NOT1_2276 (N8073, N8061);
  not NOT1_2277 (N8074, N8064);
  not NOT1_2306 (N8127, N8125);
  not NOT1_2307 (N8128, N8126);
  or OR2_199 (N2350, N1067, N514);
  or OR2_413 (N2984, N242, N514);
  or OR2_623 (N3664, N2831, N3401);
  or OR2_624 (N3665, N2832, N3402);
  or OR2_625 (N3666, N2833, N3403);
  or OR2_626 (N3667, N2834, N3404);
  or OR2_631 (N3672, N2847, N3409);
  or OR2_632 (N3673, N2848, N3410);
  or OR2_633 (N3674, N2849, N3411);
  or OR2_634 (N3675, N2850, N3412);
  or OR2_650 (N3700, N2907, N3444);
  or OR2_651 (N3701, N2908, N3445);
  or OR2_652 (N3702, N2909, N3446);
  or OR2_655 (N3705, N2910, N3447);
  or OR2_656 (N3708, N2919, N3450);
  or OR2_657 (N3709, N2921, N3451);
  or OR2_658 (N3710, N2922, N3452);
  or OR2_662 (N3715, N2934, N3459);
  or OR2_663 (N3716, N2935, N3460);
  or OR2_664 (N3717, N2936, N3461);
  or OR2_665 (N3718, N2937, N3462);
  or OR2_679 (N3732, N2942, N2958);
  or OR2_684 (N3742, N2979, N3481);
  or OR2_685 (N3743, N2981, N3483);
  or OR2_686 (N3744, N2982, N3484);
  or OR2_699 (N3757, N3013, N3502);
  or OR2_705 (N3763, N3023, N3504);
  or OR2_706 (N3764, N3024, N3505);
  or OR2_707 (N3765, N3025, N3506);
  or OR2_708 (N3766, N3026, N3507);
  or OR2_746 (N3828, N3739, N2970);
  or OR2_747 (N3829, N3740, N2971);
  or OR2_749 (N3831, N3738, N2969);
  or OR2_758 (N3842, N3681, N2868);
  or OR2_759 (N3849, N3682, N2869);
  or OR2_760 (N3855, N3683, N2870);
  or OR2_761 (N3861, N3684, N2871);
  or OR2_762 (N3867, N3685, N2872);
  or OR2_763 (N3873, N3686, N2873);
  or OR2_764 (N3881, N3687, N2874);
  or OR2_765 (N3887, N3688, N2875);
  or OR2_766 (N3893, N3689, N2876);
  or OR2_777 (N3921, N3724, N2955);
  or OR2_778 (N3927, N3725, N2956);
  or OR2_779 (N3933, N3726, N2957);
  or OR2_780 (N3942, N3727, N2959);
  or OR2_781 (N3948, N3728, N2960);
  or OR2_782 (N3956, N3729, N2961);
  or OR2_783 (N3962, N3730, N2962);
  or OR2_784 (N3968, N3731, N2963);
  or OR2_801 (N4008, N3723, N2954);
  or OR2_802 (N4011, N3680, N2867);
  or OR2_834 (N4183, N3758, N3980);
  or OR2_1223 (N5346, N3921, N5119);
  or OR2_1493 (N6419, N4305, N6105);
  or OR2_1498 (N6445, N4400, N6162);
  or OR2_1519 (N6512, N4310, N6107);
  or OR2_1637 (N6817, N6397, N6664);
  or OR2_1657 (N6844, N6427, N6693);
  or OR2_1679 (N6881, N6411, N6089);
  or OR2_1685 (N6891, N6419, N6138);
  or OR2_1691 (N6901, N6437, N6147);
  or OR2_1695 (N6909, N6445, N6194);
  or OR2_1704 (N6924, N6382, N6801);
  or OR2_1705 (N6925, N6386, N6802);
  or OR2_1736 (N6979, N6879, N6880);
  or OR2_1857 (N7236, N7173, N7125);
  or OR2_1858 (N7239, N7174, N7126);
  or OR2_1859 (N7242, N7175, N7127);
  or OR2_1860 (N7245, N7176, N7040);
  or OR2_1861 (N7250, N7178, N7139);
  or OR2_1862 (N7257, N7179, N7140);
  or OR2_1863 (N7260, N7180, N7141);
  or OR2_1864 (N7263, N7181, N7064);
  or OR2_2065 (N7698, N7624, N7625);
  or OR2_2264 (N8045, N8043, N8041);
  or OR2_2265 (N8048, N8044, N8035);
  or OR2_2282 (N8079, N7530, N8077);
  or OR2_2283 (N8082, N7479, N8078);
  or OR2_2288 (N8093, N8089, N3071);
  or OR2_2289 (N8096, N8090, N3072);
  or OR3_627 (N3668, N2835, N3405, N457);
  or OR3_628 (N3669, N2836, N3406, N468);
  or OR3_629 (N3670, N2837, N3407, N422);
  or OR3_630 (N3671, N2838, N3408, N435);
  or OR3_635 (N3676, N2851, N3413, N389);
  or OR3_636 (N3677, N2852, N3414, N400);
  or OR3_637 (N3678, N2853, N3415, N411);
  or OR3_638 (N3679, N2854, N3416, N374);
  or OR3_653 (N3703, N2911, N3448, N479);
  or OR3_654 (N3704, N2912, N3449, N490);
  or OR3_659 (N3711, N2923, N3453, N503);
  or OR3_660 (N3712, N2924, N3454, N523);
  or OR3_661 (N3713, N2925, N3455, N534);
  or OR3_666 (N3719, N2938, N3463, N389);
  or OR3_667 (N3720, N2939, N3464, N400);
  or OR3_668 (N3721, N2940, N3465, N411);
  or OR3_669 (N3722, N2941, N3466, N374);
  or OR3_687 (N3745, N2983, N3485, N503);
  or OR3_688 (N3746, N2985, N3486, N523);
  or OR3_689 (N3747, N2986, N3487, N534);
  or OR3_709 (N3767, N3027, N3508, N457);
  or OR3_710 (N3768, N3028, N3509, N468);
  or OR3_711 (N3769, N3029, N3510, N422);
  or OR3_712 (N3770, N3030, N3511, N435);
  or OR3_836 (N4185, N3761, N3982, N446);
  or OR3_1514 (N6490, N4284, N6088, N6089);
  or OR3_1518 (N6508, N4305, N6105, N6106);
  or OR3_1528 (N6572, N4379, N6146, N6147);
  or OR3_1532 (N6587, N4400, N6162, N6163);
  or OR3_1670 (N6866, N4197, N6718, N3785);
  or OR3_1837 (N7190, N4956, N7146, N3781);
  or OR3_1840 (N7198, N4960, N7147, N3786);
  or OR3_1867 (N7270, N4957, N7187, N3782);
  or OR3_1868 (N7276, N4958, N7188, N3783);
  or OR3_1869 (N7282, N4959, N7189, N3784);
  or OR3_1870 (N7288, N4961, N7196, N3787);
  or OR3_1871 (N7294, N3998, N7197, N3788);
  or OR3_1874 (N7304, N4980, N7207, N3800);
  or OR3_1875 (N7310, N4984, N7208, N3805);
  or OR3_1998 (N7531, N4981, N7481, N3801);
  or OR3_1999 (N7537, N4982, N7482, N3802);
  or OR3_2000 (N7543, N4983, N7483, N3803);
  or OR3_2001 (N7549, N5165, N7484, N3804);
  or OR3_2002 (N7555, N4985, N7485, N3806);
  or OR3_2003 (N7561, N4986, N7486, N3807);
  or OR3_2004 (N7567, N4547, N7487, N3808);
  or OR3_2005 (N7573, N4987, N7488, N3809);
  or OR4_873 (N4273, N4032, N4033, N3614, N3615);
  or OR4_874 (N4274, N4034, N4035, N3614, N3615);
  or OR4_876 (N4276, N4037, N4038, N3614, N3615);
  or OR4_877 (N4277, N4039, N4040, N3614, N3615);
  or OR4_1486 (N6382, N4268, N6071, N6072, N6073);
  or OR4_1487 (N6386, N3968, N5065, N5066, N6074);
  or OR4_1512 (N6482, N4280, N6083, N6084, N6085);
  or OR4_1517 (N6504, N4301, N6102, N6103, N6104);
  or OR4_1522 (N6536, N4301, N6102, N6103, N6133);
  or OR4_1526 (N6566, N3962, N5117, N6143, N6144);
  or OR4_1531 (N6584, N4396, N6159, N6160, N6161);
  or OR4_1535 (N6606, N4396, N6159, N6160, N6189);
  or OR4_1916 (N7435, N7011, N7338, N3621, N2591);
  or OR4_1924 (N7443, N7012, N7340, N3632, N2600);
  or OR4_1930 (N7449, N7013, N7342, N3641, N2605);
  or OR4_1950 (N7469, N7016, N7364, N3660, N2626);
  or OR4_1974 (N7505, N7433, N7434, N3616, N2585);
  or OR4_1976 (N7507, N7339, N7436, N3622, N2592);
  or OR4_1977 (N7508, N7437, N7438, N3623, N2593);
  or OR4_1978 (N7509, N7439, N7440, N3624, N2594);
  or OR4_1979 (N7510, N7441, N7442, N3627, N2595);
  or OR4_1981 (N7512, N7341, N7444, N3633, N2601);
  or OR4_1982 (N7513, N7445, N7446, N3634, N2602);
  or OR4_1983 (N7514, N7447, N7448, N3635, N2603);
  or OR4_1984 (N7515, N7450, N7451, N3646, N2610);
  or OR4_1985 (N7516, N7452, N7453, N3647, N2611);
  or OR4_1986 (N7517, N7454, N7455, N3648, N2612);
  or OR4_1987 (N7518, N7349, N7456, N3649, N2613);
  or OR4_1988 (N7519, N7457, N7458, N3654, N2618);
  or OR4_1989 (N7520, N7459, N7460, N3655, N2619);
  or OR4_1990 (N7521, N7461, N7462, N3656, N2620);
  or OR4_1991 (N7522, N7357, N7463, N3657, N2621);
  or OR4_1992 (N7525, N4741, N7114, N2624, N7464);
  or OR4_2088 (N7727, N7666, N7667, N3617, N2586);
  or OR4_2089 (N7728, N7668, N7669, N3618, N2587);
  or OR4_2090 (N7729, N7670, N7671, N3619, N2588);
  or OR4_2091 (N7730, N7672, N7673, N3620, N2589);
  or OR4_2092 (N7731, N7674, N7675, N3628, N2596);
  or OR4_2093 (N7732, N7676, N7677, N3629, N2597);
  or OR4_2094 (N7733, N7678, N7679, N3630, N2598);
  or OR4_2095 (N7734, N7680, N7681, N3631, N2599);
  or OR4_2096 (N7735, N7682, N7683, N3638, N2604);
  or OR4_2097 (N7736, N7684, N7685, N3642, N2606);
  or OR4_2098 (N7737, N7686, N7687, N3643, N2607);
  or OR4_2099 (N7738, N7688, N7689, N3644, N2608);
  or OR4_2100 (N7739, N7690, N7691, N3645, N2609);
  or OR4_2101 (N7740, N7692, N7693, N3651, N2615);
  or OR4_2102 (N7741, N7694, N7695, N3652, N2616);
  or OR4_2103 (N7742, N7696, N7697, N3653, N2617);
  or OR4_2241 (N8013, N7988, N7989, N7990, N7991);
  or OR4_2242 (N8017, N7994, N7995, N7996, N7997);
  or OR4_2278 (N8075, N7526, N8071, N3659, N2625);
  or OR4_2279 (N8076, N7636, N8072, N3661, N2625);
  or OR4_2300 (N8121, N8117, N8118, N3662, N2703);
  or OR4_2301 (N8122, N8119, N8120, N3663, N2778);
  or OR4_2302 (N8123, N8113, N8114, N3650, N2614);
  or OR4_2303 (N8124, N8115, N8116, N3658, N2622);
  and g2 (N6117, N5441, N5431, N5424, N6138);
  and g3 (n_303, N5264, N4405);
  and g4 (N6149, N5595, N5579, N5606, n_303);
  and g6 (N6175, N5595, N5264, N5579, N6194);
  and g7 (n_305, N5431, N5462);
  and g8 (N6091, N5441, N5424, N5452, n_305);
  or g9 (n_306, N4297, N6094);
  or g10 (N6397, N6095, N6096, N6097, n_306);
  and g11 (n_307, N5452, N5441);
  and g12 (N6097, N5424, N4310, N5431, n_307);
  or g13 (n_308, N4392, N6152);
  or g14 (N6427, N6153, N6154, N6155, n_308);
  and g15 (n_309, N5606, N5595);
  and g16 (N6155, N5579, N3921, N5264, n_309);
  or g25 (n_314, N4067, N5954);
  or g26 (N6580, N6156, N6157, N6158, n_314);
  and g28 (N6158, N5595, N5606, N5264, N5119);
  or g29 (n_316, N4298, N6098);
  or g30 (N6500, N6099, N6100, N6101, n_316);
  and g32 (N6101, N5441, N5452, N5431, N6107);
  nor g33 (n_318, N6932, N7037, N7034);
  nor g34 (n_319, N7031, N7028);
  nor g35 (n_320, N7245, N7242);
  nor g36 (n_321, N7239, N7236);
  and g37 (N7503, n_318, n_319, n_320, n_321);
  nor g38 (n_323, N6164, N6967, N7060);
  nor g39 (n_324, N7057, N7054);
  nor g40 (n_325, N7263, N7260);
  and g41 (n_326, n_322, N7432);
  not g42 (n_322, N7257);
  and g43 (N7504, n_323, n_324, n_325, n_326);
  nor g44 (n_328, N7474, N7476, N6716);
  and g45 (n_329, n_327, N386, N559);
  not g46 (n_327, N6877);
  and g47 (n_330, N556, N552);
  and g48 (n_331, N562, N245);
  and g49 (N7703, n_328, n_329, n_330, n_331);
  or g51 (N6609, N6156, N6157, N6184, n_314);
  or g53 (N6539, N6099, N6100, N6127, n_316);
  not g54 (N5365, N5065);
endmodule

