
module memctrl(pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006,
     pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014,
     pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022,
     pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030,
     pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038,
     pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046,
     pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054,
     pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
     pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
     pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078,
     pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086,
     pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094,
     pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102,
     pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110,
     pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118,
     pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126,
     pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
     pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
     pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150,
     pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158,
     pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166,
     pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174,
     pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182,
     pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190,
     pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198,
     pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
     pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
     pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222,
     pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230,
     pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238,
     pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246,
     pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254,
     pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262,
     pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270,
     pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
     pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
     pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294,
     pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302,
     pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310,
     pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318,
     pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326,
     pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334,
     pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342,
     pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
     pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
     pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366,
     pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374,
     pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382,
     pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390,
     pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398,
     pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406,
     pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414,
     pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
     pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
     pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438,
     pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446,
     pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454,
     pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462,
     pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470,
     pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478,
     pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486,
     pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
     pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
     pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510,
     pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518,
     pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526,
     pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534,
     pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542,
     pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550,
     pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558,
     pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
     pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
     pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582,
     pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590,
     pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598,
     pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606,
     pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614,
     pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622,
     pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630,
     pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
     pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
     pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654,
     pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662,
     pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670,
     pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678,
     pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686,
     pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694,
     pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702,
     pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
     pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
     pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726,
     pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734,
     pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742,
     pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750,
     pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758,
     pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766,
     pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774,
     pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
     pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
     pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798,
     pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806,
     pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814,
     pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822,
     pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830,
     pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838,
     pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846,
     pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
     pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
     pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870,
     pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878,
     pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886,
     pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894,
     pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902,
     pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910,
     pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918,
     pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
     pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
     pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942,
     pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950,
     pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958,
     pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966,
     pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974,
     pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982,
     pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990,
     pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
     pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
     pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014,
     pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022,
     pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030,
     pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038,
     pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046,
     pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054,
     pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062,
     pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
     pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
     pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086,
     pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094,
     pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102,
     pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110,
     pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118,
     pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126,
     pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134,
     pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
     pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
     pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158,
     pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166,
     pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174,
     pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182,
     pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190,
     pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198,
     pi1199, pi1200, pi1201, pi1202, pi1203, po0000, po0001, po0002,
     po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010,
     po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018,
     po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
     po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
     po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042,
     po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050,
     po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058,
     po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066,
     po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074,
     po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082,
     po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090,
     po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
     po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
     po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114,
     po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122,
     po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130,
     po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138,
     po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146,
     po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154,
     po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162,
     po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
     po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
     po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186,
     po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194,
     po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202,
     po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210,
     po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218,
     po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226,
     po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234,
     po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
     po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
     po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258,
     po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266,
     po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274,
     po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282,
     po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290,
     po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298,
     po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306,
     po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
     po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
     po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330,
     po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338,
     po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346,
     po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354,
     po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362,
     po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370,
     po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378,
     po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
     po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
     po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402,
     po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410,
     po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418,
     po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426,
     po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434,
     po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442,
     po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450,
     po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
     po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
     po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474,
     po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482,
     po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490,
     po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498,
     po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506,
     po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514,
     po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522,
     po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
     po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
     po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546,
     po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554,
     po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562,
     po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570,
     po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578,
     po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586,
     po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594,
     po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
     po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
     po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618,
     po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626,
     po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634,
     po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642,
     po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650,
     po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658,
     po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666,
     po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
     po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
     po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690,
     po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698,
     po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706,
     po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714,
     po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722,
     po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730,
     po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738,
     po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
     po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
     po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762,
     po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770,
     po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778,
     po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786,
     po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794,
     po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802,
     po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810,
     po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
     po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
     po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834,
     po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842,
     po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850,
     po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858,
     po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866,
     po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874,
     po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882,
     po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
     po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
     po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906,
     po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914,
     po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922,
     po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930,
     po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938,
     po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946,
     po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954,
     po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
     po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
     po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978,
     po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986,
     po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994,
     po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002,
     po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010,
     po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018,
     po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026,
     po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
     po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
     po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050,
     po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058,
     po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066,
     po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074,
     po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082,
     po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090,
     po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098,
     po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
     po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
     po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122,
     po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130,
     po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138,
     po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146,
     po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154,
     po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162,
     po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170,
     po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
     po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
     po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194,
     po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202,
     po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210,
     po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218,
     po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226,
     po1227, po1228, po1229, po1230);
  input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
       pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015,
       pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023,
       pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031,
       pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039,
       pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047,
       pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055,
       pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063,
       pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
       pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
       pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087,
       pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095,
       pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103,
       pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111,
       pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119,
       pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127,
       pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135,
       pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
       pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
       pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159,
       pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167,
       pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175,
       pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183,
       pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191,
       pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199,
       pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207,
       pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
       pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
       pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231,
       pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239,
       pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247,
       pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255,
       pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263,
       pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271,
       pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279,
       pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
       pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
       pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303,
       pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311,
       pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319,
       pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327,
       pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335,
       pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343,
       pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351,
       pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
       pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
       pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375,
       pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383,
       pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391,
       pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399,
       pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407,
       pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415,
       pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423,
       pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
       pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
       pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447,
       pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455,
       pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463,
       pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471,
       pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479,
       pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487,
       pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495,
       pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
       pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
       pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519,
       pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527,
       pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535,
       pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543,
       pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551,
       pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559,
       pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567,
       pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
       pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
       pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591,
       pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599,
       pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607,
       pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615,
       pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623,
       pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631,
       pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639,
       pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
       pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
       pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663,
       pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671,
       pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679,
       pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687,
       pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695,
       pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703,
       pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711,
       pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
       pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
       pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735,
       pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743,
       pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751,
       pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759,
       pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767,
       pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775,
       pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783,
       pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
       pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
       pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807,
       pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815,
       pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823,
       pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831,
       pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839,
       pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847,
       pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855,
       pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
       pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
       pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879,
       pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887,
       pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895,
       pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903,
       pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911,
       pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919,
       pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927,
       pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
       pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
       pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951,
       pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959,
       pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967,
       pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975,
       pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983,
       pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991,
       pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999,
       pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
       pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
       pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023,
       pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031,
       pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039,
       pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047,
       pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055,
       pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063,
       pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071,
       pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
       pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
       pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095,
       pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103,
       pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111,
       pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119,
       pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127,
       pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135,
       pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143,
       pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
       pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
       pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167,
       pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175,
       pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183,
       pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191,
       pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199,
       pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006,
       po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014,
       po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022,
       po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030,
       po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038,
       po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046,
       po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054,
       po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
       po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
       po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078,
       po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086,
       po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094,
       po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102,
       po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110,
       po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118,
       po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126,
       po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
       po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
       po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150,
       po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158,
       po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166,
       po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174,
       po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182,
       po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190,
       po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198,
       po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
       po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
       po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222,
       po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230,
       po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238,
       po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246,
       po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254,
       po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262,
       po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270,
       po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
       po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
       po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294,
       po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302,
       po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310,
       po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318,
       po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326,
       po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334,
       po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342,
       po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
       po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
       po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366,
       po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374,
       po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382,
       po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390,
       po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398,
       po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406,
       po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414,
       po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
       po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
       po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438,
       po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446,
       po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454,
       po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462,
       po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470,
       po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478,
       po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486,
       po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
       po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
       po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510,
       po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518,
       po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526,
       po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534,
       po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542,
       po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550,
       po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558,
       po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
       po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
       po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582,
       po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590,
       po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598,
       po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606,
       po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614,
       po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622,
       po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630,
       po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
       po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
       po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654,
       po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662,
       po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670,
       po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678,
       po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686,
       po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694,
       po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702,
       po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
       po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
       po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726,
       po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734,
       po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742,
       po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750,
       po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758,
       po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766,
       po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774,
       po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
       po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
       po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798,
       po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806,
       po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814,
       po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822,
       po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830,
       po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838,
       po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846,
       po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
       po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
       po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870,
       po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878,
       po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886,
       po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894,
       po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902,
       po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910,
       po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918,
       po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
       po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
       po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942,
       po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950,
       po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958,
       po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966,
       po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974,
       po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982,
       po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990,
       po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
       po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
       po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014,
       po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022,
       po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030,
       po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038,
       po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046,
       po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054,
       po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062,
       po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
       po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
       po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086,
       po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094,
       po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102,
       po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110,
       po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118,
       po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126,
       po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134,
       po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
       po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
       po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158,
       po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166,
       po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174,
       po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182,
       po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190,
       po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198,
       po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206,
       po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
       po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
       po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
       pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015,
       pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023,
       pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031,
       pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039,
       pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047,
       pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055,
       pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063,
       pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
       pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
       pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087,
       pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095,
       pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103,
       pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111,
       pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119,
       pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127,
       pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135,
       pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
       pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
       pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159,
       pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167,
       pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175,
       pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183,
       pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191,
       pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199,
       pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207,
       pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
       pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
       pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231,
       pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239,
       pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247,
       pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255,
       pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263,
       pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271,
       pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279,
       pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
       pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
       pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303,
       pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311,
       pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319,
       pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327,
       pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335,
       pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343,
       pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351,
       pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
       pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
       pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375,
       pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383,
       pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391,
       pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399,
       pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407,
       pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415,
       pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423,
       pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
       pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
       pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447,
       pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455,
       pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463,
       pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471,
       pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479,
       pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487,
       pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495,
       pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
       pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
       pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519,
       pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527,
       pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535,
       pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543,
       pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551,
       pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559,
       pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567,
       pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
       pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
       pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591,
       pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599,
       pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607,
       pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615,
       pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623,
       pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631,
       pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639,
       pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
       pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
       pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663,
       pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671,
       pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679,
       pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687,
       pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695,
       pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703,
       pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711,
       pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
       pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
       pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735,
       pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743,
       pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751,
       pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759,
       pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767,
       pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775,
       pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783,
       pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
       pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
       pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807,
       pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815,
       pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823,
       pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831,
       pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839,
       pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847,
       pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855,
       pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
       pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
       pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879,
       pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887,
       pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895,
       pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903,
       pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911,
       pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919,
       pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927,
       pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
       pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
       pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951,
       pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959,
       pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967,
       pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975,
       pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983,
       pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991,
       pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999,
       pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
       pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
       pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023,
       pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031,
       pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039,
       pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047,
       pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055,
       pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063,
       pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071,
       pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
       pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
       pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095,
       pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103,
       pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111,
       pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119,
       pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127,
       pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135,
       pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143,
       pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
       pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
       pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167,
       pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175,
       pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183,
       pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191,
       pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199,
       pi1200, pi1201, pi1202, pi1203;
  wire po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
       po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015,
       po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023,
       po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031,
       po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039,
       po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047,
       po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055,
       po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063,
       po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
       po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
       po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087,
       po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095,
       po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103,
       po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111,
       po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119,
       po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127,
       po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135,
       po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
       po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
       po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159,
       po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167,
       po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175,
       po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183,
       po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191,
       po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199,
       po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207,
       po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
       po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
       po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231,
       po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239,
       po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247,
       po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255,
       po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263,
       po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271,
       po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279,
       po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
       po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
       po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303,
       po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311,
       po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319,
       po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327,
       po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335,
       po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343,
       po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351,
       po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
       po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
       po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375,
       po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383,
       po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391,
       po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399,
       po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407,
       po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415,
       po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423,
       po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
       po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
       po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447,
       po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455,
       po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463,
       po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471,
       po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479,
       po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487,
       po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495,
       po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
       po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
       po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519,
       po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527,
       po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535,
       po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543,
       po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551,
       po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559,
       po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567,
       po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
       po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
       po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591,
       po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599,
       po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607,
       po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615,
       po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623,
       po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631,
       po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639,
       po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
       po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
       po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663,
       po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671,
       po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679,
       po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687,
       po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695,
       po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703,
       po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711,
       po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
       po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
       po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735,
       po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743,
       po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751,
       po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759,
       po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767,
       po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775,
       po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783,
       po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
       po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
       po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807,
       po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815,
       po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823,
       po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831,
       po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839,
       po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847,
       po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855,
       po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
       po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
       po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879,
       po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887,
       po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895,
       po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903,
       po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911,
       po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919,
       po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927,
       po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
       po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
       po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951,
       po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959,
       po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967,
       po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975,
       po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983,
       po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991,
       po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999,
       po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
       po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
       po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023,
       po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031,
       po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039,
       po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047,
       po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055,
       po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063,
       po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071,
       po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
       po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
       po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095,
       po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103,
       po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111,
       po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119,
       po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127,
       po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135,
       po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143,
       po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
       po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
       po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167,
       po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175,
       po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183,
       po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191,
       po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199,
       po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207,
       po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215,
       po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
       po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444;
  wire n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452;
  wire n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460;
  wire n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468;
  wire n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476;
  wire n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484;
  wire n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492;
  wire n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500;
  wire n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508;
  wire n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516;
  wire n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524;
  wire n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532;
  wire n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540;
  wire n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548;
  wire n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556;
  wire n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564;
  wire n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572;
  wire n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580;
  wire n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588;
  wire n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596;
  wire n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604;
  wire n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612;
  wire n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620;
  wire n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628;
  wire n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636;
  wire n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644;
  wire n2645, n2646, n2647, n2648, n2649, n2652, n2653, n2654;
  wire n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662;
  wire n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670;
  wire n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678;
  wire n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686;
  wire n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694;
  wire n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702;
  wire n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710;
  wire n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718;
  wire n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726;
  wire n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734;
  wire n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742;
  wire n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
  wire n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758;
  wire n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766;
  wire n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774;
  wire n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782;
  wire n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790;
  wire n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798;
  wire n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806;
  wire n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814;
  wire n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822;
  wire n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830;
  wire n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838;
  wire n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846;
  wire n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854;
  wire n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862;
  wire n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870;
  wire n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878;
  wire n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886;
  wire n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894;
  wire n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902;
  wire n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910;
  wire n2911, n2912, n2913, n2914, n2915, n2916, n2920, n2921;
  wire n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929;
  wire n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937;
  wire n2938, n2939, n2942, n2943, n2944, n2945, n2946, n2947;
  wire n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955;
  wire n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963;
  wire n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971;
  wire n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979;
  wire n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987;
  wire n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995;
  wire n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003;
  wire n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011;
  wire n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019;
  wire n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027;
  wire n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035;
  wire n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043;
  wire n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051;
  wire n3052, n3053, n3054, n3055, n3059, n3060, n3061, n3062;
  wire n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070;
  wire n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078;
  wire n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086;
  wire n3087, n3088, n3089, n3092, n3093, n3094, n3095, n3096;
  wire n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104;
  wire n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112;
  wire n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120;
  wire n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128;
  wire n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136;
  wire n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144;
  wire n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152;
  wire n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160;
  wire n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168;
  wire n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176;
  wire n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184;
  wire n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192;
  wire n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200;
  wire n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208;
  wire n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216;
  wire n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224;
  wire n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232;
  wire n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240;
  wire n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248;
  wire n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256;
  wire n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264;
  wire n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272;
  wire n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280;
  wire n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288;
  wire n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296;
  wire n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304;
  wire n3305, n3306, n3307, n3309, n3310, n3311, n3312, n3313;
  wire n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321;
  wire n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329;
  wire n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337;
  wire n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345;
  wire n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353;
  wire n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361;
  wire n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369;
  wire n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377;
  wire n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385;
  wire n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393;
  wire n3394, n3398, n3399, n3400, n3401, n3402, n3403, n3404;
  wire n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412;
  wire n3413, n3414, n3415, n3416, n3417, n3418, n3421, n3422;
  wire n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430;
  wire n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438;
  wire n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446;
  wire n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454;
  wire n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462;
  wire n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470;
  wire n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478;
  wire n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486;
  wire n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494;
  wire n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502;
  wire n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510;
  wire n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518;
  wire n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526;
  wire n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534;
  wire n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3543;
  wire n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551;
  wire n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559;
  wire n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567;
  wire n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575;
  wire n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583;
  wire n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591;
  wire n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599;
  wire n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607;
  wire n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615;
  wire n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623;
  wire n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631;
  wire n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639;
  wire n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647;
  wire n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655;
  wire n3656, n3659, n3660, n3661, n3662, n3663, n3664, n3665;
  wire n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673;
  wire n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681;
  wire n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689;
  wire n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697;
  wire n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705;
  wire n3708, n3709, n3710, n3711, n3712, n3714, n3715, n3716;
  wire n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724;
  wire n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732;
  wire n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740;
  wire n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748;
  wire n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756;
  wire n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764;
  wire n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772;
  wire n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780;
  wire n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788;
  wire n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796;
  wire n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804;
  wire n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812;
  wire n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820;
  wire n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828;
  wire n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836;
  wire n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844;
  wire n3845, n3846, n3847, n3848, n3849, n3850, n3853, n3854;
  wire n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862;
  wire n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870;
  wire n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878;
  wire n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886;
  wire n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894;
  wire n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902;
  wire n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910;
  wire n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918;
  wire n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926;
  wire n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934;
  wire n3935, n3938, n3939, n3940, n3941, n3942, n3944, n3945;
  wire n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953;
  wire n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961;
  wire n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969;
  wire n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977;
  wire n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985;
  wire n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993;
  wire n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001;
  wire n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009;
  wire n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017;
  wire n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025;
  wire n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033;
  wire n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041;
  wire n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049;
  wire n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057;
  wire n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065;
  wire n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073;
  wire n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081;
  wire n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089;
  wire n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097;
  wire n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105;
  wire n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113;
  wire n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121;
  wire n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129;
  wire n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137;
  wire n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145;
  wire n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153;
  wire n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161;
  wire n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169;
  wire n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178;
  wire n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186;
  wire n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194;
  wire n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202;
  wire n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210;
  wire n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218;
  wire n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226;
  wire n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234;
  wire n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242;
  wire n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250;
  wire n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258;
  wire n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266;
  wire n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274;
  wire n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282;
  wire n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290;
  wire n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298;
  wire n4299, n4300, n4301, n4304, n4305, n4306, n4307, n4308;
  wire n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316;
  wire n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324;
  wire n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332;
  wire n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340;
  wire n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348;
  wire n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356;
  wire n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364;
  wire n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372;
  wire n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380;
  wire n4381, n4382, n4383, n4384, n4385, n4388, n4389, n4390;
  wire n4391, n4392, n4394, n4395, n4396, n4397, n4398, n4399;
  wire n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407;
  wire n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415;
  wire n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423;
  wire n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431;
  wire n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439;
  wire n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447;
  wire n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455;
  wire n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463;
  wire n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471;
  wire n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479;
  wire n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487;
  wire n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495;
  wire n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503;
  wire n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511;
  wire n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519;
  wire n4520, n4521, n4522, n4523, n4524, n4527, n4528, n4529;
  wire n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537;
  wire n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545;
  wire n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553;
  wire n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561;
  wire n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569;
  wire n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577;
  wire n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585;
  wire n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593;
  wire n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601;
  wire n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4611;
  wire n4612, n4613, n4614, n4615, n4617, n4618, n4619, n4620;
  wire n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628;
  wire n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636;
  wire n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644;
  wire n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652;
  wire n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660;
  wire n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668;
  wire n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676;
  wire n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684;
  wire n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692;
  wire n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700;
  wire n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708;
  wire n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716;
  wire n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724;
  wire n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732;
  wire n4733, n4734, n4735, n4736, n4737, n4740, n4741, n4742;
  wire n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750;
  wire n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758;
  wire n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766;
  wire n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774;
  wire n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782;
  wire n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790;
  wire n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798;
  wire n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806;
  wire n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814;
  wire n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822;
  wire n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830;
  wire n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838;
  wire n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846;
  wire n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855;
  wire n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863;
  wire n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871;
  wire n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879;
  wire n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887;
  wire n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895;
  wire n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903;
  wire n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911;
  wire n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919;
  wire n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927;
  wire n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935;
  wire n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943;
  wire n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951;
  wire n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959;
  wire n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967;
  wire n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975;
  wire n4976, n4977, n4978, n4981, n4982, n4983, n4984, n4985;
  wire n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993;
  wire n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001;
  wire n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009;
  wire n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017;
  wire n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025;
  wire n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033;
  wire n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041;
  wire n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049;
  wire n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057;
  wire n5058, n5059, n5060, n5061, n5062, n5065, n5066, n5067;
  wire n5068, n5069, n5071, n5072, n5073, n5074, n5075, n5076;
  wire n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084;
  wire n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092;
  wire n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100;
  wire n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108;
  wire n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116;
  wire n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124;
  wire n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132;
  wire n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140;
  wire n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148;
  wire n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156;
  wire n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164;
  wire n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172;
  wire n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180;
  wire n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188;
  wire n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196;
  wire n5197, n5198, n5199, n5200, n5201, n5204, n5205, n5206;
  wire n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214;
  wire n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222;
  wire n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230;
  wire n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238;
  wire n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246;
  wire n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254;
  wire n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262;
  wire n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270;
  wire n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278;
  wire n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5288;
  wire n5289, n5290, n5291, n5292, n5294, n5295, n5296, n5297;
  wire n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305;
  wire n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313;
  wire n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321;
  wire n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329;
  wire n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337;
  wire n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345;
  wire n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353;
  wire n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361;
  wire n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369;
  wire n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377;
  wire n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385;
  wire n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393;
  wire n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401;
  wire n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409;
  wire n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417;
  wire n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425;
  wire n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433;
  wire n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441;
  wire n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449;
  wire n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457;
  wire n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465;
  wire n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473;
  wire n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481;
  wire n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489;
  wire n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497;
  wire n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505;
  wire n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513;
  wire n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521;
  wire n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5530;
  wire n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538;
  wire n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546;
  wire n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554;
  wire n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562;
  wire n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570;
  wire n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578;
  wire n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586;
  wire n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594;
  wire n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602;
  wire n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610;
  wire n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618;
  wire n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626;
  wire n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634;
  wire n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642;
  wire n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650;
  wire n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658;
  wire n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666;
  wire n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674;
  wire n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682;
  wire n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690;
  wire n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698;
  wire n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706;
  wire n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714;
  wire n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722;
  wire n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730;
  wire n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738;
  wire n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746;
  wire n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754;
  wire n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762;
  wire n5763, n5765, n5766, n5767, n5768, n5769, n5770, n5771;
  wire n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779;
  wire n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787;
  wire n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795;
  wire n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803;
  wire n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811;
  wire n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819;
  wire n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827;
  wire n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835;
  wire n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843;
  wire n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851;
  wire n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859;
  wire n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867;
  wire n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875;
  wire n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883;
  wire n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891;
  wire n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899;
  wire n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907;
  wire n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915;
  wire n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923;
  wire n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931;
  wire n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939;
  wire n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947;
  wire n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955;
  wire n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963;
  wire n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971;
  wire n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979;
  wire n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987;
  wire n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995;
  wire n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003;
  wire n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011;
  wire n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019;
  wire n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027;
  wire n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035;
  wire n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043;
  wire n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051;
  wire n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059;
  wire n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067;
  wire n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075;
  wire n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083;
  wire n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091;
  wire n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099;
  wire n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107;
  wire n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115;
  wire n6116, n6117, n6118, n6120, n6121, n6122, n6123, n6124;
  wire n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132;
  wire n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140;
  wire n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148;
  wire n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156;
  wire n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164;
  wire n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172;
  wire n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180;
  wire n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188;
  wire n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6197;
  wire n6198, n6205, n6206, n6207, n6208, n6209, n6210, n6211;
  wire n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219;
  wire n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227;
  wire n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235;
  wire n6236, n6241, n6242, n6243, n6244, n6245, n6246, n6247;
  wire n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255;
  wire n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263;
  wire n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271;
  wire n6272, n6273, n6275, n6276, n6277, n6279, n6280, n6281;
  wire n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289;
  wire n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297;
  wire n6298, n6299, n6300, n6301, n6302, n6304, n6305, n6306;
  wire n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314;
  wire n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322;
  wire n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330;
  wire n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338;
  wire n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346;
  wire n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354;
  wire n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362;
  wire n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370;
  wire n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380;
  wire n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388;
  wire n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396;
  wire n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404;
  wire n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412;
  wire n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420;
  wire n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428;
  wire n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436;
  wire n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445;
  wire n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453;
  wire n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461;
  wire n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469;
  wire n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477;
  wire n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485;
  wire n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493;
  wire n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501;
  wire n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509;
  wire n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517;
  wire n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6527;
  wire n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535;
  wire n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543;
  wire n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551;
  wire n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559;
  wire n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567;
  wire n6568, n6569, n6570, n6572, n6573, n6574, n6575, n6576;
  wire n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584;
  wire n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592;
  wire n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600;
  wire n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608;
  wire n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616;
  wire n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624;
  wire n6625, n6628, n6629, n6630, n6631, n6632, n6633, n6634;
  wire n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642;
  wire n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650;
  wire n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658;
  wire n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666;
  wire n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674;
  wire n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682;
  wire n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690;
  wire n6691, n6692, n6693, n6695, n6696, n6697, n6698, n6699;
  wire n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707;
  wire n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715;
  wire n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723;
  wire n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731;
  wire n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739;
  wire n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747;
  wire n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755;
  wire n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763;
  wire n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771;
  wire n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779;
  wire n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787;
  wire n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795;
  wire n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803;
  wire n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811;
  wire n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819;
  wire n6820, n6821, n6822, n6823, n6825, n6826, n6827, n6828;
  wire n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836;
  wire n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844;
  wire n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852;
  wire n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860;
  wire n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868;
  wire n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876;
  wire n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884;
  wire n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892;
  wire n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900;
  wire n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908;
  wire n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916;
  wire n6917, n6918, n6919, n6921, n6922, n6923, n6924, n6925;
  wire n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933;
  wire n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941;
  wire n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949;
  wire n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957;
  wire n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965;
  wire n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973;
  wire n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981;
  wire n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989;
  wire n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997;
  wire n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005;
  wire n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013;
  wire n7014, n7015, n7017, n7018, n7019, n7020, n7021, n7022;
  wire n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030;
  wire n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038;
  wire n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046;
  wire n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054;
  wire n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062;
  wire n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070;
  wire n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078;
  wire n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086;
  wire n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094;
  wire n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102;
  wire n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110;
  wire n7111, n7113, n7114, n7115, n7116, n7117, n7118, n7119;
  wire n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127;
  wire n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135;
  wire n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143;
  wire n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151;
  wire n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159;
  wire n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167;
  wire n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175;
  wire n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183;
  wire n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191;
  wire n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199;
  wire n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207;
  wire n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216;
  wire n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224;
  wire n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232;
  wire n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240;
  wire n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248;
  wire n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256;
  wire n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264;
  wire n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272;
  wire n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280;
  wire n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288;
  wire n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296;
  wire n7297, n7298, n7299, n7301, n7302, n7303, n7304, n7305;
  wire n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313;
  wire n7314, n7315, n7316, n7317, n7320, n7321, n7322, n7323;
  wire n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333;
  wire n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341;
  wire n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349;
  wire n7350, n7351, n7353, n7354, n7356, n7357, n7358, n7359;
  wire n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367;
  wire n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375;
  wire n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383;
  wire n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391;
  wire n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399;
  wire n7400, n7401, n7402, n7403, n7404, n7406, n7407, n7408;
  wire n7409, n7411, n7413, n7415, n7417, n7418, n7419, n7420;
  wire n7421, n7422, n7423, n7424, n7425, n7427, n7428, n7429;
  wire n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437;
  wire n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445;
  wire n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453;
  wire n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461;
  wire n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469;
  wire n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477;
  wire n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485;
  wire n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493;
  wire n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501;
  wire n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509;
  wire n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517;
  wire n7518, n7519, n7520, n7521, n7522, n7526, n7527, n7528;
  wire n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536;
  wire n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544;
  wire n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552;
  wire n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560;
  wire n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568;
  wire n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576;
  wire n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584;
  wire n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592;
  wire n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600;
  wire n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608;
  wire n7609, n7610, n7611, n7612, n7613, n7614, n7617, n7618;
  wire n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626;
  wire n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634;
  wire n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642;
  wire n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650;
  wire n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658;
  wire n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666;
  wire n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674;
  wire n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682;
  wire n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690;
  wire n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698;
  wire n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706;
  wire n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714;
  wire n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722;
  wire n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730;
  wire n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738;
  wire n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746;
  wire n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754;
  wire n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762;
  wire n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770;
  wire n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778;
  wire n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786;
  wire n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794;
  wire n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802;
  wire n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810;
  wire n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818;
  wire n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826;
  wire n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834;
  wire n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842;
  wire n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850;
  wire n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858;
  wire n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866;
  wire n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874;
  wire n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882;
  wire n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890;
  wire n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898;
  wire n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906;
  wire n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914;
  wire n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922;
  wire n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930;
  wire n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938;
  wire n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946;
  wire n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954;
  wire n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962;
  wire n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970;
  wire n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978;
  wire n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986;
  wire n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994;
  wire n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002;
  wire n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010;
  wire n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018;
  wire n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026;
  wire n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034;
  wire n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042;
  wire n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050;
  wire n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058;
  wire n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066;
  wire n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074;
  wire n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082;
  wire n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090;
  wire n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098;
  wire n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106;
  wire n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114;
  wire n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122;
  wire n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130;
  wire n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138;
  wire n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146;
  wire n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154;
  wire n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162;
  wire n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170;
  wire n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178;
  wire n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186;
  wire n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194;
  wire n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202;
  wire n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210;
  wire n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218;
  wire n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226;
  wire n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234;
  wire n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242;
  wire n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250;
  wire n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258;
  wire n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266;
  wire n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274;
  wire n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282;
  wire n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290;
  wire n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298;
  wire n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306;
  wire n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314;
  wire n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322;
  wire n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330;
  wire n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338;
  wire n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346;
  wire n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354;
  wire n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362;
  wire n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370;
  wire n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378;
  wire n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386;
  wire n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394;
  wire n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402;
  wire n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410;
  wire n8414, n8415, n8416, n8417, n8418, n8419, n8422, n8423;
  wire n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431;
  wire n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439;
  wire n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447;
  wire n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455;
  wire n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463;
  wire n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471;
  wire n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479;
  wire n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487;
  wire n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495;
  wire n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503;
  wire n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511;
  wire n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519;
  wire n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527;
  wire n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535;
  wire n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543;
  wire n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551;
  wire n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559;
  wire n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567;
  wire n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575;
  wire n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583;
  wire n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591;
  wire n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599;
  wire n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607;
  wire n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615;
  wire n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623;
  wire n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631;
  wire n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639;
  wire n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647;
  wire n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655;
  wire n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663;
  wire n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671;
  wire n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679;
  wire n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687;
  wire n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695;
  wire n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703;
  wire n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711;
  wire n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719;
  wire n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727;
  wire n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735;
  wire n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743;
  wire n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751;
  wire n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759;
  wire n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767;
  wire n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775;
  wire n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783;
  wire n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791;
  wire n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799;
  wire n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807;
  wire n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815;
  wire n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823;
  wire n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831;
  wire n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839;
  wire n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847;
  wire n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855;
  wire n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863;
  wire n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871;
  wire n8872, n8873, n8874, n8875, n8876, n8878, n8879, n8880;
  wire n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888;
  wire n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896;
  wire n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904;
  wire n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913;
  wire n8914, n8915, n8916, n8919, n8920, n8921, n8922, n8930;
  wire n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938;
  wire n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950;
  wire n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958;
  wire n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966;
  wire n8967, n8971, n8972, n8974, n8975, n8976, n8977, n8978;
  wire n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986;
  wire n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994;
  wire n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002;
  wire n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010;
  wire n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018;
  wire n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026;
  wire n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034;
  wire n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042;
  wire n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050;
  wire n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058;
  wire n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066;
  wire n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074;
  wire n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082;
  wire n9083, n9088, n9089, n9090, n9091, n9092, n9093, n9094;
  wire n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102;
  wire n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110;
  wire n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118;
  wire n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126;
  wire n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134;
  wire n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142;
  wire n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150;
  wire n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158;
  wire n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166;
  wire n9167, n9168, n9171, n9172, n9173, n9174, n9175, n9176;
  wire n9177, n9178, n9181, n9182, n9183, n9184, n9185, n9186;
  wire n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194;
  wire n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202;
  wire n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210;
  wire n9211, n9212, n9215, n9216, n9217, n9218, n9219, n9220;
  wire n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228;
  wire n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236;
  wire n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244;
  wire n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252;
  wire n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260;
  wire n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268;
  wire n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276;
  wire n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284;
  wire n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292;
  wire n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300;
  wire n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308;
  wire n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316;
  wire n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324;
  wire n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332;
  wire n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340;
  wire n9341, n9342, n9345, n9346, n9347, n9348, n9349, n9350;
  wire n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358;
  wire n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366;
  wire n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374;
  wire n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382;
  wire n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390;
  wire n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398;
  wire n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406;
  wire n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414;
  wire n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422;
  wire n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430;
  wire n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438;
  wire n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446;
  wire n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454;
  wire n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462;
  wire n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470;
  wire n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478;
  wire n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486;
  wire n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494;
  wire n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502;
  wire n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510;
  wire n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518;
  wire n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526;
  wire n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534;
  wire n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542;
  wire n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550;
  wire n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558;
  wire n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566;
  wire n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574;
  wire n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582;
  wire n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590;
  wire n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598;
  wire n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606;
  wire n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614;
  wire n9615, n9616, n9617, n9618, n9621, n9622, n9623, n9624;
  wire n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632;
  wire n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640;
  wire n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648;
  wire n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656;
  wire n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664;
  wire n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672;
  wire n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680;
  wire n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688;
  wire n9689, n9691, n9692, n9693, n9694, n9695, n9696, n9697;
  wire n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705;
  wire n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713;
  wire n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721;
  wire n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729;
  wire n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737;
  wire n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745;
  wire n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753;
  wire n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761;
  wire n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769;
  wire n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777;
  wire n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785;
  wire n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793;
  wire n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801;
  wire n9802, n9803, n9804, n9805, n9808, n9809, n9810, n9811;
  wire n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819;
  wire n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827;
  wire n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835;
  wire n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843;
  wire n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851;
  wire n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859;
  wire n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9870;
  wire n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878;
  wire n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886;
  wire n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894;
  wire n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902;
  wire n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910;
  wire n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918;
  wire n9919, n9920, n9923, n9924, n9925, n9926, n9927, n9928;
  wire n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936;
  wire n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944;
  wire n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952;
  wire n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960;
  wire n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968;
  wire n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976;
  wire n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984;
  wire n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992;
  wire n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000;
  wire n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008;
  wire n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016;
  wire n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024;
  wire n10025, n10026, n10027, n10028, n10029, n10032, n10033, n10034;
  wire n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042;
  wire n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050;
  wire n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058;
  wire n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10067;
  wire n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075;
  wire n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083;
  wire n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091;
  wire n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099;
  wire n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109;
  wire n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117;
  wire n10120, n10121, n10122, n10123, n10126, n10127, n10130, n10131;
  wire n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139;
  wire n10140, n10143, n10144, n10145, n10147, n10150, n10151, n10152;
  wire n10153, n10157, n10158, n10159, n10160, n10161, n10162, n10163;
  wire n10164, n10165, n10166, n10167, n10169, n10170, n10171, n10172;
  wire n10173, n10174, n10181, n10182, n10183, n10184, n10185, n10186;
  wire n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198;
  wire n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207;
  wire n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215;
  wire n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223;
  wire n10224, n10225, n10226, n10227, n10228, n10229, n10232, n10233;
  wire n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241;
  wire n10242, n10243, n10244, n10245, n10246, n10247, n10256, n10259;
  wire n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10269;
  wire n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277;
  wire n10278, n10279, n10286, n10287, n10288, n10289, n10290, n10291;
  wire n10292, n10293, n10295, n10296, n10297, n10298, n10299, n10300;
  wire n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308;
  wire n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316;
  wire n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324;
  wire n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332;
  wire n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340;
  wire n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348;
  wire n10349, n10350, n10353, n10354, n10355, n10356, n10357, n10358;
  wire n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366;
  wire n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374;
  wire n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10384;
  wire n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10394;
  wire n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402;
  wire n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410;
  wire n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418;
  wire n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426;
  wire n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434;
  wire n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442;
  wire n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450;
  wire n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458;
  wire n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466;
  wire n10467, n10470, n10471, n10472, n10473, n10474, n10475, n10476;
  wire n10477, n10478, n10479, n10482, n10484, n10485, n10486, n10487;
  wire n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495;
  wire n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503;
  wire n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511;
  wire n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519;
  wire n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527;
  wire n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535;
  wire n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543;
  wire n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551;
  wire n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559;
  wire n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567;
  wire n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575;
  wire n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583;
  wire n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591;
  wire n10592, n10595, n10596, n10597, n10598, n10599, n10600, n10601;
  wire n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609;
  wire n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617;
  wire n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625;
  wire n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633;
  wire n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641;
  wire n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649;
  wire n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657;
  wire n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665;
  wire n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673;
  wire n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681;
  wire n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689;
  wire n10690, n10691, n10692, n10695, n10696, n10697, n10698, n10699;
  wire n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707;
  wire n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715;
  wire n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723;
  wire n10724, n10725, n10726, n10727, n10729, n10730, n10731, n10732;
  wire n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740;
  wire n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748;
  wire n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756;
  wire n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764;
  wire n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772;
  wire n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780;
  wire n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788;
  wire n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796;
  wire n10797, n10798, n10801, n10802, n10803, n10804, n10805, n10806;
  wire n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814;
  wire n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822;
  wire n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830;
  wire n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840;
  wire n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848;
  wire n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856;
  wire n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10866;
  wire n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874;
  wire n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882;
  wire n10883, n10884, n10885, n10886, n10887, n10888, n10891, n10892;
  wire n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900;
  wire n10901, n10902, n10903, n10904, n10905, n10907, n10908, n10909;
  wire n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917;
  wire n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925;
  wire n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933;
  wire n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941;
  wire n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949;
  wire n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957;
  wire n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965;
  wire n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975;
  wire n10976, n10977, n10978, n10979, n10980, n10982, n10983, n10984;
  wire n10986, n10987, n10988, n10989, n11000, n11001, n11002, n11003;
  wire n11004, n11006, n11010, n11011, n11012, n11013, n11014, n11017;
  wire n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025;
  wire n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033;
  wire n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041;
  wire n11042, n11043, n11044, n11045, n11046, n11047, n11051, n11052;
  wire n11057, n11058, n11059, n11060, n11061, n11066, n11067, n11068;
  wire n11069, n11070, n11071, n11072, n11076, n11077, n11078, n11079;
  wire n11080, n11081, n11082, n11085, n11086, n11090, n11091, n11092;
  wire n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100;
  wire n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11110;
  wire n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118;
  wire n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126;
  wire n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134;
  wire n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142;
  wire n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150;
  wire n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158;
  wire n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166;
  wire n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174;
  wire n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182;
  wire n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190;
  wire n11191, n11192, n11193, n11194, n11197, n11198, n11199, n11200;
  wire n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208;
  wire n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216;
  wire n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224;
  wire n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232;
  wire n11233, n11234, n11235, n11238, n11239, n11240, n11241, n11242;
  wire n11243, n11244, n11245, n11246, n11247, n11250, n11251, n11252;
  wire n11255, n11256, n11257, n11258, n11259, n11261, n11262, n11263;
  wire n11264, n11267, n11268, n11269, n11273, n11281, n11282, n11283;
  wire n11284, n11287, n11288, n11289, n11290, n11291, n11293, n11294;
  wire n11295, n11299, n11300, n11301, n11302, n11303, n11304, n11305;
  wire n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11315;
  wire n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323;
  wire n11325, n11326, n11328, n11329, n11330, n11331, n11332, n11337;
  wire n11340, n11341, n11343, n11344, n11345, n11346, n11348, n11349;
  wire n11350, n11351, n11353, n11354, n11355, n11356, n11357, n11359;
  wire n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367;
  wire n11369, n11373, n11374, n11375, n11376, n11379, n11382, n11383;
  wire n11384, n11385, n11386, n11387, n11388, n11395, n11396, n11397;
  wire n11398, n11399, n11400, n11401, n11403, n11404, n11405, n11409;
  wire n11413, n11414, n11416, n11417, n11418, n11419, n11420, n11421;
  wire n11422, n11423, n11424, n11425, n11426, n11427, n11430, n11431;
  wire n11432, n11433, n11434, n11436, n11437, n11438, n11439, n11440;
  wire n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448;
  wire n11452, n11455, n11456, n11458, n11459, n11460, n11463, n11464;
  wire n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11473;
  wire n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481;
  wire n11482, n11483, n11485, n11486, n11487, n11488, n11489, n11490;
  wire n11491, n11497, n11498, n11500, n11501, n11502, n11503, n11504;
  wire n11505, n11506, n11507, n11508, n11510, n11511, n11512, n11513;
  wire n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521;
  wire n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529;
  wire n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537;
  wire n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545;
  wire n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553;
  wire n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561;
  wire n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569;
  wire n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577;
  wire n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585;
  wire n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593;
  wire n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601;
  wire n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609;
  wire n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617;
  wire n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625;
  wire n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633;
  wire n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641;
  wire n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649;
  wire n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657;
  wire n11658, n11659, n11660, n11661, n11663, n11664, n11665, n11666;
  wire n11667, n11668, n11669, n11670, n11671, n11673, n11675, n11676;
  wire n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684;
  wire n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692;
  wire n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700;
  wire n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708;
  wire n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716;
  wire n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724;
  wire n11725, n11726, n11727, n11728, n11729, n11730, n11733, n11734;
  wire n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742;
  wire n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750;
  wire n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11760;
  wire n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768;
  wire n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776;
  wire n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784;
  wire n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794;
  wire n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802;
  wire n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810;
  wire n11811, n11812, n11813, n11814, n11815, n11818, n11819, n11820;
  wire n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828;
  wire n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839;
  wire n11840, n11841, n11842, n11845, n11846, n11847, n11848, n11849;
  wire n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857;
  wire n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865;
  wire n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11875;
  wire n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883;
  wire n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891;
  wire n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899;
  wire n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907;
  wire n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915;
  wire n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923;
  wire n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931;
  wire n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939;
  wire n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947;
  wire n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955;
  wire n11956, n11959, n11960, n11961, n11962, n11963, n11964, n11965;
  wire n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973;
  wire n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981;
  wire n11982, n11983, n11984, n11987, n11988, n11989, n11990, n11991;
  wire n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999;
  wire n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007;
  wire n12008, n12011, n12012, n12013, n12014, n12015, n12016, n12017;
  wire n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025;
  wire n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035;
  wire n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043;
  wire n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051;
  wire n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059;
  wire n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067;
  wire n12068, n12069, n12070, n12071, n12072, n12073, n12077, n12078;
  wire n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086;
  wire n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094;
  wire n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102;
  wire n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110;
  wire n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118;
  wire n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126;
  wire n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134;
  wire n12135, n12136, n12137, n12138, n12139, n12140, n12144, n12145;
  wire n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153;
  wire n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161;
  wire n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169;
  wire n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12178;
  wire n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186;
  wire n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194;
  wire n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202;
  wire n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210;
  wire n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218;
  wire n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226;
  wire n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234;
  wire n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242;
  wire n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250;
  wire n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258;
  wire n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266;
  wire n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274;
  wire n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282;
  wire n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290;
  wire n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298;
  wire n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306;
  wire n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314;
  wire n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322;
  wire n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330;
  wire n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338;
  wire n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346;
  wire n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354;
  wire n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362;
  wire n12363, n12366, n12367, n12368, n12369, n12370, n12371, n12372;
  wire n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380;
  wire n12381, n12385, n12386, n12387, n12388, n12389, n12390, n12391;
  wire n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399;
  wire n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407;
  wire n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415;
  wire n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423;
  wire n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431;
  wire n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439;
  wire n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447;
  wire n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455;
  wire n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463;
  wire n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471;
  wire n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479;
  wire n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487;
  wire n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495;
  wire n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503;
  wire n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511;
  wire n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519;
  wire n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527;
  wire n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535;
  wire n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543;
  wire n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551;
  wire n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559;
  wire n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567;
  wire n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575;
  wire n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583;
  wire n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591;
  wire n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599;
  wire n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607;
  wire n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615;
  wire n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623;
  wire n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631;
  wire n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639;
  wire n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647;
  wire n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655;
  wire n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663;
  wire n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671;
  wire n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679;
  wire n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687;
  wire n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695;
  wire n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703;
  wire n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711;
  wire n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719;
  wire n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727;
  wire n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735;
  wire n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743;
  wire n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751;
  wire n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759;
  wire n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767;
  wire n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775;
  wire n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783;
  wire n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791;
  wire n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799;
  wire n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807;
  wire n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815;
  wire n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823;
  wire n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831;
  wire n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839;
  wire n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847;
  wire n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855;
  wire n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863;
  wire n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871;
  wire n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879;
  wire n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887;
  wire n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895;
  wire n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903;
  wire n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911;
  wire n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919;
  wire n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927;
  wire n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935;
  wire n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943;
  wire n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951;
  wire n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959;
  wire n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967;
  wire n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975;
  wire n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983;
  wire n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991;
  wire n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999;
  wire n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007;
  wire n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015;
  wire n13016, n13017, n13018, n13019, n13020, n13021, n13024, n13025;
  wire n13026, n13027, n13029, n13030, n13031, n13036, n13037, n13039;
  wire n13040, n13043, n13044, n13045, n13047, n13048, n13049, n13050;
  wire n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058;
  wire n13059, n13061, n13062, n13063, n13064, n13065, n13067, n13068;
  wire n13069, n13070, n13072, n13073, n13074, n13076, n13077, n13078;
  wire n13080, n13085, n13086, n13087, n13088, n13089, n13090, n13091;
  wire n13092, n13093, n13096, n13097, n13098, n13102, n13103, n13104;
  wire n13105, n13106, n13110, n13111, n13115, n13116, n13117, n13118;
  wire n13122, n13123, n13124, n13125, n13127, n13128, n13129, n13130;
  wire n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13139;
  wire n13140, n13141, n13142, n13143, n13144, n13146, n13147, n13148;
  wire n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156;
  wire n13157, n13158, n13159, n13160, n13161, n13162, n13164, n13165;
  wire n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173;
  wire n13174, n13175, n13176, n13177, n13178, n13180, n13181, n13182;
  wire n13186, n13187, n13188, n13189, n13193, n13194, n13195, n13198;
  wire n13199, n13201, n13202, n13206, n13207, n13208, n13211, n13212;
  wire n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220;
  wire n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228;
  wire n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236;
  wire n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244;
  wire n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252;
  wire n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260;
  wire n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13270;
  wire n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278;
  wire n13279, n13280, n13281, n13283, n13284, n13285, n13286, n13287;
  wire n13288, n13289, n13290, n13293, n13296, n13297, n13298, n13300;
  wire n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308;
  wire n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316;
  wire n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324;
  wire n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332;
  wire n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340;
  wire n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348;
  wire n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356;
  wire n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364;
  wire n13365, n13368, n13369, n13370, n13371, n13372, n13373, n13374;
  wire n13375, n13376, n13377, n13378, n13379, n13381, n13383, n13384;
  wire n13385, n13386, n13387, n13388, n13389, n13391, n13392, n13393;
  wire n13394, n13395, n13398, n13399, n13402, n13403, n13404, n13405;
  wire n13406, n13407, n13409, n13410, n13411, n13412, n13413, n13414;
  wire n13415, n13416, n13417, n13419, n13421, n13422, n13423, n13424;
  wire n13425, n13426, n13429, n13430, n13431, n13432, n13433, n13434;
  wire n13435, n13436, n13437, n13439, n13446, n13447, n13448, n13449;
  wire n13450, n13452, n13453, n13454, n13455, n13456, n13459, n13460;
  wire n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468;
  wire n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476;
  wire n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484;
  wire n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492;
  wire n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500;
  wire n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508;
  wire n13509, n13510, n13512, n13513, n13514, n13515, n13516, n13517;
  wire n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525;
  wire n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533;
  wire n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541;
  wire n13542, n13543, n13544, n13545, n13548, n13549, n13550, n13551;
  wire n13552, n13553, n13555, n13556, n13557, n13558, n13559, n13560;
  wire n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568;
  wire n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576;
  wire n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584;
  wire n13585, n13586, n13587, n13590, n13591, n13592, n13593, n13594;
  wire n13595, n13597, n13598, n13599, n13600, n13601, n13602, n13603;
  wire n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611;
  wire n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619;
  wire n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627;
  wire n13628, n13629, n13630, n13633, n13634, n13635, n13636, n13637;
  wire n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645;
  wire n13646, n13648, n13649, n13650, n13651, n13652, n13653, n13654;
  wire n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662;
  wire n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671;
  wire n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679;
  wire n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687;
  wire n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695;
  wire n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703;
  wire n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711;
  wire n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719;
  wire n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727;
  wire n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735;
  wire n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743;
  wire n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751;
  wire n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759;
  wire n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767;
  wire n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775;
  wire n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783;
  wire n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791;
  wire n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799;
  wire n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807;
  wire n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815;
  wire n13816, n13817, n13820, n13821, n13822, n13823, n13824, n13825;
  wire n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833;
  wire n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841;
  wire n13842, n13843, n13844, n13847, n13848, n13849, n13850, n13851;
  wire n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859;
  wire n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867;
  wire n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875;
  wire n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883;
  wire n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891;
  wire n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899;
  wire n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907;
  wire n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915;
  wire n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923;
  wire n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931;
  wire n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939;
  wire n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947;
  wire n13948, n13953, n13954, n13955, n13956, n13957, n13958, n13959;
  wire n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967;
  wire n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976;
  wire n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984;
  wire n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992;
  wire n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002;
  wire n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010;
  wire n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018;
  wire n14019, n14020, n14021, n14022, n14024, n14025, n14026, n14027;
  wire n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035;
  wire n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043;
  wire n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051;
  wire n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059;
  wire n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067;
  wire n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075;
  wire n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083;
  wire n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091;
  wire n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099;
  wire n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107;
  wire n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115;
  wire n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123;
  wire n14124, n14125, n14126, n14127, n14128, n14131, n14132, n14133;
  wire n14134, n14135, n14138, n14139, n14140, n14141, n14142, n14143;
  wire n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151;
  wire n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159;
  wire n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167;
  wire n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175;
  wire n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183;
  wire n14184, n14192, n14193, n14194, n14195, n14196, n14197, n14198;
  wire n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206;
  wire n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214;
  wire n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222;
  wire n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230;
  wire n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238;
  wire n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246;
  wire n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254;
  wire n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262;
  wire n14263, n14264, n14265, n14268, n14269, n14270, n14271, n14274;
  wire n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282;
  wire n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290;
  wire n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298;
  wire n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306;
  wire n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314;
  wire n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322;
  wire n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330;
  wire n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338;
  wire n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346;
  wire n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354;
  wire n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362;
  wire n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370;
  wire n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378;
  wire n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386;
  wire n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394;
  wire n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402;
  wire n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410;
  wire n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418;
  wire n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14427;
  wire n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435;
  wire n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443;
  wire n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451;
  wire n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459;
  wire n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467;
  wire n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475;
  wire n14476, n14477, n14478, n14479, n14480, n14483, n14484, n14485;
  wire n14486, n14487, n14490, n14491, n14492, n14493, n14494, n14495;
  wire n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503;
  wire n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511;
  wire n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519;
  wire n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527;
  wire n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535;
  wire n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543;
  wire n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551;
  wire n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559;
  wire n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567;
  wire n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575;
  wire n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583;
  wire n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591;
  wire n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599;
  wire n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607;
  wire n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615;
  wire n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623;
  wire n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631;
  wire n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639;
  wire n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647;
  wire n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655;
  wire n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663;
  wire n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671;
  wire n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679;
  wire n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687;
  wire n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695;
  wire n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703;
  wire n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711;
  wire n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719;
  wire n14720, n14723, n14724, n14725, n14726, n14727, n14728, n14729;
  wire n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737;
  wire n14738, n14741, n14742, n14743, n14744, n14745, n14746, n14747;
  wire n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755;
  wire n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763;
  wire n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771;
  wire n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779;
  wire n14780, n14781, n14784, n14785, n14786, n14787, n14788, n14789;
  wire n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797;
  wire n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805;
  wire n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813;
  wire n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821;
  wire n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829;
  wire n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837;
  wire n14838, n14839, n14840, n14843, n14844, n14845, n14847, n14848;
  wire n14849, n14850, n14851, n14852, n14853, n14857, n14858, n14859;
  wire n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867;
  wire n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875;
  wire n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883;
  wire n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891;
  wire n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899;
  wire n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907;
  wire n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916;
  wire n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924;
  wire n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932;
  wire n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940;
  wire n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948;
  wire n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956;
  wire n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964;
  wire n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972;
  wire n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980;
  wire n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988;
  wire n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996;
  wire n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004;
  wire n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012;
  wire n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020;
  wire n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028;
  wire n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036;
  wire n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15046;
  wire n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054;
  wire n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062;
  wire n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070;
  wire n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078;
  wire n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086;
  wire n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094;
  wire n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102;
  wire n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110;
  wire n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118;
  wire n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126;
  wire n15127, n15128, n15129, n15130, n15131, n15134, n15135, n15136;
  wire n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144;
  wire n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152;
  wire n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160;
  wire n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168;
  wire n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176;
  wire n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184;
  wire n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15194;
  wire n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202;
  wire n15203, n15204, n15207, n15208, n15209, n15210, n15211, n15212;
  wire n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220;
  wire n15221, n15222, n15223, n15224, n15225, n15226, n15229, n15230;
  wire n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238;
  wire n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246;
  wire n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254;
  wire n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262;
  wire n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270;
  wire n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278;
  wire n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286;
  wire n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294;
  wire n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302;
  wire n15303, n15304, n15305, n15306, n15307, n15308, n15311, n15312;
  wire n15313, n15315, n15316, n15317, n15318, n15319, n15320, n15321;
  wire n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329;
  wire n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337;
  wire n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345;
  wire n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353;
  wire n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361;
  wire n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369;
  wire n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377;
  wire n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385;
  wire n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393;
  wire n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401;
  wire n15402, n15403, n15404, n15405, n15408, n15409, n15410, n15411;
  wire n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419;
  wire n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427;
  wire n15428, n15429, n15430, n15431, n15432, n15435, n15436, n15437;
  wire n15438, n15439, n15440, n15441, n15442, n15445, n15446, n15447;
  wire n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455;
  wire n15456, n15457, n15460, n15461, n15462, n15463, n15464, n15465;
  wire n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473;
  wire n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481;
  wire n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489;
  wire n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497;
  wire n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505;
  wire n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513;
  wire n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521;
  wire n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531;
  wire n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15541;
  wire n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549;
  wire n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557;
  wire n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565;
  wire n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573;
  wire n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581;
  wire n15582, n15583, n15584, n15587, n15588, n15589, n15590, n15591;
  wire n15592, n15593, n15596, n15597, n15598, n15599, n15600, n15601;
  wire n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609;
  wire n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15618;
  wire n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626;
  wire n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634;
  wire n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642;
  wire n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650;
  wire n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658;
  wire n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666;
  wire n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674;
  wire n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682;
  wire n15683, n15684, n15687, n15688, n15689, n15690, n15691, n15692;
  wire n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700;
  wire n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708;
  wire n15709, n15710, n15712, n15713, n15714, n15715, n15718, n15719;
  wire n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727;
  wire n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735;
  wire n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744;
  wire n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752;
  wire n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760;
  wire n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768;
  wire n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15778;
  wire n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788;
  wire n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796;
  wire n15797, n15798, n15799, n15802, n15803, n15804, n15805, n15806;
  wire n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814;
  wire n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822;
  wire n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830;
  wire n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838;
  wire n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846;
  wire n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854;
  wire n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862;
  wire n15863, n15864, n15865, n15866, n15867, n15870, n15872, n15873;
  wire n15874, n15875, n15876, n15877, n15878, n15880, n15881, n15882;
  wire n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890;
  wire n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898;
  wire n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906;
  wire n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914;
  wire n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922;
  wire n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930;
  wire n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938;
  wire n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946;
  wire n15947, n15948, n15949, n15950, n15953, n15954, n15955, n15956;
  wire n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964;
  wire n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972;
  wire n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980;
  wire n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988;
  wire n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996;
  wire n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004;
  wire n16005, n16006, n16007, n16008, n16011, n16012, n16013, n16014;
  wire n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022;
  wire n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030;
  wire n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038;
  wire n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046;
  wire n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054;
  wire n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062;
  wire n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070;
  wire n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078;
  wire n16079, n16082, n16083, n16084, n16085, n16086, n16089, n16092;
  wire n16093, n16094, n16096, n16097, n16098, n16099, n16100, n16101;
  wire n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109;
  wire n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117;
  wire n16118, n16119, n16120, n16121, n16122, n16123, n16126, n16127;
  wire n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135;
  wire n16136, n16137, n16138, n16139, n16140, n16143, n16146, n16147;
  wire n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155;
  wire n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164;
  wire n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172;
  wire n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180;
  wire n16181, n16182, n16183, n16184, n16185, n16188, n16189, n16190;
  wire n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198;
  wire n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206;
  wire n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214;
  wire n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222;
  wire n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230;
  wire n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238;
  wire n16239, n16240, n16241, n16242, n16245, n16246, n16247, n16248;
  wire n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256;
  wire n16257, n16258, n16261, n16262, n16263, n16264, n16265, n16266;
  wire n16267, n16268, n16269, n16271, n16272, n16273, n16274, n16275;
  wire n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283;
  wire n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291;
  wire n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299;
  wire n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307;
  wire n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315;
  wire n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323;
  wire n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331;
  wire n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339;
  wire n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347;
  wire n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355;
  wire n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363;
  wire n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371;
  wire n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379;
  wire n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387;
  wire n16388, n16390, n16391, n16392, n16393, n16394, n16395, n16396;
  wire n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404;
  wire n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412;
  wire n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420;
  wire n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428;
  wire n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436;
  wire n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444;
  wire n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452;
  wire n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460;
  wire n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468;
  wire n16469, n16470, n16471, n16472, n16473, n16474, n16476, n16477;
  wire n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485;
  wire n16486, n16487, n16489, n16490, n16491, n16492, n16493, n16494;
  wire n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502;
  wire n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510;
  wire n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518;
  wire n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526;
  wire n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534;
  wire n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542;
  wire n16543, n16544, n16545, n16546, n16549, n16550, n16551, n16552;
  wire n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560;
  wire n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568;
  wire n16569, n16570, n16571, n16572, n16574, n16575, n16576, n16577;
  wire n16578, n16581, n16582, n16583, n16584, n16585, n16586, n16587;
  wire n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595;
  wire n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603;
  wire n16604, n16607, n16608, n16609, n16610, n16611, n16612, n16613;
  wire n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621;
  wire n16622, n16623, n16624, n16625, n16626, n16628, n16629, n16630;
  wire n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638;
  wire n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646;
  wire n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654;
  wire n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662;
  wire n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670;
  wire n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678;
  wire n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686;
  wire n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694;
  wire n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702;
  wire n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710;
  wire n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718;
  wire n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726;
  wire n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734;
  wire n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742;
  wire n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750;
  wire n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758;
  wire n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766;
  wire n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774;
  wire n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782;
  wire n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790;
  wire n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798;
  wire n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806;
  wire n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814;
  wire n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822;
  wire n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830;
  wire n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838;
  wire n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846;
  wire n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854;
  wire n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862;
  wire n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870;
  wire n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878;
  wire n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886;
  wire n16887, n16889, n16890, n16891, n16892, n16893, n16894, n16895;
  wire n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903;
  wire n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911;
  wire n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919;
  wire n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927;
  wire n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935;
  wire n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943;
  wire n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951;
  wire n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959;
  wire n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967;
  wire n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975;
  wire n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983;
  wire n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991;
  wire n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999;
  wire n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007;
  wire n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015;
  wire n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023;
  wire n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031;
  wire n17032, n17033, n17036, n17037, n17038, n17039, n17040, n17041;
  wire n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049;
  wire n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057;
  wire n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065;
  wire n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073;
  wire n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081;
  wire n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089;
  wire n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097;
  wire n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105;
  wire n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113;
  wire n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121;
  wire n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129;
  wire n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137;
  wire n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145;
  wire n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153;
  wire n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161;
  wire n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169;
  wire n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177;
  wire n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185;
  wire n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193;
  wire n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201;
  wire n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209;
  wire n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217;
  wire n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225;
  wire n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233;
  wire n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241;
  wire n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249;
  wire n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257;
  wire n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265;
  wire n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273;
  wire n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281;
  wire n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289;
  wire n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297;
  wire n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305;
  wire n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313;
  wire n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321;
  wire n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329;
  wire n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337;
  wire n17338, n17339, n17340, n17343, n17344, n17345, n17346, n17347;
  wire n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355;
  wire n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363;
  wire n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371;
  wire n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379;
  wire n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387;
  wire n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395;
  wire n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403;
  wire n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411;
  wire n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419;
  wire n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427;
  wire n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435;
  wire n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443;
  wire n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451;
  wire n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459;
  wire n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467;
  wire n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475;
  wire n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483;
  wire n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491;
  wire n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499;
  wire n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507;
  wire n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515;
  wire n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523;
  wire n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531;
  wire n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539;
  wire n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547;
  wire n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555;
  wire n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563;
  wire n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571;
  wire n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579;
  wire n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587;
  wire n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595;
  wire n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603;
  wire n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611;
  wire n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619;
  wire n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627;
  wire n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635;
  wire n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643;
  wire n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651;
  wire n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659;
  wire n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667;
  wire n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675;
  wire n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683;
  wire n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691;
  wire n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699;
  wire n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707;
  wire n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715;
  wire n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723;
  wire n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731;
  wire n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739;
  wire n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747;
  wire n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755;
  wire n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763;
  wire n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771;
  wire n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779;
  wire n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787;
  wire n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795;
  wire n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803;
  wire n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811;
  wire n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819;
  wire n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827;
  wire n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835;
  wire n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843;
  wire n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851;
  wire n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859;
  wire n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867;
  wire n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875;
  wire n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883;
  wire n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891;
  wire n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899;
  wire n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907;
  wire n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915;
  wire n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923;
  wire n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931;
  wire n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939;
  wire n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947;
  wire n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955;
  wire n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963;
  wire n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971;
  wire n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979;
  wire n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987;
  wire n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995;
  wire n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003;
  wire n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011;
  wire n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019;
  wire n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027;
  wire n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035;
  wire n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043;
  wire n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051;
  wire n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059;
  wire n18060, n18061, n18062, n18063, n18064, n18066, n18067, n18068;
  wire n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076;
  wire n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084;
  wire n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092;
  wire n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100;
  wire n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108;
  wire n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116;
  wire n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124;
  wire n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132;
  wire n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140;
  wire n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148;
  wire n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156;
  wire n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164;
  wire n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172;
  wire n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180;
  wire n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188;
  wire n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196;
  wire n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204;
  wire n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212;
  wire n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220;
  wire n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228;
  wire n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236;
  wire n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244;
  wire n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252;
  wire n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260;
  wire n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268;
  wire n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276;
  wire n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284;
  wire n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292;
  wire n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300;
  wire n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308;
  wire n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316;
  wire n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324;
  wire n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332;
  wire n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340;
  wire n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348;
  wire n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356;
  wire n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364;
  wire n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372;
  wire n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380;
  wire n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388;
  wire n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396;
  wire n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404;
  wire n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412;
  wire n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420;
  wire n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428;
  wire n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436;
  wire n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444;
  wire n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452;
  wire n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460;
  wire n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468;
  wire n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476;
  wire n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484;
  wire n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492;
  wire n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500;
  wire n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508;
  wire n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516;
  wire n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524;
  wire n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532;
  wire n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540;
  wire n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548;
  wire n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556;
  wire n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564;
  wire n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572;
  wire n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580;
  wire n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588;
  wire n18589, n18591, n18592, n18593, n18594, n18595, n18596, n18597;
  wire n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605;
  wire n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613;
  wire n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621;
  wire n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629;
  wire n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637;
  wire n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645;
  wire n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653;
  wire n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661;
  wire n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669;
  wire n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677;
  wire n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685;
  wire n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693;
  wire n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701;
  wire n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709;
  wire n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717;
  wire n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725;
  wire n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733;
  wire n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741;
  wire n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749;
  wire n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757;
  wire n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765;
  wire n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773;
  wire n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781;
  wire n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789;
  wire n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797;
  wire n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805;
  wire n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813;
  wire n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821;
  wire n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829;
  wire n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837;
  wire n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845;
  wire n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853;
  wire n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861;
  wire n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869;
  wire n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877;
  wire n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885;
  wire n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893;
  wire n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901;
  wire n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909;
  wire n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917;
  wire n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925;
  wire n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933;
  wire n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941;
  wire n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949;
  wire n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957;
  wire n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965;
  wire n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973;
  wire n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981;
  wire n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989;
  wire n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997;
  wire n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005;
  wire n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013;
  wire n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021;
  wire n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029;
  wire n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037;
  wire n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045;
  wire n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053;
  wire n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061;
  wire n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069;
  wire n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077;
  wire n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085;
  wire n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093;
  wire n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101;
  wire n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109;
  wire n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117;
  wire n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125;
  wire n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133;
  wire n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141;
  wire n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149;
  wire n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157;
  wire n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165;
  wire n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173;
  wire n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181;
  wire n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189;
  wire n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197;
  wire n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205;
  wire n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213;
  wire n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221;
  wire n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229;
  wire n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237;
  wire n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245;
  wire n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253;
  wire n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261;
  wire n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269;
  wire n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277;
  wire n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285;
  wire n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293;
  wire n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301;
  wire n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309;
  wire n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317;
  wire n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325;
  wire n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333;
  wire n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341;
  wire n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349;
  wire n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357;
  wire n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19366;
  wire n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374;
  wire n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382;
  wire n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390;
  wire n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398;
  wire n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406;
  wire n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414;
  wire n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422;
  wire n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430;
  wire n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438;
  wire n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446;
  wire n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454;
  wire n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462;
  wire n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470;
  wire n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478;
  wire n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488;
  wire n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496;
  wire n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504;
  wire n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512;
  wire n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520;
  wire n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528;
  wire n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536;
  wire n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544;
  wire n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552;
  wire n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560;
  wire n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568;
  wire n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576;
  wire n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584;
  wire n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592;
  wire n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600;
  wire n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608;
  wire n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616;
  wire n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624;
  wire n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632;
  wire n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640;
  wire n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648;
  wire n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656;
  wire n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664;
  wire n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672;
  wire n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680;
  wire n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688;
  wire n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696;
  wire n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704;
  wire n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712;
  wire n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720;
  wire n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728;
  wire n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736;
  wire n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744;
  wire n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752;
  wire n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760;
  wire n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768;
  wire n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776;
  wire n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784;
  wire n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792;
  wire n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800;
  wire n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808;
  wire n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816;
  wire n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824;
  wire n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832;
  wire n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840;
  wire n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848;
  wire n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856;
  wire n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864;
  wire n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872;
  wire n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880;
  wire n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888;
  wire n19889, n19890, n19892, n19893, n19894, n19895, n19896, n19897;
  wire n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905;
  wire n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913;
  wire n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921;
  wire n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929;
  wire n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937;
  wire n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945;
  wire n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953;
  wire n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961;
  wire n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969;
  wire n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977;
  wire n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985;
  wire n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993;
  wire n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001;
  wire n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009;
  wire n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017;
  wire n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025;
  wire n20026, n20027, n20028, n20029, n20030, n20033, n20034, n20035;
  wire n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043;
  wire n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051;
  wire n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059;
  wire n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067;
  wire n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075;
  wire n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083;
  wire n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091;
  wire n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099;
  wire n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107;
  wire n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115;
  wire n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123;
  wire n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131;
  wire n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139;
  wire n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147;
  wire n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155;
  wire n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163;
  wire n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171;
  wire n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179;
  wire n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187;
  wire n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195;
  wire n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203;
  wire n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211;
  wire n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219;
  wire n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227;
  wire n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235;
  wire n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243;
  wire n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251;
  wire n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259;
  wire n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267;
  wire n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275;
  wire n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283;
  wire n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291;
  wire n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299;
  wire n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307;
  wire n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315;
  wire n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323;
  wire n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331;
  wire n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339;
  wire n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347;
  wire n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355;
  wire n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363;
  wire n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371;
  wire n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379;
  wire n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387;
  wire n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395;
  wire n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403;
  wire n20404, n20405, n20406, n20407, n20408, n20409, n20411, n20412;
  wire n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420;
  wire n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428;
  wire n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436;
  wire n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444;
  wire n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452;
  wire n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460;
  wire n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468;
  wire n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476;
  wire n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484;
  wire n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492;
  wire n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500;
  wire n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508;
  wire n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516;
  wire n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524;
  wire n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532;
  wire n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540;
  wire n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548;
  wire n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556;
  wire n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564;
  wire n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572;
  wire n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580;
  wire n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588;
  wire n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596;
  wire n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604;
  wire n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612;
  wire n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620;
  wire n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628;
  wire n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636;
  wire n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644;
  wire n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652;
  wire n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660;
  wire n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668;
  wire n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676;
  wire n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684;
  wire n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692;
  wire n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700;
  wire n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708;
  wire n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716;
  wire n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724;
  wire n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732;
  wire n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740;
  wire n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748;
  wire n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756;
  wire n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764;
  wire n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772;
  wire n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780;
  wire n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788;
  wire n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796;
  wire n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804;
  wire n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812;
  wire n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820;
  wire n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828;
  wire n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836;
  wire n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844;
  wire n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852;
  wire n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860;
  wire n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868;
  wire n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876;
  wire n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884;
  wire n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892;
  wire n20893, n20894, n20895, n20896, n20897, n20899, n20900, n20901;
  wire n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909;
  wire n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917;
  wire n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925;
  wire n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933;
  wire n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941;
  wire n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949;
  wire n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957;
  wire n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965;
  wire n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973;
  wire n20974, n20975, n20976, n20977, n20978, n20980, n20981, n20982;
  wire n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990;
  wire n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998;
  wire n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006;
  wire n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014;
  wire n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022;
  wire n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030;
  wire n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038;
  wire n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046;
  wire n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054;
  wire n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062;
  wire n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070;
  wire n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078;
  wire n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086;
  wire n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094;
  wire n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102;
  wire n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110;
  wire n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118;
  wire n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126;
  wire n21127, n21129, n21130, n21131, n21132, n21133, n21134, n21135;
  wire n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143;
  wire n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151;
  wire n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159;
  wire n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167;
  wire n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175;
  wire n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183;
  wire n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191;
  wire n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200;
  wire n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208;
  wire n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216;
  wire n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224;
  wire n21225, n21226, n21227, n21228, n21229, n21230, n21233, n21234;
  wire n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242;
  wire n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250;
  wire n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259;
  wire n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267;
  wire n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275;
  wire n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283;
  wire n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291;
  wire n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299;
  wire n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21308;
  wire n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316;
  wire n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324;
  wire n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332;
  wire n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340;
  wire n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348;
  wire n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356;
  wire n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364;
  wire n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372;
  wire n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380;
  wire n21381, n21382, n21383, n21384, n21386, n21387, n21388, n21389;
  wire n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397;
  wire n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405;
  wire n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413;
  wire n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421;
  wire n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429;
  wire n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437;
  wire n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445;
  wire n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453;
  wire n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461;
  wire n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469;
  wire n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477;
  wire n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485;
  wire n21486, n21487, n21489, n21490, n21491, n21492, n21493, n21494;
  wire n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502;
  wire n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510;
  wire n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518;
  wire n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526;
  wire n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534;
  wire n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542;
  wire n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550;
  wire n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558;
  wire n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566;
  wire n21567, n21568, n21570, n21571, n21572, n21573, n21574, n21575;
  wire n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583;
  wire n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591;
  wire n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599;
  wire n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607;
  wire n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615;
  wire n21616, n21617, n21618, n21619, n21620, n21622, n21623, n21624;
  wire n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632;
  wire n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640;
  wire n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648;
  wire n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656;
  wire n21657, n21658, n21659, n21660, n21662, n21663, n21664, n21665;
  wire n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673;
  wire n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681;
  wire n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689;
  wire n21690, n21692, n21693, n21694, n21695, n21696, n21697, n21698;
  wire n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706;
  wire n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714;
  wire n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722;
  wire n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730;
  wire n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738;
  wire n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746;
  wire n21747, n21749, n21750, n21751, n21752, n21753, n21754, n21755;
  wire n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763;
  wire n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771;
  wire n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779;
  wire n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787;
  wire n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795;
  wire n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803;
  wire n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812;
  wire n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820;
  wire n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828;
  wire n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836;
  wire n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844;
  wire n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852;
  wire n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21861;
  wire n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869;
  wire n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877;
  wire n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885;
  wire n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893;
  wire n21894, n21895, n21896, n21897, n21898, n21899, n21902, n21903;
  wire n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911;
  wire n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21920;
  wire n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928;
  wire n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936;
  wire n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944;
  wire n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952;
  wire n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960;
  wire n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968;
  wire n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976;
  wire n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984;
  wire n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992;
  wire n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000;
  wire n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008;
  wire n22009, n22010, n22011, n22012, n22013, n22015, n22016, n22017;
  wire n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025;
  wire n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033;
  wire n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041;
  wire n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049;
  wire n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057;
  wire n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065;
  wire n22066, n22067, n22068, n22070, n22071, n22072, n22073, n22074;
  wire n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082;
  wire n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090;
  wire n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098;
  wire n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106;
  wire n22107, n22110, n22111, n22112, n22113, n22114, n22115, n22116;
  wire n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124;
  wire n22125, n22126, n22128, n22129, n22130, n22131, n22132, n22133;
  wire n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141;
  wire n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149;
  wire n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157;
  wire n22158, n22159, n22162, n22163, n22164, n22165, n22166, n22168;
  wire n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176;
  wire n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184;
  wire n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192;
  wire n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22202;
  wire n22203, n22204, n22205, n22206, n22208, n22209, n22210, n22211;
  wire n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219;
  wire n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227;
  wire n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235;
  wire n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243;
  wire n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251;
  wire n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259;
  wire n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267;
  wire n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275;
  wire n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283;
  wire n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291;
  wire n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299;
  wire n22300, n22301, n22302, n22303, n22305, n22306, n22307, n22308;
  wire n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316;
  wire n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324;
  wire n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332;
  wire n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340;
  wire n22341, n22342, n22343, n22344, n22345, n22346, n22348, n22349;
  wire n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357;
  wire n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365;
  wire n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373;
  wire n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381;
  wire n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389;
  wire n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397;
  wire n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405;
  wire n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413;
  wire n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421;
  wire n22422, n22423, n22424, n22425, n22426, n22427, n22429, n22430;
  wire n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438;
  wire n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446;
  wire n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454;
  wire n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462;
  wire n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470;
  wire n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478;
  wire n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486;
  wire n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494;
  wire n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502;
  wire n22503, n22504, n22505, n22506, n22507, n22508, n22510, n22511;
  wire n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519;
  wire n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527;
  wire n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535;
  wire n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543;
  wire n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551;
  wire n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559;
  wire n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567;
  wire n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575;
  wire n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583;
  wire n22584, n22585, n22586, n22587, n22588, n22590, n22591, n22592;
  wire n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600;
  wire n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608;
  wire n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616;
  wire n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624;
  wire n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632;
  wire n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640;
  wire n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648;
  wire n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656;
  wire n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664;
  wire n22665, n22666, n22667, n22668, n22669, n22671, n22672, n22673;
  wire n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681;
  wire n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689;
  wire n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697;
  wire n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705;
  wire n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713;
  wire n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721;
  wire n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729;
  wire n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737;
  wire n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745;
  wire n22746, n22747, n22748, n22749, n22750, n22752, n22753, n22754;
  wire n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762;
  wire n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770;
  wire n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778;
  wire n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786;
  wire n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794;
  wire n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802;
  wire n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810;
  wire n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818;
  wire n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826;
  wire n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834;
  wire n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842;
  wire n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850;
  wire n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858;
  wire n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866;
  wire n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874;
  wire n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882;
  wire n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890;
  wire n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898;
  wire n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906;
  wire n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914;
  wire n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922;
  wire n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930;
  wire n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938;
  wire n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946;
  wire n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954;
  wire n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962;
  wire n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970;
  wire n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978;
  wire n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986;
  wire n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994;
  wire n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002;
  wire n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010;
  wire n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018;
  wire n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026;
  wire n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034;
  wire n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042;
  wire n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050;
  wire n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058;
  wire n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066;
  wire n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074;
  wire n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082;
  wire n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090;
  wire n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098;
  wire n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106;
  wire n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114;
  wire n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122;
  wire n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130;
  wire n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138;
  wire n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146;
  wire n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154;
  wire n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162;
  wire n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170;
  wire n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178;
  wire n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186;
  wire n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194;
  wire n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202;
  wire n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210;
  wire n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218;
  wire n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23227;
  wire n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235;
  wire n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243;
  wire n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251;
  wire n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259;
  wire n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267;
  wire n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275;
  wire n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283;
  wire n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291;
  wire n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299;
  wire n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307;
  wire n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315;
  wire n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323;
  wire n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331;
  wire n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339;
  wire n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347;
  wire n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355;
  wire n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23365;
  wire n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373;
  wire n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381;
  wire n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389;
  wire n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397;
  wire n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405;
  wire n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413;
  wire n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421;
  wire n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429;
  wire n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437;
  wire n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445;
  wire n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453;
  wire n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461;
  wire n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469;
  wire n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477;
  wire n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485;
  wire n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493;
  wire n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501;
  wire n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509;
  wire n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517;
  wire n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525;
  wire n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533;
  wire n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541;
  wire n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549;
  wire n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557;
  wire n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565;
  wire n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573;
  wire n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581;
  wire n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589;
  wire n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597;
  wire n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605;
  wire n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613;
  wire n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621;
  wire n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629;
  wire n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637;
  wire n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645;
  wire n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653;
  wire n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661;
  wire n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669;
  wire n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677;
  wire n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685;
  wire n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693;
  wire n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701;
  wire n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709;
  wire n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718;
  wire n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726;
  wire n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734;
  wire n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742;
  wire n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750;
  wire n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758;
  wire n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766;
  wire n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774;
  wire n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782;
  wire n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790;
  wire n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798;
  wire n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806;
  wire n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814;
  wire n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822;
  wire n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830;
  wire n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838;
  wire n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846;
  wire n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854;
  wire n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862;
  wire n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870;
  wire n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878;
  wire n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886;
  wire n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894;
  wire n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902;
  wire n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910;
  wire n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918;
  wire n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926;
  wire n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934;
  wire n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942;
  wire n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950;
  wire n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958;
  wire n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966;
  wire n23967, n23968, n23969, n23970, n23971, n23972, n23975, n23976;
  wire n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984;
  wire n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992;
  wire n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000;
  wire n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008;
  wire n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016;
  wire n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024;
  wire n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032;
  wire n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040;
  wire n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048;
  wire n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056;
  wire n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064;
  wire n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072;
  wire n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080;
  wire n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088;
  wire n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096;
  wire n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104;
  wire n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112;
  wire n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120;
  wire n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128;
  wire n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136;
  wire n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144;
  wire n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152;
  wire n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160;
  wire n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168;
  wire n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176;
  wire n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184;
  wire n24185, n24186, n24187, n24189, n24190, n24191, n24192, n24193;
  wire n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201;
  wire n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209;
  wire n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217;
  wire n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225;
  wire n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233;
  wire n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241;
  wire n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249;
  wire n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257;
  wire n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265;
  wire n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273;
  wire n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281;
  wire n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289;
  wire n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297;
  wire n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305;
  wire n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313;
  wire n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321;
  wire n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329;
  wire n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337;
  wire n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345;
  wire n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353;
  wire n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361;
  wire n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369;
  wire n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377;
  wire n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385;
  wire n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393;
  wire n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401;
  wire n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409;
  wire n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417;
  wire n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425;
  wire n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433;
  wire n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441;
  wire n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449;
  wire n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457;
  wire n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465;
  wire n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473;
  wire n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481;
  wire n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489;
  wire n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497;
  wire n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505;
  wire n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513;
  wire n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521;
  wire n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529;
  wire n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537;
  wire n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545;
  wire n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553;
  wire n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561;
  wire n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569;
  wire n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577;
  wire n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585;
  wire n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593;
  wire n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601;
  wire n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609;
  wire n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617;
  wire n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625;
  wire n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633;
  wire n24634, n24635, n24636, n24637, n24639, n24640, n24641, n24642;
  wire n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650;
  wire n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658;
  wire n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666;
  wire n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674;
  wire n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682;
  wire n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690;
  wire n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698;
  wire n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706;
  wire n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714;
  wire n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722;
  wire n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730;
  wire n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738;
  wire n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746;
  wire n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754;
  wire n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762;
  wire n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770;
  wire n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778;
  wire n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786;
  wire n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794;
  wire n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802;
  wire n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810;
  wire n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818;
  wire n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826;
  wire n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834;
  wire n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842;
  wire n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850;
  wire n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858;
  wire n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866;
  wire n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874;
  wire n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882;
  wire n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890;
  wire n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898;
  wire n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906;
  wire n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914;
  wire n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922;
  wire n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930;
  wire n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938;
  wire n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946;
  wire n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954;
  wire n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962;
  wire n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970;
  wire n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978;
  wire n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986;
  wire n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994;
  wire n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002;
  wire n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010;
  wire n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018;
  wire n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026;
  wire n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034;
  wire n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042;
  wire n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050;
  wire n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058;
  wire n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066;
  wire n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074;
  wire n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082;
  wire n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090;
  wire n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098;
  wire n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106;
  wire n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114;
  wire n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25123;
  wire n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131;
  wire n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139;
  wire n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147;
  wire n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155;
  wire n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163;
  wire n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171;
  wire n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179;
  wire n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187;
  wire n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195;
  wire n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203;
  wire n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211;
  wire n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219;
  wire n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227;
  wire n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235;
  wire n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243;
  wire n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251;
  wire n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259;
  wire n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267;
  wire n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275;
  wire n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283;
  wire n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291;
  wire n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299;
  wire n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307;
  wire n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315;
  wire n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323;
  wire n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331;
  wire n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339;
  wire n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347;
  wire n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355;
  wire n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363;
  wire n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371;
  wire n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379;
  wire n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387;
  wire n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395;
  wire n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403;
  wire n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411;
  wire n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419;
  wire n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427;
  wire n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435;
  wire n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443;
  wire n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451;
  wire n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459;
  wire n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467;
  wire n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475;
  wire n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483;
  wire n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491;
  wire n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499;
  wire n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507;
  wire n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515;
  wire n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523;
  wire n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531;
  wire n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539;
  wire n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547;
  wire n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555;
  wire n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563;
  wire n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571;
  wire n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579;
  wire n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587;
  wire n25588, n25589, n25590, n25591, n25592, n25594, n25595, n25596;
  wire n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604;
  wire n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612;
  wire n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620;
  wire n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628;
  wire n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636;
  wire n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644;
  wire n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652;
  wire n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25662;
  wire n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670;
  wire n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678;
  wire n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686;
  wire n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694;
  wire n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702;
  wire n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710;
  wire n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718;
  wire n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726;
  wire n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734;
  wire n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742;
  wire n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750;
  wire n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758;
  wire n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766;
  wire n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774;
  wire n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782;
  wire n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790;
  wire n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798;
  wire n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806;
  wire n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814;
  wire n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822;
  wire n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830;
  wire n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838;
  wire n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846;
  wire n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854;
  wire n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862;
  wire n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870;
  wire n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878;
  wire n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886;
  wire n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894;
  wire n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902;
  wire n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910;
  wire n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918;
  wire n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926;
  wire n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934;
  wire n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942;
  wire n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950;
  wire n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958;
  wire n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966;
  wire n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974;
  wire n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982;
  wire n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990;
  wire n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998;
  wire n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006;
  wire n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014;
  wire n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022;
  wire n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030;
  wire n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038;
  wire n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046;
  wire n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054;
  wire n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062;
  wire n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070;
  wire n26071, n26072, n26073, n26074, n26076, n26077, n26078, n26079;
  wire n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087;
  wire n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095;
  wire n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103;
  wire n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111;
  wire n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119;
  wire n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127;
  wire n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135;
  wire n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143;
  wire n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151;
  wire n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159;
  wire n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167;
  wire n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175;
  wire n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183;
  wire n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191;
  wire n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199;
  wire n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207;
  wire n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215;
  wire n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223;
  wire n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231;
  wire n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239;
  wire n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247;
  wire n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255;
  wire n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263;
  wire n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271;
  wire n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279;
  wire n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287;
  wire n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295;
  wire n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303;
  wire n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311;
  wire n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319;
  wire n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327;
  wire n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335;
  wire n26336, n26337, n26338, n26341, n26342, n26343, n26344, n26345;
  wire n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353;
  wire n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361;
  wire n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369;
  wire n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377;
  wire n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385;
  wire n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393;
  wire n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401;
  wire n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409;
  wire n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417;
  wire n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425;
  wire n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433;
  wire n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441;
  wire n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449;
  wire n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457;
  wire n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465;
  wire n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473;
  wire n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481;
  wire n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489;
  wire n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497;
  wire n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505;
  wire n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513;
  wire n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521;
  wire n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529;
  wire n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537;
  wire n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545;
  wire n26546, n26547, n26548, n26549, n26550, n26551, n26553, n26554;
  wire n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562;
  wire n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570;
  wire n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578;
  wire n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586;
  wire n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594;
  wire n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602;
  wire n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610;
  wire n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618;
  wire n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626;
  wire n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634;
  wire n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642;
  wire n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650;
  wire n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658;
  wire n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666;
  wire n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674;
  wire n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682;
  wire n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690;
  wire n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698;
  wire n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706;
  wire n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714;
  wire n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722;
  wire n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730;
  wire n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738;
  wire n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746;
  wire n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754;
  wire n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762;
  wire n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770;
  wire n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778;
  wire n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786;
  wire n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794;
  wire n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802;
  wire n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810;
  wire n26811, n26812, n26813, n26814, n26815, n26818, n26819, n26820;
  wire n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828;
  wire n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836;
  wire n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844;
  wire n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852;
  wire n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860;
  wire n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868;
  wire n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876;
  wire n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884;
  wire n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892;
  wire n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900;
  wire n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908;
  wire n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916;
  wire n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924;
  wire n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932;
  wire n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940;
  wire n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948;
  wire n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956;
  wire n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964;
  wire n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972;
  wire n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980;
  wire n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988;
  wire n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996;
  wire n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004;
  wire n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012;
  wire n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020;
  wire n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028;
  wire n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037;
  wire n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045;
  wire n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053;
  wire n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061;
  wire n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069;
  wire n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077;
  wire n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085;
  wire n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093;
  wire n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101;
  wire n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109;
  wire n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117;
  wire n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125;
  wire n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133;
  wire n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141;
  wire n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149;
  wire n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157;
  wire n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165;
  wire n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173;
  wire n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181;
  wire n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189;
  wire n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197;
  wire n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205;
  wire n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213;
  wire n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221;
  wire n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229;
  wire n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237;
  wire n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245;
  wire n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253;
  wire n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261;
  wire n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269;
  wire n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277;
  wire n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285;
  wire n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293;
  wire n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301;
  wire n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309;
  wire n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317;
  wire n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325;
  wire n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333;
  wire n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341;
  wire n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349;
  wire n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357;
  wire n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365;
  wire n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373;
  wire n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381;
  wire n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389;
  wire n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397;
  wire n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405;
  wire n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413;
  wire n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421;
  wire n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429;
  wire n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437;
  wire n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445;
  wire n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453;
  wire n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461;
  wire n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469;
  wire n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477;
  wire n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485;
  wire n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493;
  wire n27494, n27495, n27496, n27497, n27498, n27499, n27501, n27502;
  wire n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510;
  wire n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518;
  wire n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526;
  wire n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534;
  wire n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542;
  wire n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550;
  wire n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558;
  wire n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566;
  wire n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574;
  wire n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582;
  wire n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590;
  wire n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598;
  wire n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606;
  wire n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614;
  wire n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622;
  wire n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630;
  wire n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638;
  wire n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646;
  wire n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654;
  wire n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662;
  wire n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670;
  wire n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678;
  wire n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686;
  wire n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694;
  wire n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702;
  wire n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710;
  wire n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718;
  wire n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726;
  wire n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734;
  wire n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742;
  wire n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750;
  wire n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758;
  wire n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766;
  wire n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774;
  wire n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782;
  wire n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790;
  wire n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798;
  wire n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806;
  wire n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814;
  wire n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822;
  wire n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830;
  wire n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838;
  wire n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846;
  wire n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854;
  wire n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862;
  wire n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870;
  wire n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878;
  wire n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886;
  wire n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894;
  wire n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902;
  wire n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910;
  wire n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918;
  wire n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926;
  wire n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934;
  wire n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942;
  wire n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950;
  wire n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958;
  wire n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966;
  wire n27967, n27968, n27969, n27970, n27972, n27973, n27974, n27975;
  wire n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983;
  wire n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991;
  wire n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999;
  wire n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007;
  wire n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015;
  wire n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023;
  wire n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031;
  wire n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039;
  wire n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047;
  wire n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055;
  wire n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063;
  wire n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071;
  wire n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079;
  wire n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087;
  wire n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095;
  wire n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103;
  wire n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111;
  wire n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119;
  wire n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127;
  wire n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135;
  wire n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143;
  wire n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151;
  wire n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159;
  wire n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167;
  wire n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175;
  wire n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183;
  wire n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191;
  wire n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199;
  wire n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207;
  wire n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215;
  wire n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223;
  wire n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231;
  wire n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239;
  wire n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247;
  wire n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255;
  wire n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263;
  wire n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271;
  wire n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279;
  wire n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287;
  wire n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295;
  wire n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303;
  wire n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311;
  wire n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319;
  wire n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327;
  wire n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335;
  wire n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343;
  wire n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351;
  wire n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359;
  wire n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367;
  wire n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375;
  wire n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383;
  wire n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391;
  wire n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399;
  wire n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407;
  wire n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415;
  wire n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423;
  wire n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431;
  wire n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439;
  wire n28440, n28441, n28443, n28444, n28445, n28446, n28447, n28448;
  wire n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456;
  wire n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464;
  wire n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472;
  wire n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480;
  wire n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488;
  wire n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496;
  wire n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504;
  wire n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512;
  wire n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520;
  wire n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528;
  wire n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536;
  wire n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544;
  wire n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552;
  wire n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560;
  wire n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568;
  wire n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576;
  wire n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584;
  wire n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592;
  wire n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600;
  wire n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608;
  wire n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616;
  wire n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624;
  wire n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632;
  wire n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640;
  wire n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648;
  wire n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656;
  wire n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664;
  wire n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672;
  wire n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680;
  wire n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688;
  wire n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696;
  wire n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704;
  wire n28705, n28708, n28709, n28710, n28711, n28712, n28713, n28714;
  wire n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722;
  wire n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730;
  wire n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738;
  wire n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746;
  wire n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754;
  wire n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762;
  wire n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770;
  wire n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778;
  wire n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786;
  wire n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794;
  wire n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802;
  wire n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810;
  wire n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818;
  wire n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826;
  wire n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834;
  wire n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842;
  wire n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850;
  wire n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858;
  wire n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866;
  wire n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874;
  wire n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882;
  wire n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890;
  wire n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898;
  wire n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906;
  wire n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914;
  wire n28915, n28916, n28917, n28918, n28920, n28921, n28922, n28923;
  wire n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931;
  wire n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939;
  wire n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947;
  wire n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955;
  wire n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963;
  wire n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971;
  wire n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979;
  wire n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987;
  wire n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995;
  wire n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003;
  wire n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011;
  wire n29012, n29013, n29016, n29017, n29018, n29019, n29020, n29021;
  wire n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029;
  wire n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037;
  wire n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045;
  wire n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053;
  wire n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061;
  wire n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069;
  wire n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077;
  wire n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085;
  wire n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093;
  wire n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101;
  wire n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109;
  wire n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117;
  wire n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125;
  wire n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133;
  wire n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141;
  wire n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149;
  wire n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157;
  wire n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165;
  wire n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173;
  wire n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181;
  wire n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189;
  wire n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197;
  wire n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205;
  wire n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213;
  wire n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221;
  wire n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229;
  wire n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237;
  wire n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245;
  wire n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253;
  wire n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261;
  wire n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269;
  wire n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277;
  wire n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285;
  wire n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293;
  wire n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301;
  wire n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309;
  wire n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317;
  wire n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325;
  wire n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333;
  wire n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341;
  wire n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349;
  wire n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357;
  wire n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365;
  wire n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373;
  wire n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381;
  wire n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389;
  wire n29390, n29391, n29392, n29393, n29395, n29396, n29397, n29398;
  wire n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406;
  wire n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414;
  wire n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422;
  wire n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430;
  wire n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438;
  wire n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446;
  wire n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454;
  wire n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462;
  wire n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470;
  wire n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478;
  wire n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486;
  wire n29487, n29488, n29491, n29492, n29493, n29494, n29495, n29496;
  wire n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504;
  wire n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512;
  wire n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520;
  wire n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528;
  wire n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536;
  wire n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544;
  wire n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552;
  wire n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560;
  wire n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568;
  wire n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576;
  wire n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584;
  wire n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592;
  wire n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600;
  wire n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608;
  wire n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616;
  wire n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624;
  wire n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632;
  wire n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640;
  wire n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648;
  wire n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656;
  wire n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664;
  wire n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672;
  wire n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680;
  wire n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688;
  wire n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696;
  wire n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704;
  wire n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712;
  wire n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720;
  wire n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728;
  wire n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736;
  wire n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744;
  wire n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752;
  wire n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760;
  wire n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768;
  wire n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776;
  wire n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784;
  wire n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792;
  wire n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800;
  wire n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808;
  wire n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816;
  wire n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824;
  wire n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832;
  wire n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840;
  wire n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848;
  wire n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856;
  wire n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864;
  wire n29865, n29866, n29867, n29868, n29870, n29871, n29872, n29873;
  wire n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881;
  wire n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889;
  wire n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897;
  wire n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905;
  wire n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913;
  wire n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921;
  wire n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929;
  wire n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937;
  wire n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945;
  wire n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953;
  wire n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961;
  wire n29962, n29963, n29966, n29967, n29968, n29969, n29970, n29971;
  wire n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979;
  wire n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987;
  wire n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995;
  wire n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003;
  wire n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011;
  wire n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019;
  wire n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027;
  wire n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035;
  wire n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043;
  wire n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051;
  wire n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059;
  wire n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067;
  wire n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075;
  wire n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083;
  wire n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091;
  wire n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099;
  wire n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107;
  wire n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115;
  wire n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123;
  wire n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131;
  wire n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139;
  wire n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147;
  wire n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155;
  wire n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163;
  wire n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171;
  wire n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179;
  wire n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187;
  wire n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195;
  wire n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203;
  wire n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211;
  wire n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219;
  wire n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227;
  wire n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235;
  wire n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243;
  wire n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251;
  wire n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259;
  wire n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267;
  wire n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275;
  wire n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283;
  wire n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291;
  wire n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299;
  wire n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307;
  wire n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315;
  wire n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323;
  wire n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331;
  wire n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339;
  wire n30340, n30341, n30342, n30343, n30345, n30346, n30347, n30348;
  wire n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356;
  wire n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364;
  wire n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372;
  wire n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380;
  wire n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388;
  wire n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396;
  wire n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404;
  wire n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412;
  wire n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420;
  wire n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428;
  wire n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436;
  wire n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444;
  wire n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452;
  wire n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460;
  wire n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468;
  wire n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476;
  wire n30477, n30478, n30479, n30480, n30483, n30484, n30485, n30486;
  wire n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494;
  wire n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502;
  wire n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510;
  wire n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518;
  wire n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526;
  wire n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534;
  wire n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542;
  wire n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550;
  wire n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558;
  wire n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566;
  wire n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574;
  wire n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582;
  wire n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590;
  wire n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598;
  wire n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606;
  wire n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614;
  wire n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622;
  wire n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630;
  wire n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638;
  wire n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646;
  wire n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654;
  wire n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662;
  wire n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670;
  wire n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678;
  wire n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686;
  wire n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694;
  wire n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702;
  wire n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710;
  wire n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718;
  wire n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726;
  wire n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734;
  wire n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742;
  wire n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750;
  wire n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758;
  wire n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766;
  wire n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774;
  wire n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782;
  wire n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790;
  wire n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798;
  wire n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806;
  wire n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814;
  wire n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822;
  wire n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831;
  wire n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839;
  wire n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847;
  wire n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855;
  wire n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863;
  wire n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871;
  wire n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879;
  wire n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887;
  wire n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895;
  wire n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903;
  wire n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911;
  wire n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919;
  wire n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927;
  wire n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935;
  wire n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943;
  wire n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951;
  wire n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959;
  wire n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967;
  wire n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975;
  wire n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983;
  wire n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991;
  wire n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999;
  wire n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007;
  wire n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015;
  wire n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023;
  wire n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031;
  wire n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039;
  wire n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047;
  wire n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055;
  wire n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063;
  wire n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071;
  wire n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079;
  wire n31080, n31081, n31082, n31083, n31084, n31085, n31088, n31089;
  wire n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097;
  wire n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105;
  wire n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113;
  wire n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121;
  wire n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129;
  wire n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137;
  wire n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145;
  wire n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153;
  wire n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161;
  wire n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169;
  wire n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177;
  wire n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185;
  wire n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193;
  wire n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201;
  wire n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209;
  wire n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217;
  wire n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225;
  wire n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233;
  wire n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241;
  wire n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249;
  wire n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257;
  wire n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265;
  wire n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273;
  wire n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281;
  wire n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289;
  wire n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297;
  wire n31298, n31299, n31301, n31302, n31303, n31304, n31305, n31306;
  wire n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314;
  wire n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322;
  wire n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330;
  wire n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338;
  wire n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346;
  wire n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354;
  wire n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362;
  wire n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370;
  wire n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378;
  wire n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386;
  wire n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394;
  wire n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402;
  wire n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410;
  wire n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418;
  wire n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426;
  wire n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434;
  wire n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442;
  wire n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450;
  wire n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458;
  wire n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466;
  wire n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474;
  wire n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482;
  wire n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490;
  wire n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498;
  wire n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506;
  wire n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514;
  wire n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522;
  wire n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530;
  wire n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538;
  wire n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546;
  wire n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554;
  wire n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562;
  wire n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572;
  wire n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580;
  wire n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588;
  wire n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596;
  wire n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604;
  wire n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612;
  wire n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620;
  wire n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628;
  wire n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636;
  wire n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644;
  wire n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652;
  wire n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660;
  wire n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668;
  wire n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676;
  wire n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684;
  wire n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692;
  wire n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700;
  wire n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708;
  wire n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716;
  wire n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724;
  wire n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732;
  wire n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740;
  wire n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748;
  wire n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756;
  wire n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764;
  wire n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772;
  wire n31773, n31774, n31775, n31776, n31778, n31779, n31780, n31781;
  wire n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789;
  wire n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797;
  wire n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805;
  wire n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813;
  wire n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821;
  wire n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829;
  wire n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837;
  wire n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845;
  wire n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853;
  wire n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861;
  wire n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869;
  wire n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877;
  wire n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885;
  wire n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893;
  wire n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901;
  wire n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909;
  wire n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917;
  wire n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925;
  wire n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933;
  wire n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941;
  wire n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949;
  wire n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957;
  wire n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965;
  wire n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973;
  wire n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981;
  wire n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989;
  wire n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997;
  wire n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005;
  wire n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013;
  wire n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021;
  wire n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029;
  wire n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037;
  wire n32038, n32039, n32042, n32043, n32044, n32045, n32046, n32047;
  wire n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055;
  wire n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063;
  wire n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071;
  wire n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079;
  wire n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087;
  wire n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095;
  wire n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103;
  wire n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111;
  wire n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119;
  wire n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127;
  wire n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135;
  wire n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143;
  wire n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151;
  wire n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159;
  wire n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167;
  wire n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175;
  wire n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183;
  wire n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191;
  wire n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199;
  wire n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207;
  wire n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215;
  wire n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223;
  wire n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231;
  wire n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239;
  wire n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247;
  wire n32248, n32249, n32250, n32251, n32252, n32253, n32255, n32256;
  wire n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264;
  wire n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272;
  wire n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280;
  wire n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288;
  wire n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296;
  wire n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304;
  wire n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312;
  wire n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320;
  wire n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328;
  wire n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336;
  wire n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344;
  wire n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352;
  wire n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360;
  wire n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368;
  wire n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376;
  wire n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384;
  wire n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392;
  wire n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400;
  wire n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408;
  wire n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416;
  wire n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424;
  wire n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432;
  wire n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440;
  wire n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448;
  wire n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456;
  wire n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464;
  wire n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472;
  wire n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480;
  wire n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488;
  wire n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496;
  wire n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504;
  wire n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512;
  wire n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520;
  wire n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528;
  wire n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536;
  wire n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544;
  wire n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552;
  wire n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560;
  wire n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568;
  wire n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576;
  wire n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584;
  wire n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592;
  wire n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600;
  wire n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608;
  wire n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616;
  wire n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624;
  wire n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632;
  wire n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640;
  wire n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648;
  wire n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656;
  wire n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664;
  wire n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672;
  wire n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680;
  wire n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688;
  wire n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696;
  wire n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704;
  wire n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712;
  wire n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720;
  wire n32721, n32722, n32723, n32724, n32725, n32727, n32728, n32729;
  wire n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737;
  wire n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745;
  wire n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753;
  wire n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761;
  wire n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769;
  wire n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777;
  wire n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785;
  wire n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793;
  wire n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801;
  wire n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809;
  wire n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817;
  wire n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825;
  wire n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833;
  wire n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841;
  wire n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849;
  wire n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857;
  wire n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865;
  wire n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873;
  wire n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881;
  wire n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889;
  wire n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897;
  wire n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905;
  wire n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913;
  wire n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921;
  wire n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929;
  wire n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937;
  wire n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945;
  wire n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953;
  wire n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961;
  wire n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969;
  wire n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977;
  wire n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985;
  wire n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993;
  wire n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001;
  wire n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009;
  wire n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017;
  wire n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025;
  wire n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033;
  wire n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041;
  wire n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049;
  wire n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057;
  wire n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065;
  wire n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073;
  wire n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081;
  wire n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089;
  wire n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097;
  wire n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105;
  wire n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113;
  wire n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121;
  wire n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129;
  wire n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137;
  wire n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145;
  wire n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153;
  wire n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161;
  wire n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169;
  wire n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177;
  wire n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185;
  wire n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193;
  wire n33195, n33196, n33197, n33198, n33199, n33200, n33203, n33204;
  wire n33205, n33206, n33207, n33208, n33211, n33212, n33213, n33214;
  wire n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222;
  wire n33223, n33224, n33225, n33226, n33227, n33228, n33231, n33232;
  wire n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240;
  wire n33241, n33242, n33243, n33245, n33246, n33247, n33248, n33249;
  wire n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257;
  wire n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265;
  wire n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273;
  wire n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281;
  wire n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289;
  wire n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297;
  wire n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305;
  wire n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33314;
  wire n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322;
  wire n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330;
  wire n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338;
  wire n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346;
  wire n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354;
  wire n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362;
  wire n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370;
  wire n33371, n33372, n33373, n33375, n33376, n33377, n33378, n33379;
  wire n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387;
  wire n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395;
  wire n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403;
  wire n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411;
  wire n33412, n33413, n33416, n33417, n33418, n33419, n33420, n33421;
  wire n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429;
  wire n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437;
  wire n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445;
  wire n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453;
  wire n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461;
  wire n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469;
  wire n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477;
  wire n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485;
  wire n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493;
  wire n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501;
  wire n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509;
  wire n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517;
  wire n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525;
  wire n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533;
  wire n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541;
  wire n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549;
  wire n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557;
  wire n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565;
  wire n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573;
  wire n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581;
  wire n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589;
  wire n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597;
  wire n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605;
  wire n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613;
  wire n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621;
  wire n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629;
  wire n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637;
  wire n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645;
  wire n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653;
  wire n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661;
  wire n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669;
  wire n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677;
  wire n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685;
  wire n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693;
  wire n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701;
  wire n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709;
  wire n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717;
  wire n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725;
  wire n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733;
  wire n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741;
  wire n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749;
  wire n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757;
  wire n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33767;
  wire n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775;
  wire n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783;
  wire n33784, n33787, n33788, n33789, n33790, n33791, n33792, n33793;
  wire n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801;
  wire n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809;
  wire n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817;
  wire n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825;
  wire n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833;
  wire n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841;
  wire n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849;
  wire n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857;
  wire n33858, n33859, n33862, n33863, n33864, n33865, n33866, n33867;
  wire n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875;
  wire n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883;
  wire n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891;
  wire n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899;
  wire n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907;
  wire n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915;
  wire n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923;
  wire n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931;
  wire n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939;
  wire n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947;
  wire n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955;
  wire n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963;
  wire n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971;
  wire n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979;
  wire n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987;
  wire n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995;
  wire n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003;
  wire n34004, n34005, n34006, n34007, n34008, n34009, n34011, n34012;
  wire n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020;
  wire n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028;
  wire n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036;
  wire n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044;
  wire n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052;
  wire n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060;
  wire n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068;
  wire n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076;
  wire n34077, n34078, n34079, n34080, n34081, n34084, n34085, n34086;
  wire n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094;
  wire n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102;
  wire n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110;
  wire n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118;
  wire n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126;
  wire n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134;
  wire n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142;
  wire n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150;
  wire n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158;
  wire n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166;
  wire n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174;
  wire n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182;
  wire n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190;
  wire n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198;
  wire n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206;
  wire n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214;
  wire n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222;
  wire n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230;
  wire n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238;
  wire n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246;
  wire n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254;
  wire n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262;
  wire n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270;
  wire n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278;
  wire n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286;
  wire n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294;
  wire n34295, n34296, n34297, n34298, n34299, n34300, n34302, n34303;
  wire n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311;
  wire n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319;
  wire n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327;
  wire n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335;
  wire n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343;
  wire n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351;
  wire n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359;
  wire n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367;
  wire n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375;
  wire n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383;
  wire n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391;
  wire n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399;
  wire n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407;
  wire n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415;
  wire n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423;
  wire n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431;
  wire n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439;
  wire n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447;
  wire n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455;
  wire n34456, n34460, n34461, n34462, n34463, n34464, n34465, n34466;
  wire n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474;
  wire n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482;
  wire n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490;
  wire n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498;
  wire n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506;
  wire n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514;
  wire n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522;
  wire n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530;
  wire n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538;
  wire n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546;
  wire n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554;
  wire n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562;
  wire n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570;
  wire n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578;
  wire n34579, n34580, n34581, n34583, n34584, n34585, n34586, n34587;
  wire n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595;
  wire n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603;
  wire n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611;
  wire n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619;
  wire n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627;
  wire n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635;
  wire n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643;
  wire n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651;
  wire n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659;
  wire n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667;
  wire n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675;
  wire n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683;
  wire n34684, n34685, n34686, n34687, n34688, n34689, n34692, n34693;
  wire n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701;
  wire n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709;
  wire n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717;
  wire n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725;
  wire n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733;
  wire n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741;
  wire n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749;
  wire n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757;
  wire n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765;
  wire n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773;
  wire n34774, n34775, n34776, n34778, n34779, n34780, n34781, n34782;
  wire n34783, n34784, n34786, n34787, n34788, n34789, n34790, n34791;
  wire n34792, n34794, n34795, n34796, n34797, n34798, n34799, n34800;
  wire n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808;
  wire n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816;
  wire n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824;
  wire n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832;
  wire n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840;
  wire n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848;
  wire n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856;
  wire n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864;
  wire n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872;
  wire n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880;
  wire n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888;
  wire n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896;
  wire n34897, n34898, n34899, n34900, n34901, n34903, n34904, n34905;
  wire n34906, n34907, n34908, n34910, n34911, n34912, n34913, n34914;
  wire n34915, n34916, n34918, n34919, n34920, n34921, n34922, n34923;
  wire n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931;
  wire n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939;
  wire n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947;
  wire n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955;
  wire n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963;
  wire n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971;
  wire n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979;
  wire n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987;
  wire n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995;
  wire n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003;
  wire n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011;
  wire n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019;
  wire n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027;
  wire n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035;
  wire n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043;
  wire n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051;
  wire n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059;
  wire n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067;
  wire n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075;
  wire n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083;
  wire n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091;
  wire n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099;
  wire n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107;
  wire n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115;
  wire n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123;
  wire n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131;
  wire n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139;
  wire n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147;
  wire n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155;
  wire n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163;
  wire n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171;
  wire n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179;
  wire n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187;
  wire n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195;
  wire n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203;
  wire n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211;
  wire n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219;
  wire n35222, n35223, n35224, n35227, n35228, n35229, n35230, n35231;
  wire n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239;
  wire n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247;
  wire n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255;
  wire n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263;
  wire n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271;
  wire n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279;
  wire n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287;
  wire n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295;
  wire n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303;
  wire n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311;
  wire n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319;
  wire n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327;
  wire n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335;
  wire n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343;
  wire n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351;
  wire n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359;
  wire n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367;
  wire n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375;
  wire n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383;
  wire n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391;
  wire n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399;
  wire n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407;
  wire n35408, n35410, n35411, n35412, n35413, n35414, n35415, n35416;
  wire n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424;
  wire n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432;
  wire n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440;
  wire n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448;
  wire n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456;
  wire n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464;
  wire n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472;
  wire n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480;
  wire n35481, n35482, n35483, n35485, n35486, n35487, n35488, n35489;
  wire n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497;
  wire n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505;
  wire n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513;
  wire n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521;
  wire n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529;
  wire n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537;
  wire n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545;
  wire n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553;
  wire n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561;
  wire n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569;
  wire n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577;
  wire n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585;
  wire n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593;
  wire n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601;
  wire n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609;
  wire n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617;
  wire n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625;
  wire n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633;
  wire n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35643;
  wire n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652;
  wire n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660;
  wire n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668;
  wire n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676;
  wire n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684;
  wire n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692;
  wire n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700;
  wire n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708;
  wire n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716;
  wire n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724;
  wire n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732;
  wire n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740;
  wire n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748;
  wire n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756;
  wire n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764;
  wire n35765, n35766, n35767, n35768, n35769, n35771, n35772, n35773;
  wire n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781;
  wire n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789;
  wire n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35798;
  wire n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806;
  wire n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814;
  wire n35815, n35816, n35817, n35819, n35820, n35821, n35822, n35823;
  wire n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831;
  wire n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35840;
  wire n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848;
  wire n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856;
  wire n35857, n35858, n35859, n35861, n35862, n35863, n35864, n35865;
  wire n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873;
  wire n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881;
  wire n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889;
  wire n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897;
  wire n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905;
  wire n35906, n35909, n35910, n35911, n35912, n35913, n35914, n35915;
  wire n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923;
  wire n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931;
  wire n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939;
  wire n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947;
  wire n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955;
  wire n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963;
  wire n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971;
  wire n35972, n35973, n35974, n35975, n35977, n35978, n35979, n35980;
  wire n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988;
  wire n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996;
  wire n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004;
  wire n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012;
  wire n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020;
  wire n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028;
  wire n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036;
  wire n36037, n36038, n36039, n36042, n36043, n36044, n36045, n36046;
  wire n36047, n36048, n36049, n36052, n36053, n36054, n36055, n36056;
  wire n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064;
  wire n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072;
  wire n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082;
  wire n36083, n36084, n36085, n36086, n36088, n36089, n36090, n36091;
  wire n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099;
  wire n36100, n36101, n36102, n36103, n36104, n36105, n36107, n36108;
  wire n36109, n36110, n36111, n36112, n36114, n36115, n36116, n36117;
  wire n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125;
  wire n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133;
  wire n36135, n36136, n36137, n36138, n36139, n36140, n36142, n36143;
  wire n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151;
  wire n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159;
  wire n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167;
  wire n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175;
  wire n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183;
  wire n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191;
  wire n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199;
  wire n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207;
  wire n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215;
  wire n36216, n36219, n36220, n36221, n36222, n36223, n36224, n36225;
  wire n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233;
  wire n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243;
  wire n36244, n36245, n36246, n36247, n36248, n36249, n36251, n36252;
  wire n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260;
  wire n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268;
  wire n36269, n36272, n36273, n36274, n36275, n36278, n36279, n36280;
  wire n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288;
  wire n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296;
  wire n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304;
  wire n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312;
  wire n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320;
  wire n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328;
  wire n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336;
  wire n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344;
  wire n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352;
  wire n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360;
  wire n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368;
  wire n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376;
  wire n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384;
  wire n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392;
  wire n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400;
  wire n36401, n36402, n36403, n36404, n36405, n36406, n36409, n36410;
  wire n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418;
  wire n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426;
  wire n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434;
  wire n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442;
  wire n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450;
  wire n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458;
  wire n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466;
  wire n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474;
  wire n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482;
  wire n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490;
  wire n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498;
  wire n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506;
  wire n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514;
  wire n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522;
  wire n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530;
  wire n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538;
  wire n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546;
  wire n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554;
  wire n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562;
  wire n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570;
  wire n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578;
  wire n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586;
  wire n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594;
  wire n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602;
  wire n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610;
  wire n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618;
  wire n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626;
  wire n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634;
  wire n36635, n36636, n36637, n36638, n36639, n36642, n36643, n36644;
  wire n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652;
  wire n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660;
  wire n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668;
  wire n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676;
  wire n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684;
  wire n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692;
  wire n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700;
  wire n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708;
  wire n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716;
  wire n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724;
  wire n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732;
  wire n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740;
  wire n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748;
  wire n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756;
  wire n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764;
  wire n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772;
  wire n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780;
  wire n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788;
  wire n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796;
  wire n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804;
  wire n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812;
  wire n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820;
  wire n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828;
  wire n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836;
  wire n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844;
  wire n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852;
  wire n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860;
  wire n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868;
  wire n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36877;
  wire n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885;
  wire n36886, n36887, n36888, n36889, n36890, n36893, n36894, n36895;
  wire n36896, n36899, n36900, n36901, n36902, n36903, n36904, n36905;
  wire n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913;
  wire n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921;
  wire n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929;
  wire n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937;
  wire n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945;
  wire n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953;
  wire n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961;
  wire n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969;
  wire n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977;
  wire n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985;
  wire n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993;
  wire n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001;
  wire n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009;
  wire n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017;
  wire n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025;
  wire n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033;
  wire n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041;
  wire n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049;
  wire n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057;
  wire n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065;
  wire n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073;
  wire n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081;
  wire n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089;
  wire n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097;
  wire n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105;
  wire n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113;
  wire n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121;
  wire n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129;
  wire n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137;
  wire n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145;
  wire n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153;
  wire n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161;
  wire n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169;
  wire n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177;
  wire n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185;
  wire n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193;
  wire n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201;
  wire n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209;
  wire n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217;
  wire n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225;
  wire n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233;
  wire n37234, n37235, n37236, n37239, n37240, n37241, n37242, n37243;
  wire n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251;
  wire n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37261;
  wire n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269;
  wire n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277;
  wire n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37287;
  wire n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295;
  wire n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303;
  wire n37304, n37307, n37308, n37309, n37310, n37311, n37312, n37313;
  wire n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321;
  wire n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331;
  wire n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339;
  wire n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347;
  wire n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355;
  wire n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363;
  wire n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371;
  wire n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379;
  wire n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387;
  wire n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395;
  wire n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403;
  wire n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411;
  wire n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419;
  wire n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427;
  wire n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435;
  wire n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443;
  wire n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451;
  wire n37452, n37453, n37454, n37455, n37456, n37457, n37459, n37460;
  wire n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468;
  wire n37469, n37472, n37473, n37474, n37475, n37478, n37479, n37480;
  wire n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488;
  wire n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496;
  wire n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506;
  wire n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514;
  wire n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522;
  wire n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530;
  wire n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538;
  wire n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546;
  wire n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554;
  wire n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562;
  wire n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570;
  wire n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578;
  wire n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586;
  wire n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594;
  wire n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602;
  wire n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610;
  wire n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618;
  wire n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626;
  wire n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634;
  wire n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642;
  wire n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650;
  wire n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658;
  wire n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666;
  wire n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674;
  wire n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682;
  wire n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690;
  wire n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698;
  wire n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708;
  wire n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716;
  wire n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724;
  wire n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732;
  wire n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740;
  wire n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748;
  wire n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756;
  wire n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764;
  wire n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772;
  wire n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780;
  wire n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788;
  wire n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796;
  wire n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804;
  wire n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812;
  wire n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820;
  wire n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828;
  wire n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836;
  wire n37837, n37838, n37841, n37842, n37843, n37844, n37845, n37846;
  wire n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854;
  wire n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862;
  wire n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870;
  wire n37871, n37872, n37873, n37874, n37875, n37878, n37879, n37880;
  wire n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888;
  wire n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896;
  wire n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904;
  wire n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912;
  wire n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920;
  wire n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928;
  wire n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936;
  wire n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944;
  wire n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952;
  wire n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960;
  wire n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968;
  wire n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976;
  wire n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984;
  wire n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992;
  wire n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000;
  wire n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008;
  wire n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016;
  wire n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024;
  wire n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032;
  wire n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040;
  wire n38041, n38042, n38043, n38044, n38045, n38046, n38048, n38049;
  wire n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057;
  wire n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065;
  wire n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073;
  wire n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081;
  wire n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089;
  wire n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097;
  wire n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105;
  wire n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113;
  wire n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121;
  wire n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129;
  wire n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137;
  wire n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145;
  wire n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153;
  wire n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161;
  wire n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169;
  wire n38170, n38171, n38173, n38174, n38175, n38176, n38177, n38178;
  wire n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186;
  wire n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194;
  wire n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202;
  wire n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210;
  wire n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218;
  wire n38219, n38220, n38221, n38222, n38223, n38224, n38226, n38227;
  wire n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235;
  wire n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243;
  wire n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251;
  wire n38252, n38253, n38254, n38255, n38257, n38258, n38259, n38260;
  wire n38261, n38265, n38266, n38267, n38269, n38270, n38271, n38272;
  wire n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280;
  wire n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288;
  wire n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296;
  wire n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304;
  wire n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312;
  wire n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320;
  wire n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328;
  wire n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336;
  wire n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344;
  wire n38345, n38346, n38347, n38348, n38349, n38350, n38352, n38353;
  wire n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361;
  wire n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369;
  wire n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377;
  wire n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385;
  wire n38386, n38387, n38389, n38390, n38391, n38392, n38393, n38394;
  wire n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402;
  wire n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410;
  wire n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419;
  wire n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427;
  wire n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435;
  wire n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443;
  wire n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451;
  wire n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459;
  wire n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467;
  wire n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475;
  wire n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483;
  wire n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491;
  wire n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499;
  wire n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507;
  wire n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515;
  wire n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523;
  wire n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531;
  wire n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539;
  wire n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547;
  wire n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555;
  wire n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563;
  wire n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571;
  wire n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579;
  wire n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587;
  wire n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595;
  wire n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603;
  wire n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611;
  wire n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619;
  wire n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627;
  wire n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635;
  wire n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643;
  wire n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651;
  wire n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659;
  wire n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667;
  wire n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675;
  wire n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683;
  wire n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691;
  wire n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699;
  wire n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707;
  wire n38708, n38709, n38712, n38715, n38716, n38717, n38718, n38719;
  wire n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727;
  wire n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735;
  wire n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743;
  wire n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751;
  wire n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759;
  wire n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767;
  wire n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775;
  wire n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783;
  wire n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791;
  wire n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799;
  wire n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807;
  wire n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815;
  wire n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38824;
  wire n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832;
  wire n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840;
  wire n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848;
  wire n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856;
  wire n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864;
  wire n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872;
  wire n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880;
  wire n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888;
  wire n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896;
  wire n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904;
  wire n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912;
  wire n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920;
  wire n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928;
  wire n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936;
  wire n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944;
  wire n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952;
  wire n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960;
  wire n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968;
  wire n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976;
  wire n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984;
  wire n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992;
  wire n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000;
  wire n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008;
  wire n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016;
  wire n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024;
  wire n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032;
  wire n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040;
  wire n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048;
  wire n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056;
  wire n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064;
  wire n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072;
  wire n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080;
  wire n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088;
  wire n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096;
  wire n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104;
  wire n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112;
  wire n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120;
  wire n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128;
  wire n39129, n39130, n39131, n39132, n39133, n39136, n39137, n39138;
  wire n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146;
  wire n39147, n39148, n39149, n39150, n39153, n39154, n39155, n39156;
  wire n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165;
  wire n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175;
  wire n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183;
  wire n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191;
  wire n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199;
  wire n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207;
  wire n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215;
  wire n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223;
  wire n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231;
  wire n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239;
  wire n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247;
  wire n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255;
  wire n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263;
  wire n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271;
  wire n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279;
  wire n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287;
  wire n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295;
  wire n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303;
  wire n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311;
  wire n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319;
  wire n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327;
  wire n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335;
  wire n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343;
  wire n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351;
  wire n39352, n39353, n39354, n39356, n39357, n39358, n39359, n39360;
  wire n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39369;
  wire n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377;
  wire n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385;
  wire n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393;
  wire n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401;
  wire n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409;
  wire n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417;
  wire n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425;
  wire n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433;
  wire n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441;
  wire n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449;
  wire n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457;
  wire n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465;
  wire n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473;
  wire n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481;
  wire n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489;
  wire n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497;
  wire n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505;
  wire n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513;
  wire n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521;
  wire n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529;
  wire n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537;
  wire n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545;
  wire n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553;
  wire n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561;
  wire n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569;
  wire n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577;
  wire n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585;
  wire n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593;
  wire n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601;
  wire n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609;
  wire n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617;
  wire n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625;
  wire n39626, n39627, n39628, n39629, n39631, n39632, n39633, n39634;
  wire n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642;
  wire n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650;
  wire n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658;
  wire n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666;
  wire n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674;
  wire n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682;
  wire n39683, n39684, n39685, n39686, n39687, n39688, n39691, n39692;
  wire n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700;
  wire n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708;
  wire n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716;
  wire n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724;
  wire n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732;
  wire n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740;
  wire n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748;
  wire n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756;
  wire n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764;
  wire n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774;
  wire n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782;
  wire n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790;
  wire n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798;
  wire n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806;
  wire n39807, n39808, n39809, n39810, n39811, n39812, n39815, n39816;
  wire n39817, n39820, n39821, n39822, n39823, n39824, n39825, n39826;
  wire n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834;
  wire n39835, n39836, n39839, n39840, n39841, n39842, n39843, n39844;
  wire n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852;
  wire n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860;
  wire n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868;
  wire n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876;
  wire n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884;
  wire n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892;
  wire n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39902;
  wire n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910;
  wire n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918;
  wire n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926;
  wire n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934;
  wire n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942;
  wire n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950;
  wire n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958;
  wire n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966;
  wire n39967, n39969, n39970, n39971, n39972, n39973, n39974, n39975;
  wire n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983;
  wire n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991;
  wire n39992, n39993, n39994, n39997, n39998, n39999, n40000, n40001;
  wire n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009;
  wire n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017;
  wire n40018, n40019, n40020, n40021, n40024, n40027, n40028, n40029;
  wire n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037;
  wire n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045;
  wire n40046, n40047, n40048, n40049, n40050, n40051, n40052, n40053;
  wire n40054, n40055, n40056, n40057, n40058, n40060, n40061, n40062;
  wire n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070;
  wire n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078;
  wire n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086;
  wire n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094;
  wire n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102;
  wire n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110;
  wire n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118;
  wire n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126;
  wire n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134;
  wire n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142;
  wire n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150;
  wire n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158;
  wire n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166;
  wire n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174;
  wire n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182;
  wire n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190;
  wire n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198;
  wire n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206;
  wire n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214;
  wire n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222;
  wire n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230;
  wire n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238;
  wire n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246;
  wire n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254;
  wire n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262;
  wire n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270;
  wire n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278;
  wire n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286;
  wire n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294;
  wire n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302;
  wire n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310;
  wire n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318;
  wire n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326;
  wire n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334;
  wire n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342;
  wire n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350;
  wire n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358;
  wire n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366;
  wire n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374;
  wire n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382;
  wire n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390;
  wire n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398;
  wire n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406;
  wire n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414;
  wire n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422;
  wire n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430;
  wire n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438;
  wire n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446;
  wire n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454;
  wire n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462;
  wire n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470;
  wire n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478;
  wire n40479, n40481, n40482, n40483, n40484, n40485, n40486, n40487;
  wire n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495;
  wire n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503;
  wire n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511;
  wire n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519;
  wire n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527;
  wire n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535;
  wire n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543;
  wire n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551;
  wire n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559;
  wire n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567;
  wire n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575;
  wire n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583;
  wire n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591;
  wire n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599;
  wire n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607;
  wire n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615;
  wire n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623;
  wire n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631;
  wire n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639;
  wire n40640, n40641, n40642, n40645, n40646, n40647, n40648, n40649;
  wire n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657;
  wire n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665;
  wire n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673;
  wire n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681;
  wire n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689;
  wire n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697;
  wire n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705;
  wire n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713;
  wire n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721;
  wire n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729;
  wire n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737;
  wire n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745;
  wire n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753;
  wire n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761;
  wire n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40770;
  wire n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778;
  wire n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786;
  wire n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794;
  wire n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802;
  wire n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810;
  wire n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818;
  wire n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826;
  wire n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834;
  wire n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842;
  wire n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850;
  wire n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40859;
  wire n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867;
  wire n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875;
  wire n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883;
  wire n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891;
  wire n40892, n40893, n40896, n40897, n40898, n40899, n40900, n40901;
  wire n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909;
  wire n40910, n40911, n40912, n40913, n40914, n40915, n40916, n40917;
  wire n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925;
  wire n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933;
  wire n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941;
  wire n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949;
  wire n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957;
  wire n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965;
  wire n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973;
  wire n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983;
  wire n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991;
  wire n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999;
  wire n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007;
  wire n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015;
  wire n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023;
  wire n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031;
  wire n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039;
  wire n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047;
  wire n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055;
  wire n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063;
  wire n41064, n41067, n41068, n41069, n41070, n41071, n41072, n41073;
  wire n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081;
  wire n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089;
  wire n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097;
  wire n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105;
  wire n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113;
  wire n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121;
  wire n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129;
  wire n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137;
  wire n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145;
  wire n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153;
  wire n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161;
  wire n41162, n41163, n41166, n41167, n41168, n41170, n41171, n41172;
  wire n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180;
  wire n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188;
  wire n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41198;
  wire n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208;
  wire n41209, n41212, n41213, n41214, n41215, n41216, n41217, n41218;
  wire n41219, n41220, n41221, n41223, n41224, n41225, n41226, n41227;
  wire n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235;
  wire n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243;
  wire n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251;
  wire n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259;
  wire n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267;
  wire n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275;
  wire n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283;
  wire n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291;
  wire n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299;
  wire n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307;
  wire n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315;
  wire n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323;
  wire n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331;
  wire n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339;
  wire n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347;
  wire n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355;
  wire n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363;
  wire n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371;
  wire n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379;
  wire n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387;
  wire n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395;
  wire n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403;
  wire n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411;
  wire n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419;
  wire n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427;
  wire n41428, n41429, n41432, n41433, n41434, n41435, n41436, n41437;
  wire n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445;
  wire n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453;
  wire n41454, n41455, n41456, n41457, n41458, n41461, n41462, n41463;
  wire n41464, n41465, n41466, n41467, n41468, n41470, n41471, n41472;
  wire n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480;
  wire n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488;
  wire n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496;
  wire n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504;
  wire n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512;
  wire n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520;
  wire n41521, n41522, n41523, n41524, n41525, n41526, n41530, n41531;
  wire n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539;
  wire n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547;
  wire n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555;
  wire n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563;
  wire n41564, n41565, n41566, n41567, n41568, n41571, n41572, n41573;
  wire n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581;
  wire n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589;
  wire n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597;
  wire n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605;
  wire n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613;
  wire n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621;
  wire n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629;
  wire n41630, n41631, n41632, n41635, n41636, n41637, n41638, n41639;
  wire n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647;
  wire n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655;
  wire n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663;
  wire n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671;
  wire n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679;
  wire n41680, n41681, n41682, n41683, n41686, n41687, n41688, n41689;
  wire n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697;
  wire n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707;
  wire n41710, n41711, n41712, n41713, n41717, n41718, n41719, n41720;
  wire n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728;
  wire n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738;
  wire n41739, n41740, n41741, n41742, n41744, n41745, n41746, n41747;
  wire n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755;
  wire n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763;
  wire n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771;
  wire n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779;
  wire n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787;
  wire n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795;
  wire n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803;
  wire n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811;
  wire n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819;
  wire n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827;
  wire n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835;
  wire n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843;
  wire n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851;
  wire n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859;
  wire n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867;
  wire n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875;
  wire n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883;
  wire n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891;
  wire n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899;
  wire n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907;
  wire n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915;
  wire n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923;
  wire n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931;
  wire n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939;
  wire n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947;
  wire n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955;
  wire n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963;
  wire n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971;
  wire n41972, n41974, n41975, n41976, n41977, n41978, n41979, n41980;
  wire n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988;
  wire n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996;
  wire n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004;
  wire n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012;
  wire n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020;
  wire n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028;
  wire n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036;
  wire n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044;
  wire n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052;
  wire n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060;
  wire n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068;
  wire n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076;
  wire n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084;
  wire n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092;
  wire n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100;
  wire n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108;
  wire n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116;
  wire n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124;
  wire n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132;
  wire n42133, n42134, n42135, n42137, n42138, n42139, n42140, n42141;
  wire n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149;
  wire n42150, n42151, n42152, n42155, n42156, n42157, n42158, n42159;
  wire n42160, n42161, n42162, n42163, n42164, n42165, n42166, n42167;
  wire n42168, n42171, n42172, n42173, n42174, n42175, n42176, n42177;
  wire n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185;
  wire n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193;
  wire n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42203;
  wire n42204, n42205, n42206, n42207, n42208, n42209, n42212, n42213;
  wire n42214, n42215, n42216, n42217, n42218, n42219, n42220, n42221;
  wire n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229;
  wire n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237;
  wire n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245;
  wire n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253;
  wire n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261;
  wire n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269;
  wire n42270, n42271, n42272, n42273, n42274, n42275, n42276, n42277;
  wire n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285;
  wire n42286, n42287, n42288, n42289, n42290, n42291, n42292, n42293;
  wire n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301;
  wire n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309;
  wire n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317;
  wire n42318, n42319, n42320, n42321, n42322, n42323, n42325, n42326;
  wire n42327, n42328, n42329, n42333, n42334, n42335, n42336, n42337;
  wire n42338, n42339, n42340, n42341, n42343, n42344, n42345, n42346;
  wire n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354;
  wire n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362;
  wire n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370;
  wire n42371, n42372, n42373, n42378, n42379, n42380, n42381, n42382;
  wire n42383, n42385, n42386, n42387, n42388, n42389, n42390, n42391;
  wire n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399;
  wire n42400, n42401, n42402, n42403, n42404, n42407, n42408, n42409;
  wire n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417;
  wire n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425;
  wire n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433;
  wire n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441;
  wire n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449;
  wire n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459;
  wire n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467;
  wire n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475;
  wire n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483;
  wire n42484, n42485, n42486, n42487, n42488, n42489, n42492, n42493;
  wire n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501;
  wire n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509;
  wire n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517;
  wire n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525;
  wire n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533;
  wire n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541;
  wire n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42549;
  wire n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557;
  wire n42558, n42559, n42560, n42561, n42562, n42563, n42564, n42565;
  wire n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573;
  wire n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581;
  wire n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589;
  wire n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597;
  wire n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605;
  wire n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613;
  wire n42614, n42615, n42616, n42617, n42618, n42619, n42621, n42622;
  wire n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630;
  wire n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638;
  wire n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646;
  wire n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654;
  wire n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662;
  wire n42663, n42664, n42667, n42668, n42669, n42670, n42671, n42672;
  wire n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680;
  wire n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688;
  wire n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696;
  wire n42697, n42698, n42699, n42700, n42703, n42704, n42705, n42706;
  wire n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714;
  wire n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722;
  wire n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730;
  wire n42731, n42732, n42733, n42734, n42735, n42738, n42739, n42742;
  wire n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750;
  wire n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758;
  wire n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766;
  wire n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774;
  wire n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782;
  wire n42783, n42784, n42787, n42788, n42789, n42790, n42791, n42792;
  wire n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800;
  wire n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808;
  wire n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816;
  wire n42817, n42818, n42821, n42822, n42823, n42824, n42825, n42826;
  wire n42827, n42828, n42829, n42830, n42833, n42834, n42835, n42836;
  wire n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844;
  wire n42845, n42847, n42848, n42849, n42850, n42851, n42853, n42854;
  wire n42855, n42856, n42857, n42859, n42860, n42861, n42862, n42863;
  wire n42865, n42866, n42867, n42868, n42869, n42871, n42872, n42873;
  wire n42874, n42875, n42877, n42878, n42879, n42880, n42881, n42882;
  wire n42884, n42885, n42886, n42887, n42888, n42889, n42891, n42892;
  wire n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900;
  wire n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908;
  wire n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916;
  wire n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42925;
  wire n42926, n42927, n42928, n42929, n42930, n42931, n42932, n42933;
  wire n42934, n42935, n42936, n42939, n42942, n42943, n42944, n42945;
  wire n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953;
  wire n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961;
  wire n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969;
  wire n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977;
  wire n42978, n42979, n42980, n42981, n42984, n42985, n42986, n42987;
  wire n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995;
  wire n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003;
  wire n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011;
  wire n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019;
  wire n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027;
  wire n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035;
  wire n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043;
  wire n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051;
  wire n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059;
  wire n43060, n43061, n43062, n43065, n43066, n43067, n43068, n43069;
  wire n43070, n43071, n43072, n43073, n43074, n43075, n43076, n43077;
  wire n43078, n43079, n43080, n43083, n43084, n43085, n43086, n43087;
  wire n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095;
  wire n43096, n43097, n43098, n43099, n43100, n43101, n43102, n43103;
  wire n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111;
  wire n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119;
  wire n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127;
  wire n43128, n43129, n43130, n43131, n43132, n43133, n43135, n43136;
  wire n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144;
  wire n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152;
  wire n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160;
  wire n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168;
  wire n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176;
  wire n43177, n43178, n43180, n43181, n43182, n43183, n43184, n43185;
  wire n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193;
  wire n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201;
  wire n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209;
  wire n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217;
  wire n43218, n43219, n43221, n43222, n43223, n43224, n43225, n43226;
  wire n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234;
  wire n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242;
  wire n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250;
  wire n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258;
  wire n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266;
  wire n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274;
  wire n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282;
  wire n43283, n43284, n43285, n43286, n43288, n43289, n43290, n43291;
  wire n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299;
  wire n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307;
  wire n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315;
  wire n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323;
  wire n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331;
  wire n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339;
  wire n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347;
  wire n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355;
  wire n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363;
  wire n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371;
  wire n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379;
  wire n43380, n43383, n43384, n43385, n43386, n43389, n43390, n43391;
  wire n43392, n43395, n43396, n43397, n43398, n43399, n43400, n43401;
  wire n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409;
  wire n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417;
  wire n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425;
  wire n43426, n43427, n43428, n43429, n43430, n43433, n43434, n43435;
  wire n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443;
  wire n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451;
  wire n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459;
  wire n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467;
  wire n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475;
  wire n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483;
  wire n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491;
  wire n43492, n43493, n43495, n43496, n43497, n43498, n43499, n43500;
  wire n43501, n43502, n43503, n43504, n43505, n43506, n43507, n43508;
  wire n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516;
  wire n43517, n43520, n43521, n43522, n43523, n43524, n43525, n43526;
  wire n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534;
  wire n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542;
  wire n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550;
  wire n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558;
  wire n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566;
  wire n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574;
  wire n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582;
  wire n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590;
  wire n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598;
  wire n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606;
  wire n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614;
  wire n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622;
  wire n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630;
  wire n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638;
  wire n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646;
  wire n43647, n43648, n43649, n43650, n43652, n43653, n43654, n43655;
  wire n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663;
  wire n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671;
  wire n43672, n43673, n43674, n43675, n43676, n43677, n43678, n43679;
  wire n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687;
  wire n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695;
  wire n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704;
  wire n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712;
  wire n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720;
  wire n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728;
  wire n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736;
  wire n43737, n43738, n43739, n43741, n43742, n43743, n43744, n43745;
  wire n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753;
  wire n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761;
  wire n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769;
  wire n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777;
  wire n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785;
  wire n43786, n43787, n43788, n43790, n43791, n43792, n43793, n43794;
  wire n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802;
  wire n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810;
  wire n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818;
  wire n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826;
  wire n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834;
  wire n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842;
  wire n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850;
  wire n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858;
  wire n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866;
  wire n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874;
  wire n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882;
  wire n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43891;
  wire n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899;
  wire n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907;
  wire n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915;
  wire n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923;
  wire n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931;
  wire n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939;
  wire n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947;
  wire n43948, n43949, n43950, n43951, n43952, n43954, n43955, n43956;
  wire n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964;
  wire n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972;
  wire n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980;
  wire n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988;
  wire n43989, n43990, n43991, n43992, n43993, n43995, n43996, n43997;
  wire n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005;
  wire n44006, n44007, n44008, n44009, n44010, n44011, n44012, n44013;
  wire n44014, n44015, n44016, n44017, n44018, n44019, n44020, n44021;
  wire n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029;
  wire n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037;
  wire n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045;
  wire n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053;
  wire n44054, n44055, n44056, n44057, n44058, n44059, n44060, n44061;
  wire n44062, n44063, n44064, n44065, n44066, n44067, n44069, n44070;
  wire n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078;
  wire n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086;
  wire n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094;
  wire n44095, n44096, n44098, n44099, n44100, n44101, n44102, n44103;
  wire n44104, n44105, n44106, n44107, n44108, n44109, n44110, n44111;
  wire n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119;
  wire n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127;
  wire n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135;
  wire n44136, n44137, n44138, n44139, n44141, n44142, n44143, n44144;
  wire n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152;
  wire n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160;
  wire n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168;
  wire n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176;
  wire n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184;
  wire n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192;
  wire n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200;
  wire n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208;
  wire n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217;
  wire n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225;
  wire n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233;
  wire n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241;
  wire n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249;
  wire n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257;
  wire n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265;
  wire n44266, n44267, n44269, n44270, n44271, n44272, n44273, n44274;
  wire n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282;
  wire n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290;
  wire n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298;
  wire n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306;
  wire n44307, n44308, n44309, n44310, n44311, n44313, n44314, n44315;
  wire n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323;
  wire n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331;
  wire n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339;
  wire n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347;
  wire n44348, n44349, n44350, n44352, n44353, n44354, n44355, n44356;
  wire n44357, n44358, n44359, n44360, n44361, n44362, n44363, n44364;
  wire n44365, n44366, n44367, n44368, n44369, n44370, n44371, n44372;
  wire n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380;
  wire n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388;
  wire n44389, n44391, n44392, n44393, n44394, n44395, n44396, n44397;
  wire n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405;
  wire n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413;
  wire n44414, n44415, n44416, n44417, n44418, n44419, n44420, n44421;
  wire n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429;
  wire n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437;
  wire n44438, n44439, n44440, n44441, n44442, n44443, n44444, n44445;
  wire n44446, n44447, n44448, n44450, n44451, n44452, n44454, n44455;
  wire n44456, n44457, n44458, n44459, n44460, n44461, n44462, n44463;
  wire n44464, n44465, n44466, n44467, n44468, n44469, n44470, n44472;
  wire n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480;
  wire n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488;
  wire n44490, n44492, n44493, n44495, n44496, n44497, n44499, n44500;
  wire n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508;
  wire n44509, n44510, n44511, n44512, n44514, n44515, n44517, n44518;
  wire n44520, n44521, n44523, n44524, n44526, n44527, n44529, n44530;
  wire n44532, n44533, n44535, n44536, n44538, n44539, n44541, n44542;
  wire n44543, n44544, n44545, n44546, n44547, n44549, n44550, n44551;
  wire n44552, n44553, n44554, n44556, n44557, n44558, n44560, n44561;
  wire n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569;
  wire n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577;
  wire n44578, n44582, n44583, n44585, n44586, n44588, n44589, n44591;
  wire n44592, n44594, n44595, n44597, n44598, n44600, n44601, n44603;
  wire n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611;
  wire n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619;
  wire n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44630;
  wire n44631, n44632, n44634, n44635, n44637, n44638, n44639, n44641;
  wire n44642, n44644, n44645, n44646, n44647, n44648, n44649, n44650;
  wire n44651, n44652, n44653, n44654, n44656, n44657, n44658, n44659;
  wire n44661, n44662, n44664, n44665, n44666, n44668, n44669, n44670;
  wire n44671, n44673, n44674, n44676, n44677, n44679, n44680, n44682;
  wire n44683, n44685, n44686, n44688, n44689, n44691, n44692, n44694;
  wire n44695, n44697, n44698, n44700, n44701, n44703, n44704, n44706;
  wire n44707, n44708, n44709, n44710, n44711, n44712, n44714, n44715;
  wire n44716, n44717, n44719, n44720, n44721, n44722, n44723, n44724;
  wire n44725, n44726, n44727, n44728, n44729, n44731, n44732, n44734;
  wire n44735, n44737, n44738, n44740, n44741, n44743, n44744, n44746;
  wire n44747, n44749, n44750, n44752, n44753, n44754, n44755, n44756;
  wire n44758, n44759, n44761, n44762, n44764, n44765, n44767, n44768;
  wire n44770, n44771, n44773, n44774, n44776, n44777, n44779, n44780;
  wire n44782, n44783, n44785, n44786, n44788, n44789, n44791, n44792;
  wire n44794, n44795, n44797, n44798, n44800, n44801, n44803, n44804;
  wire n44806, n44807, n44809, n44810, n44812, n44813, n44815, n44816;
  wire n44818, n44819, n44821, n44822, n44824, n44825, n44827, n44828;
  wire n44830, n44831, n44833, n44834, n44836, n44837, n44839, n44840;
  wire n44842, n44843, n44845, n44846, n44848, n44849, n44851, n44852;
  wire n44854, n44855, n44857, n44858, n44860, n44861, n44863, n44864;
  wire n44866, n44867, n44869, n44870, n44872, n44873, n44875, n44876;
  wire n44878, n44879, n44881, n44882, n44884, n44885, n44887, n44888;
  wire n44890, n44891, n44893, n44894, n44896, n44897, n44899, n44900;
  wire n44902, n44903, n44905, n44906, n44908, n44909, n44911, n44912;
  wire n44914, n44915, n44917, n44918, n44920, n44921, n44923, n44924;
  wire n44926, n44927, n44929, n44930, n44932, n44933, n44935, n44936;
  wire n44938, n44939, n44941, n44942, n44944, n44945, n44947, n44948;
  wire n44950, n44951, n44953, n44954, n44956, n44957, n44959, n44960;
  wire n44962, n44963, n44965, n44966, n44968, n44969, n44971, n44972;
  wire n44974, n44975, n44977, n44978, n44979, n44981, n44982, n44984;
  wire n44985, n44987, n44988, n44990, n44991, n44993, n44994, n44996;
  wire n44997, n44999, n45000, n45002, n45003, n45005, n45006, n45008;
  wire n45009, n45011, n45012, n45014, n45015, n45017, n45018, n45020;
  wire n45021, n45023, n45024, n45026, n45027, n45029, n45030, n45032;
  wire n45033, n45035, n45036, n45038, n45039, n45041, n45042, n45044;
  wire n45045, n45047, n45048, n45050, n45051, n45053, n45054, n45056;
  wire n45057, n45059, n45060, n45062, n45063, n45065, n45066, n45068;
  wire n45069, n45071, n45072, n45074, n45075, n45077, n45078, n45080;
  wire n45081, n45083, n45084, n45086, n45087, n45089, n45090, n45092;
  wire n45093, n45095, n45096, n45098, n45099, n45101, n45102, n45104;
  wire n45105, n45107, n45108, n45109, n45110, n45111, n45112, n45113;
  wire n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121;
  wire n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129;
  wire n45131, n45132, n45134, n45135, n45137, n45138, n45140, n45141;
  wire n45143, n45144, n45146, n45147, n45149, n45150, n45152, n45153;
  wire n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161;
  wire n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169;
  wire n45170, n45171, n45172, n45175, n45177, n45178, n45179, n45180;
  wire n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188;
  wire n45189, n45190, n45191, n45195, n45196, n45197, n45198, n45199;
  wire n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210;
  wire n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218;
  wire n45219, n45220, n45221, n45222, n45223, n45225, n45228, n45229;
  wire n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238;
  wire n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246;
  wire n45249, n45251, n45252, n45253, n45254, n45255, n45256, n45257;
  wire n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265;
  wire n45266, n45269, n45271, n45272, n45273, n45274, n45275, n45276;
  wire n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284;
  wire n45285, n45286, n45289, n45291, n45292, n45293, n45294, n45295;
  wire n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303;
  wire n45304, n45305, n45306, n45309, n45311, n45312, n45313, n45314;
  wire n45315, n45316, n45317, n45318, n45322, n45323, n45324, n45325;
  wire n45326, n45327, n45328, n45329, n45333, n45334, n45335, n45336;
  wire n45337, n45338, n45339, n45340, n45344, n45345, n45346, n45347;
  wire n45348, n45349, n45352, n45353, n45354, n45357, n45358, n45360;
  wire n45361, n45363, n45364, n45366, n45367, n45369, n45370, n45372;
  wire n45373, n45375, n45376, n45378, n45379, n45381, n45382, n45384;
  wire n45385, n45387, n45388, n45390, n45391, n45393, n45394, n45396;
  wire n45397, n45399, n45400, n45402, n45403, n45405, n45406, n45408;
  wire n45409, n45411, n45412, n45414, n45415, n45417, n45418, n45420;
  wire n45421, n45423, n45424, n45426, n45427, n45429, n45430, n45431;
  wire n45432, n45433, n45434, n45435, n45436, n45438, n45439, n45441;
  wire n45442, n45444, n45445, n45447, n45448, n45450, n45451, n45453;
  wire n45454, n45455, n45456, n45457, n45459, n45460, n45462, n45463;
  wire n45465, n45466, n45468, n45469, n45471, n45472, n45474, n45475;
  wire n45477, n45478, n45479, n45480, n45481, n45483, n45484, n45486;
  wire n45487, n45489, n45490, n45492, n45493, n45495, n45496, n45497;
  wire n45498, n45500, n45501, n45503, n45504, n45506, n45507, n45509;
  wire n45510, n45512, n45513, n45515, n45516, n45518, n45519, n45521;
  wire n45522, n45524, n45525, n45527, n45528, n45530, n45531, n45533;
  wire n45534, n45536, n45537, n45539, n45540, n45542, n45543, n45545;
  wire n45546, n45548, n45549, n45551, n45552, n45554, n45555, n45557;
  wire n45558, n45560, n45561, n45562, n45563, n45565, n45566, n45568;
  wire n45569, n45571, n45572, n45574, n45575, n45577, n45578, n45580;
  wire n45581, n45583, n45584, n45586, n45587, n45589, n45590, n45592;
  wire n45593, n45595, n45596, n45598, n45599, n45601, n45602, n45603;
  wire n45604, n45606, n45607, n45609, n45610, n45612, n45613, n45615;
  wire n45616, n45618, n45619, n45621, n45622, n45624, n45625, n45627;
  wire n45628, n45630, n45631, n45633, n45634, n45638, n45639, n45640;
  wire n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648;
  wire n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656;
  wire n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664;
  wire n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672;
  wire n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680;
  wire n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688;
  wire n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696;
  wire n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704;
  wire n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712;
  wire n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720;
  wire n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728;
  wire n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736;
  wire n45737, n45738, n45739, n45740, n45741, n45742, n45744, n45745;
  wire n45747, n45748, n45750, n45751, n45752, n45753, n45755, n45756;
  wire n45758, n45759, n45761, n45762, n45764, n45765, n45767, n45768;
  wire n45770, n45771, n45773, n45774, n45776, n45777, n45779, n45780;
  wire n45782, n45783, n45785, n45786, n45788, n45789, n45791, n45792;
  wire n45794, n45795, n45797, n45798, n45800, n45805, n45807, n45808;
  wire n45809, n45810, n45812, n45813, n45814, n45815, n45816, n45817;
  wire n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825;
  wire n45826, n45827, n45828, n45829, n45830, n45831, n45833, n45834;
  wire n45835, n45837, n45838, n45839, n45841, n45842, n45843, n45845;
  wire n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853;
  wire n45854, n45855, n45856, n45864, n45865, n45866, n45867, n45868;
  wire n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876;
  wire n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884;
  wire n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892;
  wire n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900;
  wire n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908;
  wire n45909, n45910, n45915, n45916, n45917, n45918, n45919, n45920;
  wire n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928;
  wire n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936;
  wire n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944;
  wire n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952;
  wire n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960;
  wire n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968;
  wire n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976;
  wire n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984;
  wire n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992;
  wire n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000;
  wire n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008;
  wire n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016;
  wire n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024;
  wire n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032;
  wire n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040;
  wire n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048;
  wire n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056;
  wire n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064;
  wire n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072;
  wire n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080;
  wire n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088;
  wire n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096;
  wire n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104;
  wire n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112;
  wire n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120;
  wire n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128;
  wire n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136;
  wire n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144;
  wire n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152;
  wire n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160;
  wire n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168;
  wire n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176;
  wire n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184;
  wire n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192;
  wire n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200;
  wire n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208;
  wire n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216;
  wire n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224;
  wire n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232;
  wire n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240;
  wire n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248;
  wire n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256;
  wire n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264;
  wire n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272;
  wire n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280;
  wire n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288;
  wire n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296;
  wire n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304;
  wire n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312;
  wire n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320;
  wire n46321, n46322, n46323, n46327, n46328, n46329, n46330, n46331;
  wire n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339;
  wire n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347;
  wire n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355;
  wire n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363;
  wire n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46374;
  wire n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382;
  wire n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390;
  wire n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398;
  wire n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406;
  wire n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414;
  wire n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422;
  wire n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430;
  wire n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438;
  wire n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446;
  wire n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454;
  wire n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462;
  wire n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470;
  wire n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478;
  wire n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486;
  wire n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494;
  wire n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502;
  wire n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510;
  wire n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518;
  wire n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526;
  wire n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534;
  wire n46535, n46536, n46537, n46538, n46539, n46549, n46550, n46551;
  wire n46552, n46553, n46554, n46555, n46556, n46557, n46558, n46559;
  wire n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567;
  wire n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575;
  wire n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583;
  wire n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591;
  wire n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46605;
  wire n46606, n46609, n46610, n46611, n46612, n46613, n46614, n46615;
  wire n46616, n46617, n46618, n46619, n46620, n46621, n46622, n46623;
  wire n46624, n46625, n46626, n46627, n46628, n46629, n46630, n46631;
  wire n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639;
  wire n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647;
  wire n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655;
  wire n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663;
  wire n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671;
  wire n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679;
  wire n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687;
  wire n46688, n46689, n46690, n46691, n46692, n46693, n46694, n46695;
  wire n46696, n46697, n46698, n46699, n46700, n46701, n46702, n46703;
  wire n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711;
  wire n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719;
  wire n46720, n46721, n46722, n46724, n46725, n46726, n46727, n46728;
  wire n46729, n46731, n46732, n46733, n46734, n46735, n46737, n46738;
  wire n46739, n46740, n46741, n46743, n46744, n46745, n46747, n46748;
  wire n46749, n46750, n46751, n46753, n46754, n46755, n46757, n46758;
  wire n46760, n46761, n46762, n46764, n46765, n46766, n46767, n46768;
  wire n46774, n46776, n46777, n46778, n46779, n46780, n46781, n46782;
  wire n46783, n46785, n46786, n46787, n46788, n46790, n46791, n46792;
  wire n46793, n46794, n46795, n46797, n46798, n46800, n46801, n46802;
  wire n46803, n46804, n46806, n46807, n46808, n46810, n46811, n46812;
  wire n46814, n46815, n46816, n46818, n46819, n46820, n46822, n46823;
  wire n46824, n46826, n46827, n46828, n46830, n46831, n46832, n46834;
  wire n46835, n46836, n46837, n46839, n46840, n46841, n46842, n46844;
  wire n46845, n46846, n46847, n46849, n46850, n46851, n46852, n46853;
  wire n46855, n46856, n46857, n46859, n46860, n46861, n46863, n46864;
  wire n46865, n46867, n46868, n46869, n46871, n46872, n46873, n46875;
  wire n46876, n46877, n46879, n46880, n46881, n46882, n46883, n46888;
  wire n46890, n46891, n46892, n46894, n46895, n46896, n46898, n46899;
  wire n46900, n46902, n46903, n46904, n46906, n46907, n46908, n46910;
  wire n46911, n46912, n46914, n46915, n46916, n46918, n46919, n46920;
  wire n46922, n46923, n46924, n46926, n46927, n46928, n46930, n46931;
  wire n46932, n46934, n46935, n46936, n46938, n46939, n46940, n46942;
  wire n46943, n46944, n46946, n46947, n46948, n46950, n46951, n46952;
  wire n46954, n46955, n46956, n46958, n46959, n46960, n46962, n46963;
  wire n46964, n46966, n46967, n46968, n46970, n46971, n46972, n46974;
  wire n46975, n46976, n46978, n46979, n46980, n46982, n46983, n46984;
  wire n46986, n46987, n46988, n46990, n46991, n46992, n46994, n46995;
  wire n46996, n46998, n46999, n47000, n47002, n47003, n47004, n47006;
  wire n47007, n47008, n47010, n47011, n47012, n47014, n47015, n47016;
  wire n47018, n47019, n47020, n47022, n47023, n47024, n47026, n47027;
  wire n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47036;
  wire n47038, n47039, n47040, n47042, n47043, n47044, n47046, n47047;
  wire n47048, n47050, n47051, n47052, n47053, n47054, n47055, n47056;
  wire n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064;
  wire n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072;
  wire n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080;
  wire n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088;
  wire n47089, n47090, n47091, n47092, n47095, n47096, n47097, n47099;
  wire n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107;
  wire n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115;
  wire n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123;
  wire n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131;
  wire n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139;
  wire n47141, n47142, n47143, n47145, n47146, n47147, n47148, n47149;
  wire n47150, n47151, n47152, n47153, n47154, n47155, n47156, n47157;
  wire n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167;
  wire n47168, n47169, n47170, n47171, n47172, n47173, n47174, n47175;
  wire n47176, n47177, n47178, n47179, n47181, n47182, n47183, n47184;
  wire n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192;
  wire n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200;
  wire n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208;
  wire n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216;
  wire n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225;
  wire n47226, n47227, n47228, n47229, n47230, n47233, n47234, n47235;
  wire n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243;
  wire n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251;
  wire n47252, n47254, n47255, n47256, n47258, n47259, n47260, n47261;
  wire n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269;
  wire n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277;
  wire n47278, n47281, n47282, n47283, n47284, n47287, n47288, n47289;
  wire n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298;
  wire n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306;
  wire n47307, n47308, n47309, n47310, n47311, n47314, n47315, n47316;
  wire n47319, n47320, n47321, n47323, n47324, n47325, n47326, n47327;
  wire n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335;
  wire n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345;
  wire n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353;
  wire n47354, n47355, n47356, n47357, n47359, n47360, n47361, n47362;
  wire n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370;
  wire n47371, n47374, n47375, n47376, n47377, n47378, n47379, n47380;
  wire n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388;
  wire n47389, n47390, n47391, n47392, n47393, n47395, n47396, n47397;
  wire n47398, n47399, n47400, n47401, n47402, n47403, n47404, n47405;
  wire n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413;
  wire n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421;
  wire n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429;
  wire n47430, n47431, n47433, n47434, n47435, n47436, n47437, n47438;
  wire n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446;
  wire n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454;
  wire n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462;
  wire n47463, n47464, n47465, n47466, n47467, n47469, n47470, n47471;
  wire n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479;
  wire n47480, n47481, n47484, n47485, n47486, n47487, n47488, n47489;
  wire n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497;
  wire n47498, n47499, n47500, n47501, n47502, n47503, n47505, n47506;
  wire n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514;
  wire n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522;
  wire n47523, n47524, n47525, n47528, n47529, n47530, n47533, n47534;
  wire n47535, n47537, n47538, n47539, n47540, n47541, n47542, n47543;
  wire n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551;
  wire n47552, n47553, n47554, n47555, n47556, n47557, n47560, n47561;
  wire n47562, n47565, n47566, n47567, n47569, n47570, n47571, n47572;
  wire n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580;
  wire n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588;
  wire n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596;
  wire n47597, n47598, n47599, n47602, n47603, n47604, n47606, n47607;
  wire n47608, n47610, n47611, n47612, n47614, n47615, n47616, n47617;
  wire n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625;
  wire n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633;
  wire n47634, n47637, n47638, n47639, n47642, n47643, n47644, n47647;
  wire n47648, n47649, n47651, n47652, n47653, n47654, n47655, n47656;
  wire n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664;
  wire n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672;
  wire n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680;
  wire n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688;
  wire n47689, n47691, n47692, n47693, n47695, n47696, n47697, n47699;
  wire n47700, n47701, n47703, n47704, n47705, n47706, n47707, n47708;
  wire n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716;
  wire n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724;
  wire n47725, n47726, n47727, n47728, n47729, n47730, n47733, n47734;
  wire n47735, n47737, n47738, n47739, n47741, n47742, n47743, n47745;
  wire n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753;
  wire n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761;
  wire n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769;
  wire n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777;
  wire n47778, n47780, n47781, n47782, n47784, n47785, n47786, n47788;
  wire n47789, n47790, n47792, n47793, n47794, n47796, n47797, n47798;
  wire n47800, n47801, n47802, n47804, n47805, n47806, n47808, n47809;
  wire n47810, n47812, n47813, n47814, n47816, n47817, n47818, n47820;
  wire n47821, n47822, n47824, n47825, n47826, n47828, n47829, n47830;
  wire n47832, n47833, n47834, n47836, n47837, n47838, n47839, n47840;
  wire n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848;
  wire n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856;
  wire n47857, n47858, n47859, n47862, n47863, n47864, n47865, n47868;
  wire n47869, n47870, n47872, n47873, n47874, n47875, n47876, n47877;
  wire n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885;
  wire n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47895;
  wire n47896, n47897, n47900, n47901, n47902, n47903, n47904, n47908;
  wire n47909, n47910, n47912, n47913, n47914, n47916, n47917, n47918;
  wire n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927;
  wire n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935;
  wire n47936, n47937, n47938, n47939, n47940, n47941, n47944, n47945;
  wire n47946, n47947, n47950, n47951, n47952, n47954, n47955, n47956;
  wire n47960, n47961, n47962, n47965, n47966, n47967, n47968, n47969;
  wire n47970, n47973, n47974, n47975, n47976, n47977, n47978, n47979;
  wire n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987;
  wire n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996;
  wire n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004;
  wire n48005, n48006, n48007, n48008, n48009, n48010, n48013, n48014;
  wire n48015, n48016, n48019, n48020, n48021, n48023, n48024, n48025;
  wire n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033;
  wire n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041;
  wire n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049;
  wire n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48058;
  wire n48059, n48060, n48062, n48063, n48064, n48065, n48066, n48067;
  wire n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075;
  wire n48076, n48077, n48078, n48079, n48082, n48083, n48084, n48087;
  wire n48088, n48089, n48090, n48094, n48095, n48096, n48098, n48099;
  wire n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107;
  wire n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115;
  wire n48116, n48117, n48121, n48122, n48123, n48124, n48125, n48126;
  wire n48127, n48128, n48129, n48130, n48132, n48133, n48134, n48135;
  wire n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143;
  wire n48144, n48145, n48146, n48147, n48148, n48149, n48152, n48153;
  wire n48154, n48157, n48158, n48159, n48160, n48164, n48165, n48166;
  wire n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175;
  wire n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183;
  wire n48184, n48185, n48186, n48187, n48191, n48192, n48193, n48194;
  wire n48195, n48196, n48197, n48198, n48199, n48200, n48202, n48203;
  wire n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211;
  wire n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219;
  wire n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227;
  wire n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235;
  wire n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244;
  wire n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252;
  wire n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260;
  wire n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268;
  wire n48269, n48270, n48271, n48272, n48275, n48276, n48277, n48278;
  wire n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286;
  wire n48287, n48288, n48289, n48290, n48291, n48293, n48294, n48295;
  wire n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303;
  wire n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311;
  wire n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319;
  wire n48320, n48321, n48324, n48325, n48326, n48328, n48329, n48330;
  wire n48332, n48333, n48334, n48336, n48337, n48338, n48340, n48341;
  wire n48342, n48344, n48345, n48346, n48348, n48349, n48350, n48352;
  wire n48353, n48354, n48356, n48357, n48358, n48360, n48361, n48362;
  wire n48363, n48364, n48365, n48366, n48367, n48371, n48372, n48373;
  wire n48374, n48375, n48377, n48378, n48379, n48381, n48382, n48383;
  wire n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391;
  wire n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48401;
  wire n48402, n48403, n48406, n48407, n48408, n48409, n48413, n48414;
  wire n48415, n48417, n48418, n48419, n48421, n48422, n48423, n48425;
  wire n48426, n48427, n48429, n48430, n48431, n48433, n48434, n48435;
  wire n48437, n48438, n48440, n48441, n48442, n48444, n48445, n48446;
  wire n48448, n48449, n48450, n48452, n48453, n48454, n48456, n48457;
  wire n48458, n48460, n48461, n48462, n48464, n48465, n48466, n48468;
  wire n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48478;
  wire n48479, n48481, n48482, n48483, n48485, n48486, n48487, n48489;
  wire n48490, n48491, n48493, n48494, n48495, n48497, n48498, n48499;
  wire n48501, n48502, n48503, n48505, n48506, n48507, n48509, n48510;
  wire n48511, n48513, n48514, n48515, n48517, n48518, n48519, n48521;
  wire n48522, n48523, n48525, n48526, n48527, n48529, n48530, n48531;
  wire n48533, n48534, n48535, n48537, n48538, n48539, n48541, n48542;
  wire n48543, n48545, n48546, n48547, n48550, n48551, n48552, n48555;
  wire n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563;
  wire n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571;
  wire n48573, n48574, n48575, n48577, n48578, n48579, n48581, n48582;
  wire n48583, n48588, n48589, n48590, n48591, n48592, n48593, n48594;
  wire n48595, n48596, n48597, n48598, n48599, n48600, n48602, n48603;
  wire n48604, n48606, n48607, n48608, n48609, n48611, n48612, n48613;
  wire n48614, n48616, n48617, n48618, n48620, n48621, n48622, n48623;
  wire n48624, n48625, n48626, n48628, n48629, n48630, n48632, n48633;
  wire n48634, n48635, n48640, n48641, n48642, n48643, n48644, n48645;
  wire n48646, n48647, n48649, n48650, n48651, n48653, n48654, n48655;
  wire n48660, n48661, n48662, n48663, n48667, n48668, n48670, n48672;
  wire n48673, n48675, n48676, n48678, n48679, n48681, n48682, n48684;
  wire n48685, n48687, n48688, n48690, n48691, n48693, n48694, n48696;
  wire n48697, n48699, n48700, n48702, n48703, n48704, n48706, n48707;
  wire n48712, n48713, n48714, n48715, n48716, n48718, n48719, n48721;
  wire n48722, n48724, n48725, n48727, n48728, n48730, n48731, n48733;
  wire n48734, n48736, n48737, n48738, n48740, n48741, n48743, n48744;
  wire n48746, n48747, n48749, n48750, n48752, n48753, n48755, n48756;
  wire n48758, n48759, n48761, n48762, n48764, n48765, n48767, n48768;
  wire n48770, n48772, n48774, n48776, n48779, n48780, n48781, n48783;
  wire n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791;
  wire n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799;
  wire n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807;
  wire n48808, n48809, n48810, n48812, n48813, n48814, n48815, n48816;
  wire n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824;
  wire n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832;
  wire n48833, n48834, n48835, n48836, n48837, n48838, n48840, n48841;
  wire n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849;
  wire n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857;
  wire n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865;
  wire n48866, n48868, n48869, n48870, n48871, n48872, n48873, n48874;
  wire n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882;
  wire n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890;
  wire n48891, n48892, n48893, n48894, n48896, n48897, n48899, n48904;
  wire n48907, n48909, n48910, n48912, n48913, n48915, n48916, n48918;
  wire n48919, n48922, n48923, n48925, n48926, n48928, n48929, n48931;
  wire n48932, n48934, n48935, n48937, n48938, n48940, n48941, n48943;
  wire n48944, n48946, n48947, n48949, n48950, n48952, n48953, n48955;
  wire n48956, n48958, n48959, n48961, n48962, n48964, n48965, n48967;
  wire n48968, n48970, n48971, n48973, n48974, n48976, n48977, n48979;
  wire n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48988;
  wire n48989, n48991, n48992, n48994, n48995, n48997, n48998, n49000;
  wire n49001, n49003, n49004, n49006, n49007, n49009, n49010, n49011;
  wire n49012, n49013, n49014, n49015, n49016, n49018, n49019, n49021;
  wire n49022, n49024, n49025, n49027, n49028, n49030, n49031, n49033;
  wire n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49042;
  wire n49043, n49045, n49046, n49047, n49048, n49049, n49050, n49051;
  wire n49052, n49054, n49055, n49056, n49057, n49058, n49059, n49060;
  wire n49061, n49063, n49064, n49065, n49066, n49067, n49068, n49069;
  wire n49070, n49072, n49073, n49075, n49076, n49078, n49080, n49081;
  wire n49083, n49084, n49086, n49087, n49089, n49091, n49092, n49094;
  wire n49095, n49097, n49098, n49100, n49101, n49103, n49104, n49106;
  wire n49107, n49109, n49110, n49112, n49113, n49115, n49116, n49118;
  wire n49120, n49121, n49123, n49124, n49126, n49127, n49129, n49131;
  wire n49133, n49134, n49136, n49137, n49138, n49139, n49140, n49141;
  wire n49142, n49143, n49144, n49145, n49147, n49149, n49150, n49152;
  wire n49153, n49155, n49156, n49158, n49160, n49161, n49163, n49165;
  wire n49166, n49168, n49170, n49171, n49173, n49174, n49176, n49177;
  wire n49179, n49180, n49182, n49184, n49185, n49187, n49188, n49193;
  wire n49194, n49196, n49197, n49199, n49200, n49202, n49204, n49205;
  wire n49207, n49208, n49210, n49211, n49213, n49215, n49217, n49218;
  wire n49220, n49222, n49223, n49225, n49226, n49228, n49230, n49231;
  wire n49233, n49235, n49236, n49238, n49239, n49241, n49242, n49244;
  wire n49245, n49248, n49250, n49252, n49253, n49256, n_4, n_5;
  wire n_7, n_10, n_15, n_17, n_19, n_20, n_21, n_22;
  wire n_23, n_24, n_26, n_27, n_29, n_31, n_32, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_42, n_43;
  wire n_46, n_47, n_49, n_51, n_53, n_56, n_57, n_60;
  wire n_61, n_64, n_65, n_68, n_69, n_72, n_73, n_76;
  wire n_77, n_79, n_81, n_83, n_85, n_87, n_90, n_91;
  wire n_94, n_95, n_97, n_100, n_101, n_103, n_105, n_108;
  wire n_109, n_112, n_113, n_116, n_117, n_119, n_122, n_123;
  wire n_125, n_127, n_130, n_131, n_134, n_135, n_138, n_139;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_152, n_153, n_154, n_157, n_158, n_161, n_162;
  wire n_164, n_167, n_168, n_171, n_172, n_174, n_176, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_219, n_221;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_263, n_264;
  wire n_266, n_268, n_269, n_271, n_272, n_273, n_274, n_275;
  wire n_276, n_277, n_278, n_280, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_298, n_299, n_301, n_302, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_329, n_330, n_331;
  wire n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339;
  wire n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347;
  wire n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475;
  wire n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_484;
  wire n_485, n_486, n_489, n_494, n_495, n_497, n_498, n_499;
  wire n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523;
  wire n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555;
  wire n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672;
  wire n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704;
  wire n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_780, n_781, n_782, n_783, n_784;
  wire n_785, n_786, n_787, n_788, n_789, n_790, n_791, n_792;
  wire n_793, n_794, n_796, n_797, n_798, n_799, n_800, n_803;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837;
  wire n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845;
  wire n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853;
  wire n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861;
  wire n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869;
  wire n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877;
  wire n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885;
  wire n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893;
  wire n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901;
  wire n_902, n_903, n_904, n_906, n_907, n_908, n_909, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934;
  wire n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_942;
  wire n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_974;
  wire n_975, n_976, n_977, n_978, n_981, n_983, n_984, n_985;
  wire n_986, n_988, n_989, n_990, n_991, n_992, n_993, n_994;
  wire n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002;
  wire n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010;
  wire n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018;
  wire n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026;
  wire n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034;
  wire n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042;
  wire n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050;
  wire n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093;
  wire n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101;
  wire n_1102, n_1103, n_1104, n_1105, n_1106, n_1109, n_1110, n_1111;
  wire n_1112, n_1115, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131;
  wire n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139;
  wire n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147;
  wire n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171;
  wire n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179;
  wire n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187;
  wire n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195;
  wire n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219;
  wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1226, n_1229, n_1230;
  wire n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246;
  wire n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254;
  wire n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262;
  wire n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278;
  wire n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286;
  wire n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1295, n_1296;
  wire n_1297, n_1298, n_1301, n_1304, n_1305, n_1306, n_1307, n_1308;
  wire n_1309, n_1310, n_1311, n_1313, n_1314, n_1315, n_1316, n_1317;
  wire n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325;
  wire n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
  wire n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446;
  wire n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
  wire n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462;
  wire n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470;
  wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478;
  wire n_1479, n_1480, n_1481, n_1482, n_1483, n_1486, n_1489, n_1490;
  wire n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523;
  wire n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531;
  wire n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539;
  wire n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563;
  wire n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571;
  wire n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579;
  wire n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587;
  wire n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1595, n_1598;
  wire n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606;
  wire n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614;
  wire n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622;
  wire n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638;
  wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654;
  wire n_1655, n_1656, n_1657, n_1660, n_1661, n_1662, n_1663, n_1666;
  wire n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
  wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
  wire n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765;
  wire n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1774;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
  wire n_1833, n_1834, n_1835, n_1836, n_1839, n_1840, n_1841, n_1842;
  wire n_1844, n_1846, n_1847, n_1848, n_1849, n_1851, n_1853, n_1854;
  wire n_1855, n_1856, n_1857, n_1859, n_1860, n_1861, n_1862, n_1863;
  wire n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871;
  wire n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879;
  wire n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887;
  wire n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895;
  wire n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903;
  wire n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911;
  wire n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919;
  wire n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927;
  wire n_1928, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937;
  wire n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945;
  wire n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953;
  wire n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962;
  wire n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970;
  wire n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978;
  wire n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986;
  wire n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994;
  wire n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002;
  wire n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010;
  wire n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2020;
  wire n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030;
  wire n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039;
  wire n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079;
  wire n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087;
  wire n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
  wire n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103;
  wire n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111;
  wire n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
  wire n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2128;
  wire n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138;
  wire n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146;
  wire n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154;
  wire n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162;
  wire n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170;
  wire n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186;
  wire n_2187, n_2188, n_2189, n_2190, n_2193, n_2194, n_2195, n_2196;
  wire n_2199, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217;
  wire n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225;
  wire n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233;
  wire n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241;
  wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249;
  wire n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257;
  wire n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265;
  wire n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273;
  wire n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281;
  wire n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289;
  wire n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297;
  wire n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305;
  wire n_2307, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316;
  wire n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324;
  wire n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332;
  wire n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356;
  wire n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364;
  wire n_2365, n_2366, n_2367, n_2368, n_2369, n_2372, n_2373, n_2374;
  wire n_2375, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385;
  wire n_2386, n_2387, n_2388, n_2390, n_2391, n_2392, n_2393, n_2394;
  wire n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402;
  wire n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410;
  wire n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418;
  wire n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426;
  wire n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434;
  wire n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442;
  wire n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450;
  wire n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458;
  wire n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466;
  wire n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474;
  wire n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482;
  wire n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490;
  wire n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2498, n_2499;
  wire n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507;
  wire n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515;
  wire n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523;
  wire n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531;
  wire n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539;
  wire n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547;
  wire n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555;
  wire n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563;
  wire n_2564, n_2565, n_2566, n_2567, n_2568, n_2572, n_2573, n_2574;
  wire n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2583;
  wire n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591;
  wire n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599;
  wire n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607;
  wire n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615;
  wire n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623;
  wire n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631;
  wire n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639;
  wire n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647;
  wire n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655;
  wire n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663;
  wire n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671;
  wire n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679;
  wire n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2688;
  wire n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696;
  wire n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704;
  wire n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712;
  wire n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744;
  wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
  wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
  wire n_2761, n_2763, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770;
  wire n_2771, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779;
  wire n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787;
  wire n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795;
  wire n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803;
  wire n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811;
  wire n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819;
  wire n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827;
  wire n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835;
  wire n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843;
  wire n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851;
  wire n_2852, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860;
  wire n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868;
  wire n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2876;
  wire n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884;
  wire n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892;
  wire n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900;
  wire n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908;
  wire n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916;
  wire n_2917, n_2918, n_2919, n_2921, n_2922, n_2923, n_2924, n_2925;
  wire n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933;
  wire n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941;
  wire n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949;
  wire n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957;
  wire n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965;
  wire n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973;
  wire n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981;
  wire n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989;
  wire n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997;
  wire n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005;
  wire n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013;
  wire n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021;
  wire n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, n_3029;
  wire n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037;
  wire n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045;
  wire n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053;
  wire n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061;
  wire n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, n_3069;
  wire n_3070, n_3071, n_3072, n_3073, n_3074, n_3078, n_3080, n_3081;
  wire n_3082, n_3084, n_3087, n_3090, n_3091, n_3093, n_3096, n_3098;
  wire n_3100, n_3102, n_3105, n_3106, n_3119, n_3120, n_3121, n_3122;
  wire n_3123, n_3124, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131;
  wire n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139;
  wire n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3148, n_3149;
  wire n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169;
  wire n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177;
  wire n_3178, n_3181, n_3182, n_3184, n_3187, n_3188, n_3190, n_3193;
  wire n_3194, n_3197, n_3198, n_3200, n_3202, n_3206, n_3208, n_3209;
  wire n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217;
  wire n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225;
  wire n_3226, n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233;
  wire n_3234, n_3235, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242;
  wire n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250;
  wire n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258;
  wire n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266;
  wire n_3267, n_3268, n_3269, n_3270, n_3271, n_3274, n_3275, n_3276;
  wire n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284;
  wire n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292;
  wire n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300;
  wire n_3301, n_3302, n_3307, n_3308, n_3310, n_3311, n_3312, n_3313;
  wire n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321;
  wire n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330;
  wire n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338;
  wire n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346;
  wire n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354;
  wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362;
  wire n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370;
  wire n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378;
  wire n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386;
  wire n_3387, n_3388, n_3389, n_3390, n_3391, n_3396, n_3397, n_3398;
  wire n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3407;
  wire n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415;
  wire n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423;
  wire n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431;
  wire n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439;
  wire n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447;
  wire n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455;
  wire n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463;
  wire n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471;
  wire n_3472, n_3473, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482;
  wire n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490;
  wire n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498;
  wire n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, n_3506;
  wire n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514;
  wire n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522;
  wire n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530;
  wire n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537, n_3538;
  wire n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, n_3546;
  wire n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554;
  wire n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562;
  wire n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570;
  wire n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578;
  wire n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586;
  wire n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594;
  wire n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602;
  wire n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609, n_3610;
  wire n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, n_3618;
  wire n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626;
  wire n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634;
  wire n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642;
  wire n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, n_3650;
  wire n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658;
  wire n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666;
  wire n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674;
  wire n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681, n_3682;
  wire n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690;
  wire n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698;
  wire n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706;
  wire n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714;
  wire n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722;
  wire n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730;
  wire n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738;
  wire n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746;
  wire n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753, n_3754;
  wire n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762;
  wire n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770;
  wire n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778;
  wire n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786;
  wire n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794;
  wire n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802;
  wire n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810;
  wire n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818;
  wire n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826;
  wire n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834;
  wire n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842;
  wire n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850;
  wire n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858;
  wire n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866;
  wire n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874;
  wire n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882;
  wire n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890;
  wire n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897, n_3898;
  wire n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, n_3906;
  wire n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914;
  wire n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922;
  wire n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930;
  wire n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, n_3938;
  wire n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946;
  wire n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953, n_3954;
  wire n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961, n_3962;
  wire n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970;
  wire n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978;
  wire n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985, n_3986;
  wire n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993, n_3994;
  wire n_3995, n_3996, n_3997, n_3998, n_4000, n_4001, n_4005, n_4006;
  wire n_4007, n_4008, n_4009, n_4010, n_4011, n_4012, n_4013, n_4014;
  wire n_4015, n_4016, n_4017, n_4018, n_4019, n_4020, n_4021, n_4022;
  wire n_4023, n_4024, n_4025, n_4026, n_4027, n_4028, n_4032, n_4034;
  wire n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041, n_4042;
  wire n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049, n_4050;
  wire n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057, n_4058;
  wire n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065, n_4066;
  wire n_4067, n_4068, n_4069, n_4070, n_4073, n_4074, n_4075, n_4076;
  wire n_4081, n_4085, n_4086, n_4088, n_4090, n_4091, n_4093, n_4094;
  wire n_4095, n_4096, n_4097, n_4098, n_4099, n_4100, n_4101, n_4102;
  wire n_4103, n_4104, n_4105, n_4106, n_4107, n_4108, n_4109, n_4110;
  wire n_4111, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118;
  wire n_4119, n_4120, n_4121, n_4122, n_4123, n_4124, n_4125, n_4126;
  wire n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133, n_4134;
  wire n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141, n_4142;
  wire n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150;
  wire n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157, n_4158;
  wire n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165, n_4166;
  wire n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173, n_4174;
  wire n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181, n_4182;
  wire n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4189, n_4190;
  wire n_4191, n_4192, n_4193, n_4194, n_4195, n_4196, n_4197, n_4198;
  wire n_4199, n_4200, n_4201, n_4202, n_4203, n_4204, n_4205, n_4206;
  wire n_4208, n_4209, n_4210, n_4211, n_4212, n_4213, n_4214, n_4215;
  wire n_4216, n_4217, n_4218, n_4219, n_4220, n_4221, n_4222, n_4223;
  wire n_4224, n_4225, n_4226, n_4227, n_4228, n_4230, n_4231, n_4234;
  wire n_4235, n_4237, n_4239, n_4242, n_4243, n_4244, n_4245, n_4247;
  wire n_4248, n_4249, n_4250, n_4253, n_4254, n_4255, n_4256, n_4259;
  wire n_4260, n_4261, n_4262, n_4264, n_4265, n_4266, n_4267, n_4269;
  wire n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276, n_4277;
  wire n_4278, n_4279, n_4280, n_4282, n_4285, n_4286, n_4287, n_4288;
  wire n_4291, n_4292, n_4293, n_4294, n_4297, n_4298, n_4299, n_4300;
  wire n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309, n_4310;
  wire n_4311, n_4312, n_4313, n_4314, n_4316, n_4317, n_4318, n_4319;
  wire n_4320, n_4321, n_4323, n_4324, n_4325, n_4326, n_4327, n_4330;
  wire n_4331, n_4332, n_4333, n_4336, n_4337, n_4338, n_4339, n_4341;
  wire n_4342, n_4343, n_4344, n_4347, n_4348, n_4349, n_4350, n_4352;
  wire n_4353, n_4354, n_4355, n_4356, n_4357, n_4358, n_4359, n_4360;
  wire n_4361, n_4362, n_4363, n_4365, n_4366, n_4367, n_4368, n_4369;
  wire n_4370, n_4371, n_4373, n_4374, n_4375, n_4377, n_4380, n_4381;
  wire n_4382, n_4383, n_4385, n_4386, n_4387, n_4388, n_4391, n_4392;
  wire n_4393, n_4394, n_4396, n_4397, n_4398, n_4399, n_4401, n_4402;
  wire n_4403, n_4404, n_4406, n_4407, n_4408, n_4409, n_4411, n_4412;
  wire n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420;
  wire n_4421, n_4423, n_4424, n_4428, n_4429, n_4430, n_4431, n_4433;
  wire n_4434, n_4435, n_4436, n_4439, n_4440, n_4441, n_4442, n_4443;
  wire n_4444, n_4445, n_4446, n_4449, n_4450, n_4451, n_4452, n_4455;
  wire n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462, n_4463;
  wire n_4464, n_4465, n_4466, n_4469, n_4470, n_4471, n_4472, n_4474;
  wire n_4475, n_4476, n_4477, n_4480, n_4481, n_4482, n_4483, n_4485;
  wire n_4486, n_4487, n_4488, n_4491, n_4492, n_4493, n_4494, n_4495;
  wire n_4496, n_4497, n_4498, n_4500, n_4501, n_4502, n_4503, n_4504;
  wire n_4505, n_4506, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512;
  wire n_4513, n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520;
  wire n_4523, n_4524, n_4525, n_4526, n_4529, n_4530, n_4531, n_4532;
  wire n_4534, n_4535, n_4536, n_4537, n_4540, n_4541, n_4542, n_4543;
  wire n_4545, n_4546, n_4547, n_4548, n_4549, n_4550, n_4551, n_4552;
  wire n_4553, n_4554, n_4555, n_4556, n_4558, n_4559, n_4560, n_4561;
  wire n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568, n_4569;
  wire n_4570, n_4571, n_4572, n_4573, n_4575, n_4576, n_4577, n_4578;
  wire n_4579, n_4580, n_4581, n_4582, n_4583, n_4585, n_4586, n_4587;
  wire n_4588, n_4589, n_4590, n_4591, n_4593, n_4594, n_4595, n_4596;
  wire n_4597, n_4600, n_4601, n_4602, n_4603, n_4606, n_4607, n_4608;
  wire n_4609, n_4610, n_4611, n_4612, n_4613, n_4615, n_4616, n_4617;
  wire n_4618, n_4619, n_4620, n_4621, n_4622, n_4623, n_4624, n_4625;
  wire n_4626, n_4628, n_4629, n_4630, n_4633, n_4634, n_4635, n_4636;
  wire n_4639, n_4640, n_4641, n_4642, n_4644, n_4645, n_4646, n_4647;
  wire n_4650, n_4651, n_4652, n_4653, n_4656, n_4657, n_4658, n_4659;
  wire n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667;
  wire n_4668, n_4669, n_4670, n_4671, n_4672, n_4675, n_4676, n_4677;
  wire n_4678, n_4681, n_4682, n_4683, n_4684, n_4686, n_4687, n_4688;
  wire n_4689, n_4692, n_4693, n_4694, n_4695, n_4697, n_4698, n_4699;
  wire n_4700, n_4701, n_4702, n_4703, n_4704, n_4705, n_4706, n_4707;
  wire n_4708, n_4710, n_4711, n_4712, n_4713, n_4714, n_4715, n_4716;
  wire n_4717, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724;
  wire n_4725, n_4726, n_4728, n_4729, n_4732, n_4733, n_4734, n_4735;
  wire n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4745;
  wire n_4748, n_4749, n_4750, n_4751, n_4753, n_4754, n_4755, n_4756;
  wire n_4758, n_4759, n_4760, n_4761, n_4763, n_4764, n_4765, n_4766;
  wire n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774;
  wire n_4775, n_4776, n_4778, n_4779, n_4780, n_4781, n_4782, n_4783;
  wire n_4785, n_4786, n_4787, n_4788, n_4789, n_4790, n_4791, n_4793;
  wire n_4794, n_4795, n_4796, n_4797, n_4800, n_4801, n_4802, n_4803;
  wire n_4806, n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813;
  wire n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822;
  wire n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830;
  wire n_4832, n_4833, n_4834, n_4837, n_4838, n_4839, n_4840, n_4842;
  wire n_4843, n_4844, n_4845, n_4848, n_4849, n_4850, n_4851, n_4852;
  wire n_4853, n_4854, n_4855, n_4858, n_4859, n_4860, n_4861, n_4864;
  wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4872;
  wire n_4873, n_4874, n_4875, n_4878, n_4879, n_4880, n_4881, n_4884;
  wire n_4885, n_4886, n_4887, n_4888, n_4889, n_4890, n_4891, n_4894;
  wire n_4895, n_4896, n_4897, n_4900, n_4901, n_4902, n_4903, n_4904;
  wire n_4905, n_4906, n_4907, n_4908, n_4909, n_4910, n_4911, n_4913;
  wire n_4914, n_4915, n_4916, n_4917, n_4918, n_4921, n_4922, n_4923;
  wire n_4924, n_4927, n_4928, n_4929, n_4930, n_4933, n_4934, n_4935;
  wire n_4936, n_4937, n_4938, n_4939, n_4940, n_4941, n_4942, n_4943;
  wire n_4944, n_4947, n_4948, n_4949, n_4950, n_4952, n_4953, n_4954;
  wire n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4964;
  wire n_4965, n_4966, n_4967, n_4969, n_4970, n_4971, n_4972, n_4974;
  wire n_4976, n_4977, n_4978, n_4980, n_4981, n_4982, n_4983, n_4985;
  wire n_4986, n_4987, n_4988, n_4990, n_4991, n_4992, n_4993, n_4995;
  wire n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003;
  wire n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011;
  wire n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019;
  wire n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027;
  wire n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035;
  wire n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043;
  wire n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051;
  wire n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5058, n_5059;
  wire n_5060, n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067;
  wire n_5068, n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075;
  wire n_5076, n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083;
  wire n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091;
  wire n_5092, n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099;
  wire n_5100, n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107;
  wire n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115;
  wire n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123;
  wire n_5124, n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131;
  wire n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139;
  wire n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147;
  wire n_5148, n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155;
  wire n_5156, n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163;
  wire n_5164, n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171;
  wire n_5172, n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179;
  wire n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187;
  wire n_5188, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195;
  wire n_5196, n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203;
  wire n_5204, n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211;
  wire n_5212, n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219;
  wire n_5220, n_5221, n_5222, n_5226, n_5227, n_5228, n_5231, n_5232;
  wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
  wire n_5241, n_5242, n_5243, n_5244, n_5245, n_5246, n_5247, n_5248;
  wire n_5249, n_5250, n_5251, n_5252, n_5253, n_5254, n_5255, n_5256;
  wire n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263, n_5264;
  wire n_5265, n_5266, n_5267, n_5268, n_5269, n_5270, n_5271, n_5272;
  wire n_5273, n_5274, n_5275, n_5276, n_5277, n_5278, n_5279, n_5280;
  wire n_5281, n_5282, n_5283, n_5284, n_5285, n_5286, n_5287, n_5288;
  wire n_5289, n_5290, n_5291, n_5292, n_5293, n_5294, n_5295, n_5296;
  wire n_5297, n_5298, n_5299, n_5300, n_5301, n_5302, n_5303, n_5304;
  wire n_5305, n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312;
  wire n_5313, n_5314, n_5315, n_5316, n_5317, n_5318, n_5319, n_5320;
  wire n_5321, n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5328;
  wire n_5329, n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336;
  wire n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5343, n_5344;
  wire n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5351, n_5352;
  wire n_5353, n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5360;
  wire n_5361, n_5362, n_5363, n_5364, n_5365, n_5366, n_5367, n_5368;
  wire n_5369, n_5370, n_5371, n_5372, n_5373, n_5374, n_5375, n_5376;
  wire n_5377, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383, n_5384;
  wire n_5385, n_5386, n_5387, n_5388, n_5389, n_5390, n_5391, n_5392;
  wire n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5399, n_5400;
  wire n_5401, n_5402, n_5403, n_5404, n_5405, n_5406, n_5407, n_5408;
  wire n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416;
  wire n_5417, n_5418, n_5419, n_5420, n_5421, n_5422, n_5423, n_5424;
  wire n_5425, n_5426, n_5427, n_5428, n_5429, n_5430, n_5431, n_5432;
  wire n_5433, n_5434, n_5435, n_5436, n_5437, n_5438, n_5439, n_5440;
  wire n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447, n_5448;
  wire n_5449, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456;
  wire n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464;
  wire n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472;
  wire n_5473, n_5474, n_5475, n_5476, n_5477, n_5478, n_5479, n_5480;
  wire n_5481, n_5482, n_5483, n_5484, n_5485, n_5486, n_5487, n_5488;
  wire n_5489, n_5490, n_5491, n_5492, n_5493, n_5494, n_5495, n_5496;
  wire n_5497, n_5498, n_5499, n_5500, n_5501, n_5502, n_5503, n_5504;
  wire n_5505, n_5506, n_5507, n_5508, n_5509, n_5510, n_5511, n_5512;
  wire n_5513, n_5514, n_5515, n_5516, n_5517, n_5518, n_5519, n_5520;
  wire n_5521, n_5522, n_5523, n_5524, n_5525, n_5526, n_5527, n_5528;
  wire n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536;
  wire n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544;
  wire n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552;
  wire n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560;
  wire n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
  wire n_5569, n_5570, n_5571, n_5572, n_5573, n_5574, n_5575, n_5576;
  wire n_5577, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584;
  wire n_5585, n_5586, n_5587, n_5588, n_5589, n_5590, n_5591, n_5592;
  wire n_5593, n_5594, n_5595, n_5596, n_5597, n_5598, n_5599, n_5600;
  wire n_5601, n_5602, n_5603, n_5604, n_5605, n_5606, n_5607, n_5608;
  wire n_5609, n_5610, n_5611, n_5612, n_5613, n_5614, n_5615, n_5616;
  wire n_5617, n_5618, n_5619, n_5620, n_5621, n_5622, n_5623, n_5624;
  wire n_5625, n_5626, n_5627, n_5629, n_5630, n_5631, n_5632, n_5633;
  wire n_5634, n_5636, n_5637, n_5638, n_5639, n_5640, n_5641, n_5642;
  wire n_5643, n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652;
  wire n_5653, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660;
  wire n_5661, n_5662, n_5663, n_5664, n_5665, n_5668, n_5669, n_5671;
  wire n_5673, n_5675, n_5677, n_5679, n_5681, n_5682, n_5685, n_5686;
  wire n_5687, n_5688, n_5689, n_5690, n_5691, n_5693, n_5694, n_5695;
  wire n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703;
  wire n_5704, n_5705, n_5708, n_5709, n_5710, n_5711, n_5712, n_5713;
  wire n_5714, n_5715, n_5716, n_5717, n_5719, n_5720, n_5721, n_5722;
  wire n_5723, n_5724, n_5726, n_5727, n_5728, n_5729, n_5730, n_5731;
  wire n_5732, n_5733, n_5734, n_5735, n_5736, n_5737, n_5738, n_5739;
  wire n_5740, n_5742, n_5743, n_5744, n_5745, n_5746, n_5747, n_5748;
  wire n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5756;
  wire n_5757, n_5758, n_5759, n_5760, n_5761, n_5762, n_5763, n_5764;
  wire n_5765, n_5766, n_5767, n_5768, n_5769, n_5770, n_5771, n_5772;
  wire n_5773, n_5774, n_5775, n_5776, n_5777, n_5778, n_5779, n_5780;
  wire n_5781, n_5782, n_5783, n_5785, n_5786, n_5787, n_5788, n_5789;
  wire n_5790, n_5791, n_5792, n_5793, n_5794, n_5795, n_5796, n_5797;
  wire n_5798, n_5801, n_5802, n_5803, n_5804, n_5805, n_5806, n_5810;
  wire n_5811, n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818;
  wire n_5819, n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826;
  wire n_5827, n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834;
  wire n_5835, n_5836, n_5837, n_5838, n_5839, n_5840, n_5841, n_5842;
  wire n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5850;
  wire n_5851, n_5852, n_5853, n_5854, n_5855, n_5856, n_5857, n_5858;
  wire n_5859, n_5860, n_5861, n_5862, n_5863, n_5864, n_5865, n_5866;
  wire n_5867, n_5868, n_5869, n_5870, n_5871, n_5872, n_5873, n_5874;
  wire n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881, n_5882;
  wire n_5883, n_5884, n_5885, n_5886, n_5887, n_5888, n_5889, n_5890;
  wire n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897, n_5898;
  wire n_5899, n_5900, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906;
  wire n_5907, n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914;
  wire n_5915, n_5916, n_5917, n_5918, n_5919, n_5920, n_5923, n_5924;
  wire n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931, n_5932;
  wire n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939, n_5940;
  wire n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947, n_5948;
  wire n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955, n_5956;
  wire n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963, n_5964;
  wire n_5965, n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972;
  wire n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980;
  wire n_5981, n_5982, n_5983, n_5984, n_5985, n_5986, n_5987, n_5988;
  wire n_5989, n_5990, n_5991, n_5992, n_5993, n_5994, n_5995, n_5996;
  wire n_5997, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004;
  wire n_6005, n_6006, n_6007, n_6008, n_6009, n_6010, n_6011, n_6012;
  wire n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020;
  wire n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027, n_6028;
  wire n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036;
  wire n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044;
  wire n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052;
  wire n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060;
  wire n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068;
  wire n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076;
  wire n_6077, n_6078, n_6079, n_6080, n_6081, n_6082, n_6083, n_6084;
  wire n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092;
  wire n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100;
  wire n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107, n_6108;
  wire n_6109, n_6110, n_6111, n_6112, n_6113, n_6114, n_6115, n_6116;
  wire n_6117, n_6118, n_6119, n_6120, n_6121, n_6122, n_6123, n_6124;
  wire n_6125, n_6126, n_6127, n_6128, n_6129, n_6130, n_6131, n_6132;
  wire n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6139, n_6140;
  wire n_6141, n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148;
  wire n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6157, n_6158;
  wire n_6159, n_6160, n_6161, n_6162, n_6163, n_6164, n_6165, n_6166;
  wire n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6174;
  wire n_6175, n_6176, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182;
  wire n_6183, n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190;
  wire n_6191, n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198;
  wire n_6199, n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206;
  wire n_6207, n_6208, n_6209, n_6210, n_6211, n_6212, n_6213, n_6214;
  wire n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6221, n_6223;
  wire n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231;
  wire n_6232, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240;
  wire n_6241, n_6242, n_6244, n_6245, n_6246, n_6247, n_6248, n_6249;
  wire n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256, n_6258;
  wire n_6259, n_6260, n_6261, n_6262, n_6263, n_6264, n_6266, n_6267;
  wire n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275;
  wire n_6276, n_6277, n_6278, n_6280, n_6281, n_6282, n_6283, n_6284;
  wire n_6285, n_6286, n_6287, n_6288, n_6290, n_6291, n_6292, n_6293;
  wire n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300, n_6301;
  wire n_6302, n_6303, n_6304, n_6305, n_6306, n_6307, n_6308, n_6309;
  wire n_6310, n_6311, n_6312, n_6313, n_6314, n_6315, n_6319, n_6320;
  wire n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328;
  wire n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336;
  wire n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344;
  wire n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6352;
  wire n_6353, n_6354, n_6355, n_6356, n_6357, n_6358, n_6359, n_6360;
  wire n_6361, n_6362, n_6363, n_6364, n_6365, n_6366, n_6367, n_6368;
  wire n_6369, n_6370, n_6371, n_6372, n_6373, n_6374, n_6375, n_6376;
  wire n_6377, n_6378, n_6379, n_6380, n_6381, n_6382, n_6383, n_6384;
  wire n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391, n_6392;
  wire n_6393, n_6394, n_6395, n_6396, n_6397, n_6398, n_6399, n_6400;
  wire n_6401, n_6402, n_6403, n_6404, n_6405, n_6406, n_6407, n_6408;
  wire n_6409, n_6410, n_6411, n_6412, n_6413, n_6414, n_6415, n_6416;
  wire n_6417, n_6420, n_6421, n_6422, n_6423, n_6424, n_6425, n_6426;
  wire n_6427, n_6428, n_6429, n_6430, n_6431, n_6432, n_6433, n_6434;
  wire n_6435, n_6436, n_6437, n_6438, n_6439, n_6440, n_6441, n_6442;
  wire n_6443, n_6444, n_6445, n_6446, n_6447, n_6448, n_6449, n_6450;
  wire n_6451, n_6452, n_6453, n_6454, n_6455, n_6456, n_6457, n_6458;
  wire n_6459, n_6460, n_6461, n_6462, n_6463, n_6464, n_6465, n_6466;
  wire n_6467, n_6468, n_6469, n_6470, n_6471, n_6472, n_6473, n_6474;
  wire n_6475, n_6476, n_6477, n_6478, n_6479, n_6480, n_6481, n_6482;
  wire n_6483, n_6484, n_6485, n_6486, n_6487, n_6488, n_6489, n_6490;
  wire n_6491, n_6492, n_6493, n_6494, n_6495, n_6496, n_6497, n_6498;
  wire n_6499, n_6500, n_6501, n_6504, n_6505, n_6506, n_6507, n_6508;
  wire n_6509, n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6516;
  wire n_6517, n_6518, n_6519, n_6520, n_6521, n_6522, n_6523, n_6524;
  wire n_6525, n_6526, n_6527, n_6528, n_6529, n_6530, n_6531, n_6532;
  wire n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539, n_6540;
  wire n_6541, n_6542, n_6543, n_6544, n_6545, n_6546, n_6547, n_6548;
  wire n_6549, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555, n_6556;
  wire n_6557, n_6558, n_6559, n_6560, n_6561, n_6562, n_6563, n_6564;
  wire n_6565, n_6566, n_6567, n_6570, n_6572, n_6576, n_6579, n_6580;
  wire n_6581, n_6582, n_6583, n_6584, n_6585, n_6586, n_6587, n_6590;
  wire n_6591, n_6592, n_6593, n_6594, n_6595, n_6596, n_6598, n_6599;
  wire n_6600, n_6601, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608;
  wire n_6609, n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616;
  wire n_6617, n_6618, n_6619, n_6620, n_6621, n_6622, n_6624, n_6625;
  wire n_6626, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6634;
  wire n_6635, n_6638, n_6639, n_6640, n_6641, n_6642, n_6643, n_6644;
  wire n_6645, n_6646, n_6647, n_6648, n_6649, n_6650, n_6651, n_6652;
  wire n_6653, n_6654, n_6655, n_6656, n_6657, n_6658, n_6659, n_6660;
  wire n_6661, n_6662, n_6663, n_6664, n_6665, n_6666, n_6667, n_6668;
  wire n_6669, n_6670, n_6671, n_6672, n_6673, n_6674, n_6675, n_6676;
  wire n_6677, n_6678, n_6679, n_6680, n_6681, n_6682, n_6683, n_6684;
  wire n_6685, n_6686, n_6689, n_6690, n_6691, n_6692, n_6693, n_6694;
  wire n_6695, n_6696, n_6697, n_6698, n_6699, n_6700, n_6701, n_6702;
  wire n_6703, n_6704, n_6705, n_6708, n_6710, n_6712, n_6713, n_6715;
  wire n_6716, n_6717, n_6718, n_6721, n_6722, n_6723, n_6724, n_6725;
  wire n_6726, n_6727, n_6728, n_6729, n_6730, n_6731, n_6732, n_6733;
  wire n_6734, n_6735, n_6736, n_6737, n_6738, n_6739, n_6740, n_6741;
  wire n_6742, n_6743, n_6744, n_6745, n_6746, n_6747, n_6748, n_6749;
  wire n_6750, n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757;
  wire n_6758, n_6759, n_6760, n_6761, n_6762, n_6763, n_6764, n_6765;
  wire n_6766, n_6767, n_6768, n_6769, n_6770, n_6771, n_6772, n_6773;
  wire n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783, n_6785;
  wire n_6786, n_6791, n_6792, n_6795, n_6796, n_6797, n_6798, n_6799;
  wire n_6800, n_6801, n_6802, n_6803, n_6804, n_6805, n_6806, n_6807;
  wire n_6808, n_6810, n_6811, n_6812, n_6813, n_6814, n_6815, n_6816;
  wire n_6817, n_6818, n_6819, n_6820, n_6821, n_6822, n_6823, n_6824;
  wire n_6825, n_6826, n_6827, n_6828, n_6829, n_6830, n_6831, n_6832;
  wire n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6839, n_6840;
  wire n_6841, n_6842, n_6843, n_6844, n_6845, n_6846, n_6847, n_6848;
  wire n_6849, n_6850, n_6851, n_6852, n_6853, n_6854, n_6855, n_6856;
  wire n_6857, n_6858, n_6859, n_6860, n_6863, n_6864, n_6865, n_6866;
  wire n_6867, n_6868, n_6869, n_6870, n_6871, n_6872, n_6873, n_6874;
  wire n_6875, n_6876, n_6877, n_6878, n_6879, n_6880, n_6881, n_6882;
  wire n_6883, n_6884, n_6885, n_6886, n_6887, n_6888, n_6889, n_6890;
  wire n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6898;
  wire n_6899, n_6900, n_6901, n_6903, n_6904, n_6905, n_6906, n_6907;
  wire n_6908, n_6909, n_6910, n_6911, n_6912, n_6913, n_6914, n_6915;
  wire n_6916, n_6917, n_6918, n_6919, n_6920, n_6921, n_6922, n_6923;
  wire n_6924, n_6925, n_6926, n_6927, n_6928, n_6929, n_6930, n_6931;
  wire n_6932, n_6933, n_6934, n_6935, n_6936, n_6937, n_6938, n_6939;
  wire n_6940, n_6941, n_6942, n_6943, n_6947, n_6948, n_6949, n_6950;
  wire n_6951, n_6952, n_6953, n_6954, n_6955, n_6956, n_6957, n_6958;
  wire n_6959, n_6960, n_6961, n_6962, n_6963, n_6964, n_6965, n_6966;
  wire n_6967, n_6968, n_6969, n_6970, n_6971, n_6972, n_6973, n_6974;
  wire n_6975, n_6976, n_6977, n_6978, n_6979, n_6980, n_6981, n_6982;
  wire n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6989, n_6990;
  wire n_6991, n_6992, n_6993, n_6994, n_6995, n_6996, n_6997, n_6998;
  wire n_6999, n_7000, n_7001, n_7002, n_7003, n_7004, n_7005, n_7006;
  wire n_7007, n_7008, n_7009, n_7010, n_7011, n_7012, n_7013, n_7014;
  wire n_7015, n_7016, n_7017, n_7018, n_7019, n_7020, n_7021, n_7022;
  wire n_7023, n_7024, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030;
  wire n_7031, n_7032, n_7033, n_7034, n_7038, n_7039, n_7040, n_7041;
  wire n_7042, n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049;
  wire n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7056, n_7057;
  wire n_7058, n_7059, n_7060, n_7061, n_7065, n_7066, n_7067, n_7068;
  wire n_7069, n_7070, n_7071, n_7072, n_7073, n_7074, n_7075, n_7076;
  wire n_7077, n_7078, n_7079, n_7080, n_7081, n_7082, n_7083, n_7084;
  wire n_7085, n_7086, n_7087, n_7088, n_7089, n_7090, n_7094, n_7095;
  wire n_7096, n_7097, n_7098, n_7099, n_7100, n_7101, n_7102, n_7103;
  wire n_7104, n_7105, n_7106, n_7107, n_7111, n_7112, n_7113, n_7114;
  wire n_7115, n_7116, n_7117, n_7118, n_7119, n_7120, n_7121, n_7122;
  wire n_7123, n_7124, n_7125, n_7126, n_7127, n_7128, n_7129, n_7130;
  wire n_7131, n_7132, n_7133, n_7134, n_7135, n_7136, n_7137, n_7138;
  wire n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145, n_7146;
  wire n_7147, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153, n_7154;
  wire n_7155, n_7156, n_7157, n_7158, n_7159, n_7160, n_7161, n_7162;
  wire n_7163, n_7164, n_7165, n_7166, n_7170, n_7171, n_7172, n_7173;
  wire n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181;
  wire n_7182, n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190;
  wire n_7191, n_7192, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198;
  wire n_7199, n_7200, n_7201, n_7202, n_7206, n_7209, n_7210, n_7211;
  wire n_7212, n_7213, n_7217, n_7218, n_7219, n_7220, n_7221, n_7222;
  wire n_7223, n_7224, n_7225, n_7226, n_7227, n_7228, n_7229, n_7230;
  wire n_7231, n_7232, n_7233, n_7234, n_7235, n_7236, n_7237, n_7238;
  wire n_7239, n_7240, n_7241, n_7242, n_7243, n_7244, n_7245, n_7246;
  wire n_7247, n_7248, n_7249, n_7250, n_7251, n_7252, n_7253, n_7254;
  wire n_7255, n_7256, n_7257, n_7258, n_7259, n_7260, n_7261, n_7262;
  wire n_7263, n_7264, n_7265, n_7266, n_7267, n_7268, n_7269, n_7270;
  wire n_7271, n_7272, n_7273, n_7274, n_7275, n_7276, n_7277, n_7278;
  wire n_7279, n_7280, n_7281, n_7282, n_7283, n_7287, n_7288, n_7289;
  wire n_7290, n_7291, n_7292, n_7293, n_7294, n_7295, n_7296, n_7297;
  wire n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304, n_7305;
  wire n_7306, n_7307, n_7308, n_7309, n_7310, n_7311, n_7312, n_7316;
  wire n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7325, n_7326;
  wire n_7327, n_7328, n_7332, n_7333, n_7334, n_7335, n_7336, n_7337;
  wire n_7339, n_7340, n_7341, n_7342, n_7343, n_7344, n_7345, n_7346;
  wire n_7347, n_7348, n_7349, n_7350, n_7351, n_7352, n_7354, n_7355;
  wire n_7356, n_7357, n_7358, n_7359, n_7360, n_7361, n_7362, n_7363;
  wire n_7364, n_7365, n_7366, n_7367, n_7368, n_7369, n_7370, n_7371;
  wire n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379, n_7380;
  wire n_7381, n_7384, n_7385, n_7386, n_7387, n_7388, n_7389, n_7390;
  wire n_7391, n_7392, n_7394, n_7395, n_7396, n_7398, n_7399, n_7402;
  wire n_7403, n_7404, n_7405, n_7406, n_7407, n_7408, n_7409, n_7410;
  wire n_7411, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418, n_7419;
  wire n_7420, n_7421, n_7422, n_7423, n_7425, n_7426, n_7427, n_7428;
  wire n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7437, n_7438;
  wire n_7439, n_7440, n_7441, n_7442, n_7443, n_7444, n_7445, n_7446;
  wire n_7447, n_7448, n_7449, n_7450, n_7451, n_7452, n_7453, n_7454;
  wire n_7455, n_7456, n_7457, n_7458, n_7459, n_7460, n_7461, n_7462;
  wire n_7463, n_7464, n_7465, n_7466, n_7467, n_7468, n_7469, n_7470;
  wire n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477, n_7478;
  wire n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485, n_7486;
  wire n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494;
  wire n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502;
  wire n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510;
  wire n_7511, n_7512, n_7513, n_7514, n_7515, n_7516, n_7517, n_7518;
  wire n_7519, n_7520, n_7521, n_7522, n_7523, n_7524, n_7525, n_7526;
  wire n_7527, n_7528, n_7529, n_7530, n_7531, n_7532, n_7533, n_7534;
  wire n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541, n_7542;
  wire n_7543, n_7544, n_7545, n_7546, n_7547, n_7548, n_7549, n_7550;
  wire n_7551, n_7552, n_7553, n_7554, n_7555, n_7556, n_7557, n_7558;
  wire n_7559, n_7560, n_7561, n_7562, n_7563, n_7564, n_7565, n_7566;
  wire n_7567, n_7568, n_7569, n_7570, n_7571, n_7572, n_7573, n_7574;
  wire n_7575, n_7576, n_7577, n_7578, n_7579, n_7580, n_7581, n_7582;
  wire n_7583, n_7584, n_7585, n_7586, n_7587, n_7588, n_7589, n_7591;
  wire n_7592, n_7593, n_7594, n_7595, n_7596, n_7597, n_7599, n_7600;
  wire n_7601, n_7602, n_7603, n_7604, n_7605, n_7606, n_7607, n_7608;
  wire n_7609, n_7610, n_7611, n_7612, n_7613, n_7614, n_7615, n_7617;
  wire n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625;
  wire n_7627, n_7628, n_7629, n_7630, n_7631, n_7632, n_7633, n_7634;
  wire n_7636, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643, n_7644;
  wire n_7645, n_7646, n_7647, n_7648, n_7649, n_7650, n_7651, n_7652;
  wire n_7653, n_7654, n_7655, n_7656, n_7658, n_7659, n_7660, n_7662;
  wire n_7663, n_7664, n_7665, n_7666, n_7667, n_7668, n_7669, n_7670;
  wire n_7671, n_7672, n_7675, n_7676, n_7677, n_7678, n_7679, n_7680;
  wire n_7681, n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7688;
  wire n_7689, n_7690, n_7691, n_7692, n_7693, n_7694, n_7697, n_7698;
  wire n_7699, n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, n_7708;
  wire n_7709, n_7710, n_7711, n_7712, n_7713, n_7714, n_7715, n_7718;
  wire n_7719, n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7726;
  wire n_7727, n_7728, n_7729, n_7730, n_7731, n_7732, n_7733, n_7734;
  wire n_7735, n_7736, n_7737, n_7738, n_7739, n_7740, n_7741, n_7742;
  wire n_7743, n_7744, n_7745, n_7746, n_7747, n_7748, n_7749, n_7750;
  wire n_7751, n_7752, n_7753, n_7754, n_7755, n_7756, n_7757, n_7758;
  wire n_7759, n_7760, n_7761, n_7762, n_7763, n_7764, n_7765, n_7766;
  wire n_7767, n_7768, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774;
  wire n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781, n_7782;
  wire n_7783, n_7784, n_7785, n_7786, n_7787, n_7788, n_7789, n_7790;
  wire n_7791, n_7792, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798;
  wire n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7807, n_7808;
  wire n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816;
  wire n_7817, n_7818, n_7819, n_7820, n_7821, n_7822, n_7823, n_7824;
  wire n_7825, n_7826, n_7830, n_7831, n_7832, n_7833, n_7834, n_7835;
  wire n_7836, n_7837, n_7838, n_7839, n_7840, n_7841, n_7842, n_7844;
  wire n_7846, n_7847, n_7848, n_7849, n_7850, n_7851, n_7852, n_7853;
  wire n_7854, n_7855, n_7856, n_7859, n_7860, n_7861, n_7862, n_7863;
  wire n_7864, n_7865, n_7866, n_7867, n_7868, n_7869, n_7870, n_7871;
  wire n_7872, n_7873, n_7874, n_7875, n_7876, n_7877, n_7878, n_7879;
  wire n_7880, n_7881, n_7882, n_7883, n_7884, n_7885, n_7886, n_7887;
  wire n_7888, n_7889, n_7890, n_7891, n_7892, n_7893, n_7894, n_7895;
  wire n_7898, n_7899, n_7900, n_7901, n_7902, n_7903, n_7904, n_7905;
  wire n_7906, n_7907, n_7908, n_7909, n_7910, n_7911, n_7912, n_7913;
  wire n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920, n_7921;
  wire n_7922, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928, n_7929;
  wire n_7930, n_7931, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937;
  wire n_7938, n_7939, n_7940, n_7941, n_7944, n_7945, n_7946, n_7947;
  wire n_7948, n_7949, n_7950, n_7951, n_7952, n_7953, n_7954, n_7955;
  wire n_7956, n_7957, n_7958, n_7959, n_7960, n_7961, n_7962, n_7963;
  wire n_7964, n_7965, n_7966, n_7967, n_7968, n_7969, n_7970, n_7971;
  wire n_7972, n_7973, n_7974, n_7975, n_7977, n_7978, n_7979, n_7980;
  wire n_7981, n_7982, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988;
  wire n_7989, n_7990, n_7991, n_7992, n_7993, n_7994, n_7995, n_7996;
  wire n_7997, n_7998, n_7999, n_8000, n_8001, n_8002, n_8003, n_8004;
  wire n_8005, n_8006, n_8007, n_8008, n_8009, n_8010, n_8011, n_8012;
  wire n_8013, n_8014, n_8015, n_8016, n_8017, n_8018, n_8019, n_8020;
  wire n_8021, n_8022, n_8023, n_8024, n_8025, n_8026, n_8027, n_8028;
  wire n_8029, n_8030, n_8031, n_8032, n_8033, n_8034, n_8035, n_8036;
  wire n_8037, n_8038, n_8039, n_8040, n_8041, n_8042, n_8043, n_8044;
  wire n_8045, n_8046, n_8047, n_8048, n_8049, n_8050, n_8051, n_8052;
  wire n_8053, n_8054, n_8055, n_8056, n_8057, n_8058, n_8059, n_8060;
  wire n_8061, n_8062, n_8063, n_8064, n_8065, n_8066, n_8067, n_8068;
  wire n_8069, n_8070, n_8071, n_8072, n_8073, n_8074, n_8075, n_8076;
  wire n_8077, n_8078, n_8079, n_8080, n_8081, n_8082, n_8083, n_8084;
  wire n_8085, n_8086, n_8087, n_8088, n_8089, n_8090, n_8091, n_8092;
  wire n_8093, n_8094, n_8095, n_8096, n_8097, n_8098, n_8099, n_8100;
  wire n_8101, n_8102, n_8103, n_8104, n_8105, n_8106, n_8107, n_8108;
  wire n_8109, n_8110, n_8111, n_8112, n_8113, n_8114, n_8115, n_8116;
  wire n_8117, n_8118, n_8119, n_8120, n_8121, n_8122, n_8123, n_8124;
  wire n_8125, n_8126, n_8127, n_8128, n_8129, n_8130, n_8131, n_8134;
  wire n_8135, n_8136, n_8139, n_8140, n_8141, n_8142, n_8143, n_8144;
  wire n_8145, n_8146, n_8147, n_8148, n_8149, n_8150, n_8151, n_8152;
  wire n_8153, n_8154, n_8155, n_8156, n_8157, n_8158, n_8159, n_8160;
  wire n_8161, n_8162, n_8163, n_8164, n_8165, n_8166, n_8167, n_8168;
  wire n_8169, n_8170, n_8171, n_8172, n_8173, n_8174, n_8175, n_8176;
  wire n_8177, n_8178, n_8179, n_8180, n_8181, n_8182, n_8183, n_8184;
  wire n_8185, n_8186, n_8187, n_8188, n_8189, n_8190, n_8191, n_8192;
  wire n_8193, n_8194, n_8195, n_8196, n_8197, n_8198, n_8199, n_8200;
  wire n_8201, n_8202, n_8203, n_8204, n_8205, n_8206, n_8207, n_8208;
  wire n_8209, n_8210, n_8211, n_8212, n_8213, n_8214, n_8215, n_8216;
  wire n_8217, n_8218, n_8219, n_8220, n_8221, n_8222, n_8223, n_8224;
  wire n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8231, n_8232;
  wire n_8233, n_8234, n_8235, n_8236, n_8237, n_8238, n_8239, n_8240;
  wire n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248;
  wire n_8249, n_8250, n_8251, n_8252, n_8253, n_8254, n_8255, n_8256;
  wire n_8257, n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264;
  wire n_8265, n_8266, n_8267, n_8268, n_8269, n_8270, n_8271, n_8272;
  wire n_8273, n_8274, n_8275, n_8276, n_8277, n_8278, n_8279, n_8280;
  wire n_8281, n_8282, n_8283, n_8284, n_8285, n_8286, n_8287, n_8288;
  wire n_8289, n_8290, n_8291, n_8292, n_8293, n_8294, n_8295, n_8296;
  wire n_8297, n_8298, n_8299, n_8300, n_8301, n_8302, n_8303, n_8304;
  wire n_8305, n_8306, n_8307, n_8308, n_8309, n_8310, n_8311, n_8312;
  wire n_8313, n_8314, n_8315, n_8316, n_8317, n_8318, n_8319, n_8320;
  wire n_8321, n_8322, n_8323, n_8324, n_8325, n_8326, n_8327, n_8328;
  wire n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335, n_8336;
  wire n_8337, n_8338, n_8339, n_8340, n_8341, n_8342, n_8343, n_8344;
  wire n_8345, n_8346, n_8347, n_8348, n_8349, n_8350, n_8351, n_8352;
  wire n_8353, n_8354, n_8355, n_8356, n_8357, n_8358, n_8359, n_8360;
  wire n_8361, n_8362, n_8363, n_8364, n_8365, n_8366, n_8367, n_8368;
  wire n_8369, n_8370, n_8371, n_8372, n_8373, n_8374, n_8375, n_8376;
  wire n_8377, n_8378, n_8379, n_8380, n_8381, n_8382, n_8383, n_8384;
  wire n_8385, n_8386, n_8387, n_8388, n_8389, n_8390, n_8391, n_8392;
  wire n_8393, n_8394, n_8395, n_8396, n_8397, n_8398, n_8399, n_8400;
  wire n_8401, n_8402, n_8403, n_8404, n_8405, n_8406, n_8407, n_8408;
  wire n_8409, n_8410, n_8411, n_8412, n_8413, n_8414, n_8415, n_8416;
  wire n_8417, n_8418, n_8419, n_8420, n_8421, n_8422, n_8423, n_8424;
  wire n_8425, n_8426, n_8427, n_8428, n_8429, n_8430, n_8431, n_8432;
  wire n_8433, n_8434, n_8435, n_8436, n_8437, n_8438, n_8439, n_8440;
  wire n_8441, n_8442, n_8443, n_8444, n_8445, n_8446, n_8447, n_8448;
  wire n_8449, n_8450, n_8451, n_8452, n_8453, n_8454, n_8455, n_8456;
  wire n_8457, n_8458, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464;
  wire n_8465, n_8466, n_8467, n_8468, n_8469, n_8470, n_8471, n_8472;
  wire n_8473, n_8474, n_8475, n_8476, n_8477, n_8478, n_8479, n_8480;
  wire n_8481, n_8482, n_8483, n_8484, n_8485, n_8486, n_8487, n_8488;
  wire n_8489, n_8490, n_8491, n_8492, n_8493, n_8494, n_8495, n_8496;
  wire n_8497, n_8498, n_8499, n_8500, n_8501, n_8502, n_8503, n_8504;
  wire n_8505, n_8506, n_8507, n_8508, n_8509, n_8510, n_8511, n_8512;
  wire n_8513, n_8514, n_8515, n_8516, n_8517, n_8518, n_8519, n_8520;
  wire n_8521, n_8522, n_8523, n_8524, n_8525, n_8526, n_8527, n_8528;
  wire n_8529, n_8530, n_8531, n_8532, n_8533, n_8534, n_8535, n_8536;
  wire n_8537, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544;
  wire n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552;
  wire n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560;
  wire n_8561, n_8562, n_8563, n_8564, n_8565, n_8566, n_8567, n_8568;
  wire n_8569, n_8570, n_8571, n_8572, n_8573, n_8574, n_8575, n_8576;
  wire n_8577, n_8578, n_8579, n_8580, n_8581, n_8582, n_8583, n_8584;
  wire n_8585, n_8586, n_8587, n_8588, n_8589, n_8590, n_8591, n_8592;
  wire n_8593, n_8594, n_8595, n_8596, n_8597, n_8598, n_8599, n_8600;
  wire n_8601, n_8602, n_8603, n_8604, n_8605, n_8606, n_8607, n_8608;
  wire n_8609, n_8610, n_8611, n_8612, n_8613, n_8614, n_8615, n_8616;
  wire n_8617, n_8618, n_8619, n_8620, n_8621, n_8622, n_8623, n_8624;
  wire n_8625, n_8626, n_8627, n_8628, n_8629, n_8630, n_8631, n_8632;
  wire n_8633, n_8634, n_8635, n_8636, n_8637, n_8638, n_8639, n_8640;
  wire n_8641, n_8642, n_8643, n_8644, n_8645, n_8646, n_8647, n_8648;
  wire n_8649, n_8650, n_8651, n_8652, n_8653, n_8654, n_8655, n_8656;
  wire n_8657, n_8658, n_8659, n_8660, n_8661, n_8662, n_8663, n_8664;
  wire n_8665, n_8666, n_8667, n_8668, n_8669, n_8672, n_8673, n_8674;
  wire n_8675, n_8676, n_8677, n_8678, n_8679, n_8680, n_8681, n_8682;
  wire n_8683, n_8684, n_8685, n_8686, n_8687, n_8688, n_8689, n_8690;
  wire n_8691, n_8692, n_8693, n_8694, n_8695, n_8696, n_8697, n_8698;
  wire n_8701, n_8702, n_8703, n_8704, n_8705, n_8708, n_8709, n_8711;
  wire n_8712, n_8713, n_8714, n_8715, n_8716, n_8717, n_8718, n_8719;
  wire n_8720, n_8721, n_8722, n_8723, n_8724, n_8725, n_8726, n_8727;
  wire n_8728, n_8729, n_8730, n_8731, n_8732, n_8733, n_8734, n_8735;
  wire n_8736, n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743;
  wire n_8744, n_8745, n_8746, n_8747, n_8749, n_8750, n_8751, n_8752;
  wire n_8753, n_8754, n_8755, n_8757, n_8758, n_8759, n_8760, n_8761;
  wire n_8763, n_8764, n_8765, n_8766, n_8767, n_8768, n_8769, n_8770;
  wire n_8771, n_8772, n_8773, n_8774, n_8775, n_8776, n_8777, n_8778;
  wire n_8779, n_8780, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786;
  wire n_8787, n_8788, n_8789, n_8790, n_8791, n_8792, n_8793, n_8794;
  wire n_8795, n_8796, n_8797, n_8798, n_8799, n_8800, n_8801, n_8802;
  wire n_8803, n_8804, n_8805, n_8806, n_8807, n_8808, n_8812, n_8813;
  wire n_8814, n_8815, n_8816, n_8817, n_8818, n_8819, n_8820, n_8821;
  wire n_8822, n_8823, n_8824, n_8825, n_8826, n_8827, n_8828, n_8829;
  wire n_8831, n_8832, n_8833, n_8834, n_8835, n_8836, n_8837, n_8838;
  wire n_8839, n_8840, n_8841, n_8842, n_8843, n_8844, n_8845, n_8846;
  wire n_8847, n_8848, n_8849, n_8850, n_8851, n_8852, n_8853, n_8854;
  wire n_8855, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861, n_8862;
  wire n_8863, n_8864, n_8865, n_8866, n_8867, n_8868, n_8869, n_8870;
  wire n_8871, n_8872, n_8873, n_8874, n_8875, n_8876, n_8877, n_8878;
  wire n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888, n_8889;
  wire n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896, n_8897;
  wire n_8898, n_8899, n_8901, n_8904, n_8905, n_8906, n_8907, n_8908;
  wire n_8909, n_8910, n_8911, n_8912, n_8913, n_8914, n_8915, n_8916;
  wire n_8917, n_8918, n_8919, n_8920, n_8921, n_8922, n_8925, n_8926;
  wire n_8927, n_8928, n_8929, n_8930, n_8931, n_8932, n_8933, n_8934;
  wire n_8935, n_8937, n_8938, n_8939, n_8940, n_8941, n_8942, n_8943;
  wire n_8944, n_8945, n_8946, n_8947, n_8948, n_8949, n_8950, n_8951;
  wire n_8952, n_8953, n_8954, n_8955, n_8956, n_8957, n_8958, n_8959;
  wire n_8960, n_8961, n_8962, n_8963, n_8964, n_8965, n_8966, n_8967;
  wire n_8968, n_8969, n_8970, n_8971, n_8972, n_8973, n_8974, n_8975;
  wire n_8976, n_8977, n_8978, n_8979, n_8980, n_8981, n_8982, n_8983;
  wire n_8984, n_8985, n_8986, n_8987, n_8988, n_8989, n_8990, n_8991;
  wire n_8992, n_8993, n_8994, n_8995, n_8996, n_8997, n_8998, n_8999;
  wire n_9000, n_9001, n_9002, n_9003, n_9004, n_9005, n_9006, n_9007;
  wire n_9011, n_9012, n_9013, n_9014, n_9015, n_9016, n_9017, n_9018;
  wire n_9019, n_9020, n_9021, n_9022, n_9023, n_9024, n_9025, n_9026;
  wire n_9027, n_9028, n_9029, n_9030, n_9031, n_9032, n_9033, n_9034;
  wire n_9035, n_9036, n_9037, n_9038, n_9039, n_9043, n_9044, n_9045;
  wire n_9046, n_9047, n_9048, n_9049, n_9050, n_9051, n_9052, n_9053;
  wire n_9054, n_9055, n_9056, n_9057, n_9058, n_9059, n_9060, n_9061;
  wire n_9062, n_9063, n_9064, n_9065, n_9066, n_9067, n_9068, n_9069;
  wire n_9070, n_9071, n_9072, n_9073, n_9074, n_9075, n_9076, n_9077;
  wire n_9080, n_9081, n_9082, n_9083, n_9084, n_9085, n_9086, n_9087;
  wire n_9088, n_9089, n_9090, n_9091, n_9092, n_9093, n_9094, n_9095;
  wire n_9096, n_9097, n_9098, n_9099, n_9100, n_9101, n_9102, n_9103;
  wire n_9104, n_9105, n_9106, n_9107, n_9109, n_9110, n_9111, n_9112;
  wire n_9113, n_9114, n_9116, n_9117, n_9118, n_9119, n_9120, n_9121;
  wire n_9122, n_9123, n_9124, n_9125, n_9126, n_9127, n_9128, n_9129;
  wire n_9131, n_9132, n_9133, n_9134, n_9135, n_9136, n_9137, n_9138;
  wire n_9139, n_9141, n_9142, n_9143, n_9144, n_9145, n_9146, n_9147;
  wire n_9148, n_9149, n_9150, n_9151, n_9152, n_9153, n_9154, n_9155;
  wire n_9156, n_9157, n_9158, n_9159, n_9160, n_9161, n_9162, n_9163;
  wire n_9164, n_9165, n_9166, n_9167, n_9168, n_9169, n_9170, n_9171;
  wire n_9172, n_9173, n_9174, n_9175, n_9176, n_9177, n_9178, n_9179;
  wire n_9180, n_9181, n_9183, n_9184, n_9185, n_9186, n_9187, n_9188;
  wire n_9189, n_9190, n_9192, n_9193, n_9194, n_9195, n_9196, n_9197;
  wire n_9198, n_9199, n_9200, n_9201, n_9202, n_9203, n_9204, n_9205;
  wire n_9206, n_9207, n_9208, n_9209, n_9210, n_9211, n_9212, n_9213;
  wire n_9214, n_9215, n_9216, n_9217, n_9218, n_9219, n_9220, n_9223;
  wire n_9224, n_9225, n_9226, n_9227, n_9228, n_9229, n_9230, n_9231;
  wire n_9232, n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9239;
  wire n_9240, n_9241, n_9242, n_9243, n_9244, n_9245, n_9246, n_9249;
  wire n_9250, n_9251, n_9252, n_9253, n_9254, n_9255, n_9256, n_9257;
  wire n_9258, n_9259, n_9260, n_9261, n_9262, n_9263, n_9264, n_9265;
  wire n_9266, n_9267, n_9268, n_9269, n_9270, n_9271, n_9272, n_9273;
  wire n_9274, n_9275, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281;
  wire n_9282, n_9283, n_9284, n_9285, n_9286, n_9287, n_9288, n_9289;
  wire n_9290, n_9291, n_9292, n_9293, n_9294, n_9295, n_9296, n_9297;
  wire n_9298, n_9299, n_9300, n_9301, n_9302, n_9303, n_9304, n_9305;
  wire n_9306, n_9307, n_9308, n_9309, n_9310, n_9311, n_9312, n_9313;
  wire n_9314, n_9315, n_9316, n_9317, n_9318, n_9319, n_9320, n_9321;
  wire n_9322, n_9323, n_9324, n_9325, n_9326, n_9327, n_9329, n_9330;
  wire n_9331, n_9332, n_9333, n_9334, n_9335, n_9336, n_9337, n_9338;
  wire n_9339, n_9340, n_9341, n_9343, n_9344, n_9345, n_9346, n_9347;
  wire n_9348, n_9349, n_9350, n_9351, n_9352, n_9353, n_9354, n_9355;
  wire n_9356, n_9357, n_9358, n_9359, n_9361, n_9362, n_9363, n_9364;
  wire n_9365, n_9366, n_9367, n_9368, n_9369, n_9370, n_9371, n_9372;
  wire n_9373, n_9374, n_9375, n_9376, n_9377, n_9378, n_9379, n_9380;
  wire n_9381, n_9382, n_9383, n_9384, n_9385, n_9387, n_9389, n_9390;
  wire n_9391, n_9392, n_9393, n_9394, n_9395, n_9396, n_9397, n_9398;
  wire n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405, n_9406;
  wire n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413, n_9414;
  wire n_9415, n_9416, n_9417, n_9418, n_9419, n_9420, n_9421, n_9422;
  wire n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430;
  wire n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438;
  wire n_9439, n_9440, n_9441, n_9442, n_9443, n_9444, n_9445, n_9446;
  wire n_9447, n_9448, n_9449, n_9450, n_9451, n_9452, n_9453, n_9454;
  wire n_9455, n_9456, n_9457, n_9458, n_9459, n_9460, n_9461, n_9462;
  wire n_9465, n_9468, n_9469, n_9470, n_9471, n_9472, n_9473, n_9474;
  wire n_9475, n_9476, n_9477, n_9478, n_9479, n_9480, n_9481, n_9482;
  wire n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489, n_9490;
  wire n_9491, n_9492, n_9493, n_9494, n_9495, n_9496, n_9499, n_9500;
  wire n_9501, n_9502, n_9503, n_9504, n_9505, n_9506, n_9507, n_9508;
  wire n_9509, n_9510, n_9511, n_9512, n_9513, n_9514, n_9515, n_9516;
  wire n_9517, n_9518, n_9519, n_9520, n_9521, n_9522, n_9523, n_9524;
  wire n_9525, n_9526, n_9527, n_9528, n_9529, n_9530, n_9531, n_9532;
  wire n_9533, n_9534, n_9535, n_9536, n_9537, n_9538, n_9539, n_9540;
  wire n_9541, n_9542, n_9543, n_9544, n_9545, n_9546, n_9547, n_9548;
  wire n_9549, n_9550, n_9551, n_9552, n_9553, n_9554, n_9555, n_9556;
  wire n_9557, n_9558, n_9560, n_9562, n_9563, n_9564, n_9565, n_9566;
  wire n_9567, n_9568, n_9569, n_9570, n_9571, n_9572, n_9573, n_9574;
  wire n_9575, n_9576, n_9577, n_9578, n_9579, n_9580, n_9581, n_9582;
  wire n_9583, n_9584, n_9585, n_9586, n_9587, n_9588, n_9589, n_9590;
  wire n_9591, n_9592, n_9593, n_9594, n_9595, n_9596, n_9597, n_9598;
  wire n_9599, n_9600, n_9601, n_9602, n_9603, n_9604, n_9605, n_9606;
  wire n_9607, n_9608, n_9609, n_9610, n_9611, n_9612, n_9613, n_9614;
  wire n_9615, n_9616, n_9617, n_9618, n_9619, n_9620, n_9621, n_9622;
  wire n_9623, n_9624, n_9625, n_9626, n_9627, n_9628, n_9629, n_9630;
  wire n_9631, n_9632, n_9633, n_9634, n_9635, n_9636, n_9637, n_9638;
  wire n_9639, n_9640, n_9641, n_9642, n_9643, n_9644, n_9645, n_9646;
  wire n_9647, n_9648, n_9649, n_9650, n_9651, n_9652, n_9653, n_9654;
  wire n_9655, n_9656, n_9657, n_9658, n_9659, n_9660, n_9661, n_9662;
  wire n_9663, n_9664, n_9665, n_9666, n_9667, n_9668, n_9669, n_9670;
  wire n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677, n_9678;
  wire n_9679, n_9680, n_9681, n_9682, n_9683, n_9684, n_9685, n_9686;
  wire n_9687, n_9688, n_9689, n_9690, n_9691, n_9692, n_9693, n_9694;
  wire n_9695, n_9696, n_9697, n_9698, n_9701, n_9702, n_9704, n_9706;
  wire n_9708, n_9710, n_9712, n_9715, n_9716, n_9717, n_9718, n_9719;
  wire n_9720, n_9721, n_9722, n_9723, n_9724, n_9725, n_9726, n_9727;
  wire n_9728, n_9729, n_9730, n_9731, n_9732, n_9733, n_9734, n_9735;
  wire n_9736, n_9737, n_9738, n_9739, n_9740, n_9741, n_9742, n_9743;
  wire n_9744, n_9745, n_9746, n_9747, n_9748, n_9749, n_9750, n_9751;
  wire n_9752, n_9753, n_9754, n_9755, n_9756, n_9757, n_9758, n_9759;
  wire n_9760, n_9761, n_9762, n_9763, n_9764, n_9765, n_9766, n_9767;
  wire n_9768, n_9769, n_9770, n_9771, n_9772, n_9773, n_9774, n_9775;
  wire n_9776, n_9777, n_9778, n_9779, n_9780, n_9781, n_9782, n_9783;
  wire n_9784, n_9785, n_9786, n_9787, n_9788, n_9789, n_9790, n_9791;
  wire n_9792, n_9793, n_9794, n_9795, n_9796, n_9797, n_9798, n_9799;
  wire n_9800, n_9801, n_9802, n_9803, n_9804, n_9805, n_9806, n_9807;
  wire n_9808, n_9809, n_9810, n_9811, n_9812, n_9813, n_9814, n_9815;
  wire n_9816, n_9817, n_9818, n_9819, n_9820, n_9821, n_9822, n_9823;
  wire n_9824, n_9825, n_9826, n_9827, n_9828, n_9829, n_9830, n_9831;
  wire n_9832, n_9833, n_9834, n_9835, n_9836, n_9837, n_9838, n_9839;
  wire n_9840, n_9841, n_9842, n_9843, n_9844, n_9845, n_9846, n_9847;
  wire n_9848, n_9849, n_9850, n_9851, n_9852, n_9853, n_9854, n_9855;
  wire n_9856, n_9857, n_9858, n_9859, n_9860, n_9861, n_9862, n_9863;
  wire n_9864, n_9865, n_9866, n_9867, n_9868, n_9869, n_9870, n_9871;
  wire n_9872, n_9873, n_9874, n_9875, n_9876, n_9877, n_9878, n_9879;
  wire n_9880, n_9881, n_9882, n_9883, n_9884, n_9885, n_9886, n_9887;
  wire n_9888, n_9889, n_9890, n_9891, n_9892, n_9893, n_9894, n_9895;
  wire n_9896, n_9897, n_9898, n_9899, n_9900, n_9901, n_9902, n_9903;
  wire n_9904, n_9905, n_9906, n_9907, n_9908, n_9909, n_9910, n_9911;
  wire n_9912, n_9913, n_9914, n_9915, n_9916, n_9917, n_9918, n_9919;
  wire n_9920, n_9921, n_9922, n_9923, n_9924, n_9925, n_9926, n_9927;
  wire n_9928, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937, n_9938;
  wire n_9939, n_9940, n_9941, n_9942, n_9943, n_9944, n_9945, n_9948;
  wire n_9949, n_9950, n_9951, n_9952, n_9953, n_9954, n_9955, n_9956;
  wire n_9957, n_9958, n_9959, n_9960, n_9961, n_9962, n_9963, n_9964;
  wire n_9965, n_9966, n_9967, n_9968, n_9969, n_9970, n_9971, n_9972;
  wire n_9973, n_9977, n_9978, n_9979, n_9980, n_9981, n_9982, n_9983;
  wire n_9984, n_9985, n_9986, n_9987, n_9988, n_9989, n_9990, n_9991;
  wire n_9992, n_9993, n_9994, n_9995, n_9996, n_9997, n_9998, n_9999;
  wire n_10000, n_10001, n_10002, n_10003, n_10004, n_10005, n_10006,
       n_10007;
  wire n_10008, n_10009, n_10010, n_10011, n_10012, n_10013, n_10014,
       n_10015;
  wire n_10016, n_10017, n_10020, n_10021, n_10022, n_10023, n_10024,
       n_10025;
  wire n_10027, n_10028, n_10029, n_10030, n_10031, n_10032, n_10033,
       n_10034;
  wire n_10035, n_10036, n_10037, n_10038, n_10039, n_10040, n_10041,
       n_10042;
  wire n_10043, n_10044, n_10045, n_10046, n_10047, n_10048, n_10049,
       n_10050;
  wire n_10051, n_10052, n_10053, n_10054, n_10055, n_10056, n_10057,
       n_10058;
  wire n_10059, n_10060, n_10061, n_10062, n_10063, n_10064, n_10065,
       n_10066;
  wire n_10067, n_10068, n_10069, n_10070, n_10071, n_10072, n_10073,
       n_10074;
  wire n_10075, n_10076, n_10077, n_10078, n_10079, n_10080, n_10081,
       n_10082;
  wire n_10083, n_10084, n_10085, n_10086, n_10087, n_10088, n_10089,
       n_10090;
  wire n_10091, n_10092, n_10093, n_10094, n_10095, n_10096, n_10097,
       n_10098;
  wire n_10099, n_10100, n_10101, n_10102, n_10103, n_10104, n_10105,
       n_10106;
  wire n_10107, n_10108, n_10109, n_10110, n_10111, n_10112, n_10113,
       n_10114;
  wire n_10115, n_10116, n_10117, n_10118, n_10119, n_10120, n_10121,
       n_10122;
  wire n_10123, n_10124, n_10125, n_10126, n_10127, n_10128, n_10129,
       n_10130;
  wire n_10131, n_10132, n_10133, n_10134, n_10135, n_10136, n_10137,
       n_10138;
  wire n_10139, n_10140, n_10141, n_10142, n_10143, n_10144, n_10145,
       n_10146;
  wire n_10147, n_10148, n_10149, n_10150, n_10151, n_10152, n_10153,
       n_10154;
  wire n_10155, n_10156, n_10157, n_10158, n_10159, n_10160, n_10161,
       n_10162;
  wire n_10163, n_10164, n_10165, n_10168, n_10169, n_10170, n_10171,
       n_10172;
  wire n_10173, n_10174, n_10175, n_10176, n_10177, n_10178, n_10179,
       n_10180;
  wire n_10181, n_10182, n_10183, n_10184, n_10185, n_10186, n_10187,
       n_10188;
  wire n_10189, n_10190, n_10191, n_10192, n_10193, n_10194, n_10195,
       n_10196;
  wire n_10197, n_10198, n_10199, n_10200, n_10201, n_10202, n_10203,
       n_10204;
  wire n_10205, n_10206, n_10207, n_10208, n_10209, n_10210, n_10211,
       n_10212;
  wire n_10213, n_10214, n_10215, n_10216, n_10217, n_10218, n_10219,
       n_10220;
  wire n_10221, n_10222, n_10223, n_10224, n_10225, n_10226, n_10227,
       n_10228;
  wire n_10229, n_10230, n_10231, n_10232, n_10233, n_10236, n_10237,
       n_10238;
  wire n_10239, n_10240, n_10241, n_10242, n_10243, n_10244, n_10245,
       n_10246;
  wire n_10247, n_10248, n_10249, n_10250, n_10251, n_10252, n_10253,
       n_10254;
  wire n_10255, n_10256, n_10257, n_10258, n_10259, n_10260, n_10261,
       n_10262;
  wire n_10263, n_10264, n_10265, n_10266, n_10267, n_10268, n_10269,
       n_10270;
  wire n_10271, n_10272, n_10273, n_10277, n_10278, n_10279, n_10280,
       n_10281;
  wire n_10282, n_10283, n_10284, n_10287, n_10288, n_10289, n_10290,
       n_10291;
  wire n_10292, n_10293, n_10294, n_10295, n_10296, n_10299, n_10300,
       n_10301;
  wire n_10302, n_10303, n_10304, n_10305, n_10306, n_10307, n_10308,
       n_10309;
  wire n_10310, n_10311, n_10312, n_10313, n_10314, n_10315, n_10316,
       n_10317;
  wire n_10318, n_10319, n_10320, n_10321, n_10322, n_10323, n_10324,
       n_10325;
  wire n_10326, n_10327, n_10328, n_10329, n_10330, n_10331, n_10332,
       n_10333;
  wire n_10334, n_10335, n_10336, n_10337, n_10338, n_10339, n_10340,
       n_10341;
  wire n_10342, n_10343, n_10344, n_10345, n_10346, n_10347, n_10348,
       n_10349;
  wire n_10350, n_10351, n_10352, n_10353, n_10354, n_10355, n_10356,
       n_10357;
  wire n_10358, n_10359, n_10360, n_10361, n_10362, n_10365, n_10366,
       n_10367;
  wire n_10368, n_10369, n_10370, n_10371, n_10372, n_10373, n_10374,
       n_10375;
  wire n_10376, n_10377, n_10378, n_10379, n_10380, n_10381, n_10382,
       n_10383;
  wire n_10384, n_10385, n_10386, n_10387, n_10388, n_10389, n_10390,
       n_10391;
  wire n_10392, n_10393, n_10394, n_10395, n_10396, n_10397, n_10398,
       n_10399;
  wire n_10400, n_10401, n_10402, n_10403, n_10404, n_10405, n_10406,
       n_10407;
  wire n_10408, n_10409, n_10410, n_10411, n_10412, n_10413, n_10414,
       n_10415;
  wire n_10416, n_10417, n_10418, n_10419, n_10420, n_10421, n_10422,
       n_10423;
  wire n_10424, n_10425, n_10426, n_10427, n_10428, n_10429, n_10430,
       n_10431;
  wire n_10432, n_10433, n_10434, n_10437, n_10438, n_10439, n_10440,
       n_10441;
  wire n_10442, n_10443, n_10444, n_10445, n_10446, n_10447, n_10448,
       n_10449;
  wire n_10450, n_10451, n_10452, n_10456, n_10457, n_10458, n_10459,
       n_10460;
  wire n_10461, n_10462, n_10466, n_10467, n_10468, n_10469, n_10470,
       n_10471;
  wire n_10472, n_10473, n_10474, n_10479, n_10480, n_10481, n_10482,
       n_10483;
  wire n_10484, n_10485, n_10486, n_10487, n_10488, n_10489, n_10490,
       n_10491;
  wire n_10492, n_10493, n_10494, n_10495, n_10496, n_10497, n_10498,
       n_10499;
  wire n_10500, n_10501, n_10502, n_10503, n_10504, n_10505, n_10506,
       n_10507;
  wire n_10508, n_10509, n_10510, n_10511, n_10512, n_10513, n_10514,
       n_10515;
  wire n_10516, n_10517, n_10518, n_10519, n_10520, n_10521, n_10522,
       n_10523;
  wire n_10524, n_10525, n_10526, n_10529, n_10530, n_10531, n_10532,
       n_10533;
  wire n_10534, n_10535, n_10536, n_10537, n_10538, n_10541, n_10542,
       n_10543;
  wire n_10544, n_10545, n_10546, n_10547, n_10548, n_10549, n_10550,
       n_10551;
  wire n_10552, n_10553, n_10554, n_10555, n_10556, n_10557, n_10558,
       n_10559;
  wire n_10560, n_10561, n_10562, n_10563, n_10564, n_10565, n_10566,
       n_10567;
  wire n_10568, n_10569, n_10570, n_10571, n_10572, n_10577, n_10578,
       n_10579;
  wire n_10580, n_10581, n_10582, n_10586, n_10587, n_10588, n_10589,
       n_10590;
  wire n_10591, n_10592, n_10593, n_10594, n_10595, n_10596, n_10597,
       n_10598;
  wire n_10599, n_10600, n_10601, n_10602, n_10603, n_10604, n_10605,
       n_10606;
  wire n_10607, n_10608, n_10609, n_10610, n_10611, n_10612, n_10613,
       n_10614;
  wire n_10615, n_10616, n_10617, n_10618, n_10619, n_10620, n_10621,
       n_10622;
  wire n_10623, n_10624, n_10625, n_10626, n_10627, n_10628, n_10629,
       n_10630;
  wire n_10631, n_10632, n_10633, n_10634, n_10635, n_10636, n_10637,
       n_10638;
  wire n_10640, n_10641, n_10642, n_10643, n_10644, n_10645, n_10646,
       n_10647;
  wire n_10648, n_10649, n_10650, n_10651, n_10652, n_10653, n_10654,
       n_10655;
  wire n_10656, n_10657, n_10658, n_10660, n_10661, n_10662, n_10663,
       n_10664;
  wire n_10665, n_10666, n_10667, n_10668, n_10669, n_10670, n_10671,
       n_10672;
  wire n_10673, n_10674, n_10675, n_10676, n_10677, n_10678, n_10679,
       n_10680;
  wire n_10681, n_10682, n_10683, n_10684, n_10685, n_10688, n_10689,
       n_10690;
  wire n_10691, n_10692, n_10693, n_10694, n_10695, n_10696, n_10697,
       n_10698;
  wire n_10699, n_10700, n_10701, n_10702, n_10703, n_10704, n_10705,
       n_10706;
  wire n_10707, n_10708, n_10709, n_10710, n_10711, n_10712, n_10713,
       n_10714;
  wire n_10715, n_10716, n_10717, n_10718, n_10719, n_10720, n_10721,
       n_10722;
  wire n_10723, n_10724, n_10725, n_10726, n_10727, n_10728, n_10734,
       n_10735;
  wire n_10736, n_10737, n_10738, n_10739, n_10740, n_10741, n_10742,
       n_10743;
  wire n_10744, n_10745, n_10746, n_10747, n_10750, n_10751, n_10752,
       n_10753;
  wire n_10754, n_10755, n_10756, n_10757, n_10758, n_10759, n_10760,
       n_10761;
  wire n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768,
       n_10769;
  wire n_10770, n_10771, n_10772, n_10773, n_10774, n_10775, n_10776,
       n_10777;
  wire n_10778, n_10779, n_10780, n_10781, n_10782, n_10783, n_10784,
       n_10785;
  wire n_10786, n_10787, n_10788, n_10789, n_10790, n_10791, n_10792,
       n_10793;
  wire n_10794, n_10795, n_10796, n_10797, n_10798, n_10799, n_10800,
       n_10804;
  wire n_10805, n_10806, n_10807, n_10808, n_10809, n_10810, n_10811,
       n_10812;
  wire n_10813, n_10814, n_10815, n_10816, n_10817, n_10818, n_10819,
       n_10820;
  wire n_10821, n_10822, n_10823, n_10824, n_10825, n_10826, n_10827,
       n_10828;
  wire n_10829, n_10830, n_10831, n_10832, n_10833, n_10834, n_10835,
       n_10836;
  wire n_10837, n_10838, n_10839, n_10840, n_10841, n_10842, n_10843,
       n_10844;
  wire n_10845, n_10846, n_10847, n_10848, n_10849, n_10850, n_10851,
       n_10852;
  wire n_10853, n_10854, n_10855, n_10856, n_10857, n_10861, n_10862,
       n_10863;
  wire n_10864, n_10865, n_10866, n_10867, n_10868, n_10869, n_10870,
       n_10871;
  wire n_10872, n_10873, n_10874, n_10875, n_10876, n_10877, n_10878,
       n_10879;
  wire n_10880, n_10881, n_10882, n_10883, n_10884, n_10885, n_10886,
       n_10887;
  wire n_10888, n_10889, n_10890, n_10891, n_10892, n_10893, n_10894,
       n_10895;
  wire n_10896, n_10897, n_10898, n_10899, n_10900, n_10901, n_10902,
       n_10903;
  wire n_10904, n_10905, n_10908, n_10909, n_10910, n_10911, n_10912,
       n_10913;
  wire n_10914, n_10915, n_10916, n_10917, n_10918, n_10919, n_10920,
       n_10921;
  wire n_10922, n_10923, n_10924, n_10925, n_10926, n_10927, n_10928,
       n_10929;
  wire n_10930, n_10931, n_10932, n_10933, n_10934, n_10935, n_10936,
       n_10937;
  wire n_10938, n_10939, n_10940, n_10941, n_10942, n_10943, n_10944,
       n_10945;
  wire n_10946, n_10947, n_10948, n_10949, n_10950, n_10951, n_10952,
       n_10953;
  wire n_10954, n_10955, n_10959, n_10960, n_10961, n_10962, n_10963,
       n_10967;
  wire n_10968, n_10969, n_10970, n_10971, n_10972, n_10973, n_10974,
       n_10975;
  wire n_10976, n_10977, n_10978, n_10979, n_10980, n_10981, n_10982,
       n_10983;
  wire n_10984, n_10985, n_10986, n_10987, n_10988, n_10989, n_10990,
       n_10993;
  wire n_10994, n_10995, n_10996, n_10997, n_10998, n_10999, n_11000,
       n_11001;
  wire n_11002, n_11008, n_11009, n_11010, n_11011, n_11012, n_11013,
       n_11014;
  wire n_11015, n_11016, n_11017, n_11018, n_11020, n_11021, n_11022,
       n_11023;
  wire n_11024, n_11025, n_11026, n_11027, n_11028, n_11029, n_11030,
       n_11031;
  wire n_11032, n_11033, n_11034, n_11037, n_11038, n_11039, n_11040,
       n_11041;
  wire n_11042, n_11043, n_11044, n_11045, n_11046, n_11047, n_11048,
       n_11049;
  wire n_11050, n_11051, n_11052, n_11053, n_11054, n_11055, n_11056,
       n_11057;
  wire n_11058, n_11059, n_11060, n_11061, n_11062, n_11063, n_11064,
       n_11065;
  wire n_11066, n_11067, n_11068, n_11069, n_11070, n_11071, n_11072,
       n_11073;
  wire n_11074, n_11075, n_11076, n_11077, n_11078, n_11079, n_11080,
       n_11081;
  wire n_11082, n_11083, n_11084, n_11085, n_11086, n_11089, n_11090,
       n_11091;
  wire n_11092, n_11093, n_11094, n_11095, n_11096, n_11097, n_11098,
       n_11101;
  wire n_11102, n_11103, n_11104, n_11105, n_11106, n_11107, n_11108,
       n_11109;
  wire n_11110, n_11111, n_11113, n_11114, n_11115, n_11116, n_11117,
       n_11118;
  wire n_11119, n_11120, n_11121, n_11122, n_11123, n_11124, n_11125,
       n_11126;
  wire n_11127, n_11128, n_11129, n_11130, n_11131, n_11132, n_11133,
       n_11134;
  wire n_11135, n_11136, n_11137, n_11138, n_11139, n_11140, n_11141,
       n_11142;
  wire n_11143, n_11144, n_11145, n_11146, n_11147, n_11148, n_11149,
       n_11150;
  wire n_11151, n_11152, n_11153, n_11154, n_11155, n_11156, n_11157,
       n_11158;
  wire n_11159, n_11160, n_11161, n_11162, n_11163, n_11164, n_11165,
       n_11166;
  wire n_11167, n_11168, n_11169, n_11170, n_11171, n_11172, n_11173,
       n_11174;
  wire n_11175, n_11176, n_11177, n_11178, n_11179, n_11180, n_11181,
       n_11182;
  wire n_11183, n_11184, n_11185, n_11186, n_11187, n_11188, n_11189,
       n_11190;
  wire n_11191, n_11192, n_11193, n_11194, n_11195, n_11196, n_11197,
       n_11198;
  wire n_11199, n_11200, n_11201, n_11202, n_11203, n_11204, n_11205,
       n_11206;
  wire n_11207, n_11208, n_11209, n_11210, n_11211, n_11212, n_11213,
       n_11214;
  wire n_11215, n_11216, n_11217, n_11218, n_11219, n_11220, n_11221,
       n_11222;
  wire n_11223, n_11224, n_11225, n_11226, n_11227, n_11228, n_11229,
       n_11230;
  wire n_11231, n_11232, n_11233, n_11234, n_11235, n_11236, n_11237,
       n_11238;
  wire n_11239, n_11240, n_11241, n_11242, n_11243, n_11244, n_11245,
       n_11246;
  wire n_11247, n_11248, n_11249, n_11250, n_11251, n_11252, n_11253,
       n_11254;
  wire n_11255, n_11256, n_11257, n_11258, n_11259, n_11260, n_11261,
       n_11262;
  wire n_11263, n_11264, n_11265, n_11266, n_11267, n_11268, n_11269,
       n_11270;
  wire n_11271, n_11272, n_11273, n_11274, n_11275, n_11276, n_11277,
       n_11278;
  wire n_11279, n_11280, n_11281, n_11282, n_11283, n_11284, n_11285,
       n_11286;
  wire n_11287, n_11288, n_11289, n_11290, n_11291, n_11292, n_11293,
       n_11294;
  wire n_11295, n_11296, n_11297, n_11298, n_11299, n_11300, n_11301,
       n_11302;
  wire n_11303, n_11304, n_11305, n_11306, n_11307, n_11308, n_11309,
       n_11310;
  wire n_11311, n_11312, n_11313, n_11314, n_11315, n_11316, n_11317,
       n_11318;
  wire n_11319, n_11320, n_11321, n_11322, n_11323, n_11327, n_11328,
       n_11329;
  wire n_11330, n_11331, n_11332, n_11333, n_11334, n_11335, n_11336,
       n_11337;
  wire n_11338, n_11339, n_11340, n_11341, n_11342, n_11343, n_11344,
       n_11345;
  wire n_11346, n_11347, n_11348, n_11349, n_11350, n_11354, n_11355,
       n_11356;
  wire n_11357, n_11358, n_11359, n_11360, n_11361, n_11362, n_11363,
       n_11364;
  wire n_11365, n_11366, n_11367, n_11368, n_11369, n_11370, n_11374,
       n_11375;
  wire n_11376, n_11377, n_11378, n_11379, n_11380, n_11381, n_11382,
       n_11383;
  wire n_11384, n_11385, n_11386, n_11387, n_11388, n_11389, n_11390,
       n_11391;
  wire n_11392, n_11393, n_11395, n_11397, n_11398, n_11399, n_11401,
       n_11403;
  wire n_11405, n_11406, n_11407, n_11409, n_11412, n_11413, n_11415,
       n_11416;
  wire n_11417, n_11418, n_11420, n_11421, n_11422, n_11423, n_11424,
       n_11425;
  wire n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432,
       n_11433;
  wire n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440,
       n_11441;
  wire n_11442, n_11443, n_11444, n_11445, n_11446, n_11447, n_11448,
       n_11449;
  wire n_11450, n_11451, n_11452, n_11453, n_11454, n_11455, n_11456,
       n_11457;
  wire n_11458, n_11459, n_11460, n_11461, n_11462, n_11463, n_11464,
       n_11465;
  wire n_11466, n_11467, n_11468, n_11469, n_11470, n_11471, n_11472,
       n_11473;
  wire n_11474, n_11475, n_11476, n_11477, n_11478, n_11479, n_11480,
       n_11481;
  wire n_11482, n_11483, n_11484, n_11485, n_11486, n_11487, n_11488,
       n_11489;
  wire n_11490, n_11491, n_11492, n_11493, n_11494, n_11495, n_11496,
       n_11497;
  wire n_11498, n_11499, n_11500, n_11501, n_11502, n_11503, n_11504,
       n_11505;
  wire n_11506, n_11507, n_11508, n_11509, n_11510, n_11511, n_11512,
       n_11513;
  wire n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520,
       n_11521;
  wire n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528,
       n_11529;
  wire n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536,
       n_11537;
  wire n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544,
       n_11545;
  wire n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552,
       n_11553;
  wire n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560,
       n_11561;
  wire n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568,
       n_11569;
  wire n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576,
       n_11577;
  wire n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584,
       n_11585;
  wire n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592,
       n_11593;
  wire n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600,
       n_11601;
  wire n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11609,
       n_11610;
  wire n_11611, n_11612, n_11613, n_11614, n_11615, n_11616, n_11617,
       n_11618;
  wire n_11619, n_11620, n_11621, n_11622, n_11623, n_11624, n_11625,
       n_11626;
  wire n_11627, n_11628, n_11629, n_11630, n_11631, n_11632, n_11633,
       n_11634;
  wire n_11635, n_11636, n_11637, n_11638, n_11639, n_11640, n_11641,
       n_11642;
  wire n_11643, n_11644, n_11645, n_11646, n_11647, n_11648, n_11649,
       n_11650;
  wire n_11651, n_11652, n_11653, n_11654, n_11655, n_11656, n_11657,
       n_11658;
  wire n_11659, n_11660, n_11661, n_11662, n_11663, n_11664, n_11665,
       n_11667;
  wire n_11668, n_11669, n_11670, n_11671, n_11672, n_11673, n_11674,
       n_11675;
  wire n_11676, n_11677, n_11678, n_11679, n_11680, n_11681, n_11682,
       n_11683;
  wire n_11684, n_11685, n_11686, n_11687, n_11688, n_11689, n_11690,
       n_11691;
  wire n_11692, n_11693, n_11694, n_11695, n_11696, n_11697, n_11698,
       n_11699;
  wire n_11700, n_11701, n_11702, n_11703, n_11704, n_11705, n_11706,
       n_11707;
  wire n_11708, n_11709, n_11710, n_11711, n_11712, n_11713, n_11714,
       n_11715;
  wire n_11716, n_11717, n_11718, n_11719, n_11720, n_11721, n_11722,
       n_11723;
  wire n_11725, n_11726, n_11727, n_11728, n_11729, n_11730, n_11731,
       n_11732;
  wire n_11733, n_11734, n_11735, n_11736, n_11737, n_11738, n_11739,
       n_11740;
  wire n_11741, n_11742, n_11743, n_11744, n_11745, n_11746, n_11747,
       n_11749;
  wire n_11750, n_11751, n_11753, n_11755, n_11756, n_11757, n_11758,
       n_11759;
  wire n_11760, n_11761, n_11762, n_11763, n_11764, n_11767, n_11768,
       n_11770;
  wire n_11771, n_11772, n_11773, n_11774, n_11775, n_11776, n_11777,
       n_11778;
  wire n_11779, n_11780, n_11781, n_11782, n_11783, n_11784, n_11785,
       n_11787;
  wire n_11789, n_11790, n_11792, n_11793, n_11794, n_11795, n_11796,
       n_11797;
  wire n_11798, n_11799, n_11800, n_11801, n_11803, n_11804, n_11806,
       n_11808;
  wire n_11809, n_11810, n_11811, n_11812, n_11813, n_11814, n_11815,
       n_11816;
  wire n_11817, n_11819, n_11821, n_11823, n_11824, n_11825, n_11826,
       n_11828;
  wire n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835,
       n_11836;
  wire n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843,
       n_11844;
  wire n_11845, n_11846, n_11847, n_11848, n_11849, n_11850, n_11851,
       n_11852;
  wire n_11853, n_11854, n_11855, n_11856, n_11857, n_11858, n_11859,
       n_11860;
  wire n_11861, n_11862, n_11863, n_11864, n_11865, n_11866, n_11867,
       n_11868;
  wire n_11869, n_11870, n_11871, n_11872, n_11873, n_11874, n_11875,
       n_11876;
  wire n_11877, n_11878, n_11879, n_11880, n_11881, n_11882, n_11883,
       n_11884;
  wire n_11885, n_11886, n_11887, n_11888, n_11889, n_11890, n_11891,
       n_11892;
  wire n_11893, n_11894, n_11895, n_11896, n_11897, n_11898, n_11899,
       n_11900;
  wire n_11901, n_11902, n_11903, n_11904, n_11905, n_11906, n_11907,
       n_11908;
  wire n_11909, n_11910, n_11912, n_11913, n_11914, n_11915, n_11916,
       n_11917;
  wire n_11918, n_11919, n_11920, n_11921, n_11922, n_11923, n_11924,
       n_11925;
  wire n_11926, n_11927, n_11928, n_11929, n_11930, n_11931, n_11932,
       n_11933;
  wire n_11934, n_11935, n_11936, n_11937, n_11938, n_11939, n_11940,
       n_11941;
  wire n_11942, n_11943, n_11944, n_11945, n_11946, n_11947, n_11948,
       n_11949;
  wire n_11950, n_11951, n_11952, n_11953, n_11954, n_11955, n_11956,
       n_11957;
  wire n_11958, n_11959, n_11960, n_11961, n_11962, n_11963, n_11964,
       n_11965;
  wire n_11967, n_11968, n_11969, n_11970, n_11971, n_11972, n_11973,
       n_11974;
  wire n_11975, n_11976, n_11977, n_11978, n_11979, n_11980, n_11981,
       n_11982;
  wire n_11984, n_11985, n_11986, n_11987, n_11988, n_11989, n_11990,
       n_11991;
  wire n_11992, n_11993, n_11994, n_11995, n_11996, n_11997, n_11998,
       n_11999;
  wire n_12000, n_12001, n_12002, n_12003, n_12004, n_12005, n_12006,
       n_12007;
  wire n_12008, n_12009, n_12010, n_12011, n_12012, n_12013, n_12014,
       n_12015;
  wire n_12016, n_12017, n_12018, n_12019, n_12020, n_12021, n_12022,
       n_12023;
  wire n_12024, n_12025, n_12026, n_12027, n_12028, n_12029, n_12030,
       n_12031;
  wire n_12032, n_12033, n_12034, n_12035, n_12036, n_12037, n_12038,
       n_12039;
  wire n_12040, n_12041, n_12042, n_12043, n_12044, n_12045, n_12046,
       n_12047;
  wire n_12048, n_12049, n_12050, n_12051, n_12052, n_12053, n_12054,
       n_12055;
  wire n_12056, n_12057, n_12058, n_12059, n_12060, n_12061, n_12062,
       n_12063;
  wire n_12064, n_12065, n_12066, n_12067, n_12068, n_12069, n_12070,
       n_12071;
  wire n_12072, n_12073, n_12074, n_12075, n_12076, n_12077, n_12078,
       n_12079;
  wire n_12080, n_12081, n_12082, n_12083, n_12084, n_12085, n_12086,
       n_12087;
  wire n_12088, n_12089, n_12090, n_12091, n_12092, n_12093, n_12094,
       n_12095;
  wire n_12096, n_12097, n_12098, n_12099, n_12100, n_12101, n_12102,
       n_12103;
  wire n_12104, n_12105, n_12106, n_12107, n_12108, n_12109, n_12110,
       n_12111;
  wire n_12112, n_12113, n_12114, n_12115, n_12116, n_12117, n_12118,
       n_12119;
  wire n_12120, n_12121, n_12122, n_12123, n_12124, n_12125, n_12126,
       n_12127;
  wire n_12128, n_12129, n_12130, n_12131, n_12132, n_12133, n_12134,
       n_12135;
  wire n_12136, n_12137, n_12138, n_12139, n_12140, n_12141, n_12142,
       n_12143;
  wire n_12144, n_12145, n_12146, n_12147, n_12148, n_12149, n_12150,
       n_12151;
  wire n_12152, n_12153, n_12154, n_12155, n_12156, n_12157, n_12158,
       n_12159;
  wire n_12160, n_12161, n_12162, n_12163, n_12164, n_12165, n_12166,
       n_12167;
  wire n_12168, n_12169, n_12170, n_12171, n_12172, n_12173, n_12174,
       n_12175;
  wire n_12176, n_12177, n_12178, n_12179, n_12180, n_12181, n_12182,
       n_12183;
  wire n_12184, n_12185, n_12186, n_12187, n_12188, n_12189, n_12190,
       n_12191;
  wire n_12192, n_12193, n_12194, n_12195, n_12196, n_12197, n_12198,
       n_12199;
  wire n_12200, n_12201, n_12202, n_12203, n_12204, n_12205, n_12206,
       n_12207;
  wire n_12208, n_12209, n_12210, n_12211, n_12212, n_12213, n_12214,
       n_12215;
  wire n_12216, n_12217, n_12218, n_12219, n_12220, n_12221, n_12222,
       n_12223;
  wire n_12224, n_12225, n_12226, n_12227, n_12228, n_12229, n_12230,
       n_12231;
  wire n_12232, n_12233, n_12234, n_12235, n_12236, n_12237, n_12238,
       n_12239;
  wire n_12240, n_12241, n_12242, n_12243, n_12244, n_12245, n_12246,
       n_12247;
  wire n_12248, n_12249, n_12250, n_12251, n_12252, n_12253, n_12254,
       n_12255;
  wire n_12256, n_12257, n_12258, n_12259, n_12260, n_12261, n_12262,
       n_12263;
  wire n_12264, n_12265, n_12266, n_12267, n_12268, n_12269, n_12270,
       n_12271;
  wire n_12272, n_12273, n_12274, n_12275, n_12276, n_12277, n_12278,
       n_12279;
  wire n_12280, n_12281, n_12282, n_12283, n_12284, n_12285, n_12286,
       n_12287;
  wire n_12288, n_12289, n_12290, n_12291, n_12292, n_12293, n_12294,
       n_12295;
  wire n_12296, n_12297, n_12298, n_12299, n_12300, n_12301, n_12302,
       n_12303;
  wire n_12304, n_12305, n_12306, n_12307, n_12308, n_12309, n_12310,
       n_12311;
  wire n_12312, n_12313, n_12314, n_12315, n_12316, n_12317, n_12318,
       n_12320;
  wire n_12321, n_12322, n_12323, n_12324, n_12325, n_12326, n_12327,
       n_12328;
  wire n_12329, n_12330, n_12331, n_12332, n_12333, n_12334, n_12335,
       n_12336;
  wire n_12337, n_12338, n_12339, n_12340, n_12341, n_12342, n_12343,
       n_12344;
  wire n_12345, n_12346, n_12347, n_12348, n_12349, n_12350, n_12351,
       n_12352;
  wire n_12354, n_12355, n_12356, n_12357, n_12358, n_12359, n_12360,
       n_12361;
  wire n_12362, n_12363, n_12364, n_12365, n_12366, n_12367, n_12368,
       n_12369;
  wire n_12370, n_12371, n_12372, n_12373, n_12375, n_12376, n_12377,
       n_12378;
  wire n_12379, n_12380, n_12381, n_12382, n_12383, n_12384, n_12385,
       n_12387;
  wire n_12388, n_12389, n_12390, n_12391, n_12392, n_12393, n_12394,
       n_12395;
  wire n_12396, n_12397, n_12399, n_12400, n_12401, n_12402, n_12403,
       n_12404;
  wire n_12405, n_12406, n_12407, n_12409, n_12410, n_12411, n_12412,
       n_12413;
  wire n_12415, n_12416, n_12417, n_12418, n_12419, n_12420, n_12421,
       n_12422;
  wire n_12423, n_12424, n_12425, n_12426, n_12427, n_12428, n_12429,
       n_12430;
  wire n_12431, n_12432, n_12433, n_12434, n_12435, n_12436, n_12437,
       n_12438;
  wire n_12439, n_12440, n_12441, n_12442, n_12443, n_12444, n_12445,
       n_12446;
  wire n_12447, n_12448, n_12449, n_12450, n_12451, n_12452, n_12453,
       n_12454;
  wire n_12455, n_12456, n_12457, n_12458, n_12459, n_12460, n_12461,
       n_12462;
  wire n_12463, n_12464, n_12465, n_12466, n_12467, n_12468, n_12469,
       n_12470;
  wire n_12471, n_12472, n_12473, n_12474, n_12475, n_12476, n_12477,
       n_12478;
  wire n_12479, n_12480, n_12481, n_12482, n_12483, n_12484, n_12485,
       n_12486;
  wire n_12487, n_12488, n_12489, n_12490, n_12491, n_12492, n_12493,
       n_12494;
  wire n_12495, n_12496, n_12497, n_12498, n_12499, n_12500, n_12501,
       n_12502;
  wire n_12503, n_12504, n_12505, n_12506, n_12507, n_12508, n_12509,
       n_12510;
  wire n_12511, n_12512, n_12513, n_12514, n_12515, n_12516, n_12517,
       n_12518;
  wire n_12519, n_12520, n_12521, n_12522, n_12523, n_12524, n_12525,
       n_12526;
  wire n_12527, n_12528, n_12529, n_12530, n_12531, n_12532, n_12533,
       n_12534;
  wire n_12535, n_12536, n_12537, n_12538, n_12539, n_12540, n_12541,
       n_12542;
  wire n_12543, n_12544, n_12545, n_12546, n_12547, n_12548, n_12549,
       n_12550;
  wire n_12551, n_12552, n_12553, n_12554, n_12555, n_12556, n_12557,
       n_12558;
  wire n_12559, n_12560, n_12561, n_12562, n_12563, n_12564, n_12565,
       n_12566;
  wire n_12567, n_12568, n_12569, n_12570, n_12571, n_12572, n_12573,
       n_12574;
  wire n_12575, n_12576, n_12577, n_12578, n_12579, n_12580, n_12581,
       n_12582;
  wire n_12583, n_12584, n_12585, n_12586, n_12587, n_12588, n_12589,
       n_12590;
  wire n_12591, n_12592, n_12593, n_12594, n_12595, n_12596, n_12597,
       n_12598;
  wire n_12599, n_12600, n_12601, n_12602, n_12603, n_12604, n_12605,
       n_12606;
  wire n_12607, n_12608, n_12609, n_12610, n_12612, n_12613, n_12614,
       n_12615;
  wire n_12616, n_12617, n_12618, n_12619, n_12620, n_12621, n_12622,
       n_12623;
  wire n_12624, n_12625, n_12626, n_12627, n_12628, n_12629, n_12630,
       n_12631;
  wire n_12632, n_12633, n_12634, n_12635, n_12636, n_12637, n_12638,
       n_12639;
  wire n_12640, n_12641, n_12642, n_12643, n_12644, n_12645, n_12646,
       n_12647;
  wire n_12648, n_12649, n_12650, n_12651, n_12652, n_12653, n_12654,
       n_12655;
  wire n_12656, n_12657, n_12659, n_12660, n_12661, n_12662, n_12663,
       n_12664;
  wire n_12665, n_12666, n_12667, n_12668, n_12669, n_12670, n_12671,
       n_12672;
  wire n_12673, n_12674, n_12675, n_12676, n_12677, n_12678, n_12679,
       n_12680;
  wire n_12681, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687,
       n_12688;
  wire n_12689, n_12690, n_12691, n_12692, n_12693, n_12694, n_12695,
       n_12696;
  wire n_12697, n_12698, n_12699, n_12700, n_12701, n_12702, n_12703,
       n_12704;
  wire n_12705, n_12706, n_12707, n_12708, n_12709, n_12710, n_12711,
       n_12712;
  wire n_12713, n_12714, n_12715, n_12716, n_12717, n_12718, n_12719,
       n_12720;
  wire n_12721, n_12722, n_12723, n_12724, n_12725, n_12726, n_12727,
       n_12728;
  wire n_12729, n_12730, n_12731, n_12732, n_12733, n_12734, n_12735,
       n_12736;
  wire n_12737, n_12738, n_12739, n_12740, n_12741, n_12742, n_12743,
       n_12744;
  wire n_12745, n_12746, n_12747, n_12748, n_12749, n_12750, n_12751,
       n_12752;
  wire n_12753, n_12754, n_12755, n_12756, n_12757, n_12758, n_12759,
       n_12760;
  wire n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767,
       n_12768;
  wire n_12769, n_12770, n_12771, n_12772, n_12773, n_12774, n_12775,
       n_12776;
  wire n_12777, n_12778, n_12779, n_12780, n_12781, n_12782, n_12783,
       n_12784;
  wire n_12785, n_12786, n_12787, n_12788, n_12789, n_12790, n_12791,
       n_12792;
  wire n_12793, n_12794, n_12795, n_12796, n_12797, n_12798, n_12799,
       n_12800;
  wire n_12801, n_12802, n_12803, n_12804, n_12805, n_12806, n_12807,
       n_12808;
  wire n_12809, n_12810, n_12811, n_12812, n_12813, n_12814, n_12815,
       n_12816;
  wire n_12817, n_12818, n_12819, n_12820, n_12821, n_12822, n_12823,
       n_12824;
  wire n_12825, n_12826, n_12827, n_12828, n_12829, n_12830, n_12831,
       n_12832;
  wire n_12833, n_12834, n_12835, n_12836, n_12837, n_12838, n_12839,
       n_12840;
  wire n_12841, n_12842, n_12843, n_12844, n_12845, n_12846, n_12847,
       n_12848;
  wire n_12849, n_12850, n_12851, n_12852, n_12853, n_12854, n_12855,
       n_12856;
  wire n_12857, n_12858, n_12859, n_12860, n_12861, n_12862, n_12863,
       n_12864;
  wire n_12865, n_12866, n_12867, n_12868, n_12869, n_12870, n_12871,
       n_12872;
  wire n_12873, n_12874, n_12875, n_12876, n_12877, n_12878, n_12879,
       n_12880;
  wire n_12881, n_12882, n_12883, n_12884, n_12885, n_12886, n_12887,
       n_12888;
  wire n_12889, n_12890, n_12891, n_12892, n_12893, n_12894, n_12895,
       n_12896;
  wire n_12897, n_12898, n_12899, n_12900, n_12901, n_12902, n_12903,
       n_12904;
  wire n_12905, n_12906, n_12907, n_12908, n_12909, n_12910, n_12911,
       n_12912;
  wire n_12913, n_12914, n_12915, n_12916, n_12917, n_12918, n_12919,
       n_12920;
  wire n_12921, n_12922, n_12923, n_12924, n_12925, n_12926, n_12927,
       n_12928;
  wire n_12929, n_12930, n_12931, n_12932, n_12933, n_12934, n_12935,
       n_12936;
  wire n_12937, n_12938, n_12939, n_12940, n_12941, n_12942, n_12943,
       n_12944;
  wire n_12945, n_12946, n_12947, n_12948, n_12949, n_12950, n_12951,
       n_12952;
  wire n_12953, n_12954, n_12955, n_12956, n_12957, n_12958, n_12959,
       n_12960;
  wire n_12961, n_12962, n_12963, n_12964, n_12965, n_12966, n_12967,
       n_12968;
  wire n_12969, n_12970, n_12971, n_12972, n_12973, n_12974, n_12975,
       n_12976;
  wire n_12977, n_12978, n_12979, n_12980, n_12981, n_12982, n_12983,
       n_12984;
  wire n_12985, n_12986, n_12987, n_12988, n_12989, n_12990, n_12991,
       n_12992;
  wire n_12993, n_12994, n_12995, n_12996, n_12997, n_12998, n_12999,
       n_13000;
  wire n_13001, n_13002, n_13003, n_13004, n_13005, n_13006, n_13007,
       n_13008;
  wire n_13009, n_13010, n_13011, n_13012, n_13013, n_13014, n_13015,
       n_13016;
  wire n_13017, n_13018, n_13019, n_13020, n_13021, n_13022, n_13023,
       n_13024;
  wire n_13025, n_13026, n_13027, n_13028, n_13029, n_13030, n_13031,
       n_13032;
  wire n_13033, n_13034, n_13035, n_13036, n_13037, n_13039, n_13040,
       n_13041;
  wire n_13042, n_13043, n_13044, n_13045, n_13046, n_13047, n_13048,
       n_13049;
  wire n_13050, n_13051, n_13052, n_13053, n_13054, n_13055, n_13056,
       n_13057;
  wire n_13058, n_13059, n_13060, n_13061, n_13062, n_13063, n_13064,
       n_13065;
  wire n_13066, n_13067, n_13068, n_13069, n_13070, n_13071, n_13072,
       n_13073;
  wire n_13074, n_13075, n_13076, n_13077, n_13078, n_13079, n_13080,
       n_13081;
  wire n_13082, n_13083, n_13084, n_13085, n_13086, n_13087, n_13088,
       n_13089;
  wire n_13090, n_13091, n_13092, n_13093, n_13094, n_13095, n_13096,
       n_13097;
  wire n_13098, n_13099, n_13100, n_13101, n_13102, n_13103, n_13104,
       n_13105;
  wire n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13112,
       n_13113;
  wire n_13114, n_13115, n_13116, n_13117, n_13118, n_13119, n_13120,
       n_13121;
  wire n_13122, n_13123, n_13124, n_13125, n_13126, n_13127, n_13128,
       n_13129;
  wire n_13130, n_13131, n_13132, n_13133, n_13134, n_13135, n_13137,
       n_13138;
  wire n_13139, n_13140, n_13141, n_13142, n_13143, n_13144, n_13145,
       n_13146;
  wire n_13147, n_13148, n_13149, n_13150, n_13151, n_13152, n_13153,
       n_13154;
  wire n_13155, n_13156, n_13157, n_13158, n_13159, n_13160, n_13161,
       n_13162;
  wire n_13163, n_13164, n_13165, n_13166, n_13167, n_13168, n_13169,
       n_13170;
  wire n_13171, n_13172, n_13173, n_13174, n_13175, n_13176, n_13177,
       n_13178;
  wire n_13179, n_13180, n_13181, n_13182, n_13183, n_13184, n_13185,
       n_13186;
  wire n_13187, n_13188, n_13189, n_13190, n_13191, n_13192, n_13193,
       n_13194;
  wire n_13195, n_13196, n_13197, n_13198, n_13199, n_13200, n_13201,
       n_13202;
  wire n_13203, n_13204, n_13205, n_13206, n_13207, n_13208, n_13209,
       n_13210;
  wire n_13211, n_13212, n_13213, n_13214, n_13215, n_13216, n_13217,
       n_13218;
  wire n_13219, n_13220, n_13221, n_13222, n_13223, n_13224, n_13225,
       n_13226;
  wire n_13227, n_13228, n_13229, n_13230, n_13231, n_13232, n_13233,
       n_13234;
  wire n_13235, n_13236, n_13237, n_13238, n_13239, n_13240, n_13241,
       n_13242;
  wire n_13243, n_13244, n_13245, n_13246, n_13247, n_13248, n_13249,
       n_13250;
  wire n_13251, n_13252, n_13253, n_13254, n_13255, n_13256, n_13257,
       n_13258;
  wire n_13259, n_13260, n_13261, n_13262, n_13263, n_13264, n_13265,
       n_13266;
  wire n_13267, n_13268, n_13269, n_13270, n_13271, n_13272, n_13273,
       n_13274;
  wire n_13275, n_13276, n_13277, n_13278, n_13279, n_13280, n_13281,
       n_13282;
  wire n_13283, n_13284, n_13285, n_13286, n_13287, n_13288, n_13289,
       n_13290;
  wire n_13291, n_13292, n_13293, n_13294, n_13295, n_13296, n_13297,
       n_13298;
  wire n_13299, n_13300, n_13301, n_13302, n_13303, n_13304, n_13305,
       n_13306;
  wire n_13307, n_13308, n_13309, n_13310, n_13311, n_13312, n_13313,
       n_13314;
  wire n_13315, n_13316, n_13317, n_13318, n_13319, n_13320, n_13321,
       n_13322;
  wire n_13323, n_13324, n_13325, n_13326, n_13327, n_13328, n_13329,
       n_13330;
  wire n_13331, n_13332, n_13333, n_13334, n_13335, n_13336, n_13337,
       n_13338;
  wire n_13339, n_13340, n_13341, n_13342, n_13343, n_13344, n_13345,
       n_13346;
  wire n_13347, n_13348, n_13349, n_13350, n_13351, n_13352, n_13353,
       n_13354;
  wire n_13355, n_13356, n_13357, n_13358, n_13359, n_13360, n_13361,
       n_13362;
  wire n_13363, n_13364, n_13365, n_13366, n_13367, n_13368, n_13369,
       n_13370;
  wire n_13371, n_13372, n_13373, n_13374, n_13375, n_13376, n_13377,
       n_13378;
  wire n_13379, n_13380, n_13381, n_13382, n_13383, n_13384, n_13385,
       n_13386;
  wire n_13387, n_13388, n_13389, n_13390, n_13391, n_13392, n_13393,
       n_13394;
  wire n_13395, n_13396, n_13397, n_13398, n_13399, n_13400, n_13401,
       n_13402;
  wire n_13403, n_13404, n_13405, n_13406, n_13407, n_13408, n_13409,
       n_13410;
  wire n_13411, n_13412, n_13413, n_13414, n_13415, n_13416, n_13417,
       n_13418;
  wire n_13419, n_13420, n_13421, n_13422, n_13423, n_13424, n_13425,
       n_13426;
  wire n_13427, n_13428, n_13429, n_13430, n_13431, n_13432, n_13433,
       n_13434;
  wire n_13435, n_13436, n_13437, n_13438, n_13439, n_13440, n_13441,
       n_13442;
  wire n_13443, n_13444, n_13445, n_13446, n_13447, n_13448, n_13449,
       n_13450;
  wire n_13451, n_13452, n_13453, n_13454, n_13455, n_13456, n_13457,
       n_13458;
  wire n_13459, n_13460, n_13461, n_13462, n_13463, n_13464, n_13465,
       n_13466;
  wire n_13467, n_13468, n_13469, n_13470, n_13471, n_13472, n_13473,
       n_13474;
  wire n_13475, n_13476, n_13477, n_13478, n_13479, n_13480, n_13481,
       n_13482;
  wire n_13483, n_13484, n_13485, n_13486, n_13487, n_13488, n_13489,
       n_13490;
  wire n_13491, n_13492, n_13493, n_13494, n_13495, n_13496, n_13497,
       n_13498;
  wire n_13499, n_13500, n_13501, n_13502, n_13503, n_13504, n_13505,
       n_13506;
  wire n_13507, n_13508, n_13509, n_13510, n_13511, n_13512, n_13513,
       n_13514;
  wire n_13515, n_13516, n_13517, n_13518, n_13519, n_13520, n_13521,
       n_13522;
  wire n_13523, n_13524, n_13525, n_13526, n_13527, n_13528, n_13529,
       n_13530;
  wire n_13531, n_13532, n_13533, n_13534, n_13535, n_13536, n_13537,
       n_13538;
  wire n_13539, n_13540, n_13541, n_13542, n_13543, n_13544, n_13545,
       n_13546;
  wire n_13547, n_13548, n_13549, n_13550, n_13551, n_13552, n_13553,
       n_13554;
  wire n_13555, n_13556, n_13557, n_13558, n_13559, n_13560, n_13561,
       n_13562;
  wire n_13563, n_13564, n_13565, n_13566, n_13567, n_13568, n_13569,
       n_13570;
  wire n_13571, n_13572, n_13573, n_13574, n_13575, n_13576, n_13577,
       n_13578;
  wire n_13579, n_13580, n_13581, n_13582, n_13583, n_13584, n_13585,
       n_13586;
  wire n_13587, n_13588, n_13589, n_13590, n_13591, n_13592, n_13593,
       n_13594;
  wire n_13595, n_13596, n_13597, n_13598, n_13599, n_13600, n_13601,
       n_13602;
  wire n_13603, n_13604, n_13605, n_13606, n_13607, n_13608, n_13609,
       n_13610;
  wire n_13611, n_13612, n_13613, n_13614, n_13615, n_13616, n_13617,
       n_13618;
  wire n_13620, n_13621, n_13622, n_13623, n_13624, n_13625, n_13626,
       n_13627;
  wire n_13628, n_13629, n_13630, n_13631, n_13632, n_13633, n_13634,
       n_13635;
  wire n_13636, n_13637, n_13638, n_13639, n_13640, n_13641, n_13642,
       n_13643;
  wire n_13644, n_13645, n_13646, n_13647, n_13648, n_13649, n_13650,
       n_13651;
  wire n_13652, n_13653, n_13654, n_13655, n_13656, n_13657, n_13658,
       n_13659;
  wire n_13660, n_13661, n_13662, n_13663, n_13664, n_13665, n_13666,
       n_13667;
  wire n_13668, n_13670, n_13671, n_13672, n_13673, n_13674, n_13675,
       n_13676;
  wire n_13677, n_13678, n_13679, n_13680, n_13681, n_13682, n_13683,
       n_13684;
  wire n_13685, n_13686, n_13687, n_13688, n_13689, n_13690, n_13691,
       n_13692;
  wire n_13693, n_13694, n_13695, n_13696, n_13697, n_13698, n_13699,
       n_13700;
  wire n_13701, n_13702, n_13703, n_13704, n_13705, n_13706, n_13707,
       n_13708;
  wire n_13709, n_13710, n_13711, n_13714, n_13715, n_13716, n_13717,
       n_13718;
  wire n_13719, n_13720, n_13721, n_13722, n_13723, n_13724, n_13725,
       n_13726;
  wire n_13727, n_13728, n_13729, n_13730, n_13731, n_13732, n_13733,
       n_13734;
  wire n_13735, n_13736, n_13737, n_13738, n_13739, n_13740, n_13741,
       n_13742;
  wire n_13743, n_13744, n_13745, n_13746, n_13747, n_13748, n_13749,
       n_13750;
  wire n_13751, n_13752, n_13753, n_13754, n_13755, n_13756, n_13757,
       n_13758;
  wire n_13759, n_13760, n_13761, n_13762, n_13763, n_13764, n_13765,
       n_13766;
  wire n_13767, n_13768, n_13769, n_13770, n_13771, n_13772, n_13773,
       n_13774;
  wire n_13775, n_13776, n_13777, n_13778, n_13779, n_13780, n_13781,
       n_13782;
  wire n_13783, n_13784, n_13785, n_13786, n_13787, n_13788, n_13789,
       n_13790;
  wire n_13791, n_13792, n_13793, n_13794, n_13795, n_13796, n_13797,
       n_13798;
  wire n_13799, n_13800, n_13801, n_13802, n_13803, n_13804, n_13805,
       n_13806;
  wire n_13807, n_13808, n_13809, n_13810, n_13811, n_13812, n_13813,
       n_13814;
  wire n_13815, n_13816, n_13817, n_13818, n_13819, n_13820, n_13821,
       n_13822;
  wire n_13823, n_13824, n_13825, n_13826, n_13827, n_13828, n_13829,
       n_13830;
  wire n_13831, n_13832, n_13833, n_13834, n_13835, n_13836, n_13837,
       n_13838;
  wire n_13839, n_13840, n_13841, n_13842, n_13843, n_13844, n_13845,
       n_13846;
  wire n_13847, n_13848, n_13849, n_13850, n_13851, n_13852, n_13853,
       n_13854;
  wire n_13855, n_13856, n_13857, n_13858, n_13859, n_13860, n_13861,
       n_13862;
  wire n_13863, n_13864, n_13865, n_13866, n_13867, n_13868, n_13869,
       n_13870;
  wire n_13871, n_13872, n_13873, n_13874, n_13875, n_13876, n_13877,
       n_13878;
  wire n_13879, n_13880, n_13881, n_13882, n_13883, n_13884, n_13885,
       n_13886;
  wire n_13887, n_13888, n_13889, n_13890, n_13891, n_13892, n_13893,
       n_13894;
  wire n_13895, n_13896, n_13897, n_13898, n_13899, n_13900, n_13901,
       n_13902;
  wire n_13903, n_13904, n_13905, n_13906, n_13907, n_13908, n_13909,
       n_13910;
  wire n_13911, n_13912, n_13913, n_13914, n_13915, n_13916, n_13917,
       n_13918;
  wire n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925,
       n_13926;
  wire n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933,
       n_13934;
  wire n_13935, n_13936, n_13937, n_13938, n_13939, n_13940, n_13941,
       n_13942;
  wire n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949,
       n_13950;
  wire n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957,
       n_13958;
  wire n_13959, n_13960, n_13961, n_13962, n_13963, n_13964, n_13965,
       n_13966;
  wire n_13967, n_13968, n_13969, n_13970, n_13971, n_13972, n_13973,
       n_13974;
  wire n_13975, n_13976, n_13977, n_13978, n_13979, n_13980, n_13981,
       n_13982;
  wire n_13983, n_13984, n_13985, n_13986, n_13987, n_13988, n_13989,
       n_13990;
  wire n_13991, n_13992, n_13993, n_13994, n_13995, n_13996, n_13997,
       n_13998;
  wire n_13999, n_14000, n_14001, n_14002, n_14003, n_14004, n_14005,
       n_14006;
  wire n_14007, n_14008, n_14009, n_14010, n_14011, n_14012, n_14013,
       n_14014;
  wire n_14015, n_14016, n_14017, n_14018, n_14019, n_14020, n_14021,
       n_14022;
  wire n_14023, n_14024, n_14025, n_14026, n_14027, n_14028, n_14029,
       n_14030;
  wire n_14031, n_14032, n_14034, n_14035, n_14036, n_14037, n_14038,
       n_14039;
  wire n_14040, n_14041, n_14042, n_14043, n_14044, n_14045, n_14046,
       n_14047;
  wire n_14048, n_14049, n_14050, n_14051, n_14052, n_14053, n_14054,
       n_14055;
  wire n_14056, n_14057, n_14058, n_14059, n_14060, n_14061, n_14062,
       n_14063;
  wire n_14064, n_14065, n_14066, n_14067, n_14068, n_14069, n_14070,
       n_14071;
  wire n_14072, n_14073, n_14074, n_14075, n_14076, n_14077, n_14078,
       n_14079;
  wire n_14080, n_14081, n_14083, n_14084, n_14085, n_14086, n_14087,
       n_14088;
  wire n_14089, n_14090, n_14091, n_14092, n_14093, n_14094, n_14095,
       n_14096;
  wire n_14097, n_14098, n_14099, n_14100, n_14101, n_14102, n_14103,
       n_14104;
  wire n_14105, n_14106, n_14107, n_14108, n_14109, n_14110, n_14111,
       n_14112;
  wire n_14113, n_14114, n_14115, n_14116, n_14117, n_14118, n_14119,
       n_14120;
  wire n_14121, n_14122, n_14123, n_14124, n_14125, n_14126, n_14127,
       n_14128;
  wire n_14129, n_14130, n_14131, n_14132, n_14133, n_14134, n_14135,
       n_14136;
  wire n_14137, n_14138, n_14139, n_14140, n_14142, n_14143, n_14144,
       n_14145;
  wire n_14146, n_14147, n_14148, n_14149, n_14150, n_14151, n_14152,
       n_14153;
  wire n_14154, n_14155, n_14156, n_14157, n_14158, n_14159, n_14160,
       n_14161;
  wire n_14162, n_14163, n_14164, n_14165, n_14166, n_14167, n_14168,
       n_14169;
  wire n_14170, n_14171, n_14172, n_14173, n_14174, n_14175, n_14176,
       n_14177;
  wire n_14178, n_14179, n_14180, n_14181, n_14182, n_14183, n_14184,
       n_14185;
  wire n_14186, n_14187, n_14188, n_14189, n_14190, n_14191, n_14192,
       n_14193;
  wire n_14194, n_14195, n_14196, n_14197, n_14198, n_14199, n_14200,
       n_14201;
  wire n_14202, n_14203, n_14204, n_14205, n_14206, n_14207, n_14208,
       n_14209;
  wire n_14210, n_14211, n_14212, n_14213, n_14214, n_14215, n_14216,
       n_14217;
  wire n_14218, n_14219, n_14220, n_14221, n_14222, n_14223, n_14224,
       n_14225;
  wire n_14226, n_14227, n_14228, n_14229, n_14230, n_14231, n_14232,
       n_14233;
  wire n_14234, n_14235, n_14236, n_14237, n_14238, n_14239, n_14240,
       n_14241;
  wire n_14242, n_14243, n_14244, n_14245, n_14246, n_14247, n_14248,
       n_14249;
  wire n_14250, n_14251, n_14252, n_14253, n_14254, n_14255, n_14256,
       n_14257;
  wire n_14258, n_14259, n_14260, n_14261, n_14262, n_14263, n_14264,
       n_14265;
  wire n_14266, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272,
       n_14273;
  wire n_14274, n_14275, n_14276, n_14277, n_14278, n_14279, n_14280,
       n_14281;
  wire n_14282, n_14283, n_14284, n_14285, n_14286, n_14287, n_14288,
       n_14289;
  wire n_14290, n_14291, n_14292, n_14293, n_14294, n_14295, n_14296,
       n_14297;
  wire n_14298, n_14299, n_14300, n_14301, n_14302, n_14303, n_14304,
       n_14305;
  wire n_14306, n_14307, n_14308, n_14309, n_14310, n_14311, n_14312,
       n_14313;
  wire n_14314, n_14315, n_14316, n_14317, n_14318, n_14319, n_14320,
       n_14321;
  wire n_14322, n_14323, n_14324, n_14325, n_14326, n_14327, n_14328,
       n_14329;
  wire n_14330, n_14331, n_14332, n_14333, n_14334, n_14335, n_14336,
       n_14337;
  wire n_14338, n_14339, n_14340, n_14341, n_14342, n_14343, n_14344,
       n_14345;
  wire n_14346, n_14347, n_14348, n_14349, n_14350, n_14351, n_14352,
       n_14353;
  wire n_14354, n_14355, n_14356, n_14357, n_14358, n_14359, n_14360,
       n_14361;
  wire n_14362, n_14363, n_14364, n_14365, n_14366, n_14367, n_14368,
       n_14369;
  wire n_14370, n_14371, n_14372, n_14373, n_14374, n_14375, n_14376,
       n_14377;
  wire n_14378, n_14379, n_14380, n_14381, n_14382, n_14383, n_14384,
       n_14385;
  wire n_14386, n_14387, n_14388, n_14389, n_14390, n_14391, n_14392,
       n_14393;
  wire n_14394, n_14395, n_14396, n_14397, n_14398, n_14399, n_14400,
       n_14401;
  wire n_14402, n_14403, n_14404, n_14405, n_14406, n_14407, n_14408,
       n_14409;
  wire n_14410, n_14411, n_14412, n_14413, n_14414, n_14415, n_14416,
       n_14417;
  wire n_14418, n_14419, n_14420, n_14421, n_14422, n_14424, n_14425,
       n_14426;
  wire n_14427, n_14428, n_14429, n_14430, n_14431, n_14432, n_14433,
       n_14434;
  wire n_14435, n_14436, n_14437, n_14438, n_14439, n_14440, n_14441,
       n_14442;
  wire n_14443, n_14444, n_14445, n_14446, n_14447, n_14448, n_14449,
       n_14450;
  wire n_14451, n_14452, n_14453, n_14454, n_14455, n_14456, n_14457,
       n_14458;
  wire n_14459, n_14460, n_14461, n_14462, n_14463, n_14464, n_14465,
       n_14466;
  wire n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, n_14473,
       n_14474;
  wire n_14475, n_14476, n_14478, n_14479, n_14480, n_14481, n_14482,
       n_14483;
  wire n_14484, n_14485, n_14486, n_14487, n_14488, n_14489, n_14490,
       n_14491;
  wire n_14492, n_14493, n_14494, n_14495, n_14496, n_14497, n_14498,
       n_14499;
  wire n_14500, n_14501, n_14502, n_14503, n_14504, n_14505, n_14506,
       n_14507;
  wire n_14508, n_14509, n_14510, n_14511, n_14512, n_14513, n_14514,
       n_14515;
  wire n_14516, n_14517, n_14518, n_14519, n_14520, n_14521, n_14522,
       n_14523;
  wire n_14524, n_14525, n_14526, n_14527, n_14528, n_14529, n_14530,
       n_14531;
  wire n_14532, n_14533, n_14534, n_14535, n_14536, n_14537, n_14538,
       n_14539;
  wire n_14540, n_14541, n_14542, n_14543, n_14544, n_14545, n_14546,
       n_14547;
  wire n_14548, n_14549, n_14550, n_14551, n_14552, n_14553, n_14554,
       n_14555;
  wire n_14556, n_14557, n_14558, n_14559, n_14560, n_14561, n_14562,
       n_14563;
  wire n_14564, n_14565, n_14566, n_14567, n_14568, n_14569, n_14570,
       n_14571;
  wire n_14572, n_14573, n_14574, n_14575, n_14576, n_14577, n_14578,
       n_14579;
  wire n_14580, n_14581, n_14582, n_14583, n_14584, n_14585, n_14586,
       n_14587;
  wire n_14588, n_14589, n_14590, n_14591, n_14592, n_14593, n_14594,
       n_14595;
  wire n_14596, n_14597, n_14598, n_14599, n_14600, n_14601, n_14602,
       n_14603;
  wire n_14604, n_14605, n_14606, n_14607, n_14608, n_14609, n_14610,
       n_14611;
  wire n_14612, n_14613, n_14614, n_14615, n_14616, n_14617, n_14618,
       n_14619;
  wire n_14620, n_14621, n_14622, n_14623, n_14624, n_14625, n_14626,
       n_14627;
  wire n_14628, n_14629, n_14630, n_14631, n_14632, n_14633, n_14634,
       n_14635;
  wire n_14636, n_14637, n_14638, n_14639, n_14640, n_14641, n_14642,
       n_14643;
  wire n_14644, n_14645, n_14646, n_14647, n_14648, n_14649, n_14650,
       n_14651;
  wire n_14652, n_14653, n_14654, n_14655, n_14656, n_14657, n_14658,
       n_14659;
  wire n_14660, n_14661, n_14662, n_14663, n_14664, n_14665, n_14666,
       n_14667;
  wire n_14668, n_14669, n_14670, n_14671, n_14672, n_14673, n_14674,
       n_14675;
  wire n_14676, n_14677, n_14678, n_14679, n_14680, n_14681, n_14682,
       n_14683;
  wire n_14684, n_14685, n_14686, n_14687, n_14688, n_14689, n_14690,
       n_14691;
  wire n_14692, n_14693, n_14694, n_14695, n_14696, n_14697, n_14698,
       n_14699;
  wire n_14700, n_14701, n_14702, n_14703, n_14704, n_14705, n_14706,
       n_14707;
  wire n_14708, n_14709, n_14710, n_14711, n_14712, n_14713, n_14714,
       n_14715;
  wire n_14716, n_14717, n_14718, n_14719, n_14720, n_14721, n_14722,
       n_14723;
  wire n_14724, n_14725, n_14726, n_14727, n_14728, n_14729, n_14730,
       n_14731;
  wire n_14732, n_14733, n_14734, n_14735, n_14736, n_14737, n_14738,
       n_14739;
  wire n_14740, n_14741, n_14742, n_14743, n_14744, n_14745, n_14746,
       n_14747;
  wire n_14748, n_14749, n_14750, n_14751, n_14752, n_14753, n_14754,
       n_14755;
  wire n_14756, n_14757, n_14758, n_14759, n_14760, n_14761, n_14762,
       n_14763;
  wire n_14764, n_14765, n_14766, n_14767, n_14768, n_14769, n_14770,
       n_14771;
  wire n_14772, n_14773, n_14774, n_14775, n_14776, n_14777, n_14778,
       n_14779;
  wire n_14780, n_14781, n_14782, n_14783, n_14784, n_14785, n_14786,
       n_14787;
  wire n_14788, n_14789, n_14790, n_14791, n_14792, n_14793, n_14794,
       n_14795;
  wire n_14796, n_14797, n_14798, n_14799, n_14800, n_14801, n_14802,
       n_14803;
  wire n_14804, n_14805, n_14806, n_14807, n_14808, n_14809, n_14810,
       n_14811;
  wire n_14812, n_14813, n_14814, n_14815, n_14816, n_14817, n_14818,
       n_14819;
  wire n_14820, n_14821, n_14822, n_14823, n_14824, n_14825, n_14826,
       n_14827;
  wire n_14828, n_14829, n_14830, n_14831, n_14832, n_14833, n_14834,
       n_14835;
  wire n_14836, n_14837, n_14838, n_14839, n_14840, n_14841, n_14842,
       n_14843;
  wire n_14844, n_14845, n_14846, n_14847, n_14848, n_14849, n_14850,
       n_14851;
  wire n_14852, n_14853, n_14854, n_14855, n_14856, n_14857, n_14858,
       n_14859;
  wire n_14860, n_14861, n_14862, n_14863, n_14864, n_14865, n_14866,
       n_14867;
  wire n_14868, n_14869, n_14870, n_14871, n_14872, n_14873, n_14875,
       n_14877;
  wire n_14878, n_14879, n_14880, n_14881, n_14882, n_14883, n_14884,
       n_14885;
  wire n_14886, n_14887, n_14888, n_14889, n_14890, n_14891, n_14892,
       n_14893;
  wire n_14894, n_14895, n_14896, n_14897, n_14898, n_14899, n_14900,
       n_14901;
  wire n_14902, n_14903, n_14904, n_14905, n_14906, n_14907, n_14908,
       n_14909;
  wire n_14910, n_14911, n_14912, n_14913, n_14914, n_14915, n_14916,
       n_14917;
  wire n_14918, n_14919, n_14920, n_14921, n_14922, n_14923, n_14924,
       n_14925;
  wire n_14926, n_14927, n_14928, n_14929, n_14930, n_14931, n_14932,
       n_14933;
  wire n_14934, n_14935, n_14936, n_14937, n_14938, n_14939, n_14940,
       n_14941;
  wire n_14942, n_14943, n_14944, n_14945, n_14946, n_14947, n_14948,
       n_14949;
  wire n_14950, n_14951, n_14952, n_14953, n_14954, n_14955, n_14956,
       n_14957;
  wire n_14958, n_14959, n_14960, n_14961, n_14962, n_14963, n_14964,
       n_14965;
  wire n_14966, n_14967, n_14968, n_14969, n_14970, n_14971, n_14972,
       n_14973;
  wire n_14974, n_14975, n_14976, n_14977, n_14978, n_14979, n_14980,
       n_14981;
  wire n_14982, n_14983, n_14984, n_14985, n_14986, n_14987, n_14988,
       n_14989;
  wire n_14990, n_14991, n_14992, n_14993, n_14994, n_14995, n_14996,
       n_14997;
  wire n_14998, n_14999, n_15000, n_15001, n_15002, n_15003, n_15004,
       n_15005;
  wire n_15006, n_15007, n_15008, n_15009, n_15010, n_15011, n_15012,
       n_15013;
  wire n_15014, n_15015, n_15016, n_15017, n_15018, n_15019, n_15020,
       n_15021;
  wire n_15022, n_15023, n_15024, n_15025, n_15026, n_15027, n_15028,
       n_15029;
  wire n_15030, n_15031, n_15032, n_15034, n_15036, n_15037, n_15038,
       n_15039;
  wire n_15040, n_15041, n_15042, n_15043, n_15044, n_15045, n_15046,
       n_15047;
  wire n_15048, n_15049, n_15050, n_15051, n_15052, n_15053, n_15054,
       n_15055;
  wire n_15056, n_15057, n_15058, n_15059, n_15062, n_15063, n_15064,
       n_15065;
  wire n_15066, n_15067, n_15068, n_15069, n_15070, n_15071, n_15072,
       n_15073;
  wire n_15074, n_15075, n_15076, n_15077, n_15078, n_15080, n_15081,
       n_15082;
  wire n_15083, n_15084, n_15085, n_15086, n_15087, n_15088, n_15089,
       n_15090;
  wire n_15091, n_15092, n_15093, n_15095, n_15096, n_15097, n_15098,
       n_15099;
  wire n_15100, n_15101, n_15102, n_15103, n_15104, n_15105, n_15106,
       n_15107;
  wire n_15108, n_15109, n_15110, n_15111, n_15112, n_15113, n_15114,
       n_15115;
  wire n_15116, n_15117, n_15118, n_15119, n_15120, n_15121, n_15122,
       n_15123;
  wire n_15125, n_15127, n_15128, n_15129, n_15130, n_15131, n_15132,
       n_15133;
  wire n_15134, n_15135, n_15136, n_15137, n_15138, n_15139, n_15140,
       n_15141;
  wire n_15142, n_15143, n_15144, n_15145, n_15146, n_15147, n_15148,
       n_15149;
  wire n_15150, n_15151, n_15152, n_15153, n_15154, n_15155, n_15156,
       n_15157;
  wire n_15158, n_15159, n_15160, n_15161, n_15162, n_15163, n_15164,
       n_15165;
  wire n_15166, n_15167, n_15168, n_15169, n_15170, n_15171, n_15172,
       n_15173;
  wire n_15174, n_15175, n_15176, n_15177, n_15178, n_15179, n_15180,
       n_15181;
  wire n_15182, n_15183, n_15184, n_15185, n_15186, n_15187, n_15188,
       n_15189;
  wire n_15191, n_15192, n_15193, n_15194, n_15195, n_15196, n_15197,
       n_15198;
  wire n_15199, n_15200, n_15201, n_15202, n_15203, n_15204, n_15205,
       n_15206;
  wire n_15207, n_15208, n_15209, n_15210, n_15211, n_15212, n_15213,
       n_15214;
  wire n_15215, n_15216, n_15217, n_15218, n_15219, n_15220, n_15221,
       n_15222;
  wire n_15223, n_15224, n_15225, n_15226, n_15227, n_15228, n_15229,
       n_15230;
  wire n_15231, n_15232, n_15233, n_15235, n_15236, n_15237, n_15238,
       n_15239;
  wire n_15240, n_15241, n_15242, n_15243, n_15244, n_15245, n_15246,
       n_15247;
  wire n_15248, n_15249, n_15250, n_15251, n_15252, n_15253, n_15254,
       n_15255;
  wire n_15256, n_15257, n_15258, n_15259, n_15260, n_15261, n_15262,
       n_15263;
  wire n_15264, n_15266, n_15268, n_15269, n_15270, n_15271, n_15272,
       n_15273;
  wire n_15274, n_15275, n_15276, n_15277, n_15278, n_15279, n_15280,
       n_15281;
  wire n_15282, n_15283, n_15284, n_15285, n_15286, n_15287, n_15288,
       n_15289;
  wire n_15290, n_15291, n_15292, n_15293, n_15294, n_15295, n_15296,
       n_15297;
  wire n_15298, n_15299, n_15300, n_15301, n_15302, n_15303, n_15304,
       n_15305;
  wire n_15306, n_15307, n_15308, n_15309, n_15310, n_15311, n_15312,
       n_15313;
  wire n_15314, n_15315, n_15316, n_15317, n_15318, n_15319, n_15320,
       n_15321;
  wire n_15322, n_15323, n_15324, n_15325, n_15327, n_15329, n_15330,
       n_15331;
  wire n_15332, n_15333, n_15334, n_15335, n_15336, n_15337, n_15338,
       n_15339;
  wire n_15340, n_15341, n_15342, n_15343, n_15344, n_15345, n_15346,
       n_15347;
  wire n_15348, n_15349, n_15350, n_15351, n_15352, n_15353, n_15354,
       n_15355;
  wire n_15356, n_15357, n_15358, n_15359, n_15360, n_15361, n_15362,
       n_15363;
  wire n_15364, n_15365, n_15366, n_15367, n_15368, n_15369, n_15370,
       n_15371;
  wire n_15373, n_15375, n_15376, n_15377, n_15378, n_15379, n_15380,
       n_15381;
  wire n_15382, n_15383, n_15384, n_15385, n_15386, n_15387, n_15388,
       n_15389;
  wire n_15390, n_15391, n_15392, n_15393, n_15394, n_15395, n_15396,
       n_15397;
  wire n_15398, n_15399, n_15400, n_15401, n_15402, n_15403, n_15404,
       n_15405;
  wire n_15406, n_15407, n_15408, n_15409, n_15410, n_15412, n_15414,
       n_15415;
  wire n_15416, n_15417, n_15418, n_15419, n_15420, n_15421, n_15422,
       n_15423;
  wire n_15424, n_15425, n_15426, n_15427, n_15428, n_15429, n_15430,
       n_15431;
  wire n_15432, n_15433, n_15434, n_15435, n_15436, n_15437, n_15438,
       n_15439;
  wire n_15440, n_15442, n_15444, n_15445, n_15446, n_15447, n_15448,
       n_15449;
  wire n_15450, n_15451, n_15452, n_15453, n_15454, n_15455, n_15456,
       n_15457;
  wire n_15458, n_15459, n_15460, n_15461, n_15462, n_15463, n_15464,
       n_15465;
  wire n_15466, n_15467, n_15468, n_15469, n_15470, n_15471, n_15472,
       n_15473;
  wire n_15474, n_15475, n_15476, n_15477, n_15478, n_15479, n_15480,
       n_15481;
  wire n_15482, n_15483, n_15484, n_15485, n_15486, n_15488, n_15489,
       n_15490;
  wire n_15491, n_15492, n_15493, n_15494, n_15495, n_15496, n_15497,
       n_15498;
  wire n_15499, n_15500, n_15501, n_15503, n_15504, n_15505, n_15506,
       n_15507;
  wire n_15508, n_15509, n_15510, n_15511, n_15512, n_15513, n_15514,
       n_15515;
  wire n_15516, n_15517, n_15518, n_15519, n_15520, n_15521, n_15522,
       n_15523;
  wire n_15524, n_15525, n_15526, n_15527, n_15528, n_15529, n_15530,
       n_15531;
  wire n_15533, n_15534, n_15535, n_15536, n_15537, n_15538, n_15539,
       n_15540;
  wire n_15541, n_15542, n_15543, n_15544, n_15545, n_15546, n_15548,
       n_15549;
  wire n_15550, n_15551, n_15552, n_15553, n_15554, n_15555, n_15556,
       n_15557;
  wire n_15558, n_15559, n_15560, n_15561, n_15562, n_15563, n_15564,
       n_15565;
  wire n_15566, n_15567, n_15568, n_15569, n_15570, n_15571, n_15572,
       n_15573;
  wire n_15574, n_15575, n_15576, n_15578, n_15580, n_15581, n_15582,
       n_15583;
  wire n_15584, n_15585, n_15586, n_15587, n_15588, n_15589, n_15590,
       n_15591;
  wire n_15592, n_15593, n_15594, n_15595, n_15596, n_15597, n_15598,
       n_15599;
  wire n_15600, n_15601, n_15602, n_15603, n_15606, n_15607, n_15608,
       n_15609;
  wire n_15610, n_15611, n_15612, n_15613, n_15614, n_15615, n_15616,
       n_15617;
  wire n_15618, n_15619, n_15620, n_15621, n_15622, n_15623, n_15624,
       n_15625;
  wire n_15626, n_15627, n_15628, n_15629, n_15630, n_15631, n_15632,
       n_15633;
  wire n_15634, n_15635, n_15636, n_15637, n_15638, n_15639, n_15640,
       n_15641;
  wire n_15642, n_15643, n_15644, n_15645, n_15646, n_15647, n_15648,
       n_15649;
  wire n_15650, n_15651, n_15652, n_15653, n_15654, n_15655, n_15656,
       n_15657;
  wire n_15658, n_15659, n_15660, n_15661, n_15662, n_15663, n_15664,
       n_15665;
  wire n_15666, n_15667, n_15668, n_15669, n_15670, n_15671, n_15672,
       n_15673;
  wire n_15674, n_15675, n_15676, n_15677, n_15678, n_15679, n_15680,
       n_15681;
  wire n_15682, n_15683, n_15684, n_15685, n_15686, n_15687, n_15688,
       n_15689;
  wire n_15690, n_15691, n_15692, n_15693, n_15694, n_15695, n_15696,
       n_15697;
  wire n_15698, n_15699, n_15700, n_15701, n_15702, n_15703, n_15704,
       n_15705;
  wire n_15706, n_15707, n_15708, n_15709, n_15710, n_15711, n_15712,
       n_15713;
  wire n_15714, n_15715, n_15716, n_15717, n_15718, n_15719, n_15720,
       n_15721;
  wire n_15722, n_15723, n_15724, n_15725, n_15726, n_15727, n_15728,
       n_15730;
  wire n_15732, n_15733, n_15734, n_15735, n_15736, n_15737, n_15738,
       n_15739;
  wire n_15740, n_15741, n_15742, n_15743, n_15744, n_15745, n_15746,
       n_15747;
  wire n_15748, n_15749, n_15750, n_15751, n_15752, n_15753, n_15754,
       n_15755;
  wire n_15758, n_15759, n_15760, n_15761, n_15762, n_15763, n_15764,
       n_15765;
  wire n_15766, n_15767, n_15768, n_15769, n_15770, n_15771, n_15772,
       n_15773;
  wire n_15774, n_15776, n_15778, n_15779, n_15780, n_15781, n_15782,
       n_15783;
  wire n_15784, n_15785, n_15786, n_15787, n_15788, n_15789, n_15790,
       n_15791;
  wire n_15792, n_15793, n_15794, n_15795, n_15796, n_15797, n_15798,
       n_15802;
  wire n_15803, n_15804, n_15805, n_15806, n_15807, n_15808, n_15809,
       n_15810;
  wire n_15811, n_15812, n_15813, n_15814, n_15815, n_15816, n_15817,
       n_15818;
  wire n_15819, n_15820, n_15821, n_15822, n_15823, n_15824, n_15825,
       n_15826;
  wire n_15827, n_15828, n_15832, n_15833, n_15834, n_15835, n_15836,
       n_15837;
  wire n_15838, n_15840, n_15841, n_15842, n_15843, n_15844, n_15845,
       n_15846;
  wire n_15847, n_15848, n_15849, n_15850, n_15851, n_15852, n_15853,
       n_15854;
  wire n_15855, n_15856, n_15857, n_15858, n_15859, n_15860, n_15861,
       n_15862;
  wire n_15863, n_15864, n_15865, n_15866, n_15867, n_15868, n_15870,
       n_15871;
  wire n_15872, n_15873, n_15874, n_15875, n_15876, n_15877, n_15878,
       n_15879;
  wire n_15880, n_15881, n_15882, n_15883, n_15884, n_15885, n_15886,
       n_15887;
  wire n_15888, n_15889, n_15890, n_15891, n_15892, n_15893, n_15894,
       n_15895;
  wire n_15896, n_15897, n_15898, n_15899, n_15900, n_15901, n_15902,
       n_15903;
  wire n_15904, n_15905, n_15906, n_15907, n_15908, n_15909, n_15911,
       n_15913;
  wire n_15914, n_15915, n_15916, n_15917, n_15918, n_15919, n_15920,
       n_15921;
  wire n_15922, n_15923, n_15924, n_15925, n_15926, n_15927, n_15928,
       n_15929;
  wire n_15930, n_15931, n_15932, n_15933, n_15934, n_15935, n_15936,
       n_15937;
  wire n_15938, n_15939, n_15940, n_15941, n_15942, n_15943, n_15944,
       n_15946;
  wire n_15948, n_15949, n_15950, n_15951, n_15952, n_15953, n_15954,
       n_15955;
  wire n_15956, n_15957, n_15958, n_15959, n_15960, n_15961, n_15962,
       n_15963;
  wire n_15964, n_15965, n_15966, n_15967, n_15968, n_15969, n_15970,
       n_15971;
  wire n_15972, n_15973, n_15974, n_15975, n_15976, n_15977, n_15978,
       n_15979;
  wire n_15980, n_15981, n_15982, n_15983, n_15984, n_15985, n_15986,
       n_15987;
  wire n_15988, n_15989, n_15990, n_15991, n_15992, n_15993, n_15994,
       n_15995;
  wire n_15996, n_15997, n_15998, n_15999, n_16000, n_16001, n_16002,
       n_16003;
  wire n_16004, n_16006, n_16008, n_16009, n_16010, n_16011, n_16012,
       n_16013;
  wire n_16014, n_16015, n_16016, n_16017, n_16018, n_16019, n_16020,
       n_16021;
  wire n_16022, n_16023, n_16024, n_16025, n_16026, n_16027, n_16028,
       n_16029;
  wire n_16030, n_16031, n_16032, n_16033, n_16034, n_16035, n_16036,
       n_16037;
  wire n_16038, n_16039, n_16040, n_16041, n_16042, n_16043, n_16044,
       n_16045;
  wire n_16046, n_16047, n_16048, n_16049, n_16050, n_16051, n_16052,
       n_16053;
  wire n_16054, n_16055, n_16056, n_16057, n_16058, n_16059, n_16060,
       n_16061;
  wire n_16062, n_16063, n_16064, n_16067, n_16068, n_16069, n_16070,
       n_16071;
  wire n_16072, n_16073, n_16074, n_16075, n_16076, n_16077, n_16078,
       n_16079;
  wire n_16080, n_16081, n_16082, n_16083, n_16084, n_16085, n_16086,
       n_16087;
  wire n_16088, n_16089, n_16090, n_16091, n_16092, n_16093, n_16094,
       n_16095;
  wire n_16096, n_16097, n_16098, n_16099, n_16100, n_16101, n_16102,
       n_16103;
  wire n_16104, n_16105, n_16106, n_16107, n_16108, n_16109, n_16110,
       n_16111;
  wire n_16112, n_16113, n_16114, n_16115, n_16116, n_16117, n_16118,
       n_16119;
  wire n_16120, n_16121, n_16122, n_16123, n_16124, n_16125, n_16127,
       n_16129;
  wire n_16130, n_16131, n_16132, n_16133, n_16134, n_16135, n_16136,
       n_16137;
  wire n_16138, n_16139, n_16140, n_16141, n_16142, n_16143, n_16144,
       n_16145;
  wire n_16146, n_16147, n_16148, n_16149, n_16150, n_16151, n_16152,
       n_16153;
  wire n_16154, n_16155, n_16156, n_16157, n_16158, n_16159, n_16160,
       n_16161;
  wire n_16162, n_16163, n_16164, n_16165, n_16166, n_16167, n_16168,
       n_16169;
  wire n_16170, n_16171, n_16172, n_16173, n_16174, n_16175, n_16176,
       n_16177;
  wire n_16178, n_16179, n_16180, n_16181, n_16182, n_16183, n_16184,
       n_16185;
  wire n_16187, n_16189, n_16190, n_16191, n_16192, n_16193, n_16194,
       n_16195;
  wire n_16196, n_16197, n_16198, n_16199, n_16200, n_16201, n_16202,
       n_16203;
  wire n_16204, n_16205, n_16206, n_16207, n_16208, n_16209, n_16210,
       n_16211;
  wire n_16212, n_16213, n_16214, n_16215, n_16216, n_16217, n_16218,
       n_16219;
  wire n_16220, n_16221, n_16222, n_16223, n_16224, n_16225, n_16226,
       n_16227;
  wire n_16228, n_16229, n_16230, n_16231, n_16232, n_16233, n_16234,
       n_16235;
  wire n_16236, n_16237, n_16238, n_16239, n_16240, n_16241, n_16242,
       n_16243;
  wire n_16244, n_16245, n_16246, n_16247, n_16248, n_16249, n_16250,
       n_16251;
  wire n_16252, n_16253, n_16254, n_16255, n_16256, n_16257, n_16258,
       n_16259;
  wire n_16260, n_16261, n_16262, n_16263, n_16264, n_16265, n_16266,
       n_16267;
  wire n_16268, n_16269, n_16270, n_16271, n_16272, n_16273, n_16274,
       n_16275;
  wire n_16276, n_16277, n_16278, n_16279, n_16280, n_16281, n_16282,
       n_16283;
  wire n_16284, n_16285, n_16286, n_16287, n_16288, n_16289, n_16290,
       n_16291;
  wire n_16292, n_16293, n_16294, n_16295, n_16296, n_16297, n_16298,
       n_16299;
  wire n_16300, n_16301, n_16302, n_16303, n_16304, n_16305, n_16306,
       n_16307;
  wire n_16308, n_16309, n_16310, n_16311, n_16312, n_16313, n_16314,
       n_16315;
  wire n_16316, n_16317, n_16318, n_16319, n_16320, n_16321, n_16322,
       n_16323;
  wire n_16324, n_16325, n_16326, n_16327, n_16328, n_16329, n_16330,
       n_16331;
  wire n_16332, n_16333, n_16334, n_16335, n_16336, n_16337, n_16338,
       n_16339;
  wire n_16340, n_16341, n_16342, n_16343, n_16344, n_16345, n_16346,
       n_16347;
  wire n_16348, n_16349, n_16350, n_16351, n_16352, n_16353, n_16354,
       n_16355;
  wire n_16356, n_16357, n_16358, n_16359, n_16360, n_16361, n_16362,
       n_16363;
  wire n_16364, n_16365, n_16366, n_16367, n_16368, n_16369, n_16370,
       n_16371;
  wire n_16372, n_16373, n_16374, n_16375, n_16376, n_16377, n_16378,
       n_16379;
  wire n_16380, n_16381, n_16382, n_16383, n_16384, n_16385, n_16386,
       n_16387;
  wire n_16388, n_16389, n_16390, n_16391, n_16392, n_16393, n_16394,
       n_16395;
  wire n_16396, n_16397, n_16398, n_16399, n_16400, n_16401, n_16402,
       n_16403;
  wire n_16404, n_16405, n_16406, n_16407, n_16408, n_16409, n_16410,
       n_16411;
  wire n_16412, n_16413, n_16414, n_16415, n_16416, n_16417, n_16418,
       n_16419;
  wire n_16420, n_16421, n_16422, n_16423, n_16424, n_16425, n_16426,
       n_16427;
  wire n_16428, n_16429, n_16430, n_16431, n_16432, n_16433, n_16434,
       n_16435;
  wire n_16436, n_16437, n_16438, n_16439, n_16440, n_16441, n_16442,
       n_16443;
  wire n_16444, n_16445, n_16446, n_16447, n_16448, n_16449, n_16450,
       n_16451;
  wire n_16452, n_16453, n_16454, n_16455, n_16456, n_16457, n_16458,
       n_16459;
  wire n_16460, n_16461, n_16462, n_16463, n_16464, n_16465, n_16466,
       n_16467;
  wire n_16468, n_16469, n_16470, n_16471, n_16472, n_16473, n_16474,
       n_16475;
  wire n_16476, n_16477, n_16478, n_16479, n_16480, n_16481, n_16482,
       n_16483;
  wire n_16484, n_16485, n_16486, n_16487, n_16488, n_16489, n_16490,
       n_16491;
  wire n_16492, n_16493, n_16494, n_16495, n_16496, n_16497, n_16498,
       n_16499;
  wire n_16500, n_16501, n_16502, n_16503, n_16504, n_16505, n_16506,
       n_16507;
  wire n_16508, n_16509, n_16510, n_16511, n_16512, n_16513, n_16514,
       n_16515;
  wire n_16516, n_16517, n_16518, n_16519, n_16520, n_16521, n_16522,
       n_16523;
  wire n_16524, n_16525, n_16526, n_16527, n_16528, n_16529, n_16530,
       n_16531;
  wire n_16532, n_16533, n_16534, n_16535, n_16536, n_16537, n_16538,
       n_16539;
  wire n_16540, n_16541, n_16542, n_16543, n_16544, n_16545, n_16546,
       n_16547;
  wire n_16548, n_16549, n_16550, n_16551, n_16552, n_16553, n_16554,
       n_16555;
  wire n_16556, n_16557, n_16558, n_16559, n_16560, n_16561, n_16562,
       n_16563;
  wire n_16564, n_16565, n_16566, n_16567, n_16568, n_16569, n_16570,
       n_16571;
  wire n_16572, n_16573, n_16574, n_16575, n_16576, n_16577, n_16578,
       n_16579;
  wire n_16580, n_16581, n_16582, n_16583, n_16584, n_16585, n_16586,
       n_16587;
  wire n_16588, n_16589, n_16590, n_16591, n_16592, n_16593, n_16594,
       n_16595;
  wire n_16596, n_16597, n_16598, n_16599, n_16600, n_16601, n_16602,
       n_16603;
  wire n_16604, n_16605, n_16606, n_16607, n_16608, n_16609, n_16610,
       n_16611;
  wire n_16612, n_16613, n_16614, n_16615, n_16616, n_16617, n_16618,
       n_16619;
  wire n_16620, n_16621, n_16622, n_16623, n_16624, n_16625, n_16626,
       n_16627;
  wire n_16628, n_16629, n_16630, n_16631, n_16632, n_16633, n_16634,
       n_16635;
  wire n_16636, n_16637, n_16638, n_16639, n_16640, n_16641, n_16642,
       n_16643;
  wire n_16644, n_16645, n_16646, n_16647, n_16648, n_16649, n_16650,
       n_16651;
  wire n_16652, n_16653, n_16654, n_16655, n_16656, n_16657, n_16658,
       n_16659;
  wire n_16660, n_16661, n_16662, n_16663, n_16664, n_16665, n_16666,
       n_16667;
  wire n_16668, n_16669, n_16670, n_16671, n_16672, n_16673, n_16674,
       n_16675;
  wire n_16676, n_16677, n_16678, n_16679, n_16680, n_16681, n_16682,
       n_16683;
  wire n_16684, n_16685, n_16686, n_16687, n_16688, n_16689, n_16690,
       n_16691;
  wire n_16692, n_16693, n_16694, n_16695, n_16696, n_16697, n_16698,
       n_16699;
  wire n_16700, n_16701, n_16702, n_16703, n_16704, n_16705, n_16706,
       n_16707;
  wire n_16708, n_16709, n_16710, n_16711, n_16712, n_16713, n_16714,
       n_16715;
  wire n_16716, n_16717, n_16718, n_16719, n_16720, n_16721, n_16722,
       n_16723;
  wire n_16724, n_16725, n_16726, n_16727, n_16729, n_16730, n_16731,
       n_16732;
  wire n_16733, n_16734, n_16735, n_16736, n_16737, n_16738, n_16739,
       n_16740;
  wire n_16741, n_16742, n_16743, n_16744, n_16745, n_16746, n_16747,
       n_16748;
  wire n_16749, n_16750, n_16751, n_16752, n_16753, n_16754, n_16755,
       n_16756;
  wire n_16757, n_16758, n_16759, n_16760, n_16761, n_16762, n_16763,
       n_16764;
  wire n_16765, n_16766, n_16767, n_16768, n_16769, n_16770, n_16771,
       n_16772;
  wire n_16773, n_16774, n_16775, n_16776, n_16777, n_16778, n_16779,
       n_16780;
  wire n_16781, n_16782, n_16783, n_16784, n_16785, n_16786, n_16787,
       n_16788;
  wire n_16789, n_16790, n_16791, n_16792, n_16793, n_16794, n_16795,
       n_16796;
  wire n_16797, n_16798, n_16799, n_16800, n_16801, n_16802, n_16803,
       n_16804;
  wire n_16805, n_16806, n_16807, n_16808, n_16809, n_16810, n_16811,
       n_16812;
  wire n_16813, n_16814, n_16815, n_16816, n_16817, n_16818, n_16819,
       n_16820;
  wire n_16821, n_16822, n_16823, n_16824, n_16825, n_16826, n_16827,
       n_16828;
  wire n_16829, n_16830, n_16831, n_16832, n_16833, n_16834, n_16835,
       n_16836;
  wire n_16837, n_16838, n_16839, n_16840, n_16841, n_16842, n_16843,
       n_16844;
  wire n_16845, n_16846, n_16847, n_16848, n_16849, n_16850, n_16851,
       n_16852;
  wire n_16853, n_16854, n_16855, n_16856, n_16857, n_16858, n_16859,
       n_16860;
  wire n_16861, n_16862, n_16863, n_16864, n_16865, n_16866, n_16867,
       n_16868;
  wire n_16869, n_16870, n_16871, n_16872, n_16873, n_16874, n_16875,
       n_16876;
  wire n_16877, n_16878, n_16879, n_16880, n_16881, n_16882, n_16883,
       n_16884;
  wire n_16885, n_16886, n_16887, n_16888, n_16889, n_16890, n_16891,
       n_16892;
  wire n_16893, n_16894, n_16895, n_16896, n_16897, n_16898, n_16899,
       n_16900;
  wire n_16901, n_16902, n_16903, n_16904, n_16905, n_16906, n_16907,
       n_16908;
  wire n_16909, n_16910, n_16911, n_16912, n_16913, n_16914, n_16915,
       n_16916;
  wire n_16917, n_16918, n_16919, n_16920, n_16921, n_16922, n_16923,
       n_16924;
  wire n_16925, n_16926, n_16927, n_16928, n_16929, n_16930, n_16931,
       n_16932;
  wire n_16933, n_16934, n_16935, n_16936, n_16937, n_16938, n_16939,
       n_16940;
  wire n_16941, n_16942, n_16943, n_16944, n_16945, n_16946, n_16947,
       n_16948;
  wire n_16949, n_16950, n_16951, n_16952, n_16953, n_16954, n_16955,
       n_16956;
  wire n_16957, n_16958, n_16959, n_16960, n_16961, n_16962, n_16963,
       n_16964;
  wire n_16965, n_16966, n_16967, n_16968, n_16969, n_16970, n_16971,
       n_16972;
  wire n_16973, n_16974, n_16975, n_16976, n_16977, n_16978, n_16979,
       n_16980;
  wire n_16981, n_16982, n_16983, n_16984, n_16985, n_16986, n_16987,
       n_16988;
  wire n_16989, n_16990, n_16991, n_16992, n_16993, n_16994, n_16995,
       n_16996;
  wire n_16997, n_16998, n_16999, n_17000, n_17001, n_17002, n_17003,
       n_17004;
  wire n_17005, n_17006, n_17007, n_17008, n_17009, n_17010, n_17011,
       n_17012;
  wire n_17013, n_17014, n_17015, n_17016, n_17017, n_17018, n_17019,
       n_17020;
  wire n_17021, n_17022, n_17023, n_17024, n_17025, n_17026, n_17027,
       n_17028;
  wire n_17029, n_17030, n_17031, n_17032, n_17033, n_17034, n_17035,
       n_17036;
  wire n_17037, n_17038, n_17039, n_17040, n_17041, n_17042, n_17043,
       n_17044;
  wire n_17045, n_17046, n_17047, n_17048, n_17049, n_17050, n_17051,
       n_17052;
  wire n_17053, n_17054, n_17055, n_17056, n_17057, n_17058, n_17059,
       n_17060;
  wire n_17061, n_17062, n_17063, n_17064, n_17065, n_17066, n_17067,
       n_17068;
  wire n_17069, n_17070, n_17071, n_17072, n_17073, n_17074, n_17075,
       n_17076;
  wire n_17077, n_17078, n_17079, n_17080, n_17081, n_17082, n_17083,
       n_17084;
  wire n_17085, n_17086, n_17087, n_17088, n_17089, n_17090, n_17091,
       n_17092;
  wire n_17093, n_17094, n_17095, n_17096, n_17097, n_17098, n_17099,
       n_17100;
  wire n_17101, n_17102, n_17103, n_17104, n_17105, n_17106, n_17107,
       n_17108;
  wire n_17109, n_17110, n_17111, n_17112, n_17113, n_17114, n_17115,
       n_17116;
  wire n_17117, n_17118, n_17119, n_17120, n_17121, n_17122, n_17123,
       n_17124;
  wire n_17125, n_17126, n_17127, n_17128, n_17129, n_17130, n_17131,
       n_17132;
  wire n_17133, n_17134, n_17135, n_17136, n_17137, n_17138, n_17139,
       n_17140;
  wire n_17141, n_17142, n_17143, n_17144, n_17145, n_17146, n_17147,
       n_17148;
  wire n_17149, n_17150, n_17151, n_17152, n_17153, n_17154, n_17155,
       n_17156;
  wire n_17157, n_17158, n_17159, n_17160, n_17161, n_17162, n_17163,
       n_17164;
  wire n_17165, n_17166, n_17167, n_17168, n_17169, n_17170, n_17171,
       n_17172;
  wire n_17173, n_17174, n_17175, n_17176, n_17177, n_17178, n_17179,
       n_17180;
  wire n_17181, n_17182, n_17183, n_17184, n_17185, n_17186, n_17187,
       n_17188;
  wire n_17189, n_17190, n_17191, n_17192, n_17193, n_17194, n_17195,
       n_17199;
  wire n_17200, n_17201, n_17202, n_17203, n_17204, n_17205, n_17206,
       n_17207;
  wire n_17208, n_17209, n_17210, n_17211, n_17212, n_17213, n_17214,
       n_17215;
  wire n_17216, n_17217, n_17218, n_17219, n_17220, n_17221, n_17222,
       n_17223;
  wire n_17224, n_17225, n_17226, n_17227, n_17228, n_17229, n_17230,
       n_17231;
  wire n_17232, n_17233, n_17234, n_17235, n_17236, n_17237, n_17238,
       n_17239;
  wire n_17240, n_17241, n_17242, n_17243, n_17244, n_17245, n_17246,
       n_17247;
  wire n_17248, n_17249, n_17250, n_17251, n_17252, n_17253, n_17254,
       n_17255;
  wire n_17256, n_17257, n_17258, n_17259, n_17260, n_17261, n_17262,
       n_17263;
  wire n_17264, n_17265, n_17266, n_17267, n_17268, n_17269, n_17270,
       n_17271;
  wire n_17272, n_17273, n_17274, n_17275, n_17276, n_17277, n_17278,
       n_17279;
  wire n_17280, n_17281, n_17282, n_17283, n_17284, n_17285, n_17286,
       n_17287;
  wire n_17288, n_17289, n_17290, n_17291, n_17292, n_17293, n_17294,
       n_17295;
  wire n_17296, n_17297, n_17298, n_17299, n_17300, n_17301, n_17302,
       n_17303;
  wire n_17304, n_17305, n_17306, n_17307, n_17308, n_17309, n_17310,
       n_17311;
  wire n_17312, n_17313, n_17314, n_17315, n_17316, n_17317, n_17318,
       n_17319;
  wire n_17320, n_17321, n_17322, n_17323, n_17324, n_17325, n_17326,
       n_17327;
  wire n_17328, n_17329, n_17330, n_17331, n_17332, n_17333, n_17334,
       n_17335;
  wire n_17336, n_17337, n_17338, n_17339, n_17340, n_17341, n_17342,
       n_17343;
  wire n_17344, n_17345, n_17346, n_17347, n_17348, n_17349, n_17350,
       n_17351;
  wire n_17352, n_17353, n_17354, n_17355, n_17356, n_17357, n_17358,
       n_17359;
  wire n_17360, n_17361, n_17362, n_17363, n_17364, n_17365, n_17366,
       n_17367;
  wire n_17368, n_17369, n_17370, n_17371, n_17372, n_17373, n_17374,
       n_17375;
  wire n_17376, n_17377, n_17378, n_17379, n_17380, n_17381, n_17382,
       n_17383;
  wire n_17384, n_17385, n_17386, n_17387, n_17388, n_17389, n_17390,
       n_17391;
  wire n_17392, n_17393, n_17394, n_17395, n_17396, n_17397, n_17398,
       n_17399;
  wire n_17400, n_17401, n_17402, n_17403, n_17404, n_17405, n_17406,
       n_17407;
  wire n_17408, n_17409, n_17410, n_17411, n_17412, n_17413, n_17414,
       n_17415;
  wire n_17416, n_17417, n_17418, n_17419, n_17420, n_17421, n_17422,
       n_17423;
  wire n_17424, n_17425, n_17426, n_17427, n_17428, n_17429, n_17430,
       n_17431;
  wire n_17432, n_17433, n_17434, n_17435, n_17436, n_17437, n_17438,
       n_17439;
  wire n_17440, n_17441, n_17442, n_17443, n_17444, n_17445, n_17446,
       n_17447;
  wire n_17448, n_17449, n_17450, n_17451, n_17452, n_17453, n_17454,
       n_17455;
  wire n_17456, n_17457, n_17458, n_17459, n_17460, n_17461, n_17462,
       n_17463;
  wire n_17464, n_17465, n_17466, n_17467, n_17468, n_17469, n_17470,
       n_17471;
  wire n_17472, n_17473, n_17474, n_17475, n_17476, n_17477, n_17478,
       n_17479;
  wire n_17480, n_17481, n_17482, n_17483, n_17484, n_17485, n_17486,
       n_17487;
  wire n_17488, n_17489, n_17490, n_17491, n_17492, n_17493, n_17494,
       n_17495;
  wire n_17496, n_17497, n_17498, n_17499, n_17500, n_17501, n_17502,
       n_17503;
  wire n_17504, n_17505, n_17506, n_17507, n_17508, n_17509, n_17510,
       n_17511;
  wire n_17512, n_17513, n_17514, n_17515, n_17516, n_17517, n_17518,
       n_17519;
  wire n_17520, n_17521, n_17522, n_17523, n_17524, n_17525, n_17526,
       n_17527;
  wire n_17528, n_17529, n_17530, n_17531, n_17532, n_17533, n_17534,
       n_17535;
  wire n_17536, n_17537, n_17538, n_17539, n_17540, n_17541, n_17542,
       n_17543;
  wire n_17544, n_17545, n_17546, n_17547, n_17548, n_17549, n_17550,
       n_17551;
  wire n_17552, n_17553, n_17554, n_17555, n_17556, n_17557, n_17558,
       n_17559;
  wire n_17560, n_17561, n_17562, n_17563, n_17564, n_17565, n_17566,
       n_17567;
  wire n_17568, n_17569, n_17570, n_17571, n_17572, n_17573, n_17574,
       n_17575;
  wire n_17576, n_17577, n_17578, n_17579, n_17580, n_17581, n_17582,
       n_17583;
  wire n_17584, n_17585, n_17586, n_17587, n_17588, n_17589, n_17590,
       n_17591;
  wire n_17592, n_17593, n_17594, n_17595, n_17596, n_17597, n_17598,
       n_17599;
  wire n_17600, n_17601, n_17602, n_17603, n_17604, n_17605, n_17606,
       n_17607;
  wire n_17608, n_17609, n_17610, n_17611, n_17612, n_17613, n_17614,
       n_17615;
  wire n_17616, n_17617, n_17618, n_17619, n_17620, n_17621, n_17622,
       n_17623;
  wire n_17624, n_17625, n_17626, n_17627, n_17628, n_17629, n_17630,
       n_17631;
  wire n_17632, n_17633, n_17634, n_17635, n_17636, n_17637, n_17638,
       n_17639;
  wire n_17640, n_17641, n_17642, n_17643, n_17644, n_17645, n_17646,
       n_17647;
  wire n_17648, n_17649, n_17650, n_17651, n_17652, n_17653, n_17654,
       n_17655;
  wire n_17656, n_17657, n_17658, n_17659, n_17660, n_17661, n_17662,
       n_17663;
  wire n_17664, n_17665, n_17666, n_17667, n_17668, n_17669, n_17670,
       n_17671;
  wire n_17672, n_17673, n_17674, n_17675, n_17676, n_17677, n_17678,
       n_17679;
  wire n_17680, n_17681, n_17682, n_17683, n_17684, n_17685, n_17686,
       n_17687;
  wire n_17688, n_17689, n_17690, n_17691, n_17692, n_17693, n_17694,
       n_17695;
  wire n_17696, n_17697, n_17698, n_17699, n_17700, n_17701, n_17702,
       n_17703;
  wire n_17704, n_17705, n_17706, n_17707, n_17708, n_17709, n_17710,
       n_17711;
  wire n_17712, n_17713, n_17714, n_17715, n_17716, n_17717, n_17718,
       n_17719;
  wire n_17720, n_17721, n_17722, n_17723, n_17724, n_17725, n_17726,
       n_17727;
  wire n_17728, n_17729, n_17730, n_17731, n_17732, n_17733, n_17734,
       n_17735;
  wire n_17736, n_17737, n_17738, n_17739, n_17740, n_17741, n_17742,
       n_17743;
  wire n_17744, n_17745, n_17746, n_17747, n_17748, n_17749, n_17750,
       n_17751;
  wire n_17752, n_17753, n_17754, n_17755, n_17756, n_17757, n_17758,
       n_17759;
  wire n_17760, n_17761, n_17762, n_17763, n_17764, n_17765, n_17766,
       n_17767;
  wire n_17768, n_17769, n_17770, n_17771, n_17772, n_17773, n_17774,
       n_17775;
  wire n_17776, n_17777, n_17778, n_17779, n_17780, n_17781, n_17782,
       n_17783;
  wire n_17784, n_17785, n_17786, n_17787, n_17788, n_17789, n_17790,
       n_17791;
  wire n_17792, n_17793, n_17794, n_17795, n_17796, n_17797, n_17798,
       n_17799;
  wire n_17800, n_17801, n_17802, n_17803, n_17804, n_17805, n_17806,
       n_17807;
  wire n_17808, n_17809, n_17810, n_17811, n_17812, n_17813, n_17814,
       n_17815;
  wire n_17816, n_17817, n_17818, n_17819, n_17820, n_17821, n_17822,
       n_17823;
  wire n_17824, n_17825, n_17826, n_17827, n_17828, n_17829, n_17830,
       n_17831;
  wire n_17832, n_17833, n_17834, n_17835, n_17836, n_17837, n_17838,
       n_17839;
  wire n_17840, n_17841, n_17842, n_17843, n_17844, n_17845, n_17846,
       n_17847;
  wire n_17848, n_17849, n_17850, n_17851, n_17852, n_17853, n_17854,
       n_17855;
  wire n_17856, n_17857, n_17858, n_17859, n_17860, n_17861, n_17862,
       n_17863;
  wire n_17864, n_17865, n_17866, n_17867, n_17868, n_17869, n_17870,
       n_17871;
  wire n_17872, n_17873, n_17874, n_17875, n_17876, n_17877, n_17878,
       n_17879;
  wire n_17880, n_17881, n_17882, n_17883, n_17884, n_17885, n_17886,
       n_17887;
  wire n_17888, n_17889, n_17890, n_17891, n_17892, n_17893, n_17894,
       n_17895;
  wire n_17896, n_17897, n_17898, n_17899, n_17900, n_17901, n_17902,
       n_17903;
  wire n_17904, n_17905, n_17906, n_17907, n_17908, n_17909, n_17910,
       n_17911;
  wire n_17912, n_17913, n_17914, n_17915, n_17916, n_17917, n_17918,
       n_17919;
  wire n_17920, n_17921, n_17922, n_17923, n_17924, n_17925, n_17926,
       n_17927;
  wire n_17928, n_17929, n_17930, n_17931, n_17932, n_17933, n_17934,
       n_17935;
  wire n_17936, n_17937, n_17938, n_17939, n_17940, n_17941, n_17942,
       n_17943;
  wire n_17944, n_17945, n_17946, n_17947, n_17948, n_17949, n_17950,
       n_17951;
  wire n_17952, n_17953, n_17954, n_17955, n_17956, n_17957, n_17958,
       n_17959;
  wire n_17960, n_17961, n_17962, n_17963, n_17964, n_17965, n_17966,
       n_17967;
  wire n_17968, n_17969, n_17970, n_17971, n_17972, n_17973, n_17974,
       n_17975;
  wire n_17976, n_17977, n_17978, n_17979, n_17980, n_17981, n_17982,
       n_17983;
  wire n_17984, n_17985, n_17986, n_17987, n_17988, n_17989, n_17990,
       n_17991;
  wire n_17992, n_17993, n_17994, n_17995, n_17996, n_17997, n_17998,
       n_17999;
  wire n_18000, n_18001, n_18002, n_18003, n_18004, n_18005, n_18006,
       n_18007;
  wire n_18008, n_18009, n_18010, n_18011, n_18012, n_18013, n_18014,
       n_18015;
  wire n_18016, n_18017, n_18018, n_18019, n_18020, n_18021, n_18022,
       n_18023;
  wire n_18024, n_18025, n_18026, n_18027, n_18028, n_18029, n_18030,
       n_18031;
  wire n_18032, n_18033, n_18034, n_18035, n_18036, n_18037, n_18038,
       n_18039;
  wire n_18040, n_18041, n_18042, n_18043, n_18044, n_18045, n_18046,
       n_18047;
  wire n_18048, n_18049, n_18050, n_18051, n_18052, n_18053, n_18054,
       n_18055;
  wire n_18056, n_18057, n_18058, n_18059, n_18060, n_18061, n_18062,
       n_18063;
  wire n_18064, n_18065, n_18066, n_18067, n_18068, n_18069, n_18070,
       n_18071;
  wire n_18072, n_18073, n_18074, n_18075, n_18076, n_18077, n_18078,
       n_18079;
  wire n_18080, n_18081, n_18082, n_18083, n_18084, n_18085, n_18086,
       n_18087;
  wire n_18088, n_18089, n_18090, n_18091, n_18092, n_18093, n_18094,
       n_18095;
  wire n_18096, n_18097, n_18098, n_18099, n_18100, n_18101, n_18102,
       n_18103;
  wire n_18104, n_18105, n_18106, n_18107, n_18108, n_18109, n_18110,
       n_18111;
  wire n_18112, n_18113, n_18114, n_18115, n_18116, n_18117, n_18118,
       n_18119;
  wire n_18120, n_18121, n_18122, n_18123, n_18124, n_18125, n_18126,
       n_18127;
  wire n_18128, n_18129, n_18130, n_18131, n_18132, n_18133, n_18134,
       n_18135;
  wire n_18136, n_18137, n_18138, n_18139, n_18140, n_18141, n_18142,
       n_18143;
  wire n_18144, n_18145, n_18146, n_18147, n_18148, n_18149, n_18150,
       n_18151;
  wire n_18152, n_18153, n_18154, n_18155, n_18156, n_18157, n_18158,
       n_18159;
  wire n_18160, n_18161, n_18162, n_18163, n_18164, n_18165, n_18166,
       n_18167;
  wire n_18168, n_18169, n_18170, n_18171, n_18172, n_18173, n_18174,
       n_18175;
  wire n_18176, n_18177, n_18178, n_18179, n_18180, n_18181, n_18182,
       n_18183;
  wire n_18184, n_18185, n_18186, n_18187, n_18188, n_18189, n_18190,
       n_18191;
  wire n_18192, n_18193, n_18194, n_18195, n_18196, n_18197, n_18198,
       n_18199;
  wire n_18200, n_18201, n_18202, n_18203, n_18204, n_18205, n_18206,
       n_18207;
  wire n_18208, n_18209, n_18210, n_18211, n_18212, n_18213, n_18214,
       n_18215;
  wire n_18216, n_18217, n_18218, n_18219, n_18220, n_18221, n_18222,
       n_18223;
  wire n_18224, n_18225, n_18226, n_18227, n_18228, n_18229, n_18230,
       n_18231;
  wire n_18232, n_18233, n_18234, n_18235, n_18236, n_18237, n_18238,
       n_18239;
  wire n_18240, n_18241, n_18242, n_18243, n_18244, n_18245, n_18246,
       n_18247;
  wire n_18248, n_18249, n_18250, n_18251, n_18252, n_18253, n_18254,
       n_18255;
  wire n_18256, n_18257, n_18258, n_18259, n_18260, n_18261, n_18262,
       n_18263;
  wire n_18264, n_18265, n_18266, n_18267, n_18268, n_18269, n_18270,
       n_18271;
  wire n_18272, n_18273, n_18274, n_18275, n_18276, n_18277, n_18278,
       n_18279;
  wire n_18280, n_18281, n_18282, n_18283, n_18284, n_18285, n_18286,
       n_18287;
  wire n_18288, n_18289, n_18290, n_18291, n_18292, n_18293, n_18294,
       n_18295;
  wire n_18296, n_18297, n_18298, n_18299, n_18300, n_18301, n_18302,
       n_18303;
  wire n_18304, n_18305, n_18306, n_18307, n_18308, n_18309, n_18310,
       n_18311;
  wire n_18312, n_18313, n_18314, n_18315, n_18316, n_18317, n_18318,
       n_18319;
  wire n_18320, n_18321, n_18322, n_18323, n_18324, n_18325, n_18326,
       n_18327;
  wire n_18328, n_18329, n_18330, n_18331, n_18332, n_18333, n_18334,
       n_18335;
  wire n_18336, n_18337, n_18338, n_18339, n_18340, n_18341, n_18342,
       n_18343;
  wire n_18344, n_18345, n_18346, n_18347, n_18348, n_18349, n_18350,
       n_18351;
  wire n_18352, n_18353, n_18354, n_18355, n_18356, n_18357, n_18358,
       n_18359;
  wire n_18360, n_18361, n_18362, n_18363, n_18364, n_18365, n_18366,
       n_18367;
  wire n_18368, n_18369, n_18370, n_18371, n_18372, n_18373, n_18374,
       n_18375;
  wire n_18376, n_18377, n_18378, n_18379, n_18380, n_18381, n_18382,
       n_18383;
  wire n_18384, n_18385, n_18386, n_18387, n_18388, n_18389, n_18390,
       n_18391;
  wire n_18392, n_18393, n_18394, n_18395, n_18396, n_18397, n_18398,
       n_18399;
  wire n_18400, n_18401, n_18402, n_18403, n_18404, n_18405, n_18406,
       n_18407;
  wire n_18408, n_18409, n_18410, n_18411, n_18412, n_18413, n_18414,
       n_18415;
  wire n_18416, n_18417, n_18418, n_18419, n_18420, n_18421, n_18422,
       n_18423;
  wire n_18424, n_18425, n_18426, n_18427, n_18428, n_18429, n_18430,
       n_18431;
  wire n_18432, n_18433, n_18434, n_18435, n_18436, n_18437, n_18438,
       n_18439;
  wire n_18440, n_18441, n_18442, n_18443, n_18444, n_18445, n_18446,
       n_18447;
  wire n_18448, n_18449, n_18450, n_18451, n_18452, n_18453, n_18454,
       n_18455;
  wire n_18456, n_18457, n_18458, n_18459, n_18460, n_18461, n_18462,
       n_18463;
  wire n_18464, n_18465, n_18466, n_18467, n_18468, n_18469, n_18470,
       n_18471;
  wire n_18472, n_18473, n_18474, n_18475, n_18476, n_18477, n_18478,
       n_18479;
  wire n_18480, n_18481, n_18482, n_18483, n_18484, n_18485, n_18486,
       n_18487;
  wire n_18488, n_18489, n_18490, n_18491, n_18492, n_18493, n_18494,
       n_18495;
  wire n_18496, n_18497, n_18498, n_18499, n_18500, n_18501, n_18502,
       n_18503;
  wire n_18504, n_18505, n_18506, n_18507, n_18508, n_18509, n_18510,
       n_18511;
  wire n_18512, n_18513, n_18514, n_18515, n_18516, n_18517, n_18518,
       n_18519;
  wire n_18520, n_18521, n_18522, n_18523, n_18524, n_18525, n_18526,
       n_18527;
  wire n_18528, n_18529, n_18530, n_18531, n_18532, n_18533, n_18534,
       n_18535;
  wire n_18536, n_18537, n_18538, n_18539, n_18540, n_18541, n_18542,
       n_18543;
  wire n_18544, n_18545, n_18546, n_18547, n_18548, n_18549, n_18550,
       n_18551;
  wire n_18552, n_18553, n_18554, n_18555, n_18556, n_18557, n_18558,
       n_18559;
  wire n_18560, n_18561, n_18562, n_18563, n_18564, n_18565, n_18566,
       n_18567;
  wire n_18568, n_18569, n_18570, n_18571, n_18572, n_18573, n_18574,
       n_18575;
  wire n_18576, n_18577, n_18578, n_18579, n_18580, n_18581, n_18582,
       n_18583;
  wire n_18584, n_18585, n_18586, n_18587, n_18588, n_18589, n_18590,
       n_18591;
  wire n_18592, n_18593, n_18594, n_18595, n_18596, n_18597, n_18598,
       n_18599;
  wire n_18600, n_18601, n_18602, n_18603, n_18604, n_18605, n_18606,
       n_18607;
  wire n_18608, n_18609, n_18610, n_18611, n_18612, n_18613, n_18614,
       n_18615;
  wire n_18616, n_18617, n_18618, n_18619, n_18620, n_18621, n_18622,
       n_18623;
  wire n_18624, n_18625, n_18626, n_18627, n_18628, n_18629, n_18630,
       n_18631;
  wire n_18632, n_18633, n_18634, n_18635, n_18636, n_18637, n_18638,
       n_18639;
  wire n_18640, n_18641, n_18642, n_18643, n_18644, n_18645, n_18646,
       n_18647;
  wire n_18648, n_18649, n_18650, n_18651, n_18652, n_18653, n_18654,
       n_18655;
  wire n_18656, n_18657, n_18658, n_18659, n_18660, n_18661, n_18662,
       n_18663;
  wire n_18664, n_18665, n_18666, n_18667, n_18668, n_18669, n_18670,
       n_18671;
  wire n_18672, n_18673, n_18674, n_18675, n_18676, n_18677, n_18678,
       n_18679;
  wire n_18680, n_18681, n_18682, n_18683, n_18684, n_18685, n_18686,
       n_18687;
  wire n_18688, n_18689, n_18690, n_18691, n_18692, n_18693, n_18694,
       n_18695;
  wire n_18696, n_18697, n_18698, n_18699, n_18700, n_18701, n_18702,
       n_18703;
  wire n_18704, n_18705, n_18706, n_18707, n_18708, n_18709, n_18710,
       n_18711;
  wire n_18712, n_18713, n_18714, n_18715, n_18716, n_18717, n_18718,
       n_18719;
  wire n_18720, n_18721, n_18722, n_18723, n_18724, n_18725, n_18726,
       n_18727;
  wire n_18728, n_18729, n_18730, n_18731, n_18732, n_18733, n_18734,
       n_18735;
  wire n_18736, n_18737, n_18738, n_18739, n_18740, n_18741, n_18742,
       n_18743;
  wire n_18744, n_18745, n_18746, n_18747, n_18748, n_18749, n_18750,
       n_18751;
  wire n_18752, n_18753, n_18754, n_18755, n_18756, n_18757, n_18758,
       n_18759;
  wire n_18760, n_18761, n_18762, n_18763, n_18764, n_18765, n_18766,
       n_18767;
  wire n_18768, n_18769, n_18770, n_18771, n_18772, n_18773, n_18774,
       n_18775;
  wire n_18776, n_18777, n_18778, n_18779, n_18780, n_18781, n_18782,
       n_18783;
  wire n_18784, n_18785, n_18786, n_18787, n_18788, n_18789, n_18790,
       n_18791;
  wire n_18792, n_18793, n_18794, n_18795, n_18796, n_18797, n_18798,
       n_18799;
  wire n_18800, n_18801, n_18802, n_18803, n_18804, n_18805, n_18806,
       n_18807;
  wire n_18808, n_18809, n_18810, n_18811, n_18812, n_18813, n_18814,
       n_18815;
  wire n_18816, n_18817, n_18818, n_18819, n_18820, n_18821, n_18822,
       n_18823;
  wire n_18824, n_18825, n_18826, n_18827, n_18828, n_18829, n_18830,
       n_18831;
  wire n_18832, n_18833, n_18834, n_18835, n_18836, n_18837, n_18838,
       n_18839;
  wire n_18840, n_18841, n_18842, n_18843, n_18844, n_18845, n_18846,
       n_18847;
  wire n_18848, n_18849, n_18850, n_18851, n_18852, n_18853, n_18854,
       n_18855;
  wire n_18856, n_18857, n_18858, n_18859, n_18860, n_18861, n_18862,
       n_18863;
  wire n_18864, n_18865, n_18866, n_18867, n_18868, n_18869, n_18870,
       n_18871;
  wire n_18872, n_18873, n_18874, n_18875, n_18876, n_18877, n_18878,
       n_18879;
  wire n_18880, n_18881, n_18882, n_18883, n_18884, n_18885, n_18886,
       n_18887;
  wire n_18888, n_18889, n_18890, n_18891, n_18892, n_18893, n_18894,
       n_18895;
  wire n_18896, n_18897, n_18898, n_18899, n_18900, n_18901, n_18902,
       n_18903;
  wire n_18904, n_18905, n_18906, n_18907, n_18908, n_18909, n_18910,
       n_18911;
  wire n_18912, n_18913, n_18914, n_18915, n_18916, n_18917, n_18918,
       n_18919;
  wire n_18920, n_18921, n_18922, n_18923, n_18924, n_18925, n_18926,
       n_18927;
  wire n_18928, n_18929, n_18930, n_18931, n_18932, n_18933, n_18934,
       n_18935;
  wire n_18936, n_18937, n_18938, n_18939, n_18940, n_18941, n_18942,
       n_18943;
  wire n_18944, n_18945, n_18946, n_18947, n_18948, n_18949, n_18950,
       n_18951;
  wire n_18952, n_18953, n_18954, n_18955, n_18956, n_18957, n_18958,
       n_18959;
  wire n_18960, n_18961, n_18962, n_18963, n_18964, n_18965, n_18966,
       n_18967;
  wire n_18968, n_18969, n_18970, n_18971, n_18972, n_18973, n_18974,
       n_18975;
  wire n_18976, n_18977, n_18978, n_18979, n_18980, n_18981, n_18982,
       n_18983;
  wire n_18984, n_18985, n_18986, n_18987, n_18988, n_18989, n_18990,
       n_18991;
  wire n_18992, n_18993, n_18994, n_18995, n_18996, n_18997, n_18998,
       n_18999;
  wire n_19000, n_19001, n_19002, n_19003, n_19004, n_19005, n_19006,
       n_19007;
  wire n_19008, n_19009, n_19010, n_19011, n_19012, n_19013, n_19014,
       n_19015;
  wire n_19016, n_19017, n_19018, n_19019, n_19020, n_19021, n_19022,
       n_19023;
  wire n_19024, n_19025, n_19026, n_19027, n_19028, n_19029, n_19030,
       n_19031;
  wire n_19032, n_19033, n_19034, n_19035, n_19036, n_19037, n_19038,
       n_19039;
  wire n_19040, n_19041, n_19042, n_19043, n_19044, n_19045, n_19046,
       n_19047;
  wire n_19048, n_19049, n_19050, n_19051, n_19052, n_19053, n_19054,
       n_19055;
  wire n_19056, n_19057, n_19058, n_19059, n_19060, n_19061, n_19062,
       n_19063;
  wire n_19064, n_19065, n_19066, n_19067, n_19068, n_19073, n_19074,
       n_19075;
  wire n_19076, n_19077, n_19078, n_19079, n_19080, n_19081, n_19082,
       n_19083;
  wire n_19084, n_19085, n_19086, n_19087, n_19088, n_19089, n_19090,
       n_19091;
  wire n_19092, n_19093, n_19094, n_19095, n_19096, n_19097, n_19098,
       n_19099;
  wire n_19100, n_19101, n_19102, n_19103, n_19104, n_19105, n_19106,
       n_19107;
  wire n_19108, n_19109, n_19110, n_19111, n_19112, n_19113, n_19114,
       n_19115;
  wire n_19116, n_19117, n_19118, n_19119, n_19120, n_19121, n_19122,
       n_19123;
  wire n_19124, n_19125, n_19126, n_19127, n_19128, n_19129, n_19130,
       n_19131;
  wire n_19132, n_19133, n_19134, n_19135, n_19136, n_19137, n_19138,
       n_19139;
  wire n_19140, n_19141, n_19142, n_19143, n_19144, n_19145, n_19146,
       n_19147;
  wire n_19148, n_19149, n_19150, n_19151, n_19152, n_19153, n_19154,
       n_19155;
  wire n_19156, n_19157, n_19158, n_19159, n_19160, n_19161, n_19162,
       n_19163;
  wire n_19164, n_19165, n_19166, n_19167, n_19168, n_19169, n_19170,
       n_19171;
  wire n_19172, n_19173, n_19174, n_19175, n_19176, n_19177, n_19178,
       n_19179;
  wire n_19180, n_19181, n_19182, n_19183, n_19184, n_19185, n_19186,
       n_19187;
  wire n_19188, n_19189, n_19190, n_19191, n_19192, n_19193, n_19194,
       n_19195;
  wire n_19196, n_19197, n_19198, n_19199, n_19200, n_19201, n_19202,
       n_19203;
  wire n_19204, n_19205, n_19206, n_19207, n_19208, n_19209, n_19210,
       n_19211;
  wire n_19212, n_19213, n_19214, n_19215, n_19216, n_19217, n_19218,
       n_19219;
  wire n_19220, n_19221, n_19222, n_19223, n_19224, n_19225, n_19226,
       n_19227;
  wire n_19228, n_19229, n_19230, n_19231, n_19232, n_19233, n_19234,
       n_19235;
  wire n_19236, n_19237, n_19238, n_19239, n_19240, n_19241, n_19242,
       n_19243;
  wire n_19244, n_19245, n_19246, n_19247, n_19248, n_19249, n_19250,
       n_19251;
  wire n_19252, n_19253, n_19254, n_19255, n_19256, n_19257, n_19258,
       n_19259;
  wire n_19260, n_19261, n_19262, n_19263, n_19264, n_19265, n_19266,
       n_19267;
  wire n_19268, n_19269, n_19270, n_19271, n_19272, n_19273, n_19274,
       n_19275;
  wire n_19276, n_19277, n_19278, n_19279, n_19280, n_19281, n_19282,
       n_19283;
  wire n_19284, n_19285, n_19286, n_19287, n_19288, n_19289, n_19290,
       n_19291;
  wire n_19292, n_19293, n_19294, n_19295, n_19296, n_19297, n_19298,
       n_19299;
  wire n_19300, n_19301, n_19302, n_19303, n_19304, n_19305, n_19306,
       n_19307;
  wire n_19308, n_19309, n_19310, n_19311, n_19312, n_19313, n_19314,
       n_19315;
  wire n_19316, n_19317, n_19318, n_19319, n_19320, n_19321, n_19322,
       n_19323;
  wire n_19324, n_19325, n_19326, n_19327, n_19328, n_19329, n_19330,
       n_19331;
  wire n_19332, n_19333, n_19334, n_19335, n_19336, n_19337, n_19338,
       n_19339;
  wire n_19340, n_19341, n_19342, n_19343, n_19344, n_19345, n_19346,
       n_19347;
  wire n_19348, n_19349, n_19350, n_19351, n_19352, n_19353, n_19354,
       n_19355;
  wire n_19356, n_19357, n_19358, n_19359, n_19360, n_19361, n_19362,
       n_19363;
  wire n_19364, n_19365, n_19366, n_19367, n_19368, n_19369, n_19370,
       n_19371;
  wire n_19372, n_19373, n_19374, n_19375, n_19376, n_19377, n_19378,
       n_19379;
  wire n_19380, n_19381, n_19382, n_19383, n_19384, n_19385, n_19386,
       n_19387;
  wire n_19388, n_19389, n_19390, n_19391, n_19392, n_19393, n_19394,
       n_19395;
  wire n_19396, n_19397, n_19398, n_19399, n_19400, n_19401, n_19402,
       n_19403;
  wire n_19404, n_19405, n_19406, n_19407, n_19408, n_19409, n_19410,
       n_19411;
  wire n_19412, n_19413, n_19414, n_19415, n_19416, n_19417, n_19418,
       n_19419;
  wire n_19420, n_19421, n_19422, n_19423, n_19424, n_19425, n_19426,
       n_19427;
  wire n_19428, n_19429, n_19430, n_19431, n_19432, n_19433, n_19434,
       n_19435;
  wire n_19436, n_19437, n_19438, n_19439, n_19440, n_19441, n_19442,
       n_19443;
  wire n_19444, n_19445, n_19446, n_19447, n_19448, n_19453, n_19454,
       n_19455;
  wire n_19456, n_19457, n_19458, n_19459, n_19460, n_19461, n_19462,
       n_19463;
  wire n_19464, n_19465, n_19466, n_19467, n_19468, n_19469, n_19470,
       n_19471;
  wire n_19472, n_19473, n_19474, n_19475, n_19476, n_19477, n_19478,
       n_19479;
  wire n_19480, n_19481, n_19482, n_19483, n_19484, n_19485, n_19486,
       n_19487;
  wire n_19488, n_19489, n_19490, n_19491, n_19492, n_19493, n_19494,
       n_19495;
  wire n_19496, n_19497, n_19498, n_19499, n_19500, n_19501, n_19502,
       n_19503;
  wire n_19504, n_19505, n_19506, n_19507, n_19508, n_19509, n_19510,
       n_19511;
  wire n_19512, n_19513, n_19514, n_19515, n_19516, n_19517, n_19518,
       n_19519;
  wire n_19520, n_19521, n_19522, n_19523, n_19524, n_19525, n_19526,
       n_19527;
  wire n_19528, n_19529, n_19530, n_19531, n_19532, n_19533, n_19534,
       n_19535;
  wire n_19536, n_19537, n_19538, n_19539, n_19540, n_19541, n_19542,
       n_19543;
  wire n_19544, n_19545, n_19546, n_19547, n_19548, n_19549, n_19550,
       n_19551;
  wire n_19552, n_19553, n_19554, n_19555, n_19556, n_19557, n_19558,
       n_19559;
  wire n_19560, n_19561, n_19562, n_19563, n_19564, n_19565, n_19566,
       n_19567;
  wire n_19568, n_19569, n_19570, n_19571, n_19572, n_19573, n_19574,
       n_19575;
  wire n_19576, n_19577, n_19578, n_19579, n_19580, n_19581, n_19582,
       n_19583;
  wire n_19584, n_19585, n_19586, n_19587, n_19588, n_19589, n_19590,
       n_19591;
  wire n_19592, n_19593, n_19594, n_19595, n_19596, n_19597, n_19598,
       n_19599;
  wire n_19600, n_19601, n_19602, n_19603, n_19604, n_19605, n_19606,
       n_19607;
  wire n_19608, n_19609, n_19610, n_19611, n_19612, n_19613, n_19614,
       n_19615;
  wire n_19616, n_19617, n_19618, n_19619, n_19620, n_19621, n_19622,
       n_19623;
  wire n_19624, n_19625, n_19626, n_19627, n_19628, n_19629, n_19630,
       n_19631;
  wire n_19632, n_19633, n_19634, n_19635, n_19636, n_19637, n_19638,
       n_19639;
  wire n_19640, n_19641, n_19642, n_19643, n_19644, n_19645, n_19646,
       n_19647;
  wire n_19648, n_19649, n_19650, n_19651, n_19652, n_19653, n_19654,
       n_19655;
  wire n_19656, n_19657, n_19658, n_19659, n_19660, n_19661, n_19662,
       n_19663;
  wire n_19664, n_19665, n_19666, n_19667, n_19668, n_19669, n_19670,
       n_19671;
  wire n_19672, n_19673, n_19674, n_19675, n_19676, n_19677, n_19678,
       n_19679;
  wire n_19680, n_19681, n_19682, n_19683, n_19684, n_19685, n_19686,
       n_19687;
  wire n_19688, n_19689, n_19690, n_19691, n_19692, n_19693, n_19694,
       n_19695;
  wire n_19696, n_19697, n_19698, n_19699, n_19700, n_19701, n_19702,
       n_19703;
  wire n_19704, n_19705, n_19706, n_19707, n_19708, n_19709, n_19710,
       n_19711;
  wire n_19712, n_19713, n_19714, n_19715, n_19716, n_19717, n_19718,
       n_19719;
  wire n_19720, n_19721, n_19722, n_19723, n_19724, n_19725, n_19726,
       n_19727;
  wire n_19728, n_19729, n_19730, n_19731, n_19732, n_19733, n_19734,
       n_19735;
  wire n_19736, n_19737, n_19738, n_19739, n_19740, n_19741, n_19742,
       n_19743;
  wire n_19744, n_19745, n_19746, n_19747, n_19748, n_19749, n_19750,
       n_19751;
  wire n_19752, n_19753, n_19754, n_19755, n_19756, n_19757, n_19758,
       n_19759;
  wire n_19760, n_19761, n_19762, n_19763, n_19764, n_19765, n_19766,
       n_19767;
  wire n_19768, n_19769, n_19770, n_19771, n_19772, n_19773, n_19774,
       n_19775;
  wire n_19776, n_19777, n_19778, n_19779, n_19780, n_19781, n_19782,
       n_19783;
  wire n_19784, n_19785, n_19786, n_19787, n_19788, n_19789, n_19790,
       n_19791;
  wire n_19792, n_19793, n_19794, n_19795, n_19796, n_19797, n_19798,
       n_19799;
  wire n_19800, n_19801, n_19802, n_19803, n_19804, n_19805, n_19806,
       n_19807;
  wire n_19808, n_19809, n_19810, n_19811, n_19812, n_19813, n_19814,
       n_19815;
  wire n_19816, n_19817, n_19818, n_19819, n_19820, n_19821, n_19822,
       n_19823;
  wire n_19824, n_19825, n_19826, n_19827, n_19828, n_19829, n_19830,
       n_19831;
  wire n_19832, n_19833, n_19834, n_19835, n_19836, n_19837, n_19838,
       n_19839;
  wire n_19840, n_19841, n_19842, n_19843, n_19844, n_19845, n_19846,
       n_19847;
  wire n_19848, n_19849, n_19850, n_19851, n_19852, n_19853, n_19854,
       n_19855;
  wire n_19856, n_19857, n_19858, n_19859, n_19860, n_19861, n_19862,
       n_19863;
  wire n_19864, n_19865, n_19866, n_19867, n_19868, n_19869, n_19870,
       n_19871;
  wire n_19872, n_19873, n_19874, n_19875, n_19876, n_19877, n_19878,
       n_19879;
  wire n_19880, n_19881, n_19882, n_19883, n_19884, n_19885, n_19886,
       n_19887;
  wire n_19888, n_19889, n_19890, n_19891, n_19892, n_19893, n_19894,
       n_19895;
  wire n_19896, n_19897, n_19898, n_19899, n_19900, n_19901, n_19902,
       n_19903;
  wire n_19904, n_19905, n_19906, n_19907, n_19908, n_19909, n_19910,
       n_19911;
  wire n_19912, n_19913, n_19914, n_19915, n_19916, n_19917, n_19918,
       n_19919;
  wire n_19920, n_19921, n_19922, n_19923, n_19924, n_19925, n_19926,
       n_19927;
  wire n_19928, n_19929, n_19930, n_19931, n_19932, n_19933, n_19934,
       n_19935;
  wire n_19936, n_19937, n_19938, n_19939, n_19940, n_19941, n_19942,
       n_19943;
  wire n_19944, n_19945, n_19946, n_19947, n_19948, n_19949, n_19950,
       n_19951;
  wire n_19952, n_19953, n_19954, n_19955, n_19956, n_19957, n_19958,
       n_19959;
  wire n_19960, n_19961, n_19962, n_19963, n_19964, n_19965, n_19966,
       n_19967;
  wire n_19968, n_19969, n_19970, n_19971, n_19972, n_19973, n_19974,
       n_19975;
  wire n_19976, n_19977, n_19978, n_19979, n_19980, n_19981, n_19982,
       n_19983;
  wire n_19984, n_19985, n_19986, n_19987, n_19988, n_19989, n_19990,
       n_19991;
  wire n_19992, n_19993, n_19994, n_19995, n_19996, n_19997, n_19998,
       n_19999;
  wire n_20000, n_20001, n_20002, n_20003, n_20004, n_20005, n_20006,
       n_20007;
  wire n_20008, n_20009, n_20010, n_20011, n_20012, n_20013, n_20014,
       n_20015;
  wire n_20016, n_20017, n_20018, n_20019, n_20020, n_20021, n_20022,
       n_20023;
  wire n_20024, n_20025, n_20026, n_20027, n_20028, n_20029, n_20030,
       n_20031;
  wire n_20032, n_20033, n_20034, n_20035, n_20036, n_20037, n_20038,
       n_20039;
  wire n_20040, n_20041, n_20042, n_20043, n_20044, n_20045, n_20046,
       n_20047;
  wire n_20048, n_20049, n_20050, n_20051, n_20052, n_20053, n_20054,
       n_20055;
  wire n_20056, n_20057, n_20058, n_20059, n_20060, n_20061, n_20062,
       n_20063;
  wire n_20064, n_20065, n_20066, n_20067, n_20068, n_20069, n_20070,
       n_20071;
  wire n_20072, n_20073, n_20074, n_20075, n_20076, n_20077, n_20078,
       n_20079;
  wire n_20080, n_20081, n_20082, n_20083, n_20084, n_20085, n_20086,
       n_20087;
  wire n_20088, n_20089, n_20090, n_20091, n_20092, n_20093, n_20094,
       n_20095;
  wire n_20096, n_20097, n_20098, n_20099, n_20100, n_20101, n_20102,
       n_20103;
  wire n_20104, n_20105, n_20106, n_20107, n_20108, n_20109, n_20110,
       n_20111;
  wire n_20112, n_20113, n_20114, n_20115, n_20116, n_20117, n_20118,
       n_20119;
  wire n_20120, n_20121, n_20122, n_20123, n_20124, n_20125, n_20126,
       n_20127;
  wire n_20128, n_20129, n_20130, n_20131, n_20132, n_20133, n_20134,
       n_20135;
  wire n_20136, n_20137, n_20138, n_20139, n_20140, n_20141, n_20142,
       n_20143;
  wire n_20144, n_20145, n_20146, n_20147, n_20148, n_20149, n_20150,
       n_20151;
  wire n_20152, n_20153, n_20154, n_20155, n_20156, n_20157, n_20158,
       n_20159;
  wire n_20160, n_20161, n_20162, n_20163, n_20164, n_20165, n_20166,
       n_20167;
  wire n_20168, n_20169, n_20170, n_20171, n_20172, n_20173, n_20174,
       n_20175;
  wire n_20176, n_20177, n_20178, n_20179, n_20180, n_20181, n_20182,
       n_20183;
  wire n_20184, n_20185, n_20186, n_20187, n_20188, n_20189, n_20190,
       n_20191;
  wire n_20192, n_20193, n_20194, n_20195, n_20196, n_20197, n_20198,
       n_20199;
  wire n_20200, n_20201, n_20202, n_20203, n_20204, n_20205, n_20206,
       n_20207;
  wire n_20208, n_20209, n_20210, n_20211, n_20212, n_20213, n_20214,
       n_20215;
  wire n_20216, n_20217, n_20218, n_20219, n_20220, n_20221, n_20222,
       n_20223;
  wire n_20224, n_20225, n_20226, n_20227, n_20228, n_20229, n_20230,
       n_20231;
  wire n_20232, n_20233, n_20234, n_20235, n_20236, n_20237, n_20238,
       n_20239;
  wire n_20240, n_20241, n_20242, n_20243, n_20244, n_20245, n_20246,
       n_20247;
  wire n_20248, n_20249, n_20250, n_20251, n_20252, n_20253, n_20254,
       n_20255;
  wire n_20256, n_20257, n_20258, n_20259, n_20260, n_20261, n_20262,
       n_20263;
  wire n_20264, n_20265, n_20266, n_20267, n_20268, n_20269, n_20270,
       n_20271;
  wire n_20272, n_20273, n_20274, n_20275, n_20276, n_20277, n_20278,
       n_20279;
  wire n_20280, n_20281, n_20282, n_20283, n_20284, n_20285, n_20286,
       n_20287;
  wire n_20288, n_20289, n_20290, n_20291, n_20292, n_20293, n_20294,
       n_20295;
  wire n_20296, n_20297, n_20298, n_20299, n_20300, n_20301, n_20302,
       n_20303;
  wire n_20304, n_20305, n_20306, n_20307, n_20308, n_20309, n_20310,
       n_20311;
  wire n_20312, n_20313, n_20314, n_20315, n_20316, n_20317, n_20318,
       n_20319;
  wire n_20320, n_20321, n_20322, n_20323, n_20324, n_20325, n_20326,
       n_20327;
  wire n_20328, n_20329, n_20330, n_20331, n_20332, n_20333, n_20334,
       n_20335;
  wire n_20336, n_20337, n_20338, n_20339, n_20340, n_20341, n_20342,
       n_20343;
  wire n_20344, n_20345, n_20346, n_20347, n_20348, n_20349, n_20350,
       n_20351;
  wire n_20352, n_20353, n_20354, n_20355, n_20356, n_20357, n_20358,
       n_20359;
  wire n_20360, n_20361, n_20362, n_20363, n_20364, n_20365, n_20366,
       n_20367;
  wire n_20368, n_20369, n_20370, n_20371, n_20372, n_20373, n_20374,
       n_20375;
  wire n_20376, n_20377, n_20378, n_20379, n_20380, n_20381, n_20382,
       n_20383;
  wire n_20384, n_20385, n_20386, n_20387, n_20388, n_20389, n_20390,
       n_20391;
  wire n_20392, n_20393, n_20394, n_20395, n_20396, n_20397, n_20398,
       n_20399;
  wire n_20400, n_20401, n_20402, n_20403, n_20404, n_20405, n_20406,
       n_20407;
  wire n_20408, n_20409, n_20410, n_20411, n_20412, n_20413, n_20414,
       n_20415;
  wire n_20416, n_20417, n_20418, n_20419, n_20420, n_20421, n_20422,
       n_20423;
  wire n_20424, n_20425, n_20426, n_20427, n_20428, n_20429, n_20430,
       n_20431;
  wire n_20432, n_20433, n_20434, n_20435, n_20436, n_20437, n_20438,
       n_20439;
  wire n_20440, n_20441, n_20442, n_20443, n_20444, n_20445, n_20446,
       n_20447;
  wire n_20448, n_20449, n_20450, n_20451, n_20452, n_20453, n_20454,
       n_20455;
  wire n_20456, n_20457, n_20458, n_20459, n_20460, n_20461, n_20462,
       n_20463;
  wire n_20464, n_20465, n_20466, n_20467, n_20468, n_20469, n_20470,
       n_20471;
  wire n_20472, n_20473, n_20474, n_20475, n_20476, n_20477, n_20478,
       n_20479;
  wire n_20480, n_20481, n_20482, n_20483, n_20484, n_20485, n_20486,
       n_20487;
  wire n_20488, n_20489, n_20490, n_20491, n_20492, n_20493, n_20494,
       n_20495;
  wire n_20496, n_20497, n_20498, n_20499, n_20500, n_20501, n_20502,
       n_20503;
  wire n_20504, n_20505, n_20506, n_20507, n_20508, n_20509, n_20510,
       n_20511;
  wire n_20512, n_20513, n_20514, n_20515, n_20516, n_20517, n_20518,
       n_20519;
  wire n_20520, n_20521, n_20522, n_20523, n_20524, n_20525, n_20526,
       n_20527;
  wire n_20528, n_20529, n_20530, n_20531, n_20532, n_20533, n_20534,
       n_20535;
  wire n_20536, n_20537, n_20538, n_20539, n_20540, n_20541, n_20542,
       n_20543;
  wire n_20544, n_20545, n_20546, n_20547, n_20548, n_20549, n_20550,
       n_20551;
  wire n_20552, n_20553, n_20554, n_20555, n_20556, n_20557, n_20558,
       n_20559;
  wire n_20560, n_20561, n_20562, n_20563, n_20564, n_20565, n_20566,
       n_20567;
  wire n_20568, n_20569, n_20570, n_20571, n_20572, n_20573, n_20574,
       n_20575;
  wire n_20576, n_20577, n_20578, n_20579, n_20580, n_20581, n_20582,
       n_20583;
  wire n_20584, n_20585, n_20586, n_20587, n_20588, n_20589, n_20590,
       n_20591;
  wire n_20592, n_20593, n_20594, n_20595, n_20596, n_20597, n_20598,
       n_20599;
  wire n_20600, n_20601, n_20602, n_20603, n_20604, n_20605, n_20606,
       n_20607;
  wire n_20608, n_20609, n_20610, n_20611, n_20612, n_20613, n_20614,
       n_20615;
  wire n_20616, n_20617, n_20618, n_20619, n_20620, n_20621, n_20622,
       n_20623;
  wire n_20624, n_20625, n_20626, n_20627, n_20628, n_20629, n_20630,
       n_20631;
  wire n_20632, n_20633, n_20634, n_20635, n_20636, n_20637, n_20638,
       n_20639;
  wire n_20640, n_20641, n_20642, n_20643, n_20644, n_20645, n_20646,
       n_20647;
  wire n_20648, n_20649, n_20650, n_20651, n_20652, n_20653, n_20654,
       n_20655;
  wire n_20656, n_20657, n_20658, n_20659, n_20660, n_20661, n_20662,
       n_20663;
  wire n_20664, n_20665, n_20666, n_20667, n_20668, n_20669, n_20670,
       n_20671;
  wire n_20672, n_20673, n_20674, n_20675, n_20676, n_20677, n_20678,
       n_20679;
  wire n_20680, n_20681, n_20682, n_20683, n_20684, n_20685, n_20686,
       n_20687;
  wire n_20688, n_20689, n_20690, n_20691, n_20692, n_20693, n_20694,
       n_20695;
  wire n_20696, n_20697, n_20698, n_20699, n_20700, n_20701, n_20702,
       n_20703;
  wire n_20704, n_20705, n_20706, n_20707, n_20708, n_20709, n_20710,
       n_20711;
  wire n_20712, n_20713, n_20714, n_20715, n_20716, n_20717, n_20718,
       n_20719;
  wire n_20720, n_20721, n_20722, n_20723, n_20724, n_20725, n_20726,
       n_20727;
  wire n_20728, n_20729, n_20730, n_20731, n_20732, n_20733, n_20734,
       n_20735;
  wire n_20736, n_20737, n_20738, n_20739, n_20740, n_20741, n_20742,
       n_20743;
  wire n_20744, n_20745, n_20746, n_20747, n_20748, n_20749, n_20750,
       n_20751;
  wire n_20752, n_20753, n_20754, n_20755, n_20756, n_20757, n_20758,
       n_20759;
  wire n_20760, n_20761, n_20762, n_20763, n_20764, n_20765, n_20766,
       n_20767;
  wire n_20768, n_20769, n_20770, n_20771, n_20772, n_20773, n_20774,
       n_20775;
  wire n_20776, n_20777, n_20778, n_20779, n_20780, n_20781, n_20782,
       n_20783;
  wire n_20784, n_20785, n_20786, n_20787, n_20788, n_20789, n_20790,
       n_20791;
  wire n_20792, n_20793, n_20794, n_20795, n_20796, n_20797, n_20798,
       n_20799;
  wire n_20800, n_20801, n_20802, n_20803, n_20804, n_20805, n_20806,
       n_20807;
  wire n_20808, n_20809, n_20810, n_20811, n_20812, n_20813, n_20814,
       n_20815;
  wire n_20816, n_20817, n_20818, n_20819, n_20820, n_20821, n_20822,
       n_20823;
  wire n_20824, n_20825, n_20826, n_20827, n_20828, n_20829, n_20830,
       n_20831;
  wire n_20832, n_20833, n_20834, n_20835, n_20836, n_20837, n_20838,
       n_20839;
  wire n_20840, n_20841, n_20842, n_20843, n_20844, n_20845, n_20846,
       n_20847;
  wire n_20848, n_20849, n_20850, n_20851, n_20852, n_20853, n_20854,
       n_20855;
  wire n_20856, n_20857, n_20858, n_20859, n_20860, n_20861, n_20862,
       n_20863;
  wire n_20864, n_20865, n_20866, n_20867, n_20868, n_20869, n_20870,
       n_20871;
  wire n_20872, n_20873, n_20874, n_20875, n_20876, n_20877, n_20878,
       n_20879;
  wire n_20880, n_20881, n_20882, n_20883, n_20884, n_20885, n_20886,
       n_20887;
  wire n_20888, n_20889, n_20890, n_20891, n_20892, n_20893, n_20894,
       n_20895;
  wire n_20896, n_20897, n_20898, n_20899, n_20900, n_20901, n_20902,
       n_20903;
  wire n_20904, n_20905, n_20906, n_20907, n_20908, n_20909, n_20910,
       n_20911;
  wire n_20912, n_20913, n_20914, n_20915, n_20916, n_20917, n_20918,
       n_20919;
  wire n_20920, n_20921, n_20922, n_20923, n_20924, n_20925, n_20926,
       n_20927;
  wire n_20928, n_20929, n_20930, n_20931, n_20932, n_20933, n_20934,
       n_20935;
  wire n_20936, n_20937, n_20938, n_20939, n_20940, n_20941, n_20942,
       n_20943;
  wire n_20944, n_20945, n_20946, n_20947, n_20948, n_20949, n_20950,
       n_20951;
  wire n_20952, n_20953, n_20954, n_20955, n_20956, n_20961, n_20962,
       n_20963;
  wire n_20964, n_20965, n_20966, n_20967, n_20968, n_20969, n_20970,
       n_20971;
  wire n_20972, n_20973, n_20974, n_20975, n_20976, n_20977, n_20978,
       n_20979;
  wire n_20980, n_20981, n_20982, n_20983, n_20984, n_20985, n_20986,
       n_20987;
  wire n_20988, n_20989, n_20990, n_20991, n_20992, n_20993, n_20994,
       n_20995;
  wire n_20996, n_20997, n_20998, n_20999, n_21000, n_21001, n_21002,
       n_21003;
  wire n_21004, n_21005, n_21006, n_21007, n_21008, n_21009, n_21010,
       n_21011;
  wire n_21012, n_21013, n_21014, n_21015, n_21016, n_21017, n_21018,
       n_21019;
  wire n_21020, n_21021, n_21022, n_21023, n_21024, n_21025, n_21026,
       n_21027;
  wire n_21028, n_21029, n_21030, n_21031, n_21032, n_21033, n_21034,
       n_21035;
  wire n_21036, n_21037, n_21038, n_21039, n_21040, n_21041, n_21042,
       n_21043;
  wire n_21044, n_21045, n_21046, n_21047, n_21048, n_21049, n_21050,
       n_21051;
  wire n_21052, n_21053, n_21054, n_21055, n_21056, n_21057, n_21058,
       n_21059;
  wire n_21060, n_21061, n_21062, n_21063, n_21064, n_21065, n_21066,
       n_21067;
  wire n_21068, n_21069, n_21070, n_21071, n_21072, n_21073, n_21074,
       n_21075;
  wire n_21076, n_21077, n_21078, n_21079, n_21080, n_21081, n_21082,
       n_21083;
  wire n_21084, n_21085, n_21086, n_21087, n_21088, n_21089, n_21090,
       n_21091;
  wire n_21092, n_21093, n_21094, n_21095, n_21096, n_21097, n_21098,
       n_21099;
  wire n_21100, n_21101, n_21102, n_21103, n_21104, n_21105, n_21106,
       n_21107;
  wire n_21108, n_21109, n_21110, n_21111, n_21112, n_21113, n_21114,
       n_21115;
  wire n_21116, n_21117, n_21118, n_21119, n_21120, n_21121, n_21122,
       n_21123;
  wire n_21124, n_21125, n_21126, n_21127, n_21128, n_21129, n_21130,
       n_21131;
  wire n_21132, n_21133, n_21134, n_21135, n_21136, n_21137, n_21138,
       n_21139;
  wire n_21140, n_21141, n_21142, n_21143, n_21144, n_21145, n_21146,
       n_21147;
  wire n_21148, n_21149, n_21150, n_21151, n_21152, n_21153, n_21154,
       n_21155;
  wire n_21156, n_21157, n_21158, n_21159, n_21160, n_21161, n_21162,
       n_21163;
  wire n_21164, n_21165, n_21166, n_21167, n_21168, n_21169, n_21170,
       n_21171;
  wire n_21172, n_21173, n_21174, n_21175, n_21176, n_21177, n_21178,
       n_21179;
  wire n_21180, n_21181, n_21182, n_21183, n_21184, n_21185, n_21186,
       n_21187;
  wire n_21188, n_21189, n_21190, n_21191, n_21192, n_21193, n_21194,
       n_21195;
  wire n_21196, n_21197, n_21198, n_21199, n_21200, n_21201, n_21202,
       n_21203;
  wire n_21204, n_21205, n_21208, n_21209, n_21210, n_21211, n_21212,
       n_21213;
  wire n_21214, n_21215, n_21216, n_21217, n_21218, n_21219, n_21220,
       n_21221;
  wire n_21222, n_21223, n_21224, n_21225, n_21226, n_21227, n_21228,
       n_21229;
  wire n_21230, n_21231, n_21232, n_21233, n_21234, n_21235, n_21236,
       n_21237;
  wire n_21238, n_21239, n_21240, n_21241, n_21242, n_21243, n_21244,
       n_21245;
  wire n_21246, n_21247, n_21248, n_21249, n_21250, n_21251, n_21252,
       n_21253;
  wire n_21254, n_21255, n_21256, n_21257, n_21258, n_21259, n_21260,
       n_21261;
  wire n_21262, n_21263, n_21264, n_21265, n_21266, n_21267, n_21268,
       n_21269;
  wire n_21270, n_21271, n_21272, n_21273, n_21274, n_21275, n_21276,
       n_21277;
  wire n_21278, n_21279, n_21280, n_21281, n_21282, n_21283, n_21284,
       n_21285;
  wire n_21286, n_21287, n_21288, n_21289, n_21290, n_21291, n_21292,
       n_21293;
  wire n_21294, n_21295, n_21296, n_21297, n_21298, n_21299, n_21300,
       n_21301;
  wire n_21302, n_21303, n_21304, n_21305, n_21306, n_21307, n_21308,
       n_21309;
  wire n_21310, n_21311, n_21312, n_21313, n_21314, n_21315, n_21316,
       n_21317;
  wire n_21318, n_21319, n_21320, n_21321, n_21322, n_21323, n_21324,
       n_21325;
  wire n_21326, n_21327, n_21328, n_21329, n_21330, n_21331, n_21332,
       n_21333;
  wire n_21334, n_21335, n_21336, n_21337, n_21338, n_21339, n_21340,
       n_21341;
  wire n_21342, n_21343, n_21344, n_21345, n_21346, n_21347, n_21348,
       n_21349;
  wire n_21350, n_21351, n_21352, n_21353, n_21354, n_21355, n_21356,
       n_21357;
  wire n_21358, n_21359, n_21360, n_21361, n_21362, n_21363, n_21364,
       n_21365;
  wire n_21366, n_21367, n_21368, n_21369, n_21370, n_21371, n_21372,
       n_21373;
  wire n_21374, n_21375, n_21376, n_21377, n_21378, n_21379, n_21380,
       n_21381;
  wire n_21382, n_21383, n_21384, n_21385, n_21386, n_21387, n_21388,
       n_21389;
  wire n_21390, n_21391, n_21392, n_21393, n_21394, n_21395, n_21396,
       n_21397;
  wire n_21398, n_21399, n_21400, n_21401, n_21402, n_21403, n_21404,
       n_21405;
  wire n_21406, n_21407, n_21408, n_21409, n_21410, n_21411, n_21412,
       n_21413;
  wire n_21414, n_21415, n_21416, n_21417, n_21418, n_21419, n_21420,
       n_21421;
  wire n_21422, n_21423, n_21424, n_21425, n_21426, n_21427, n_21428,
       n_21429;
  wire n_21430, n_21431, n_21432, n_21433, n_21434, n_21435, n_21436,
       n_21437;
  wire n_21438, n_21439, n_21440, n_21441, n_21442, n_21443, n_21444,
       n_21445;
  wire n_21446, n_21447, n_21448, n_21449, n_21450, n_21451, n_21452,
       n_21453;
  wire n_21454, n_21455, n_21456, n_21457, n_21458, n_21459, n_21460,
       n_21461;
  wire n_21462, n_21463, n_21464, n_21465, n_21466, n_21467, n_21468,
       n_21469;
  wire n_21470, n_21471, n_21472, n_21473, n_21474, n_21475, n_21476,
       n_21477;
  wire n_21478, n_21479, n_21480, n_21481, n_21482, n_21483, n_21484,
       n_21485;
  wire n_21486, n_21487, n_21488, n_21489, n_21490, n_21491, n_21492,
       n_21493;
  wire n_21494, n_21495, n_21496, n_21497, n_21498, n_21499, n_21500,
       n_21501;
  wire n_21502, n_21503, n_21504, n_21505, n_21506, n_21507, n_21508,
       n_21509;
  wire n_21510, n_21511, n_21512, n_21513, n_21514, n_21515, n_21516,
       n_21517;
  wire n_21518, n_21519, n_21520, n_21521, n_21522, n_21523, n_21524,
       n_21525;
  wire n_21526, n_21527, n_21528, n_21529, n_21530, n_21531, n_21532,
       n_21533;
  wire n_21534, n_21535, n_21536, n_21537, n_21538, n_21539, n_21540,
       n_21541;
  wire n_21542, n_21543, n_21544, n_21545, n_21546, n_21547, n_21548,
       n_21549;
  wire n_21550, n_21551, n_21552, n_21553, n_21554, n_21555, n_21556,
       n_21557;
  wire n_21558, n_21559, n_21560, n_21561, n_21562, n_21563, n_21564,
       n_21565;
  wire n_21566, n_21567, n_21568, n_21569, n_21570, n_21571, n_21572,
       n_21573;
  wire n_21576, n_21577, n_21578, n_21579, n_21580, n_21581, n_21582,
       n_21583;
  wire n_21584, n_21585, n_21586, n_21587, n_21588, n_21589, n_21590,
       n_21591;
  wire n_21592, n_21593, n_21594, n_21595, n_21596, n_21597, n_21598,
       n_21599;
  wire n_21600, n_21601, n_21602, n_21603, n_21604, n_21605, n_21606,
       n_21607;
  wire n_21608, n_21609, n_21610, n_21611, n_21612, n_21613, n_21614,
       n_21615;
  wire n_21616, n_21617, n_21618, n_21619, n_21620, n_21621, n_21622,
       n_21623;
  wire n_21624, n_21625, n_21626, n_21627, n_21628, n_21629, n_21630,
       n_21631;
  wire n_21632, n_21633, n_21634, n_21635, n_21636, n_21637, n_21638,
       n_21639;
  wire n_21640, n_21641, n_21642, n_21643, n_21644, n_21645, n_21646,
       n_21647;
  wire n_21648, n_21649, n_21650, n_21651, n_21652, n_21653, n_21654,
       n_21655;
  wire n_21656, n_21657, n_21658, n_21659, n_21660, n_21661, n_21662,
       n_21663;
  wire n_21664, n_21665, n_21666, n_21667, n_21668, n_21669, n_21670,
       n_21671;
  wire n_21672, n_21673, n_21674, n_21675, n_21676, n_21677, n_21678,
       n_21679;
  wire n_21680, n_21681, n_21682, n_21683, n_21684, n_21685, n_21686,
       n_21687;
  wire n_21688, n_21689, n_21690, n_21691, n_21692, n_21693, n_21694,
       n_21695;
  wire n_21696, n_21697, n_21698, n_21699, n_21700, n_21701, n_21702,
       n_21703;
  wire n_21704, n_21705, n_21706, n_21707, n_21708, n_21709, n_21710,
       n_21711;
  wire n_21712, n_21713, n_21714, n_21715, n_21716, n_21717, n_21718,
       n_21719;
  wire n_21720, n_21721, n_21722, n_21723, n_21724, n_21725, n_21726,
       n_21727;
  wire n_21728, n_21729, n_21730, n_21731, n_21732, n_21733, n_21734,
       n_21735;
  wire n_21736, n_21737, n_21738, n_21739, n_21740, n_21741, n_21742,
       n_21743;
  wire n_21744, n_21745, n_21746, n_21747, n_21748, n_21749, n_21750,
       n_21751;
  wire n_21752, n_21753, n_21754, n_21755, n_21756, n_21757, n_21758,
       n_21759;
  wire n_21760, n_21761, n_21762, n_21763, n_21764, n_21765, n_21766,
       n_21767;
  wire n_21768, n_21769, n_21770, n_21771, n_21772, n_21773, n_21774,
       n_21775;
  wire n_21776, n_21777, n_21778, n_21779, n_21780, n_21781, n_21782,
       n_21783;
  wire n_21784, n_21785, n_21786, n_21787, n_21788, n_21789, n_21790,
       n_21791;
  wire n_21792, n_21793, n_21794, n_21795, n_21796, n_21797, n_21798,
       n_21799;
  wire n_21800, n_21801, n_21802, n_21803, n_21804, n_21805, n_21806,
       n_21807;
  wire n_21808, n_21809, n_21810, n_21811, n_21812, n_21813, n_21814,
       n_21815;
  wire n_21816, n_21817, n_21818, n_21819, n_21820, n_21821, n_21822,
       n_21823;
  wire n_21824, n_21825, n_21826, n_21827, n_21828, n_21829, n_21830,
       n_21831;
  wire n_21832, n_21833, n_21834, n_21835, n_21836, n_21837, n_21838,
       n_21839;
  wire n_21840, n_21841, n_21842, n_21843, n_21844, n_21845, n_21846,
       n_21847;
  wire n_21848, n_21849, n_21850, n_21851, n_21852, n_21853, n_21854,
       n_21855;
  wire n_21856, n_21857, n_21858, n_21859, n_21860, n_21861, n_21862,
       n_21863;
  wire n_21864, n_21865, n_21866, n_21867, n_21868, n_21869, n_21870,
       n_21871;
  wire n_21872, n_21873, n_21874, n_21875, n_21876, n_21877, n_21878,
       n_21879;
  wire n_21880, n_21881, n_21882, n_21883, n_21884, n_21885, n_21886,
       n_21887;
  wire n_21888, n_21889, n_21890, n_21891, n_21892, n_21893, n_21894,
       n_21895;
  wire n_21896, n_21897, n_21898, n_21899, n_21900, n_21901, n_21902,
       n_21903;
  wire n_21904, n_21905, n_21906, n_21907, n_21908, n_21909, n_21910,
       n_21911;
  wire n_21912, n_21913, n_21914, n_21915, n_21916, n_21917, n_21918,
       n_21919;
  wire n_21920, n_21921, n_21922, n_21923, n_21924, n_21925, n_21926,
       n_21927;
  wire n_21928, n_21929, n_21930, n_21931, n_21932, n_21933, n_21934,
       n_21935;
  wire n_21936, n_21937, n_21938, n_21939, n_21940, n_21941, n_21942,
       n_21943;
  wire n_21946, n_21947, n_21948, n_21949, n_21950, n_21951, n_21952,
       n_21953;
  wire n_21954, n_21955, n_21956, n_21957, n_21958, n_21959, n_21960,
       n_21961;
  wire n_21962, n_21963, n_21964, n_21965, n_21966, n_21967, n_21968,
       n_21969;
  wire n_21970, n_21971, n_21972, n_21973, n_21974, n_21975, n_21976,
       n_21977;
  wire n_21978, n_21979, n_21980, n_21981, n_21982, n_21983, n_21984,
       n_21985;
  wire n_21986, n_21987, n_21988, n_21989, n_21990, n_21991, n_21992,
       n_21993;
  wire n_21994, n_21995, n_21996, n_21997, n_21998, n_21999, n_22000,
       n_22001;
  wire n_22002, n_22003, n_22004, n_22005, n_22006, n_22007, n_22008,
       n_22009;
  wire n_22010, n_22011, n_22012, n_22013, n_22014, n_22015, n_22016,
       n_22017;
  wire n_22018, n_22019, n_22020, n_22021, n_22022, n_22023, n_22024,
       n_22025;
  wire n_22026, n_22027, n_22028, n_22029, n_22030, n_22031, n_22032,
       n_22033;
  wire n_22034, n_22035, n_22036, n_22037, n_22038, n_22039, n_22040,
       n_22041;
  wire n_22042, n_22043, n_22044, n_22045, n_22046, n_22047, n_22048,
       n_22049;
  wire n_22050, n_22051, n_22052, n_22053, n_22054, n_22055, n_22056,
       n_22057;
  wire n_22058, n_22059, n_22060, n_22061, n_22062, n_22063, n_22064,
       n_22065;
  wire n_22066, n_22067, n_22068, n_22069, n_22070, n_22071, n_22072,
       n_22073;
  wire n_22074, n_22075, n_22076, n_22077, n_22078, n_22079, n_22080,
       n_22081;
  wire n_22082, n_22083, n_22084, n_22085, n_22086, n_22087, n_22088,
       n_22089;
  wire n_22090, n_22091, n_22092, n_22093, n_22094, n_22095, n_22096,
       n_22097;
  wire n_22098, n_22099, n_22100, n_22101, n_22102, n_22103, n_22104,
       n_22105;
  wire n_22106, n_22107, n_22108, n_22109, n_22110, n_22111, n_22112,
       n_22113;
  wire n_22114, n_22115, n_22116, n_22117, n_22118, n_22119, n_22120,
       n_22121;
  wire n_22122, n_22123, n_22124, n_22125, n_22126, n_22127, n_22128,
       n_22129;
  wire n_22130, n_22131, n_22132, n_22133, n_22134, n_22135, n_22136,
       n_22137;
  wire n_22138, n_22139, n_22140, n_22141, n_22142, n_22143, n_22144,
       n_22145;
  wire n_22146, n_22147, n_22148, n_22149, n_22150, n_22151, n_22152,
       n_22153;
  wire n_22154, n_22155, n_22156, n_22157, n_22158, n_22159, n_22160,
       n_22161;
  wire n_22162, n_22163, n_22164, n_22165, n_22166, n_22167, n_22168,
       n_22169;
  wire n_22170, n_22171, n_22172, n_22173, n_22174, n_22175, n_22176,
       n_22177;
  wire n_22178, n_22179, n_22180, n_22181, n_22182, n_22183, n_22184,
       n_22185;
  wire n_22186, n_22187, n_22188, n_22189, n_22190, n_22191, n_22192,
       n_22193;
  wire n_22194, n_22195, n_22196, n_22197, n_22198, n_22199, n_22200,
       n_22201;
  wire n_22202, n_22203, n_22204, n_22205, n_22206, n_22207, n_22208,
       n_22209;
  wire n_22210, n_22211, n_22212, n_22213, n_22214, n_22215, n_22216,
       n_22217;
  wire n_22218, n_22219, n_22220, n_22221, n_22222, n_22223, n_22224,
       n_22225;
  wire n_22226, n_22227, n_22228, n_22229, n_22230, n_22231, n_22232,
       n_22233;
  wire n_22234, n_22235, n_22236, n_22237, n_22238, n_22239, n_22240,
       n_22241;
  wire n_22242, n_22243, n_22244, n_22245, n_22246, n_22247, n_22248,
       n_22249;
  wire n_22250, n_22251, n_22252, n_22253, n_22254, n_22255, n_22256,
       n_22257;
  wire n_22258, n_22259, n_22260, n_22261, n_22262, n_22263, n_22264,
       n_22265;
  wire n_22266, n_22267, n_22268, n_22269, n_22270, n_22271, n_22272,
       n_22273;
  wire n_22274, n_22275, n_22276, n_22277, n_22278, n_22279, n_22280,
       n_22281;
  wire n_22282, n_22283, n_22284, n_22285, n_22286, n_22287, n_22288,
       n_22289;
  wire n_22290, n_22291, n_22292, n_22293, n_22294, n_22295, n_22296,
       n_22297;
  wire n_22298, n_22299, n_22300, n_22301, n_22302, n_22303, n_22304,
       n_22305;
  wire n_22306, n_22307, n_22308, n_22309, n_22310, n_22311, n_22312,
       n_22313;
  wire n_22314, n_22315, n_22316, n_22317, n_22318, n_22319, n_22320,
       n_22321;
  wire n_22322, n_22323, n_22324, n_22325, n_22326, n_22327, n_22328,
       n_22329;
  wire n_22330, n_22331, n_22332, n_22333, n_22334, n_22335, n_22336,
       n_22337;
  wire n_22338, n_22339, n_22340, n_22341, n_22342, n_22343, n_22345,
       n_22346;
  wire n_22347, n_22348, n_22349, n_22350, n_22351, n_22352, n_22353,
       n_22354;
  wire n_22355, n_22356, n_22357, n_22358, n_22359, n_22360, n_22361,
       n_22362;
  wire n_22363, n_22364, n_22365, n_22366, n_22367, n_22368, n_22369,
       n_22370;
  wire n_22371, n_22372, n_22373, n_22374, n_22375, n_22376, n_22377,
       n_22378;
  wire n_22379, n_22380, n_22381, n_22382, n_22383, n_22384, n_22385,
       n_22386;
  wire n_22387, n_22388, n_22389, n_22390, n_22391, n_22392, n_22393,
       n_22394;
  wire n_22395, n_22396, n_22397, n_22398, n_22399, n_22400, n_22401,
       n_22402;
  wire n_22403, n_22404, n_22405, n_22406, n_22407, n_22408, n_22409,
       n_22410;
  wire n_22411, n_22412, n_22413, n_22414, n_22415, n_22416, n_22417,
       n_22418;
  wire n_22419, n_22420, n_22421, n_22422, n_22423, n_22424, n_22425,
       n_22426;
  wire n_22427, n_22428, n_22429, n_22430, n_22431, n_22432, n_22433,
       n_22434;
  wire n_22435, n_22436, n_22437, n_22438, n_22439, n_22440, n_22441,
       n_22442;
  wire n_22443, n_22444, n_22445, n_22446, n_22447, n_22448, n_22449,
       n_22450;
  wire n_22451, n_22452, n_22453, n_22454, n_22455, n_22456, n_22457,
       n_22458;
  wire n_22459, n_22460, n_22461, n_22462, n_22463, n_22464, n_22465,
       n_22466;
  wire n_22467, n_22468, n_22469, n_22470, n_22471, n_22472, n_22473,
       n_22474;
  wire n_22475, n_22476, n_22477, n_22478, n_22479, n_22480, n_22481,
       n_22482;
  wire n_22483, n_22484, n_22485, n_22486, n_22487, n_22488, n_22489,
       n_22490;
  wire n_22491, n_22492, n_22493, n_22494, n_22495, n_22496, n_22497,
       n_22498;
  wire n_22499, n_22500, n_22501, n_22502, n_22503, n_22504, n_22505,
       n_22506;
  wire n_22507, n_22508, n_22509, n_22510, n_22511, n_22512, n_22513,
       n_22514;
  wire n_22515, n_22516, n_22517, n_22518, n_22519, n_22520, n_22521,
       n_22522;
  wire n_22523, n_22524, n_22525, n_22526, n_22527, n_22528, n_22529,
       n_22530;
  wire n_22531, n_22532, n_22533, n_22534, n_22535, n_22536, n_22537,
       n_22538;
  wire n_22539, n_22540, n_22541, n_22542, n_22543, n_22544, n_22545,
       n_22546;
  wire n_22547, n_22548, n_22549, n_22550, n_22551, n_22552, n_22553,
       n_22554;
  wire n_22555, n_22556, n_22557, n_22558, n_22559, n_22560, n_22561,
       n_22562;
  wire n_22563, n_22564, n_22565, n_22566, n_22567, n_22568, n_22569,
       n_22570;
  wire n_22571, n_22572, n_22573, n_22574, n_22575, n_22576, n_22577,
       n_22578;
  wire n_22579, n_22580, n_22581, n_22582, n_22583, n_22584, n_22585,
       n_22586;
  wire n_22587, n_22588, n_22589, n_22590, n_22591, n_22592, n_22593,
       n_22594;
  wire n_22595, n_22596, n_22597, n_22598, n_22599, n_22600, n_22601,
       n_22602;
  wire n_22603, n_22604, n_22605, n_22606, n_22607, n_22608, n_22609,
       n_22610;
  wire n_22611, n_22612, n_22613, n_22614, n_22615, n_22616, n_22617,
       n_22618;
  wire n_22619, n_22620, n_22621, n_22622, n_22623, n_22624, n_22625,
       n_22626;
  wire n_22627, n_22628, n_22629, n_22630, n_22631, n_22632, n_22633,
       n_22634;
  wire n_22635, n_22636, n_22637, n_22638, n_22639, n_22640, n_22641,
       n_22642;
  wire n_22643, n_22644, n_22645, n_22646, n_22647, n_22648, n_22649,
       n_22650;
  wire n_22651, n_22652, n_22653, n_22654, n_22655, n_22656, n_22657,
       n_22658;
  wire n_22659, n_22660, n_22661, n_22662, n_22663, n_22664, n_22665,
       n_22666;
  wire n_22667, n_22668, n_22669, n_22670, n_22671, n_22672, n_22673,
       n_22674;
  wire n_22675, n_22676, n_22677, n_22678, n_22679, n_22680, n_22681,
       n_22682;
  wire n_22683, n_22684, n_22685, n_22686, n_22687, n_22688, n_22689,
       n_22690;
  wire n_22691, n_22692, n_22693, n_22694, n_22695, n_22696, n_22697,
       n_22698;
  wire n_22699, n_22700, n_22701, n_22702, n_22703, n_22704, n_22705,
       n_22706;
  wire n_22707, n_22708, n_22709, n_22710, n_22711, n_22712, n_22713,
       n_22714;
  wire n_22715, n_22716, n_22717, n_22718, n_22719, n_22720, n_22721,
       n_22722;
  wire n_22723, n_22724, n_22725, n_22726, n_22727, n_22728, n_22729,
       n_22730;
  wire n_22731, n_22732, n_22733, n_22734, n_22735, n_22736, n_22737,
       n_22738;
  wire n_22739, n_22740, n_22741, n_22742, n_22743, n_22744, n_22745,
       n_22746;
  wire n_22747, n_22748, n_22749, n_22750, n_22751, n_22752, n_22753,
       n_22754;
  wire n_22755, n_22756, n_22757, n_22758, n_22759, n_22760, n_22761,
       n_22762;
  wire n_22763, n_22764, n_22765, n_22766, n_22767, n_22768, n_22769,
       n_22770;
  wire n_22771, n_22772, n_22773, n_22774, n_22775, n_22776, n_22777,
       n_22778;
  wire n_22779, n_22780, n_22781, n_22782, n_22783, n_22784, n_22785,
       n_22786;
  wire n_22787, n_22788, n_22789, n_22790, n_22791, n_22792, n_22793,
       n_22794;
  wire n_22795, n_22796, n_22797, n_22798, n_22799, n_22800, n_22801,
       n_22802;
  wire n_22803, n_22804, n_22805, n_22806, n_22810, n_22811, n_22812,
       n_22813;
  wire n_22814, n_22815, n_22816, n_22817, n_22818, n_22819, n_22820,
       n_22821;
  wire n_22822, n_22823, n_22824, n_22825, n_22826, n_22827, n_22828,
       n_22829;
  wire n_22830, n_22831, n_22832, n_22833, n_22834, n_22835, n_22836,
       n_22837;
  wire n_22838, n_22839, n_22840, n_22841, n_22842, n_22843, n_22844,
       n_22845;
  wire n_22846, n_22847, n_22848, n_22849, n_22850, n_22851, n_22852,
       n_22853;
  wire n_22854, n_22855, n_22856, n_22857, n_22858, n_22859, n_22860,
       n_22861;
  wire n_22862, n_22863, n_22864, n_22865, n_22866, n_22867, n_22868,
       n_22869;
  wire n_22870, n_22871, n_22872, n_22873, n_22874, n_22875, n_22876,
       n_22877;
  wire n_22878, n_22879, n_22880, n_22881, n_22882, n_22883, n_22884,
       n_22885;
  wire n_22886, n_22887, n_22888, n_22889, n_22890, n_22891, n_22892,
       n_22893;
  wire n_22894, n_22895, n_22896, n_22897, n_22898, n_22899, n_22900,
       n_22901;
  wire n_22902, n_22903, n_22904, n_22905, n_22906, n_22907, n_22908,
       n_22909;
  wire n_22910, n_22911, n_22912, n_22913, n_22914, n_22915, n_22916,
       n_22917;
  wire n_22918, n_22919, n_22920, n_22921, n_22922, n_22923, n_22924,
       n_22925;
  wire n_22926, n_22927, n_22928, n_22929, n_22930, n_22931, n_22932,
       n_22933;
  wire n_22934, n_22935, n_22936, n_22937, n_22938, n_22939, n_22940,
       n_22941;
  wire n_22942, n_22943, n_22944, n_22945, n_22946, n_22947, n_22948,
       n_22949;
  wire n_22950, n_22951, n_22952, n_22953, n_22954, n_22955, n_22956,
       n_22957;
  wire n_22958, n_22959, n_22960, n_22961, n_22962, n_22963, n_22964,
       n_22965;
  wire n_22966, n_22967, n_22968, n_22969, n_22970, n_22971, n_22972,
       n_22973;
  wire n_22974, n_22975, n_22976, n_22977, n_22978, n_22979, n_22980,
       n_22981;
  wire n_22982, n_22983, n_22984, n_22985, n_22986, n_22987, n_22988,
       n_22989;
  wire n_22990, n_22991, n_22992, n_22993, n_22994, n_22995, n_22996,
       n_22997;
  wire n_22998, n_22999, n_23000, n_23001, n_23002, n_23003, n_23004,
       n_23005;
  wire n_23006, n_23007, n_23008, n_23009, n_23010, n_23011, n_23012,
       n_23013;
  wire n_23014, n_23015, n_23016, n_23017, n_23018, n_23019, n_23020,
       n_23021;
  wire n_23022, n_23023, n_23024, n_23025, n_23026, n_23027, n_23028,
       n_23029;
  wire n_23030, n_23031, n_23032, n_23033, n_23034, n_23035, n_23036,
       n_23037;
  wire n_23038, n_23039, n_23040, n_23041, n_23042, n_23043, n_23044,
       n_23045;
  wire n_23046, n_23047, n_23048, n_23049, n_23050, n_23051, n_23052,
       n_23053;
  wire n_23054, n_23055, n_23056, n_23057, n_23058, n_23059, n_23060,
       n_23061;
  wire n_23062, n_23063, n_23064, n_23065, n_23066, n_23067, n_23068,
       n_23069;
  wire n_23070, n_23071, n_23072, n_23073, n_23074, n_23075, n_23076,
       n_23077;
  wire n_23078, n_23079, n_23080, n_23081, n_23082, n_23083, n_23084,
       n_23085;
  wire n_23086, n_23087, n_23088, n_23089, n_23090, n_23091, n_23092,
       n_23093;
  wire n_23094, n_23095, n_23096, n_23097, n_23098, n_23099, n_23100,
       n_23101;
  wire n_23102, n_23103, n_23104, n_23105, n_23106, n_23107, n_23108,
       n_23109;
  wire n_23110, n_23111, n_23112, n_23113, n_23114, n_23115, n_23116,
       n_23117;
  wire n_23118, n_23119, n_23120, n_23121, n_23122, n_23123, n_23124,
       n_23125;
  wire n_23126, n_23127, n_23128, n_23129, n_23130, n_23131, n_23132,
       n_23133;
  wire n_23134, n_23135, n_23136, n_23137, n_23138, n_23139, n_23140,
       n_23141;
  wire n_23142, n_23143, n_23144, n_23145, n_23146, n_23147, n_23148,
       n_23149;
  wire n_23150, n_23151, n_23152, n_23153, n_23154, n_23155, n_23156,
       n_23157;
  wire n_23158, n_23159, n_23160, n_23161, n_23162, n_23163, n_23164,
       n_23165;
  wire n_23166, n_23167, n_23168, n_23169, n_23170, n_23171, n_23172,
       n_23173;
  wire n_23174, n_23175, n_23176, n_23177, n_23178, n_23179, n_23180,
       n_23181;
  wire n_23182, n_23183, n_23184, n_23188, n_23189, n_23190, n_23191,
       n_23192;
  wire n_23193, n_23194, n_23195, n_23196, n_23197, n_23198, n_23199,
       n_23200;
  wire n_23201, n_23202, n_23203, n_23204, n_23205, n_23206, n_23207,
       n_23208;
  wire n_23209, n_23210, n_23211, n_23212, n_23213, n_23214, n_23215,
       n_23216;
  wire n_23217, n_23218, n_23219, n_23220, n_23221, n_23222, n_23223,
       n_23224;
  wire n_23225, n_23226, n_23227, n_23228, n_23229, n_23230, n_23231,
       n_23232;
  wire n_23233, n_23234, n_23235, n_23236, n_23237, n_23238, n_23239,
       n_23240;
  wire n_23241, n_23242, n_23243, n_23244, n_23245, n_23246, n_23247,
       n_23248;
  wire n_23249, n_23250, n_23251, n_23252, n_23253, n_23254, n_23255,
       n_23256;
  wire n_23257, n_23258, n_23259, n_23260, n_23261, n_23262, n_23263,
       n_23264;
  wire n_23265, n_23266, n_23267, n_23268, n_23269, n_23270, n_23271,
       n_23272;
  wire n_23273, n_23274, n_23275, n_23276, n_23277, n_23278, n_23279,
       n_23280;
  wire n_23281, n_23282, n_23283, n_23284, n_23285, n_23286, n_23287,
       n_23288;
  wire n_23289, n_23290, n_23291, n_23292, n_23293, n_23294, n_23295,
       n_23296;
  wire n_23297, n_23298, n_23299, n_23300, n_23301, n_23302, n_23303,
       n_23304;
  wire n_23305, n_23306, n_23307, n_23308, n_23309, n_23310, n_23311,
       n_23312;
  wire n_23313, n_23314, n_23315, n_23316, n_23317, n_23318, n_23319,
       n_23320;
  wire n_23321, n_23322, n_23323, n_23324, n_23325, n_23326, n_23327,
       n_23328;
  wire n_23329, n_23330, n_23331, n_23332, n_23333, n_23334, n_23335,
       n_23336;
  wire n_23337, n_23338, n_23339, n_23340, n_23341, n_23342, n_23343,
       n_23344;
  wire n_23345, n_23346, n_23347, n_23348, n_23349, n_23350, n_23351,
       n_23352;
  wire n_23353, n_23354, n_23355, n_23356, n_23357, n_23358, n_23359,
       n_23360;
  wire n_23361, n_23362, n_23363, n_23364, n_23365, n_23366, n_23367,
       n_23368;
  wire n_23369, n_23370, n_23371, n_23372, n_23373, n_23374, n_23375,
       n_23376;
  wire n_23377, n_23378, n_23379, n_23380, n_23381, n_23382, n_23383,
       n_23384;
  wire n_23385, n_23386, n_23387, n_23388, n_23389, n_23390, n_23391,
       n_23392;
  wire n_23393, n_23394, n_23395, n_23396, n_23397, n_23398, n_23399,
       n_23400;
  wire n_23401, n_23402, n_23403, n_23404, n_23405, n_23406, n_23407,
       n_23408;
  wire n_23409, n_23410, n_23411, n_23412, n_23413, n_23414, n_23415,
       n_23416;
  wire n_23417, n_23418, n_23419, n_23420, n_23421, n_23422, n_23423,
       n_23424;
  wire n_23425, n_23426, n_23427, n_23428, n_23429, n_23430, n_23431,
       n_23432;
  wire n_23433, n_23434, n_23435, n_23436, n_23437, n_23438, n_23439,
       n_23440;
  wire n_23441, n_23442, n_23443, n_23444, n_23445, n_23446, n_23447,
       n_23448;
  wire n_23449, n_23450, n_23451, n_23452, n_23453, n_23454, n_23455,
       n_23456;
  wire n_23457, n_23458, n_23459, n_23460, n_23461, n_23462, n_23463,
       n_23464;
  wire n_23465, n_23466, n_23467, n_23468, n_23469, n_23470, n_23471,
       n_23472;
  wire n_23473, n_23474, n_23475, n_23476, n_23477, n_23478, n_23479,
       n_23480;
  wire n_23481, n_23482, n_23483, n_23484, n_23485, n_23486, n_23487,
       n_23488;
  wire n_23489, n_23490, n_23491, n_23492, n_23493, n_23494, n_23495,
       n_23496;
  wire n_23497, n_23498, n_23499, n_23500, n_23501, n_23502, n_23503,
       n_23504;
  wire n_23505, n_23506, n_23507, n_23508, n_23509, n_23510, n_23511,
       n_23512;
  wire n_23513, n_23514, n_23515, n_23516, n_23517, n_23518, n_23519,
       n_23520;
  wire n_23521, n_23522, n_23523, n_23524, n_23525, n_23526, n_23527,
       n_23528;
  wire n_23529, n_23530, n_23531, n_23532, n_23533, n_23534, n_23535,
       n_23536;
  wire n_23537, n_23538, n_23539, n_23540, n_23541, n_23542, n_23543,
       n_23544;
  wire n_23545, n_23546, n_23547, n_23548, n_23549, n_23550, n_23551,
       n_23552;
  wire n_23553, n_23554, n_23555, n_23556, n_23557, n_23558, n_23559,
       n_23560;
  wire n_23561, n_23562, n_23566, n_23567, n_23568, n_23569, n_23570,
       n_23571;
  wire n_23572, n_23573, n_23574, n_23575, n_23576, n_23577, n_23578,
       n_23579;
  wire n_23580, n_23581, n_23582, n_23583, n_23584, n_23585, n_23586,
       n_23587;
  wire n_23588, n_23589, n_23590, n_23591, n_23592, n_23593, n_23594,
       n_23595;
  wire n_23596, n_23597, n_23598, n_23599, n_23600, n_23601, n_23602,
       n_23603;
  wire n_23604, n_23605, n_23606, n_23607, n_23608, n_23609, n_23610,
       n_23611;
  wire n_23612, n_23613, n_23614, n_23615, n_23616, n_23617, n_23618,
       n_23619;
  wire n_23620, n_23621, n_23622, n_23623, n_23624, n_23625, n_23626,
       n_23627;
  wire n_23628, n_23629, n_23630, n_23631, n_23632, n_23633, n_23634,
       n_23635;
  wire n_23636, n_23637, n_23638, n_23639, n_23640, n_23641, n_23642,
       n_23643;
  wire n_23644, n_23645, n_23646, n_23647, n_23648, n_23649, n_23650,
       n_23651;
  wire n_23652, n_23653, n_23654, n_23655, n_23656, n_23657, n_23658,
       n_23659;
  wire n_23660, n_23661, n_23662, n_23663, n_23664, n_23665, n_23666,
       n_23667;
  wire n_23668, n_23669, n_23670, n_23671, n_23672, n_23673, n_23674,
       n_23675;
  wire n_23676, n_23677, n_23678, n_23679, n_23680, n_23681, n_23682,
       n_23683;
  wire n_23684, n_23685, n_23686, n_23687, n_23688, n_23689, n_23690,
       n_23691;
  wire n_23692, n_23693, n_23694, n_23695, n_23696, n_23697, n_23698,
       n_23699;
  wire n_23700, n_23701, n_23702, n_23703, n_23704, n_23705, n_23706,
       n_23707;
  wire n_23708, n_23709, n_23710, n_23711, n_23712, n_23713, n_23714,
       n_23715;
  wire n_23716, n_23717, n_23718, n_23719, n_23720, n_23721, n_23722,
       n_23723;
  wire n_23724, n_23725, n_23726, n_23727, n_23728, n_23729, n_23730,
       n_23731;
  wire n_23732, n_23733, n_23734, n_23735, n_23736, n_23737, n_23738,
       n_23739;
  wire n_23740, n_23741, n_23742, n_23743, n_23744, n_23745, n_23746,
       n_23747;
  wire n_23748, n_23749, n_23750, n_23751, n_23752, n_23753, n_23754,
       n_23755;
  wire n_23756, n_23757, n_23758, n_23759, n_23760, n_23761, n_23762,
       n_23763;
  wire n_23764, n_23765, n_23766, n_23767, n_23768, n_23769, n_23770,
       n_23771;
  wire n_23772, n_23773, n_23774, n_23775, n_23776, n_23777, n_23778,
       n_23779;
  wire n_23780, n_23781, n_23782, n_23783, n_23784, n_23785, n_23786,
       n_23787;
  wire n_23788, n_23789, n_23790, n_23791, n_23792, n_23793, n_23794,
       n_23795;
  wire n_23796, n_23797, n_23798, n_23799, n_23800, n_23801, n_23802,
       n_23803;
  wire n_23804, n_23805, n_23806, n_23807, n_23808, n_23809, n_23810,
       n_23811;
  wire n_23812, n_23813, n_23814, n_23815, n_23816, n_23817, n_23818,
       n_23819;
  wire n_23820, n_23821, n_23822, n_23823, n_23824, n_23825, n_23826,
       n_23827;
  wire n_23828, n_23829, n_23830, n_23831, n_23832, n_23833, n_23834,
       n_23835;
  wire n_23836, n_23837, n_23838, n_23839, n_23840, n_23841, n_23842,
       n_23843;
  wire n_23844, n_23845, n_23846, n_23847, n_23848, n_23849, n_23850,
       n_23851;
  wire n_23852, n_23853, n_23854, n_23855, n_23856, n_23857, n_23858,
       n_23859;
  wire n_23860, n_23861, n_23862, n_23863, n_23864, n_23865, n_23866,
       n_23867;
  wire n_23868, n_23869, n_23870, n_23871, n_23872, n_23873, n_23874,
       n_23875;
  wire n_23876, n_23877, n_23878, n_23879, n_23880, n_23881, n_23882,
       n_23883;
  wire n_23884, n_23885, n_23886, n_23887, n_23888, n_23889, n_23890,
       n_23891;
  wire n_23892, n_23893, n_23894, n_23895, n_23896, n_23897, n_23898,
       n_23899;
  wire n_23900, n_23901, n_23902, n_23903, n_23904, n_23905, n_23906,
       n_23907;
  wire n_23908, n_23909, n_23910, n_23911, n_23912, n_23913, n_23914,
       n_23915;
  wire n_23916, n_23917, n_23918, n_23919, n_23920, n_23921, n_23922,
       n_23923;
  wire n_23924, n_23925, n_23926, n_23927, n_23928, n_23929, n_23930,
       n_23931;
  wire n_23932, n_23933, n_23934, n_23935, n_23936, n_23937, n_23938,
       n_23939;
  wire n_23940, n_23941, n_23942, n_23943, n_23944, n_23945, n_23946,
       n_23947;
  wire n_23948, n_23949, n_23950, n_23951, n_23952, n_23953, n_23954,
       n_23955;
  wire n_23956, n_23957, n_23958, n_23959, n_23960, n_23961, n_23962,
       n_23963;
  wire n_23964, n_23965, n_23966, n_23967, n_23968, n_23969, n_23970,
       n_23971;
  wire n_23972, n_23973, n_23974, n_23975, n_23976, n_23977, n_23978,
       n_23979;
  wire n_23980, n_23981, n_23982, n_23983, n_23984, n_23985, n_23986,
       n_23987;
  wire n_23988, n_23989, n_23990, n_23991, n_23992, n_23993, n_23994,
       n_23995;
  wire n_23996, n_23997, n_23998, n_23999, n_24000, n_24001, n_24002,
       n_24003;
  wire n_24004, n_24005, n_24006, n_24007, n_24008, n_24009, n_24010,
       n_24011;
  wire n_24012, n_24013, n_24014, n_24015, n_24016, n_24017, n_24018,
       n_24019;
  wire n_24020, n_24021, n_24022, n_24023, n_24024, n_24025, n_24026,
       n_24027;
  wire n_24028, n_24029, n_24030, n_24031, n_24032, n_24033, n_24034,
       n_24035;
  wire n_24036, n_24037, n_24038, n_24039, n_24040, n_24041, n_24042,
       n_24043;
  wire n_24044, n_24045, n_24046, n_24047, n_24048, n_24049, n_24050,
       n_24051;
  wire n_24052, n_24053, n_24054, n_24055, n_24056, n_24057, n_24058,
       n_24059;
  wire n_24060, n_24061, n_24062, n_24063, n_24064, n_24065, n_24066,
       n_24067;
  wire n_24068, n_24069, n_24070, n_24071, n_24072, n_24073, n_24074,
       n_24075;
  wire n_24076, n_24077, n_24078, n_24079, n_24080, n_24081, n_24082,
       n_24083;
  wire n_24084, n_24085, n_24086, n_24087, n_24088, n_24089, n_24090,
       n_24091;
  wire n_24092, n_24093, n_24094, n_24095, n_24096, n_24097, n_24098,
       n_24099;
  wire n_24100, n_24101, n_24102, n_24103, n_24104, n_24105, n_24106,
       n_24107;
  wire n_24108, n_24109, n_24110, n_24111, n_24112, n_24113, n_24114,
       n_24115;
  wire n_24116, n_24117, n_24118, n_24119, n_24120, n_24121, n_24122,
       n_24123;
  wire n_24124, n_24125, n_24126, n_24127, n_24128, n_24129, n_24130,
       n_24131;
  wire n_24132, n_24133, n_24134, n_24135, n_24136, n_24137, n_24138,
       n_24139;
  wire n_24140, n_24141, n_24142, n_24143, n_24144, n_24145, n_24146,
       n_24147;
  wire n_24148, n_24149, n_24150, n_24151, n_24152, n_24153, n_24154,
       n_24155;
  wire n_24156, n_24157, n_24158, n_24159, n_24160, n_24161, n_24162,
       n_24163;
  wire n_24164, n_24165, n_24166, n_24167, n_24168, n_24169, n_24170,
       n_24171;
  wire n_24172, n_24173, n_24174, n_24175, n_24176, n_24177, n_24178,
       n_24179;
  wire n_24180, n_24181, n_24182, n_24183, n_24184, n_24185, n_24186,
       n_24187;
  wire n_24188, n_24189, n_24190, n_24191, n_24192, n_24193, n_24194,
       n_24195;
  wire n_24196, n_24197, n_24198, n_24199, n_24200, n_24201, n_24202,
       n_24203;
  wire n_24204, n_24205, n_24206, n_24207, n_24208, n_24209, n_24210,
       n_24211;
  wire n_24212, n_24213, n_24214, n_24215, n_24216, n_24217, n_24218,
       n_24219;
  wire n_24220, n_24221, n_24222, n_24223, n_24224, n_24225, n_24226,
       n_24227;
  wire n_24228, n_24229, n_24230, n_24231, n_24232, n_24233, n_24234,
       n_24235;
  wire n_24236, n_24237, n_24238, n_24239, n_24240, n_24241, n_24242,
       n_24243;
  wire n_24244, n_24245, n_24246, n_24247, n_24248, n_24249, n_24250,
       n_24251;
  wire n_24252, n_24253, n_24254, n_24255, n_24256, n_24257, n_24258,
       n_24259;
  wire n_24260, n_24261, n_24262, n_24263, n_24264, n_24265, n_24266,
       n_24267;
  wire n_24268, n_24269, n_24270, n_24271, n_24272, n_24273, n_24274,
       n_24275;
  wire n_24276, n_24277, n_24278, n_24279, n_24280, n_24281, n_24282,
       n_24283;
  wire n_24284, n_24285, n_24286, n_24287, n_24288, n_24289, n_24290,
       n_24291;
  wire n_24292, n_24293, n_24294, n_24295, n_24296, n_24297, n_24298,
       n_24299;
  wire n_24300, n_24301, n_24302, n_24303, n_24304, n_24305, n_24306,
       n_24307;
  wire n_24308, n_24309, n_24310, n_24311, n_24312, n_24313, n_24314,
       n_24315;
  wire n_24316, n_24317, n_24318, n_24319, n_24320, n_24321, n_24322,
       n_24323;
  wire n_24324, n_24325, n_24326, n_24327, n_24328, n_24329, n_24330,
       n_24331;
  wire n_24332, n_24333, n_24334, n_24335, n_24336, n_24337, n_24338,
       n_24339;
  wire n_24340, n_24341, n_24342, n_24343, n_24344, n_24345, n_24346,
       n_24347;
  wire n_24348, n_24349, n_24350, n_24351, n_24352, n_24353, n_24354,
       n_24355;
  wire n_24356, n_24357, n_24358, n_24359, n_24360, n_24361, n_24362,
       n_24363;
  wire n_24364, n_24365, n_24366, n_24367, n_24368, n_24369, n_24370,
       n_24371;
  wire n_24372, n_24373, n_24374, n_24375, n_24376, n_24377, n_24378,
       n_24379;
  wire n_24380, n_24381, n_24382, n_24383, n_24384, n_24385, n_24386,
       n_24387;
  wire n_24388, n_24389, n_24390, n_24391, n_24392, n_24393, n_24394,
       n_24395;
  wire n_24396, n_24397, n_24398, n_24399, n_24400, n_24401, n_24402,
       n_24403;
  wire n_24404, n_24405, n_24406, n_24407, n_24408, n_24409, n_24410,
       n_24411;
  wire n_24412, n_24413, n_24414, n_24415, n_24416, n_24417, n_24418,
       n_24419;
  wire n_24420, n_24421, n_24422, n_24423, n_24424, n_24425, n_24426,
       n_24427;
  wire n_24428, n_24429, n_24430, n_24431, n_24432, n_24433, n_24434,
       n_24435;
  wire n_24436, n_24437, n_24438, n_24439, n_24440, n_24441, n_24442,
       n_24443;
  wire n_24444, n_24445, n_24446, n_24447, n_24448, n_24449, n_24450,
       n_24451;
  wire n_24452, n_24453, n_24454, n_24455, n_24456, n_24457, n_24458,
       n_24459;
  wire n_24460, n_24461, n_24462, n_24463, n_24464, n_24465, n_24466,
       n_24467;
  wire n_24468, n_24469, n_24470, n_24471, n_24472, n_24473, n_24474,
       n_24475;
  wire n_24476, n_24477, n_24478, n_24482, n_24483, n_24484, n_24485,
       n_24489;
  wire n_24490, n_24491, n_24492, n_24493, n_24494, n_24495, n_24496,
       n_24497;
  wire n_24498, n_24499, n_24500, n_24504, n_24505, n_24506, n_24507,
       n_24508;
  wire n_24509, n_24510, n_24511, n_24512, n_24513, n_24514, n_24515,
       n_24516;
  wire n_24517, n_24518, n_24519, n_24520, n_24521, n_24522, n_24523,
       n_24524;
  wire n_24525, n_24526, n_24527, n_24528, n_24529, n_24530, n_24531,
       n_24532;
  wire n_24533, n_24534, n_24535, n_24536, n_24537, n_24538, n_24539,
       n_24540;
  wire n_24541, n_24542, n_24543, n_24544, n_24545, n_24546, n_24547,
       n_24548;
  wire n_24549, n_24550, n_24551, n_24552, n_24553, n_24554, n_24555,
       n_24556;
  wire n_24557, n_24558, n_24559, n_24560, n_24561, n_24562, n_24563,
       n_24564;
  wire n_24565, n_24566, n_24567, n_24568, n_24569, n_24570, n_24571,
       n_24572;
  wire n_24573, n_24574, n_24575, n_24576, n_24577, n_24578, n_24579,
       n_24580;
  wire n_24581, n_24582, n_24583, n_24584, n_24585, n_24586, n_24587,
       n_24588;
  wire n_24589, n_24590, n_24591, n_24592, n_24593, n_24594, n_24595,
       n_24596;
  wire n_24597, n_24598, n_24599, n_24600, n_24601, n_24602, n_24603,
       n_24604;
  wire n_24605, n_24606, n_24607, n_24608, n_24609, n_24610, n_24611,
       n_24612;
  wire n_24613, n_24614, n_24615, n_24616, n_24617, n_24618, n_24619,
       n_24620;
  wire n_24621, n_24622, n_24623, n_24624, n_24625, n_24626, n_24627,
       n_24628;
  wire n_24629, n_24630, n_24631, n_24632, n_24633, n_24634, n_24635,
       n_24636;
  wire n_24637, n_24638, n_24639, n_24640, n_24641, n_24642, n_24643,
       n_24644;
  wire n_24645, n_24646, n_24649, n_24650, n_24651, n_24652, n_24653,
       n_24655;
  wire n_24656, n_24657, n_24658, n_24659, n_24660, n_24661, n_24662,
       n_24663;
  wire n_24664, n_24665, n_24666, n_24667, n_24668, n_24669, n_24670,
       n_24671;
  wire n_24672, n_24673, n_24674, n_24675, n_24676, n_24677, n_24678,
       n_24679;
  wire n_24680, n_24681, n_24682, n_24683, n_24684, n_24685, n_24686,
       n_24687;
  wire n_24688, n_24689, n_24690, n_24691, n_24692, n_24693, n_24694,
       n_24695;
  wire n_24696, n_24697, n_24698, n_24699, n_24700, n_24701, n_24702,
       n_24703;
  wire n_24704, n_24705, n_24706, n_24707, n_24708, n_24709, n_24710,
       n_24711;
  wire n_24712, n_24713, n_24714, n_24715, n_24716, n_24717, n_24718,
       n_24719;
  wire n_24720, n_24721, n_24722, n_24723, n_24724, n_24725, n_24726,
       n_24727;
  wire n_24728, n_24729, n_24730, n_24731, n_24732, n_24733, n_24734,
       n_24735;
  wire n_24736, n_24737, n_24738, n_24739, n_24740, n_24741, n_24742,
       n_24743;
  wire n_24744, n_24745, n_24746, n_24747, n_24748, n_24749, n_24750,
       n_24751;
  wire n_24752, n_24753, n_24754, n_24755, n_24756, n_24757, n_24758,
       n_24759;
  wire n_24760, n_24761, n_24762, n_24763, n_24764, n_24765, n_24766,
       n_24767;
  wire n_24769, n_24770, n_24771, n_24772, n_24773, n_24774, n_24775,
       n_24776;
  wire n_24777, n_24778, n_24779, n_24780, n_24781, n_24782, n_24783,
       n_24784;
  wire n_24785, n_24786, n_24787, n_24788, n_24789, n_24790, n_24791,
       n_24792;
  wire n_24793, n_24794, n_24795, n_24796, n_24797, n_24798, n_24799,
       n_24800;
  wire n_24801, n_24802, n_24803, n_24804, n_24805, n_24806, n_24807,
       n_24808;
  wire n_24809, n_24810, n_24811, n_24812, n_24813, n_24814, n_24815,
       n_24816;
  wire n_24817, n_24818, n_24819, n_24820, n_24821, n_24822, n_24823,
       n_24824;
  wire n_24825, n_24826, n_24827, n_24828, n_24829, n_24830, n_24831,
       n_24832;
  wire n_24833, n_24834, n_24835, n_24836, n_24837, n_24838, n_24839,
       n_24840;
  wire n_24841, n_24842, n_24843, n_24844, n_24845, n_24846, n_24847,
       n_24848;
  wire n_24849, n_24850, n_24851, n_24852, n_24853, n_24854, n_24855,
       n_24856;
  wire n_24857, n_24858, n_24859, n_24860, n_24861, n_24862, n_24863,
       n_24864;
  wire n_24865, n_24866, n_24867, n_24868, n_24869, n_24870, n_24871,
       n_24872;
  wire n_24873, n_24874, n_24875, n_24876, n_24877, n_24878, n_24879,
       n_24880;
  wire n_24881, n_24882, n_24883, n_24884, n_24885, n_24886, n_24887,
       n_24888;
  wire n_24889, n_24890, n_24891, n_24892, n_24893, n_24894, n_24895,
       n_24896;
  wire n_24897, n_24898, n_24899, n_24900, n_24901, n_24902, n_24903,
       n_24904;
  wire n_24905, n_24906, n_24907, n_24908, n_24909, n_24910, n_24911,
       n_24912;
  wire n_24913, n_24914, n_24915, n_24916, n_24917, n_24918, n_24919,
       n_24920;
  wire n_24922, n_24923, n_24924, n_24925, n_24926, n_24927, n_24928,
       n_24929;
  wire n_24930, n_24931, n_24932, n_24933, n_24936, n_24937, n_24938,
       n_24939;
  wire n_24940, n_24941, n_24942, n_24943, n_24944, n_24945, n_24946,
       n_24947;
  wire n_24948, n_24949, n_24950, n_24951, n_24952, n_24953, n_24954,
       n_24955;
  wire n_24956, n_24957, n_24958, n_24959, n_24960, n_24961, n_24962,
       n_24963;
  wire n_24964, n_24965, n_24966, n_24967, n_24968, n_24969, n_24970,
       n_24971;
  wire n_24972, n_24973, n_24974, n_24975, n_24976, n_24977, n_24978,
       n_24979;
  wire n_24980, n_24981, n_24982, n_24983, n_24984, n_24985, n_24986,
       n_24987;
  wire n_24988, n_24989, n_24990, n_24991, n_24992, n_24993, n_24994,
       n_24998;
  wire n_24999, n_25000, n_25001, n_25002, n_25003, n_25004, n_25005,
       n_25006;
  wire n_25007, n_25008, n_25009, n_25010, n_25011, n_25012, n_25013,
       n_25014;
  wire n_25015, n_25016, n_25017, n_25018, n_25019, n_25020, n_25021,
       n_25022;
  wire n_25023, n_25024, n_25025, n_25026, n_25027, n_25028, n_25029,
       n_25030;
  wire n_25031, n_25032, n_25033, n_25034, n_25035, n_25036, n_25037,
       n_25038;
  wire n_25039, n_25040, n_25041, n_25042, n_25043, n_25044, n_25045,
       n_25046;
  wire n_25047, n_25048, n_25049, n_25050, n_25051, n_25052, n_25053,
       n_25054;
  wire n_25055, n_25056, n_25057, n_25058, n_25059, n_25060, n_25061,
       n_25062;
  wire n_25063, n_25064, n_25065, n_25066, n_25067, n_25068, n_25069,
       n_25070;
  wire n_25071, n_25072, n_25073, n_25074, n_25075, n_25076, n_25077,
       n_25078;
  wire n_25079, n_25080, n_25081, n_25082, n_25083, n_25084, n_25085,
       n_25086;
  wire n_25087, n_25088, n_25089, n_25090, n_25091, n_25092, n_25093,
       n_25094;
  wire n_25095, n_25096, n_25097, n_25098, n_25099, n_25100, n_25101,
       n_25102;
  wire n_25103, n_25104, n_25105, n_25106, n_25107, n_25108, n_25109,
       n_25110;
  wire n_25111, n_25112, n_25113, n_25114, n_25115, n_25117, n_25118,
       n_25119;
  wire n_25120, n_25121, n_25122, n_25123, n_25124, n_25125, n_25126,
       n_25127;
  wire n_25128, n_25129, n_25130, n_25131, n_25132, n_25133, n_25134,
       n_25135;
  wire n_25136, n_25137, n_25138, n_25139, n_25140, n_25141, n_25142,
       n_25143;
  wire n_25144, n_25145, n_25146, n_25147, n_25148, n_25149, n_25150,
       n_25151;
  wire n_25152, n_25153, n_25155, n_25156, n_25157, n_25158, n_25159,
       n_25160;
  wire n_25161, n_25162, n_25163, n_25164, n_25165, n_25166, n_25167,
       n_25168;
  wire n_25169, n_25170, n_25171, n_25172, n_25173, n_25176, n_25177,
       n_25178;
  wire n_25179, n_25180, n_25181, n_25182, n_25183, n_25184, n_25185,
       n_25186;
  wire n_25187, n_25188, n_25189, n_25190, n_25191, n_25192, n_25193,
       n_25194;
  wire n_25195, n_25196, n_25197, n_25198, n_25199, n_25200, n_25201,
       n_25202;
  wire n_25203, n_25204, n_25205, n_25206, n_25207, n_25208, n_25209,
       n_25210;
  wire n_25211, n_25212, n_25213, n_25214, n_25215, n_25216, n_25217,
       n_25218;
  wire n_25219, n_25220, n_25221, n_25222, n_25223, n_25224, n_25225,
       n_25226;
  wire n_25227, n_25228, n_25229, n_25230, n_25231, n_25232, n_25233,
       n_25234;
  wire n_25235, n_25236, n_25237, n_25238, n_25239, n_25240, n_25241,
       n_25242;
  wire n_25243, n_25244, n_25245, n_25246, n_25247, n_25248, n_25249,
       n_25250;
  wire n_25251, n_25252, n_25253, n_25254, n_25255, n_25256, n_25257,
       n_25258;
  wire n_25259, n_25260, n_25261, n_25262, n_25263, n_25264, n_25265,
       n_25266;
  wire n_25267, n_25268, n_25269, n_25270, n_25271, n_25272, n_25273,
       n_25274;
  wire n_25275, n_25276, n_25277, n_25278, n_25279, n_25280, n_25281,
       n_25282;
  wire n_25283, n_25284, n_25285, n_25286, n_25287, n_25288, n_25289,
       n_25290;
  wire n_25291, n_25292, n_25293, n_25294, n_25295, n_25296, n_25297,
       n_25298;
  wire n_25299, n_25300, n_25301, n_25302, n_25303, n_25304, n_25305,
       n_25306;
  wire n_25307, n_25308, n_25309, n_25310, n_25311, n_25312, n_25313,
       n_25314;
  wire n_25315, n_25316, n_25317, n_25318, n_25319, n_25320, n_25321,
       n_25322;
  wire n_25323, n_25324, n_25325, n_25326, n_25327, n_25328, n_25329,
       n_25330;
  wire n_25331, n_25332, n_25333, n_25334, n_25335, n_25336, n_25337,
       n_25338;
  wire n_25339, n_25340, n_25341, n_25343, n_25344, n_25345, n_25346,
       n_25347;
  wire n_25348, n_25349, n_25350, n_25351, n_25352, n_25353, n_25354,
       n_25355;
  wire n_25356, n_25357, n_25358, n_25359, n_25360, n_25361, n_25362,
       n_25363;
  wire n_25364, n_25365, n_25366, n_25367, n_25368, n_25369, n_25370,
       n_25371;
  wire n_25372, n_25373, n_25374, n_25375, n_25376, n_25377, n_25378,
       n_25379;
  wire n_25380, n_25381, n_25382, n_25383, n_25384, n_25385, n_25386,
       n_25387;
  wire n_25388, n_25389, n_25390, n_25391, n_25392, n_25393, n_25394,
       n_25395;
  wire n_25396, n_25397, n_25398, n_25400, n_25401, n_25402, n_25403,
       n_25404;
  wire n_25405, n_25406, n_25407, n_25408, n_25409, n_25410, n_25411,
       n_25412;
  wire n_25413, n_25414, n_25415, n_25416, n_25417, n_25418, n_25419,
       n_25420;
  wire n_25421, n_25422, n_25423, n_25424, n_25425, n_25426, n_25427,
       n_25428;
  wire n_25429, n_25430, n_25431, n_25432, n_25433, n_25434, n_25435,
       n_25436;
  wire n_25437, n_25438, n_25439, n_25440, n_25441, n_25442, n_25443,
       n_25444;
  wire n_25445, n_25446, n_25447, n_25448, n_25449, n_25450, n_25451,
       n_25452;
  wire n_25453, n_25454, n_25455, n_25456, n_25457, n_25458, n_25459,
       n_25460;
  wire n_25461, n_25462, n_25463, n_25464, n_25465, n_25469, n_25470,
       n_25471;
  wire n_25472, n_25473, n_25474, n_25475, n_25476, n_25477, n_25478,
       n_25479;
  wire n_25480, n_25481, n_25482, n_25483, n_25484, n_25485, n_25486,
       n_25487;
  wire n_25488, n_25489, n_25490, n_25491, n_25492, n_25493, n_25494,
       n_25495;
  wire n_25496, n_25497, n_25498, n_25499, n_25500, n_25501, n_25502,
       n_25503;
  wire n_25504, n_25505, n_25506, n_25507, n_25508, n_25509, n_25510,
       n_25511;
  wire n_25512, n_25513, n_25514, n_25515, n_25516, n_25517, n_25518,
       n_25519;
  wire n_25520, n_25521, n_25522, n_25523, n_25524, n_25525, n_25526,
       n_25527;
  wire n_25528, n_25529, n_25530, n_25531, n_25532, n_25533, n_25534,
       n_25535;
  wire n_25536, n_25537, n_25538, n_25539, n_25540, n_25541, n_25542,
       n_25543;
  wire n_25544, n_25545, n_25546, n_25547, n_25548, n_25549, n_25550,
       n_25551;
  wire n_25552, n_25553, n_25554, n_25555, n_25556, n_25557, n_25558,
       n_25559;
  wire n_25560, n_25561, n_25562, n_25563, n_25564, n_25565, n_25568,
       n_25569;
  wire n_25570, n_25571, n_25572, n_25573, n_25574, n_25575, n_25576,
       n_25577;
  wire n_25578, n_25579, n_25580, n_25581, n_25582, n_25583, n_25584,
       n_25585;
  wire n_25586, n_25587, n_25588, n_25589, n_25590, n_25591, n_25592,
       n_25593;
  wire n_25594, n_25595, n_25596, n_25597, n_25598, n_25599, n_25600,
       n_25601;
  wire n_25602, n_25603, n_25604, n_25605, n_25606, n_25607, n_25608,
       n_25609;
  wire n_25610, n_25611, n_25612, n_25613, n_25614, n_25615, n_25616,
       n_25617;
  wire n_25618, n_25619, n_25620, n_25621, n_25622, n_25623, n_25624,
       n_25625;
  wire n_25626, n_25627, n_25628, n_25629, n_25630, n_25631, n_25632,
       n_25633;
  wire n_25634, n_25635, n_25636, n_25637, n_25638, n_25639, n_25640,
       n_25641;
  wire n_25644, n_25645, n_25646, n_25647, n_25648, n_25649, n_25650,
       n_25651;
  wire n_25652, n_25653, n_25654, n_25655, n_25656, n_25657, n_25658,
       n_25659;
  wire n_25660, n_25661, n_25662, n_25663, n_25664, n_25665, n_25666,
       n_25667;
  wire n_25668, n_25669, n_25670, n_25671, n_25672, n_25673, n_25674,
       n_25675;
  wire n_25676, n_25677, n_25678, n_25679, n_25680, n_25681, n_25682,
       n_25683;
  wire n_25684, n_25685, n_25686, n_25687, n_25688, n_25689, n_25690,
       n_25691;
  wire n_25692, n_25693, n_25694, n_25695, n_25696, n_25697, n_25698,
       n_25699;
  wire n_25700, n_25701, n_25702, n_25703, n_25704, n_25705, n_25706,
       n_25707;
  wire n_25709, n_25710, n_25711, n_25712, n_25713, n_25714, n_25715,
       n_25716;
  wire n_25717, n_25718, n_25719, n_25720, n_25721, n_25722, n_25723,
       n_25725;
  wire n_25726, n_25727, n_25728, n_25729, n_25730, n_25731, n_25732,
       n_25733;
  wire n_25735, n_25736, n_25737, n_25738, n_25739, n_25740, n_25741,
       n_25742;
  wire n_25743, n_25744, n_25745, n_25746, n_25747, n_25748, n_25749,
       n_25750;
  wire n_25751, n_25752, n_25753, n_25754, n_25755, n_25756, n_25757,
       n_25758;
  wire n_25759, n_25760, n_25761, n_25762, n_25763, n_25764, n_25765,
       n_25766;
  wire n_25767, n_25768, n_25769, n_25770, n_25771, n_25772, n_25773,
       n_25774;
  wire n_25775, n_25776, n_25777, n_25778, n_25779, n_25780, n_25781,
       n_25782;
  wire n_25783, n_25784, n_25785, n_25786, n_25787, n_25788, n_25789,
       n_25790;
  wire n_25791, n_25792, n_25793, n_25794, n_25795, n_25796, n_25797,
       n_25798;
  wire n_25799, n_25800, n_25801, n_25802, n_25803, n_25804, n_25805,
       n_25806;
  wire n_25807, n_25808, n_25809, n_25810, n_25811, n_25812, n_25813,
       n_25814;
  wire n_25815, n_25816, n_25817, n_25818, n_25819, n_25820, n_25822,
       n_25823;
  wire n_25824, n_25825, n_25826, n_25827, n_25828, n_25829, n_25830,
       n_25831;
  wire n_25832, n_25834, n_25835, n_25836, n_25837, n_25838, n_25839,
       n_25840;
  wire n_25841, n_25843, n_25844, n_25845, n_25846, n_25847, n_25848,
       n_25849;
  wire n_25850, n_25851, n_25852, n_25853, n_25854, n_25855, n_25856,
       n_25857;
  wire n_25858, n_25859, n_25860, n_25861, n_25862, n_25863, n_25864,
       n_25865;
  wire n_25866, n_25867, n_25868, n_25869, n_25870, n_25871, n_25872,
       n_25873;
  wire n_25874, n_25875, n_25876, n_25878, n_25879, n_25880, n_25881,
       n_25882;
  wire n_25883, n_25884, n_25885, n_25886, n_25887, n_25888, n_25889,
       n_25890;
  wire n_25891, n_25892, n_25893, n_25894, n_25895, n_25896, n_25897,
       n_25898;
  wire n_25899, n_25900, n_25901, n_25902, n_25903, n_25904, n_25905,
       n_25906;
  wire n_25907, n_25908, n_25909, n_25910, n_25911, n_25912, n_25913,
       n_25914;
  wire n_25915, n_25916, n_25917, n_25918, n_25919, n_25920, n_25921,
       n_25922;
  wire n_25923, n_25924, n_25925, n_25926, n_25927, n_25928, n_25929,
       n_25930;
  wire n_25931, n_25932, n_25933, n_25934, n_25936, n_25937, n_25938,
       n_25939;
  wire n_25940, n_25941, n_25942, n_25943, n_25944, n_25945, n_25946,
       n_25947;
  wire n_25948, n_25949, n_25950, n_25951, n_25952, n_25953, n_25954,
       n_25955;
  wire n_25956, n_25957, n_25958, n_25959, n_25960, n_25961, n_25962,
       n_25963;
  wire n_25964, n_25965, n_25966, n_25967, n_25968, n_25969, n_25970,
       n_25971;
  wire n_25972, n_25973, n_25974, n_25975, n_25976, n_25977, n_25978,
       n_25979;
  wire n_25980, n_25981, n_25982, n_25983, n_25984, n_25985, n_25986,
       n_25987;
  wire n_25988, n_25989, n_25990, n_25991, n_25992, n_25993, n_25994,
       n_25995;
  wire n_25996, n_25997, n_25998, n_25999, n_26000, n_26001, n_26002,
       n_26003;
  wire n_26004, n_26005, n_26006, n_26007, n_26008, n_26009, n_26010,
       n_26011;
  wire n_26012, n_26013, n_26014, n_26015, n_26016, n_26017, n_26018,
       n_26019;
  wire n_26020, n_26021, n_26022, n_26023, n_26024, n_26025, n_26026,
       n_26027;
  wire n_26028, n_26029, n_26030, n_26031, n_26032, n_26033, n_26034,
       n_26035;
  wire n_26036, n_26037, n_26038, n_26039, n_26040, n_26041, n_26042,
       n_26043;
  wire n_26044, n_26045, n_26046, n_26047, n_26048, n_26049, n_26050,
       n_26051;
  wire n_26052, n_26053, n_26054, n_26055, n_26056, n_26057, n_26058,
       n_26059;
  wire n_26060, n_26061, n_26062, n_26063, n_26064, n_26065, n_26066,
       n_26067;
  wire n_26068, n_26069, n_26070, n_26071, n_26072, n_26073, n_26074,
       n_26075;
  wire n_26076, n_26077, n_26078, n_26079, n_26080, n_26081, n_26082,
       n_26083;
  wire n_26084, n_26085, n_26086, n_26087, n_26088, n_26089, n_26090,
       n_26091;
  wire n_26092, n_26093, n_26094, n_26099, n_26100, n_26101, n_26102,
       n_26103;
  wire n_26104, n_26105, n_26106, n_26107, n_26108, n_26109, n_26110,
       n_26111;
  wire n_26112, n_26113, n_26114, n_26115, n_26116, n_26117, n_26118,
       n_26119;
  wire n_26120, n_26121, n_26122, n_26123, n_26124, n_26125, n_26126,
       n_26127;
  wire n_26128, n_26129, n_26130, n_26131, n_26132, n_26133, n_26134,
       n_26135;
  wire n_26136, n_26137, n_26138, n_26139, n_26140, n_26141, n_26142,
       n_26143;
  wire n_26144, n_26145, n_26146, n_26147, n_26148, n_26149, n_26150,
       n_26151;
  wire n_26152, n_26153, n_26154, n_26155, n_26156, n_26157, n_26158,
       n_26159;
  wire n_26160, n_26161, n_26162, n_26163, n_26164, n_26165, n_26166,
       n_26167;
  wire n_26168, n_26169, n_26170, n_26171, n_26172, n_26173, n_26174,
       n_26175;
  wire n_26176, n_26177, n_26178, n_26179, n_26180, n_26181, n_26182,
       n_26183;
  wire n_26184, n_26185, n_26186, n_26187, n_26188, n_26189, n_26190,
       n_26191;
  wire n_26192, n_26193, n_26194, n_26195, n_26196, n_26197, n_26198,
       n_26199;
  wire n_26200, n_26201, n_26202, n_26203, n_26204, n_26205, n_26206,
       n_26207;
  wire n_26208, n_26209, n_26210, n_26211, n_26212, n_26213, n_26214,
       n_26215;
  wire n_26216, n_26217, n_26218, n_26219, n_26220, n_26221, n_26222,
       n_26223;
  wire n_26224, n_26225, n_26226, n_26227, n_26228, n_26229, n_26230,
       n_26231;
  wire n_26232, n_26233, n_26234, n_26235, n_26236, n_26237, n_26238,
       n_26239;
  wire n_26240, n_26241, n_26242, n_26243, n_26244, n_26246, n_26247,
       n_26248;
  wire n_26249, n_26250, n_26251, n_26252, n_26253, n_26254, n_26255,
       n_26256;
  wire n_26257, n_26258, n_26259, n_26260, n_26262, n_26263, n_26264,
       n_26265;
  wire n_26266, n_26267, n_26268, n_26269, n_26270, n_26271, n_26272,
       n_26273;
  wire n_26274, n_26275, n_26276, n_26277, n_26278, n_26279, n_26280,
       n_26281;
  wire n_26282, n_26283, n_26284, n_26285, n_26286, n_26287, n_26288,
       n_26289;
  wire n_26290, n_26291, n_26292, n_26293, n_26294, n_26295, n_26296,
       n_26297;
  wire n_26298, n_26299, n_26300, n_26301, n_26303, n_26304, n_26305,
       n_26306;
  wire n_26307, n_26308, n_26309, n_26310, n_26311, n_26312, n_26313,
       n_26314;
  wire n_26315, n_26316, n_26317, n_26318, n_26319, n_26320, n_26321,
       n_26322;
  wire n_26323, n_26324, n_26325, n_26326, n_26327, n_26328, n_26329,
       n_26330;
  wire n_26331, n_26332, n_26333, n_26334, n_26336, n_26337, n_26338,
       n_26339;
  wire n_26340, n_26341, n_26342, n_26343, n_26344, n_26345, n_26346,
       n_26347;
  wire n_26348, n_26349, n_26350, n_26351, n_26352, n_26353, n_26354,
       n_26355;
  wire n_26356, n_26357, n_26358, n_26359, n_26360, n_26361, n_26362,
       n_26363;
  wire n_26364, n_26365, n_26366, n_26367, n_26368, n_26369, n_26370,
       n_26372;
  wire n_26373, n_26374, n_26375, n_26376, n_26377, n_26378, n_26379,
       n_26380;
  wire n_26381, n_26382, n_26383, n_26384, n_26385, n_26386, n_26387,
       n_26388;
  wire n_26389, n_26390, n_26391, n_26392, n_26393, n_26394, n_26395,
       n_26396;
  wire n_26397, n_26398, n_26399, n_26400, n_26401, n_26402, n_26403,
       n_26404;
  wire n_26405, n_26406, n_26407, n_26408, n_26409, n_26410, n_26411,
       n_26412;
  wire n_26413, n_26414, n_26415, n_26416, n_26417, n_26421, n_26422,
       n_26423;
  wire n_26424, n_26425, n_26426, n_26427, n_26428, n_26429, n_26430,
       n_26431;
  wire n_26432, n_26433, n_26434, n_26435, n_26436, n_26437, n_26438,
       n_26439;
  wire n_26440, n_26441, n_26442, n_26443, n_26444, n_26445, n_26446,
       n_26447;
  wire n_26448, n_26449, n_26450, n_26451, n_26452, n_26453, n_26454,
       n_26455;
  wire n_26456, n_26457, n_26458, n_26459, n_26460, n_26461, n_26462,
       n_26463;
  wire n_26464, n_26465, n_26466, n_26467, n_26468, n_26469, n_26470,
       n_26471;
  wire n_26472, n_26473, n_26474, n_26475, n_26476, n_26477, n_26478,
       n_26479;
  wire n_26480, n_26481, n_26482, n_26483, n_26484, n_26485, n_26486,
       n_26487;
  wire n_26488, n_26489, n_26490, n_26491, n_26492, n_26493, n_26494,
       n_26495;
  wire n_26496, n_26497, n_26498, n_26499, n_26500, n_26501, n_26502,
       n_26503;
  wire n_26504, n_26505, n_26506, n_26507, n_26508, n_26509, n_26510,
       n_26511;
  wire n_26512, n_26513, n_26514, n_26515, n_26516, n_26517, n_26518,
       n_26519;
  wire n_26520, n_26521, n_26522, n_26523, n_26524, n_26525, n_26526,
       n_26527;
  wire n_26528, n_26529, n_26530, n_26531, n_26532, n_26533, n_26534,
       n_26535;
  wire n_26536, n_26537, n_26538, n_26539, n_26540, n_26541, n_26542,
       n_26543;
  wire n_26544, n_26546, n_26547, n_26548, n_26549, n_26550, n_26551,
       n_26552;
  wire n_26553, n_26554, n_26555, n_26556, n_26557, n_26558, n_26559,
       n_26560;
  wire n_26561, n_26562, n_26563, n_26564, n_26565, n_26566, n_26567,
       n_26568;
  wire n_26569, n_26570, n_26571, n_26572, n_26573, n_26574, n_26575,
       n_26576;
  wire n_26577, n_26578, n_26579, n_26580, n_26581, n_26582, n_26583,
       n_26584;
  wire n_26585, n_26586, n_26587, n_26588, n_26589, n_26590, n_26591,
       n_26592;
  wire n_26593, n_26594, n_26595, n_26596, n_26597, n_26598, n_26599,
       n_26600;
  wire n_26602, n_26604, n_26605, n_26606, n_26607, n_26608, n_26609,
       n_26610;
  wire n_26611, n_26612, n_26613, n_26614, n_26615, n_26616, n_26617,
       n_26618;
  wire n_26619, n_26620, n_26621, n_26622, n_26623, n_26624, n_26625,
       n_26626;
  wire n_26627, n_26628, n_26629, n_26630, n_26631, n_26632, n_26633,
       n_26634;
  wire n_26635, n_26636, n_26637, n_26638, n_26639, n_26640, n_26641,
       n_26642;
  wire n_26643, n_26644, n_26645, n_26646, n_26647, n_26648, n_26649,
       n_26650;
  wire n_26651, n_26652, n_26653, n_26654, n_26655, n_26656, n_26657,
       n_26658;
  wire n_26659, n_26660, n_26661, n_26662, n_26663, n_26664, n_26665,
       n_26666;
  wire n_26667, n_26668, n_26669, n_26670, n_26671, n_26672, n_26673,
       n_26674;
  wire n_26675, n_26676, n_26677, n_26678, n_26679, n_26680, n_26681,
       n_26682;
  wire n_26683, n_26684, n_26685, n_26686, n_26687, n_26688, n_26689,
       n_26690;
  wire n_26691, n_26692, n_26693, n_26694, n_26695, n_26696, n_26697,
       n_26698;
  wire n_26699, n_26700, n_26701, n_26702, n_26705, n_26706, n_26707,
       n_26708;
  wire n_26709, n_26710, n_26711, n_26712, n_26713, n_26714, n_26715,
       n_26716;
  wire n_26717, n_26718, n_26719, n_26721, n_26722, n_26723, n_26724,
       n_26725;
  wire n_26726, n_26727, n_26728, n_26729, n_26730, n_26731, n_26732,
       n_26733;
  wire n_26735, n_26736, n_26737, n_26738, n_26739, n_26740, n_26742,
       n_26743;
  wire n_26744, n_26745, n_26746, n_26747, n_26748, n_26749, n_26750,
       n_26751;
  wire n_26752, n_26753, n_26754, n_26756, n_26757, n_26758, n_26759,
       n_26760;
  wire n_26761, n_26762, n_26763, n_26764, n_26765, n_26766, n_26767,
       n_26768;
  wire n_26769, n_26770, n_26771, n_26772, n_26773, n_26774, n_26776,
       n_26777;
  wire n_26778, n_26779, n_26780, n_26781, n_26782, n_26783, n_26784,
       n_26785;
  wire n_26786, n_26787, n_26788, n_26789, n_26790, n_26791, n_26792,
       n_26793;
  wire n_26794, n_26795, n_26796, n_26797, n_26798, n_26799, n_26800,
       n_26801;
  wire n_26802, n_26803, n_26804, n_26805, n_26806, n_26807, n_26808,
       n_26809;
  wire n_26810, n_26811, n_26812, n_26813, n_26814, n_26815, n_26816,
       n_26817;
  wire n_26818, n_26819, n_26820, n_26821, n_26822, n_26823, n_26824,
       n_26825;
  wire n_26826, n_26827, n_26828, n_26829, n_26830, n_26831, n_26832,
       n_26833;
  wire n_26834, n_26837, n_26838, n_26839, n_26840, n_26841, n_26842,
       n_26843;
  wire n_26844, n_26845, n_26846, n_26847, n_26848, n_26849, n_26850,
       n_26851;
  wire n_26852, n_26853, n_26854, n_26855, n_26856, n_26857, n_26858,
       n_26859;
  wire n_26860, n_26861, n_26862, n_26863, n_26864, n_26865, n_26866,
       n_26867;
  wire n_26868, n_26869, n_26870, n_26871, n_26872, n_26873, n_26880,
       n_26881;
  wire n_26882, n_26883, n_26884, n_26885, n_26886, n_26887, n_26888,
       n_26889;
  wire n_26890, n_26891, n_26892, n_26893, n_26894, n_26895, n_26896,
       n_26897;
  wire n_26898, n_26899, n_26900, n_26901, n_26902, n_26903, n_26904,
       n_26905;
  wire n_26906, n_26907, n_26908, n_26909, n_26910, n_26911, n_26912,
       n_26913;
  wire n_26914, n_26915, n_26916, n_26917, n_26918, n_26919, n_26920,
       n_26921;
  wire n_26922, n_26923, n_26924, n_26925, n_26926, n_26927, n_26928,
       n_26929;
  wire n_26930, n_26931, n_26932, n_26933, n_26934, n_26935, n_26936,
       n_26937;
  wire n_26938, n_26939, n_26940, n_26941, n_26942, n_26943, n_26944,
       n_26945;
  wire n_26946, n_26947, n_26948, n_26949, n_26950, n_26951, n_26952,
       n_26953;
  wire n_26954, n_26955, n_26956, n_26957, n_26958, n_26959, n_26960,
       n_26961;
  wire n_26962, n_26963, n_26964, n_26965, n_26966, n_26967, n_26968,
       n_26969;
  wire n_26970, n_26971, n_26972, n_26973, n_26974, n_26975, n_26976,
       n_26977;
  wire n_26978, n_26982, n_26983, n_26984, n_26985, n_26986, n_26987,
       n_26988;
  wire n_26989, n_26990, n_26991, n_26992, n_26993, n_26994, n_26995,
       n_26996;
  wire n_26997, n_26998, n_26999, n_27000, n_27001, n_27002, n_27003,
       n_27004;
  wire n_27005, n_27006, n_27007, n_27008, n_27009, n_27010, n_27011,
       n_27012;
  wire n_27013, n_27014, n_27015, n_27016, n_27017, n_27018, n_27019,
       n_27020;
  wire n_27021, n_27022, n_27023, n_27024, n_27025, n_27026, n_27027,
       n_27028;
  wire n_27029, n_27030, n_27031, n_27032, n_27033, n_27034, n_27035,
       n_27036;
  wire n_27037, n_27038, n_27039, n_27040, n_27041, n_27042, n_27043,
       n_27044;
  wire n_27045, n_27046, n_27047, n_27048, n_27049, n_27050, n_27051,
       n_27052;
  wire n_27053, n_27054, n_27055, n_27056, n_27057, n_27058, n_27059,
       n_27060;
  wire n_27061, n_27062, n_27063, n_27064, n_27065, n_27066, n_27067,
       n_27068;
  wire n_27069, n_27070, n_27071, n_27072, n_27073, n_27074, n_27075,
       n_27076;
  wire n_27077, n_27078, n_27079, n_27080, n_27081, n_27082, n_27083,
       n_27084;
  wire n_27085, n_27086, n_27087, n_27088, n_27089, n_27090, n_27091,
       n_27092;
  wire n_27093, n_27094, n_27095, n_27096, n_27097, n_27098, n_27099,
       n_27100;
  wire n_27101, n_27102, n_27103, n_27104, n_27105, n_27106, n_27107,
       n_27108;
  wire n_27109, n_27110, n_27111, n_27112, n_27113, n_27114, n_27115,
       n_27116;
  wire n_27117, n_27118, n_27119, n_27120, n_27121, n_27122, n_27123,
       n_27124;
  wire n_27125, n_27126, n_27127, n_27128, n_27129, n_27130, n_27131,
       n_27132;
  wire n_27133, n_27134, n_27135, n_27136, n_27137, n_27138, n_27139,
       n_27140;
  wire n_27141, n_27142, n_27143, n_27144, n_27145, n_27146, n_27147,
       n_27148;
  wire n_27149, n_27150, n_27151, n_27152, n_27153, n_27156, n_27157,
       n_27158;
  wire n_27159, n_27160, n_27161, n_27162, n_27163, n_27164, n_27165,
       n_27166;
  wire n_27167, n_27168, n_27169, n_27170, n_27171, n_27172, n_27173,
       n_27174;
  wire n_27175, n_27176, n_27177, n_27178, n_27179, n_27180, n_27181,
       n_27182;
  wire n_27183, n_27184, n_27185, n_27186, n_27187, n_27188, n_27189,
       n_27190;
  wire n_27191, n_27192, n_27193, n_27194, n_27195, n_27196, n_27197,
       n_27198;
  wire n_27199, n_27200, n_27201, n_27202, n_27203, n_27204, n_27205,
       n_27206;
  wire n_27207, n_27208, n_27209, n_27210, n_27211, n_27212, n_27213,
       n_27214;
  wire n_27215, n_27216, n_27217, n_27218, n_27219, n_27220, n_27221,
       n_27222;
  wire n_27223, n_27224, n_27225, n_27226, n_27227, n_27228, n_27229,
       n_27230;
  wire n_27231, n_27232, n_27233, n_27234, n_27235, n_27236, n_27237,
       n_27238;
  wire n_27239, n_27240, n_27241, n_27242, n_27243, n_27244, n_27245,
       n_27246;
  wire n_27247, n_27248, n_27249, n_27250, n_27251, n_27252, n_27253,
       n_27254;
  wire n_27255, n_27256, n_27257, n_27258, n_27259, n_27260, n_27261,
       n_27262;
  wire n_27263, n_27264, n_27265, n_27266, n_27267, n_27268, n_27269,
       n_27270;
  wire n_27271, n_27272, n_27273, n_27274, n_27275, n_27276, n_27277,
       n_27278;
  wire n_27279, n_27280, n_27281, n_27282, n_27283, n_27284, n_27285,
       n_27286;
  wire n_27287, n_27288, n_27289, n_27290, n_27291, n_27292, n_27293,
       n_27294;
  wire n_27295, n_27296, n_27297, n_27298, n_27299, n_27300, n_27301,
       n_27302;
  wire n_27303, n_27304, n_27305, n_27306, n_27307, n_27308, n_27309,
       n_27310;
  wire n_27311, n_27312, n_27313, n_27314, n_27315, n_27316, n_27317,
       n_27318;
  wire n_27319, n_27320, n_27321, n_27322, n_27323, n_27324, n_27325,
       n_27326;
  wire n_27327, n_27328, n_27329, n_27330, n_27331, n_27332, n_27333,
       n_27334;
  wire n_27335, n_27336, n_27337, n_27338, n_27339, n_27340, n_27341,
       n_27342;
  wire n_27349, n_27350, n_27351, n_27352, n_27353, n_27354, n_27355,
       n_27356;
  wire n_27357, n_27358, n_27359, n_27360, n_27361, n_27362, n_27363,
       n_27364;
  wire n_27365, n_27366, n_27367, n_27368, n_27369, n_27370, n_27371,
       n_27372;
  wire n_27373, n_27374, n_27375, n_27376, n_27377, n_27378, n_27379,
       n_27380;
  wire n_27381, n_27382, n_27383, n_27384, n_27385, n_27386, n_27387,
       n_27388;
  wire n_27389, n_27390, n_27391, n_27392, n_27393, n_27394, n_27395,
       n_27396;
  wire n_27397, n_27398, n_27399, n_27400, n_27401, n_27402, n_27403,
       n_27404;
  wire n_27405, n_27406, n_27407, n_27408, n_27409, n_27410, n_27411,
       n_27412;
  wire n_27413, n_27414, n_27415, n_27416, n_27417, n_27418, n_27419,
       n_27420;
  wire n_27421, n_27422, n_27423, n_27424, n_27425, n_27426, n_27427,
       n_27428;
  wire n_27429, n_27430, n_27431, n_27432, n_27433, n_27434, n_27435,
       n_27436;
  wire n_27437, n_27438, n_27439, n_27440, n_27441, n_27442, n_27443,
       n_27444;
  wire n_27445, n_27446, n_27447, n_27448, n_27449, n_27450, n_27451,
       n_27452;
  wire n_27453, n_27454, n_27455, n_27456, n_27457, n_27458, n_27459,
       n_27460;
  wire n_27461, n_27462, n_27463, n_27464, n_27465, n_27466, n_27467,
       n_27468;
  wire n_27469, n_27470, n_27471, n_27472, n_27473, n_27474, n_27475,
       n_27476;
  wire n_27477, n_27478, n_27479, n_27480, n_27481, n_27482, n_27483,
       n_27484;
  wire n_27485, n_27486, n_27487, n_27488, n_27489, n_27490, n_27491,
       n_27492;
  wire n_27493, n_27494, n_27495, n_27496, n_27497, n_27498, n_27499,
       n_27500;
  wire n_27501, n_27502, n_27503, n_27504, n_27505, n_27506, n_27507,
       n_27508;
  wire n_27509, n_27510, n_27511, n_27512, n_27513, n_27514, n_27515,
       n_27516;
  wire n_27517, n_27518, n_27519, n_27520, n_27521, n_27522, n_27523,
       n_27524;
  wire n_27525, n_27526, n_27527, n_27528, n_27529, n_27530, n_27531,
       n_27532;
  wire n_27533, n_27534, n_27535, n_27536, n_27537, n_27538, n_27539,
       n_27540;
  wire n_27541, n_27542, n_27543, n_27544, n_27545, n_27546, n_27547,
       n_27548;
  wire n_27549, n_27550, n_27551, n_27552, n_27553, n_27554, n_27555,
       n_27556;
  wire n_27557, n_27558, n_27559, n_27560, n_27561, n_27562, n_27563,
       n_27564;
  wire n_27565, n_27566, n_27567, n_27568, n_27569, n_27570, n_27571,
       n_27572;
  wire n_27573, n_27574, n_27575, n_27576, n_27577, n_27578, n_27579,
       n_27580;
  wire n_27581, n_27582, n_27583, n_27584, n_27585, n_27586, n_27587,
       n_27588;
  wire n_27589, n_27590, n_27591, n_27592, n_27593, n_27594, n_27595,
       n_27596;
  wire n_27598, n_27599, n_27600, n_27601, n_27602, n_27603, n_27604,
       n_27605;
  wire n_27606, n_27607, n_27608, n_27609, n_27610, n_27611, n_27614,
       n_27615;
  wire n_27616, n_27617, n_27618, n_27619, n_27620, n_27621, n_27622,
       n_27623;
  wire n_27624, n_27625, n_27626, n_27627, n_27628, n_27632, n_27633,
       n_27634;
  wire n_27635, n_27636, n_27637, n_27638, n_27639, n_27640, n_27641,
       n_27642;
  wire n_27643, n_27644, n_27648, n_27649, n_27650, n_27651, n_27652,
       n_27653;
  wire n_27654, n_27655, n_27656, n_27657, n_27658, n_27661, n_27662,
       n_27663;
  wire n_27664, n_27665, n_27666, n_27667, n_27668, n_27669, n_27670,
       n_27671;
  wire n_27672, n_27673, n_27674, n_27675, n_27676, n_27677, n_27678,
       n_27679;
  wire n_27680, n_27681, n_27682, n_27683, n_27684, n_27685, n_27686,
       n_27687;
  wire n_27688, n_27689, n_27690, n_27691, n_27692, n_27693, n_27694,
       n_27695;
  wire n_27696, n_27697, n_27698, n_27699, n_27700, n_27701, n_27702,
       n_27703;
  wire n_27704, n_27705, n_27706, n_27707, n_27708, n_27709, n_27710,
       n_27711;
  wire n_27712, n_27713, n_27714, n_27715, n_27716, n_27717, n_27718,
       n_27719;
  wire n_27720, n_27721, n_27722, n_27723, n_27724, n_27725, n_27726,
       n_27727;
  wire n_27728, n_27729, n_27730, n_27731, n_27732, n_27733, n_27734,
       n_27735;
  wire n_27736, n_27737, n_27738, n_27739, n_27740, n_27741, n_27742,
       n_27743;
  wire n_27744, n_27745, n_27746, n_27747, n_27748, n_27749, n_27750,
       n_27751;
  wire n_27752, n_27753, n_27754, n_27755, n_27756, n_27757, n_27758,
       n_27759;
  wire n_27760, n_27761, n_27762, n_27763, n_27764, n_27765, n_27766,
       n_27767;
  wire n_27768, n_27769, n_27770, n_27771, n_27772, n_27779, n_27780,
       n_27781;
  wire n_27782, n_27783, n_27784, n_27785, n_27786, n_27787, n_27788,
       n_27789;
  wire n_27793, n_27794, n_27795, n_27796, n_27797, n_27798, n_27799,
       n_27800;
  wire n_27801, n_27802, n_27803, n_27804, n_27805, n_27806, n_27807,
       n_27808;
  wire n_27809, n_27810, n_27811, n_27812, n_27813, n_27814, n_27815,
       n_27816;
  wire n_27817, n_27818, n_27819, n_27820, n_27821, n_27822, n_27823,
       n_27824;
  wire n_27825, n_27826, n_27827, n_27828, n_27829, n_27830, n_27831,
       n_27832;
  wire n_27833, n_27834, n_27835, n_27836, n_27837, n_27838, n_27839,
       n_27840;
  wire n_27841, n_27842, n_27843, n_27844, n_27845, n_27846, n_27847,
       n_27848;
  wire n_27849, n_27850, n_27851, n_27852, n_27853, n_27854, n_27855,
       n_27856;
  wire n_27857, n_27858, n_27859, n_27860, n_27861, n_27862, n_27863,
       n_27864;
  wire n_27865, n_27866, n_27867, n_27868, n_27869, n_27870, n_27871,
       n_27872;
  wire n_27873, n_27874, n_27875, n_27876, n_27877, n_27878, n_27879,
       n_27880;
  wire n_27881, n_27882, n_27883, n_27884, n_27885, n_27886, n_27887,
       n_27888;
  wire n_27889, n_27890, n_27891, n_27892, n_27893, n_27894, n_27895,
       n_27896;
  wire n_27897, n_27898, n_27899, n_27900, n_27901, n_27902, n_27903,
       n_27904;
  wire n_27905, n_27906, n_27907, n_27908, n_27909, n_27910, n_27911,
       n_27912;
  wire n_27913, n_27914, n_27915, n_27916, n_27917, n_27918, n_27919,
       n_27920;
  wire n_27921, n_27922, n_27923, n_27924, n_27925, n_27926, n_27927,
       n_27928;
  wire n_27929, n_27930, n_27931, n_27932, n_27933, n_27934, n_27935,
       n_27939;
  wire n_27940, n_27941, n_27942, n_27943, n_27944, n_27945, n_27946,
       n_27947;
  wire n_27948, n_27949, n_27950, n_27951, n_27952, n_27953, n_27954,
       n_27955;
  wire n_27956, n_27957, n_27958, n_27959, n_27960, n_27961, n_27962,
       n_27963;
  wire n_27964, n_27965, n_27966, n_27967, n_27968, n_27969, n_27970,
       n_27971;
  wire n_27972, n_27973, n_27974, n_27975, n_27976, n_27977, n_27978,
       n_27979;
  wire n_27980, n_27981, n_27982, n_27983, n_27984, n_27985, n_27986,
       n_27987;
  wire n_27988, n_27989, n_27990, n_27991, n_27992, n_27993, n_27994,
       n_27995;
  wire n_27996, n_27997, n_27998, n_27999, n_28000, n_28001, n_28002,
       n_28003;
  wire n_28004, n_28005, n_28006, n_28007, n_28008, n_28009, n_28010,
       n_28011;
  wire n_28012, n_28013, n_28014, n_28015, n_28016, n_28017, n_28018,
       n_28019;
  wire n_28020, n_28021, n_28022, n_28023, n_28024, n_28025, n_28026,
       n_28027;
  wire n_28028, n_28029, n_28030, n_28031, n_28032, n_28033, n_28034,
       n_28035;
  wire n_28036, n_28037, n_28038, n_28039, n_28040, n_28041, n_28042,
       n_28043;
  wire n_28044, n_28045, n_28046, n_28047, n_28048, n_28049, n_28050,
       n_28051;
  wire n_28055, n_28056, n_28057, n_28058, n_28059, n_28060, n_28061,
       n_28062;
  wire n_28063, n_28064, n_28065, n_28066, n_28067, n_28068, n_28069,
       n_28070;
  wire n_28071, n_28072, n_28073, n_28074, n_28075, n_28076, n_28077,
       n_28080;
  wire n_28081, n_28082, n_28083, n_28084, n_28085, n_28086, n_28087,
       n_28088;
  wire n_28089, n_28090, n_28091, n_28092, n_28093, n_28094, n_28095,
       n_28096;
  wire n_28097, n_28098, n_28099, n_28100, n_28101, n_28102, n_28103,
       n_28104;
  wire n_28105, n_28106, n_28107, n_28108, n_28109, n_28110, n_28111,
       n_28112;
  wire n_28113, n_28114, n_28115, n_28116, n_28117, n_28118, n_28119,
       n_28120;
  wire n_28121, n_28122, n_28123, n_28124, n_28125, n_28126, n_28127,
       n_28128;
  wire n_28129, n_28130, n_28131, n_28132, n_28133, n_28134, n_28135,
       n_28136;
  wire n_28137, n_28138, n_28139, n_28140, n_28141, n_28142, n_28143,
       n_28144;
  wire n_28145, n_28146, n_28147, n_28148, n_28149, n_28150, n_28151,
       n_28152;
  wire n_28153, n_28154, n_28155, n_28156, n_28157, n_28158, n_28159,
       n_28160;
  wire n_28161, n_28162, n_28163, n_28164, n_28165, n_28166, n_28167,
       n_28168;
  wire n_28169, n_28170, n_28171, n_28172, n_28173, n_28174, n_28175,
       n_28176;
  wire n_28177, n_28178, n_28179, n_28180, n_28181, n_28182, n_28183,
       n_28184;
  wire n_28185, n_28186, n_28187, n_28188, n_28189, n_28190, n_28191,
       n_28192;
  wire n_28193, n_28194, n_28195, n_28196, n_28197, n_28198, n_28199,
       n_28200;
  wire n_28201, n_28202, n_28203, n_28204, n_28205, n_28206, n_28207,
       n_28208;
  wire n_28209, n_28210, n_28211, n_28212, n_28213, n_28214, n_28215,
       n_28216;
  wire n_28217, n_28218, n_28219, n_28220, n_28221, n_28222, n_28223,
       n_28224;
  wire n_28225, n_28226, n_28227, n_28228, n_28229, n_28230, n_28231,
       n_28232;
  wire n_28233, n_28234, n_28235, n_28236, n_28237, n_28238, n_28239,
       n_28240;
  wire n_28241, n_28242, n_28243, n_28244, n_28245, n_28246, n_28247,
       n_28248;
  wire n_28249, n_28250, n_28251, n_28252, n_28253, n_28254, n_28255,
       n_28256;
  wire n_28257, n_28258, n_28259, n_28260, n_28261, n_28262, n_28263,
       n_28264;
  wire n_28265, n_28266, n_28267, n_28268, n_28269, n_28270, n_28271,
       n_28272;
  wire n_28273, n_28274, n_28275, n_28276, n_28277, n_28278, n_28279,
       n_28280;
  wire n_28281, n_28282, n_28283, n_28284, n_28285, n_28286, n_28287,
       n_28288;
  wire n_28289, n_28290, n_28291, n_28292, n_28293, n_28294, n_28295,
       n_28296;
  wire n_28297, n_28298, n_28299, n_28300, n_28301, n_28302, n_28303,
       n_28304;
  wire n_28305, n_28306, n_28307, n_28308, n_28309, n_28311, n_28312,
       n_28313;
  wire n_28314, n_28315, n_28316, n_28317, n_28318, n_28319, n_28320,
       n_28321;
  wire n_28322, n_28323, n_28324, n_28325, n_28326, n_28327, n_28328,
       n_28329;
  wire n_28330, n_28331, n_28332, n_28333, n_28334, n_28335, n_28336,
       n_28337;
  wire n_28338, n_28339, n_28340, n_28341, n_28342, n_28343, n_28344,
       n_28345;
  wire n_28346, n_28347, n_28348, n_28349, n_28350, n_28351, n_28352,
       n_28353;
  wire n_28354, n_28355, n_28356, n_28357, n_28358, n_28359, n_28360,
       n_28361;
  wire n_28362, n_28363, n_28364, n_28365, n_28366, n_28367, n_28368,
       n_28369;
  wire n_28370, n_28371, n_28372, n_28373, n_28374, n_28375, n_28376,
       n_28377;
  wire n_28378, n_28379, n_28380, n_28381, n_28383, n_28384, n_28385,
       n_28386;
  wire n_28387, n_28388, n_28389, n_28390, n_28391, n_28392, n_28393,
       n_28394;
  wire n_28395, n_28396, n_28397, n_28398, n_28399, n_28400, n_28401,
       n_28402;
  wire n_28403, n_28404, n_28405, n_28406, n_28407, n_28408, n_28409,
       n_28410;
  wire n_28411, n_28412, n_28413, n_28414, n_28415, n_28416, n_28417,
       n_28418;
  wire n_28419, n_28420, n_28421, n_28422, n_28423, n_28424, n_28425,
       n_28426;
  wire n_28427, n_28428, n_28429, n_28430, n_28431, n_28432, n_28433,
       n_28434;
  wire n_28435, n_28436, n_28437, n_28438, n_28439, n_28440, n_28441,
       n_28442;
  wire n_28443, n_28444, n_28445, n_28446, n_28447, n_28448, n_28449,
       n_28450;
  wire n_28451, n_28452, n_28453, n_28454, n_28455, n_28456, n_28457,
       n_28458;
  wire n_28459, n_28460, n_28461, n_28462, n_28463, n_28464, n_28465,
       n_28466;
  wire n_28467, n_28468, n_28469, n_28470, n_28471, n_28472, n_28473,
       n_28474;
  wire n_28475, n_28476, n_28477, n_28478, n_28479, n_28480, n_28481,
       n_28482;
  wire n_28483, n_28484, n_28485, n_28487, n_28488, n_28489, n_28490,
       n_28491;
  wire n_28492, n_28493, n_28494, n_28495, n_28496, n_28497, n_28498,
       n_28499;
  wire n_28500, n_28501, n_28502, n_28503, n_28504, n_28505, n_28506,
       n_28507;
  wire n_28508, n_28510, n_28511, n_28512, n_28513, n_28514, n_28515,
       n_28516;
  wire n_28517, n_28518, n_28519, n_28520, n_28521, n_28522, n_28523,
       n_28524;
  wire n_28525, n_28526, n_28527, n_28528, n_28529, n_28530, n_28531,
       n_28532;
  wire n_28533, n_28534, n_28535, n_28536, n_28537, n_28538, n_28539,
       n_28540;
  wire n_28541, n_28542, n_28543, n_28544, n_28545, n_28546, n_28547,
       n_28548;
  wire n_28549, n_28550, n_28551, n_28552, n_28553, n_28554, n_28555,
       n_28556;
  wire n_28557, n_28558, n_28559, n_28560, n_28561, n_28562, n_28563,
       n_28564;
  wire n_28565, n_28566, n_28567, n_28568, n_28569, n_28570, n_28571,
       n_28572;
  wire n_28573, n_28574, n_28575, n_28576, n_28577, n_28578, n_28579,
       n_28580;
  wire n_28581, n_28582, n_28583, n_28584, n_28585, n_28586, n_28587,
       n_28588;
  wire n_28589, n_28590, n_28591, n_28592, n_28593, n_28594, n_28595,
       n_28596;
  wire n_28597, n_28598, n_28599, n_28600, n_28601, n_28602, n_28603,
       n_28604;
  wire n_28605, n_28606, n_28607, n_28608, n_28609, n_28610, n_28611,
       n_28612;
  wire n_28613, n_28614, n_28615, n_28616, n_28617, n_28618, n_28619,
       n_28620;
  wire n_28621, n_28622, n_28623, n_28624, n_28625, n_28626, n_28627,
       n_28628;
  wire n_28629, n_28630, n_28631, n_28632, n_28633, n_28634, n_28635,
       n_28636;
  wire n_28637, n_28638, n_28639, n_28640, n_28641, n_28642, n_28643,
       n_28644;
  wire n_28645, n_28646, n_28647, n_28648, n_28649, n_28650, n_28651,
       n_28652;
  wire n_28653, n_28654, n_28655, n_28656, n_28657, n_28658, n_28659,
       n_28660;
  wire n_28661, n_28662, n_28663, n_28664, n_28665, n_28666, n_28667,
       n_28668;
  wire n_28669, n_28670, n_28671, n_28672, n_28673, n_28674, n_28675,
       n_28676;
  wire n_28677, n_28678, n_28679, n_28680, n_28681, n_28682, n_28683,
       n_28684;
  wire n_28685, n_28686, n_28687, n_28688, n_28689, n_28690, n_28691,
       n_28692;
  wire n_28693, n_28694, n_28695, n_28696, n_28697, n_28698, n_28699,
       n_28700;
  wire n_28701, n_28702, n_28703, n_28704, n_28705, n_28706, n_28707,
       n_28708;
  wire n_28709, n_28710, n_28711, n_28712, n_28713, n_28714, n_28715,
       n_28716;
  wire n_28717, n_28718, n_28719, n_28720, n_28721, n_28722, n_28723,
       n_28724;
  wire n_28725, n_28726, n_28727, n_28728, n_28729, n_28730, n_28731,
       n_28732;
  wire n_28733, n_28734, n_28735, n_28741, n_28742, n_28743, n_28744,
       n_28745;
  wire n_28746, n_28747, n_28748, n_28749, n_28750, n_28751, n_28752,
       n_28753;
  wire n_28754, n_28755, n_28756, n_28757, n_28758, n_28759, n_28760,
       n_28761;
  wire n_28762, n_28763, n_28764, n_28765, n_28766, n_28767, n_28768,
       n_28769;
  wire n_28770, n_28771, n_28772, n_28773, n_28774, n_28775, n_28776,
       n_28777;
  wire n_28778, n_28779, n_28780, n_28781, n_28782, n_28783, n_28784,
       n_28785;
  wire n_28786, n_28787, n_28788, n_28789, n_28790, n_28791, n_28792,
       n_28793;
  wire n_28794, n_28795, n_28796, n_28797, n_28798, n_28799, n_28800,
       n_28801;
  wire n_28802, n_28803, n_28804, n_28805, n_28806, n_28807, n_28808,
       n_28809;
  wire n_28810, n_28811, n_28812, n_28813, n_28814, n_28815, n_28816,
       n_28817;
  wire n_28818, n_28819, n_28820, n_28821, n_28822, n_28823, n_28824,
       n_28825;
  wire n_28826, n_28827, n_28828, n_28829, n_28830, n_28831, n_28832,
       n_28833;
  wire n_28834, n_28835, n_28836, n_28837, n_28838, n_28839, n_28840,
       n_28841;
  wire n_28842, n_28843, n_28844, n_28845, n_28846, n_28847, n_28848,
       n_28849;
  wire n_28850, n_28851, n_28852, n_28853, n_28854, n_28855, n_28856,
       n_28857;
  wire n_28858, n_28859, n_28860, n_28861, n_28862, n_28863, n_28864,
       n_28865;
  wire n_28866, n_28867, n_28868, n_28869, n_28870, n_28871, n_28873,
       n_28874;
  wire n_28875, n_28876, n_28877, n_28878, n_28879, n_28880, n_28881,
       n_28882;
  wire n_28883, n_28884, n_28885, n_28886, n_28887, n_28888, n_28889,
       n_28890;
  wire n_28891, n_28892, n_28893, n_28894, n_28895, n_28896, n_28897,
       n_28898;
  wire n_28899, n_28900, n_28901, n_28902, n_28903, n_28904, n_28905,
       n_28906;
  wire n_28907, n_28908, n_28909, n_28910, n_28911, n_28912, n_28913,
       n_28914;
  wire n_28915, n_28916, n_28917, n_28918, n_28919, n_28920, n_28921,
       n_28922;
  wire n_28923, n_28924, n_28925, n_28926, n_28927, n_28928, n_28929,
       n_28930;
  wire n_28931, n_28932, n_28933, n_28934, n_28935, n_28936, n_28937,
       n_28938;
  wire n_28939, n_28940, n_28941, n_28942, n_28943, n_28944, n_28945,
       n_28946;
  wire n_28947, n_28948, n_28949, n_28950, n_28951, n_28952, n_28953,
       n_28954;
  wire n_28955, n_28956, n_28957, n_28958, n_28959, n_28960, n_28961,
       n_28962;
  wire n_28963, n_28964, n_28965, n_28966, n_28967, n_28968, n_28969,
       n_28970;
  wire n_28971, n_28972, n_28973, n_28974, n_28975, n_28976, n_28977,
       n_28978;
  wire n_28979, n_28980, n_28981, n_28982, n_28983, n_28984, n_28985,
       n_28986;
  wire n_28987, n_28988, n_28989, n_28990, n_28991, n_28992, n_28993,
       n_28994;
  wire n_28995, n_28996, n_28997, n_28998, n_28999, n_29000, n_29001,
       n_29002;
  wire n_29003, n_29004, n_29005, n_29006, n_29007, n_29008, n_29009,
       n_29010;
  wire n_29011, n_29012, n_29013, n_29014, n_29015, n_29016, n_29017,
       n_29018;
  wire n_29019, n_29020, n_29021, n_29022, n_29023, n_29024, n_29025,
       n_29026;
  wire n_29027, n_29028, n_29029, n_29030, n_29031, n_29032, n_29033,
       n_29034;
  wire n_29035, n_29036, n_29037, n_29038, n_29039, n_29040, n_29041,
       n_29042;
  wire n_29043, n_29044, n_29045, n_29046, n_29047, n_29048, n_29049,
       n_29050;
  wire n_29051, n_29052, n_29053, n_29054, n_29055, n_29056, n_29057,
       n_29058;
  wire n_29059, n_29060, n_29061, n_29062, n_29066, n_29067, n_29068,
       n_29069;
  wire n_29070, n_29071, n_29072, n_29073, n_29074, n_29075, n_29076,
       n_29077;
  wire n_29078, n_29079, n_29081, n_29082, n_29083, n_29084, n_29085,
       n_29086;
  wire n_29087, n_29088, n_29089, n_29090, n_29092, n_29093, n_29094,
       n_29095;
  wire n_29096, n_29097, n_29098, n_29099, n_29100, n_29101, n_29102,
       n_29103;
  wire n_29104, n_29105, n_29106, n_29107, n_29108, n_29109, n_29110,
       n_29111;
  wire n_29112, n_29113, n_29114, n_29115, n_29116, n_29117, n_29118,
       n_29119;
  wire n_29120, n_29121, n_29122, n_29123, n_29124, n_29125, n_29126,
       n_29127;
  wire n_29128, n_29129, n_29130, n_29131, n_29132, n_29133, n_29134,
       n_29135;
  wire n_29136, n_29137, n_29138, n_29139, n_29140, n_29141, n_29142,
       n_29143;
  wire n_29144, n_29145, n_29146, n_29147, n_29148, n_29149, n_29150,
       n_29151;
  wire n_29152, n_29153, n_29154, n_29155, n_29156, n_29157, n_29158,
       n_29159;
  wire n_29160, n_29161, n_29162, n_29163, n_29164, n_29165, n_29166,
       n_29167;
  wire n_29168, n_29169, n_29170, n_29171, n_29172, n_29173, n_29174,
       n_29175;
  wire n_29176, n_29177, n_29178, n_29179, n_29180, n_29181, n_29182,
       n_29183;
  wire n_29184, n_29185, n_29186, n_29187, n_29188, n_29189, n_29190,
       n_29191;
  wire n_29192, n_29193, n_29194, n_29195, n_29196, n_29197, n_29198,
       n_29199;
  wire n_29200, n_29201, n_29202, n_29203, n_29204, n_29205, n_29206,
       n_29207;
  wire n_29208, n_29209, n_29210, n_29211, n_29212, n_29213, n_29214,
       n_29215;
  wire n_29216, n_29217, n_29218, n_29219, n_29220, n_29221, n_29222,
       n_29223;
  wire n_29224, n_29225, n_29226, n_29227, n_29228, n_29229, n_29230,
       n_29231;
  wire n_29232, n_29233, n_29234, n_29235, n_29236, n_29237, n_29238,
       n_29239;
  wire n_29240, n_29241, n_29242, n_29243, n_29244, n_29245, n_29246,
       n_29247;
  wire n_29248, n_29249, n_29250, n_29251, n_29252, n_29253, n_29254,
       n_29255;
  wire n_29256, n_29257, n_29258, n_29259, n_29260, n_29261, n_29262,
       n_29263;
  wire n_29264, n_29265, n_29266, n_29267, n_29268, n_29269, n_29270,
       n_29271;
  wire n_29272, n_29273, n_29274, n_29275, n_29276, n_29277, n_29278,
       n_29279;
  wire n_29280, n_29281, n_29282, n_29283, n_29284, n_29285, n_29286,
       n_29287;
  wire n_29288, n_29289, n_29290, n_29291, n_29292, n_29293, n_29294,
       n_29295;
  wire n_29296, n_29297, n_29298, n_29299, n_29300, n_29301, n_29302,
       n_29303;
  wire n_29304, n_29305, n_29306, n_29307, n_29308, n_29309, n_29310,
       n_29311;
  wire n_29312, n_29313, n_29314, n_29315, n_29316, n_29317, n_29318,
       n_29319;
  wire n_29320, n_29321, n_29322, n_29323, n_29324, n_29325, n_29326,
       n_29327;
  wire n_29328, n_29329, n_29330, n_29331, n_29332, n_29333, n_29334,
       n_29335;
  wire n_29336, n_29337, n_29338, n_29339, n_29340, n_29341, n_29342,
       n_29343;
  wire n_29344, n_29345, n_29346, n_29347, n_29348, n_29349, n_29350,
       n_29351;
  wire n_29352, n_29353, n_29354, n_29355, n_29356, n_29357, n_29358,
       n_29359;
  wire n_29360, n_29361, n_29362, n_29363, n_29364, n_29365, n_29366,
       n_29367;
  wire n_29368, n_29369, n_29370, n_29371, n_29372, n_29373, n_29374,
       n_29375;
  wire n_29376, n_29377, n_29378, n_29379, n_29380, n_29381, n_29382,
       n_29383;
  wire n_29384, n_29385, n_29386, n_29387, n_29388, n_29389, n_29390,
       n_29391;
  wire n_29392, n_29393, n_29394, n_29395, n_29396, n_29397, n_29398,
       n_29399;
  wire n_29400, n_29401, n_29402, n_29403, n_29404, n_29405, n_29406,
       n_29407;
  wire n_29408, n_29409, n_29410, n_29411, n_29412, n_29413, n_29414,
       n_29415;
  wire n_29416, n_29417, n_29418, n_29419, n_29420, n_29421, n_29422,
       n_29423;
  wire n_29424, n_29425, n_29426, n_29427, n_29428, n_29429, n_29430,
       n_29431;
  wire n_29432, n_29433, n_29434, n_29435, n_29436, n_29437, n_29438,
       n_29439;
  wire n_29440, n_29441, n_29442, n_29443, n_29444, n_29445, n_29446,
       n_29447;
  wire n_29448, n_29449, n_29450, n_29451, n_29452, n_29453, n_29454,
       n_29455;
  wire n_29456, n_29457, n_29458, n_29459, n_29460, n_29461, n_29462,
       n_29463;
  wire n_29464, n_29465, n_29466, n_29468, n_29469, n_29470, n_29471,
       n_29472;
  wire n_29473, n_29474, n_29475, n_29476, n_29477, n_29478, n_29479,
       n_29480;
  wire n_29481, n_29482, n_29483, n_29484, n_29485, n_29486, n_29487,
       n_29488;
  wire n_29489, n_29490, n_29491, n_29492, n_29493, n_29494, n_29495,
       n_29496;
  wire n_29497, n_29498, n_29499, n_29500, n_29501, n_29502, n_29503,
       n_29504;
  wire n_29505, n_29506, n_29507, n_29508, n_29512, n_29513, n_29514,
       n_29515;
  wire n_29516, n_29517, n_29518, n_29519, n_29520, n_29521, n_29522,
       n_29523;
  wire n_29524, n_29525, n_29526, n_29527, n_29528, n_29529, n_29530,
       n_29531;
  wire n_29532, n_29533, n_29534, n_29535, n_29536, n_29537, n_29538,
       n_29539;
  wire n_29540, n_29541, n_29542, n_29543, n_29544, n_29545, n_29546,
       n_29547;
  wire n_29548, n_29549, n_29550, n_29551, n_29552, n_29553, n_29554,
       n_29555;
  wire n_29556, n_29557, n_29558, n_29559, n_29560, n_29561, n_29562,
       n_29563;
  wire n_29564, n_29565, n_29566, n_29567, n_29571, n_29572, n_29573,
       n_29574;
  wire n_29575, n_29576, n_29577, n_29578, n_29579, n_29580, n_29581,
       n_29582;
  wire n_29583, n_29584, n_29585, n_29586, n_29587, n_29588, n_29589,
       n_29590;
  wire n_29591, n_29592, n_29593, n_29594, n_29595, n_29596, n_29597,
       n_29598;
  wire n_29599, n_29600, n_29604, n_29605, n_29606, n_29607, n_29610,
       n_29611;
  wire n_29612, n_29613, n_29614, n_29615, n_29616, n_29617, n_29618,
       n_29619;
  wire n_29620, n_29623, n_29624, n_29625, n_29626, n_29627, n_29628,
       n_29629;
  wire n_29630, n_29631, n_29632, n_29633, n_29634, n_29635, n_29636,
       n_29637;
  wire n_29638, n_29639, n_29640, n_29641, n_29642, n_29643, n_29644,
       n_29645;
  wire n_29646, n_29647, n_29648, n_29649, n_29650, n_29651, n_29652,
       n_29653;
  wire n_29654, n_29655, n_29656, n_29657, n_29658, n_29659, n_29660,
       n_29661;
  wire n_29662, n_29663, n_29664, n_29665, n_29669, n_29670, n_29671,
       n_29672;
  wire n_29673, n_29674, n_29675, n_29676, n_29677, n_29678, n_29679,
       n_29680;
  wire n_29681, n_29682, n_29683, n_29684, n_29685, n_29686, n_29687,
       n_29688;
  wire n_29689, n_29690, n_29691, n_29692, n_29693, n_29694, n_29695,
       n_29696;
  wire n_29697, n_29698, n_29699, n_29700, n_29701, n_29702, n_29703,
       n_29704;
  wire n_29705, n_29706, n_29707, n_29708, n_29709, n_29710, n_29711,
       n_29712;
  wire n_29713, n_29714, n_29715, n_29716, n_29717, n_29718, n_29719,
       n_29720;
  wire n_29721, n_29722, n_29723, n_29724, n_29725, n_29726, n_29727,
       n_29728;
  wire n_29729, n_29730, n_29731, n_29732, n_29733, n_29734, n_29735,
       n_29736;
  wire n_29737, n_29738, n_29739, n_29740, n_29741, n_29742, n_29743,
       n_29746;
  wire n_29747, n_29748, n_29749, n_29750, n_29751, n_29752, n_29753,
       n_29754;
  wire n_29755, n_29756, n_29757, n_29758, n_29759, n_29760, n_29761,
       n_29762;
  wire n_29768, n_29769, n_29770, n_29771, n_29772, n_29773, n_29774,
       n_29775;
  wire n_29776, n_29777, n_29778, n_29779, n_29780, n_29781, n_29782,
       n_29783;
  wire n_29784, n_29785, n_29786, n_29787, n_29788, n_29789, n_29790,
       n_29791;
  wire n_29792, n_29793, n_29794, n_29795, n_29796, n_29797, n_29798,
       n_29799;
  wire n_29800, n_29801, n_29802, n_29803, n_29804, n_29805, n_29806,
       n_29807;
  wire n_29808, n_29810, n_29811, n_29812, n_29813, n_29814, n_29815,
       n_29817;
  wire n_29818, n_29819, n_29820, n_29821, n_29822, n_29823, n_29824,
       n_29825;
  wire n_29826, n_29827, n_29828, n_29829, n_29830, n_29831, n_29832,
       n_29833;
  wire n_29834, n_29835, n_29836, n_29837, n_29838, n_29839, n_29840,
       n_29841;
  wire n_29842, n_29843, n_29844, n_29845, n_29846, n_29847, n_29848,
       n_29849;
  wire n_29850, n_29851, n_29852, n_29853, n_29854, n_29856, n_29857,
       n_29858;
  wire n_29859, n_29860, n_29861, n_29862, n_29863, n_29864, n_29865,
       n_29866;
  wire n_29867, n_29868, n_29869, n_29870, n_29871, n_29872, n_29873,
       n_29874;
  wire n_29875, n_29876, n_29877, n_29878, n_29879, n_29880, n_29881,
       n_29882;
  wire n_29883, n_29884, n_29885, n_29886, n_29887, n_29888, n_29889,
       n_29890;
  wire n_29891, n_29892, n_29893, n_29894, n_29895, n_29896, n_29897,
       n_29898;
  wire n_29899, n_29900, n_29901, n_29902, n_29903, n_29904, n_29905,
       n_29906;
  wire n_29907, n_29908, n_29909, n_29910, n_29911, n_29912, n_29913,
       n_29914;
  wire n_29915, n_29916, n_29917, n_29918, n_29919, n_29920, n_29921,
       n_29922;
  wire n_29923, n_29924, n_29925, n_29926, n_29927, n_29928, n_29929,
       n_29930;
  wire n_29931, n_29932, n_29933, n_29934, n_29935, n_29936, n_29937,
       n_29938;
  wire n_29939, n_29940, n_29941, n_29942, n_29943, n_29944, n_29945,
       n_29946;
  wire n_29947, n_29948, n_29949, n_29950, n_29951, n_29952, n_29953,
       n_29954;
  wire n_29955, n_29956, n_29957, n_29958, n_29959, n_29960, n_29961,
       n_29962;
  wire n_29963, n_29964, n_29965, n_29966, n_29967, n_29968, n_29969,
       n_29970;
  wire n_29971, n_29972, n_29973, n_29974, n_29975, n_29976, n_29977,
       n_29978;
  wire n_29979, n_29980, n_29981, n_29982, n_29983, n_29984, n_29985,
       n_29986;
  wire n_29987, n_29988, n_29989, n_29990, n_29991, n_29992, n_29993,
       n_29994;
  wire n_29995, n_29996, n_29997, n_29998, n_29999, n_30000, n_30001,
       n_30002;
  wire n_30003, n_30004, n_30005, n_30006, n_30007, n_30008, n_30009,
       n_30010;
  wire n_30011, n_30012, n_30013, n_30014, n_30015, n_30016, n_30017,
       n_30018;
  wire n_30019, n_30020, n_30021, n_30022, n_30023, n_30024, n_30025,
       n_30026;
  wire n_30027, n_30028, n_30029, n_30030, n_30031, n_30032, n_30033,
       n_30034;
  wire n_30035, n_30036, n_30037, n_30038, n_30039, n_30040, n_30041,
       n_30042;
  wire n_30043, n_30044, n_30045, n_30046, n_30047, n_30048, n_30049,
       n_30050;
  wire n_30051, n_30052, n_30053, n_30054, n_30055, n_30056, n_30057,
       n_30058;
  wire n_30059, n_30060, n_30061, n_30062, n_30063, n_30064, n_30065,
       n_30066;
  wire n_30067, n_30068, n_30069, n_30070, n_30071, n_30072, n_30073,
       n_30074;
  wire n_30075, n_30076, n_30077, n_30078, n_30079, n_30080, n_30081,
       n_30082;
  wire n_30083, n_30084, n_30085, n_30086, n_30087, n_30088, n_30089,
       n_30090;
  wire n_30091, n_30092, n_30093, n_30094, n_30095, n_30096, n_30097,
       n_30098;
  wire n_30099, n_30100, n_30101, n_30102, n_30103, n_30104, n_30105,
       n_30106;
  wire n_30107, n_30108, n_30109, n_30110, n_30111, n_30112, n_30113,
       n_30114;
  wire n_30115, n_30116, n_30117, n_30118, n_30119, n_30120, n_30121,
       n_30122;
  wire n_30123, n_30124, n_30125, n_30126, n_30127, n_30128, n_30129,
       n_30130;
  wire n_30131, n_30133, n_30134, n_30135, n_30136, n_30137, n_30138,
       n_30139;
  wire n_30140, n_30141, n_30142, n_30143, n_30144, n_30145, n_30146,
       n_30147;
  wire n_30148, n_30149, n_30150, n_30151, n_30152, n_30153, n_30154,
       n_30155;
  wire n_30156, n_30157, n_30158, n_30159, n_30160, n_30161, n_30162,
       n_30163;
  wire n_30164, n_30165, n_30166, n_30167, n_30168, n_30169, n_30170,
       n_30171;
  wire n_30172, n_30173, n_30174, n_30175, n_30176, n_30177, n_30178,
       n_30179;
  wire n_30180, n_30181, n_30182, n_30183, n_30184, n_30185, n_30186,
       n_30187;
  wire n_30188, n_30189, n_30190, n_30191, n_30192, n_30193, n_30194,
       n_30195;
  wire n_30196, n_30197, n_30198, n_30199, n_30200, n_30201, n_30202,
       n_30203;
  wire n_30204, n_30205, n_30206, n_30207, n_30208, n_30209, n_30210,
       n_30211;
  wire n_30212, n_30213, n_30214, n_30215, n_30216, n_30217, n_30218,
       n_30219;
  wire n_30220, n_30221, n_30222, n_30223, n_30224, n_30225, n_30226,
       n_30227;
  wire n_30228, n_30229, n_30230, n_30231, n_30232, n_30233, n_30234,
       n_30235;
  wire n_30236, n_30237, n_30238, n_30239, n_30240, n_30241, n_30242,
       n_30243;
  wire n_30244, n_30245, n_30246, n_30247, n_30248, n_30249, n_30250,
       n_30251;
  wire n_30252, n_30253, n_30254, n_30255, n_30256, n_30257, n_30258,
       n_30259;
  wire n_30260, n_30261, n_30262, n_30263, n_30264, n_30265, n_30266,
       n_30267;
  wire n_30268, n_30269, n_30270, n_30271, n_30272, n_30273, n_30274,
       n_30275;
  wire n_30276, n_30277, n_30278, n_30279, n_30280, n_30281, n_30282,
       n_30283;
  wire n_30284, n_30285, n_30286, n_30287, n_30288, n_30289, n_30290,
       n_30291;
  wire n_30292, n_30293, n_30294, n_30295, n_30296, n_30297, n_30298,
       n_30299;
  wire n_30300, n_30301, n_30302, n_30303, n_30304, n_30305, n_30306,
       n_30307;
  wire n_30308, n_30309, n_30310, n_30311, n_30312, n_30313, n_30314,
       n_30315;
  wire n_30316, n_30317, n_30318, n_30319, n_30320, n_30321, n_30322,
       n_30323;
  wire n_30324, n_30325, n_30326, n_30327, n_30328, n_30329, n_30330,
       n_30331;
  wire n_30332, n_30333, n_30334, n_30335, n_30336, n_30337, n_30338,
       n_30339;
  wire n_30340, n_30341, n_30342, n_30343, n_30344, n_30345, n_30346,
       n_30347;
  wire n_30348, n_30349, n_30350, n_30351, n_30352, n_30353, n_30354,
       n_30355;
  wire n_30356, n_30357, n_30358, n_30359, n_30360, n_30361, n_30362,
       n_30363;
  wire n_30364, n_30365, n_30366, n_30367, n_30368, n_30369, n_30370,
       n_30371;
  wire n_30372, n_30373, n_30374, n_30375, n_30376, n_30377, n_30378,
       n_30379;
  wire n_30380, n_30381, n_30382, n_30383, n_30384, n_30385, n_30386,
       n_30387;
  wire n_30388, n_30389, n_30390, n_30391, n_30392, n_30393, n_30394,
       n_30395;
  wire n_30396, n_30397, n_30398, n_30399, n_30400, n_30401, n_30402,
       n_30403;
  wire n_30404, n_30405, n_30406, n_30407, n_30408, n_30409, n_30410,
       n_30411;
  wire n_30412, n_30417, n_30418, n_30423, n_30424, n_30425, n_30426,
       n_30427;
  wire n_30428, n_30429, n_30430, n_30431, n_30432, n_30433, n_30434,
       n_30435;
  wire n_30436, n_30440, n_30441, n_30442, n_30443, n_30444, n_30445,
       n_30446;
  wire n_30447, n_30448, n_30449, n_30450, n_30451, n_30452, n_30457,
       n_30458;
  wire n_30459, n_30460, n_30461, n_30462, n_30463, n_30464, n_30465,
       n_30466;
  wire n_30467, n_30468, n_30469, n_30470, n_30471, n_30472, n_30473,
       n_30474;
  wire n_30475, n_30476, n_30477, n_30478, n_30479, n_30480, n_30481,
       n_30482;
  wire n_30483, n_30484, n_30485, n_30486, n_30487, n_30488, n_30489,
       n_30490;
  wire n_30491, n_30492, n_30493, n_30494, n_30495, n_30496, n_30497,
       n_30498;
  wire n_30499, n_30500, n_30501, n_30505, n_30506, n_30507, n_30508,
       n_30509;
  wire n_30510, n_30511, n_30512, n_30513, n_30514, n_30515, n_30516,
       n_30517;
  wire n_30518, n_30519, n_30520, n_30521, n_30522, n_30523, n_30524,
       n_30525;
  wire n_30526, n_30527, n_30528, n_30529, n_30530, n_30531, n_30532,
       n_30533;
  wire n_30534, n_30535, n_30536, n_30537, n_30538, n_30539, n_30540,
       n_30541;
  wire n_30542, n_30543, n_30544, n_30545, n_30546, n_30547, n_30548,
       n_30549;
  wire n_30550, n_30551, n_30552, n_30553, n_30554, n_30555, n_30556,
       n_30557;
  wire n_30558, n_30559, n_30560, n_30561, n_30562, n_30563, n_30564,
       n_30565;
  wire n_30566, n_30567, n_30568, n_30569, n_30570, n_30571, n_30572,
       n_30573;
  wire n_30577, n_30578, n_30579, n_30580, n_30581, n_30582, n_30583,
       n_30584;
  wire n_30585, n_30586, n_30587, n_30588, n_30589, n_30590, n_30591,
       n_30592;
  wire n_30593, n_30594, n_30595, n_30596, n_30597, n_30598, n_30599,
       n_30600;
  wire n_30601, n_30602, n_30603, n_30604, n_30605, n_30606, n_30607,
       n_30608;
  wire n_30609, n_30610, n_30611, n_30612, n_30613, n_30614, n_30615,
       n_30616;
  wire n_30617, n_30618, n_30619, n_30620, n_30621, n_30622, n_30623,
       n_30624;
  wire n_30625, n_30626, n_30627, n_30628, n_30629, n_30630, n_30631,
       n_30632;
  wire n_30633, n_30634, n_30635, n_30636, n_30637, n_30638, n_30639,
       n_30640;
  wire n_30641, n_30642, n_30643, n_30644, n_30645, n_30646, n_30647,
       n_30648;
  wire n_30649, n_30652, n_30653, n_30654, n_30655, n_30656, n_30657,
       n_30658;
  wire n_30659, n_30660, n_30661, n_30662, n_30663, n_30664, n_30665,
       n_30666;
  wire n_30667, n_30668, n_30669, n_30670, n_30671, n_30672, n_30677,
       n_30678;
  wire n_30679, n_30680, n_30681, n_30682, n_30683, n_30687, n_30688,
       n_30689;
  wire n_30690, n_30691, n_30692, n_30693, n_30694, n_30695, n_30696,
       n_30697;
  wire n_30698, n_30699, n_30700, n_30701, n_30702, n_30703, n_30704,
       n_30705;
  wire n_30706, n_30707, n_30708, n_30709, n_30710, n_30711, n_30712,
       n_30713;
  wire n_30714, n_30715, n_30716, n_30717, n_30718, n_30719, n_30720,
       n_30721;
  wire n_30722, n_30723, n_30724, n_30725, n_30726, n_30727, n_30728,
       n_30729;
  wire n_30730, n_30731, n_30732, n_30733, n_30734, n_30735, n_30736,
       n_30737;
  wire n_30738, n_30739, n_30740, n_30741, n_30742, n_30743, n_30744,
       n_30745;
  wire n_30746, n_30747, n_30748, n_30749, n_30750, n_30751, n_30752,
       n_30753;
  wire n_30754, n_30755, n_30756, n_30757, n_30758, n_30759, n_30760,
       n_30761;
  wire n_30762, n_30763, n_30764, n_30765, n_30766, n_30767, n_30768,
       n_30769;
  wire n_30770, n_30771, n_30772, n_30773, n_30774, n_30775, n_30776,
       n_30777;
  wire n_30778, n_30779, n_30780, n_30781, n_30782, n_30783, n_30784,
       n_30785;
  wire n_30786, n_30787, n_30788, n_30789, n_30790, n_30791, n_30792,
       n_30793;
  wire n_30794, n_30795, n_30796, n_30797, n_30798, n_30799, n_30800,
       n_30801;
  wire n_30802, n_30803, n_30804, n_30805, n_30806, n_30807, n_30808,
       n_30809;
  wire n_30810, n_30811, n_30812, n_30813, n_30814, n_30815, n_30816,
       n_30817;
  wire n_30818, n_30819, n_30820, n_30821, n_30822, n_30823, n_30824,
       n_30825;
  wire n_30826, n_30827, n_30828, n_30829, n_30830, n_30831, n_30832,
       n_30833;
  wire n_30834, n_30835, n_30836, n_30837, n_30838, n_30839, n_30840,
       n_30841;
  wire n_30842, n_30843, n_30844, n_30845, n_30846, n_30847, n_30848,
       n_30849;
  wire n_30850, n_30851, n_30852, n_30853, n_30854, n_30855, n_30856,
       n_30859;
  wire n_30860, n_30861, n_30862, n_30863, n_30864, n_30865, n_30866,
       n_30867;
  wire n_30868, n_30869, n_30870, n_30871, n_30872, n_30873, n_30874,
       n_30875;
  wire n_30876, n_30877, n_30878, n_30879, n_30882, n_30883, n_30884,
       n_30885;
  wire n_30886, n_30887, n_30888, n_30889, n_30890, n_30891, n_30892,
       n_30893;
  wire n_30894, n_30895, n_30896, n_30897, n_30898, n_30899, n_30900,
       n_30901;
  wire n_30902, n_30903, n_30904, n_30905, n_30906, n_30907, n_30908,
       n_30909;
  wire n_30910, n_30911, n_30912, n_30913, n_30914, n_30915, n_30916,
       n_30917;
  wire n_30918, n_30919, n_30920, n_30921, n_30922, n_30923, n_30924,
       n_30925;
  wire n_30926, n_30927, n_30928, n_30929, n_30930, n_30931, n_30932,
       n_30933;
  wire n_30934, n_30935, n_30938, n_30939, n_30940, n_30941, n_30942,
       n_30943;
  wire n_30944, n_30945, n_30946, n_30947, n_30948, n_30949, n_30950,
       n_30951;
  wire n_30952, n_30953, n_30954, n_30955, n_30956, n_30957, n_30958,
       n_30959;
  wire n_30960, n_30961, n_30962, n_30963, n_30964, n_30965, n_30966,
       n_30967;
  wire n_30968, n_30970, n_30971, n_30972, n_30973, n_30974, n_30975,
       n_30976;
  wire n_30977, n_30978, n_30979, n_30980, n_30981, n_30982, n_30983,
       n_30984;
  wire n_30985, n_30986, n_30987, n_30988, n_30989, n_30990, n_30991,
       n_30992;
  wire n_30993, n_30994, n_30995, n_30996, n_30997, n_30998, n_30999,
       n_31000;
  wire n_31001, n_31002, n_31003, n_31004, n_31005, n_31006, n_31007,
       n_31008;
  wire n_31009, n_31010, n_31011, n_31012, n_31013, n_31014, n_31015,
       n_31016;
  wire n_31017, n_31018, n_31021, n_31022, n_31023, n_31024, n_31025,
       n_31026;
  wire n_31027, n_31028, n_31029, n_31030, n_31031, n_31032, n_31033,
       n_31034;
  wire n_31035, n_31036, n_31037, n_31038, n_31039, n_31040, n_31041,
       n_31042;
  wire n_31043, n_31044, n_31045, n_31046, n_31047, n_31048, n_31049,
       n_31050;
  wire n_31051, n_31052, n_31053, n_31054, n_31055, n_31056, n_31057,
       n_31058;
  wire n_31059, n_31060, n_31063, n_31064, n_31065, n_31066, n_31067,
       n_31068;
  wire n_31069, n_31072, n_31073, n_31074, n_31075, n_31076, n_31080,
       n_31081;
  wire n_31082, n_31083, n_31084, n_31085, n_31086, n_31087, n_31090,
       n_31091;
  wire n_31092, n_31093, n_31094, n_31095, n_31096, n_31097, n_31098,
       n_31099;
  wire n_31100, n_31101, n_31102, n_31103, n_31104, n_31105, n_31106,
       n_31107;
  wire n_31108, n_31109, n_31110, n_31111, n_31112, n_31113, n_31114,
       n_31115;
  wire n_31116, n_31117, n_31118, n_31119, n_31120, n_31121, n_31122,
       n_31123;
  wire n_31124, n_31125, n_31126, n_31127, n_31128, n_31129, n_31130,
       n_31131;
  wire n_31132, n_31133, n_31134, n_31135, n_31136, n_31137, n_31138,
       n_31139;
  wire n_31140, n_31141, n_31142, n_31143, n_31144, n_31145, n_31146,
       n_31147;
  wire n_31148, n_31149, n_31150, n_31151, n_31152, n_31153, n_31154,
       n_31155;
  wire n_31156, n_31157, n_31158, n_31159, n_31160, n_31161, n_31162,
       n_31163;
  wire n_31164, n_31165, n_31166, n_31167, n_31168, n_31169, n_31170,
       n_31171;
  wire n_31172, n_31173, n_31174, n_31175, n_31176, n_31177, n_31178,
       n_31179;
  wire n_31180, n_31181, n_31182, n_31183, n_31184, n_31185, n_31186,
       n_31187;
  wire n_31188, n_31189, n_31190, n_31191, n_31192, n_31193, n_31194,
       n_31195;
  wire n_31196, n_31197, n_31198, n_31199, n_31200, n_31201, n_31202,
       n_31203;
  wire n_31204, n_31205, n_31206, n_31207, n_31208, n_31209, n_31210,
       n_31211;
  wire n_31212, n_31213, n_31214, n_31215, n_31216, n_31217, n_31218,
       n_31219;
  wire n_31220, n_31221, n_31222, n_31223, n_31224, n_31225, n_31226,
       n_31227;
  wire n_31228, n_31229, n_31230, n_31231, n_31232, n_31233, n_31234,
       n_31235;
  wire n_31236, n_31237, n_31238, n_31239, n_31240, n_31241, n_31242,
       n_31243;
  wire n_31244, n_31245, n_31246, n_31247, n_31248, n_31249, n_31250,
       n_31251;
  wire n_31252, n_31253, n_31254, n_31255, n_31256, n_31257, n_31258,
       n_31259;
  wire n_31260, n_31261, n_31262, n_31263, n_31264, n_31265, n_31266,
       n_31267;
  wire n_31268, n_31269, n_31270, n_31271, n_31272, n_31273, n_31274,
       n_31275;
  wire n_31276, n_31277, n_31278, n_31279, n_31280, n_31281, n_31282,
       n_31283;
  wire n_31284, n_31285, n_31286, n_31287, n_31288, n_31289, n_31290,
       n_31291;
  wire n_31292, n_31293, n_31294, n_31295, n_31296, n_31297, n_31298,
       n_31299;
  wire n_31300, n_31301, n_31302, n_31303, n_31304, n_31305, n_31306,
       n_31307;
  wire n_31308, n_31309, n_31310, n_31311, n_31312, n_31313, n_31314,
       n_31315;
  wire n_31316, n_31317, n_31318, n_31319, n_31320, n_31321, n_31322,
       n_31323;
  wire n_31324, n_31325, n_31326, n_31327, n_31328, n_31329, n_31330,
       n_31331;
  wire n_31332, n_31333, n_31334, n_31335, n_31336, n_31337, n_31338,
       n_31339;
  wire n_31340, n_31341, n_31342, n_31343, n_31344, n_31345, n_31346,
       n_31347;
  wire n_31348, n_31349, n_31350, n_31351, n_31352, n_31353, n_31354,
       n_31355;
  wire n_31356, n_31357, n_31358, n_31359, n_31360, n_31361, n_31362,
       n_31363;
  wire n_31364, n_31365, n_31366, n_31367, n_31368, n_31369, n_31370,
       n_31371;
  wire n_31372, n_31373, n_31374, n_31375, n_31376, n_31377, n_31378,
       n_31379;
  wire n_31380, n_31381, n_31382, n_31383, n_31384, n_31385, n_31387,
       n_31388;
  wire n_31389, n_31390, n_31391, n_31392, n_31393, n_31394, n_31396,
       n_31397;
  wire n_31398, n_31399, n_31400, n_31401, n_31402, n_31403, n_31404,
       n_31405;
  wire n_31406, n_31407, n_31408, n_31409, n_31410, n_31411, n_31412,
       n_31413;
  wire n_31414, n_31415, n_31416, n_31417, n_31420, n_31421, n_31422,
       n_31425;
  wire n_31426, n_31427, n_31428, n_31429, n_31430, n_31431, n_31432,
       n_31433;
  wire n_31434, n_31435, n_31436, n_31437, n_31438, n_31439, n_31440,
       n_31441;
  wire n_31442, n_31443, n_31444, n_31445, n_31446, n_31447, n_31448,
       n_31449;
  wire n_31450, n_31451, n_31452, n_31453, n_31454, n_31455, n_31456,
       n_31457;
  wire n_31458, n_31459, n_31460, n_31461, n_31462, n_31463, n_31464,
       n_31465;
  wire n_31466, n_31467, n_31468, n_31469, n_31470, n_31471, n_31472,
       n_31473;
  wire n_31474, n_31475, n_31476, n_31477, n_31478, n_31479, n_31480,
       n_31481;
  wire n_31482, n_31483, n_31484, n_31485, n_31486, n_31487, n_31488,
       n_31489;
  wire n_31490, n_31491, n_31492, n_31493, n_31494, n_31495, n_31496,
       n_31497;
  wire n_31498, n_31499, n_31500, n_31501, n_31502, n_31503, n_31504,
       n_31505;
  wire n_31506, n_31507, n_31508, n_31509, n_31510, n_31511, n_31512,
       n_31513;
  wire n_31514, n_31515, n_31516, n_31517, n_31518, n_31519, n_31520,
       n_31521;
  wire n_31522, n_31526, n_31527, n_31528, n_31531, n_31532, n_31533,
       n_31534;
  wire n_31536, n_31537, n_31538, n_31539, n_31540, n_31541, n_31542,
       n_31543;
  wire n_31544, n_31545, n_31546, n_31547, n_31548, n_31549, n_31550,
       n_31551;
  wire n_31552, n_31553, n_31554, n_31555, n_31556, n_31557, n_31558,
       n_31559;
  wire n_31560, n_31561, n_31562, n_31563, n_31564, n_31565, n_31566,
       n_31567;
  wire n_31568, n_31569, n_31570, n_31571, n_31572, n_31573, n_31574,
       n_31575;
  wire n_31576, n_31577, n_31579, n_31580, n_31581, n_31582, n_31583,
       n_31584;
  wire n_31585, n_31586, n_31587, n_31588, n_31589, n_31590, n_31591,
       n_31592;
  wire n_31593, n_31594, n_31595, n_31596, n_31597, n_31598, n_31599,
       n_31600;
  wire n_31601, n_31602, n_31603, n_31604, n_31605, n_31606, n_31607,
       n_31610;
  wire n_31611, n_31612, n_31613, n_31614, n_31615, n_31616, n_31617,
       n_31618;
  wire n_31619, n_31620, n_31621, n_31622, n_31623, n_31624, n_31625,
       n_31626;
  wire n_31627, n_31628, n_31629, n_31630, n_31631, n_31632, n_31633,
       n_31634;
  wire n_31635, n_31639, n_31640, n_31641, n_31642, n_31643, n_31644,
       n_31645;
  wire n_31646, n_31647, n_31648, n_31649, n_31650, n_31651, n_31652,
       n_31653;
  wire n_31654, n_31655, n_31656, n_31657, n_31658, n_31659, n_31660,
       n_31661;
  wire n_31662, n_31663, n_31664, n_31665, n_31666, n_31667, n_31668,
       n_31669;
  wire n_31670, n_31671, n_31672, n_31673, n_31674, n_31675, n_31676,
       n_31677;
  wire n_31678, n_31679, n_31680, n_31681, n_31682, n_31683, n_31684,
       n_31685;
  wire n_31686, n_31687, n_31688, n_31689, n_31690, n_31691, n_31692,
       n_31693;
  wire n_31694, n_31695, n_31696, n_31697, n_31698, n_31699, n_31700,
       n_31701;
  wire n_31702, n_31703, n_31704, n_31705, n_31706, n_31707, n_31708,
       n_31709;
  wire n_31710, n_31711, n_31712, n_31713, n_31714, n_31715, n_31716,
       n_31717;
  wire n_31718, n_31719, n_31720, n_31721, n_31722, n_31723, n_31724,
       n_31725;
  wire n_31726, n_31727, n_31728, n_31729, n_31730, n_31731, n_31732,
       n_31733;
  wire n_31734, n_31735, n_31736, n_31737, n_31738, n_31739, n_31740,
       n_31741;
  wire n_31742, n_31743, n_31744, n_31745, n_31746, n_31747, n_31748,
       n_31749;
  wire n_31750, n_31751, n_31752, n_31753, n_31754, n_31755, n_31756,
       n_31757;
  wire n_31758, n_31759, n_31760, n_31761, n_31762, n_31763, n_31764,
       n_31765;
  wire n_31766, n_31767, n_31768, n_31769, n_31770, n_31771, n_31772,
       n_31773;
  wire n_31774, n_31775, n_31776, n_31777, n_31778, n_31779, n_31780,
       n_31781;
  wire n_31782, n_31783, n_31784, n_31785, n_31786, n_31787, n_31788,
       n_31789;
  wire n_31790, n_31791, n_31792, n_31793, n_31794, n_31795, n_31796,
       n_31799;
  wire n_31800, n_31801, n_31802, n_31803, n_31804, n_31805, n_31806,
       n_31807;
  wire n_31808, n_31809, n_31810, n_31811, n_31812, n_31813, n_31814,
       n_31815;
  wire n_31816, n_31817, n_31818, n_31819, n_31820, n_31821, n_31822,
       n_31823;
  wire n_31825, n_31826, n_31828, n_31829, n_31830, n_31831, n_31832,
       n_31833;
  wire n_31834, n_31835, n_31836, n_31837, n_31838, n_31839, n_31840,
       n_31841;
  wire n_31842, n_31843, n_31844, n_31845, n_31846, n_31847, n_31848,
       n_31849;
  wire n_31850, n_31851, n_31852, n_31853, n_31854, n_31855, n_31859,
       n_31860;
  wire n_31861, n_31862, n_31863, n_31864, n_31865, n_31866, n_31867,
       n_31868;
  wire n_31869, n_31870, n_31871, n_31872, n_31873, n_31874, n_31875,
       n_31876;
  wire n_31877, n_31878, n_31879, n_31880, n_31881, n_31882, n_31883,
       n_31884;
  wire n_31885, n_31889, n_31890, n_31891, n_31892, n_31896, n_31897,
       n_31898;
  wire n_31899, n_31900, n_31901, n_31902, n_31903, n_31904, n_31905,
       n_31906;
  wire n_31907, n_31908, n_31909, n_31910, n_31913, n_31914, n_31916,
       n_31917;
  wire n_31918, n_31921, n_31922, n_31924, n_31925, n_31926, n_31929,
       n_31930;
  wire n_31932, n_31933, n_31934, n_31937, n_31938, n_31940, n_31941,
       n_31942;
  wire n_31945, n_31946, n_31948, n_31949, n_31950, n_31953, n_31954,
       n_31955;
  wire n_31959, n_31960, n_31961, n_31963, n_31964, n_31965, n_31967,
       n_31968;
  wire n_31969, n_31970, n_31971, n_31972, n_31973, n_31974, n_31975,
       n_31976;
  wire n_31977, n_31978, n_31979, n_31980, n_31981, n_31982, n_31983,
       n_31984;
  wire n_31985, n_31986, n_31987, n_31988, n_31989, n_31990, n_31991,
       n_31992;
  wire n_31993, n_31994, n_31995, n_31996, n_31997, n_31998, n_31999,
       n_32005;
  wire n_32006, n_32007, n_32008, n_32009, n_32010, n_32011, n_32012,
       n_32013;
  wire n_32014, n_32015, n_32016, n_32017, n_32018, n_32019, n_32020,
       n_32021;
  wire n_32022, n_32023, n_32024, n_32025, n_32026, n_32027, n_32028,
       n_32029;
  wire n_32030, n_32031, n_32032, n_32033, n_32034, n_32035, n_32038,
       n_32039;
  wire n_32040, n_32041, n_32042, n_32043, n_32044, n_32045, n_32046,
       n_32047;
  wire n_32048, n_32049, n_32050, n_32051, n_32052, n_32053, n_32054,
       n_32055;
  wire n_32056, n_32057, n_32058, n_32059, n_32060, n_32061, n_32062,
       n_32063;
  wire n_32064, n_32065, n_32066, n_32067, n_32068, n_32069, n_32070,
       n_32071;
  wire n_32072, n_32073, n_32074, n_32075, n_32076, n_32077, n_32078,
       n_32079;
  wire n_32080, n_32081, n_32082, n_32083, n_32084, n_32085, n_32086,
       n_32087;
  wire n_32088, n_32089, n_32090, n_32091, n_32092, n_32093, n_32097,
       n_32098;
  wire n_32099, n_32100, n_32101, n_32102, n_32103, n_32104, n_32105,
       n_32106;
  wire n_32107, n_32108, n_32112, n_32113, n_32114, n_32115, n_32116,
       n_32117;
  wire n_32118, n_32119, n_32120, n_32121, n_32122, n_32123, n_32124,
       n_32125;
  wire n_32126, n_32127, n_32128, n_32129, n_32130, n_32131, n_32132,
       n_32133;
  wire n_32134, n_32135, n_32136, n_32137, n_32138, n_32139, n_32140,
       n_32141;
  wire n_32142, n_32143, n_32144, n_32145, n_32146, n_32147, n_32148,
       n_32149;
  wire n_32150, n_32151, n_32152, n_32153, n_32155, n_32156, n_32157,
       n_32158;
  wire n_32159, n_32160, n_32161, n_32162, n_32163, n_32164, n_32165,
       n_32166;
  wire n_32167, n_32168, n_32169, n_32170, n_32171, n_32172, n_32173,
       n_32174;
  wire n_32175, n_32176, n_32177, n_32178, n_32179, n_32180, n_32181,
       n_32182;
  wire n_32183, n_32184, n_32185, n_32186, n_32187, n_32188, n_32189,
       n_32190;
  wire n_32192, n_32193, n_32194, n_32195, n_32196, n_32197, n_32198,
       n_32199;
  wire n_32200, n_32201, n_32202, n_32203, n_32204, n_32205, n_32206,
       n_32207;
  wire n_32208, n_32209, n_32210, n_32211, n_32212, n_32213, n_32214,
       n_32215;
  wire n_32216, n_32217, n_32218, n_32219, n_32220, n_32221, n_32222,
       n_32223;
  wire n_32224, n_32225, n_32226, n_32227, n_32228, n_32229, n_32230,
       n_32231;
  wire n_32232, n_32233, n_32235, n_32236, n_32237, n_32238, n_32239,
       n_32240;
  wire n_32241, n_32242, n_32243, n_32244, n_32245, n_32246, n_32247,
       n_32248;
  wire n_32249, n_32250, n_32251, n_32252, n_32253, n_32254, n_32255,
       n_32256;
  wire n_32257, n_32258, n_32259, n_32260, n_32261, n_32262, n_32263,
       n_32264;
  wire n_32265, n_32266, n_32267, n_32268, n_32269, n_32270, n_32271,
       n_32272;
  wire n_32273, n_32274, n_32275, n_32276, n_32277, n_32278, n_32279,
       n_32280;
  wire n_32281, n_32282, n_32283, n_32284, n_32285, n_32286, n_32287,
       n_32288;
  wire n_32289, n_32290, n_32291, n_32292, n_32293, n_32294, n_32295,
       n_32296;
  wire n_32297, n_32298, n_32299, n_32300, n_32301, n_32302, n_32303,
       n_32304;
  wire n_32305, n_32306, n_32307, n_32308, n_32309, n_32310, n_32311,
       n_32312;
  wire n_32313, n_32314, n_32315, n_32316, n_32317, n_32318, n_32319,
       n_32320;
  wire n_32321, n_32322, n_32323, n_32324, n_32325, n_32326, n_32327,
       n_32328;
  wire n_32329, n_32330, n_32331, n_32332, n_32333, n_32334, n_32335,
       n_32336;
  wire n_32337, n_32338, n_32339, n_32340, n_32341, n_32342, n_32343,
       n_32344;
  wire n_32345, n_32346, n_32350, n_32351, n_32352, n_32353, n_32354,
       n_32355;
  wire n_32356, n_32357, n_32358, n_32359, n_32360, n_32361, n_32362,
       n_32363;
  wire n_32364, n_32365, n_32366, n_32367, n_32368, n_32369, n_32370,
       n_32371;
  wire n_32372, n_32373, n_32374, n_32375, n_32376, n_32378, n_32379,
       n_32380;
  wire n_32381, n_32382, n_32383, n_32384, n_32385, n_32386, n_32387,
       n_32388;
  wire n_32389, n_32390, n_32391, n_32392, n_32393, n_32394, n_32395,
       n_32396;
  wire n_32397, n_32398, n_32399, n_32400, n_32401, n_32402, n_32403,
       n_32404;
  wire n_32405, n_32406, n_32407, n_32408, n_32409, n_32410, n_32411,
       n_32412;
  wire n_32413, n_32414, n_32415, n_32416, n_32417, n_32418, n_32419,
       n_32420;
  wire n_32421, n_32422, n_32423, n_32424, n_32425, n_32426, n_32427,
       n_32428;
  wire n_32429, n_32430, n_32431, n_32432, n_32433, n_32434, n_32435,
       n_32436;
  wire n_32437, n_32438, n_32439, n_32440, n_32441, n_32442, n_32443,
       n_32444;
  wire n_32448, n_32449, n_32450, n_32451, n_32452, n_32453, n_32454,
       n_32455;
  wire n_32456, n_32457, n_32458, n_32459, n_32460, n_32461, n_32462,
       n_32463;
  wire n_32464, n_32465, n_32466, n_32467, n_32468, n_32469, n_32470,
       n_32471;
  wire n_32472, n_32473, n_32474, n_32475, n_32476, n_32477, n_32478,
       n_32479;
  wire n_32480, n_32481, n_32482, n_32483, n_32484, n_32485, n_32486,
       n_32487;
  wire n_32488, n_32489, n_32490, n_32491, n_32492, n_32493, n_32494,
       n_32495;
  wire n_32496, n_32497, n_32498, n_32499, n_32500, n_32501, n_32502,
       n_32503;
  wire n_32504, n_32505, n_32506, n_32507, n_32508, n_32509, n_32510,
       n_32511;
  wire n_32512, n_32513, n_32514, n_32515, n_32516, n_32517, n_32518,
       n_32519;
  wire n_32520, n_32521, n_32522, n_32523, n_32524, n_32525, n_32526,
       n_32527;
  wire n_32528, n_32529, n_32530, n_32531, n_32532, n_32533, n_32534,
       n_32535;
  wire n_32536, n_32537, n_32538, n_32539, n_32540, n_32541, n_32542,
       n_32543;
  wire n_32544, n_32545, n_32546, n_32547, n_32548, n_32549, n_32550,
       n_32551;
  wire n_32552, n_32553, n_32554, n_32555, n_32556, n_32557, n_32558,
       n_32559;
  wire n_32560, n_32561, n_32562, n_32563, n_32564, n_32565, n_32566,
       n_32567;
  wire n_32568, n_32569, n_32570, n_32571, n_32572, n_32573, n_32574,
       n_32575;
  wire n_32577, n_32578, n_32579, n_32580, n_32581, n_32582, n_32583,
       n_32584;
  wire n_32585, n_32586, n_32587, n_32588, n_32589, n_32590, n_32591,
       n_32592;
  wire n_32593, n_32594, n_32596, n_32597, n_32598, n_32599, n_32600,
       n_32601;
  wire n_32602, n_32603, n_32604, n_32605, n_32606, n_32607, n_32608,
       n_32609;
  wire n_32610, n_32611, n_32612, n_32613, n_32614, n_32615, n_32616,
       n_32617;
  wire n_32618, n_32619, n_32620, n_32621, n_32622, n_32623, n_32624,
       n_32625;
  wire n_32626, n_32627, n_32628, n_32629, n_32630, n_32631, n_32632,
       n_32633;
  wire n_32634, n_32635, n_32636, n_32637, n_32638, n_32639, n_32640,
       n_32641;
  wire n_32642, n_32643, n_32644, n_32645, n_32646, n_32647, n_32648,
       n_32649;
  wire n_32650, n_32651, n_32652, n_32653, n_32654, n_32655, n_32656,
       n_32657;
  wire n_32658, n_32659, n_32660, n_32661, n_32662, n_32663, n_32664,
       n_32665;
  wire n_32666, n_32667, n_32668, n_32669, n_32670, n_32671, n_32672,
       n_32673;
  wire n_32674, n_32675, n_32676, n_32677, n_32678, n_32679, n_32680,
       n_32681;
  wire n_32682, n_32683, n_32684, n_32685, n_32686, n_32687, n_32688,
       n_32689;
  wire n_32690, n_32691, n_32692, n_32693, n_32694, n_32695, n_32696,
       n_32697;
  wire n_32698, n_32699, n_32700, n_32701, n_32702, n_32703, n_32704,
       n_32705;
  wire n_32706, n_32707, n_32708, n_32709, n_32710, n_32711, n_32712,
       n_32713;
  wire n_32714, n_32715, n_32716, n_32717, n_32718, n_32719, n_32720,
       n_32721;
  wire n_32722, n_32723, n_32724, n_32725, n_32726, n_32727, n_32728,
       n_32729;
  wire n_32730, n_32731, n_32732, n_32733, n_32734, n_32735, n_32736,
       n_32737;
  wire n_32738, n_32739, n_32740, n_32741, n_32742, n_32743, n_32744,
       n_32745;
  wire n_32746, n_32747, n_32748, n_32749, n_32750, n_32751, n_32752,
       n_32753;
  wire n_32754, n_32755, n_32756, n_32757, n_32758, n_32759, n_32760,
       n_32761;
  wire n_32762, n_32763, n_32764, n_32765, n_32766, n_32767, n_32768,
       n_32769;
  wire n_32770, n_32771, n_32772, n_32773, n_32774, n_32775, n_32776,
       n_32777;
  wire n_32778, n_32779, n_32780, n_32781, n_32782, n_32783, n_32784,
       n_32785;
  wire n_32786, n_32787, n_32788, n_32789, n_32790, n_32791, n_32792,
       n_32793;
  wire n_32794, n_32795, n_32796, n_32797, n_32798, n_32799, n_32800,
       n_32801;
  wire n_32802, n_32803, n_32804, n_32805, n_32806, n_32807, n_32809,
       n_32810;
  wire n_32811, n_32812, n_32813, n_32814, n_32815, n_32816, n_32817,
       n_32818;
  wire n_32819, n_32820, n_32821, n_32822, n_32823, n_32824, n_32825,
       n_32826;
  wire n_32827, n_32828, n_32829, n_32830, n_32831, n_32832, n_32833,
       n_32834;
  wire n_32835, n_32836, n_32837, n_32838, n_32839, n_32840, n_32841,
       n_32842;
  wire n_32843, n_32844, n_32845, n_32846, n_32847, n_32848, n_32849,
       n_32850;
  wire n_32851, n_32852, n_32853, n_32854, n_32855, n_32856, n_32857,
       n_32858;
  wire n_32859, n_32860, n_32861, n_32862, n_32863, n_32864, n_32865,
       n_32866;
  wire n_32867, n_32868, n_32869, n_32870, n_32871, n_32872, n_32873,
       n_32874;
  wire n_32875, n_32876, n_32877, n_32878, n_32879, n_32880, n_32881,
       n_32882;
  wire n_32883, n_32884, n_32885, n_32886, n_32887, n_32888, n_32889,
       n_32890;
  wire n_32891, n_32892, n_32893, n_32894, n_32895, n_32896, n_32897,
       n_32898;
  wire n_32899, n_32900, n_32901, n_32902, n_32903, n_32904, n_32905,
       n_32906;
  wire n_32907, n_32908, n_32909, n_32910, n_32911, n_32912, n_32913,
       n_32914;
  wire n_32915, n_32917, n_32918, n_32919, n_32920, n_32921, n_32922,
       n_32923;
  wire n_32924, n_32925, n_32926, n_32927, n_32928, n_32929, n_32930,
       n_32931;
  wire n_32932, n_32933, n_32934, n_32935, n_32936, n_32937, n_32938,
       n_32939;
  wire n_32940, n_32941, n_32942, n_32943, n_32944, n_32945, n_32946,
       n_32947;
  wire n_32948, n_32949, n_32952, n_32953, n_32954, n_32955, n_32957,
       n_32958;
  wire n_32959, n_32960, n_32961, n_32962, n_32963, n_32964, n_32965,
       n_32967;
  wire n_32968, n_32969, n_32970, n_32971, n_32972, n_32973, n_32974,
       n_32975;
  wire n_32976, n_32977, n_32978, n_32979, n_32980, n_32981, n_32982,
       n_32983;
  wire n_32984, n_32985, n_32986, n_32987, n_32988, n_32989, n_32990,
       n_32991;
  wire n_32992, n_32993, n_32994, n_32995, n_32996, n_32997, n_32998,
       n_32999;
  wire n_33000, n_33001, n_33002, n_33003, n_33004, n_33005, n_33006,
       n_33007;
  wire n_33008, n_33009, n_33010, n_33011, n_33012, n_33013, n_33014,
       n_33016;
  wire n_33017, n_33018, n_33019, n_33020, n_33021, n_33022, n_33023,
       n_33024;
  wire n_33025, n_33026, n_33027, n_33028, n_33029, n_33030, n_33031,
       n_33032;
  wire n_33033, n_33034, n_33035, n_33036, n_33037, n_33038, n_33039,
       n_33040;
  wire n_33041, n_33042, n_33043, n_33044, n_33045, n_33046, n_33047,
       n_33048;
  wire n_33049, n_33050, n_33051, n_33052, n_33053, n_33054, n_33055,
       n_33056;
  wire n_33057, n_33058, n_33059, n_33060, n_33061, n_33062, n_33063,
       n_33064;
  wire n_33065, n_33066, n_33067, n_33069, n_33070, n_33071, n_33072,
       n_33073;
  wire n_33074, n_33075, n_33076, n_33077, n_33078, n_33079, n_33080,
       n_33081;
  wire n_33082, n_33083, n_33084, n_33085, n_33086, n_33087, n_33088,
       n_33089;
  wire n_33090, n_33091, n_33092, n_33093, n_33094, n_33095, n_33096,
       n_33097;
  wire n_33098, n_33099, n_33100, n_33101, n_33102, n_33103, n_33104,
       n_33105;
  wire n_33106, n_33107, n_33108, n_33109, n_33110, n_33111, n_33112,
       n_33114;
  wire n_33115, n_33116, n_33117, n_33118, n_33119, n_33120, n_33121,
       n_33122;
  wire n_33123, n_33124, n_33125, n_33126, n_33127, n_33128, n_33129,
       n_33130;
  wire n_33131, n_33132, n_33133, n_33134, n_33135, n_33136, n_33137,
       n_33138;
  wire n_33139, n_33140, n_33141, n_33142, n_33143, n_33144, n_33145,
       n_33146;
  wire n_33148, n_33149, n_33150, n_33151, n_33152, n_33153, n_33154,
       n_33155;
  wire n_33156, n_33157, n_33158, n_33159, n_33160, n_33161, n_33162,
       n_33163;
  wire n_33164, n_33165, n_33166, n_33167, n_33168, n_33169, n_33170,
       n_33171;
  wire n_33172, n_33173, n_33174, n_33175, n_33176, n_33177, n_33178,
       n_33179;
  wire n_33180, n_33181, n_33182, n_33183, n_33184, n_33185, n_33186,
       n_33187;
  wire n_33188, n_33189, n_33190, n_33191, n_33192, n_33193, n_33194,
       n_33195;
  wire n_33196, n_33197, n_33198, n_33199, n_33200, n_33201, n_33202,
       n_33203;
  wire n_33204, n_33205, n_33206, n_33207, n_33208, n_33209, n_33210,
       n_33211;
  wire n_33212, n_33213, n_33214, n_33215, n_33216, n_33217, n_33218,
       n_33220;
  wire n_33221, n_33222, n_33223, n_33224, n_33225, n_33226, n_33227,
       n_33228;
  wire n_33229, n_33230, n_33231, n_33232, n_33233, n_33234, n_33235,
       n_33236;
  wire n_33237, n_33239, n_33240, n_33241, n_33243, n_33244, n_33245,
       n_33246;
  wire n_33247, n_33248, n_33249, n_33250, n_33251, n_33252, n_33253,
       n_33254;
  wire n_33255, n_33257, n_33258, n_33259, n_33260, n_33262, n_33263,
       n_33264;
  wire n_33265, n_33267, n_33268, n_33269, n_33270, n_33272, n_33273,
       n_33274;
  wire n_33275, n_33277, n_33278, n_33279, n_33280, n_33282, n_33283,
       n_33284;
  wire n_33285, n_33287, n_33288, n_33289, n_33290, n_33292, n_33293,
       n_33294;
  wire n_33295, n_33297, n_33299, n_33300, n_33301, n_33302, n_33303,
       n_33305;
  wire n_33307, n_33308, n_33309, n_33310, n_33312, n_33314, n_33315,
       n_33316;
  wire n_33317, n_33318, n_33319, n_33320, n_33321, n_33322, n_33323,
       n_33324;
  wire n_33325, n_33338, n_33339, n_33340, n_33341, n_33342, n_33343,
       n_33344;
  wire n_33345, n_33346, n_33347, n_33348, n_33349, n_33350, n_33353,
       n_33354;
  wire n_33355, n_33356, n_33357, n_33358, n_33359, n_33361, n_33362,
       n_33363;
  wire n_33364, n_33365, n_33366, n_33367, n_33368, n_33369, n_33370,
       n_33371;
  wire n_33372, n_33373, n_33376, n_33377, n_33378, n_33379, n_33380,
       n_33381;
  wire n_33382, n_33383, n_33384, n_33385, n_33387, n_33388, n_33392,
       n_33393;
  wire n_33396, n_33397, n_33405, n_33406, n_33407, n_33409, n_33410,
       n_33411;
  wire n_33412, n_33413, n_33414, n_33415, n_33416, n_33417, n_33418,
       n_33419;
  wire n_33420, n_33421, n_33422, n_33423, n_33424, n_33425, n_33426,
       n_33427;
  wire n_33428, n_33429, n_33440, n_33447, n_33448, n_33450, n_33452,
       n_33454;
  wire n_33455, n_33457, n_33458, n_33459, n_33460, n_33461, n_33462,
       n_33463;
  wire n_33464, n_33465, n_33466, n_33467, n_33468, n_33470, n_33472,
       n_33473;
  wire n_33475, n_33476, n_33477, n_33478, n_33479, n_33480, n_33481,
       n_33482;
  wire n_33483, n_33484, n_33485, n_33487, n_33488, n_33489, n_33490,
       n_33491;
  wire n_33492, n_33493, n_33494, n_33495, n_33496, n_33497, n_33501,
       n_33502;
  wire n_33503, n_33504, n_33505, n_33507, n_33508, n_33509, n_33510,
       n_33511;
  wire n_33512, n_33513, n_33514, n_33515, n_33516, n_33521, n_33522,
       n_33523;
  wire n_33525, n_33526, n_33527, n_33528, n_33529, n_33530, n_33531,
       n_33532;
  wire n_33533, n_33534, n_33535, n_33536, n_33537, n_33538, n_33539,
       n_33540;
  wire n_33541, n_33542, n_33543, n_33544, n_33545, n_33546, n_33547,
       n_33549;
  wire n_33550, n_33551, n_33552, n_33553, n_33554, n_33558, n_33559,
       n_33560;
  wire n_33561, n_33563, n_33564, n_33565, n_33566, n_33567, n_33568,
       n_33572;
  wire n_33573, n_33574, n_33575, n_33577, n_33578, n_33579, n_33580,
       n_33581;
  wire n_33582, n_33586, n_33587, n_33588, n_33589, n_33591, n_33592,
       n_33593;
  wire n_33594, n_33595, n_33596, n_33600, n_33601, n_33603, n_33604,
       n_33605;
  wire n_33606, n_33612, n_33613, n_33614, n_33615, n_33621, n_33622,
       n_33623;
  wire n_33624, n_33629, n_33630, n_33632, n_33633, n_33634, n_33643,
       n_33644;
  wire n_33651, n_33652, n_33656, n_33657, n_33665, n_33666, n_33668,
       n_33669;
  wire n_33675, n_33676, n_33685, n_33686, n_33688, n_33689, n_33694,
       n_33695;
  wire n_33697, n_33698, n_33709, n_33710, n_33721, n_33722, n_33729,
       n_33730;
  wire n_33738, n_33739, n_33749, n_33750, n_33751, n_33752, n_33753,
       n_33754;
  wire n_33755, n_33756, n_33757, n_33758, n_33759, n_33760, n_33761,
       n_33762;
  wire n_33763, n_33764, n_33765, n_33766, n_33767, n_33768, n_33769,
       n_33770;
  wire n_33771, n_33772, n_33773, n_33774, n_33775, n_33776, n_33777,
       n_33778;
  wire n_33779, n_33780, n_33781, n_33782, n_33783, n_33784, n_33785,
       n_33786;
  wire n_33787, n_33788, n_33789, n_33790, n_33791, n_33792, n_33793,
       n_33794;
  wire n_33795, n_33796, n_33797, n_33798, n_33799, n_33800, n_33801,
       n_33802;
  wire n_33803, n_33804, n_33805, n_33806, n_33807, n_33808, n_33809,
       n_33810;
  wire n_33811, n_33812, n_33813, n_33814, n_33815, n_33816, n_33817,
       n_33818;
  wire n_33819, n_33820, n_33821, n_33822, n_33823, n_33824, n_33825,
       n_33826;
  wire n_33827, n_33828, n_33829, n_33832, n_33833, n_33835, n_33836,
       n_33852;
  wire n_33853, n_33854, n_33855, n_33856, n_33857, n_33858, n_33859,
       n_33860;
  wire n_33861, n_33862, n_33863, n_33864, n_33865, n_33866, n_33867,
       n_33868;
  wire n_33869, n_33870, n_33871, n_33872, n_33873, n_33874, n_33875,
       n_33876;
  wire n_33877, n_33878, n_33879, n_33880, n_33881, n_33882, n_33883,
       n_33893;
  wire n_33894, n_33895, n_33896, n_33897, n_33898, n_33899, n_33900,
       n_33901;
  wire n_33902, n_33903, n_33904, n_33905, n_33906, n_33907, n_33908,
       n_33909;
  wire n_33910, n_33911, n_33912, n_33913, n_33914, n_33915, n_33916,
       n_33917;
  wire n_33918, n_33919, n_33920, n_33921, n_33922, n_33923, n_33924,
       n_33925;
  wire n_33926, n_33927, n_33928, n_33929, n_33930, n_33931, n_33932,
       n_33933;
  wire n_33934, n_33935, n_33942, n_33943, n_33944, n_33945, n_33946,
       n_33947;
  wire n_33948, n_33949, n_33950, n_33951, n_33952, n_33953, n_33954,
       n_33955;
  wire n_33956, n_33957, n_33958, n_33959, n_33960, n_33961, n_33962,
       n_33963;
  wire n_33964, n_33965, n_33966, n_33967, n_33968, n_33969, n_33970,
       n_33971;
  wire n_33972, n_33973, n_33974, n_33975, n_33976, n_33977, n_33978,
       n_33979;
  wire n_33980, n_33981, n_33982, n_33983, n_33984, n_33985, n_33986,
       n_33987;
  wire n_33988, n_33989, n_33990, n_33991, n_33992, n_33993, n_33994,
       n_33995;
  wire n_33996, n_33997, n_33998, n_33999, n_34000, n_34001, n_34002,
       n_34003;
  wire n_34004, n_34005, n_34006, n_34007, n_34008, n_34009, n_34010,
       n_34011;
  wire n_34012, n_34013, n_34014, n_34015, n_34016, n_34017, n_34018,
       n_34019;
  wire n_34020, n_34021, n_34022, n_34023, n_34024, n_34025, n_34026,
       n_34027;
  wire n_34028, n_34029, n_34030, n_34031, n_34032, n_34033, n_34034,
       n_34035;
  wire n_34036, n_34037, n_34038, n_34039, n_34040, n_34041, n_34042,
       n_34043;
  wire n_34044, n_34045, n_34046, n_34047, n_34048, n_34049, n_34050,
       n_34051;
  wire n_34052, n_34053, n_34054, n_34055, n_34056, n_34057, n_34058,
       n_34059;
  wire n_34060, n_34061, n_34062, n_34063, n_34064, n_34065, n_34066,
       n_34067;
  wire n_34068, n_34069, n_34070, n_34071, n_34072, n_34073, n_34074,
       n_34075;
  wire n_34076, n_34077, n_34078, n_34079, n_34080, n_34081, n_34082,
       n_34083;
  wire n_34084, n_34085, n_34086, n_34087, n_34088, n_34089, n_34090,
       n_34091;
  wire n_34092, n_34093, n_34094, n_34095, n_34096, n_34097, n_34098,
       n_34099;
  wire n_34100, n_34101, n_34102, n_34103, n_34104, n_34105, n_34106,
       n_34107;
  wire n_34108, n_34109, n_34110, n_34111, n_34112, n_34113, n_34114,
       n_34115;
  wire n_34116, n_34117, n_34118, n_34119, n_34120, n_34121, n_34122,
       n_34123;
  wire n_34124, n_34125, n_34126, n_34127, n_34128, n_34129, n_34130,
       n_34131;
  wire n_34132, n_34133, n_34134, n_34135, n_34136, n_34137, n_34138,
       n_34139;
  wire n_34140, n_34141, n_34142, n_34143, n_34144, n_34145, n_34146,
       n_34147;
  wire n_34148, n_34149, n_34150, n_34151, n_34152, n_34153, n_34154,
       n_34155;
  wire n_34156, n_34157, n_34158, n_34159, n_34160, n_34161, n_34162,
       n_34163;
  wire n_34164, n_34165, n_34166, n_34167, n_34168, n_34169, n_34170,
       n_34171;
  wire n_34172, n_34173, n_34174, n_34175, n_34176, n_34177, n_34178,
       n_34179;
  wire n_34180, n_34181, n_34182, n_34183, n_34184, n_34185, n_34186,
       n_34187;
  wire n_34188, n_34189, n_34190, n_34191, n_34192, n_34193, n_34194,
       n_34195;
  wire n_34196, n_34197, n_34198, n_34199, n_34200, n_34201, n_34202,
       n_34203;
  wire n_34204, n_34205, n_34206, n_34207, n_34208, n_34209, n_34210,
       n_34211;
  wire n_34212, n_34213, n_34214, n_34215, n_34216, n_34217, n_34218,
       n_34219;
  wire n_34220, n_34221, n_34222, n_34223, n_34224, n_34225, n_34226,
       n_34227;
  wire n_34228, n_34229, n_34230, n_34231, n_34232, n_34233, n_34234,
       n_34235;
  wire n_34236, n_34237, n_34238, n_34239, n_34240, n_34241, n_34242,
       n_34243;
  wire n_34244, n_34245, n_34246, n_34247, n_34248, n_34249, n_34250,
       n_34251;
  wire n_34252, n_34253, n_34254, n_34255, n_34256, n_34257, n_34258,
       n_34259;
  wire n_34260, n_34261, n_34262, n_34263, n_34264, n_34265, n_34266,
       n_34267;
  wire n_34268, n_34269, n_34270, n_34271, n_34272, n_34273, n_34274,
       n_34275;
  wire n_34276, n_34277, n_34278, n_34279, n_34280, n_34281, n_34282,
       n_34283;
  wire n_34284, n_34285, n_34286, n_34287, n_34288, n_34289, n_34290,
       n_34291;
  wire n_34292, n_34293, n_34294, n_34295, n_34296, n_34297, n_34303,
       n_34304;
  wire n_34305, n_34306, n_34307, n_34308, n_34309, n_34310, n_34311,
       n_34312;
  wire n_34313, n_34314, n_34315, n_34316, n_34317, n_34318, n_34319,
       n_34320;
  wire n_34321, n_34322, n_34323, n_34324, n_34325, n_34326, n_34327,
       n_34328;
  wire n_34329, n_34330, n_34331, n_34332, n_34333, n_34334, n_34335,
       n_34336;
  wire n_34337, n_34338, n_34339, n_34340, n_34341, n_34342, n_34348,
       n_34349;
  wire n_34350, n_34351, n_34352, n_34353, n_34354, n_34355, n_34356,
       n_34357;
  wire n_34358, n_34359, n_34360, n_34361, n_34362, n_34363, n_34364,
       n_34365;
  wire n_34366, n_34367, n_34368, n_34369, n_34370, n_34371, n_34372,
       n_34373;
  wire n_34374, n_34375, n_34376, n_34377, n_34378, n_34379, n_34380,
       n_34381;
  wire n_34382, n_34383, n_34384, n_34385, n_34386, n_34387, n_34388,
       n_34389;
  wire n_34390, n_34391, n_34392, n_34393, n_34394, n_34395, n_34396,
       n_34397;
  wire n_34398, n_34399, n_34400, n_34401, n_34402, n_34403, n_34404,
       n_34405;
  wire n_34406, n_34407, n_34408, n_34409, n_34410, n_34411, n_34412,
       n_34413;
  wire n_34414, n_34415, n_34416, n_34417, n_34418, n_34419, n_34420,
       n_34421;
  wire n_34422, n_34423, n_34424, n_34425, n_34426, n_34427, n_34428,
       n_34429;
  wire n_34430, n_34431, n_34432, n_34433, n_34434, n_34435, n_34436,
       n_34437;
  wire n_34438, n_34439, n_34440, n_34441, n_34442, n_34443, n_34444,
       n_34445;
  wire n_34446, n_34447, n_34448, n_34449, n_34450, n_34451, n_34452,
       n_34453;
  wire n_34454, n_34455, n_34456, n_34457, n_34458, n_34459, n_34460,
       n_34461;
  wire n_34462, n_34463, n_34464, n_34465, n_34466, n_34467, n_34468,
       n_34469;
  wire n_34470, n_34471, n_34472, n_34473, n_34474, n_34475, n_34476,
       n_34477;
  wire n_34478, n_34479, n_34480, n_34481, n_34482, n_34483, n_34484,
       n_34496;
  wire n_34497, n_34498, n_34499, n_34500, n_34501, n_34502, n_34503,
       n_34504;
  wire n_34505, n_34506, n_34507, n_34508, n_34509, n_34510, n_34511,
       n_34512;
  wire n_34513, n_34514, n_34515, n_34516, n_34517, n_34518, n_34519,
       n_34520;
  wire n_34521, n_34522, n_34523, n_34524, n_34525, n_34526, n_34527,
       n_34528;
  wire n_34529, n_34530, n_34531, n_34532, n_34539, n_34540, n_34541,
       n_34542;
  wire n_34543, n_34544, n_34545, n_34547, n_34548, n_34549, n_34550,
       n_34551;
  wire n_34552, n_34553, n_34554, n_34555, n_34556, n_34557, n_34558,
       n_34559;
  wire n_34560, n_34561, n_34562, n_34563, n_34564, n_34565, n_34566,
       n_34567;
  wire n_34568, n_34569, n_34570, n_34571, n_34572, n_34573, n_34574,
       n_34575;
  wire n_34576, n_34577, n_34578, n_34579, n_34580, n_34581, n_34582,
       n_34583;
  wire n_34584, n_34585, n_34586, n_34587, n_34588, n_34589, n_34590,
       n_34591;
  wire n_34592, n_34593, n_34594, n_34595, n_34596, n_34597, n_34598,
       n_34599;
  wire n_34600, n_34601, n_34602, n_34603, n_34604, n_34605, n_34606,
       n_34607;
  wire n_34608, n_34609, n_34610, n_34611, n_34612, n_34613, n_34614,
       n_34615;
  wire n_34616, n_34617, n_34618, n_34619, n_34620, n_34621, n_34622,
       n_34623;
  wire n_34624, n_34625, n_34626, n_34627, n_34628, n_34629, n_34630,
       n_34631;
  wire n_34632, n_34633, n_34634, n_34635, n_34636, n_34637, n_34638,
       n_34639;
  wire n_34640, n_34641, n_34642, n_34643, n_34644, n_34645, n_34647,
       n_34648;
  wire n_34649, n_34650, n_34651, n_34652, n_34653, n_34654, n_34655,
       n_34656;
  wire n_34657, n_34658, n_34659, n_34660, n_34661, n_34663, n_34665,
       n_34668;
  wire n_34669, n_34670, n_34671, n_34672, n_34673, n_34675, n_34676,
       n_34677;
  wire n_34678, n_34679, n_34686, n_34688, n_34693, n_34695, n_34696,
       n_34697;
  wire n_34698, n_34699, n_34700, n_34701, n_34704, n_34707, n_34708,
       n_34709;
  wire n_34710, n_34711, n_34712, n_34714, n_34715, n_34716, n_34717,
       n_34719;
  wire n_34720, n_34721, n_34723, n_34724, n_34725, n_34727, n_34728,
       n_34729;
  wire n_34731, n_34732, n_34733, n_34735, n_34737, n_34738, n_34739,
       n_34741;
  wire n_34743, n_34744, n_34745, n_34747, n_34748, n_34749, n_34751,
       n_34753;
  wire n_34754, n_34755, n_34757, n_34758, n_34759, n_34761, n_34762,
       n_34765;
  wire n_34766, n_34767, n_34769, n_34770, n_34771, n_34772, n_34774,
       n_34775;
  wire n_34776, n_34778, n_34779, n_34780, n_34782, n_34783, n_34784,
       n_34786;
  wire n_34788, n_34789, n_34790, n_34792, n_34793, n_34794, n_34796,
       n_34797;
  wire n_34798, n_34800, n_34801, n_34802, n_34804, n_34806, n_34807,
       n_34815;
  wire n_34817, n_34819, n_34820, n_34821, n_34823, n_34824, n_34825,
       n_34826;
  wire n_34827, n_34829, n_34830, n_34831, n_34832, n_34833, n_34835,
       n_34836;
  wire n_34837, n_34839, n_34840, n_34842, n_34843, n_34845, n_34846,
       n_34847;
  wire n_34848, n_34849, n_34851, n_34852, n_34854, n_34856, n_34857,
       n_34858;
  wire n_34859, n_34860, n_34861, n_34862, n_34863, n_34864, n_34866,
       n_34868;
  wire n_34869, n_34870, n_34871, n_34872, n_34874, n_34875, n_34876,
       n_34877;
  wire n_34878, n_34880, n_34881, n_34882, n_34884, n_34886, n_34887,
       n_34888;
  wire n_34890, n_34891, n_34892, n_34893, n_34894, n_34895, n_34897,
       n_34899;
  wire n_34900, n_34902, n_34903, n_34905, n_34907, n_34908, n_34909,
       n_34911;
  wire n_34913, n_34914, n_34915, n_34917, n_34919, n_34920, n_34921,
       n_34923;
  wire n_34924, n_34926, n_34928, n_34929, n_34931, n_34932, n_34933,
       n_34935;
  wire n_34936, n_34938, n_34939, n_34940, n_34942, n_34943, n_34944,
       n_34945;
  wire n_34946, n_34947, n_34948, n_34949, n_34950, n_34952, n_34953,
       n_34954;
  wire n_34955, n_34956, n_34957, n_34958, n_34959, n_34960, n_34961,
       n_34962;
  wire n_34963, n_34964, n_34965, n_34966, n_34967, n_34968, n_34969,
       n_34970;
  wire n_34971, n_34972, n_34973, n_34974, n_34976, n_34977, n_34978,
       n_34979;
  wire n_34980, n_34981, n_34982, n_34983, n_34984, n_34986, n_34987,
       n_34991;
  wire n_34992, n_34993, n_34994, n_34995, n_34996, n_34997, n_34998,
       n_34999;
  wire n_35000, n_35001, n_35002, n_35003, n_35004, n_35005, n_35006,
       n_35007;
  wire n_35008, n_35009, n_35010, n_35011, n_35012, n_35013, n_35014,
       n_35016;
  wire n_35017, n_35018, n_35019, n_35020, n_35021, n_35022, n_35023,
       n_35024;
  wire n_35025, n_35026, n_35028, n_35029, n_35030, n_35031, n_35032,
       n_35034;
  wire n_35038, n_35039, n_35040, n_35041, n_35042, n_35043, n_35044,
       n_35045;
  wire n_35046, n_35047, n_35048, n_35049, n_35050, n_35051, n_35052,
       n_35053;
  wire n_35054, n_35055, n_35056, n_35057, n_35058, n_35059, n_35060,
       n_35061;
  wire n_35062, n_35063, n_35064, n_35065, n_35066, n_35067, n_35068,
       n_35069;
  wire n_35070, n_35071, n_35072, n_35073, n_35074, n_35076, n_35077,
       n_35078;
  wire n_35079, n_35080, n_35081, n_35082, n_35083, n_35084, n_35085,
       n_35087;
  wire n_35088, n_35089, n_35090, n_35091, n_35092, n_35096, n_35097,
       n_35098;
  wire n_35099, n_35100, n_35101, n_35102, n_35103, n_35104, n_35105,
       n_35106;
  wire n_35107, n_35108, n_35109, n_35110, n_35111, n_35112, n_35114,
       n_35115;
  wire n_35116, n_35117, n_35118, n_35119, n_35120, n_35121, n_35122,
       n_35123;
  wire n_35124, n_35125, n_35126, n_35127, n_35128, n_35129, n_35131,
       n_35137;
  wire n_35138, n_35139, n_35140, n_35141, n_35142, n_35143, n_35144,
       n_35145;
  wire n_35146, n_35147, n_35148, n_35149, n_35150, n_35151, n_35152,
       n_35153;
  wire n_35154, n_35156, n_35162, n_35163, n_35164, n_35165, n_35166,
       n_35168;
  wire n_35169, n_35170, n_35171, n_35172, n_35173, n_35177, n_35178,
       n_35179;
  wire n_35180, n_35181, n_35182, n_35183, n_35184, n_35185, n_35186,
       n_35187;
  wire n_35188, n_35189, n_35190, n_35191, n_35192, n_35193, n_35194,
       n_35195;
  wire n_35197, n_35198, n_35199, n_35200, n_35201, n_35203, n_35207,
       n_35208;
  wire n_35209, n_35210, n_35211, n_35212, n_35213, n_35214, n_35215,
       n_35216;
  wire n_35217, n_35218, n_35219, n_35220, n_35221, n_35222, n_35223,
       n_35224;
  wire n_35225, n_35226, n_35227, n_35228, n_35229, n_35230, n_35231,
       n_35232;
  wire n_35233, n_35234, n_35235, n_35236, n_35237, n_35239, n_35240,
       n_35241;
  wire n_35242, n_35243, n_35244, n_35246, n_35247, n_35248, n_35249,
       n_35250;
  wire n_35251, n_35252, n_35254, n_35255, n_35256, n_35257, n_35258,
       n_35259;
  wire n_35261, n_35262, n_35263, n_35264, n_35265, n_35266, n_35267,
       n_35268;
  wire n_35269, n_35270, n_35271, n_35272, n_35273, n_35274, n_35275,
       n_35276;
  wire n_35277, n_35278, n_35279, n_35280, n_35281, n_35282, n_35283,
       n_35284;
  wire n_35285, n_35287, n_35288, n_35289, n_35290, n_35291, n_35293,
       n_35297;
  wire n_35298, n_35299, n_35300, n_35301, n_35302, n_35303, n_35304,
       n_35305;
  wire n_35306, n_35307, n_35308, n_35309, n_35310, n_35311, n_35312,
       n_35313;
  wire n_35314, n_35315, n_35316, n_35317, n_35318, n_35319, n_35320,
       n_35321;
  wire n_35322, n_35323, n_35324, n_35325, n_35326, n_35327, n_35329,
       n_35335;
  wire n_35336, n_35337, n_35338, n_35339, n_35340, n_35341, n_35342,
       n_35343;
  wire n_35344, n_35345, n_35346, n_35347, n_35348, n_35349, n_35350,
       n_35351;
  wire n_35352, n_35354, n_35360, n_35361, n_35362, n_35363, n_35364,
       n_35365;
  wire n_35366, n_35367, n_35368, n_35369, n_35370, n_35371, n_35372,
       n_35373;
  wire n_35374, n_35375, n_35376, n_35378, n_35379, n_35380, n_35381,
       n_35382;
  wire n_35383, n_35384, n_35385, n_35387, n_35391, n_35392, n_35393,
       n_35394;
  wire n_35395, n_35396, n_35397, n_35398, n_35399, n_35400, n_35401,
       n_35402;
  wire n_35403, n_35404, n_35405, n_35406, n_35407, n_35408, n_35409,
       n_35410;
  wire n_35411, n_35412, n_35414, n_35420, n_35421, n_35422, n_35425,
       n_35426;
  wire n_35427, n_35428, n_35429, n_35430, n_35431, n_35432, n_35433,
       n_35434;
  wire n_35435, n_35436, n_35437, n_35438, n_35439, n_35440, n_35441,
       n_35445;
  wire n_35446, n_35447, n_35448, n_35449, n_35450, n_35451, n_35452,
       n_35453;
  wire n_35455, n_35456, n_35457, n_35458, n_35459, n_35460, n_35461,
       n_35462;
  wire n_35463, n_35464, n_35465, n_35466, n_35467, n_35468, n_35469,
       n_35470;
  wire n_35471, n_35472, n_35473, n_35474, n_35475, n_35476, n_35477,
       n_35478;
  wire n_35479, n_35480, n_35481, n_35483, n_35484, n_35485, n_35486,
       n_35487;
  wire n_35489, n_35493, n_35494, n_35495, n_35496, n_35497, n_35498,
       n_35499;
  wire n_35500, n_35501, n_35502, n_35503, n_35504, n_35505, n_35506,
       n_35507;
  wire n_35508, n_35509, n_35510, n_35511, n_35512, n_35513, n_35514,
       n_35516;
  wire n_35517, n_35518, n_35519, n_35521, n_35522, n_35523, n_35524,
       n_35525;
  wire n_35526, n_35528, n_35529, n_35531, n_35532, n_35533, n_35534,
       n_35535;
  wire n_35536, n_35538, n_35539, n_35540, n_35541, n_35542, n_35543,
       n_35544;
  wire n_35545, n_35546, n_35547, n_35548, n_35549, n_35550, n_35551,
       n_35552;
  wire n_35553, n_35554, n_35555, n_35556, n_35557, n_35558, n_35559,
       n_35560;
  wire n_35561, n_35562, n_35563, n_35564, n_35565, n_35566, n_35567,
       n_35568;
  wire n_35569, n_35570, n_35571, n_35572, n_35573, n_35574, n_35578,
       n_35582;
  wire n_35583, n_35584, n_35585, n_35586, n_35587, n_35588, n_35589,
       n_35590;
  wire n_35591, n_35592, n_35593, n_35594, n_35595, n_35596, n_35597,
       n_35604;
  wire n_35608, n_35609, n_35610, n_35611, n_35612, n_35613, n_35614,
       n_35615;
  wire n_35616, n_35617, n_35618, n_35619, n_35620, n_35621, n_35622,
       n_35623;
  wire n_35624, n_35625, n_35626, n_35627, n_35628, n_35629, n_35630,
       n_35631;
  wire n_35632, n_35636, n_35640, n_35641, n_35642, n_35644, n_35650,
       n_35651;
  wire n_35652, n_35656, n_35657, n_35658, n_35659, n_35660, n_35661,
       n_35662;
  wire n_35663, n_35664, n_35665, n_35666, n_35667, n_35668, n_35669,
       n_35670;
  wire n_35671, n_35672, n_35673, n_35674, n_35675, n_35676, n_35677,
       n_35678;
  wire n_35679, n_35680, n_35681, n_35682, n_35686, n_35690, n_35691,
       n_35692;
  wire n_35693, n_35694, n_35695, n_35696, n_35697, n_35698, n_35699,
       n_35700;
  wire n_35701, n_35702, n_35703, n_35704, n_35705, n_35706, n_35709,
       n_35710;
  wire n_35711, n_35712, n_35713, n_35714, n_35715, n_35717, n_35718,
       n_35719;
  wire n_35720, n_35721, n_35722, n_35723, n_35724, n_35725, n_35726,
       n_35727;
  wire n_35728, n_35729, n_35730, n_35731, n_35732, n_35733, n_35734,
       n_35735;
  wire n_35736, n_35737, n_35744, n_35748, n_35749, n_35750, n_35751,
       n_35752;
  wire n_35753, n_35754, n_35755, n_35756, n_35757, n_35758, n_35759,
       n_35760;
  wire n_35761, n_35762, n_35763, n_35764, n_35766, n_35771, n_35772,
       n_35773;
  wire n_35774, n_35775, n_35776, n_35777, n_35778, n_35779, n_35780,
       n_35781;
  wire n_35782, n_35783, n_35784, n_35785, n_35786, n_35787, n_35788,
       n_35789;
  wire n_35790, n_35791, n_35798, n_35802, n_35803, n_35804, n_35805,
       n_35806;
  wire n_35807, n_35808, n_35809, n_35810, n_35811, n_35812, n_35813,
       n_35814;
  wire n_35815, n_35816, n_35817, n_35818, n_35820, n_35825, n_35826,
       n_35827;
  wire n_35828, n_35829, n_35830, n_35831, n_35832, n_35833, n_35834,
       n_35835;
  wire n_35836, n_35837, n_35838, n_35839, n_35840, n_35841, n_35842,
       n_35843;
  wire n_35844, n_35845, n_35846, n_35849, n_35850, n_35851, n_35852,
       n_35853;
  wire n_35854, n_35855, n_35857, n_35858, n_35859, n_35860, n_35861,
       n_35862;
  wire n_35865, n_35867, n_35868, n_35869, n_35870, n_35872, n_35873,
       n_35874;
  wire n_35875, n_35877, n_35878, n_35879, n_35880, n_35882, n_35883,
       n_35884;
  wire n_35885, n_35886, n_35888, n_35889, n_35890, n_35891, n_35892,
       n_35893;
  wire n_35894, n_35895, n_35896, n_35897, n_35898, n_35899, n_35900,
       n_35901;
  wire n_35902, n_35903, n_35904, n_35905, n_35906, n_35907, n_35908,
       n_35909;
  wire n_35911, n_35913, n_35916, n_35917, n_35918, n_35919, n_35920,
       n_35921;
  wire n_35922, n_35923, n_35924, n_35925, n_35926, n_35927, n_35928,
       n_35929;
  wire n_35930, n_35931, n_35932, n_35933, n_35934, n_35935, n_35936,
       n_35937;
  wire n_35938, n_35939, n_35940, n_35941, n_35942, n_35944, n_35945,
       n_35946;
  wire n_35948, n_35949, n_35950, n_35951, n_35952, n_35956, n_35957,
       n_35958;
  wire n_35959, n_35960, n_35961, n_35962, n_35963, n_35964, n_35965,
       n_35966;
  wire n_35967, n_35968, n_35969, n_35970, n_35971, n_35972, n_35973,
       n_35974;
  wire n_35975, n_35976, n_35977, n_35978, n_35979, n_35980, n_35981,
       n_35982;
  wire n_35983, n_35984, n_35985, n_35986, n_35987, n_35988, n_35989,
       n_35990;
  wire n_35991, n_35992, n_35993, n_35994, n_35995, n_35996, n_35997,
       n_35998;
  wire n_35999, n_36000, n_36001, n_36002, n_36009, n_36013, n_36014,
       n_36015;
  wire n_36016, n_36017, n_36018, n_36019, n_36020, n_36021, n_36022,
       n_36023;
  wire n_36024, n_36025, n_36026, n_36027, n_36029, n_36030, n_36031,
       n_36032;
  wire n_36033, n_36034, n_36035, n_36036, n_36037, n_36038, n_36039,
       n_36040;
  wire n_36041, n_36042, n_36043, n_36044, n_36045, n_36046, n_36047,
       n_36049;
  wire n_36050, n_36051, n_36052, n_36053, n_36054, n_36055, n_36056,
       n_36057;
  wire n_36058, n_36059, n_36060, n_36061, n_36062, n_36063, n_36064,
       n_36065;
  wire n_36066, n_36067, n_36068, n_36069, n_36070, n_36071, n_36072,
       n_36073;
  wire n_36074, n_36075, n_36076, n_36077, n_36078, n_36079, n_36080,
       n_36081;
  wire n_36082, n_36083, n_36084, n_36085, n_36086, n_36087, n_36089,
       n_36090;
  wire n_36091, n_36092, n_36093, n_36094, n_36095, n_36096, n_36097,
       n_36098;
  wire n_36099, n_36100, n_36101, n_36102, n_36103, n_36104, n_36105,
       n_36106;
  wire n_36107, n_36108, n_36109, n_36110, n_36111, n_36112, n_36113,
       n_36114;
  wire n_36115, n_36116, n_36117, n_36118, n_36119, n_36120, n_36121,
       n_36122;
  wire n_36123, n_36124, n_36125, n_36126, n_36127, n_36128, n_36131,
       n_36132;
  wire n_36133, n_36134, n_36135, n_36136, n_36137, n_36138, n_36139,
       n_36140;
  wire n_36141, n_36142, n_36143, n_36144, n_36145, n_36146, n_36147,
       n_36148;
  wire n_36149, n_36150, n_36151, n_36152, n_36153, n_36154, n_36155,
       n_36156;
  wire n_36164, n_36165, n_36166, n_36167, n_36168, n_36169, n_36170,
       n_36171;
  wire n_36172, n_36173, n_36174, n_36175, n_36176, n_36177, n_36178,
       n_36179;
  wire n_36180, n_36181, n_36182, n_36183, n_36184, n_36185, n_36186,
       n_36187;
  wire n_36188, n_36189, n_36190, n_36191, n_36192, n_36193, n_36194,
       n_36196;
  wire n_36197, n_36198, n_36199, n_36200, n_36201, n_36202, n_36203,
       n_36204;
  wire n_36207, n_36208, n_36209, n_36210, n_36211, n_36212, n_36213,
       n_36214;
  wire n_36215, n_36216, n_36217, n_36218, n_36219, n_36220, n_36221,
       n_36222;
  wire n_36223, n_36224, n_36225, n_36226, n_36227, n_36228, n_36229,
       n_36230;
  wire n_36231, n_36234, n_36235, n_36236, n_36237, n_36238, n_36239,
       n_36240;
  wire n_36241, n_36242, n_36243, n_36244, n_36245, n_36246, n_36247,
       n_36248;
  wire n_36249, n_36250, n_36251, n_36252, n_36253, n_36254, n_36255,
       n_36256;
  wire n_36257, n_36258, n_36261, n_36262, n_36263, n_36264, n_36265,
       n_36266;
  wire n_36267, n_36268, n_36269, n_36270, n_36271, n_36272, n_36273,
       n_36274;
  wire n_36275, n_36276, n_36277, n_36278, n_36279, n_36280, n_36281,
       n_36282;
  wire n_36283, n_36284, n_36285, n_36288, n_36289, n_36290, n_36291,
       n_36292;
  wire n_36293, n_36294, n_36295, n_36296, n_36297, n_36298, n_36299,
       n_36300;
  wire n_36301, n_36302, n_36303, n_36304, n_36305, n_36306, n_36307,
       n_36308;
  wire n_36309, n_36310, n_36311, n_36312, n_36313, n_36314, n_36315,
       n_36317;
  wire n_36318, n_36320, n_36323, n_36324, n_36325, n_36326, n_36327,
       n_36330;
  wire n_36331, n_36332, n_36333, n_36334, n_36335, n_36336, n_36337,
       n_36338;
  wire n_36339, n_36340, n_36341, n_36342, n_36343, n_36344, n_36345,
       n_36346;
  wire n_36347, n_36348, n_36349, n_36350, n_36351, n_36352, n_36353,
       n_36354;
  wire n_36355, n_36356, n_36400, n_36401, n_36402, n_36403, n_36404,
       n_36405;
  wire n_36406, n_36407, n_36408, n_36409, n_36410, n_36411, n_36424,
       n_36425;
  wire n_36436, n_36437, n_36438, n_36439, n_36440, n_36441, n_36442,
       n_36443;
  wire n_36444, n_36445, n_36446, n_36447, n_36448, n_36449, n_36450,
       n_36451;
  wire n_36452, n_36453, n_36454, n_36455, n_36456, n_36457, n_36458,
       n_36459;
  wire n_36460, n_36461, n_36462, n_36463, n_36464, n_36465, n_36466,
       n_36467;
  wire n_36468, n_36469, n_36470, n_36471, n_36472, n_36473, n_36474,
       n_37592;
  wire n_37593, n_37594, n_37595, n_37596, n_37597, n_37598, n_37599,
       n_37600;
  wire n_37601, n_37602, n_37603, n_37604, n_37605, n_37606, n_37607,
       n_37608;
  wire n_37609, n_37610, n_37611, n_37612, n_37613, n_37614, n_37615,
       n_37616;
  wire n_37617, n_37618, n_37619, n_37620, n_37621, n_37622, n_37623,
       n_37624;
  wire n_37625, n_37626, n_37627, n_37628, n_37629, n_37630, n_37631,
       n_37632;
  wire n_37633, n_37634, n_37635, n_37636, n_37637, n_37638, n_37639,
       n_37640;
  wire n_37641, n_37642, n_37643, n_37644, n_37645, n_37646, n_37647,
       n_37648;
  wire n_37649, n_37650, n_37651, n_37652, n_37653, n_37654, n_37655,
       n_37656;
  wire n_37657, n_37658, n_37659, n_37660, n_37661, n_37662, n_37663,
       n_37664;
  wire n_37665, n_37666, n_37667, n_37668, n_37669, n_37670, n_37671,
       n_37672;
  wire n_37673, n_37674, n_37675, n_37676, n_37677, n_37678, n_37679,
       n_37680;
  wire n_37681, n_37682, n_37683, n_37684, n_37685, n_37686, n_37687,
       n_37688;
  wire n_37689, n_37690, n_37691, n_37692, n_37693, n_37694, n_37695,
       n_37696;
  wire n_37697, n_37698, n_37699, n_37700, n_37702, n_37703, n_37704,
       n_37705;
  wire n_37706, n_37707, n_37708, n_37709, n_37710, n_37711, n_37712,
       n_37713;
  wire n_37714, n_37715, n_37716, n_37717, n_37718, n_37719, n_37720,
       n_37721;
  wire n_37722, n_37723, n_37724, n_37725, n_37726, n_37727, n_37728,
       n_37729;
  wire n_37730, n_37731, n_37732, n_37733, n_37734, n_37735, n_37736,
       n_37737;
  wire n_37738, n_37739, n_37740, n_37741, n_37742, n_37743, n_37744,
       n_37745;
  wire n_37746, n_37747, n_37748, n_37749, n_37750, n_37751, n_37752,
       n_37753;
  wire n_37754, n_37755, n_37756, n_37757, n_37758, n_37759, n_37760,
       n_37761;
  wire n_37762, n_37763, n_37764, n_37765, n_37766, n_37767, n_37768,
       n_37769;
  wire n_37770, n_37771, n_37772, n_37773, n_37774, n_37775, n_37776,
       n_37777;
  wire n_37778, n_37779, n_37780, n_37781, n_37782, n_37783, n_37784,
       n_37785;
  wire n_37786, n_37787, n_37788, n_37789, n_37790, n_37791, n_37792,
       n_37793;
  wire n_37794, n_37795, n_37796, n_37797, n_37798, n_37799, n_37800,
       n_37801;
  wire n_37802, n_37803, n_37804, n_37805, n_37806, n_37807, n_37808,
       n_37809;
  wire n_37810, n_37811, n_37812, n_37813, n_37814, n_37815, n_37816,
       n_37817;
  wire n_37818, n_37819, n_37820, n_37821, n_37822, n_37823, n_37824,
       n_37825;
  wire n_37826, n_37827, n_37828, n_37829, n_37830, n_37831, n_37832,
       n_37833;
  wire n_37834, n_37835, n_37836, n_37837, n_37838, n_37839, n_37840,
       n_37841;
  wire n_37842, n_37843, n_37844, n_37845, n_37846, n_37847, n_37848,
       n_37849;
  wire n_37850, n_37851, n_37852, n_37853, n_37854, n_37855, n_37856,
       n_37857;
  wire n_37858, n_37859, n_37860, n_37861, n_37862, n_37863, n_37864,
       n_37865;
  wire n_37866, n_37867, n_37868, n_37869, n_37870, n_37871, n_37872,
       n_37873;
  wire n_37874, n_37875, n_37876, n_37877, n_37878, n_37879, n_37880,
       n_37881;
  wire n_37882, n_37883, n_37884, n_37885, n_37886, n_37887, n_37888,
       n_37889;
  wire n_37890, n_37891, n_37892, n_37893, n_37894, n_37895, n_37896,
       n_37897;
  wire n_37898, n_37899, n_37900, n_37901, n_37902, n_37903, n_37904,
       n_37905;
  wire n_37906, n_37907, n_37908, n_37909, n_37910, n_37911, n_37912,
       n_37913;
  wire n_37914, n_37915, n_37916, n_37917, n_37918, n_37919, n_37920,
       n_37921;
  wire n_37922, n_37923, n_37924, n_37925, n_37926, n_37927, n_37928,
       n_37929;
  wire n_37930, n_37931, n_37932, n_37933, n_37934, n_37935, n_37936,
       n_37937;
  wire n_37938, n_37939, n_37940, n_37941, n_37942, n_37943, n_37944,
       n_37945;
  wire n_37946, n_37947, n_37948, n_37949, n_37950, n_37951, n_37952,
       n_37953;
  wire n_37954, n_37955, n_37956, n_37957, n_37958, n_37959, n_37960,
       n_37961;
  wire n_37962, n_37963, n_37964, n_37965, n_37966, n_37967, n_37968,
       n_37969;
  wire n_37970, n_37971, n_37972, n_37973, n_37974, n_37975, n_37976,
       n_37977;
  wire n_37978, n_37979, n_37980, n_37981, n_37982, n_37983, n_37984,
       n_37985;
  wire n_37986, n_37987, n_37988, n_37989, n_37990, n_37991, n_37992,
       n_37993;
  wire n_37994, n_37995, n_37996, n_37997, n_37998, n_37999, n_38000,
       n_38001;
  wire n_38002, n_38003, n_38004, n_38005, n_38006, n_38007, n_38008,
       n_38009;
  wire n_38010, n_38011, n_38012, n_38013, n_38014, n_38015, n_38016,
       n_38017;
  wire n_38018, n_38019, n_38020, n_38021, n_38022, n_38023, n_38024,
       n_38025;
  wire n_38026, n_38027, n_38028, n_38029, n_38030, n_38031, n_38032,
       n_38033;
  wire n_38034, n_38035, n_38036, n_38037, n_38038, n_38039, n_38040,
       n_38041;
  wire n_38042, n_38043, n_38044, n_38045, n_38046, n_38047, n_38048,
       n_38049;
  wire n_38050, n_38051, n_38052, n_38053, n_38054, n_38055, n_38056,
       n_38057;
  wire n_38058, n_38059, n_38060, n_38061, n_38062, n_38063, n_38064,
       n_38065;
  wire n_38066, n_38067, n_38068, n_38069, n_38070, n_38071, n_38072,
       n_38073;
  wire n_38074, n_38075, n_38076, n_38077, n_38078, n_38079, n_38080,
       n_38081;
  wire n_38082, n_38083, n_38084, n_38085, n_38086, n_38087, n_38088,
       n_38089;
  wire n_38090, n_38091, n_38092, n_38093, n_38094, n_38095, n_38096,
       n_38097;
  wire n_38098, n_38099, n_38100, n_38101, n_38102, n_38103, n_38104,
       n_38105;
  wire n_38106, n_38107, n_38108, n_38109, n_38110, n_38111, n_38112,
       n_38113;
  wire n_38114, n_38115, n_38116, n_38117, n_38118, n_38119, n_38120,
       n_38121;
  wire n_38122, n_38123, n_38124, n_38125, n_38126, n_38127, n_38128,
       n_38129;
  wire n_38130, n_38131, n_38132, n_38133, n_38134, n_38135, n_38136,
       n_38137;
  wire n_38138, n_38139, n_38140, n_38141, n_38142, n_38143, n_38144,
       n_38145;
  wire n_38146, n_38147, n_38148, n_38149, n_38150, n_38151, n_38152,
       n_38153;
  wire n_38154, n_38155, n_38156, n_38157, n_38158, n_38159, n_38160,
       n_38161;
  wire n_38162, n_38163, n_38164, n_38165, n_38166, n_38167, n_38168,
       n_38169;
  wire n_38170, n_38171, n_38172, n_38173, n_38174, n_38175, n_38176,
       n_38177;
  wire n_38178, n_38179, n_38180, n_38181, n_38182, n_38183, n_38184,
       n_38185;
  wire n_38186, n_38187, n_38188, n_38189, n_38190, n_38191, n_38192,
       n_38193;
  wire n_38194, n_38195, n_38196, n_38197, n_38198, n_38199, n_38200,
       n_38201;
  wire n_38202, n_38203, n_38204, n_38205, n_38206, n_38207, n_38208,
       n_38209;
  wire n_38210, n_38211, n_38212, n_38213, n_38214, n_38215, n_38216,
       n_38217;
  wire n_38218, n_38219, n_38220, n_38221, n_38222, n_38223, n_38224,
       n_38225;
  wire n_38226, n_38227, n_38228, n_38229, n_38230, n_38231, n_38232,
       n_38233;
  wire n_38234, n_38235, n_38236, n_38237, n_38238, n_38239, n_38240,
       n_38241;
  wire n_38242, n_38243, n_38244, n_38245, n_38246, n_38247, n_38248,
       n_38249;
  wire n_38250, n_38251, n_38252, n_38253, n_38254, n_38255, n_38256,
       n_38257;
  wire n_38258, n_38259, n_38260, n_38261, n_38262, n_38263, n_38264,
       n_38265;
  wire n_38266, n_38267, n_38268, n_38269, n_38270, n_38271, n_38272,
       n_38273;
  wire n_38274, n_38275, n_38276, n_38277, n_38278, n_38279, n_38280,
       n_38281;
  wire n_38282, n_38283, n_38284, n_38285, n_38286, n_38287, n_38288,
       n_38289;
  wire n_38290, n_38291, n_38292, n_38293, n_38294, n_38295, n_38296,
       n_38297;
  wire n_38298, n_38299, n_38300, n_38301, n_38302, n_38303, n_38304,
       n_38305;
  wire n_38306, n_38307, n_38308, n_38309, n_38310, n_38311, n_38312,
       n_38313;
  wire n_38314, n_38315, n_38316, n_38317, n_38318, n_38319, n_38320,
       n_38321;
  wire n_38322, n_38323, n_38324, n_38325, n_38326, n_38327, n_38328,
       n_38329;
  wire n_38330, n_38331, n_38332, n_38333, n_38334, n_38335, n_38336,
       n_38337;
  wire n_38338, n_38339, n_38340, n_38341, n_38342;
  assign po1230 = pi1184;
  assign p-o1229 = pi1200;
  assign po1228 = pi1166;
  assign po1227 = pi1097;
  assign po1226 = pi1194;
  assign po1225 = pi1180;
  assign po1224 = pi1188;
  assign po1223 = pi1190;
  assign po1222 = pi0864;
  assign po1221 = pi1195;
  assign po1220 = pi1189;
  assign po1219 = pi0840;
  assign po1218 = pi1167;
  assign po1217 = pi1201;
  assign po1216 = pi1173;
  assign po1215 = pi1176;
  assign po1214 = pi1202;
  assign po1213 = pi1179;
  assign po1212 = pi1174;
  assign po1211 = pi1099;
  assign po1210 = pi1191;
  assign po1209 = pi1175;
  assign po1208 = pi1168;
  assign po1207 = pi1182;
  assign po1206 = pi1193;
  assign po1205 = pi0849;
  assign po1204 = pi1181;
  assign po1203 = pi1136;
  assign po1202 = pi1169;
  assign po1201 = pi0230;
  assign po1200 = pi1183;
  assign po1199 = pi1098;
  assign po1198 = pi1164;
  assign po1197 = pi1165;
  assign po1196 = pi1186;
  assign po1195 = pi1137;
  assign po1194 = pi1192;
  assign po1193 = pi1171;
  assign po1192 = pi1185;
  assign po1191 = pi1203;
  assign po1190 = pi0863;
  assign po1189 = pi1178;
  assign po1188 = pi1177;
  assign po1187 = pi1138;
  assign po1186 = pi1170;
  assign po1185 = pi1172;
  assign po1184 = pi1187;
  assign po1154 = pi1094;
  assign po1152 = pi1095;
  assign po1145 = pi0279;
  assign po1144 = pi0278;
  assign po1143 = pi0601;
  assign po1142 = pi0605;
  assign po1141 = pi0765;
  assign po1140 = pi0771;
  assign po1139 = pi1052;
  assign po1138 = pi1075;
  assign po1136 = pi0299;
  assign po1134 = pi1064;
  assign po1123 = pi1135;
  assign po1121 = pi1007;
  assign po1120 = pi1004;
  assign po1119 = pi1029;
  assign po1117 = pi1014;
  assign po1114 = pi0985;
  assign po1113 = pi0991;
  assign po1111 = pi0965;
  assign po1109 = pi0964;
  assign po1108 = pi1134;
  assign po1053 = pi0067;
  assign po0636 = pi0583;
  assign po0388 = pi0236;
  assign po0386 = pi0232;
  assign po0285 = pi0131;
  assign po0263 = pi0117;
  assign po0188 = pi0037;
  assign po0181 = po0167;
  assign po0180 = pi0023;
  assign po0179 = pi1089;
  assign po0169 = pi0022;
  assign po0168 = pi0228;
  assign po0166 = 1'b1;
  assign po0152 = pi1096;
  assign po0151 = pi0016;
  assign po0150 = pi0017;
  assign po0149 = pi0018;
  assign po0148 = pi0019;
  assign po0147 = pi0020;
  assign po0146 = pi0021;
  assign po0145 = pi0014;
  assign po0144 = pi0015;
  assign po0143 = pi0029;
  assign po0142 = pi0026;
  assign po0141 = pi0027;
  assign po0140 = pi0028;
  assign po0139 = pi0994;
  assign po0138 = pi0995;
  assign po0137 = pi1033;
  assign po0136 = pi1028;
  assign po0135 = pi0465;
  assign po0134 = pi0469;
  assign po0133 = pi0470;
  assign po0132 = pi0472;
  assign po0131 = pi0471;
  assign po0130 = pi0473;
  assign po0129 = pi0466;
  assign po0128 = pi0474;
  assign po0127 = pi0475;
  assign po0126 = pi0302;
  assign po0125 = pi0310;
  assign po0124 = pi0001;
  assign po0123 = pi0002;
  assign po0122 = pi0000;
  assign po0121 = pi0003;
  assign po0120 = pi0004;
  assign po0119 = pi0005;
  assign po0118 = pi0006;
  assign po0117 = pi0007;
  assign po0116 = pi0008;
  assign po0115 = pi0009;
  assign po0114 = pi0010;
  assign po0113 = pi0011;
  assign po0112 = pi0012;
  assign po0111 = pi0229;
  assign po0110 = pi0834;
  assign po0109 = pi0477;
  assign po0108 = pi0227;
  assign po0107 = pi0808;
  assign po0106 = pi0822;
  assign po0105 = pi0127;
  assign po0104 = pi0226;
  assign po0103 = pi0025;
  assign po0102 = pi0013;
  assign po0101 = pi0112;
  assign po0100 = pi0078;
  assign po0099 = pi0467;
  assign po0098 = pi0893;
  assign po0097 = pi0080;
  assign po0096 = pi0031;
  assign po0095 = pi0998;
  assign po0094 = pi1006;
  assign po0093 = pi1026;
  assign po0092 = pi1002;
  assign po0091 = pi1023;
  assign po0090 = pi1000;
  assign po0089 = pi1022;
  assign po0088 = pi1031;
  assign po0087 = pi1019;
  assign po0086 = pi1008;
  assign po0085 = pi1011;
  assign po0084 = pi1013;
  assign po0083 = pi0997;
  assign po0082 = pi1003;
  assign po0081 = pi1032;
  assign po0080 = pi1009;
  assign po0079 = pi1024;
  assign po0078 = pi1017;
  assign po0077 = pi1018;
  assign po0076 = pi1027;
  assign po0075 = pi1010;
  assign po0074 = pi1021;
  assign po0073 = pi1016;
  assign po0072 = pi0993;
  assign po0071 = pi1012;
  assign po0070 = pi0996;
  assign po0069 = pi1005;
  assign po0068 = pi1025;
  assign po0067 = pi1020;
  assign po0066 = pi1015;
  assign po0065 = pi1034;
  assign po0064 = pi1030;
  assign po0063 = pi0860;
  assign po0062 = pi0880;
  assign po0061 = pi0867;
  assign po0060 = pi0851;
  assign po0059 = pi0868;
  assign po0058 = pi0844;
  assign po0057 = pi0839;
  assign po0056 = pi0843;
  assign po0055 = pi0842;
  assign po0054 = pi0838;
  assign po0053 = pi0845;
  assign po0052 = pi0858;
  assign po0051 = pi0854;
  assign po0050 = pi0857;
  assign po0049 = pi0847;
  assign po0048 = pi0853;
  assign po0047 = pi0856;
  assign po0046 = pi0865;
  assign po0045 = pi0848;
  assign po0044 = pi0870;
  assign po0043 = pi0852;
  assign po0042 = pi0855;
  assign po0041 = pi0859;
  assign po0040 = pi0874;
  assign po0039 = pi0873;
  assign po0038 = pi0876;
  assign po0037 = pi0866;
  assign po0036 = pi0881;
  assign po0035 = pi0871;
  assign po0034 = pi0872;
  assign po0033 = pi0850;
  assign po0032 = pi0837;
  assign po0031 = pi0685;
  assign po0030 = pi0720;
  assign po0029 = pi0714;
  assign po0028 = pi0722;
  assign po0027 = pi0719;
  assign po0026 = pi0692;
  assign po0025 = pi0717;
  assign po0024 = pi0689;
  assign po0023 = pi0712;
  assign po0022 = pi0733;
  assign po0021 = pi0716;
  assign po0020 = pi0711;
  assign po0019 = pi0713;
  assign po0018 = pi0708;
  assign po0017 = pi0707;
  assign po0016 = pi0718;
  assign po0015 = pi0678;
  assign po0014 = pi0671;
  assign po0013 = pi0682;
  assign po0012 = pi0677;
  assign po0011 = pi0670;
  assign po0010 = pi0663;
  assign po0009 = pi0674;
  assign po0008 = pi0679;
  assign po0007 = pi0666;
  assign po0006 = pi0675;
  assign po0005 = pi0673;
  assign po0004 = pi0676;
  assign po0003 = pi0667;
  assign po0002 = pi0664;
  assign po0001 = pi0672;
  assign po0000 = pi0668;
  not g1 (n_4, pi0332);
  not g2 (n_5, pi1144);
  and g3 (n2437, n_4, n_5);
  not g4 (n_7, n2437);
  and g5 (n2438, pi0215, n_7);
  and g6 (n2439, pi0265, n_4);
  not g7 (n_10, n2439);
  and g8 (n2440, pi0216, n_10);
  and g9 (n2441, pi0105, pi0228);
  not g10 (n_15, pi0479);
  and g11 (n2442, pi0095, n_15);
  and g12 (n2443, pi0234, n2442);
  not g13 (n_17, n2443);
  and g14 (n2444, n_4, n_17);
  and g15 (n2445, n2441, n2444);
  and g16 (n2446, pi0153, n_4);
  not g17 (n_19, n2441);
  and g18 (n2447, n_19, n2446);
  not g19 (n_20, pi0216);
  not g20 (n_21, n2447);
  and g21 (n2448, n_20, n_21);
  not g22 (n_22, n2445);
  and g23 (n2449, n_22, n2448);
  not g24 (n_23, n2440);
  not g25 (n_24, n2449);
  and g26 (n2450, n_23, n_24);
  not g27 (n_26, pi0221);
  not g28 (n_27, n2450);
  and g29 (n2451, n_26, n_27);
  and g30 (n2452, n_20, pi0833);
  not g31 (n_29, n2452);
  and g32 (n2453, pi1144, n_29);
  and g33 (n2454, pi0929, n2452);
  not g34 (n_31, n2453);
  and g35 (n2455, n_4, n_31);
  not g36 (n_32, n2454);
  and g37 (n2456, n_32, n2455);
  not g38 (n_33, n2456);
  and g39 (n2457, pi0221, n_33);
  not g40 (n_34, n2451);
  not g41 (n_35, n2457);
  and g42 (n2458, n_34, n_35);
  not g43 (n_36, pi0215);
  not g44 (n_37, n2458);
  and g45 (n2459, n_36, n_37);
  not g46 (n_38, n2438);
  not g47 (n_39, n2459);
  and g48 (n2460, n_38, n_39);
  not g49 (n_42, pi0058);
  not g50 (n_43, pi0090);
  and g51 (n2461, n_42, n_43);
  not g52 (n_46, pi0088);
  not g53 (n_47, pi0098);
  and g54 (n2462, n_46, n_47);
  not g55 (n_49, pi0077);
  and g56 (n2463, n_49, n2462);
  not g57 (n_51, pi0050);
  and g58 (n2464, n_51, n2463);
  not g59 (n_53, pi0102);
  and g60 (n2465, n_53, n2464);
  not g61 (n_56, pi0065);
  not g62 (n_57, pi0071);
  and g63 (n2466, n_56, n_57);
  not g64 (n_60, pi0083);
  not g65 (n_61, pi0103);
  and g66 (n2467, n_60, n_61);
  not g67 (n_64, pi0067);
  not g68 (n_65, pi0069);
  and g69 (n2468, n_64, n_65);
  not g70 (n_68, pi0066);
  not g71 (n_69, pi0073);
  and g72 (n2469, n_68, n_69);
  not g73 (n_72, pi0061);
  not g74 (n_73, pi0076);
  and g75 (n2470, n_72, n_73);
  not g76 (n_76, pi0085);
  not g77 (n_77, pi0106);
  and g78 (n2471, n_76, n_77);
  and g79 (n2472, n2470, n2471);
  not g80 (n_79, pi0048);
  and g81 (n2473, n_79, n2472);
  not g82 (n_81, pi0089);
  and g83 (n2474, n_81, n2473);
  not g84 (n_83, pi0049);
  and g85 (n2475, n_83, n2474);
  not g86 (n_85, pi0104);
  and g87 (n2476, n_85, n2475);
  not g88 (n_87, pi0045);
  and g89 (n2477, n_87, n2476);
  not g90 (n_90, pi0068);
  not g91 (n_91, pi0084);
  and g92 (n2478, n_90, n_91);
  not g93 (n_94, pi0082);
  not g94 (n_95, pi0111);
  and g95 (n2479, n_94, n_95);
  not g96 (n_97, pi0036);
  and g97 (n2480, n_97, n2479);
  and g98 (n2481, n2478, n2480);
  and g99 (n2482, n2477, n2481);
  and g100 (n2483, n2469, n2482);
  and g101 (n2484, n2468, n2483);
  and g102 (n2485, n2467, n2484);
  and g103 (n2486, n2466, n2485);
  not g104 (n_100, pi0063);
  not g105 (n_101, pi0107);
  and g106 (n2487, n_100, n_101);
  and g107 (n2488, n2486, n2487);
  not g108 (n_103, pi0064);
  and g109 (n2489, n_103, n2488);
  not g110 (n_105, pi0081);
  and g111 (n2490, n_105, n2489);
  and g112 (n2491, n2465, n2490);
  not g113 (n_108, pi0047);
  not g114 (n_109, pi0091);
  and g115 (n2492, n_108, n_109);
  not g116 (n_112, pi0109);
  not g117 (n_113, pi0110);
  and g118 (n2493, n_112, n_113);
  not g119 (n_116, pi0053);
  not g120 (n_117, pi0060);
  and g121 (n2494, n_116, n_117);
  not g122 (n_119, pi0086);
  and g123 (n2495, n_119, n2494);
  not g124 (n_122, pi0097);
  not g125 (n_123, pi0108);
  and g126 (n2496, n_122, n_123);
  not g127 (n_125, pi0094);
  and g128 (n2497, n_125, n2496);
  not g129 (n_127, pi0046);
  and g130 (n2498, n_127, n2495);
  and g131 (n2499, n2497, n2498);
  and g132 (n2500, n2493, n2499);
  and g133 (n2501, n2492, n2500);
  and g134 (n2502, n2491, n2501);
  and g135 (n2503, n2461, n2502);
  not g136 (n_130, pi0035);
  not g137 (n_131, pi0093);
  and g138 (n2504, n_130, n_131);
  and g139 (n2505, n2503, n2504);
  not g140 (n_134, pi0072);
  not g141 (n_135, pi0096);
  and g142 (n2506, n_134, n_135);
  not g143 (n_138, pi0051);
  not g144 (n_139, pi0070);
  and g145 (n2507, n_138, n_139);
  and g146 (n2508, n2506, n2507);
  and g147 (n2509, n2505, n2508);
  not g148 (n_142, pi0032);
  not g149 (n_143, pi0040);
  and g150 (n2510, n_142, n_143);
  and g151 (n2511, n2509, n2510);
  not g152 (n_144, pi0095);
  and g153 (n2512, n_144, n2511);
  not g154 (n_145, n2442);
  not g155 (n_146, n2512);
  and g156 (n2513, n_145, n_146);
  not g157 (n_147, n2513);
  and g158 (n2514, pi0234, n_147);
  and g159 (n2515, n_139, n2505);
  and g160 (n2516, n_138, n_135);
  and g161 (n2517, n_143, n_134);
  and g162 (n2518, n_142, n_144);
  and g163 (n2519, n2517, n2518);
  and g164 (n2520, n2516, n2519);
  and g165 (n2521, n2515, n2520);
  not g166 (n_148, pi0234);
  and g167 (n2522, n_148, n2521);
  not g168 (n_149, n2514);
  not g169 (n_150, n2522);
  and g170 (n2523, n_149, n_150);
  not g171 (n_152, n2523);
  and g172 (n2524, pi0137, n_152);
  not g173 (n_153, n2524);
  and g174 (n2525, n2444, n_153);
  and g175 (n2526, n_36, n_26);
  and g176 (n2527, n2448, n2526);
  not g177 (n_154, n2525);
  and g178 (n2528, n_154, n2527);
  not g179 (n_157, pi0056);
  not g180 (n_158, pi0062);
  and g181 (n2529, n_157, n_158);
  not g182 (n_161, pi0038);
  not g183 (n_162, pi0039);
  and g184 (n2530, n_161, n_162);
  not g185 (n_164, pi0100);
  and g186 (n2531, n_164, n2530);
  not g187 (n_167, pi0054);
  not g188 (n_168, pi0074);
  and g189 (n2532, n_167, n_168);
  not g190 (n_171, pi0075);
  not g191 (n_172, pi0087);
  and g192 (n2533, n_171, n_172);
  not g193 (n_174, pi0092);
  and g194 (n2534, n_174, n2533);
  and g195 (n2535, n2532, n2534);
  not g196 (n_176, pi0055);
  and g197 (n2536, n_176, n2535);
  and g198 (n2537, n2531, n2536);
  and g199 (n2538, n2529, n2537);
  and g200 (n2539, n2528, n2538);
  and g201 (n2540, pi0059, n2460);
  not g202 (n_178, n2539);
  and g203 (n2541, n_178, n2540);
  not g204 (n_179, n2537);
  and g205 (n2542, n2460, n_179);
  not g206 (n_180, pi0105);
  not g207 (n_181, n2446);
  and g208 (n2543, n_180, n_181);
  and g209 (n2544, pi0105, n_154);
  not g210 (n_182, n2543);
  not g211 (n_183, n2544);
  and g212 (n2545, n_182, n_183);
  not g213 (n_184, n2545);
  and g214 (n2546, pi0228, n_184);
  and g215 (n2547, pi0137, n2521);
  not g216 (n_185, n2547);
  and g217 (n2548, n2446, n_185);
  and g218 (n2549, n_4, n2512);
  not g219 (n_186, pi0137);
  not g220 (n_187, pi0153);
  and g221 (n2550, n_186, n_187);
  and g222 (n2551, n2549, n2550);
  not g223 (n_188, pi0228);
  not g224 (n_189, n2548);
  and g225 (n2552, n_188, n_189);
  not g226 (n_190, n2551);
  and g227 (n2553, n_190, n2552);
  not g228 (n_191, n2546);
  not g229 (n_192, n2553);
  and g230 (n2554, n_191, n_192);
  not g231 (n_193, n2554);
  and g232 (n2555, n_20, n_193);
  not g233 (n_194, n2555);
  and g234 (n2556, n_23, n_194);
  not g235 (n_195, n2556);
  and g236 (n2557, n_26, n_195);
  not g237 (n_196, n2557);
  and g238 (n2558, n_35, n_196);
  not g239 (n_197, n2558);
  and g240 (n2559, n_36, n_197);
  not g241 (n_198, n2559);
  and g242 (n2560, n_38, n_198);
  and g243 (n2561, n2537, n2560);
  not g244 (n_199, n2542);
  not g245 (n_200, n2561);
  and g246 (n2562, n_199, n_200);
  not g247 (n_201, n2562);
  and g248 (n2563, n_157, n_201);
  and g249 (n2564, pi0056, n2460);
  not g250 (n_202, n2564);
  and g251 (n2565, pi0062, n_202);
  not g252 (n_203, n2563);
  and g253 (n2566, n_203, n2565);
  and g254 (n2567, pi0056, n_201);
  and g255 (n2568, n_172, n_164);
  and g256 (n2569, n_171, n_174);
  and g257 (n2570, n2532, n2569);
  and g258 (n2571, n2568, n2570);
  and g259 (n2572, n2530, n2571);
  not g260 (n_204, n2572);
  and g261 (n2573, n2460, n_204);
  and g262 (n2574, pi0228, n_182);
  and g263 (n2575, n_4, n2523);
  not g264 (n_205, n2575);
  and g265 (n2576, pi0105, n_205);
  not g266 (n_206, n2576);
  and g267 (n2577, n2574, n_206);
  and g268 (n2578, n_188, n2446);
  not g269 (n_207, n2521);
  and g270 (n2579, n_207, n2578);
  not g271 (n_208, n2579);
  and g272 (n2580, n_20, n_208);
  not g273 (n_209, n2577);
  and g274 (n2581, n_209, n2580);
  not g275 (n_210, n2581);
  and g276 (n2582, n_23, n_210);
  not g277 (n_211, n2582);
  and g278 (n2583, n_26, n_211);
  not g279 (n_212, n2583);
  and g280 (n2584, n_35, n_212);
  not g281 (n_213, n2584);
  and g282 (n2585, n_36, n_213);
  and g283 (n2586, n_38, n2572);
  not g284 (n_214, n2585);
  and g285 (n2587, n_214, n2586);
  not g286 (n_215, n2573);
  and g287 (n2588, pi0055, n_215);
  not g288 (n_216, n2587);
  and g289 (n2589, n_216, n2588);
  and g290 (n2590, pi0299, n2460);
  not g291 (n_219, pi0224);
  and g292 (n2591, n_219, pi0833);
  not g293 (n_221, n2591);
  and g294 (n2592, pi0222, n_221);
  not g295 (n_223, pi0223);
  not g296 (n_224, n2592);
  and g297 (n2593, n_223, n_224);
  not g298 (n_225, n2593);
  and g299 (n2594, n2437, n_225);
  and g300 (n2595, pi0224, n_10);
  not g301 (n_226, pi0222);
  not g302 (n_227, n2595);
  and g303 (n2596, n_226, n_227);
  not g304 (n_228, pi0929);
  and g305 (n2597, n_4, n_228);
  and g306 (n2598, n2591, n2597);
  not g307 (n_229, n2596);
  not g308 (n_230, n2598);
  and g309 (n2599, n_229, n_230);
  not g310 (n_231, n2599);
  and g311 (n2600, n_223, n_231);
  not g312 (n_232, n2594);
  not g313 (n_233, n2600);
  and g314 (n2601, n_232, n_233);
  not g315 (n_234, pi0299);
  not g316 (n_235, n2601);
  and g317 (n2602, n_234, n_235);
  and g318 (n2603, n_226, n_219);
  and g319 (n2604, n_223, n2603);
  not g320 (n_236, n2444);
  and g321 (n2605, n_236, n2604);
  not g322 (n_237, n2605);
  and g323 (n2606, n2602, n_237);
  not g324 (n_238, n2590);
  not g325 (n_239, n2606);
  and g326 (n2607, n_238, n_239);
  and g327 (n2608, n_161, n_164);
  and g328 (n2609, n_162, n_172);
  and g329 (n2610, n2608, n2609);
  and g330 (n2611, n2569, n2610);
  not g331 (n_240, n2611);
  and g332 (n2612, n2607, n_240);
  and g333 (n2613, n_154, n2604);
  not g334 (n_241, n2613);
  and g335 (n2614, n_235, n_241);
  not g336 (n_242, n2614);
  and g337 (n2615, n_234, n_242);
  not g338 (n_243, n2528);
  and g339 (n2616, n2460, n_243);
  not g340 (n_244, n2616);
  and g341 (n2617, pi0299, n_244);
  not g342 (n_245, n2615);
  not g343 (n_246, n2617);
  and g344 (n2618, n_245, n_246);
  not g345 (n_247, n2618);
  and g346 (n2619, n_162, n_247);
  and g347 (n2620, n_161, n2568);
  and g348 (n2621, n2569, n2620);
  and g349 (n2622, n2619, n2621);
  not g350 (n_248, n2612);
  not g351 (n_249, n2622);
  and g352 (n2623, n_248, n_249);
  and g353 (n2624, pi0054, n2623);
  and g354 (n2625, n_162, n2608);
  not g355 (n_250, n2607);
  not g356 (n_251, n2625);
  and g357 (n2626, n_250, n_251);
  not g358 (n_252, n2560);
  and g359 (n2627, pi0299, n_252);
  not g360 (n_253, n2627);
  and g361 (n2628, n_245, n_253);
  and g362 (n2629, n2625, n2628);
  not g363 (n_254, n2626);
  not g364 (n_255, n2629);
  and g365 (n2630, n_254, n_255);
  not g366 (n_256, n2630);
  and g367 (n2631, n2533, n_256);
  not g368 (n_257, n2533);
  and g369 (n2632, n_257, n_250);
  not g370 (n_258, n2632);
  and g371 (n2633, pi0092, n_258);
  not g372 (n_259, n2631);
  and g373 (n2634, n_259, n2633);
  and g374 (n2635, pi0087, n_256);
  not g375 (n_260, n2530);
  and g376 (n2636, n_260, n_250);
  and g377 (n2637, pi0095, pi0234);
  not g378 (n_263, pi0152);
  not g379 (n_264, pi0161);
  and g380 (n2638, n_263, n_264);
  not g381 (n_266, pi0166);
  and g382 (n2639, n_266, n2638);
  not g383 (n_268, pi0146);
  not g384 (n_269, n2639);
  and g385 (n2640, n_268, n_269);
  not g386 (n_271, pi0210);
  not g387 (n_272, n2640);
  and g388 (n2641, n_271, n_272);
  not g389 (n_273, n2637);
  and g390 (n2642, n_186, n_273);
  not g391 (n_274, n2641);
  and g392 (n2643, n_274, n2642);
  not g393 (n_275, n2643);
  and g394 (n2644, n_152, n_275);
  not g395 (n_276, n2644);
  and g396 (n2645, n_4, n_276);
  not g397 (n_277, n2645);
  and g398 (n2646, pi0105, n_277);
  not g399 (n_278, n2646);
  and g400 (n2647, n2574, n_278);
  and g401 (n2648, n2547, n2640);
  and g402 (n2649, n_186, pi0210);
  not g403 (n_280, pi0252);
  not g408 (n_282, n2648);
  and g409 (n2653, n2446, n_282);
  not g410 (n_283, n2652);
  and g411 (n2654, n_283, n2653);
  and g412 (n2655, pi0252, n_272);
  not g413 (n_284, n2655);
  and g414 (n2656, n_274, n_284);
  and g415 (n2657, n2551, n2656);
  not g416 (n_285, n2654);
  not g417 (n_286, n2657);
  and g418 (n2658, n_285, n_286);
  not g419 (n_287, n2658);
  and g420 (n2659, n_188, n_287);
  not g421 (n_288, n2659);
  and g422 (n2660, n_20, n_288);
  not g423 (n_289, n2647);
  and g424 (n2661, n_289, n2660);
  not g425 (n_290, n2661);
  and g426 (n2662, n_23, n_290);
  not g427 (n_291, n2662);
  and g428 (n2663, n_26, n_291);
  not g429 (n_292, n2663);
  and g430 (n2664, n_35, n_292);
  not g431 (n_293, n2664);
  and g432 (n2665, n_36, n_293);
  not g433 (n_294, n2665);
  and g434 (n2666, n_38, n_294);
  not g435 (n_295, n2666);
  and g436 (n2667, pi0299, n_295);
  not g437 (n_298, pi0144);
  not g438 (n_299, pi0174);
  and g439 (n2668, n_298, n_299);
  not g440 (n_301, pi0189);
  and g441 (n2669, n_301, n2668);
  not g442 (n_302, n2669);
  and g443 (n2670, n_223, n_302);
  not g444 (n_305, pi0198);
  and g445 (n2671, pi0142, n_305);
  not g446 (n_306, n2671);
  and g447 (n2672, n_186, n_306);
  not g448 (n_307, n2672);
  and g449 (n2673, n_152, n_307);
  not g450 (n_308, n2673);
  and g451 (n2674, n2444, n_308);
  not g452 (n_309, n2674);
  and g453 (n2675, n2670, n_309);
  and g454 (n2676, n_148, n_4);
  and g455 (n2677, n_186, pi0198);
  not g456 (n_310, n2677);
  and g457 (n2678, n2521, n_310);
  not g458 (n_311, n2678);
  and g459 (n2679, n2676, n_311);
  and g460 (n2680, n_223, n2669);
  and g461 (n2681, pi0234, n_4);
  and g462 (n2682, n_144, n2677);
  not g463 (n_312, n2682);
  and g464 (n2683, n_147, n_312);
  not g465 (n_313, n2683);
  and g466 (n2684, n2681, n_313);
  not g467 (n_314, n2679);
  and g468 (n2685, n_314, n2680);
  not g469 (n_315, n2684);
  and g470 (n2686, n_315, n2685);
  not g471 (n_316, n2675);
  not g472 (n_317, n2686);
  and g473 (n2687, n_316, n_317);
  not g474 (n_318, n2687);
  and g475 (n2688, n2603, n_318);
  not g476 (n_319, n2688);
  and g477 (n2689, n_235, n_319);
  not g478 (n_320, n2689);
  and g479 (n2690, n_234, n_320);
  not g480 (n_321, n2690);
  and g481 (n2691, n2530, n_321);
  not g482 (n_322, n2667);
  and g483 (n2692, n_322, n2691);
  not g484 (n_323, n2636);
  and g485 (n2693, pi0100, n_323);
  not g486 (n_324, n2692);
  and g487 (n2694, n_324, n2693);
  and g488 (n2695, pi0039, n2607);
  not g489 (n_325, n2695);
  and g490 (n2696, pi0038, n_325);
  not g491 (n_326, n2619);
  and g492 (n2697, n_326, n2696);
  not g493 (n_327, n2628);
  and g494 (n2698, pi0039, n_327);
  and g495 (n2699, n2491, n2499);
  and g496 (n2700, n_42, n_109);
  and g497 (n2701, n_108, n2700);
  and g498 (n2702, n2493, n2701);
  and g499 (n2703, n2699, n2702);
  and g500 (n2704, n_43, n_131);
  and g501 (n2705, n_139, n_135);
  and g502 (n2706, n_130, n_138);
  and g503 (n2707, n2705, n2706);
  and g504 (n2708, n2704, n2707);
  and g505 (n2709, n2703, n2708);
  and g506 (n2710, n2517, n2709);
  and g507 (n2711, pi0225, n2710);
  not g508 (n_329, n2711);
  and g509 (n2712, pi0032, n_329);
  not g510 (n_330, n2712);
  and g511 (n2713, n_144, n_330);
  and g512 (n2714, n_127, n2493);
  and g513 (n2715, n2492, n2496);
  and g514 (n2716, n2714, n2715);
  and g515 (n2717, n_42, n2716);
  and g516 (n2718, pi0060, n2491);
  not g517 (n_331, n2718);
  and g518 (n2719, n_116, n_331);
  and g519 (n2720, n_119, n_125);
  and g520 (n2721, n_117, n2491);
  not g521 (n_332, n2721);
  and g522 (n2722, pi0053, n_332);
  not g523 (n_333, n2722);
  and g524 (n2723, n2720, n_333);
  not g525 (n_334, n2719);
  and g526 (n2724, n_334, n2723);
  and g527 (n2725, n2704, n2717);
  and g528 (n2726, n2724, n2725);
  not g529 (n_335, n2726);
  and g530 (n2727, n_130, n_335);
  and g531 (n2728, n_131, n2503);
  not g532 (n_336, n2728);
  and g533 (n2729, pi0035, n_336);
  and g534 (n2730, pi0035, n2728);
  not g535 (n_337, pi0225);
  and g536 (n2731, n_337, n2730);
  not g537 (n_338, n2731);
  and g538 (n2732, n_139, n_338);
  and g539 (n2733, n_138, n2732);
  not g540 (n_339, n2729);
  and g541 (n2734, n_339, n2733);
  not g542 (n_340, n2727);
  and g543 (n2735, n_340, n2734);
  and g544 (n2736, n_143, n2506);
  and g545 (n2737, n2735, n2736);
  not g546 (n_341, n2737);
  and g547 (n2738, n_142, n_341);
  not g548 (n_342, n2738);
  and g549 (n2739, n2713, n_342);
  not g550 (n_343, n2739);
  and g551 (n2740, n_186, n_343);
  not g552 (n_344, n2511);
  and g553 (n2741, pi0095, n_344);
  not g554 (n_345, n2741);
  and g555 (n2742, n_145, n_345);
  and g556 (n2743, pi0040, n2509);
  not g557 (n_346, n2743);
  and g558 (n2744, n_142, n_346);
  not g559 (n_347, n2709);
  and g560 (n2745, pi0072, n_347);
  not g561 (n_348, n2745);
  and g562 (n2746, n_143, n_348);
  not g563 (n_349, n2515);
  and g564 (n2747, pi0051, n_349);
  not g565 (n_350, n2747);
  and g566 (n2748, n_135, n_350);
  and g567 (n2749, n_138, pi0070);
  not g568 (n_351, n2749);
  and g569 (n2750, n2748, n_351);
  and g570 (n2751, n_339, n_338);
  and g571 (n2752, pi0093, n2503);
  not g572 (n_352, n2752);
  and g573 (n2753, n_130, n_352);
  and g574 (n2754, n_108, n2500);
  and g575 (n2755, n2491, n2754);
  and g576 (n2756, pi0091, n2755);
  not g577 (n_353, n2756);
  and g578 (n2757, n2461, n_353);
  and g579 (n2758, n_112, n2699);
  not g580 (n_354, n2758);
  and g581 (n2759, pi0110, n_354);
  and g582 (n2760, pi0047, n2491);
  and g583 (n2761, n2500, n2760);
  not g584 (n_355, n2761);
  and g585 (n2762, pi0047, n_355);
  not g586 (n_356, n2762);
  and g587 (n2763, n_109, n_356);
  not g588 (n_357, n2759);
  and g589 (n2764, n_357, n2763);
  and g590 (n2765, n_108, n_113);
  not g591 (n_358, n2699);
  and g592 (n2766, pi0109, n_358);
  and g593 (n2767, n_53, n2490);
  and g594 (n2768, n2462, n2767);
  and g595 (n2769, n_51, n2494);
  and g596 (n2770, n_49, n2769);
  and g597 (n2771, n2720, n2770);
  and g598 (n2772, n2768, n2771);
  and g599 (n2773, n_122, n2772);
  not g600 (n_359, n2773);
  and g601 (n2774, pi0108, n_359);
  not g602 (n_360, n2774);
  and g603 (n2775, n_127, n_360);
  not g604 (n_361, n2772);
  and g605 (n2776, pi0097, n_361);
  and g606 (n2777, n2463, n2767);
  and g607 (n2778, n2769, n2777);
  and g608 (n2779, n_119, pi0094);
  and g609 (n2780, n2778, n2779);
  not g610 (n_362, n2780);
  and g611 (n2781, n_122, n_362);
  not g612 (n_363, n2778);
  and g613 (n2782, pi0086, n_363);
  not g614 (n_364, n2782);
  and g615 (n2783, n_125, n_364);
  and g616 (n2784, pi0077, n2768);
  not g617 (n_365, n2784);
  and g618 (n2785, n_51, n_365);
  not g619 (n_366, n2489);
  and g620 (n2786, pi0081, n_366);
  not g621 (n_367, n2490);
  and g622 (n2787, pi0102, n_367);
  not g623 (n_368, n2786);
  not g624 (n_369, n2787);
  and g625 (n2788, n_368, n_369);
  not g626 (n_370, n2488);
  and g627 (n2789, pi0064, n_370);
  not g628 (n_371, n2485);
  and g629 (n2790, pi0071, n_371);
  not g630 (n_372, n2790);
  and g631 (n2791, n_56, n_372);
  and g632 (n2792, n_64, n2483);
  not g633 (n_373, n2792);
  and g634 (n2793, pi0069, n_373);
  not g635 (n_374, n2484);
  and g636 (n2794, pi0083, n_374);
  not g637 (n_375, n2794);
  and g638 (n2795, n_61, n_375);
  not g639 (n_376, n2793);
  and g640 (n2796, n_376, n2795);
  and g641 (n2797, n_65, n_60);
  not g642 (n_377, n2483);
  and g643 (n2798, pi0067, n_377);
  and g644 (n2799, n2469, n2477);
  and g645 (n2800, n_91, n2799);
  and g646 (n2801, n_90, n2800);
  and g647 (n2802, n2479, n2801);
  not g648 (n_378, n2802);
  and g649 (n2803, pi0036, n_378);
  and g650 (n2804, n_97, n_64);
  and g651 (n2805, n_90, n_95);
  and g652 (n2806, pi0082, n2805);
  and g653 (n2807, n2800, n2806);
  not g654 (n_379, n2801);
  and g655 (n2808, pi0111, n_379);
  not g656 (n_380, n2808);
  and g657 (n2809, n_94, n_380);
  not g658 (n_381, n2800);
  and g659 (n2810, pi0068, n_381);
  not g660 (n_382, n2799);
  and g661 (n2811, pi0084, n_382);
  not g662 (n_383, n2475);
  and g663 (n2812, pi0104, n_383);
  and g664 (n2813, pi0085, pi0106);
  not g665 (n_384, n2813);
  and g666 (n2814, n2470, n_384);
  and g667 (n2815, pi0061, pi0076);
  not g668 (n_385, n2815);
  and g669 (n2816, n2471, n_385);
  not g670 (n_386, n2814);
  not g671 (n_387, n2816);
  and g672 (n2817, n_386, n_387);
  not g673 (n_388, n2817);
  and g674 (n2818, n_79, n_388);
  not g675 (n_389, n2472);
  not g676 (n_390, n2818);
  and g677 (n2819, n_389, n_390);
  not g678 (n_391, n2473);
  and g679 (n2820, pi0089, n_391);
  not g680 (n_392, n2820);
  and g681 (n2821, n_83, n_392);
  not g682 (n_393, n2819);
  and g683 (n2822, n_393, n2821);
  not g684 (n_394, n2474);
  not g685 (n_395, n2822);
  and g686 (n2823, n_394, n_395);
  not g687 (n_396, n2812);
  and g688 (n2824, n_87, n_396);
  not g689 (n_397, n2823);
  and g690 (n2825, n_397, n2824);
  not g691 (n_398, n2476);
  not g692 (n_399, n2825);
  and g693 (n2826, n_398, n_399);
  not g694 (n_400, n2477);
  not g695 (n_401, n2826);
  and g696 (n2827, n_400, n_401);
  not g697 (n_402, n2827);
  and g698 (n2828, n2469, n_402);
  and g699 (n2829, pi0066, pi0073);
  not g700 (n_403, n2469);
  and g701 (n2830, n_403, n_400);
  not g702 (n_404, n2829);
  not g703 (n_405, n2830);
  and g704 (n2831, n_404, n_405);
  not g705 (n_406, n2828);
  and g706 (n2832, n_406, n2831);
  not g707 (n_407, n2832);
  and g708 (n2833, n_91, n_407);
  not g709 (n_408, n2811);
  not g710 (n_409, n2833);
  and g711 (n2834, n_408, n_409);
  not g712 (n_410, n2834);
  and g713 (n2835, n2805, n_410);
  not g714 (n_411, n2810);
  and g715 (n2836, n2809, n_411);
  not g716 (n_412, n2835);
  and g717 (n2837, n_412, n2836);
  not g718 (n_413, n2807);
  and g719 (n2838, n2804, n_413);
  not g720 (n_414, n2837);
  and g721 (n2839, n_414, n2838);
  not g722 (n_415, n2798);
  not g723 (n_416, n2803);
  and g724 (n2840, n_415, n_416);
  not g725 (n_417, n2839);
  and g726 (n2841, n_417, n2840);
  not g727 (n_418, n2841);
  and g728 (n2842, n2797, n_418);
  not g729 (n_419, n2842);
  and g730 (n2843, n2796, n_419);
  and g731 (n2844, pi0103, n2797);
  and g732 (n2845, n2792, n2844);
  not g733 (n_420, n2845);
  and g734 (n2846, n_57, n_420);
  not g735 (n_421, n2843);
  and g736 (n2847, n_421, n2846);
  not g737 (n_422, n2847);
  and g738 (n2848, n2791, n_422);
  not g739 (n_423, n2848);
  and g740 (n2849, n_101, n_423);
  and g741 (n2850, pi0065, n_57);
  and g742 (n2851, n2485, n2850);
  not g743 (n_424, n2851);
  and g744 (n2852, n2849, n_424);
  not g745 (n_425, n2486);
  and g746 (n2853, pi0107, n_425);
  not g747 (n_426, n2853);
  and g748 (n2854, n_100, n_426);
  not g749 (n_427, n2852);
  and g750 (n2855, n_427, n2854);
  not g751 (n_428, n2855);
  and g752 (n2856, n_103, n_428);
  not g753 (n_429, n2789);
  not g754 (n_430, n2856);
  and g755 (n2857, n_429, n_430);
  and g756 (n2858, n_105, n_53);
  not g757 (n_431, n2857);
  and g758 (n2859, n_431, n2858);
  not g759 (n_432, n2849);
  and g760 (n2860, n_432, n2854);
  and g761 (n2861, pi0063, n_101);
  and g762 (n2862, n2486, n2861);
  not g763 (n_433, n2862);
  and g764 (n2863, n_103, n_433);
  not g765 (n_434, n2860);
  and g766 (n2864, n_434, n2863);
  not g767 (n_435, n2864);
  and g768 (n2865, n_429, n_435);
  not g769 (n_436, n2865);
  and g770 (n2866, n2859, n_436);
  not g771 (n_437, n2866);
  and g772 (n2867, n2788, n_437);
  not g773 (n_438, n2867);
  and g774 (n2868, n2462, n_438);
  not g775 (n_439, n2767);
  and g776 (n2869, pi0098, n_439);
  and g777 (n2870, n_47, n2767);
  not g778 (n_440, n2870);
  and g779 (n2871, pi0088, n_440);
  not g780 (n_441, n2869);
  and g781 (n2872, n_49, n_441);
  not g782 (n_442, n2871);
  and g783 (n2873, n_442, n2872);
  not g784 (n_443, n2868);
  and g785 (n2874, n_443, n2873);
  not g786 (n_444, n2874);
  and g787 (n2875, n2785, n_444);
  not g788 (n_445, n2777);
  and g789 (n2876, pi0050, n_445);
  not g790 (n_446, n2876);
  and g791 (n2877, n_117, n_446);
  not g792 (n_447, n2875);
  and g793 (n2878, n_447, n2877);
  not g794 (n_448, n2878);
  and g795 (n2879, n2719, n_448);
  not g796 (n_449, n2879);
  and g797 (n2880, n_333, n_449);
  not g798 (n_450, n2880);
  and g799 (n2881, n_119, n_450);
  not g800 (n_451, n2881);
  and g801 (n2882, n2783, n_451);
  not g802 (n_452, n2882);
  and g803 (n2883, n2781, n_452);
  not g804 (n_453, n2776);
  not g805 (n_454, n2883);
  and g806 (n2884, n_453, n_454);
  not g807 (n_455, n2884);
  and g808 (n2885, n_123, n_455);
  not g809 (n_456, n2885);
  and g810 (n2886, n2775, n_456);
  and g811 (n2887, pi0046, n2496);
  and g812 (n2888, n2772, n2887);
  not g813 (n_457, n2888);
  and g814 (n2889, n_112, n_457);
  not g815 (n_458, n2886);
  and g816 (n2890, n_458, n2889);
  not g817 (n_459, n2766);
  not g818 (n_460, n2890);
  and g819 (n2891, n_459, n_460);
  not g820 (n_461, n2891);
  and g821 (n2892, n2765, n_461);
  not g822 (n_462, n2892);
  and g823 (n2893, n2764, n_462);
  not g824 (n_463, n2893);
  and g825 (n2894, n2757, n_463);
  not g826 (n_464, n2502);
  and g827 (n2895, pi0058, n_464);
  not g828 (n_465, n2703);
  and g829 (n2896, pi0090, n_465);
  not g830 (n_466, n2896);
  and g831 (n2897, n_131, n_466);
  not g832 (n_467, n2895);
  and g833 (n2898, n_467, n2897);
  not g834 (n_468, n2894);
  and g835 (n2899, n_468, n2898);
  not g836 (n_469, n2899);
  and g837 (n2900, n2753, n_469);
  not g838 (n_470, n2900);
  and g839 (n2901, n2751, n_470);
  not g840 (n_471, n2901);
  and g841 (n2902, n_138, n_471);
  not g842 (n_472, n2902);
  and g843 (n2903, n2750, n_472);
  not g844 (n_473, n2903);
  and g845 (n2904, n_134, n_473);
  not g846 (n_474, n2904);
  and g847 (n2905, n2746, n_474);
  not g848 (n_475, n2905);
  and g849 (n2906, n2744, n_475);
  not g850 (n_476, n2906);
  and g851 (n2907, n_330, n_476);
  not g852 (n_477, n2907);
  and g853 (n2908, n_144, n_477);
  not g854 (n_478, n2908);
  and g855 (n2909, n2742, n_478);
  not g856 (n_479, n2909);
  and g857 (n2910, pi0137, n_479);
  not g858 (n_480, n2740);
  not g859 (n_481, n2910);
  and g860 (n2911, n_480, n_481);
  not g861 (n_482, n2911);
  and g862 (n2912, pi0210, n_482);
  and g863 (n2913, n_138, n_134);
  and g864 (n2914, pi0841, n2503);
  and g865 (n2915, n_131, n2914);
  and g866 (n2916, n2913, n2915);
  not g871 (n_484, n2920);
  and g872 (n2921, pi0032, n_484);
  not g873 (n_485, n2921);
  and g874 (n2922, n_144, n_485);
  not g875 (n_486, pi0833);
  and g876 (n2923, n_486, pi0957);
  not g877 (n_489, n2923);
  and g878 (n2924, pi1091, n_489);
  and g879 (n2925, pi0829, pi0950);
  and g880 (n2926, pi1092, pi1093);
  and g881 (n2927, n2925, n2926);
  and g882 (n2928, n2924, n2927);
  not g883 (n_494, n2928);
  and g884 (n2929, n_340, n_494);
  and g885 (n2930, pi1091, pi1093);
  and g886 (n2931, n_489, n2930);
  and g887 (n2932, pi0950, pi1092);
  and g888 (n2933, pi0829, n2932);
  and g889 (n2934, n_127, n_112);
  and g890 (n2935, n2492, n2934);
  and g891 (n2936, n_123, n_453);
  and g892 (n2937, n_113, n2936);
  and g893 (n2938, n_131, n2461);
  not g894 (n_495, n2724);
  and g895 (n2939, n_122, n_495);
  not g900 (n_497, n2942);
  and g901 (n2943, n_130, n_497);
  and g902 (n2944, n2931, n2933);
  not g903 (n_498, n2943);
  and g904 (n2945, n_498, n2944);
  not g905 (n_499, n2929);
  not g906 (n_500, n2945);
  and g907 (n2946, n_499, n_500);
  and g908 (n2947, n2734, n2736);
  not g909 (n_501, n2946);
  and g910 (n2948, n_501, n2947);
  not g911 (n_502, n2948);
  and g912 (n2949, n_142, n_502);
  not g913 (n_503, n2949);
  and g914 (n2950, n2922, n_503);
  not g915 (n_504, n2950);
  and g916 (n2951, n_186, n_504);
  and g917 (n2952, n_476, n_485);
  not g918 (n_505, n2952);
  and g919 (n2953, n_144, n_505);
  not g920 (n_506, n2953);
  and g921 (n2954, n2742, n_506);
  not g922 (n_507, n2954);
  and g923 (n2955, pi0137, n_507);
  not g924 (n_508, n2951);
  not g925 (n_509, n2955);
  and g926 (n2956, n_508, n_509);
  not g927 (n_510, n2956);
  and g928 (n2957, n_271, n_510);
  not g929 (n_511, n2912);
  not g930 (n_512, n2957);
  and g931 (n2958, n_511, n_512);
  and g932 (n2959, n_148, n2958);
  not g933 (n_513, n2735);
  and g934 (n2960, n_135, n_513);
  and g935 (n2961, n_130, n_139);
  and g936 (n2962, n_138, n2961);
  and g937 (n2963, n_109, n2938);
  and g938 (n2964, n2962, n2963);
  and g939 (n2965, n2755, n2964);
  not g940 (n_514, n2965);
  and g941 (n2966, pi0096, n_514);
  not g942 (n_515, n2966);
  and g943 (n2967, n2517, n_515);
  not g944 (n_516, n2960);
  and g945 (n2968, n_516, n2967);
  not g946 (n_517, n2968);
  and g947 (n2969, n_142, n_517);
  not g948 (n_518, n2969);
  and g949 (n2970, n2713, n_518);
  not g950 (n_519, n2970);
  and g951 (n2971, n_145, n_519);
  and g952 (n2972, n_186, n2971);
  and g953 (n2973, pi0096, n2965);
  and g954 (n2974, n_143, n2913);
  and g955 (n2975, n2505, n2974);
  and g956 (n2976, n2973, n2975);
  not g957 (n_520, n2976);
  and g958 (n2977, n2906, n_520);
  not g959 (n_521, n2977);
  and g960 (n2978, n_330, n_521);
  not g961 (n_522, n2978);
  and g962 (n2979, n_144, n_522);
  and g963 (n2980, pi0479, n2741);
  not g964 (n_523, n2979);
  not g965 (n_524, n2980);
  and g966 (n2981, n_523, n_524);
  not g967 (n_525, n2981);
  and g968 (n2982, pi0137, n_525);
  not g969 (n_526, n2972);
  not g970 (n_527, n2982);
  and g971 (n2983, n_526, n_527);
  not g972 (n_528, n2983);
  and g973 (n2984, pi0210, n_528);
  and g974 (n2985, n_485, n_521);
  not g975 (n_529, n2985);
  and g976 (n2986, n_144, n_529);
  not g977 (n_530, n2986);
  and g978 (n2987, n_524, n_530);
  not g979 (n_531, n2987);
  and g980 (n2988, pi0137, n_531);
  and g981 (n2989, pi0095, pi0479);
  and g982 (n2990, n_485, n_518);
  not g983 (n_532, n2990);
  and g984 (n2991, n_144, n_532);
  not g985 (n_533, n2989);
  not g986 (n_534, n2991);
  and g987 (n2992, n_533, n_534);
  not g988 (n_535, n2992);
  and g989 (n2993, n_186, n_535);
  not g990 (n_536, n2988);
  not g991 (n_537, n2993);
  and g992 (n2994, n_536, n_537);
  not g993 (n_538, n2924);
  and g994 (n2995, n_538, n2994);
  and g995 (n2996, n2734, n_498);
  not g996 (n_539, n2996);
  and g997 (n2997, n_135, n_539);
  not g998 (n_540, n2997);
  and g999 (n2998, n2967, n_540);
  not g1000 (n_541, n2998);
  and g1001 (n2999, n_142, n_541);
  not g1002 (n_542, n2999);
  and g1003 (n3000, n_485, n_542);
  not g1004 (n_543, n3000);
  and g1005 (n3001, n_144, n_543);
  and g1006 (n3002, n2927, n_533);
  not g1007 (n_544, n3001);
  and g1008 (n3003, n_544, n3002);
  not g1009 (n_545, n2927);
  and g1010 (n3004, n_545, n2992);
  not g1011 (n_546, n3003);
  and g1012 (n3005, n_186, n_546);
  not g1013 (n_547, n3004);
  and g1014 (n3006, n_547, n3005);
  not g1015 (n_548, n3006);
  and g1016 (n3007, n2924, n_548);
  and g1017 (n3008, n_536, n3007);
  not g1018 (n_549, n2995);
  not g1019 (n_550, n3008);
  and g1020 (n3009, n_549, n_550);
  and g1021 (n3010, n_271, n3009);
  not g1022 (n_551, n2984);
  not g1023 (n_552, n3010);
  and g1024 (n3011, n_551, n_552);
  and g1025 (n3012, pi0234, n3011);
  not g1026 (n_553, n2959);
  and g1027 (n3013, n_4, n_553);
  not g1028 (n_554, n3012);
  and g1029 (n3014, n_554, n3013);
  not g1030 (n_555, n3014);
  and g1031 (n3015, n2639, n_555);
  and g1032 (n3016, pi0146, n3011);
  not g1033 (n_556, n2994);
  and g1034 (n3017, n_271, n_556);
  and g1035 (n3018, n_268, n_551);
  not g1036 (n_557, n3017);
  and g1037 (n3019, n_557, n3018);
  not g1038 (n_558, n3019);
  and g1039 (n3020, n2681, n_558);
  not g1040 (n_559, n3016);
  and g1041 (n3021, n_559, n3020);
  and g1042 (n3022, pi0146, n2958);
  and g1043 (n3023, n_342, n2922);
  not g1044 (n_560, n3023);
  and g1045 (n3024, n_186, n_560);
  not g1046 (n_561, n3024);
  and g1047 (n3025, n_509, n_561);
  not g1048 (n_562, n3025);
  and g1049 (n3026, n_271, n_562);
  and g1050 (n3027, n_268, n_511);
  not g1051 (n_563, n3026);
  and g1052 (n3028, n_563, n3027);
  not g1053 (n_564, n3022);
  and g1054 (n3029, n2676, n_564);
  not g1055 (n_565, n3028);
  and g1056 (n3030, n_565, n3029);
  not g1057 (n_566, n3030);
  and g1058 (n3031, n_269, n_566);
  not g1059 (n_567, n3021);
  and g1060 (n3032, n_567, n3031);
  not g1061 (n_568, n3015);
  not g1062 (n_569, n3032);
  and g1063 (n3033, n_568, n_569);
  not g1064 (n_570, n3033);
  and g1065 (n3034, pi0105, n_570);
  not g1066 (n_571, n3034);
  and g1067 (n3035, n_182, n_571);
  not g1068 (n_572, n3035);
  and g1069 (n3036, pi0228, n_572);
  and g1070 (n3037, n_112, n_458);
  not g1071 (n_573, n3037);
  and g1072 (n3038, n_459, n_573);
  not g1073 (n_574, n3038);
  and g1074 (n3039, n2765, n_574);
  not g1075 (n_575, n3039);
  and g1076 (n3040, n2764, n_575);
  not g1077 (n_576, n3040);
  and g1078 (n3041, n2757, n_576);
  not g1079 (n_577, n3041);
  and g1080 (n3042, n2898, n_577);
  not g1081 (n_578, n3042);
  and g1082 (n3043, n2753, n_578);
  not g1083 (n_579, n3043);
  and g1084 (n3044, n2751, n_579);
  not g1085 (n_580, n3044);
  and g1086 (n3045, n_138, n_580);
  not g1087 (n_581, n3045);
  and g1088 (n3046, n2750, n_581);
  not g1089 (n_582, n3046);
  and g1090 (n3047, n_134, n_582);
  not g1091 (n_583, n3047);
  and g1092 (n3048, n2746, n_583);
  not g1093 (n_584, n3048);
  and g1094 (n3049, n2744, n_584);
  not g1095 (n_585, n3049);
  and g1096 (n3050, n_485, n_585);
  not g1097 (n_586, n3050);
  and g1098 (n3051, n_144, n_586);
  not g1099 (n_587, n3051);
  and g1100 (n3052, n2742, n_587);
  not g1101 (n_588, n3052);
  and g1102 (n3053, pi0137, n_588);
  and g1103 (n3054, n2640, n3024);
  and g1104 (n3055, n_272, n2951);
  and g1112 (n3060, n_330, n_585);
  not g1113 (n_592, n3060);
  and g1114 (n3061, n_144, n_592);
  not g1115 (n_593, n3061);
  and g1116 (n3062, n2742, n_593);
  not g1117 (n_594, n3062);
  and g1118 (n3063, pi0137, n_594);
  and g1119 (n3064, pi0210, n_480);
  not g1120 (n_595, n3063);
  and g1121 (n3065, n_595, n3064);
  and g1122 (n3066, n_520, n3049);
  not g1123 (n_596, n3066);
  and g1124 (n3067, n_485, n_596);
  not g1125 (n_597, n3067);
  and g1126 (n3068, n_144, n_597);
  not g1127 (n_598, n3068);
  and g1128 (n3069, n_345, n_598);
  not g1129 (n_599, n3069);
  and g1130 (n3070, pi0137, n_599);
  and g1131 (n3071, n_272, n2924);
  and g1132 (n3072, n_547, n3071);
  and g1133 (n3073, n_345, n2992);
  not g1134 (n_600, n3072);
  and g1135 (n3074, n_600, n3073);
  and g1136 (n3075, n_345, n3071);
  and g1137 (n3076, n3003, n3075);
  not g1138 (n_601, n3076);
  and g1139 (n3077, n_186, n_601);
  not g1140 (n_602, n3074);
  and g1141 (n3078, n_602, n3077);
  not g1142 (n_603, n3070);
  not g1143 (n_604, n3078);
  and g1144 (n3079, n_603, n_604);
  not g1145 (n_605, n3079);
  and g1146 (n3080, n_271, n_605);
  not g1147 (n_606, n3080);
  and g1148 (n3081, pi0234, n_606);
  not g1149 (n_607, n3059);
  not g1150 (n_608, n3065);
  and g1151 (n3082, n_607, n_608);
  not g1152 (n_609, n3081);
  and g1153 (n3083, n_609, n3082);
  and g1154 (n3084, n_186, n_345);
  not g1155 (n_610, n2971);
  and g1156 (n3085, n_610, n3084);
  and g1157 (n3086, n_330, n_596);
  not g1158 (n_611, n3086);
  and g1159 (n3087, n_144, n_611);
  and g1160 (n3088, pi0137, n_345);
  not g1161 (n_612, n3087);
  and g1162 (n3089, n_612, n3088);
  not g1168 (n_615, n3083);
  not g1169 (n_616, n3092);
  and g1170 (n3093, n_615, n_616);
  not g1171 (n_617, n3093);
  and g1172 (n3094, n2446, n_617);
  and g1173 (n3095, pi0225, pi0841);
  not g1174 (n_618, n3095);
  and g1175 (n3096, n2710, n_618);
  not g1176 (n_619, n3096);
  and g1177 (n3097, pi0032, n_619);
  not g1178 (n_620, n3097);
  and g1179 (n3098, n_144, n_620);
  not g1180 (n_621, n2505);
  and g1181 (n3099, pi0070, n_621);
  not g1182 (n_622, n3099);
  and g1183 (n3100, n2516, n_622);
  and g1184 (n3101, n2517, n3100);
  not g1185 (n_623, n2732);
  and g1186 (n3102, n_623, n3101);
  not g1187 (n_624, n3102);
  and g1188 (n3103, n_142, n_624);
  not g1189 (n_625, n3103);
  and g1190 (n3104, n3098, n_625);
  not g1191 (n_626, n3104);
  and g1192 (n3105, pi0137, n_626);
  not g1193 (n_627, n2503);
  and g1194 (n3106, pi0093, n_627);
  not g1195 (n_628, n3106);
  and g1196 (n3107, n_130, n_628);
  and g1197 (n3108, n_467, n_466);
  and g1198 (n3109, n_116, n2878);
  not g1199 (n_629, n3109);
  and g1200 (n3110, n_119, n_629);
  not g1201 (n_630, n3110);
  and g1202 (n3111, n2783, n_630);
  not g1203 (n_631, n3111);
  and g1204 (n3112, n2781, n_631);
  not g1205 (n_632, n3112);
  and g1206 (n3113, n_453, n_632);
  not g1207 (n_633, n3113);
  and g1208 (n3114, n_123, n_633);
  not g1209 (n_634, n3114);
  and g1210 (n3115, n2775, n_634);
  not g1211 (n_635, n3115);
  and g1212 (n3116, n_112, n_635);
  not g1213 (n_636, n3116);
  and g1214 (n3117, n_459, n_636);
  not g1215 (n_637, n3117);
  and g1216 (n3118, n2765, n_637);
  not g1217 (n_638, n3118);
  and g1218 (n3119, n2764, n_638);
  not g1219 (n_639, n3119);
  and g1220 (n3120, n2757, n_639);
  not g1221 (n_640, n3120);
  and g1222 (n3121, n3108, n_640);
  not g1223 (n_641, n3121);
  and g1224 (n3122, n_131, n_641);
  not g1225 (n_642, n3122);
  and g1226 (n3123, n3107, n_642);
  not g1227 (n_643, n3123);
  and g1228 (n3124, n2733, n_643);
  and g1229 (n3125, n2748, n_622);
  not g1230 (n_644, n3124);
  and g1231 (n3126, n_644, n3125);
  not g1232 (n_645, n3126);
  and g1233 (n3127, n_134, n_645);
  not g1234 (n_646, n3127);
  and g1235 (n3128, n2746, n_646);
  not g1236 (n_647, n3128);
  and g1237 (n3129, n2744, n_647);
  and g1238 (n3130, n_494, n3129);
  and g1239 (n3131, n2744, n2928);
  and g1240 (n3132, n_122, n_632);
  not g1241 (n_648, n3132);
  and g1242 (n3133, n_123, n_648);
  not g1243 (n_649, n3133);
  and g1244 (n3134, n2775, n_649);
  not g1245 (n_650, n3134);
  and g1246 (n3135, n_112, n_650);
  not g1247 (n_651, n3135);
  and g1248 (n3136, n_459, n_651);
  not g1249 (n_652, n3136);
  and g1250 (n3137, n2765, n_652);
  not g1251 (n_653, n3137);
  and g1252 (n3138, n2764, n_653);
  not g1253 (n_654, n3138);
  and g1254 (n3139, n2757, n_654);
  not g1255 (n_655, n3139);
  and g1256 (n3140, n3108, n_655);
  not g1257 (n_656, n3140);
  and g1258 (n3141, n_131, n_656);
  not g1259 (n_657, n3141);
  and g1260 (n3142, n3107, n_657);
  not g1261 (n_658, n3142);
  and g1262 (n3143, n2733, n_658);
  not g1263 (n_659, n3143);
  and g1264 (n3144, n3125, n_659);
  not g1265 (n_660, n3144);
  and g1266 (n3145, n_134, n_660);
  not g1267 (n_661, n3145);
  and g1268 (n3146, n2746, n_661);
  not g1269 (n_662, n3146);
  and g1270 (n3147, n3131, n_662);
  not g1271 (n_663, n3147);
  and g1272 (n3148, n_620, n_663);
  not g1273 (n_664, n3130);
  and g1274 (n3149, n_664, n3148);
  not g1275 (n_665, n3149);
  and g1276 (n3150, n_144, n_665);
  not g1277 (n_666, n3150);
  and g1278 (n3151, n2742, n_666);
  not g1279 (n_667, n3151);
  and g1280 (n3152, n_186, n_667);
  not g1281 (n_668, n3105);
  not g1282 (n_669, n3152);
  and g1283 (n3153, n_668, n_669);
  not g1284 (n_670, n3153);
  and g1285 (n3154, n_271, n_670);
  and g1286 (n3155, n_337, n2710);
  not g1287 (n_671, n3155);
  and g1288 (n3156, pi0032, n_671);
  not g1289 (n_672, n3156);
  and g1290 (n3157, n_144, n_672);
  and g1291 (n3158, pi0137, n3157);
  and g1292 (n3159, n_625, n3158);
  not g1293 (n_673, n3129);
  and g1294 (n3160, n_673, n_672);
  not g1295 (n_674, n3160);
  and g1296 (n3161, n_144, n_674);
  and g1297 (n3162, n_186, n2742);
  not g1298 (n_675, n3161);
  and g1299 (n3163, n_675, n3162);
  not g1300 (n_676, n3159);
  and g1301 (n3164, pi0210, n_676);
  not g1302 (n_677, n3163);
  and g1303 (n3165, n_677, n3164);
  not g1304 (n_678, n3165);
  and g1305 (n3166, n2681, n_678);
  not g1306 (n_679, n3154);
  and g1307 (n3167, n_679, n3166);
  not g1308 (n_680, n2973);
  and g1309 (n3168, n_134, n_680);
  and g1310 (n3169, n_645, n3168);
  not g1311 (n_681, n3169);
  and g1312 (n3170, n2746, n_681);
  not g1313 (n_682, n3170);
  and g1314 (n3171, n2744, n_682);
  and g1315 (n3172, n_494, n3171);
  and g1316 (n3173, n_660, n3168);
  not g1317 (n_683, n3173);
  and g1318 (n3174, n2746, n_683);
  not g1319 (n_684, n3174);
  and g1320 (n3175, n3131, n_684);
  not g1321 (n_685, n3175);
  and g1322 (n3176, n_620, n_685);
  not g1323 (n_686, n3172);
  and g1324 (n3177, n_686, n3176);
  not g1325 (n_687, n3177);
  and g1326 (n3178, n_144, n_687);
  not g1327 (n_688, n3178);
  and g1328 (n3179, n_345, n_688);
  not g1329 (n_689, n3179);
  and g1330 (n3180, n_186, n_689);
  and g1331 (n3181, n2442, n2511);
  and g1332 (n3182, n_134, n2510);
  and g1333 (n3183, n2973, n3182);
  not g1334 (n_690, n3183);
  and g1335 (n3184, n3103, n_690);
  not g1336 (n_691, n3184);
  and g1337 (n3185, n3098, n_691);
  not g1338 (n_692, n3181);
  and g1339 (n3186, pi0137, n_692);
  not g1340 (n_693, n3185);
  and g1341 (n3187, n_693, n3186);
  not g1342 (n_694, n3180);
  not g1343 (n_695, n3187);
  and g1344 (n3188, n_694, n_695);
  not g1345 (n_696, n3188);
  and g1346 (n3189, n_271, n_696);
  not g1347 (n_697, n3171);
  and g1348 (n3190, n_672, n_697);
  not g1349 (n_698, n3190);
  and g1350 (n3191, n_144, n_698);
  not g1351 (n_699, n3191);
  and g1352 (n3192, n3084, n_699);
  and g1353 (n3193, n3157, n_691);
  not g1354 (n_700, n3193);
  and g1355 (n3194, n_692, n_700);
  not g1356 (n_701, n3194);
  and g1357 (n3195, pi0137, n_701);
  not g1358 (n_702, n3195);
  and g1359 (n3196, pi0210, n_702);
  not g1360 (n_703, n3192);
  and g1361 (n3197, n_703, n3196);
  not g1362 (n_704, n3197);
  and g1363 (n3198, n2676, n_704);
  not g1364 (n_705, n3189);
  and g1365 (n3199, n_705, n3198);
  not g1366 (n_706, n3167);
  and g1367 (n3200, n2639, n_706);
  not g1368 (n_707, n3199);
  and g1369 (n3201, n_707, n3200);
  and g1370 (n3202, pi0146, n3189);
  and g1371 (n3203, n_268, n_271);
  and g1372 (n3204, n_620, n_697);
  not g1373 (n_708, n3204);
  and g1374 (n3205, n_144, n_708);
  not g1375 (n_709, n3205);
  and g1376 (n3206, n_345, n_709);
  not g1377 (n_710, n3206);
  and g1378 (n3207, n_186, n_710);
  not g1379 (n_711, n3207);
  and g1380 (n3208, n_695, n_711);
  not g1381 (n_712, n3208);
  and g1382 (n3209, n3203, n_712);
  not g1383 (n_713, n3209);
  and g1384 (n3210, n3198, n_713);
  not g1385 (n_714, n3202);
  and g1386 (n3211, n_714, n3210);
  and g1387 (n3212, n_620, n_673);
  not g1388 (n_715, n3212);
  and g1389 (n3213, n_144, n_715);
  not g1390 (n_716, n3213);
  and g1391 (n3214, n2742, n_716);
  not g1392 (n_717, n3214);
  and g1393 (n3215, n_186, n_717);
  not g1394 (n_718, n3215);
  and g1395 (n3216, n_668, n_718);
  not g1396 (n_719, n3216);
  and g1397 (n3217, n3203, n_719);
  and g1398 (n3218, pi0146, n3154);
  not g1399 (n_720, n3217);
  and g1400 (n3219, n3166, n_720);
  not g1401 (n_721, n3218);
  and g1402 (n3220, n_721, n3219);
  not g1403 (n_722, n3211);
  and g1404 (n3221, n_269, n_722);
  not g1405 (n_723, n3220);
  and g1406 (n3222, n_723, n3221);
  not g1407 (n_724, n3201);
  and g1408 (n3223, n_187, n_724);
  not g1409 (n_725, n3222);
  and g1410 (n3224, n_725, n3223);
  not g1411 (n_726, n3094);
  and g1412 (n3225, n_188, n_726);
  not g1413 (n_727, n3224);
  and g1414 (n3226, n_727, n3225);
  not g1415 (n_728, n3036);
  not g1416 (n_729, n3226);
  and g1417 (n3227, n_728, n_729);
  not g1418 (n_730, n3227);
  and g1419 (n3228, n_20, n_730);
  not g1420 (n_731, n3228);
  and g1421 (n3229, n_23, n_731);
  not g1422 (n_732, n3229);
  and g1423 (n3230, n_26, n_732);
  not g1424 (n_733, n3230);
  and g1425 (n3231, n_35, n_733);
  not g1426 (n_734, n3231);
  and g1427 (n3232, n_36, n_734);
  and g1428 (n3233, pi0299, n_38);
  not g1429 (n_735, n3232);
  and g1430 (n3234, n_735, n3233);
  and g1431 (n3235, pi0198, n_528);
  and g1432 (n3236, n_305, n3009);
  not g1433 (n_736, n3235);
  not g1434 (n_737, n3236);
  and g1435 (n3237, n_736, n_737);
  and g1436 (n3238, pi0142, n3237);
  and g1437 (n3239, n_305, n_556);
  not g1438 (n_738, pi0142);
  and g1439 (n3240, n_738, n_736);
  not g1440 (n_739, n3239);
  and g1441 (n3241, n_739, n3240);
  not g1442 (n_740, n3241);
  and g1443 (n3242, n2681, n_740);
  not g1444 (n_741, n3238);
  and g1445 (n3243, n_741, n3242);
  and g1446 (n3244, pi0198, n_482);
  and g1447 (n3245, n_305, n_510);
  not g1448 (n_742, n3244);
  not g1449 (n_743, n3245);
  and g1450 (n3246, n_742, n_743);
  and g1451 (n3247, pi0142, n3246);
  and g1452 (n3248, n_305, n_562);
  and g1453 (n3249, n_738, n_742);
  not g1454 (n_744, n3248);
  and g1455 (n3250, n_744, n3249);
  not g1456 (n_745, n3247);
  and g1457 (n3251, n2676, n_745);
  not g1458 (n_746, n3250);
  and g1459 (n3252, n_746, n3251);
  not g1460 (n_747, n3252);
  and g1461 (n3253, n2670, n_747);
  not g1462 (n_748, n3243);
  and g1463 (n3254, n_748, n3253);
  and g1464 (n3255, n_148, n3246);
  and g1465 (n3256, pi0234, n3237);
  not g1466 (n_749, n3255);
  and g1467 (n3257, n_4, n_749);
  not g1468 (n_750, n3256);
  and g1469 (n3258, n_750, n3257);
  not g1470 (n_751, n3258);
  and g1471 (n3259, n2680, n_751);
  not g1472 (n_752, n3254);
  not g1473 (n_753, n3259);
  and g1474 (n3260, n_752, n_753);
  not g1475 (n_754, n3260);
  and g1476 (n3261, n2603, n_754);
  not g1477 (n_755, n3261);
  and g1478 (n3262, n2602, n_755);
  not g1479 (n_756, n3262);
  and g1480 (n3263, n_162, n_756);
  not g1481 (n_757, n3234);
  and g1482 (n3264, n_757, n3263);
  not g1483 (n_758, n2698);
  and g1484 (n3265, n_161, n_758);
  not g1485 (n_759, n3264);
  and g1486 (n3266, n_759, n3265);
  not g1487 (n_760, n2697);
  and g1488 (n3267, n_164, n_760);
  not g1489 (n_761, n3266);
  and g1490 (n3268, n_761, n3267);
  not g1491 (n_762, n2694);
  and g1492 (n3269, n_172, n_762);
  not g1493 (n_763, n3268);
  and g1494 (n3270, n_763, n3269);
  not g1495 (n_764, n2635);
  and g1496 (n3271, n_171, n_764);
  not g1497 (n_765, n3270);
  and g1498 (n3272, n_765, n3271);
  not g1499 (n_766, n2610);
  and g1500 (n3273, n_250, n_766);
  and g1501 (n3274, n2448, n_289);
  not g1502 (n_767, n3274);
  and g1503 (n3275, n_23, n_767);
  not g1504 (n_768, n3275);
  and g1505 (n3276, n_26, n_768);
  not g1506 (n_769, n3276);
  and g1507 (n3277, n_35, n_769);
  not g1508 (n_770, n3277);
  and g1509 (n3278, n_36, n_770);
  not g1510 (n_771, n3278);
  and g1511 (n3279, n_38, n_771);
  not g1512 (n_772, n3279);
  and g1513 (n3280, pi0299, n_772);
  and g1514 (n3281, n2610, n_321);
  not g1515 (n_773, n3280);
  and g1516 (n3282, n_773, n3281);
  not g1517 (n_774, n3273);
  and g1518 (n3283, pi0075, n_774);
  not g1519 (n_775, n3282);
  and g1520 (n3284, n_775, n3283);
  not g1521 (n_776, n3272);
  not g1522 (n_777, n3284);
  and g1523 (n3285, n_776, n_777);
  not g1524 (n_778, n3285);
  and g1525 (n3286, n_174, n_778);
  not g1526 (n_779, n2634);
  and g1527 (n3287, n_167, n_779);
  not g1528 (n_780, n3286);
  and g1529 (n3288, n_780, n3287);
  not g1530 (n_781, n2624);
  and g1531 (n3289, n_168, n_781);
  not g1532 (n_782, n3288);
  and g1533 (n3290, n_782, n3289);
  and g1534 (n3291, pi0054, n_250);
  and g1535 (n3292, n_167, n2623);
  not g1536 (n_783, n3291);
  and g1537 (n3293, pi0074, n_783);
  not g1538 (n_784, n3292);
  and g1539 (n3294, n_784, n3293);
  not g1540 (n_785, n3290);
  not g1541 (n_786, n3294);
  and g1542 (n3295, n_785, n_786);
  not g1543 (n_787, n3295);
  and g1544 (n3296, n_176, n_787);
  not g1545 (n_788, n2589);
  and g1546 (n3297, n_157, n_788);
  not g1547 (n_789, n3296);
  and g1548 (n3298, n_789, n3297);
  not g1549 (n_790, n2567);
  and g1550 (n3299, n_158, n_790);
  not g1551 (n_791, n3298);
  and g1552 (n3300, n_791, n3299);
  not g1553 (n_792, pi0059);
  not g1554 (n_793, n2566);
  and g1555 (n3301, n_792, n_793);
  not g1556 (n_794, n3300);
  and g1557 (n3302, n_794, n3301);
  not g1558 (n_796, pi0057);
  not g1559 (n_797, n2541);
  and g1560 (n3303, n_796, n_797);
  not g1561 (n_798, n3302);
  and g1562 (n3304, n_798, n3303);
  and g1563 (n3305, n_792, n2539);
  not g1564 (n_799, n3305);
  and g1565 (n3306, n2460, n_799);
  not g1566 (n_800, n3306);
  and g1567 (n3307, pi0057, n_800);
  or g1568 (po0153, n3304, n3307);
  and g1569 (n3309, pi0215, pi1146);
  and g1570 (n3310, pi0216, n_26);
  and g1571 (n3311, pi0276, n3310);
  not g1572 (n_803, pi1146);
  and g1573 (n3312, n_803, n_29);
  not g1574 (n_805, pi0939);
  and g1575 (n3313, n_805, n2452);
  not g1576 (n_806, n3312);
  and g1577 (n3314, pi0221, n_806);
  not g1578 (n_807, n3313);
  and g1579 (n3315, n_807, n3314);
  not g1580 (n_808, n3311);
  not g1581 (n_809, n3315);
  and g1582 (n3316, n_808, n_809);
  not g1583 (n_810, n3316);
  and g1584 (n3317, n_36, n_810);
  not g1585 (n_811, n3309);
  not g1586 (n_812, n3317);
  and g1587 (n3318, n_811, n_812);
  not g1588 (n_814, n3318);
  and g1589 (n3319, pi0154, n_814);
  and g1590 (n3320, n_20, n_19);
  not g1591 (n_815, n3320);
  and g1592 (n3321, n_808, n_815);
  not g1593 (n_816, n3321);
  and g1594 (n3322, n_26, n_816);
  not g1595 (n_817, n3322);
  and g1596 (n3323, n_809, n_817);
  not g1597 (n_818, n3323);
  and g1598 (n3324, n_36, n_818);
  not g1599 (n_819, n3324);
  and g1600 (n3325, n_811, n_819);
  not g1601 (n_820, pi0154);
  not g1602 (n_821, n3325);
  and g1603 (n3326, n_820, n_821);
  not g1604 (n_822, n3319);
  not g1605 (n_823, n3326);
  and g1606 (n3327, n_822, n_823);
  and g1607 (n3328, n_796, n_792);
  not g1608 (n_824, n3328);
  and g1609 (n3329, n3327, n_824);
  and g1610 (n3330, n_157, n2536);
  and g1611 (n3331, n2531, n3330);
  not g1612 (n_825, n3327);
  not g1613 (n_826, n3331);
  and g1614 (n3332, n_825, n_826);
  and g1615 (n3333, n_176, n2572);
  and g1616 (n3334, n_811, n_809);
  and g1617 (n3335, n_188, n2521);
  and g1618 (n3336, n_20, n3335);
  and g1619 (n3337, n3334, n3336);
  and g1620 (n3338, n_822, n3337);
  and g1621 (n3339, n_825, n3333);
  not g1622 (n_827, n3338);
  and g1623 (n3340, n_827, n3339);
  not g1624 (n_828, n3332);
  not g1625 (n_829, n3340);
  and g1626 (n3341, n_828, n_829);
  not g1627 (n_830, n3341);
  and g1628 (n3342, pi0062, n_830);
  and g1629 (n3343, n_179, n_825);
  not g1630 (n_831, n3343);
  and g1631 (n3344, pi0056, n_831);
  and g1632 (n3345, n_829, n3344);
  and g1633 (n3346, n2572, n3338);
  and g1634 (n3347, pi0055, n_825);
  not g1635 (n_832, n3346);
  and g1636 (n3348, n_832, n3347);
  and g1637 (n3349, pi0299, n_825);
  and g1638 (n3350, pi0223, n_803);
  and g1639 (n3351, n_226, pi0224);
  and g1640 (n3352, pi0276, n3351);
  and g1641 (n3353, n_803, n_221);
  and g1642 (n3354, n_805, n2591);
  not g1643 (n_833, n3353);
  and g1644 (n3355, pi0222, n_833);
  not g1645 (n_834, n3354);
  and g1646 (n3356, n_834, n3355);
  not g1647 (n_835, n3352);
  and g1648 (n3357, n_223, n_835);
  not g1649 (n_836, n3356);
  and g1650 (n3358, n_836, n3357);
  not g1651 (n_837, n3350);
  and g1652 (n3359, n_234, n_837);
  not g1653 (n_838, n3358);
  and g1654 (n3360, n_838, n3359);
  not g1655 (n_839, n3349);
  not g1656 (n_840, n3360);
  and g1657 (n3361, n_839, n_840);
  not g1658 (n_841, n2532);
  and g1659 (n3362, n_841, n3361);
  and g1660 (n3363, pi0299, n_814);
  not g1661 (n_842, n3363);
  and g1662 (n3364, n_840, n_842);
  not g1663 (n_843, n3364);
  and g1664 (n3365, pi0154, n_843);
  and g1665 (n3366, pi0299, n_821);
  not g1666 (n_844, n3337);
  and g1667 (n3367, n_844, n3366);
  not g1668 (n_845, n3367);
  and g1669 (n3368, n_840, n_845);
  not g1670 (n_846, n3368);
  and g1671 (n3369, n_820, n_846);
  not g1672 (n_847, n3365);
  and g1673 (n3370, n2625, n_847);
  not g1674 (n_848, n3369);
  and g1675 (n3371, n_848, n3370);
  and g1676 (n3372, n2533, n3371);
  and g1677 (n3373, n2531, n2533);
  not g1678 (n_849, n3373);
  and g1679 (n3374, n3361, n_849);
  not g1680 (n_850, n3374);
  and g1681 (n3375, pi0092, n_850);
  not g1682 (n_851, n3372);
  and g1683 (n3376, n_851, n3375);
  and g1684 (n3377, pi0075, n3361);
  and g1685 (n3378, n_251, n3361);
  not g1686 (n_852, n3371);
  not g1687 (n_853, n3378);
  and g1688 (n3379, n_852, n_853);
  not g1689 (n_854, n3379);
  and g1690 (n3380, pi0087, n_854);
  and g1691 (n3381, n_161, n_20);
  and g1692 (n3382, n_188, n3381);
  and g1693 (n3383, n_820, pi0299);
  and g1694 (n3384, n_268, n_207);
  and g1695 (n3385, n_280, n2521);
  not g1696 (n_855, n3385);
  and g1697 (n3386, pi0146, n_855);
  not g1698 (n_856, n3384);
  not g1699 (n_857, n3386);
  and g1700 (n3387, n_856, n_857);
  not g1701 (n_858, n3387);
  and g1702 (n3388, pi0152, n_858);
  and g1703 (n3389, n_264, n_266);
  and g1704 (n3390, n3385, n3389);
  not g1705 (n_859, n3389);
  and g1706 (n3391, n3387, n_859);
  not g1707 (n_860, n3390);
  and g1708 (n3392, n_263, n_860);
  not g1709 (n_861, n3391);
  and g1710 (n3393, n_861, n3392);
  not g1711 (n_862, n3388);
  not g1712 (n_863, n3393);
  and g1713 (n3394, n_862, n_863);
  not g1718 (n_864, n3361);
  and g1719 (n3399, pi0100, n_864);
  not g1720 (n_865, n3398);
  and g1721 (n3400, n_865, n3399);
  and g1722 (n3401, pi0038, n3361);
  and g1723 (n3402, pi0039, n_207);
  and g1724 (n3403, n_139, n3043);
  and g1725 (n3404, n_339, n_622);
  not g1726 (n_866, n3403);
  and g1727 (n3405, n_866, n3404);
  not g1728 (n_867, n3405);
  and g1729 (n3406, n_138, n_867);
  not g1730 (n_868, n3406);
  and g1731 (n3407, n2748, n_868);
  not g1732 (n_869, n3407);
  and g1733 (n3408, n3168, n_869);
  not g1734 (n_870, n3408);
  and g1735 (n3409, n_348, n_870);
  not g1736 (n_871, n3409);
  and g1737 (n3410, n2510, n_871);
  not g1738 (n_872, n2509);
  and g1739 (n3411, pi0040, n_872);
  not g1740 (n_873, n2710);
  and g1741 (n3412, pi0032, n_873);
  not g1742 (n_874, n3411);
  not g1743 (n_875, n3412);
  and g1744 (n3413, n_874, n_875);
  not g1745 (n_876, n3410);
  and g1746 (n3414, n_876, n3413);
  not g1747 (n_877, n3414);
  and g1748 (n3415, n_144, n_877);
  not g1749 (n_878, n3415);
  and g1750 (n3416, n_345, n_878);
  not g1751 (n_879, n3416);
  and g1752 (n3417, n_162, n_879);
  not g1753 (n_880, n3402);
  not g1754 (n_881, n3417);
  and g1755 (n3418, n_880, n_881);
  not g1759 (n_882, n3421);
  and g1760 (n3422, n3366, n_882);
  not g1761 (n_883, n3422);
  and g1762 (n3423, n_840, n_883);
  not g1763 (n_884, n3423);
  and g1764 (n3424, n_820, n_884);
  and g1765 (n3425, n_161, n_847);
  not g1766 (n_885, n3424);
  and g1767 (n3426, n_885, n3425);
  not g1768 (n_886, n3401);
  and g1769 (n3427, n_164, n_886);
  not g1770 (n_887, n3426);
  and g1771 (n3428, n_887, n3427);
  not g1772 (n_888, n3400);
  and g1773 (n3429, n_172, n_888);
  not g1774 (n_889, n3428);
  and g1775 (n3430, n_889, n3429);
  not g1776 (n_890, n3380);
  not g1777 (n_891, n3430);
  and g1778 (n3431, n_890, n_891);
  not g1779 (n_892, n3431);
  and g1780 (n3432, n_171, n_892);
  not g1781 (n_893, n3377);
  and g1782 (n3433, n_174, n_893);
  not g1783 (n_894, n3432);
  and g1784 (n3434, n_894, n3433);
  not g1785 (n_895, n3376);
  and g1786 (n3435, n2532, n_895);
  not g1787 (n_896, n3434);
  and g1788 (n3436, n_896, n3435);
  not g1789 (n_897, n3362);
  and g1790 (n3437, n_176, n_897);
  not g1791 (n_898, n3436);
  and g1792 (n3438, n_898, n3437);
  not g1793 (n_899, n3348);
  and g1794 (n3439, n_157, n_899);
  not g1795 (n_900, n3438);
  and g1796 (n3440, n_900, n3439);
  not g1797 (n_901, n3345);
  and g1798 (n3441, n_158, n_901);
  not g1799 (n_902, n3440);
  and g1800 (n3442, n_902, n3441);
  not g1801 (n_903, n3342);
  and g1802 (n3443, n3328, n_903);
  not g1803 (n_904, n3442);
  and g1804 (n3444, n_904, n3443);
  not g1805 (n_906, pi0239);
  not g1806 (n_907, n3329);
  and g1807 (n3445, n_906, n_907);
  not g1808 (n_908, n3444);
  and g1809 (n3446, n_908, n3445);
  and g1810 (n3447, n2441, n2442);
  and g1811 (n3448, n_20, n_26);
  and g1812 (n3449, n_36, n3448);
  and g1813 (n3450, n3447, n3449);
  not g1814 (n_909, n3450);
  and g1815 (n3451, n3318, n_909);
  not g1816 (n_910, n3451);
  and g1817 (n3452, n_36, n_910);
  and g1818 (n3453, pi0154, n_910);
  not g1819 (n_911, n3452);
  and g1820 (n3454, n_823, n_911);
  not g1821 (n_912, n3453);
  and g1822 (n3455, n_912, n3454);
  and g1823 (n3456, n_824, n3455);
  not g1824 (n_913, n3455);
  and g1825 (n3457, n_826, n_913);
  and g1826 (n3458, n3337, n_912);
  not g1827 (n_914, n3458);
  and g1828 (n3459, n_913, n_914);
  and g1829 (n3460, n3333, n3459);
  and g1830 (n3461, n_157, n3460);
  not g1831 (n_915, n3457);
  not g1832 (n_916, n3461);
  and g1833 (n3462, n_915, n_916);
  not g1834 (n_917, n3462);
  and g1835 (n3463, pi0062, n_917);
  and g1836 (n3464, n_179, n_913);
  not g1837 (n_918, n3464);
  and g1838 (n3465, pi0056, n_918);
  not g1839 (n_919, n3460);
  and g1840 (n3466, n_919, n3465);
  and g1841 (n3467, n2572, n3458);
  and g1842 (n3468, pi0055, n_913);
  not g1843 (n_920, n3467);
  and g1844 (n3469, n_920, n3468);
  and g1845 (n3470, n_223, n_234);
  and g1846 (n3471, n2603, n3470);
  and g1847 (n3472, n2442, n3471);
  and g1848 (n3473, pi0299, n_913);
  not g1849 (n_921, n3472);
  and g1850 (n3474, n_840, n_921);
  not g1851 (n_922, n3473);
  and g1852 (n3475, n_922, n3474);
  and g1853 (n3476, n_841, n3475);
  not g1854 (n_923, n3459);
  and g1855 (n3477, pi0299, n_923);
  and g1856 (n3478, n3373, n3477);
  not g1857 (n_924, n3475);
  and g1858 (n3479, pi0092, n_924);
  not g1859 (n_925, n3478);
  and g1860 (n3480, n_925, n3479);
  and g1861 (n3481, pi0075, n3475);
  and g1862 (n3482, n2625, n3477);
  and g1863 (n3483, pi0087, n_924);
  not g1864 (n_926, n3482);
  and g1865 (n3484, n_926, n3483);
  not g1866 (n_927, n3477);
  and g1867 (n3485, n_924, n_927);
  not g1868 (n_928, n3485);
  and g1869 (n3486, pi0039, n_928);
  and g1870 (n3487, n2519, n2973);
  not g1871 (n_929, n3487);
  and g1872 (n3488, n_145, n_929);
  and g1873 (n3489, n_219, n3488);
  not g1874 (n_930, pi0276);
  and g1875 (n3490, pi0224, n_930);
  not g1876 (n_931, n3490);
  and g1877 (n3491, n_226, n_931);
  not g1878 (n_932, n3489);
  and g1879 (n3492, n_932, n3491);
  and g1880 (n3493, n_223, n_836);
  not g1881 (n_933, n3492);
  and g1882 (n3494, n_933, n3493);
  not g1883 (n_934, n3494);
  and g1884 (n3495, n_837, n_934);
  not g1885 (n_935, n3495);
  and g1886 (n3496, n_234, n_935);
  not g1887 (n_936, n3488);
  and g1888 (n3497, pi0105, n_936);
  not g1889 (n_937, n3497);
  and g1890 (n3498, pi0228, n_937);
  and g1891 (n3499, n_345, n_936);
  not g1892 (n_938, n3499);
  and g1893 (n3500, n_188, n_938);
  not g1894 (n_939, n3498);
  not g1895 (n_940, n3500);
  and g1896 (n3501, n_939, n_940);
  not g1897 (n_941, n3501);
  and g1898 (n3502, pi0154, n_941);
  and g1899 (n3503, n_134, n_869);
  not g1900 (n_942, n3503);
  and g1901 (n3504, n_348, n_942);
  not g1902 (n_943, n3504);
  and g1903 (n3505, n2510, n_943);
  not g1904 (n_944, n3505);
  and g1905 (n3506, n3413, n_944);
  not g1906 (n_945, n3506);
  and g1907 (n3507, n_144, n_945);
  not g1908 (n_946, n3507);
  and g1909 (n3508, n2742, n_946);
  and g1910 (n3509, n_188, n3508);
  and g1911 (n3510, n2441, n3488);
  not g1912 (n_947, n3509);
  not g1913 (n_948, n3510);
  and g1914 (n3511, n_947, n_948);
  not g1915 (n_949, n3511);
  and g1916 (n3512, n_820, n_949);
  not g1917 (n_950, n3502);
  and g1918 (n3513, n3449, n_950);
  not g1919 (n_951, n3512);
  and g1920 (n3514, n_951, n3513);
  and g1921 (n3515, pi0299, n3318);
  not g1922 (n_952, n3514);
  and g1923 (n3516, n_952, n3515);
  not g1924 (n_953, n3496);
  not g1925 (n_954, n3516);
  and g1926 (n3517, n_953, n_954);
  not g1927 (n_955, n3517);
  and g1928 (n3518, n_162, n_955);
  not g1929 (n_956, n3486);
  and g1930 (n3519, n2608, n_956);
  not g1931 (n_957, n3518);
  and g1932 (n3520, n_957, n3519);
  and g1933 (n3521, pi0100, n3398);
  not g1934 (n_958, n2608);
  and g1935 (n3522, n_958, n_924);
  not g1936 (n_959, n3521);
  and g1937 (n3523, n_959, n3522);
  not g1938 (n_960, n3520);
  not g1939 (n_961, n3523);
  and g1940 (n3524, n_960, n_961);
  not g1941 (n_962, n3524);
  and g1942 (n3525, n_172, n_962);
  not g1943 (n_963, n3484);
  and g1944 (n3526, n_171, n_963);
  not g1945 (n_964, n3525);
  and g1946 (n3527, n_964, n3526);
  not g1947 (n_965, n3481);
  and g1948 (n3528, n_174, n_965);
  not g1949 (n_966, n3527);
  and g1950 (n3529, n_966, n3528);
  not g1951 (n_967, n3480);
  and g1952 (n3530, n2532, n_967);
  not g1953 (n_968, n3529);
  and g1954 (n3531, n_968, n3530);
  not g1955 (n_969, n3476);
  and g1956 (n3532, n_176, n_969);
  not g1957 (n_970, n3531);
  and g1958 (n3533, n_970, n3532);
  not g1959 (n_971, n3469);
  and g1960 (n3534, n_157, n_971);
  not g1961 (n_972, n3533);
  and g1962 (n3535, n_972, n3534);
  not g1963 (n_973, n3466);
  and g1964 (n3536, n_158, n_973);
  not g1965 (n_974, n3535);
  and g1966 (n3537, n_974, n3536);
  not g1967 (n_975, n3463);
  and g1968 (n3538, n3328, n_975);
  not g1969 (n_976, n3537);
  and g1970 (n3539, n_976, n3538);
  not g1971 (n_977, n3456);
  and g1972 (n3540, pi0239, n_977);
  not g1973 (n_978, n3539);
  and g1974 (n3541, n_978, n3540);
  or g1975 (po0154, n3446, n3541);
  and g1976 (n3543, pi0215, pi1145);
  and g1977 (n3544, pi0216, pi0274);
  not g1978 (n_981, n3544);
  and g1979 (n3545, n_26, n_981);
  not g1980 (n_983, pi0151);
  and g1981 (n3546, n_983, n_19);
  not g1982 (n_984, n3546);
  and g1983 (n3547, n_20, n_984);
  not g1984 (n_985, n3547);
  and g1985 (n3548, n3545, n_985);
  not g1986 (n_986, pi1145);
  and g1987 (n3549, n_986, n_29);
  not g1988 (n_988, pi0927);
  and g1989 (n3550, n_988, n2452);
  not g1990 (n_989, n3549);
  and g1991 (n3551, pi0221, n_989);
  not g1992 (n_990, n3550);
  and g1993 (n3552, n_990, n3551);
  not g1994 (n_991, n3548);
  not g1995 (n_992, n3552);
  and g1996 (n3553, n_991, n_992);
  not g1997 (n_993, n3553);
  and g1998 (n3554, n_36, n_993);
  not g1999 (n_994, n3543);
  not g2000 (n_995, n3554);
  and g2001 (n3555, n_994, n_995);
  and g2002 (n3556, n2526, n3447);
  and g2003 (n3557, n_981, n3556);
  not g2004 (n_996, n3557);
  and g2005 (n3558, n3555, n_996);
  and g2006 (n3559, n_826, n3558);
  not g2007 (n_997, n3447);
  and g2008 (n3560, n_997, n_984);
  and g2009 (n3561, n_983, n3335);
  not g2010 (n_998, n3560);
  not g2011 (n_999, n3561);
  and g2012 (n3562, n_998, n_999);
  not g2013 (n_1000, n3562);
  and g2014 (n3563, n_20, n_1000);
  not g2015 (n_1001, n3563);
  and g2016 (n3564, n3545, n_1001);
  not g2017 (n_1002, n3564);
  and g2018 (n3565, n_992, n_1002);
  not g2019 (n_1003, n3565);
  and g2020 (n3566, n_36, n_1003);
  not g2021 (n_1004, n3566);
  and g2022 (n3567, n_994, n_1004);
  and g2023 (n3568, n3331, n3567);
  not g2024 (n_1005, n3559);
  and g2025 (n3569, pi0062, n_1005);
  not g2026 (n_1006, n3568);
  and g2027 (n3570, n_1006, n3569);
  not g2028 (n_1007, n3558);
  and g2029 (n3571, n_179, n_1007);
  not g2030 (n_1008, n3567);
  and g2031 (n3572, n2537, n_1008);
  not g2032 (n_1009, n3571);
  and g2033 (n3573, pi0056, n_1009);
  not g2034 (n_1010, n3572);
  and g2035 (n3574, n_1010, n3573);
  and g2036 (n3575, n_204, n3558);
  and g2037 (n3576, n2572, n3567);
  not g2038 (n_1011, n3575);
  and g2039 (n3577, pi0055, n_1011);
  not g2040 (n_1012, n3576);
  and g2041 (n3578, n_1012, n3577);
  and g2042 (n3579, pi0223, pi1145);
  and g2043 (n3580, n_986, n_221);
  and g2044 (n3581, n_988, n2591);
  not g2045 (n_1013, n3580);
  and g2046 (n3582, pi0222, n_1013);
  not g2047 (n_1014, n3581);
  and g2048 (n3583, n_1014, n3582);
  and g2049 (n3584, pi0224, pi0274);
  not g2050 (n_1015, n3584);
  and g2051 (n3585, n3351, n_1015);
  not g2052 (n_1016, n3583);
  not g2053 (n_1017, n3585);
  and g2054 (n3586, n_1016, n_1017);
  not g2055 (n_1018, n3586);
  and g2056 (n3587, n_223, n_1018);
  not g2057 (n_1019, n3579);
  not g2058 (n_1020, n3587);
  and g2059 (n3588, n_1019, n_1020);
  not g2060 (n_1021, n3588);
  and g2061 (n3589, n_234, n_1021);
  not g2062 (n_1022, n3589);
  and g2063 (n3590, n_921, n_1022);
  and g2064 (n3591, pi0299, n_1007);
  not g2065 (n_1023, n3591);
  and g2066 (n3592, n3590, n_1023);
  and g2067 (n3593, n_841, n3592);
  and g2068 (n3594, n_251, n3592);
  and g2069 (n3595, pi0299, n_1008);
  not g2070 (n_1024, n3595);
  and g2071 (n3596, n3590, n_1024);
  and g2072 (n3597, n2625, n3596);
  not g2073 (n_1025, n3594);
  not g2074 (n_1026, n3597);
  and g2075 (n3598, n_1025, n_1026);
  not g2076 (n_1027, n3598);
  and g2077 (n3599, n2533, n_1027);
  and g2078 (n3600, n_257, n3592);
  not g2079 (n_1028, n3600);
  and g2080 (n3601, pi0092, n_1028);
  not g2081 (n_1029, n3599);
  and g2082 (n3602, n_1029, n3601);
  and g2083 (n3603, pi0075, n3592);
  and g2084 (n3604, pi0087, n3598);
  and g2085 (n3605, pi0038, n3592);
  not g2086 (n_1030, n3596);
  and g2087 (n3606, pi0039, n_1030);
  and g2088 (n3607, n_226, n_1015);
  and g2089 (n3608, n_932, n3607);
  not g2090 (n_1031, n3608);
  and g2091 (n3609, n_1016, n_1031);
  not g2092 (n_1032, n3609);
  and g2093 (n3610, n_223, n_1032);
  and g2094 (n3611, n_234, n_1019);
  not g2095 (n_1033, n3610);
  and g2096 (n3612, n_1033, n3611);
  and g2097 (n3613, n_983, n3511);
  and g2098 (n3614, pi0151, n3501);
  not g2099 (n_1034, n3614);
  and g2100 (n3615, n_20, n_1034);
  not g2101 (n_1035, n3613);
  and g2102 (n3616, n_1035, n3615);
  not g2103 (n_1036, n3616);
  and g2104 (n3617, n3545, n_1036);
  not g2105 (n_1037, n3617);
  and g2106 (n3618, n_992, n_1037);
  not g2107 (n_1038, n3618);
  and g2108 (n3619, n_36, n_1038);
  and g2109 (n3620, pi0299, n_994);
  not g2110 (n_1039, n3619);
  and g2111 (n3621, n_1039, n3620);
  not g2112 (n_1040, n3612);
  and g2113 (n3622, n_162, n_1040);
  not g2114 (n_1041, n3621);
  and g2115 (n3623, n_1041, n3622);
  not g2116 (n_1042, n3606);
  and g2117 (n3624, n_161, n_1042);
  not g2118 (n_1043, n3623);
  and g2119 (n3625, n_1043, n3624);
  not g2120 (n_1044, n3605);
  and g2121 (n3626, n_164, n_1044);
  not g2122 (n_1045, n3625);
  and g2123 (n3627, n_1045, n3626);
  and g2124 (n3628, n_260, n3592);
  and g2125 (n3629, n_188, n3394);
  and g2126 (n3630, n2441, n_145);
  not g2127 (n_1046, n3629);
  not g2128 (n_1047, n3630);
  and g2129 (n3631, n_1046, n_1047);
  and g2130 (n3632, n_983, n3631);
  not g2131 (n_1048, n3632);
  and g2132 (n3633, n3563, n_1048);
  not g2133 (n_1049, n3633);
  and g2134 (n3634, n3545, n_1049);
  not g2135 (n_1050, n3634);
  and g2136 (n3635, n_992, n_1050);
  not g2137 (n_1051, n3635);
  and g2138 (n3636, n_36, n_1051);
  not g2139 (n_1052, n3636);
  and g2140 (n3637, n_994, n_1052);
  not g2141 (n_1053, n3637);
  and g2142 (n3638, pi0299, n_1053);
  and g2143 (n3639, n2530, n3590);
  not g2144 (n_1054, n3638);
  and g2145 (n3640, n_1054, n3639);
  not g2146 (n_1055, n3628);
  and g2147 (n3641, pi0100, n_1055);
  not g2148 (n_1056, n3640);
  and g2149 (n3642, n_1056, n3641);
  not g2150 (n_1057, n3627);
  not g2151 (n_1058, n3642);
  and g2152 (n3643, n_1057, n_1058);
  not g2153 (n_1059, n3643);
  and g2154 (n3644, n_172, n_1059);
  not g2155 (n_1060, n3604);
  and g2156 (n3645, n_171, n_1060);
  not g2157 (n_1061, n3644);
  and g2158 (n3646, n_1061, n3645);
  not g2159 (n_1062, n3603);
  and g2160 (n3647, n_174, n_1062);
  not g2161 (n_1063, n3646);
  and g2162 (n3648, n_1063, n3647);
  not g2163 (n_1064, n3602);
  and g2164 (n3649, n2532, n_1064);
  not g2165 (n_1065, n3648);
  and g2166 (n3650, n_1065, n3649);
  not g2167 (n_1066, n3593);
  and g2168 (n3651, n_176, n_1066);
  not g2169 (n_1067, n3650);
  and g2170 (n3652, n_1067, n3651);
  not g2171 (n_1068, n3578);
  and g2172 (n3653, n_157, n_1068);
  not g2173 (n_1069, n3652);
  and g2174 (n3654, n_1069, n3653);
  not g2175 (n_1070, n3574);
  and g2176 (n3655, n_158, n_1070);
  not g2177 (n_1071, n3654);
  and g2178 (n3656, n_1071, n3655);
  and g2184 (n3660, n_994, n_992);
  and g2185 (n3661, n3336, n3660);
  and g2186 (n3662, n2537, n3661);
  and g2187 (n3663, n_157, n3662);
  not g2188 (n_1075, n3555);
  and g2189 (n3664, pi0062, n_1075);
  not g2190 (n_1076, n3663);
  and g2191 (n3665, n_1076, n3664);
  not g2192 (n_1077, n3662);
  and g2193 (n3666, n_1075, n_1077);
  not g2194 (n_1078, n3666);
  and g2195 (n3667, pi0056, n_1078);
  and g2196 (n3668, n2572, n3661);
  and g2197 (n3669, pi0055, n_1075);
  not g2198 (n_1079, n3668);
  and g2199 (n3670, n_1079, n3669);
  and g2200 (n3671, pi0299, n_1075);
  not g2201 (n_1080, n3671);
  and g2202 (n3672, n_1022, n_1080);
  and g2203 (n3673, n_841, n3672);
  not g2204 (n_1081, n3661);
  and g2205 (n3674, n_1081, n3671);
  and g2206 (n3675, n2531, n_1022);
  not g2207 (n_1082, n3674);
  and g2208 (n3676, n_1082, n3675);
  and g2209 (n3677, n2533, n3676);
  and g2210 (n3678, n_849, n3672);
  not g2211 (n_1083, n3678);
  and g2212 (n3679, pi0092, n_1083);
  not g2213 (n_1084, n3677);
  and g2214 (n3680, n_1084, n3679);
  and g2215 (n3681, pi0075, n3672);
  and g2216 (n3682, n_251, n3672);
  not g2217 (n_1085, n3676);
  not g2218 (n_1086, n3682);
  and g2219 (n3683, n_1085, n_1086);
  not g2220 (n_1087, n3683);
  and g2221 (n3684, pi0087, n_1087);
  and g2222 (n3685, n_164, n3418);
  and g2223 (n3686, n_162, pi0100);
  and g2224 (n3687, n3394, n3686);
  not g2225 (n_1088, n3685);
  not g2226 (n_1089, n3687);
  and g2227 (n3688, n_1088, n_1089);
  and g2228 (n3689, n3382, n3660);
  not g2229 (n_1090, n3688);
  and g2230 (n3690, n_1090, n3689);
  not g2231 (n_1091, n3690);
  and g2232 (n3691, n3671, n_1091);
  and g2233 (n3692, n_172, n_1022);
  not g2234 (n_1092, n3691);
  and g2235 (n3693, n_1092, n3692);
  not g2236 (n_1093, n3684);
  not g2237 (n_1094, n3693);
  and g2238 (n3694, n_1093, n_1094);
  not g2239 (n_1095, n3694);
  and g2240 (n3695, n_171, n_1095);
  not g2241 (n_1096, n3681);
  and g2242 (n3696, n_174, n_1096);
  not g2243 (n_1097, n3695);
  and g2244 (n3697, n_1097, n3696);
  not g2245 (n_1098, n3680);
  and g2246 (n3698, n2532, n_1098);
  not g2247 (n_1099, n3697);
  and g2248 (n3699, n_1099, n3698);
  not g2249 (n_1100, n3673);
  and g2250 (n3700, n_176, n_1100);
  not g2251 (n_1101, n3699);
  and g2252 (n3701, n_1101, n3700);
  not g2253 (n_1102, n3670);
  and g2254 (n3702, n_157, n_1102);
  not g2255 (n_1103, n3701);
  and g2256 (n3703, n_1103, n3702);
  not g2257 (n_1104, n3667);
  and g2258 (n3704, n_158, n_1104);
  not g2259 (n_1105, n3703);
  and g2260 (n3705, n_1105, n3704);
  not g2261 (n_1106, pi0235);
  and g2267 (n3709, pi0235, n3557);
  not g2268 (n_1109, n3709);
  and g2269 (n3710, n_824, n_1109);
  and g2270 (n3711, n3555, n3710);
  not g2271 (n_1110, n3708);
  not g2272 (n_1111, n3711);
  and g2273 (n3712, n_1110, n_1111);
  not g2274 (n_1112, n3659);
  and g2275 (po0155, n_1112, n3712);
  and g2276 (n3714, pi0215, pi1143);
  and g2277 (n3715, pi0216, pi0264);
  not g2278 (n_1115, n3715);
  and g2279 (n3716, n_26, n_1115);
  and g2280 (n3717, n_180, pi0146);
  and g2281 (n3718, pi0284, n_145);
  not g2282 (n_1117, n3718);
  and g2283 (n3719, pi0105, n_1117);
  not g2284 (n_1118, n3717);
  and g2285 (n3720, pi0228, n_1118);
  not g2286 (n_1119, n3719);
  and g2287 (n3721, n_1119, n3720);
  not g2288 (n_1120, n3721);
  and g2289 (n3722, n_997, n_1120);
  and g2290 (n3723, n_268, n_188);
  not g2291 (n_1121, n3723);
  and g2292 (n3724, n3722, n_1121);
  not g2293 (n_1122, n3724);
  and g2294 (n3725, n_20, n_1122);
  not g2295 (n_1123, n3725);
  and g2296 (n3726, n3716, n_1123);
  not g2297 (n_1124, pi1143);
  and g2298 (n3727, n_1124, n_29);
  not g2299 (n_1126, pi0944);
  and g2300 (n3728, n_1126, n2452);
  not g2301 (n_1127, n3727);
  and g2302 (n3729, pi0221, n_1127);
  not g2303 (n_1128, n3728);
  and g2304 (n3730, n_1128, n3729);
  not g2305 (n_1129, n3726);
  not g2306 (n_1130, n3730);
  and g2307 (n3731, n_1129, n_1130);
  not g2308 (n_1131, n3731);
  and g2309 (n3732, n_36, n_1131);
  not g2310 (n_1132, n3714);
  not g2311 (n_1133, n3732);
  and g2312 (n3733, n_1132, n_1133);
  and g2313 (n3734, n_826, n3733);
  and g2314 (n3735, pi0284, n2521);
  not g2315 (n_1134, n3735);
  and g2316 (n3736, n_856, n_1134);
  not g2317 (n_1135, n3736);
  and g2318 (n3737, n_188, n_1135);
  not g2319 (n_1136, n3737);
  and g2320 (n3738, n3722, n_1136);
  not g2321 (n_1137, n3738);
  and g2322 (n3739, n_20, n_1137);
  not g2323 (n_1138, n3739);
  and g2324 (n3740, n3716, n_1138);
  not g2325 (n_1139, n3740);
  and g2326 (n3741, n_1130, n_1139);
  not g2327 (n_1140, n3741);
  and g2328 (n3742, n_36, n_1140);
  not g2329 (n_1141, n3742);
  and g2330 (n3743, n_1132, n_1141);
  and g2331 (n3744, n3331, n3743);
  not g2332 (n_1142, n3734);
  and g2333 (n3745, pi0062, n_1142);
  not g2334 (n_1143, n3744);
  and g2335 (n3746, n_1143, n3745);
  not g2336 (n_1144, n3733);
  and g2337 (n3747, n_179, n_1144);
  not g2338 (n_1145, n3743);
  and g2339 (n3748, n2537, n_1145);
  not g2340 (n_1146, n3747);
  and g2341 (n3749, pi0056, n_1146);
  not g2342 (n_1147, n3748);
  and g2343 (n3750, n_1147, n3749);
  and g2344 (n3751, n_204, n3733);
  and g2345 (n3752, n2572, n3743);
  not g2346 (n_1148, n3751);
  and g2347 (n3753, pi0055, n_1148);
  not g2348 (n_1149, n3752);
  and g2349 (n3754, n_1149, n3753);
  and g2350 (n3755, n2442, n2604);
  and g2351 (n3756, pi0223, pi1143);
  and g2352 (n3757, pi0224, pi0264);
  not g2353 (n_1150, n3757);
  and g2354 (n3758, n_226, n_1150);
  and g2355 (n3759, n_219, n3718);
  not g2356 (n_1151, n3759);
  and g2357 (n3760, n3758, n_1151);
  and g2358 (n3761, n_1124, n_221);
  and g2359 (n3762, n_1126, n2591);
  not g2360 (n_1152, n3761);
  and g2361 (n3763, pi0222, n_1152);
  not g2362 (n_1153, n3762);
  and g2363 (n3764, n_1153, n3763);
  not g2364 (n_1154, n3760);
  not g2365 (n_1155, n3764);
  and g2366 (n3765, n_1154, n_1155);
  not g2367 (n_1156, n3765);
  and g2368 (n3766, n_223, n_1156);
  not g2369 (n_1157, n3756);
  not g2370 (n_1158, n3766);
  and g2371 (n3767, n_1157, n_1158);
  not g2372 (n_1159, n3767);
  and g2373 (n3768, n_234, n_1159);
  not g2374 (n_1160, n3755);
  and g2375 (n3769, n_1160, n3768);
  and g2376 (n3770, pi0299, n_1144);
  not g2377 (n_1161, n3769);
  not g2378 (n_1162, n3770);
  and g2379 (n3771, n_1161, n_1162);
  and g2380 (n3772, n_841, n3771);
  and g2381 (n3773, n_251, n3771);
  and g2382 (n3774, pi0299, n_1145);
  not g2383 (n_1163, n3774);
  and g2384 (n3775, n_1161, n_1163);
  and g2385 (n3776, n2625, n3775);
  not g2386 (n_1164, n3773);
  not g2387 (n_1165, n3776);
  and g2388 (n3777, n_1164, n_1165);
  not g2389 (n_1166, n3777);
  and g2390 (n3778, n2533, n_1166);
  and g2391 (n3779, n_257, n3771);
  not g2392 (n_1167, n3779);
  and g2393 (n3780, pi0092, n_1167);
  not g2394 (n_1168, n3778);
  and g2395 (n3781, n_1168, n3780);
  and g2396 (n3782, pi0075, n3771);
  and g2397 (n3783, pi0087, n3777);
  and g2398 (n3784, pi0038, n3771);
  not g2399 (n_1169, n3775);
  and g2400 (n3785, pi0039, n_1169);
  and g2401 (n3786, n_234, n_1157);
  not g2402 (n_1170, pi0284);
  and g2403 (n3787, n_1170, n3488);
  not g2404 (n_1171, n3787);
  and g2405 (n3788, n_219, n_1171);
  not g2406 (n_1172, n3788);
  and g2407 (n3789, n3758, n_1172);
  not g2408 (n_1173, n3789);
  and g2409 (n3790, n_1155, n_1173);
  and g2410 (n3791, n3786, n3790);
  and g2411 (n3792, pi0299, n_1132);
  and g2412 (n3793, n2441, n_936);
  not g2413 (n_1174, n3508);
  and g2414 (n3794, n_268, n_1174);
  and g2415 (n3795, pi0146, n3499);
  not g2416 (n_1175, n3795);
  and g2417 (n3796, n_1170, n_1175);
  and g2418 (n3797, pi0146, pi0284);
  and g2419 (n3798, n_879, n3797);
  not g2420 (n_1176, n3796);
  not g2421 (n_1177, n3798);
  and g2422 (n3799, n_1176, n_1177);
  not g2423 (n_1178, n3794);
  not g2424 (n_1179, n3799);
  and g2425 (n3800, n_1178, n_1179);
  not g2426 (n_1180, n3800);
  and g2427 (n3801, n_188, n_1180);
  not g2428 (n_1181, n3793);
  and g2429 (n3802, n_1120, n_1181);
  not g2430 (n_1182, n3801);
  and g2431 (n3803, n_1182, n3802);
  not g2432 (n_1183, n3803);
  and g2433 (n3804, n_20, n_1183);
  not g2434 (n_1184, n3804);
  and g2435 (n3805, n3716, n_1184);
  not g2436 (n_1185, n3805);
  and g2437 (n3806, n_1130, n_1185);
  not g2438 (n_1186, n3806);
  and g2439 (n3807, n_36, n_1186);
  not g2440 (n_1187, n3807);
  and g2441 (n3808, n3792, n_1187);
  and g2442 (n3809, n_936, n3758);
  not g2443 (n_1188, n3809);
  and g2444 (n3810, n3790, n_1188);
  not g2445 (n_1189, n3810);
  and g2446 (n3811, n_223, n_1189);
  not g2447 (n_1190, n3811);
  and g2448 (n3812, n3786, n_1190);
  not g2449 (n_1191, n3812);
  and g2450 (n3813, n_162, n_1191);
  not g2451 (n_1192, n3791);
  and g2452 (n3814, n_1192, n3813);
  not g2453 (n_1193, n3808);
  and g2454 (n3815, n_1193, n3814);
  not g2455 (n_1194, n3785);
  and g2456 (n3816, n_161, n_1194);
  not g2457 (n_1195, n3815);
  and g2458 (n3817, n_1195, n3816);
  not g2459 (n_1196, n3784);
  and g2460 (n3818, n_164, n_1196);
  not g2461 (n_1197, n3817);
  and g2462 (n3819, n_1197, n3818);
  and g2463 (n3820, n_260, n3771);
  and g2464 (n3821, pi0252, n2639);
  not g2465 (n_1198, n3821);
  and g2466 (n3822, n_1170, n_1198);
  and g2467 (n3823, n2521, n3822);
  not g2468 (n_1199, n3823);
  and g2469 (n3824, n_188, n_1199);
  and g2470 (n3825, n_857, n3824);
  not g2471 (n_1200, n3825);
  and g2472 (n3826, n3722, n_1200);
  not g2473 (n_1201, n3826);
  and g2474 (n3827, n_20, n_1201);
  not g2475 (n_1202, n3827);
  and g2476 (n3828, n3716, n_1202);
  not g2477 (n_1203, n3828);
  and g2478 (n3829, n_1130, n_1203);
  not g2479 (n_1204, n3829);
  and g2480 (n3830, n_36, n_1204);
  not g2481 (n_1205, n3830);
  and g2482 (n3831, n_1132, n_1205);
  not g2483 (n_1206, n3831);
  and g2484 (n3832, pi0299, n_1206);
  and g2485 (n3833, n2530, n_1161);
  not g2486 (n_1207, n3832);
  and g2487 (n3834, n_1207, n3833);
  not g2488 (n_1208, n3820);
  and g2489 (n3835, pi0100, n_1208);
  not g2490 (n_1209, n3834);
  and g2491 (n3836, n_1209, n3835);
  not g2492 (n_1210, n3819);
  not g2493 (n_1211, n3836);
  and g2494 (n3837, n_1210, n_1211);
  not g2495 (n_1212, n3837);
  and g2496 (n3838, n_172, n_1212);
  not g2497 (n_1213, n3783);
  and g2498 (n3839, n_171, n_1213);
  not g2499 (n_1214, n3838);
  and g2500 (n3840, n_1214, n3839);
  not g2501 (n_1215, n3782);
  and g2502 (n3841, n_174, n_1215);
  not g2503 (n_1216, n3840);
  and g2504 (n3842, n_1216, n3841);
  not g2505 (n_1217, n3781);
  and g2506 (n3843, n2532, n_1217);
  not g2507 (n_1218, n3842);
  and g2508 (n3844, n_1218, n3843);
  not g2509 (n_1219, n3772);
  and g2510 (n3845, n_176, n_1219);
  not g2511 (n_1220, n3844);
  and g2512 (n3846, n_1220, n3845);
  not g2513 (n_1221, n3754);
  and g2514 (n3847, n_157, n_1221);
  not g2515 (n_1222, n3846);
  and g2516 (n3848, n_1222, n3847);
  not g2517 (n_1223, n3750);
  and g2518 (n3849, n_158, n_1223);
  not g2519 (n_1224, n3848);
  and g2520 (n3850, n_1224, n3849);
  not g2521 (n_1226, pi0238);
  and g2527 (n3854, n_1120, n_1136);
  not g2528 (n_1229, n3854);
  and g2529 (n3855, n_20, n_1229);
  not g2530 (n_1230, n3855);
  and g2531 (n3856, n3716, n_1230);
  not g2532 (n_1231, n3856);
  and g2533 (n3857, n_1130, n_1231);
  not g2534 (n_1232, n3857);
  and g2535 (n3858, n_36, n_1232);
  not g2536 (n_1233, n3858);
  and g2537 (n3859, n_1132, n_1233);
  and g2538 (n3860, n3331, n3859);
  and g2539 (n3861, n3556, n_1115);
  not g2540 (n_1234, n3861);
  and g2541 (n3862, n3733, n_1234);
  and g2542 (n3863, n_826, n3862);
  not g2543 (n_1235, n3863);
  and g2544 (n3864, pi0062, n_1235);
  not g2545 (n_1236, n3860);
  and g2546 (n3865, n_1236, n3864);
  not g2547 (n_1237, n3862);
  and g2548 (n3866, n_179, n_1237);
  not g2549 (n_1238, n3859);
  and g2550 (n3867, n2537, n_1238);
  not g2551 (n_1239, n3866);
  and g2552 (n3868, pi0056, n_1239);
  not g2553 (n_1240, n3867);
  and g2554 (n3869, n_1240, n3868);
  and g2555 (n3870, n2572, n3859);
  and g2556 (n3871, n_204, n3862);
  not g2557 (n_1241, n3871);
  and g2558 (n3872, pi0055, n_1241);
  not g2559 (n_1242, n3870);
  and g2560 (n3873, n_1242, n3872);
  and g2561 (n3874, pi0299, n_1237);
  not g2562 (n_1243, n3768);
  not g2563 (n_1244, n3874);
  and g2564 (n3875, n_1243, n_1244);
  and g2565 (n3876, n_841, n3875);
  and g2566 (n3877, n_251, n3875);
  and g2567 (n3878, pi0299, n_1238);
  not g2568 (n_1245, n3878);
  and g2569 (n3879, n_1243, n_1245);
  and g2570 (n3880, n2625, n3879);
  not g2571 (n_1246, n3877);
  not g2572 (n_1247, n3880);
  and g2573 (n3881, n_1246, n_1247);
  not g2574 (n_1248, n3881);
  and g2575 (n3882, n2533, n_1248);
  and g2576 (n3883, n_257, n3875);
  not g2577 (n_1249, n3883);
  and g2578 (n3884, pi0092, n_1249);
  not g2579 (n_1250, n3882);
  and g2580 (n3885, n_1250, n3884);
  and g2581 (n3886, pi0075, n3875);
  and g2582 (n3887, pi0087, n3881);
  and g2583 (n3888, pi0038, n3875);
  not g2584 (n_1251, n3879);
  and g2585 (n3889, pi0039, n_1251);
  and g2586 (n3890, n_937, n3721);
  and g2587 (n3891, n_268, n3499);
  and g2588 (n3892, pi0146, n_1174);
  not g2589 (n_1252, n3891);
  and g2590 (n3893, pi0284, n_1252);
  not g2591 (n_1253, n3892);
  and g2592 (n3894, n_1253, n3893);
  and g2593 (n3895, n_268, n_1170);
  and g2594 (n3896, n_879, n3895);
  not g2595 (n_1254, n3894);
  not g2596 (n_1255, n3896);
  and g2597 (n3897, n_1254, n_1255);
  not g2598 (n_1256, n3897);
  and g2599 (n3898, n_188, n_1256);
  not g2600 (n_1257, n3890);
  not g2601 (n_1258, n3898);
  and g2602 (n3899, n_1257, n_1258);
  not g2603 (n_1259, n3899);
  and g2604 (n3900, n_20, n_1259);
  not g2605 (n_1260, n3900);
  and g2606 (n3901, n3716, n_1260);
  not g2607 (n_1261, n3901);
  and g2608 (n3902, n_1130, n_1261);
  not g2609 (n_1262, n3902);
  and g2610 (n3903, n_36, n_1262);
  not g2611 (n_1263, n3903);
  and g2612 (n3904, n3792, n_1263);
  not g2613 (n_1264, n3904);
  and g2614 (n3905, n3813, n_1264);
  not g2615 (n_1265, n3889);
  and g2616 (n3906, n_161, n_1265);
  not g2617 (n_1266, n3905);
  and g2618 (n3907, n_1266, n3906);
  not g2619 (n_1267, n3888);
  and g2620 (n3908, n_164, n_1267);
  not g2621 (n_1268, n3907);
  and g2622 (n3909, n_1268, n3908);
  and g2623 (n3910, n_260, n3875);
  and g2624 (n3911, n_1120, n_1200);
  not g2625 (n_1269, n3911);
  and g2626 (n3912, n_20, n_1269);
  not g2627 (n_1270, n3912);
  and g2628 (n3913, n3716, n_1270);
  not g2629 (n_1271, n3913);
  and g2630 (n3914, n_1130, n_1271);
  not g2631 (n_1272, n3914);
  and g2632 (n3915, n_36, n_1272);
  not g2633 (n_1273, n3915);
  and g2634 (n3916, n_1132, n_1273);
  not g2635 (n_1274, n3916);
  and g2636 (n3917, pi0299, n_1274);
  and g2637 (n3918, n2530, n_1243);
  not g2638 (n_1275, n3917);
  and g2639 (n3919, n_1275, n3918);
  not g2640 (n_1276, n3910);
  and g2641 (n3920, pi0100, n_1276);
  not g2642 (n_1277, n3919);
  and g2643 (n3921, n_1277, n3920);
  not g2644 (n_1278, n3909);
  not g2645 (n_1279, n3921);
  and g2646 (n3922, n_1278, n_1279);
  not g2647 (n_1280, n3922);
  and g2648 (n3923, n_172, n_1280);
  not g2649 (n_1281, n3887);
  and g2650 (n3924, n_171, n_1281);
  not g2651 (n_1282, n3923);
  and g2652 (n3925, n_1282, n3924);
  not g2653 (n_1283, n3886);
  and g2654 (n3926, n_174, n_1283);
  not g2655 (n_1284, n3925);
  and g2656 (n3927, n_1284, n3926);
  not g2657 (n_1285, n3885);
  and g2658 (n3928, n2532, n_1285);
  not g2659 (n_1286, n3927);
  and g2660 (n3929, n_1286, n3928);
  not g2661 (n_1287, n3876);
  and g2662 (n3930, n_176, n_1287);
  not g2663 (n_1288, n3929);
  and g2664 (n3931, n_1288, n3930);
  not g2665 (n_1289, n3873);
  and g2666 (n3932, n_157, n_1289);
  not g2667 (n_1290, n3931);
  and g2668 (n3933, n_1290, n3932);
  not g2669 (n_1291, n3869);
  and g2670 (n3934, n_158, n_1291);
  not g2671 (n_1292, n3933);
  and g2672 (n3935, n_1292, n3934);
  and g2678 (n3939, pi0238, n3861);
  not g2679 (n_1295, n3939);
  and g2680 (n3940, n_824, n_1295);
  and g2681 (n3941, n3733, n3940);
  not g2682 (n_1296, n3853);
  not g2683 (n_1297, n3941);
  and g2684 (n3942, n_1296, n_1297);
  not g2685 (n_1298, n3938);
  and g2686 (po0156, n_1298, n3942);
  and g2687 (n3944, pi0215, pi1142);
  and g2688 (n3945, pi0216, pi0277);
  not g2689 (n_1301, n3945);
  and g2690 (n3946, n_26, n_1301);
  and g2691 (n3947, pi0172, n_188);
  and g2692 (n3948, n_180, pi0172);
  and g2693 (n3949, pi0262, n_145);
  and g2694 (n3950, pi0105, n3949);
  not g2695 (n_1304, n3948);
  not g2696 (n_1305, n3950);
  and g2697 (n3951, n_1304, n_1305);
  not g2698 (n_1306, n3951);
  and g2699 (n3952, pi0228, n_1306);
  not g2700 (n_1307, n3947);
  not g2701 (n_1308, n3952);
  and g2702 (n3953, n_1307, n_1308);
  not g2703 (n_1309, n3953);
  and g2704 (n3954, n_20, n_1309);
  not g2705 (n_1310, n3954);
  and g2706 (n3955, n3946, n_1310);
  not g2707 (n_1311, pi1142);
  and g2708 (n3956, n_1311, n_29);
  not g2709 (n_1313, pi0932);
  and g2710 (n3957, n_1313, n2452);
  not g2711 (n_1314, n3956);
  and g2712 (n3958, pi0221, n_1314);
  not g2713 (n_1315, n3957);
  and g2714 (n3959, n_1315, n3958);
  not g2715 (n_1316, n3955);
  not g2716 (n_1317, n3959);
  and g2717 (n3960, n_1316, n_1317);
  not g2718 (n_1318, n3960);
  and g2719 (n3961, n_36, n_1318);
  not g2720 (n_1319, n3944);
  not g2721 (n_1320, n3961);
  and g2722 (n3962, n_1319, n_1320);
  not g2723 (n_1321, n3962);
  and g2724 (n3963, n_909, n_1321);
  not g2725 (n_1322, n3963);
  and g2726 (n3964, n_824, n_1322);
  and g2727 (n3965, n_826, n_1322);
  not g2728 (n_1323, pi0262);
  and g2729 (n3966, n_1323, n2521);
  not g2730 (n_1324, n3335);
  and g2731 (n3967, n_1324, n_1307);
  not g2732 (n_1325, n3966);
  not g2733 (n_1326, n3967);
  and g2734 (n3968, n_1325, n_1326);
  and g2735 (n3969, n_997, n_1308);
  not g2736 (n_1327, n3968);
  and g2737 (n3970, n_1327, n3969);
  not g2738 (n_1328, n3970);
  and g2739 (n3971, n_20, n_1328);
  not g2740 (n_1329, n3971);
  and g2741 (n3972, n3946, n_1329);
  not g2742 (n_1330, n3972);
  and g2743 (n3973, n_1317, n_1330);
  not g2744 (n_1331, n3973);
  and g2745 (n3974, n_36, n_1331);
  not g2746 (n_1332, n3974);
  and g2747 (n3975, n_1319, n_1332);
  and g2748 (n3976, n3331, n3975);
  not g2749 (n_1333, n3965);
  and g2750 (n3977, pi0062, n_1333);
  not g2751 (n_1334, n3976);
  and g2752 (n3978, n_1334, n3977);
  not g2753 (n_1335, n3975);
  and g2754 (n3979, n2537, n_1335);
  and g2755 (n3980, n_179, n3963);
  not g2756 (n_1336, n3980);
  and g2757 (n3981, pi0056, n_1336);
  not g2758 (n_1337, n3979);
  and g2759 (n3982, n_1337, n3981);
  and g2760 (n3983, n_204, n_1322);
  and g2761 (n3984, n2572, n3975);
  not g2762 (n_1338, n3983);
  and g2763 (n3985, pi0055, n_1338);
  not g2764 (n_1339, n3984);
  and g2765 (n3986, n_1339, n3985);
  and g2766 (n3987, pi0223, pi1142);
  and g2767 (n3988, pi0224, pi0277);
  not g2768 (n_1340, n3988);
  and g2769 (n3989, n_226, n_1340);
  and g2770 (n3990, n_219, n3949);
  not g2771 (n_1341, n3990);
  and g2772 (n3991, n3989, n_1341);
  and g2773 (n3992, n_1311, n_221);
  and g2774 (n3993, n_1313, n2591);
  not g2775 (n_1342, n3992);
  and g2776 (n3994, pi0222, n_1342);
  not g2777 (n_1343, n3993);
  and g2778 (n3995, n_1343, n3994);
  not g2779 (n_1344, n3991);
  not g2780 (n_1345, n3995);
  and g2781 (n3996, n_1344, n_1345);
  not g2782 (n_1346, n3996);
  and g2783 (n3997, n_223, n_1346);
  not g2784 (n_1347, n3987);
  not g2785 (n_1348, n3997);
  and g2786 (n3998, n_1347, n_1348);
  not g2787 (n_1349, n3998);
  and g2788 (n3999, n_234, n_1349);
  and g2789 (n4000, n_1160, n3999);
  and g2790 (n4001, pi0299, n3963);
  not g2791 (n_1350, n4000);
  not g2792 (n_1351, n4001);
  and g2793 (n4002, n_1350, n_1351);
  and g2794 (n4003, n_841, n4002);
  and g2795 (n4004, n_251, n4002);
  and g2796 (n4005, pi0299, n_1335);
  not g2797 (n_1352, n4005);
  and g2798 (n4006, n_1350, n_1352);
  and g2799 (n4007, n2625, n4006);
  not g2800 (n_1353, n4004);
  not g2801 (n_1354, n4007);
  and g2802 (n4008, n_1353, n_1354);
  not g2803 (n_1355, n4008);
  and g2804 (n4009, n2533, n_1355);
  and g2805 (n4010, n_257, n4002);
  not g2806 (n_1356, n4010);
  and g2807 (n4011, pi0092, n_1356);
  not g2808 (n_1357, n4009);
  and g2809 (n4012, n_1357, n4011);
  and g2810 (n4013, pi0075, n4002);
  and g2811 (n4014, pi0087, n4008);
  and g2812 (n4015, pi0038, n4002);
  not g2813 (n_1358, n4006);
  and g2814 (n4016, pi0039, n_1358);
  and g2815 (n4017, n_234, n_1347);
  and g2816 (n4018, n_1323, n3488);
  not g2817 (n_1359, n4018);
  and g2818 (n4019, n_219, n_1359);
  not g2819 (n_1360, n4019);
  and g2820 (n4020, n3989, n_1360);
  not g2821 (n_1361, n4020);
  and g2822 (n4021, n_1345, n_1361);
  and g2823 (n4022, n4017, n4021);
  and g2824 (n4023, pi0299, n_1319);
  and g2825 (n4024, pi0262, n3416);
  and g2826 (n4025, n_1323, n3499);
  not g2827 (n_1362, pi0172);
  not g2828 (n_1363, n4025);
  and g2829 (n4026, n_1362, n_1363);
  and g2830 (n4027, pi0172, n_1323);
  and g2831 (n4028, n3508, n4027);
  not g2832 (n_1364, n4026);
  not g2833 (n_1365, n4028);
  and g2834 (n4029, n_1364, n_1365);
  not g2835 (n_1366, n4024);
  and g2836 (n4030, n_188, n_1366);
  not g2837 (n_1367, n4029);
  and g2838 (n4031, n_1367, n4030);
  and g2839 (n4032, n_929, n3950);
  and g2840 (n4033, pi0228, n_1304);
  not g2841 (n_1368, n4032);
  and g2842 (n4034, n_1368, n4033);
  and g2843 (n4035, n_937, n4034);
  not g2844 (n_1369, n4035);
  and g2845 (n4036, n_20, n_1369);
  not g2846 (n_1370, n4031);
  and g2847 (n4037, n_1370, n4036);
  not g2848 (n_1371, n4037);
  and g2849 (n4038, n3946, n_1371);
  not g2850 (n_1372, n4038);
  and g2851 (n4039, n_1317, n_1372);
  not g2852 (n_1373, n4039);
  and g2853 (n4040, n_36, n_1373);
  not g2854 (n_1374, n4040);
  and g2855 (n4041, n4023, n_1374);
  and g2856 (n4042, n_936, n3989);
  not g2857 (n_1375, n4042);
  and g2858 (n4043, n4021, n_1375);
  not g2859 (n_1376, n4043);
  and g2860 (n4044, n_223, n_1376);
  not g2861 (n_1377, n4044);
  and g2862 (n4045, n4017, n_1377);
  not g2863 (n_1378, n4045);
  and g2864 (n4046, n_162, n_1378);
  not g2865 (n_1379, n4022);
  and g2866 (n4047, n_1379, n4046);
  not g2867 (n_1380, n4041);
  and g2868 (n4048, n_1380, n4047);
  not g2869 (n_1381, n4016);
  and g2870 (n4049, n_161, n_1381);
  not g2871 (n_1382, n4048);
  and g2872 (n4050, n_1382, n4049);
  not g2873 (n_1383, n4015);
  and g2874 (n4051, n_164, n_1383);
  not g2875 (n_1384, n4050);
  and g2876 (n4052, n_1384, n4051);
  and g2877 (n4053, n_260, n4002);
  and g2878 (n4054, n_1323, n3394);
  and g2879 (n4055, n_1046, n_1307);
  not g2880 (n_1385, n4054);
  not g2881 (n_1386, n4055);
  and g2882 (n4056, n_1385, n_1386);
  not g2883 (n_1387, n4056);
  and g2884 (n4057, n3969, n_1387);
  not g2885 (n_1388, n4057);
  and g2886 (n4058, n_20, n_1388);
  not g2887 (n_1389, n4058);
  and g2888 (n4059, n3946, n_1389);
  not g2889 (n_1390, n4059);
  and g2890 (n4060, n_1317, n_1390);
  not g2891 (n_1391, n4060);
  and g2892 (n4061, n_36, n_1391);
  not g2893 (n_1392, n4061);
  and g2894 (n4062, n_1319, n_1392);
  not g2895 (n_1393, n4062);
  and g2896 (n4063, pi0299, n_1393);
  and g2897 (n4064, n2530, n_1350);
  not g2898 (n_1394, n4063);
  and g2899 (n4065, n_1394, n4064);
  not g2900 (n_1395, n4053);
  and g2901 (n4066, pi0100, n_1395);
  not g2902 (n_1396, n4065);
  and g2903 (n4067, n_1396, n4066);
  not g2904 (n_1397, n4052);
  not g2905 (n_1398, n4067);
  and g2906 (n4068, n_1397, n_1398);
  not g2907 (n_1399, n4068);
  and g2908 (n4069, n_172, n_1399);
  not g2909 (n_1400, n4014);
  and g2910 (n4070, n_171, n_1400);
  not g2911 (n_1401, n4069);
  and g2912 (n4071, n_1401, n4070);
  not g2913 (n_1402, n4013);
  and g2914 (n4072, n_174, n_1402);
  not g2915 (n_1403, n4071);
  and g2916 (n4073, n_1403, n4072);
  not g2917 (n_1404, n4012);
  and g2918 (n4074, n2532, n_1404);
  not g2919 (n_1405, n4073);
  and g2920 (n4075, n_1405, n4074);
  not g2921 (n_1406, n4003);
  and g2922 (n4076, n_176, n_1406);
  not g2923 (n_1407, n4075);
  and g2924 (n4077, n_1407, n4076);
  not g2925 (n_1408, n3986);
  and g2926 (n4078, n_157, n_1408);
  not g2927 (n_1409, n4077);
  and g2928 (n4079, n_1409, n4078);
  not g2929 (n_1410, n3982);
  and g2930 (n4080, n_158, n_1410);
  not g2931 (n_1411, n4079);
  and g2932 (n4081, n_1411, n4080);
  not g2933 (n_1412, n3978);
  and g2934 (n4082, n3328, n_1412);
  not g2935 (n_1413, n4081);
  and g2936 (n4083, n_1413, n4082);
  not g2937 (n_1415, pi0249);
  not g2938 (n_1416, n3964);
  and g2939 (n4084, n_1415, n_1416);
  not g2940 (n_1417, n4083);
  and g2941 (n4085, n_1417, n4084);
  and g2942 (n4086, n_824, n3962);
  and g2943 (n4087, n_826, n3962);
  and g2944 (n4088, n_1308, n_1327);
  not g2945 (n_1418, n4088);
  and g2946 (n4089, n_20, n_1418);
  not g2947 (n_1419, n4089);
  and g2948 (n4090, n3946, n_1419);
  not g2949 (n_1420, n4090);
  and g2950 (n4091, n_1317, n_1420);
  not g2951 (n_1421, n4091);
  and g2952 (n4092, n_36, n_1421);
  not g2953 (n_1422, n4092);
  and g2954 (n4093, n_1319, n_1422);
  and g2955 (n4094, n3331, n4093);
  not g2956 (n_1423, n4087);
  and g2957 (n4095, pi0062, n_1423);
  not g2958 (n_1424, n4094);
  and g2959 (n4096, n_1424, n4095);
  and g2960 (n4097, n_179, n_1321);
  not g2961 (n_1425, n4093);
  and g2962 (n4098, n2537, n_1425);
  not g2963 (n_1426, n4097);
  and g2964 (n4099, pi0056, n_1426);
  not g2965 (n_1427, n4098);
  and g2966 (n4100, n_1427, n4099);
  and g2967 (n4101, n_204, n3962);
  and g2968 (n4102, n2572, n4093);
  not g2969 (n_1428, n4101);
  and g2970 (n4103, pi0055, n_1428);
  not g2971 (n_1429, n4102);
  and g2972 (n4104, n_1429, n4103);
  and g2973 (n4105, pi0299, n_1321);
  not g2974 (n_1430, n3999);
  not g2975 (n_1431, n4105);
  and g2976 (n4106, n_1430, n_1431);
  and g2977 (n4107, n_841, n4106);
  and g2978 (n4108, n_251, n4106);
  and g2979 (n4109, pi0299, n_1425);
  not g2980 (n_1432, n4109);
  and g2981 (n4110, n_1430, n_1432);
  and g2982 (n4111, n2625, n4110);
  not g2983 (n_1433, n4108);
  not g2984 (n_1434, n4111);
  and g2985 (n4112, n_1433, n_1434);
  not g2986 (n_1435, n4112);
  and g2987 (n4113, n2533, n_1435);
  and g2988 (n4114, n_257, n4106);
  not g2989 (n_1436, n4114);
  and g2990 (n4115, pi0092, n_1436);
  not g2991 (n_1437, n4113);
  and g2992 (n4116, n_1437, n4115);
  and g2993 (n4117, pi0075, n4106);
  and g2994 (n4118, pi0087, n4112);
  and g2995 (n4119, pi0038, n4106);
  not g2996 (n_1438, n4110);
  and g2997 (n4120, pi0039, n_1438);
  and g2998 (n4121, pi0262, n3508);
  not g2999 (n_1439, n4121);
  and g3000 (n4122, n_1362, n_1439);
  and g3001 (n4123, pi0262, n_938);
  and g3002 (n4124, n_1323, n_879);
  not g3003 (n_1440, n4123);
  and g3004 (n4125, pi0172, n_1440);
  not g3005 (n_1441, n4124);
  and g3006 (n4126, n_1441, n4125);
  not g3007 (n_1442, n4122);
  not g3008 (n_1443, n4126);
  and g3009 (n4127, n_1442, n_1443);
  not g3010 (n_1444, n4127);
  and g3011 (n4128, n_188, n_1444);
  not g3012 (n_1445, n4034);
  and g3013 (n4129, n_20, n_1445);
  not g3014 (n_1446, n4128);
  and g3015 (n4130, n_1446, n4129);
  not g3016 (n_1447, n4130);
  and g3017 (n4131, n3946, n_1447);
  not g3018 (n_1448, n4131);
  and g3019 (n4132, n_1317, n_1448);
  not g3020 (n_1449, n4132);
  and g3021 (n4133, n_36, n_1449);
  not g3022 (n_1450, n4133);
  and g3023 (n4134, n4023, n_1450);
  not g3024 (n_1451, n4134);
  and g3025 (n4135, n4046, n_1451);
  not g3026 (n_1452, n4120);
  and g3027 (n4136, n_161, n_1452);
  not g3028 (n_1453, n4135);
  and g3029 (n4137, n_1453, n4136);
  not g3030 (n_1454, n4119);
  and g3031 (n4138, n_164, n_1454);
  not g3032 (n_1455, n4137);
  and g3033 (n4139, n_1455, n4138);
  and g3034 (n4140, n_260, n4106);
  and g3035 (n4141, n_1308, n_1387);
  not g3036 (n_1456, n4141);
  and g3037 (n4142, n_20, n_1456);
  not g3038 (n_1457, n4142);
  and g3039 (n4143, n3946, n_1457);
  not g3040 (n_1458, n4143);
  and g3041 (n4144, n_1317, n_1458);
  not g3042 (n_1459, n4144);
  and g3043 (n4145, n_36, n_1459);
  not g3044 (n_1460, n4145);
  and g3045 (n4146, n_1319, n_1460);
  not g3046 (n_1461, n4146);
  and g3047 (n4147, pi0299, n_1461);
  and g3048 (n4148, n2530, n_1430);
  not g3049 (n_1462, n4147);
  and g3050 (n4149, n_1462, n4148);
  not g3051 (n_1463, n4140);
  and g3052 (n4150, pi0100, n_1463);
  not g3053 (n_1464, n4149);
  and g3054 (n4151, n_1464, n4150);
  not g3055 (n_1465, n4139);
  not g3056 (n_1466, n4151);
  and g3057 (n4152, n_1465, n_1466);
  not g3058 (n_1467, n4152);
  and g3059 (n4153, n_172, n_1467);
  not g3060 (n_1468, n4118);
  and g3061 (n4154, n_171, n_1468);
  not g3062 (n_1469, n4153);
  and g3063 (n4155, n_1469, n4154);
  not g3064 (n_1470, n4117);
  and g3065 (n4156, n_174, n_1470);
  not g3066 (n_1471, n4155);
  and g3067 (n4157, n_1471, n4156);
  not g3068 (n_1472, n4116);
  and g3069 (n4158, n2532, n_1472);
  not g3070 (n_1473, n4157);
  and g3071 (n4159, n_1473, n4158);
  not g3072 (n_1474, n4107);
  and g3073 (n4160, n_176, n_1474);
  not g3074 (n_1475, n4159);
  and g3075 (n4161, n_1475, n4160);
  not g3076 (n_1476, n4104);
  and g3077 (n4162, n_157, n_1476);
  not g3078 (n_1477, n4161);
  and g3079 (n4163, n_1477, n4162);
  not g3080 (n_1478, n4100);
  and g3081 (n4164, n_158, n_1478);
  not g3082 (n_1479, n4163);
  and g3083 (n4165, n_1479, n4164);
  not g3084 (n_1480, n4096);
  and g3085 (n4166, n3328, n_1480);
  not g3086 (n_1481, n4165);
  and g3087 (n4167, n_1481, n4166);
  not g3088 (n_1482, n4086);
  and g3089 (n4168, pi0249, n_1482);
  not g3090 (n_1483, n4167);
  and g3091 (n4169, n_1483, n4168);
  or g3092 (po0157, n4085, n4169);
  and g3093 (n4171, pi0215, pi1141);
  and g3094 (n4172, pi0216, pi0270);
  not g3095 (n_1486, n4172);
  and g3096 (n4173, n_26, n_1486);
  and g3097 (n4174, n_180, pi0171);
  and g3098 (n4175, pi0861, n_145);
  not g3099 (n_1489, n4175);
  and g3100 (n4176, pi0105, n_1489);
  not g3101 (n_1490, n4174);
  and g3102 (n4177, pi0228, n_1490);
  not g3103 (n_1491, n4176);
  and g3104 (n4178, n_1491, n4177);
  not g3105 (n_1492, n4178);
  and g3106 (n4179, n_20, n_1492);
  not g3107 (n_1493, pi0171);
  and g3108 (n4180, n_1493, n_188);
  not g3109 (n_1494, n4180);
  and g3110 (n4181, n4179, n_1494);
  not g3111 (n_1495, n4181);
  and g3112 (n4182, n4173, n_1495);
  not g3113 (n_1496, pi1141);
  and g3114 (n4183, n_1496, n_29);
  not g3115 (n_1498, pi0935);
  and g3116 (n4184, n_1498, n2452);
  not g3117 (n_1499, n4183);
  and g3118 (n4185, pi0221, n_1499);
  not g3119 (n_1500, n4184);
  and g3120 (n4186, n_1500, n4185);
  not g3121 (n_1501, n4182);
  not g3122 (n_1502, n4186);
  and g3123 (n4187, n_1501, n_1502);
  not g3124 (n_1503, n4187);
  and g3125 (n4188, n_36, n_1503);
  not g3126 (n_1504, n4171);
  not g3127 (n_1505, n4188);
  and g3128 (n4189, n_1504, n_1505);
  and g3129 (n4190, n_826, n4189);
  not g3130 (n_1506, pi0861);
  and g3131 (n4191, n_1506, n2521);
  and g3132 (n4192, pi0171, n_207);
  not g3133 (n_1507, n4191);
  and g3134 (n4193, n_188, n_1507);
  not g3135 (n_1508, n4192);
  and g3136 (n4194, n_1508, n4193);
  not g3137 (n_1509, n4194);
  and g3138 (n4195, n4179, n_1509);
  not g3139 (n_1510, n4195);
  and g3140 (n4196, n4173, n_1510);
  not g3141 (n_1511, n4196);
  and g3142 (n4197, n_1502, n_1511);
  not g3143 (n_1512, n4197);
  and g3144 (n4198, n_36, n_1512);
  not g3145 (n_1513, n4198);
  and g3146 (n4199, n_1504, n_1513);
  and g3147 (n4200, n3331, n4199);
  not g3148 (n_1514, n4190);
  and g3149 (n4201, pi0062, n_1514);
  not g3150 (n_1515, n4200);
  and g3151 (n4202, n_1515, n4201);
  not g3152 (n_1516, n4189);
  and g3153 (n4203, n_179, n_1516);
  not g3154 (n_1517, n4199);
  and g3155 (n4204, n2537, n_1517);
  not g3156 (n_1518, n4203);
  and g3157 (n4205, pi0056, n_1518);
  not g3158 (n_1519, n4204);
  and g3159 (n4206, n_1519, n4205);
  and g3160 (n4207, n_204, n4189);
  and g3161 (n4208, n2572, n4199);
  not g3162 (n_1520, n4207);
  and g3163 (n4209, pi0055, n_1520);
  not g3164 (n_1521, n4208);
  and g3165 (n4210, n_1521, n4209);
  and g3166 (n4211, pi0223, pi1141);
  and g3167 (n4212, pi0224, pi0270);
  not g3168 (n_1522, n4212);
  and g3169 (n4213, n_226, n_1522);
  and g3170 (n4214, n_219, n_1489);
  not g3171 (n_1523, n4214);
  and g3172 (n4215, n4213, n_1523);
  and g3173 (n4216, n_1496, n_221);
  and g3174 (n4217, n_1498, n2591);
  not g3175 (n_1524, n4216);
  and g3176 (n4218, pi0222, n_1524);
  not g3177 (n_1525, n4217);
  and g3178 (n4219, n_1525, n4218);
  not g3179 (n_1526, n4215);
  not g3180 (n_1527, n4219);
  and g3181 (n4220, n_1526, n_1527);
  not g3182 (n_1528, n4220);
  and g3183 (n4221, n_223, n_1528);
  not g3184 (n_1529, n4211);
  not g3185 (n_1530, n4221);
  and g3186 (n4222, n_1529, n_1530);
  not g3187 (n_1531, n4222);
  and g3188 (n4223, n_234, n_1531);
  and g3189 (n4224, pi0299, n_1516);
  not g3190 (n_1532, n4223);
  not g3191 (n_1533, n4224);
  and g3192 (n4225, n_1532, n_1533);
  and g3193 (n4226, n_841, n4225);
  and g3194 (n4227, n_251, n4225);
  and g3195 (n4228, pi0299, n_1517);
  not g3196 (n_1534, n4228);
  and g3197 (n4229, n_1532, n_1534);
  and g3198 (n4230, n2625, n4229);
  not g3199 (n_1535, n4227);
  not g3200 (n_1536, n4230);
  and g3201 (n4231, n_1535, n_1536);
  not g3202 (n_1537, n4231);
  and g3203 (n4232, n2533, n_1537);
  and g3204 (n4233, n_257, n4225);
  not g3205 (n_1538, n4233);
  and g3206 (n4234, pi0092, n_1538);
  not g3207 (n_1539, n4232);
  and g3208 (n4235, n_1539, n4234);
  and g3209 (n4236, pi0075, n4225);
  and g3210 (n4237, pi0087, n4231);
  and g3211 (n4238, pi0038, n4225);
  not g3212 (n_1540, n4229);
  and g3213 (n4239, pi0039, n_1540);
  and g3214 (n4240, n_234, n_1529);
  and g3215 (n4241, pi0861, n3488);
  not g3216 (n_1541, n4241);
  and g3217 (n4242, n_219, n_1541);
  not g3218 (n_1542, n4242);
  and g3219 (n4243, n4213, n_1542);
  not g3220 (n_1543, n4243);
  and g3221 (n4244, n_1527, n_1543);
  and g3222 (n4245, n4240, n4244);
  and g3223 (n4246, pi0299, n_1504);
  and g3224 (n4247, pi0861, n3499);
  not g3225 (n_1544, n4247);
  and g3226 (n4248, n_1493, n_1544);
  and g3227 (n4249, pi0171, n3508);
  not g3228 (n_1545, n4248);
  not g3229 (n_1546, n4249);
  and g3230 (n4250, n_1545, n_1546);
  not g3231 (n_1547, n4250);
  and g3232 (n4251, pi0861, n_1547);
  and g3233 (n4252, n_879, n4248);
  not g3234 (n_1548, n4251);
  not g3235 (n_1549, n4252);
  and g3236 (n4253, n_1548, n_1549);
  not g3237 (n_1550, n4253);
  and g3238 (n4254, n_188, n_1550);
  and g3239 (n4255, n_937, n4178);
  not g3240 (n_1551, n4255);
  and g3241 (n4256, n_20, n_1551);
  not g3242 (n_1552, n4254);
  and g3243 (n4257, n_1552, n4256);
  not g3244 (n_1553, n4257);
  and g3245 (n4258, n4173, n_1553);
  not g3246 (n_1554, n4258);
  and g3247 (n4259, n_1502, n_1554);
  not g3248 (n_1555, n4259);
  and g3249 (n4260, n_36, n_1555);
  not g3250 (n_1556, n4260);
  and g3251 (n4261, n4246, n_1556);
  and g3252 (n4262, n_936, n4213);
  not g3253 (n_1557, n4262);
  and g3254 (n4263, n4244, n_1557);
  not g3255 (n_1558, n4263);
  and g3256 (n4264, n_223, n_1558);
  not g3257 (n_1559, n4264);
  and g3258 (n4265, n4240, n_1559);
  not g3259 (n_1560, n4265);
  and g3260 (n4266, n_162, n_1560);
  not g3261 (n_1561, n4245);
  and g3262 (n4267, n_1561, n4266);
  not g3263 (n_1562, n4261);
  and g3264 (n4268, n_1562, n4267);
  not g3265 (n_1563, n4239);
  and g3266 (n4269, n_161, n_1563);
  not g3267 (n_1564, n4268);
  and g3268 (n4270, n_1564, n4269);
  not g3269 (n_1565, n4238);
  and g3270 (n4271, n_164, n_1565);
  not g3271 (n_1566, n4270);
  and g3272 (n4272, n_1566, n4271);
  and g3273 (n4273, n_260, n4225);
  and g3274 (n4274, n_1506, n3394);
  not g3275 (n_1567, n3394);
  and g3276 (n4275, pi0171, n_1567);
  not g3277 (n_1568, n4274);
  and g3278 (n4276, n_188, n_1568);
  not g3279 (n_1569, n4275);
  and g3280 (n4277, n_1569, n4276);
  not g3281 (n_1570, n4277);
  and g3282 (n4278, n4179, n_1570);
  not g3283 (n_1571, n4278);
  and g3284 (n4279, n4173, n_1571);
  not g3285 (n_1572, n4279);
  and g3286 (n4280, n_1502, n_1572);
  not g3287 (n_1573, n4280);
  and g3288 (n4281, n_36, n_1573);
  not g3289 (n_1574, n4281);
  and g3290 (n4282, n_1504, n_1574);
  not g3291 (n_1575, n4282);
  and g3292 (n4283, pi0299, n_1575);
  and g3293 (n4284, n2530, n_1532);
  not g3294 (n_1576, n4283);
  and g3295 (n4285, n_1576, n4284);
  not g3296 (n_1577, n4273);
  and g3297 (n4286, pi0100, n_1577);
  not g3298 (n_1578, n4285);
  and g3299 (n4287, n_1578, n4286);
  not g3300 (n_1579, n4272);
  not g3301 (n_1580, n4287);
  and g3302 (n4288, n_1579, n_1580);
  not g3303 (n_1581, n4288);
  and g3304 (n4289, n_172, n_1581);
  not g3305 (n_1582, n4237);
  and g3306 (n4290, n_171, n_1582);
  not g3307 (n_1583, n4289);
  and g3308 (n4291, n_1583, n4290);
  not g3309 (n_1584, n4236);
  and g3310 (n4292, n_174, n_1584);
  not g3311 (n_1585, n4291);
  and g3312 (n4293, n_1585, n4292);
  not g3313 (n_1586, n4235);
  and g3314 (n4294, n2532, n_1586);
  not g3315 (n_1587, n4293);
  and g3316 (n4295, n_1587, n4294);
  not g3317 (n_1588, n4226);
  and g3318 (n4296, n_176, n_1588);
  not g3319 (n_1589, n4295);
  and g3320 (n4297, n_1589, n4296);
  not g3321 (n_1590, n4210);
  and g3322 (n4298, n_157, n_1590);
  not g3323 (n_1591, n4297);
  and g3324 (n4299, n_1591, n4298);
  not g3325 (n_1592, n4206);
  and g3326 (n4300, n_158, n_1592);
  not g3327 (n_1593, n4299);
  and g3328 (n4301, n_1593, n4300);
  not g3329 (n_1595, pi0241);
  and g3335 (n4305, n_997, n4179);
  and g3336 (n4306, n_1509, n4305);
  not g3337 (n_1598, n4306);
  and g3338 (n4307, n4173, n_1598);
  not g3339 (n_1599, n4307);
  and g3340 (n4308, n_1502, n_1599);
  not g3341 (n_1600, n4308);
  and g3342 (n4309, n_36, n_1600);
  not g3343 (n_1601, n4309);
  and g3344 (n4310, n_1504, n_1601);
  and g3345 (n4311, n3331, n4310);
  and g3346 (n4312, n3556, n_1486);
  not g3347 (n_1602, n4312);
  and g3348 (n4313, n4189, n_1602);
  and g3349 (n4314, n_826, n4313);
  not g3350 (n_1603, n4314);
  and g3351 (n4315, pi0062, n_1603);
  not g3352 (n_1604, n4311);
  and g3353 (n4316, n_1604, n4315);
  not g3354 (n_1605, n4313);
  and g3355 (n4317, n_179, n_1605);
  not g3356 (n_1606, n4310);
  and g3357 (n4318, n2537, n_1606);
  not g3358 (n_1607, n4317);
  and g3359 (n4319, pi0056, n_1607);
  not g3360 (n_1608, n4318);
  and g3361 (n4320, n_1608, n4319);
  and g3362 (n4321, n2572, n4310);
  and g3363 (n4322, n_204, n4313);
  not g3364 (n_1609, n4322);
  and g3365 (n4323, pi0055, n_1609);
  not g3366 (n_1610, n4321);
  and g3367 (n4324, n_1610, n4323);
  and g3368 (n4325, n_921, n_1532);
  and g3369 (n4326, pi0299, n_1605);
  not g3370 (n_1611, n4326);
  and g3371 (n4327, n4325, n_1611);
  and g3372 (n4328, n_841, n4327);
  and g3373 (n4329, n_251, n4327);
  and g3374 (n4330, pi0299, n_1606);
  not g3375 (n_1612, n4330);
  and g3376 (n4331, n4325, n_1612);
  and g3377 (n4332, n2625, n4331);
  not g3378 (n_1613, n4329);
  not g3379 (n_1614, n4332);
  and g3380 (n4333, n_1613, n_1614);
  not g3381 (n_1615, n4333);
  and g3382 (n4334, n2533, n_1615);
  and g3383 (n4335, n_257, n4327);
  not g3384 (n_1616, n4335);
  and g3385 (n4336, pi0092, n_1616);
  not g3386 (n_1617, n4334);
  and g3387 (n4337, n_1617, n4336);
  and g3388 (n4338, pi0075, n4327);
  and g3389 (n4339, pi0087, n4333);
  and g3390 (n4340, pi0038, n4327);
  not g3391 (n_1618, n4331);
  and g3392 (n4341, pi0039, n_1618);
  and g3393 (n4342, n_1506, n3508);
  not g3394 (n_1619, n4342);
  and g3395 (n4343, n_1493, n_1619);
  and g3396 (n4344, n_1506, n_938);
  and g3397 (n4345, pi0861, n_879);
  not g3398 (n_1620, n4344);
  and g3399 (n4346, pi0171, n_1620);
  not g3400 (n_1621, n4345);
  and g3401 (n4347, n_1621, n4346);
  not g3402 (n_1622, n4343);
  not g3403 (n_1623, n4347);
  and g3404 (n4348, n_1622, n_1623);
  not g3405 (n_1624, n4348);
  and g3406 (n4349, n_188, n_1624);
  and g3407 (n4350, n_1181, n4179);
  not g3408 (n_1625, n4349);
  and g3409 (n4351, n_1625, n4350);
  not g3410 (n_1626, n4351);
  and g3411 (n4352, n4173, n_1626);
  not g3412 (n_1627, n4352);
  and g3413 (n4353, n_1502, n_1627);
  not g3414 (n_1628, n4353);
  and g3415 (n4354, n_36, n_1628);
  not g3416 (n_1629, n4354);
  and g3417 (n4355, n4246, n_1629);
  not g3418 (n_1630, n4355);
  and g3419 (n4356, n4266, n_1630);
  not g3420 (n_1631, n4341);
  and g3421 (n4357, n_161, n_1631);
  not g3422 (n_1632, n4356);
  and g3423 (n4358, n_1632, n4357);
  not g3424 (n_1633, n4340);
  and g3425 (n4359, n_164, n_1633);
  not g3426 (n_1634, n4358);
  and g3427 (n4360, n_1634, n4359);
  and g3428 (n4361, n_260, n4327);
  and g3429 (n4362, n_1570, n4305);
  not g3430 (n_1635, n4362);
  and g3431 (n4363, n4173, n_1635);
  not g3432 (n_1636, n4363);
  and g3433 (n4364, n_1502, n_1636);
  not g3434 (n_1637, n4364);
  and g3435 (n4365, n_36, n_1637);
  not g3436 (n_1638, n4365);
  and g3437 (n4366, n_1504, n_1638);
  not g3438 (n_1639, n4366);
  and g3439 (n4367, pi0299, n_1639);
  and g3440 (n4368, n2530, n4325);
  not g3441 (n_1640, n4367);
  and g3442 (n4369, n_1640, n4368);
  not g3443 (n_1641, n4361);
  and g3444 (n4370, pi0100, n_1641);
  not g3445 (n_1642, n4369);
  and g3446 (n4371, n_1642, n4370);
  not g3447 (n_1643, n4360);
  not g3448 (n_1644, n4371);
  and g3449 (n4372, n_1643, n_1644);
  not g3450 (n_1645, n4372);
  and g3451 (n4373, n_172, n_1645);
  not g3452 (n_1646, n4339);
  and g3453 (n4374, n_171, n_1646);
  not g3454 (n_1647, n4373);
  and g3455 (n4375, n_1647, n4374);
  not g3456 (n_1648, n4338);
  and g3457 (n4376, n_174, n_1648);
  not g3458 (n_1649, n4375);
  and g3459 (n4377, n_1649, n4376);
  not g3460 (n_1650, n4337);
  and g3461 (n4378, n2532, n_1650);
  not g3462 (n_1651, n4377);
  and g3463 (n4379, n_1651, n4378);
  not g3464 (n_1652, n4328);
  and g3465 (n4380, n_176, n_1652);
  not g3466 (n_1653, n4379);
  and g3467 (n4381, n_1653, n4380);
  not g3468 (n_1654, n4324);
  and g3469 (n4382, n_157, n_1654);
  not g3470 (n_1655, n4381);
  and g3471 (n4383, n_1655, n4382);
  not g3472 (n_1656, n4320);
  and g3473 (n4384, n_158, n_1656);
  not g3474 (n_1657, n4383);
  and g3475 (n4385, n_1657, n4384);
  and g3481 (n4389, pi0241, n4312);
  not g3482 (n_1660, n4389);
  and g3483 (n4390, n_824, n_1660);
  and g3484 (n4391, n4189, n4390);
  not g3485 (n_1661, n4388);
  not g3486 (n_1662, n4391);
  and g3487 (n4392, n_1661, n_1662);
  not g3488 (n_1663, n4304);
  and g3489 (po0158, n_1663, n4392);
  and g3490 (n4394, pi0215, pi1140);
  and g3491 (n4395, pi0216, pi0282);
  not g3492 (n_1666, n4395);
  and g3493 (n4396, n_26, n_1666);
  and g3494 (n4397, n_180, pi0170);
  and g3495 (n4398, pi0869, n_145);
  not g3496 (n_1669, n4398);
  and g3497 (n4399, pi0105, n_1669);
  not g3498 (n_1670, n4397);
  and g3499 (n4400, pi0228, n_1670);
  not g3500 (n_1671, n4399);
  and g3501 (n4401, n_1671, n4400);
  not g3502 (n_1672, n4401);
  and g3503 (n4402, n_20, n_1672);
  not g3504 (n_1673, pi0170);
  and g3505 (n4403, n_1673, n_188);
  not g3506 (n_1674, n4403);
  and g3507 (n4404, n4402, n_1674);
  not g3508 (n_1675, n4404);
  and g3509 (n4405, n4396, n_1675);
  not g3510 (n_1676, pi1140);
  and g3511 (n4406, n_1676, n_29);
  not g3512 (n_1678, pi0921);
  and g3513 (n4407, n_1678, n2452);
  not g3514 (n_1679, n4406);
  and g3515 (n4408, pi0221, n_1679);
  not g3516 (n_1680, n4407);
  and g3517 (n4409, n_1680, n4408);
  not g3518 (n_1681, n4405);
  not g3519 (n_1682, n4409);
  and g3520 (n4410, n_1681, n_1682);
  not g3521 (n_1683, n4410);
  and g3522 (n4411, n_36, n_1683);
  not g3523 (n_1684, n4394);
  not g3524 (n_1685, n4411);
  and g3525 (n4412, n_1684, n_1685);
  and g3526 (n4413, n_826, n4412);
  not g3527 (n_1686, pi0869);
  and g3528 (n4414, n_1686, n2521);
  and g3529 (n4415, pi0170, n_207);
  not g3530 (n_1687, n4414);
  and g3531 (n4416, n_188, n_1687);
  not g3532 (n_1688, n4415);
  and g3533 (n4417, n_1688, n4416);
  not g3534 (n_1689, n4417);
  and g3535 (n4418, n4402, n_1689);
  not g3536 (n_1690, n4418);
  and g3537 (n4419, n4396, n_1690);
  not g3538 (n_1691, n4419);
  and g3539 (n4420, n_1682, n_1691);
  not g3540 (n_1692, n4420);
  and g3541 (n4421, n_36, n_1692);
  not g3542 (n_1693, n4421);
  and g3543 (n4422, n_1684, n_1693);
  and g3544 (n4423, n3331, n4422);
  not g3545 (n_1694, n4413);
  and g3546 (n4424, pi0062, n_1694);
  not g3547 (n_1695, n4423);
  and g3548 (n4425, n_1695, n4424);
  not g3549 (n_1696, n4412);
  and g3550 (n4426, n_179, n_1696);
  not g3551 (n_1697, n4422);
  and g3552 (n4427, n2537, n_1697);
  not g3553 (n_1698, n4426);
  and g3554 (n4428, pi0056, n_1698);
  not g3555 (n_1699, n4427);
  and g3556 (n4429, n_1699, n4428);
  and g3557 (n4430, n_204, n4412);
  and g3558 (n4431, n2572, n4422);
  not g3559 (n_1700, n4430);
  and g3560 (n4432, pi0055, n_1700);
  not g3561 (n_1701, n4431);
  and g3562 (n4433, n_1701, n4432);
  and g3563 (n4434, pi0223, pi1140);
  and g3564 (n4435, pi0224, pi0282);
  not g3565 (n_1702, n4435);
  and g3566 (n4436, n_226, n_1702);
  and g3567 (n4437, n_219, n_1669);
  not g3568 (n_1703, n4437);
  and g3569 (n4438, n4436, n_1703);
  and g3570 (n4439, n_1676, n_221);
  and g3571 (n4440, n_1678, n2591);
  not g3572 (n_1704, n4439);
  and g3573 (n4441, pi0222, n_1704);
  not g3574 (n_1705, n4440);
  and g3575 (n4442, n_1705, n4441);
  not g3576 (n_1706, n4438);
  not g3577 (n_1707, n4442);
  and g3578 (n4443, n_1706, n_1707);
  not g3579 (n_1708, n4443);
  and g3580 (n4444, n_223, n_1708);
  not g3581 (n_1709, n4434);
  not g3582 (n_1710, n4444);
  and g3583 (n4445, n_1709, n_1710);
  not g3584 (n_1711, n4445);
  and g3585 (n4446, n_234, n_1711);
  and g3586 (n4447, pi0299, n_1696);
  not g3587 (n_1712, n4446);
  not g3588 (n_1713, n4447);
  and g3589 (n4448, n_1712, n_1713);
  and g3590 (n4449, n_841, n4448);
  and g3591 (n4450, n_251, n4448);
  and g3592 (n4451, pi0299, n_1697);
  not g3593 (n_1714, n4451);
  and g3594 (n4452, n_1712, n_1714);
  and g3595 (n4453, n2625, n4452);
  not g3596 (n_1715, n4450);
  not g3597 (n_1716, n4453);
  and g3598 (n4454, n_1715, n_1716);
  not g3599 (n_1717, n4454);
  and g3600 (n4455, n2533, n_1717);
  and g3601 (n4456, n_257, n4448);
  not g3602 (n_1718, n4456);
  and g3603 (n4457, pi0092, n_1718);
  not g3604 (n_1719, n4455);
  and g3605 (n4458, n_1719, n4457);
  and g3606 (n4459, pi0075, n4448);
  and g3607 (n4460, pi0087, n4454);
  and g3608 (n4461, pi0038, n4448);
  not g3609 (n_1720, n4452);
  and g3610 (n4462, pi0039, n_1720);
  and g3611 (n4463, n_234, n_1709);
  and g3612 (n4464, pi0869, n3488);
  not g3613 (n_1721, n4464);
  and g3614 (n4465, n_219, n_1721);
  not g3615 (n_1722, n4465);
  and g3616 (n4466, n4436, n_1722);
  not g3617 (n_1723, n4466);
  and g3618 (n4467, n_1707, n_1723);
  and g3619 (n4468, n4463, n4467);
  and g3620 (n4469, pi0299, n_1684);
  and g3621 (n4470, pi0869, n3499);
  not g3622 (n_1724, n4470);
  and g3623 (n4471, n_1673, n_1724);
  and g3624 (n4472, pi0170, n3508);
  not g3625 (n_1725, n4471);
  not g3626 (n_1726, n4472);
  and g3627 (n4473, n_1725, n_1726);
  not g3628 (n_1727, n4473);
  and g3629 (n4474, pi0869, n_1727);
  and g3630 (n4475, n_879, n4471);
  not g3631 (n_1728, n4474);
  not g3632 (n_1729, n4475);
  and g3633 (n4476, n_1728, n_1729);
  not g3634 (n_1730, n4476);
  and g3635 (n4477, n_188, n_1730);
  and g3636 (n4478, n_937, n4401);
  not g3637 (n_1731, n4478);
  and g3638 (n4479, n_20, n_1731);
  not g3639 (n_1732, n4477);
  and g3640 (n4480, n_1732, n4479);
  not g3641 (n_1733, n4480);
  and g3642 (n4481, n4396, n_1733);
  not g3643 (n_1734, n4481);
  and g3644 (n4482, n_1682, n_1734);
  not g3645 (n_1735, n4482);
  and g3646 (n4483, n_36, n_1735);
  not g3647 (n_1736, n4483);
  and g3648 (n4484, n4469, n_1736);
  and g3649 (n4485, n_936, n4436);
  not g3650 (n_1737, n4485);
  and g3651 (n4486, n4467, n_1737);
  not g3652 (n_1738, n4486);
  and g3653 (n4487, n_223, n_1738);
  not g3654 (n_1739, n4487);
  and g3655 (n4488, n4463, n_1739);
  not g3656 (n_1740, n4488);
  and g3657 (n4489, n_162, n_1740);
  not g3658 (n_1741, n4468);
  and g3659 (n4490, n_1741, n4489);
  not g3660 (n_1742, n4484);
  and g3661 (n4491, n_1742, n4490);
  not g3662 (n_1743, n4462);
  and g3663 (n4492, n_161, n_1743);
  not g3664 (n_1744, n4491);
  and g3665 (n4493, n_1744, n4492);
  not g3666 (n_1745, n4461);
  and g3667 (n4494, n_164, n_1745);
  not g3668 (n_1746, n4493);
  and g3669 (n4495, n_1746, n4494);
  and g3670 (n4496, n_260, n4448);
  and g3671 (n4497, n_1686, n3394);
  and g3672 (n4498, pi0170, n_1567);
  not g3673 (n_1747, n4497);
  and g3674 (n4499, n_188, n_1747);
  not g3675 (n_1748, n4498);
  and g3676 (n4500, n_1748, n4499);
  not g3677 (n_1749, n4500);
  and g3678 (n4501, n4402, n_1749);
  not g3679 (n_1750, n4501);
  and g3680 (n4502, n4396, n_1750);
  not g3681 (n_1751, n4502);
  and g3682 (n4503, n_1682, n_1751);
  not g3683 (n_1752, n4503);
  and g3684 (n4504, n_36, n_1752);
  not g3685 (n_1753, n4504);
  and g3686 (n4505, n_1684, n_1753);
  not g3687 (n_1754, n4505);
  and g3688 (n4506, pi0299, n_1754);
  and g3689 (n4507, n2530, n_1712);
  not g3690 (n_1755, n4506);
  and g3691 (n4508, n_1755, n4507);
  not g3692 (n_1756, n4496);
  and g3693 (n4509, pi0100, n_1756);
  not g3694 (n_1757, n4508);
  and g3695 (n4510, n_1757, n4509);
  not g3696 (n_1758, n4495);
  not g3697 (n_1759, n4510);
  and g3698 (n4511, n_1758, n_1759);
  not g3699 (n_1760, n4511);
  and g3700 (n4512, n_172, n_1760);
  not g3701 (n_1761, n4460);
  and g3702 (n4513, n_171, n_1761);
  not g3703 (n_1762, n4512);
  and g3704 (n4514, n_1762, n4513);
  not g3705 (n_1763, n4459);
  and g3706 (n4515, n_174, n_1763);
  not g3707 (n_1764, n4514);
  and g3708 (n4516, n_1764, n4515);
  not g3709 (n_1765, n4458);
  and g3710 (n4517, n2532, n_1765);
  not g3711 (n_1766, n4516);
  and g3712 (n4518, n_1766, n4517);
  not g3713 (n_1767, n4449);
  and g3714 (n4519, n_176, n_1767);
  not g3715 (n_1768, n4518);
  and g3716 (n4520, n_1768, n4519);
  not g3717 (n_1769, n4433);
  and g3718 (n4521, n_157, n_1769);
  not g3719 (n_1770, n4520);
  and g3720 (n4522, n_1770, n4521);
  not g3721 (n_1771, n4429);
  and g3722 (n4523, n_158, n_1771);
  not g3723 (n_1772, n4522);
  and g3724 (n4524, n_1772, n4523);
  not g3725 (n_1774, pi0248);
  and g3731 (n4528, n_997, n4402);
  and g3732 (n4529, n_1689, n4528);
  not g3733 (n_1777, n4529);
  and g3734 (n4530, n4396, n_1777);
  not g3735 (n_1778, n4530);
  and g3736 (n4531, n_1682, n_1778);
  not g3737 (n_1779, n4531);
  and g3738 (n4532, n_36, n_1779);
  not g3739 (n_1780, n4532);
  and g3740 (n4533, n_1684, n_1780);
  and g3741 (n4534, n3331, n4533);
  and g3742 (n4535, n3556, n_1666);
  not g3743 (n_1781, n4535);
  and g3744 (n4536, n4412, n_1781);
  and g3745 (n4537, n_826, n4536);
  not g3746 (n_1782, n4537);
  and g3747 (n4538, pi0062, n_1782);
  not g3748 (n_1783, n4534);
  and g3749 (n4539, n_1783, n4538);
  not g3750 (n_1784, n4536);
  and g3751 (n4540, n_179, n_1784);
  not g3752 (n_1785, n4533);
  and g3753 (n4541, n2537, n_1785);
  not g3754 (n_1786, n4540);
  and g3755 (n4542, pi0056, n_1786);
  not g3756 (n_1787, n4541);
  and g3757 (n4543, n_1787, n4542);
  and g3758 (n4544, n2572, n4533);
  and g3759 (n4545, n_204, n4536);
  not g3760 (n_1788, n4545);
  and g3761 (n4546, pi0055, n_1788);
  not g3762 (n_1789, n4544);
  and g3763 (n4547, n_1789, n4546);
  and g3764 (n4548, n_921, n_1712);
  and g3765 (n4549, pi0299, n_1784);
  not g3766 (n_1790, n4549);
  and g3767 (n4550, n4548, n_1790);
  and g3768 (n4551, n_841, n4550);
  and g3769 (n4552, n_251, n4550);
  and g3770 (n4553, pi0299, n_1785);
  not g3771 (n_1791, n4553);
  and g3772 (n4554, n4548, n_1791);
  and g3773 (n4555, n2625, n4554);
  not g3774 (n_1792, n4552);
  not g3775 (n_1793, n4555);
  and g3776 (n4556, n_1792, n_1793);
  not g3777 (n_1794, n4556);
  and g3778 (n4557, n2533, n_1794);
  and g3779 (n4558, n_257, n4550);
  not g3780 (n_1795, n4558);
  and g3781 (n4559, pi0092, n_1795);
  not g3782 (n_1796, n4557);
  and g3783 (n4560, n_1796, n4559);
  and g3784 (n4561, pi0075, n4550);
  and g3785 (n4562, pi0087, n4556);
  and g3786 (n4563, pi0038, n4550);
  not g3787 (n_1797, n4554);
  and g3788 (n4564, pi0039, n_1797);
  and g3789 (n4565, n_1686, n3508);
  not g3790 (n_1798, n4565);
  and g3791 (n4566, n_1673, n_1798);
  and g3792 (n4567, n_1686, n_938);
  and g3793 (n4568, pi0869, n_879);
  not g3794 (n_1799, n4567);
  and g3795 (n4569, pi0170, n_1799);
  not g3796 (n_1800, n4568);
  and g3797 (n4570, n_1800, n4569);
  not g3798 (n_1801, n4566);
  not g3799 (n_1802, n4570);
  and g3800 (n4571, n_1801, n_1802);
  not g3801 (n_1803, n4571);
  and g3802 (n4572, n_188, n_1803);
  and g3803 (n4573, n_1181, n4402);
  not g3804 (n_1804, n4572);
  and g3805 (n4574, n_1804, n4573);
  not g3806 (n_1805, n4574);
  and g3807 (n4575, n4396, n_1805);
  not g3808 (n_1806, n4575);
  and g3809 (n4576, n_1682, n_1806);
  not g3810 (n_1807, n4576);
  and g3811 (n4577, n_36, n_1807);
  not g3812 (n_1808, n4577);
  and g3813 (n4578, n4469, n_1808);
  not g3814 (n_1809, n4578);
  and g3815 (n4579, n4489, n_1809);
  not g3816 (n_1810, n4564);
  and g3817 (n4580, n_161, n_1810);
  not g3818 (n_1811, n4579);
  and g3819 (n4581, n_1811, n4580);
  not g3820 (n_1812, n4563);
  and g3821 (n4582, n_164, n_1812);
  not g3822 (n_1813, n4581);
  and g3823 (n4583, n_1813, n4582);
  and g3824 (n4584, n_260, n4550);
  and g3825 (n4585, n_1749, n4528);
  not g3826 (n_1814, n4585);
  and g3827 (n4586, n4396, n_1814);
  not g3828 (n_1815, n4586);
  and g3829 (n4587, n_1682, n_1815);
  not g3830 (n_1816, n4587);
  and g3831 (n4588, n_36, n_1816);
  not g3832 (n_1817, n4588);
  and g3833 (n4589, n_1684, n_1817);
  not g3834 (n_1818, n4589);
  and g3835 (n4590, pi0299, n_1818);
  and g3836 (n4591, n2530, n4548);
  not g3837 (n_1819, n4590);
  and g3838 (n4592, n_1819, n4591);
  not g3839 (n_1820, n4584);
  and g3840 (n4593, pi0100, n_1820);
  not g3841 (n_1821, n4592);
  and g3842 (n4594, n_1821, n4593);
  not g3843 (n_1822, n4583);
  not g3844 (n_1823, n4594);
  and g3845 (n4595, n_1822, n_1823);
  not g3846 (n_1824, n4595);
  and g3847 (n4596, n_172, n_1824);
  not g3848 (n_1825, n4562);
  and g3849 (n4597, n_171, n_1825);
  not g3850 (n_1826, n4596);
  and g3851 (n4598, n_1826, n4597);
  not g3852 (n_1827, n4561);
  and g3853 (n4599, n_174, n_1827);
  not g3854 (n_1828, n4598);
  and g3855 (n4600, n_1828, n4599);
  not g3856 (n_1829, n4560);
  and g3857 (n4601, n2532, n_1829);
  not g3858 (n_1830, n4600);
  and g3859 (n4602, n_1830, n4601);
  not g3860 (n_1831, n4551);
  and g3861 (n4603, n_176, n_1831);
  not g3862 (n_1832, n4602);
  and g3863 (n4604, n_1832, n4603);
  not g3864 (n_1833, n4547);
  and g3865 (n4605, n_157, n_1833);
  not g3866 (n_1834, n4604);
  and g3867 (n4606, n_1834, n4605);
  not g3868 (n_1835, n4543);
  and g3869 (n4607, n_158, n_1835);
  not g3870 (n_1836, n4606);
  and g3871 (n4608, n_1836, n4607);
  and g3877 (n4612, pi0248, n4535);
  not g3878 (n_1839, n4612);
  and g3879 (n4613, n_824, n_1839);
  and g3880 (n4614, n4412, n4613);
  not g3881 (n_1840, n4611);
  not g3882 (n_1841, n4614);
  and g3883 (n4615, n_1840, n_1841);
  not g3884 (n_1842, n4527);
  and g3885 (po0159, n_1842, n4615);
  and g3886 (n4617, pi0215, pi1139);
  not g3887 (n_1844, pi1139);
  and g3888 (n4618, pi0216, n_1844);
  and g3889 (n4619, pi0833, pi0920);
  and g3890 (n4620, n_486, pi1139);
  not g3891 (n_1846, n4619);
  and g3892 (n4621, n_20, n_1846);
  not g3893 (n_1847, n4620);
  and g3894 (n4622, n_1847, n4621);
  not g3895 (n_1848, n4622);
  and g3896 (n4623, pi0221, n_1848);
  not g3897 (n_1849, n4618);
  and g3898 (n4624, n_1849, n4623);
  and g3899 (n4625, pi0216, pi0281);
  not g3900 (n_1851, n4625);
  and g3901 (n4626, n_26, n_1851);
  not g3902 (n_1853, pi0862);
  and g3903 (n4627, n_20, n_1853);
  and g3904 (n4628, n3630, n4627);
  not g3905 (n_1854, n4628);
  and g3906 (n4629, n4626, n_1854);
  not g3907 (n_1855, n4624);
  not g3908 (n_1856, n4629);
  and g3909 (n4630, n_1855, n_1856);
  not g3910 (n_1857, n4623);
  and g3911 (n4631, n_20, n_1857);
  and g3912 (n4632, pi0148, n_19);
  and g3913 (n4633, n4631, n4632);
  not g3914 (n_1859, n4633);
  and g3915 (n4634, n_36, n_1859);
  not g3916 (n_1860, n4630);
  and g3917 (n4635, n_1860, n4634);
  not g3918 (n_1861, n4617);
  not g3919 (n_1862, n4635);
  and g3920 (n4636, n_1861, n_1862);
  not g3921 (n_1863, n4636);
  and g3922 (n4637, n_909, n_1863);
  not g3923 (n_1864, n4637);
  and g3924 (n4638, n_824, n_1864);
  and g3925 (n4639, n_826, n_1864);
  not g3926 (n_1865, pi0148);
  and g3927 (n4640, n_1865, n_36);
  and g3928 (n4641, pi0862, n_997);
  and g3929 (n4642, n_19, n_1324);
  not g3930 (n_1866, n4641);
  and g3931 (n4643, n_20, n_1866);
  not g3932 (n_1867, n4642);
  and g3933 (n4644, n_1867, n4643);
  not g3934 (n_1868, n4644);
  and g3935 (n4645, n4626, n_1868);
  not g3936 (n_1869, n4645);
  and g3937 (n4646, n_1855, n_1869);
  not g3938 (n_1870, n4646);
  and g3939 (n4647, n4640, n_1870);
  and g3940 (n4648, pi0148, n_36);
  and g3941 (n4649, n_1324, n_1047);
  not g3942 (n_1871, n4649);
  and g3943 (n4650, n4627, n_1871);
  not g3944 (n_1872, n4650);
  and g3945 (n4651, n4626, n_1872);
  not g3946 (n_1873, n4651);
  and g3947 (n4652, n_1855, n_1873);
  and g3948 (n4653, n4631, n4649);
  not g3949 (n_1874, n4653);
  and g3950 (n4654, n4648, n_1874);
  not g3951 (n_1875, n4652);
  and g3952 (n4655, n_1875, n4654);
  not g3953 (n_1876, n4655);
  and g3954 (n4656, n_1861, n_1876);
  not g3955 (n_1877, n4647);
  and g3956 (n4657, n_1877, n4656);
  and g3957 (n4658, n3331, n4657);
  not g3958 (n_1878, n4639);
  and g3959 (n4659, pi0062, n_1878);
  not g3960 (n_1879, n4658);
  and g3961 (n4660, n_1879, n4659);
  not g3962 (n_1880, n4657);
  and g3963 (n4661, n2537, n_1880);
  and g3964 (n4662, n_179, n4637);
  not g3965 (n_1881, n4662);
  and g3966 (n4663, pi0056, n_1881);
  not g3967 (n_1882, n4661);
  and g3968 (n4664, n_1882, n4663);
  and g3969 (n4665, n_204, n_1864);
  and g3970 (n4666, n2572, n4657);
  not g3971 (n_1883, n4665);
  and g3972 (n4667, pi0055, n_1883);
  not g3973 (n_1884, n4666);
  and g3974 (n4668, n_1884, n4667);
  and g3975 (n4669, pi0223, pi1139);
  and g3976 (n4670, n_1844, n_221);
  not g3977 (n_1885, pi0920);
  and g3978 (n4671, n_1885, n2591);
  not g3979 (n_1886, n4670);
  and g3980 (n4672, pi0222, n_1886);
  not g3981 (n_1887, n4671);
  and g3982 (n4673, n_1887, n4672);
  not g3983 (n_1888, n4669);
  and g3984 (n4674, n_219, n_1888);
  not g3985 (n_1889, n4673);
  and g3986 (n4675, n_1889, n4674);
  and g3987 (n4676, n2442, n4675);
  and g3988 (n4677, n_1853, n4675);
  and g3989 (n4678, pi0224, pi0281);
  not g3990 (n_1890, n4678);
  and g3991 (n4679, n_226, n_1890);
  not g3992 (n_1891, n4679);
  and g3993 (n4680, n_1889, n_1891);
  not g3994 (n_1892, n4680);
  and g3995 (n4681, n_223, n_1892);
  not g3996 (n_1893, n4681);
  and g3997 (n4682, n_1888, n_1893);
  not g3998 (n_1894, n4682);
  and g3999 (n4683, n_234, n_1894);
  not g4000 (n_1895, n4677);
  and g4001 (n4684, n_1895, n4683);
  not g4002 (n_1896, n4676);
  and g4003 (n4685, n_1896, n4684);
  and g4004 (n4686, pi0299, n4637);
  not g4005 (n_1897, n4685);
  not g4006 (n_1898, n4686);
  and g4007 (n4687, n_1897, n_1898);
  and g4008 (n4688, n_841, n4687);
  and g4009 (n4689, n_251, n4687);
  and g4010 (n4690, pi0299, n_1880);
  not g4011 (n_1899, n4690);
  and g4012 (n4691, n_1897, n_1899);
  and g4013 (n4692, n2625, n4691);
  not g4014 (n_1900, n4689);
  not g4015 (n_1901, n4692);
  and g4016 (n4693, n_1900, n_1901);
  not g4017 (n_1902, n4693);
  and g4018 (n4694, n2533, n_1902);
  and g4019 (n4695, n_257, n4687);
  not g4020 (n_1903, n4695);
  and g4021 (n4696, pi0092, n_1903);
  not g4022 (n_1904, n4694);
  and g4023 (n4697, n_1904, n4696);
  and g4024 (n4698, pi0075, n4687);
  and g4025 (n4699, pi0087, n4693);
  and g4026 (n4700, n_260, n4687);
  and g4027 (n4701, n_19, n_1046);
  and g4028 (n4702, n4626, n4701);
  not g4029 (n_1905, n4702);
  and g4030 (n4703, n4646, n_1905);
  not g4031 (n_1906, n4703);
  and g4032 (n4704, n4640, n_1906);
  and g4033 (n4705, n3631, n4626);
  not g4034 (n_1907, n4705);
  and g4035 (n4706, n4652, n_1907);
  and g4036 (n4707, n3631, n4631);
  not g4037 (n_1908, n4707);
  and g4038 (n4708, n4648, n_1908);
  not g4039 (n_1909, n4706);
  and g4040 (n4709, n_1909, n4708);
  not g4041 (n_1910, n4704);
  and g4042 (n4710, n_1861, n_1910);
  not g4043 (n_1911, n4709);
  and g4044 (n4711, n_1911, n4710);
  not g4045 (n_1912, n4711);
  and g4046 (n4712, pi0299, n_1912);
  and g4047 (n4713, n2530, n_1897);
  not g4048 (n_1913, n4712);
  and g4049 (n4714, n_1913, n4713);
  not g4050 (n_1914, n4700);
  and g4051 (n4715, pi0100, n_1914);
  not g4052 (n_1915, n4714);
  and g4053 (n4716, n_1915, n4715);
  and g4054 (n4717, pi0038, n4687);
  not g4055 (n_1916, n4691);
  and g4056 (n4718, pi0039, n_1916);
  and g4057 (n4719, n_936, n4675);
  and g4058 (n4720, n_1895, n_1894);
  not g4059 (n_1917, n4719);
  and g4060 (n4721, n_1917, n4720);
  not g4061 (n_1918, n4721);
  and g4062 (n4722, n_234, n_1918);
  and g4063 (n4723, n_949, n4627);
  not g4064 (n_1919, n4723);
  and g4065 (n4724, n4626, n_1919);
  not g4066 (n_1920, n4724);
  and g4067 (n4725, n_1855, n_1920);
  and g4068 (n4726, n3511, n4631);
  not g4069 (n_1921, n4726);
  and g4070 (n4727, n4648, n_1921);
  not g4071 (n_1922, n4725);
  and g4072 (n4728, n_1922, n4727);
  and g4073 (n4729, pi0862, n_941);
  and g4074 (n4730, n_188, n3416);
  not g4075 (n_1923, n4730);
  and g4076 (n4731, n_19, n_1923);
  and g4077 (n4732, n_1853, n4731);
  not g4078 (n_1924, n4729);
  and g4079 (n4733, n_20, n_1924);
  not g4080 (n_1925, n4732);
  and g4081 (n4734, n_1925, n4733);
  not g4082 (n_1926, n4734);
  and g4083 (n4735, n4626, n_1926);
  not g4084 (n_1927, n4735);
  and g4085 (n4736, n_1855, n_1927);
  not g4086 (n_1928, n4736);
  and g4087 (n4737, n4640, n_1928);
  not g4093 (n_1931, n4722);
  and g4094 (n4741, n_162, n_1931);
  not g4095 (n_1932, n4740);
  and g4096 (n4742, n_1932, n4741);
  not g4097 (n_1933, n4718);
  and g4098 (n4743, n_161, n_1933);
  not g4099 (n_1934, n4742);
  and g4100 (n4744, n_1934, n4743);
  not g4101 (n_1935, n4717);
  and g4102 (n4745, n_164, n_1935);
  not g4103 (n_1936, n4744);
  and g4104 (n4746, n_1936, n4745);
  not g4105 (n_1937, n4716);
  not g4106 (n_1938, n4746);
  and g4107 (n4747, n_1937, n_1938);
  not g4108 (n_1939, n4747);
  and g4109 (n4748, n_172, n_1939);
  not g4110 (n_1940, n4699);
  and g4111 (n4749, n_171, n_1940);
  not g4112 (n_1941, n4748);
  and g4113 (n4750, n_1941, n4749);
  not g4114 (n_1942, n4698);
  and g4115 (n4751, n_174, n_1942);
  not g4116 (n_1943, n4750);
  and g4117 (n4752, n_1943, n4751);
  not g4118 (n_1944, n4697);
  and g4119 (n4753, n2532, n_1944);
  not g4120 (n_1945, n4752);
  and g4121 (n4754, n_1945, n4753);
  not g4122 (n_1946, n4688);
  and g4123 (n4755, n_176, n_1946);
  not g4124 (n_1947, n4754);
  and g4125 (n4756, n_1947, n4755);
  not g4126 (n_1948, n4668);
  and g4127 (n4757, n_157, n_1948);
  not g4128 (n_1949, n4756);
  and g4129 (n4758, n_1949, n4757);
  not g4130 (n_1950, n4664);
  and g4131 (n4759, n_158, n_1950);
  not g4132 (n_1951, n4758);
  and g4133 (n4760, n_1951, n4759);
  not g4134 (n_1952, n4660);
  and g4135 (n4761, n3328, n_1952);
  not g4136 (n_1953, n4760);
  and g4137 (n4762, n_1953, n4761);
  not g4138 (n_1955, pi0247);
  not g4139 (n_1956, n4638);
  and g4140 (n4763, n_1955, n_1956);
  not g4141 (n_1957, n4762);
  and g4142 (n4764, n_1957, n4763);
  and g4143 (n4765, n_824, n4636);
  and g4144 (n4766, n_826, n4636);
  and g4145 (n4767, n4634, n_1875);
  not g4146 (n_1958, n4767);
  and g4147 (n4768, n4656, n_1958);
  and g4148 (n4769, n3331, n4768);
  not g4149 (n_1959, n4766);
  and g4150 (n4770, pi0062, n_1959);
  not g4151 (n_1960, n4769);
  and g4152 (n4771, n_1960, n4770);
  and g4153 (n4772, n_179, n_1863);
  not g4154 (n_1961, n4768);
  and g4155 (n4773, n2537, n_1961);
  not g4156 (n_1962, n4772);
  and g4157 (n4774, pi0056, n_1962);
  not g4158 (n_1963, n4773);
  and g4159 (n4775, n_1963, n4774);
  and g4160 (n4776, n_204, n4636);
  and g4161 (n4777, n2572, n4768);
  not g4162 (n_1964, n4776);
  and g4163 (n4778, pi0055, n_1964);
  not g4164 (n_1965, n4777);
  and g4165 (n4779, n_1965, n4778);
  not g4166 (n_1966, n4684);
  and g4167 (n4780, n_921, n_1966);
  and g4168 (n4781, pi0299, n_1863);
  not g4169 (n_1967, n4781);
  and g4170 (n4782, n4780, n_1967);
  and g4171 (n4783, n_841, n4782);
  and g4172 (n4784, n_251, n4782);
  and g4173 (n4785, pi0299, n_1961);
  not g4174 (n_1968, n4785);
  and g4175 (n4786, n4780, n_1968);
  and g4176 (n4787, n2625, n4786);
  not g4177 (n_1969, n4784);
  not g4178 (n_1970, n4787);
  and g4179 (n4788, n_1969, n_1970);
  not g4180 (n_1971, n4788);
  and g4181 (n4789, n2533, n_1971);
  and g4182 (n4790, n_257, n4782);
  not g4183 (n_1972, n4790);
  and g4184 (n4791, pi0092, n_1972);
  not g4185 (n_1973, n4789);
  and g4186 (n4792, n_1973, n4791);
  and g4187 (n4793, pi0075, n4782);
  and g4188 (n4794, pi0087, n4788);
  and g4189 (n4795, n_260, n4782);
  and g4190 (n4796, n4640, n_1909);
  and g4191 (n4797, n_20, n_1855);
  and g4192 (n4798, n4701, n4797);
  and g4193 (n4799, n4648, n_1875);
  not g4194 (n_1974, n4798);
  and g4195 (n4800, n_1974, n4799);
  not g4196 (n_1975, n4800);
  and g4197 (n4801, n_1861, n_1975);
  not g4198 (n_1976, n4796);
  and g4199 (n4802, n_1976, n4801);
  not g4200 (n_1977, n4802);
  and g4201 (n4803, pi0299, n_1977);
  and g4202 (n4804, n2530, n4780);
  not g4203 (n_1978, n4803);
  and g4204 (n4805, n_1978, n4804);
  not g4205 (n_1979, n4795);
  and g4206 (n4806, pi0100, n_1979);
  not g4207 (n_1980, n4805);
  and g4208 (n4807, n_1980, n4806);
  and g4209 (n4808, pi0038, n4782);
  not g4210 (n_1981, n4786);
  and g4211 (n4809, pi0039, n_1981);
  and g4212 (n4810, n3488, n4677);
  not g4213 (n_1982, n4810);
  and g4214 (n4811, n4683, n_1982);
  not g4215 (n_1983, n4731);
  and g4216 (n4812, pi0862, n_1983);
  and g4217 (n4813, n_1853, n3501);
  not g4218 (n_1984, n4813);
  and g4219 (n4814, n_20, n_1984);
  not g4220 (n_1985, n4812);
  and g4221 (n4815, n_1985, n4814);
  not g4222 (n_1986, n4815);
  and g4223 (n4816, n4626, n_1986);
  not g4224 (n_1987, n4816);
  and g4225 (n4817, n_1855, n_1987);
  not g4226 (n_1988, n4817);
  and g4227 (n4818, n4648, n_1988);
  and g4228 (n4819, n4640, n_1922);
  not g4229 (n_1989, n4819);
  and g4230 (n4820, n_1861, n_1989);
  not g4231 (n_1990, n4818);
  and g4232 (n4821, n_1990, n4820);
  not g4233 (n_1991, n4821);
  and g4234 (n4822, pi0299, n_1991);
  not g4235 (n_1992, n4811);
  not g4236 (n_1993, n4822);
  and g4237 (n4823, n_1992, n_1993);
  not g4238 (n_1994, n4823);
  and g4239 (n4824, n_162, n_1994);
  not g4240 (n_1995, n4809);
  and g4241 (n4825, n_161, n_1995);
  not g4242 (n_1996, n4824);
  and g4243 (n4826, n_1996, n4825);
  not g4244 (n_1997, n4808);
  and g4245 (n4827, n_164, n_1997);
  not g4246 (n_1998, n4826);
  and g4247 (n4828, n_1998, n4827);
  not g4248 (n_1999, n4807);
  not g4249 (n_2000, n4828);
  and g4250 (n4829, n_1999, n_2000);
  not g4251 (n_2001, n4829);
  and g4252 (n4830, n_172, n_2001);
  not g4253 (n_2002, n4794);
  and g4254 (n4831, n_171, n_2002);
  not g4255 (n_2003, n4830);
  and g4256 (n4832, n_2003, n4831);
  not g4257 (n_2004, n4793);
  and g4258 (n4833, n_174, n_2004);
  not g4259 (n_2005, n4832);
  and g4260 (n4834, n_2005, n4833);
  not g4261 (n_2006, n4792);
  and g4262 (n4835, n2532, n_2006);
  not g4263 (n_2007, n4834);
  and g4264 (n4836, n_2007, n4835);
  not g4265 (n_2008, n4783);
  and g4266 (n4837, n_176, n_2008);
  not g4267 (n_2009, n4836);
  and g4268 (n4838, n_2009, n4837);
  not g4269 (n_2010, n4779);
  and g4270 (n4839, n_157, n_2010);
  not g4271 (n_2011, n4838);
  and g4272 (n4840, n_2011, n4839);
  not g4273 (n_2012, n4775);
  and g4274 (n4841, n_158, n_2012);
  not g4275 (n_2013, n4840);
  and g4276 (n4842, n_2013, n4841);
  not g4277 (n_2014, n4771);
  and g4278 (n4843, n3328, n_2014);
  not g4279 (n_2015, n4842);
  and g4280 (n4844, n_2015, n4843);
  not g4281 (n_2016, n4765);
  and g4282 (n4845, pi0247, n_2016);
  not g4283 (n_2017, n4844);
  and g4284 (n4846, n_2017, n4845);
  or g4285 (po0160, n4764, n4846);
  and g4286 (n4848, pi0215, pi1138);
  and g4287 (n4849, pi0216, pi0269);
  not g4288 (n_2020, n4849);
  and g4289 (n4850, n_26, n_2020);
  and g4290 (n4851, n_180, pi0169);
  and g4291 (n4852, pi0877, n_145);
  not g4292 (n_2023, n4852);
  and g4293 (n4853, pi0105, n_2023);
  not g4294 (n_2024, n4851);
  and g4295 (n4854, pi0228, n_2024);
  not g4296 (n_2025, n4853);
  and g4297 (n4855, n_2025, n4854);
  not g4298 (n_2026, n4855);
  and g4299 (n4856, n_20, n_2026);
  not g4300 (n_2027, pi0169);
  and g4301 (n4857, n_2027, n_188);
  not g4302 (n_2028, n4857);
  and g4303 (n4858, n4856, n_2028);
  not g4304 (n_2029, n4858);
  and g4305 (n4859, n4850, n_2029);
  not g4306 (n_2030, pi1138);
  and g4307 (n4860, n_2030, n_29);
  not g4308 (n_2032, pi0940);
  and g4309 (n4861, n_2032, n2452);
  not g4310 (n_2033, n4860);
  and g4311 (n4862, pi0221, n_2033);
  not g4312 (n_2034, n4861);
  and g4313 (n4863, n_2034, n4862);
  not g4314 (n_2035, n4859);
  not g4315 (n_2036, n4863);
  and g4316 (n4864, n_2035, n_2036);
  not g4317 (n_2037, n4864);
  and g4318 (n4865, n_36, n_2037);
  not g4319 (n_2038, n4848);
  not g4320 (n_2039, n4865);
  and g4321 (n4866, n_2038, n_2039);
  and g4322 (n4867, n_826, n4866);
  not g4323 (n_2040, pi0877);
  and g4324 (n4868, n_2040, n2521);
  and g4325 (n4869, pi0169, n_207);
  not g4326 (n_2041, n4868);
  and g4327 (n4870, n_188, n_2041);
  not g4328 (n_2042, n4869);
  and g4329 (n4871, n_2042, n4870);
  not g4330 (n_2043, n4871);
  and g4331 (n4872, n4856, n_2043);
  not g4332 (n_2044, n4872);
  and g4333 (n4873, n4850, n_2044);
  not g4334 (n_2045, n4873);
  and g4335 (n4874, n_2036, n_2045);
  not g4336 (n_2046, n4874);
  and g4337 (n4875, n_36, n_2046);
  not g4338 (n_2047, n4875);
  and g4339 (n4876, n_2038, n_2047);
  and g4340 (n4877, n3331, n4876);
  not g4341 (n_2048, n4867);
  and g4342 (n4878, pi0062, n_2048);
  not g4343 (n_2049, n4877);
  and g4344 (n4879, n_2049, n4878);
  not g4345 (n_2050, n4866);
  and g4346 (n4880, n_179, n_2050);
  not g4347 (n_2051, n4876);
  and g4348 (n4881, n2537, n_2051);
  not g4349 (n_2052, n4880);
  and g4350 (n4882, pi0056, n_2052);
  not g4351 (n_2053, n4881);
  and g4352 (n4883, n_2053, n4882);
  and g4353 (n4884, n_204, n4866);
  and g4354 (n4885, n2572, n4876);
  not g4355 (n_2054, n4884);
  and g4356 (n4886, pi0055, n_2054);
  not g4357 (n_2055, n4885);
  and g4358 (n4887, n_2055, n4886);
  and g4359 (n4888, pi0223, pi1138);
  and g4360 (n4889, pi0224, pi0269);
  not g4361 (n_2056, n4889);
  and g4362 (n4890, n_226, n_2056);
  and g4363 (n4891, n_219, n_2023);
  not g4364 (n_2057, n4891);
  and g4365 (n4892, n4890, n_2057);
  and g4366 (n4893, n_2030, n_221);
  and g4367 (n4894, n_2032, n2591);
  not g4368 (n_2058, n4893);
  and g4369 (n4895, pi0222, n_2058);
  not g4370 (n_2059, n4894);
  and g4371 (n4896, n_2059, n4895);
  not g4372 (n_2060, n4892);
  not g4373 (n_2061, n4896);
  and g4374 (n4897, n_2060, n_2061);
  not g4375 (n_2062, n4897);
  and g4376 (n4898, n_223, n_2062);
  not g4377 (n_2063, n4888);
  not g4378 (n_2064, n4898);
  and g4379 (n4899, n_2063, n_2064);
  not g4380 (n_2065, n4899);
  and g4381 (n4900, n_234, n_2065);
  and g4382 (n4901, pi0299, n_2050);
  not g4383 (n_2066, n4900);
  not g4384 (n_2067, n4901);
  and g4385 (n4902, n_2066, n_2067);
  and g4386 (n4903, n_841, n4902);
  and g4387 (n4904, n_251, n4902);
  and g4388 (n4905, pi0299, n_2051);
  not g4389 (n_2068, n4905);
  and g4390 (n4906, n_2066, n_2068);
  and g4391 (n4907, n2625, n4906);
  not g4392 (n_2069, n4904);
  not g4393 (n_2070, n4907);
  and g4394 (n4908, n_2069, n_2070);
  not g4395 (n_2071, n4908);
  and g4396 (n4909, n2533, n_2071);
  and g4397 (n4910, n_257, n4902);
  not g4398 (n_2072, n4910);
  and g4399 (n4911, pi0092, n_2072);
  not g4400 (n_2073, n4909);
  and g4401 (n4912, n_2073, n4911);
  and g4402 (n4913, pi0075, n4902);
  and g4403 (n4914, pi0087, n4908);
  and g4404 (n4915, pi0038, n4902);
  not g4405 (n_2074, n4906);
  and g4406 (n4916, pi0039, n_2074);
  and g4407 (n4917, n_234, n_2063);
  and g4408 (n4918, pi0877, n3488);
  not g4409 (n_2075, n4918);
  and g4410 (n4919, n_219, n_2075);
  not g4411 (n_2076, n4919);
  and g4412 (n4920, n4890, n_2076);
  not g4413 (n_2077, n4920);
  and g4414 (n4921, n_2061, n_2077);
  and g4415 (n4922, n4917, n4921);
  and g4416 (n4923, pi0299, n_2038);
  and g4417 (n4924, pi0877, n3499);
  not g4418 (n_2078, n4924);
  and g4419 (n4925, n_2027, n_2078);
  and g4420 (n4926, pi0169, n3508);
  not g4421 (n_2079, n4925);
  not g4422 (n_2080, n4926);
  and g4423 (n4927, n_2079, n_2080);
  not g4424 (n_2081, n4927);
  and g4425 (n4928, pi0877, n_2081);
  and g4426 (n4929, n_879, n4925);
  not g4427 (n_2082, n4928);
  not g4428 (n_2083, n4929);
  and g4429 (n4930, n_2082, n_2083);
  not g4430 (n_2084, n4930);
  and g4431 (n4931, n_188, n_2084);
  and g4432 (n4932, n_937, n4855);
  not g4433 (n_2085, n4932);
  and g4434 (n4933, n_20, n_2085);
  not g4435 (n_2086, n4931);
  and g4436 (n4934, n_2086, n4933);
  not g4437 (n_2087, n4934);
  and g4438 (n4935, n4850, n_2087);
  not g4439 (n_2088, n4935);
  and g4440 (n4936, n_2036, n_2088);
  not g4441 (n_2089, n4936);
  and g4442 (n4937, n_36, n_2089);
  not g4443 (n_2090, n4937);
  and g4444 (n4938, n4923, n_2090);
  and g4445 (n4939, n_936, n4890);
  not g4446 (n_2091, n4939);
  and g4447 (n4940, n4921, n_2091);
  not g4448 (n_2092, n4940);
  and g4449 (n4941, n_223, n_2092);
  not g4450 (n_2093, n4941);
  and g4451 (n4942, n4917, n_2093);
  not g4452 (n_2094, n4942);
  and g4453 (n4943, n_162, n_2094);
  not g4454 (n_2095, n4922);
  and g4455 (n4944, n_2095, n4943);
  not g4456 (n_2096, n4938);
  and g4457 (n4945, n_2096, n4944);
  not g4458 (n_2097, n4916);
  and g4459 (n4946, n_161, n_2097);
  not g4460 (n_2098, n4945);
  and g4461 (n4947, n_2098, n4946);
  not g4462 (n_2099, n4915);
  and g4463 (n4948, n_164, n_2099);
  not g4464 (n_2100, n4947);
  and g4465 (n4949, n_2100, n4948);
  and g4466 (n4950, n_260, n4902);
  and g4467 (n4951, n_2040, n3394);
  and g4468 (n4952, pi0169, n_1567);
  not g4469 (n_2101, n4951);
  and g4470 (n4953, n_188, n_2101);
  not g4471 (n_2102, n4952);
  and g4472 (n4954, n_2102, n4953);
  not g4473 (n_2103, n4954);
  and g4474 (n4955, n4856, n_2103);
  not g4475 (n_2104, n4955);
  and g4476 (n4956, n4850, n_2104);
  not g4477 (n_2105, n4956);
  and g4478 (n4957, n_2036, n_2105);
  not g4479 (n_2106, n4957);
  and g4480 (n4958, n_36, n_2106);
  not g4481 (n_2107, n4958);
  and g4482 (n4959, n_2038, n_2107);
  not g4483 (n_2108, n4959);
  and g4484 (n4960, pi0299, n_2108);
  and g4485 (n4961, n2530, n_2066);
  not g4486 (n_2109, n4960);
  and g4487 (n4962, n_2109, n4961);
  not g4488 (n_2110, n4950);
  and g4489 (n4963, pi0100, n_2110);
  not g4490 (n_2111, n4962);
  and g4491 (n4964, n_2111, n4963);
  not g4492 (n_2112, n4949);
  not g4493 (n_2113, n4964);
  and g4494 (n4965, n_2112, n_2113);
  not g4495 (n_2114, n4965);
  and g4496 (n4966, n_172, n_2114);
  not g4497 (n_2115, n4914);
  and g4498 (n4967, n_171, n_2115);
  not g4499 (n_2116, n4966);
  and g4500 (n4968, n_2116, n4967);
  not g4501 (n_2117, n4913);
  and g4502 (n4969, n_174, n_2117);
  not g4503 (n_2118, n4968);
  and g4504 (n4970, n_2118, n4969);
  not g4505 (n_2119, n4912);
  and g4506 (n4971, n2532, n_2119);
  not g4507 (n_2120, n4970);
  and g4508 (n4972, n_2120, n4971);
  not g4509 (n_2121, n4903);
  and g4510 (n4973, n_176, n_2121);
  not g4511 (n_2122, n4972);
  and g4512 (n4974, n_2122, n4973);
  not g4513 (n_2123, n4887);
  and g4514 (n4975, n_157, n_2123);
  not g4515 (n_2124, n4974);
  and g4516 (n4976, n_2124, n4975);
  not g4517 (n_2125, n4883);
  and g4518 (n4977, n_158, n_2125);
  not g4519 (n_2126, n4976);
  and g4520 (n4978, n_2126, n4977);
  not g4521 (n_2128, pi0246);
  and g4527 (n4982, n_997, n4856);
  and g4528 (n4983, n_2043, n4982);
  not g4529 (n_2131, n4983);
  and g4530 (n4984, n4850, n_2131);
  not g4531 (n_2132, n4984);
  and g4532 (n4985, n_2036, n_2132);
  not g4533 (n_2133, n4985);
  and g4534 (n4986, n_36, n_2133);
  not g4535 (n_2134, n4986);
  and g4536 (n4987, n_2038, n_2134);
  and g4537 (n4988, n3331, n4987);
  and g4538 (n4989, n3556, n_2020);
  not g4539 (n_2135, n4989);
  and g4540 (n4990, n4866, n_2135);
  and g4541 (n4991, n_826, n4990);
  not g4542 (n_2136, n4991);
  and g4543 (n4992, pi0062, n_2136);
  not g4544 (n_2137, n4988);
  and g4545 (n4993, n_2137, n4992);
  not g4546 (n_2138, n4990);
  and g4547 (n4994, n_179, n_2138);
  not g4548 (n_2139, n4987);
  and g4549 (n4995, n2537, n_2139);
  not g4550 (n_2140, n4994);
  and g4551 (n4996, pi0056, n_2140);
  not g4552 (n_2141, n4995);
  and g4553 (n4997, n_2141, n4996);
  and g4554 (n4998, n2572, n4987);
  and g4555 (n4999, n_204, n4990);
  not g4556 (n_2142, n4999);
  and g4557 (n5000, pi0055, n_2142);
  not g4558 (n_2143, n4998);
  and g4559 (n5001, n_2143, n5000);
  and g4560 (n5002, n_921, n_2066);
  and g4561 (n5003, pi0299, n_2138);
  not g4562 (n_2144, n5003);
  and g4563 (n5004, n5002, n_2144);
  and g4564 (n5005, n_841, n5004);
  and g4565 (n5006, n_251, n5004);
  and g4566 (n5007, pi0299, n_2139);
  not g4567 (n_2145, n5007);
  and g4568 (n5008, n5002, n_2145);
  and g4569 (n5009, n2625, n5008);
  not g4570 (n_2146, n5006);
  not g4571 (n_2147, n5009);
  and g4572 (n5010, n_2146, n_2147);
  not g4573 (n_2148, n5010);
  and g4574 (n5011, n2533, n_2148);
  and g4575 (n5012, n_257, n5004);
  not g4576 (n_2149, n5012);
  and g4577 (n5013, pi0092, n_2149);
  not g4578 (n_2150, n5011);
  and g4579 (n5014, n_2150, n5013);
  and g4580 (n5015, pi0075, n5004);
  and g4581 (n5016, pi0087, n5010);
  and g4582 (n5017, pi0038, n5004);
  not g4583 (n_2151, n5008);
  and g4584 (n5018, pi0039, n_2151);
  and g4585 (n5019, n_2040, n3508);
  not g4586 (n_2152, n5019);
  and g4587 (n5020, n_2027, n_2152);
  and g4588 (n5021, n_2040, n_938);
  and g4589 (n5022, pi0877, n_879);
  not g4590 (n_2153, n5021);
  and g4591 (n5023, pi0169, n_2153);
  not g4592 (n_2154, n5022);
  and g4593 (n5024, n_2154, n5023);
  not g4594 (n_2155, n5020);
  not g4595 (n_2156, n5024);
  and g4596 (n5025, n_2155, n_2156);
  not g4597 (n_2157, n5025);
  and g4598 (n5026, n_188, n_2157);
  and g4599 (n5027, n_1181, n4856);
  not g4600 (n_2158, n5026);
  and g4601 (n5028, n_2158, n5027);
  not g4602 (n_2159, n5028);
  and g4603 (n5029, n4850, n_2159);
  not g4604 (n_2160, n5029);
  and g4605 (n5030, n_2036, n_2160);
  not g4606 (n_2161, n5030);
  and g4607 (n5031, n_36, n_2161);
  not g4608 (n_2162, n5031);
  and g4609 (n5032, n4923, n_2162);
  not g4610 (n_2163, n5032);
  and g4611 (n5033, n4943, n_2163);
  not g4612 (n_2164, n5018);
  and g4613 (n5034, n_161, n_2164);
  not g4614 (n_2165, n5033);
  and g4615 (n5035, n_2165, n5034);
  not g4616 (n_2166, n5017);
  and g4617 (n5036, n_164, n_2166);
  not g4618 (n_2167, n5035);
  and g4619 (n5037, n_2167, n5036);
  and g4620 (n5038, n_260, n5004);
  and g4621 (n5039, n_2103, n4982);
  not g4622 (n_2168, n5039);
  and g4623 (n5040, n4850, n_2168);
  not g4624 (n_2169, n5040);
  and g4625 (n5041, n_2036, n_2169);
  not g4626 (n_2170, n5041);
  and g4627 (n5042, n_36, n_2170);
  not g4628 (n_2171, n5042);
  and g4629 (n5043, n_2038, n_2171);
  not g4630 (n_2172, n5043);
  and g4631 (n5044, pi0299, n_2172);
  and g4632 (n5045, n2530, n5002);
  not g4633 (n_2173, n5044);
  and g4634 (n5046, n_2173, n5045);
  not g4635 (n_2174, n5038);
  and g4636 (n5047, pi0100, n_2174);
  not g4637 (n_2175, n5046);
  and g4638 (n5048, n_2175, n5047);
  not g4639 (n_2176, n5037);
  not g4640 (n_2177, n5048);
  and g4641 (n5049, n_2176, n_2177);
  not g4642 (n_2178, n5049);
  and g4643 (n5050, n_172, n_2178);
  not g4644 (n_2179, n5016);
  and g4645 (n5051, n_171, n_2179);
  not g4646 (n_2180, n5050);
  and g4647 (n5052, n_2180, n5051);
  not g4648 (n_2181, n5015);
  and g4649 (n5053, n_174, n_2181);
  not g4650 (n_2182, n5052);
  and g4651 (n5054, n_2182, n5053);
  not g4652 (n_2183, n5014);
  and g4653 (n5055, n2532, n_2183);
  not g4654 (n_2184, n5054);
  and g4655 (n5056, n_2184, n5055);
  not g4656 (n_2185, n5005);
  and g4657 (n5057, n_176, n_2185);
  not g4658 (n_2186, n5056);
  and g4659 (n5058, n_2186, n5057);
  not g4660 (n_2187, n5001);
  and g4661 (n5059, n_157, n_2187);
  not g4662 (n_2188, n5058);
  and g4663 (n5060, n_2188, n5059);
  not g4664 (n_2189, n4997);
  and g4665 (n5061, n_158, n_2189);
  not g4666 (n_2190, n5060);
  and g4667 (n5062, n_2190, n5061);
  and g4673 (n5066, pi0246, n4989);
  not g4674 (n_2193, n5066);
  and g4675 (n5067, n_824, n_2193);
  and g4676 (n5068, n4866, n5067);
  not g4677 (n_2194, n5065);
  not g4678 (n_2195, n5068);
  and g4679 (n5069, n_2194, n_2195);
  not g4680 (n_2196, n4981);
  and g4681 (po0161, n_2196, n5069);
  and g4682 (n5071, pi0215, pi1137);
  and g4683 (n5072, pi0216, pi0280);
  not g4684 (n_2199, n5072);
  and g4685 (n5073, n_26, n_2199);
  and g4686 (n5074, n_180, pi0168);
  and g4687 (n5075, pi0878, n_145);
  not g4688 (n_2202, n5075);
  and g4689 (n5076, pi0105, n_2202);
  not g4690 (n_2203, n5074);
  and g4691 (n5077, pi0228, n_2203);
  not g4692 (n_2204, n5076);
  and g4693 (n5078, n_2204, n5077);
  not g4694 (n_2205, n5078);
  and g4695 (n5079, n_20, n_2205);
  not g4696 (n_2206, pi0168);
  and g4697 (n5080, n_2206, n_188);
  not g4698 (n_2207, n5080);
  and g4699 (n5081, n5079, n_2207);
  not g4700 (n_2208, n5081);
  and g4701 (n5082, n5073, n_2208);
  not g4702 (n_2209, pi1137);
  and g4703 (n5083, n_2209, n_29);
  not g4704 (n_2211, pi0933);
  and g4705 (n5084, n_2211, n2452);
  not g4706 (n_2212, n5083);
  and g4707 (n5085, pi0221, n_2212);
  not g4708 (n_2213, n5084);
  and g4709 (n5086, n_2213, n5085);
  not g4710 (n_2214, n5082);
  not g4711 (n_2215, n5086);
  and g4712 (n5087, n_2214, n_2215);
  not g4713 (n_2216, n5087);
  and g4714 (n5088, n_36, n_2216);
  not g4715 (n_2217, n5071);
  not g4716 (n_2218, n5088);
  and g4717 (n5089, n_2217, n_2218);
  and g4718 (n5090, n_826, n5089);
  not g4719 (n_2219, pi0878);
  and g4720 (n5091, n_2219, n2521);
  and g4721 (n5092, pi0168, n_207);
  not g4722 (n_2220, n5091);
  and g4723 (n5093, n_188, n_2220);
  not g4724 (n_2221, n5092);
  and g4725 (n5094, n_2221, n5093);
  not g4726 (n_2222, n5094);
  and g4727 (n5095, n5079, n_2222);
  not g4728 (n_2223, n5095);
  and g4729 (n5096, n5073, n_2223);
  not g4730 (n_2224, n5096);
  and g4731 (n5097, n_2215, n_2224);
  not g4732 (n_2225, n5097);
  and g4733 (n5098, n_36, n_2225);
  not g4734 (n_2226, n5098);
  and g4735 (n5099, n_2217, n_2226);
  and g4736 (n5100, n3331, n5099);
  not g4737 (n_2227, n5090);
  and g4738 (n5101, pi0062, n_2227);
  not g4739 (n_2228, n5100);
  and g4740 (n5102, n_2228, n5101);
  not g4741 (n_2229, n5089);
  and g4742 (n5103, n_179, n_2229);
  not g4743 (n_2230, n5099);
  and g4744 (n5104, n2537, n_2230);
  not g4745 (n_2231, n5103);
  and g4746 (n5105, pi0056, n_2231);
  not g4747 (n_2232, n5104);
  and g4748 (n5106, n_2232, n5105);
  and g4749 (n5107, n_204, n5089);
  and g4750 (n5108, n2572, n5099);
  not g4751 (n_2233, n5107);
  and g4752 (n5109, pi0055, n_2233);
  not g4753 (n_2234, n5108);
  and g4754 (n5110, n_2234, n5109);
  and g4755 (n5111, pi0223, pi1137);
  and g4756 (n5112, pi0224, pi0280);
  not g4757 (n_2235, n5112);
  and g4758 (n5113, n_226, n_2235);
  and g4759 (n5114, n_219, n_2202);
  not g4760 (n_2236, n5114);
  and g4761 (n5115, n5113, n_2236);
  and g4762 (n5116, n_2209, n_221);
  and g4763 (n5117, n_2211, n2591);
  not g4764 (n_2237, n5116);
  and g4765 (n5118, pi0222, n_2237);
  not g4766 (n_2238, n5117);
  and g4767 (n5119, n_2238, n5118);
  not g4768 (n_2239, n5115);
  not g4769 (n_2240, n5119);
  and g4770 (n5120, n_2239, n_2240);
  not g4771 (n_2241, n5120);
  and g4772 (n5121, n_223, n_2241);
  not g4773 (n_2242, n5111);
  not g4774 (n_2243, n5121);
  and g4775 (n5122, n_2242, n_2243);
  not g4776 (n_2244, n5122);
  and g4777 (n5123, n_234, n_2244);
  and g4778 (n5124, pi0299, n_2229);
  not g4779 (n_2245, n5123);
  not g4780 (n_2246, n5124);
  and g4781 (n5125, n_2245, n_2246);
  and g4782 (n5126, n_841, n5125);
  and g4783 (n5127, n_251, n5125);
  and g4784 (n5128, pi0299, n_2230);
  not g4785 (n_2247, n5128);
  and g4786 (n5129, n_2245, n_2247);
  and g4787 (n5130, n2625, n5129);
  not g4788 (n_2248, n5127);
  not g4789 (n_2249, n5130);
  and g4790 (n5131, n_2248, n_2249);
  not g4791 (n_2250, n5131);
  and g4792 (n5132, n2533, n_2250);
  and g4793 (n5133, n_257, n5125);
  not g4794 (n_2251, n5133);
  and g4795 (n5134, pi0092, n_2251);
  not g4796 (n_2252, n5132);
  and g4797 (n5135, n_2252, n5134);
  and g4798 (n5136, pi0075, n5125);
  and g4799 (n5137, pi0087, n5131);
  and g4800 (n5138, pi0038, n5125);
  not g4801 (n_2253, n5129);
  and g4802 (n5139, pi0039, n_2253);
  and g4803 (n5140, n_234, n_2242);
  and g4804 (n5141, pi0878, n3488);
  not g4805 (n_2254, n5141);
  and g4806 (n5142, n_219, n_2254);
  not g4807 (n_2255, n5142);
  and g4808 (n5143, n5113, n_2255);
  not g4809 (n_2256, n5143);
  and g4810 (n5144, n_2240, n_2256);
  and g4811 (n5145, n5140, n5144);
  and g4812 (n5146, pi0299, n_2217);
  and g4813 (n5147, pi0878, n3499);
  not g4814 (n_2257, n5147);
  and g4815 (n5148, n_2206, n_2257);
  and g4816 (n5149, pi0168, n3508);
  not g4817 (n_2258, n5148);
  not g4818 (n_2259, n5149);
  and g4819 (n5150, n_2258, n_2259);
  not g4820 (n_2260, n5150);
  and g4821 (n5151, pi0878, n_2260);
  and g4822 (n5152, n_879, n5148);
  not g4823 (n_2261, n5151);
  not g4824 (n_2262, n5152);
  and g4825 (n5153, n_2261, n_2262);
  not g4826 (n_2263, n5153);
  and g4827 (n5154, n_188, n_2263);
  and g4828 (n5155, n_937, n5078);
  not g4829 (n_2264, n5155);
  and g4830 (n5156, n_20, n_2264);
  not g4831 (n_2265, n5154);
  and g4832 (n5157, n_2265, n5156);
  not g4833 (n_2266, n5157);
  and g4834 (n5158, n5073, n_2266);
  not g4835 (n_2267, n5158);
  and g4836 (n5159, n_2215, n_2267);
  not g4837 (n_2268, n5159);
  and g4838 (n5160, n_36, n_2268);
  not g4839 (n_2269, n5160);
  and g4840 (n5161, n5146, n_2269);
  and g4841 (n5162, n_936, n5113);
  not g4842 (n_2270, n5162);
  and g4843 (n5163, n5144, n_2270);
  not g4844 (n_2271, n5163);
  and g4845 (n5164, n_223, n_2271);
  not g4846 (n_2272, n5164);
  and g4847 (n5165, n5140, n_2272);
  not g4848 (n_2273, n5165);
  and g4849 (n5166, n_162, n_2273);
  not g4850 (n_2274, n5145);
  and g4851 (n5167, n_2274, n5166);
  not g4852 (n_2275, n5161);
  and g4853 (n5168, n_2275, n5167);
  not g4854 (n_2276, n5139);
  and g4855 (n5169, n_161, n_2276);
  not g4856 (n_2277, n5168);
  and g4857 (n5170, n_2277, n5169);
  not g4858 (n_2278, n5138);
  and g4859 (n5171, n_164, n_2278);
  not g4860 (n_2279, n5170);
  and g4861 (n5172, n_2279, n5171);
  and g4862 (n5173, n_260, n5125);
  and g4863 (n5174, n_2219, n3394);
  and g4864 (n5175, pi0168, n_1567);
  not g4865 (n_2280, n5174);
  and g4866 (n5176, n_188, n_2280);
  not g4867 (n_2281, n5175);
  and g4868 (n5177, n_2281, n5176);
  not g4869 (n_2282, n5177);
  and g4870 (n5178, n5079, n_2282);
  not g4871 (n_2283, n5178);
  and g4872 (n5179, n5073, n_2283);
  not g4873 (n_2284, n5179);
  and g4874 (n5180, n_2215, n_2284);
  not g4875 (n_2285, n5180);
  and g4876 (n5181, n_36, n_2285);
  not g4877 (n_2286, n5181);
  and g4878 (n5182, n_2217, n_2286);
  not g4879 (n_2287, n5182);
  and g4880 (n5183, pi0299, n_2287);
  and g4881 (n5184, n2530, n_2245);
  not g4882 (n_2288, n5183);
  and g4883 (n5185, n_2288, n5184);
  not g4884 (n_2289, n5173);
  and g4885 (n5186, pi0100, n_2289);
  not g4886 (n_2290, n5185);
  and g4887 (n5187, n_2290, n5186);
  not g4888 (n_2291, n5172);
  not g4889 (n_2292, n5187);
  and g4890 (n5188, n_2291, n_2292);
  not g4891 (n_2293, n5188);
  and g4892 (n5189, n_172, n_2293);
  not g4893 (n_2294, n5137);
  and g4894 (n5190, n_171, n_2294);
  not g4895 (n_2295, n5189);
  and g4896 (n5191, n_2295, n5190);
  not g4897 (n_2296, n5136);
  and g4898 (n5192, n_174, n_2296);
  not g4899 (n_2297, n5191);
  and g4900 (n5193, n_2297, n5192);
  not g4901 (n_2298, n5135);
  and g4902 (n5194, n2532, n_2298);
  not g4903 (n_2299, n5193);
  and g4904 (n5195, n_2299, n5194);
  not g4905 (n_2300, n5126);
  and g4906 (n5196, n_176, n_2300);
  not g4907 (n_2301, n5195);
  and g4908 (n5197, n_2301, n5196);
  not g4909 (n_2302, n5110);
  and g4910 (n5198, n_157, n_2302);
  not g4911 (n_2303, n5197);
  and g4912 (n5199, n_2303, n5198);
  not g4913 (n_2304, n5106);
  and g4914 (n5200, n_158, n_2304);
  not g4915 (n_2305, n5199);
  and g4916 (n5201, n_2305, n5200);
  not g4917 (n_2307, pi0240);
  and g4923 (n5205, n_997, n5079);
  and g4924 (n5206, n_2222, n5205);
  not g4925 (n_2310, n5206);
  and g4926 (n5207, n5073, n_2310);
  not g4927 (n_2311, n5207);
  and g4928 (n5208, n_2215, n_2311);
  not g4929 (n_2312, n5208);
  and g4930 (n5209, n_36, n_2312);
  not g4931 (n_2313, n5209);
  and g4932 (n5210, n_2217, n_2313);
  and g4933 (n5211, n3331, n5210);
  and g4934 (n5212, n3556, n_2199);
  not g4935 (n_2314, n5212);
  and g4936 (n5213, n5089, n_2314);
  and g4937 (n5214, n_826, n5213);
  not g4938 (n_2315, n5214);
  and g4939 (n5215, pi0062, n_2315);
  not g4940 (n_2316, n5211);
  and g4941 (n5216, n_2316, n5215);
  not g4942 (n_2317, n5213);
  and g4943 (n5217, n_179, n_2317);
  not g4944 (n_2318, n5210);
  and g4945 (n5218, n2537, n_2318);
  not g4946 (n_2319, n5217);
  and g4947 (n5219, pi0056, n_2319);
  not g4948 (n_2320, n5218);
  and g4949 (n5220, n_2320, n5219);
  and g4950 (n5221, n2572, n5210);
  and g4951 (n5222, n_204, n5213);
  not g4952 (n_2321, n5222);
  and g4953 (n5223, pi0055, n_2321);
  not g4954 (n_2322, n5221);
  and g4955 (n5224, n_2322, n5223);
  and g4956 (n5225, n_921, n_2245);
  and g4957 (n5226, pi0299, n_2317);
  not g4958 (n_2323, n5226);
  and g4959 (n5227, n5225, n_2323);
  and g4960 (n5228, n_841, n5227);
  and g4961 (n5229, n_251, n5227);
  and g4962 (n5230, pi0299, n_2318);
  not g4963 (n_2324, n5230);
  and g4964 (n5231, n5225, n_2324);
  and g4965 (n5232, n2625, n5231);
  not g4966 (n_2325, n5229);
  not g4967 (n_2326, n5232);
  and g4968 (n5233, n_2325, n_2326);
  not g4969 (n_2327, n5233);
  and g4970 (n5234, n2533, n_2327);
  and g4971 (n5235, n_257, n5227);
  not g4972 (n_2328, n5235);
  and g4973 (n5236, pi0092, n_2328);
  not g4974 (n_2329, n5234);
  and g4975 (n5237, n_2329, n5236);
  and g4976 (n5238, pi0075, n5227);
  and g4977 (n5239, pi0087, n5233);
  and g4978 (n5240, pi0038, n5227);
  not g4979 (n_2330, n5231);
  and g4980 (n5241, pi0039, n_2330);
  and g4981 (n5242, n_2219, n3508);
  not g4982 (n_2331, n5242);
  and g4983 (n5243, n_2206, n_2331);
  and g4984 (n5244, n_2219, n_938);
  and g4985 (n5245, pi0878, n_879);
  not g4986 (n_2332, n5244);
  and g4987 (n5246, pi0168, n_2332);
  not g4988 (n_2333, n5245);
  and g4989 (n5247, n_2333, n5246);
  not g4990 (n_2334, n5243);
  not g4991 (n_2335, n5247);
  and g4992 (n5248, n_2334, n_2335);
  not g4993 (n_2336, n5248);
  and g4994 (n5249, n_188, n_2336);
  and g4995 (n5250, n_1181, n5079);
  not g4996 (n_2337, n5249);
  and g4997 (n5251, n_2337, n5250);
  not g4998 (n_2338, n5251);
  and g4999 (n5252, n5073, n_2338);
  not g5000 (n_2339, n5252);
  and g5001 (n5253, n_2215, n_2339);
  not g5002 (n_2340, n5253);
  and g5003 (n5254, n_36, n_2340);
  not g5004 (n_2341, n5254);
  and g5005 (n5255, n5146, n_2341);
  not g5006 (n_2342, n5255);
  and g5007 (n5256, n5166, n_2342);
  not g5008 (n_2343, n5241);
  and g5009 (n5257, n_161, n_2343);
  not g5010 (n_2344, n5256);
  and g5011 (n5258, n_2344, n5257);
  not g5012 (n_2345, n5240);
  and g5013 (n5259, n_164, n_2345);
  not g5014 (n_2346, n5258);
  and g5015 (n5260, n_2346, n5259);
  and g5016 (n5261, n_260, n5227);
  and g5017 (n5262, n_2282, n5205);
  not g5018 (n_2347, n5262);
  and g5019 (n5263, n5073, n_2347);
  not g5020 (n_2348, n5263);
  and g5021 (n5264, n_2215, n_2348);
  not g5022 (n_2349, n5264);
  and g5023 (n5265, n_36, n_2349);
  not g5024 (n_2350, n5265);
  and g5025 (n5266, n_2217, n_2350);
  not g5026 (n_2351, n5266);
  and g5027 (n5267, pi0299, n_2351);
  and g5028 (n5268, n2530, n5225);
  not g5029 (n_2352, n5267);
  and g5030 (n5269, n_2352, n5268);
  not g5031 (n_2353, n5261);
  and g5032 (n5270, pi0100, n_2353);
  not g5033 (n_2354, n5269);
  and g5034 (n5271, n_2354, n5270);
  not g5035 (n_2355, n5260);
  not g5036 (n_2356, n5271);
  and g5037 (n5272, n_2355, n_2356);
  not g5038 (n_2357, n5272);
  and g5039 (n5273, n_172, n_2357);
  not g5040 (n_2358, n5239);
  and g5041 (n5274, n_171, n_2358);
  not g5042 (n_2359, n5273);
  and g5043 (n5275, n_2359, n5274);
  not g5044 (n_2360, n5238);
  and g5045 (n5276, n_174, n_2360);
  not g5046 (n_2361, n5275);
  and g5047 (n5277, n_2361, n5276);
  not g5048 (n_2362, n5237);
  and g5049 (n5278, n2532, n_2362);
  not g5050 (n_2363, n5277);
  and g5051 (n5279, n_2363, n5278);
  not g5052 (n_2364, n5228);
  and g5053 (n5280, n_176, n_2364);
  not g5054 (n_2365, n5279);
  and g5055 (n5281, n_2365, n5280);
  not g5056 (n_2366, n5224);
  and g5057 (n5282, n_157, n_2366);
  not g5058 (n_2367, n5281);
  and g5059 (n5283, n_2367, n5282);
  not g5060 (n_2368, n5220);
  and g5061 (n5284, n_158, n_2368);
  not g5062 (n_2369, n5283);
  and g5063 (n5285, n_2369, n5284);
  and g5069 (n5289, pi0240, n5212);
  not g5070 (n_2372, n5289);
  and g5071 (n5290, n_824, n_2372);
  and g5072 (n5291, n5089, n5290);
  not g5073 (n_2373, n5288);
  not g5074 (n_2374, n5291);
  and g5075 (n5292, n_2373, n_2374);
  not g5076 (n_2375, n5204);
  and g5077 (po0162, n_2375, n5292);
  and g5078 (n5294, pi0215, pi1136);
  and g5079 (n5295, pi0216, pi0266);
  and g5080 (n5296, pi0875, n_145);
  not g5081 (n_2379, n5296);
  and g5082 (n5297, pi0105, n_2379);
  and g5083 (n5298, n_180, n_266);
  not g5084 (n_2380, n5297);
  not g5085 (n_2381, n5298);
  and g5086 (n5299, n_2380, n_2381);
  and g5087 (n5300, pi0228, n5299);
  and g5088 (n5301, pi0166, n_188);
  not g5089 (n_2382, n5300);
  not g5090 (n_2383, n5301);
  and g5091 (n5302, n_2382, n_2383);
  not g5092 (n_2384, n5302);
  and g5093 (n5303, n_20, n_2384);
  not g5094 (n_2385, n5295);
  not g5095 (n_2386, n5303);
  and g5096 (n5304, n_2385, n_2386);
  not g5097 (n_2387, n5304);
  and g5098 (n5305, n_26, n_2387);
  not g5099 (n_2388, pi1136);
  and g5100 (n5306, n_2388, n_29);
  not g5101 (n_2390, pi0928);
  and g5102 (n5307, n_2390, n2452);
  not g5103 (n_2391, n5306);
  and g5104 (n5308, pi0221, n_2391);
  not g5105 (n_2392, n5307);
  and g5106 (n5309, n_2392, n5308);
  not g5107 (n_2393, n5305);
  not g5108 (n_2394, n5309);
  and g5109 (n5310, n_2393, n_2394);
  not g5110 (n_2395, n5310);
  and g5111 (n5311, n_36, n_2395);
  not g5112 (n_2396, n5294);
  not g5113 (n_2397, n5311);
  and g5114 (n5312, n_2396, n_2397);
  and g5115 (n5313, n_824, n5312);
  and g5116 (n5314, n_826, n5312);
  and g5117 (n5315, n_266, n_207);
  not g5118 (n_2398, pi0875);
  and g5119 (n5316, n_2398, n2521);
  not g5120 (n_2399, n5315);
  and g5121 (n5317, n_188, n_2399);
  not g5122 (n_2400, n5316);
  and g5123 (n5318, n_2400, n5317);
  not g5124 (n_2401, n5318);
  and g5125 (n5319, n_2382, n_2401);
  not g5126 (n_2402, n5319);
  and g5127 (n5320, n_20, n_2402);
  not g5128 (n_2403, n5320);
  and g5129 (n5321, n_2385, n_2403);
  not g5130 (n_2404, n5321);
  and g5131 (n5322, n_26, n_2404);
  not g5132 (n_2405, n5322);
  and g5133 (n5323, n_2394, n_2405);
  not g5134 (n_2406, n5323);
  and g5135 (n5324, n_36, n_2406);
  not g5136 (n_2407, n5324);
  and g5137 (n5325, n_2396, n_2407);
  and g5138 (n5326, n3331, n5325);
  not g5139 (n_2408, n5314);
  and g5140 (n5327, pi0062, n_2408);
  not g5141 (n_2409, n5326);
  and g5142 (n5328, n_2409, n5327);
  not g5143 (n_2410, n5312);
  and g5144 (n5329, n_179, n_2410);
  not g5145 (n_2411, n5325);
  and g5146 (n5330, n2537, n_2411);
  not g5147 (n_2412, n5329);
  and g5148 (n5331, pi0056, n_2412);
  not g5149 (n_2413, n5330);
  and g5150 (n5332, n_2413, n5331);
  and g5151 (n5333, n_204, n5312);
  and g5152 (n5334, n2572, n5325);
  not g5153 (n_2414, n5333);
  and g5154 (n5335, pi0055, n_2414);
  not g5155 (n_2415, n5334);
  and g5156 (n5336, n_2415, n5335);
  and g5157 (n5337, pi0223, pi1136);
  not g5158 (n_2416, pi0266);
  and g5159 (n5338, pi0224, n_2416);
  and g5160 (n5339, n_219, n_2398);
  and g5161 (n5340, n_145, n5339);
  not g5162 (n_2417, n5338);
  and g5163 (n5341, n_226, n_2417);
  not g5164 (n_2418, n5340);
  and g5165 (n5342, n_2418, n5341);
  and g5166 (n5343, n_2388, n_221);
  and g5167 (n5344, n_2390, n2591);
  not g5168 (n_2419, n5343);
  and g5169 (n5345, pi0222, n_2419);
  not g5170 (n_2420, n5344);
  and g5171 (n5346, n_2420, n5345);
  not g5172 (n_2421, n5342);
  not g5173 (n_2422, n5346);
  and g5174 (n5347, n_2421, n_2422);
  not g5175 (n_2423, n5347);
  and g5176 (n5348, n_223, n_2423);
  not g5177 (n_2424, n5337);
  not g5178 (n_2425, n5348);
  and g5179 (n5349, n_2424, n_2425);
  not g5180 (n_2426, n5349);
  and g5181 (n5350, n_234, n_2426);
  and g5182 (n5351, n2604, n_2379);
  not g5183 (n_2427, n5351);
  and g5184 (n5352, n5350, n_2427);
  and g5185 (n5353, pi0299, n_2410);
  not g5186 (n_2428, n5352);
  not g5187 (n_2429, n5353);
  and g5188 (n5354, n_2428, n_2429);
  and g5189 (n5355, n_841, n5354);
  and g5190 (n5356, n_251, n5354);
  and g5191 (n5357, pi0299, n_2411);
  not g5192 (n_2430, n5357);
  and g5193 (n5358, n_2428, n_2430);
  and g5194 (n5359, n2625, n5358);
  not g5195 (n_2431, n5356);
  not g5196 (n_2432, n5359);
  and g5197 (n5360, n_2431, n_2432);
  not g5198 (n_2433, n5360);
  and g5199 (n5361, n2533, n_2433);
  and g5200 (n5362, n_257, n5354);
  not g5201 (n_2434, n5362);
  and g5202 (n5363, pi0092, n_2434);
  not g5203 (n_2435, n5361);
  and g5204 (n5364, n_2435, n5363);
  and g5205 (n5365, pi0075, n5354);
  and g5206 (n5366, pi0087, n5360);
  and g5207 (n5367, pi0038, n5354);
  not g5208 (n_2436, n5358);
  and g5209 (n5368, pi0039, n_2436);
  and g5210 (n5369, n2603, n_936);
  not g5211 (n_2437, n5369);
  and g5212 (n5370, n5342, n_2437);
  and g5213 (n5371, n_234, n_2424);
  and g5214 (n5372, n_2422, n5371);
  not g5215 (n_2438, n5370);
  and g5216 (n5373, n_2438, n5372);
  not g5217 (n_2439, n5299);
  and g5218 (n5374, n3498, n_2439);
  not g5219 (n_2440, n5374);
  and g5220 (n5375, n_20, n_2440);
  and g5221 (n5376, pi0166, n3499);
  and g5222 (n5377, n_266, n_1174);
  not g5223 (n_2441, n5376);
  and g5224 (n5378, pi0875, n_2441);
  not g5225 (n_2442, n5377);
  and g5226 (n5379, n_2442, n5378);
  and g5227 (n5380, pi0166, n_2398);
  and g5228 (n5381, n_879, n5380);
  not g5229 (n_2443, n5379);
  not g5230 (n_2444, n5381);
  and g5231 (n5382, n_2443, n_2444);
  not g5232 (n_2445, n5382);
  and g5233 (n5383, n_188, n_2445);
  not g5234 (n_2446, n5383);
  and g5235 (n5384, n_939, n_2446);
  not g5236 (n_2447, n5384);
  and g5237 (n5385, n5375, n_2447);
  not g5238 (n_2448, n5385);
  and g5239 (n5386, n_2385, n_2448);
  not g5240 (n_2449, n5386);
  and g5241 (n5387, n_26, n_2449);
  not g5242 (n_2450, n5387);
  and g5243 (n5388, n_2394, n_2450);
  not g5244 (n_2451, n5388);
  and g5245 (n5389, n_36, n_2451);
  and g5246 (n5390, pi0299, n_2396);
  not g5247 (n_2452, n5389);
  and g5248 (n5391, n_2452, n5390);
  and g5249 (n5392, n5347, n_2437);
  not g5250 (n_2453, n5392);
  and g5251 (n5393, n_223, n_2453);
  not g5252 (n_2454, n5393);
  and g5253 (n5394, n5371, n_2454);
  not g5254 (n_2455, n5394);
  and g5255 (n5395, n_162, n_2455);
  not g5256 (n_2456, n5373);
  and g5257 (n5396, n_2456, n5395);
  not g5258 (n_2457, n5391);
  and g5259 (n5397, n_2457, n5396);
  not g5260 (n_2458, n5368);
  and g5261 (n5398, n_161, n_2458);
  not g5262 (n_2459, n5397);
  and g5263 (n5399, n_2459, n5398);
  not g5264 (n_2460, n5367);
  and g5265 (n5400, n_164, n_2460);
  not g5266 (n_2461, n5399);
  and g5267 (n5401, n_2461, n5400);
  and g5268 (n5402, n_260, n5354);
  and g5269 (n5403, n_2398, n3387);
  not g5270 (n_2462, n5403);
  and g5271 (n5404, pi0166, n_2462);
  not g5272 (n_2463, n2638);
  and g5273 (n5405, n_2463, n_858);
  and g5274 (n5406, n2638, n_855);
  not g5275 (n_2464, n5406);
  and g5276 (n5407, pi0875, n_2464);
  not g5277 (n_2465, n5405);
  and g5278 (n5408, n_2465, n5407);
  not g5279 (n_2466, n5404);
  not g5280 (n_2467, n5408);
  and g5281 (n5409, n_2466, n_2467);
  not g5282 (n_2468, n5409);
  and g5283 (n5410, n_188, n_2468);
  not g5284 (n_2469, n5410);
  and g5285 (n5411, n_2382, n_2469);
  not g5286 (n_2470, n5411);
  and g5287 (n5412, n_20, n_2470);
  not g5288 (n_2471, n5412);
  and g5289 (n5413, n_2385, n_2471);
  not g5290 (n_2472, n5413);
  and g5291 (n5414, n_26, n_2472);
  not g5292 (n_2473, n5414);
  and g5293 (n5415, n_2394, n_2473);
  not g5294 (n_2474, n5415);
  and g5295 (n5416, n_36, n_2474);
  not g5296 (n_2475, n5416);
  and g5297 (n5417, n_2396, n_2475);
  not g5298 (n_2476, n5417);
  and g5299 (n5418, pi0299, n_2476);
  and g5300 (n5419, n2530, n_2428);
  not g5301 (n_2477, n5418);
  and g5302 (n5420, n_2477, n5419);
  not g5303 (n_2478, n5402);
  and g5304 (n5421, pi0100, n_2478);
  not g5305 (n_2479, n5420);
  and g5306 (n5422, n_2479, n5421);
  not g5307 (n_2480, n5401);
  not g5308 (n_2481, n5422);
  and g5309 (n5423, n_2480, n_2481);
  not g5310 (n_2482, n5423);
  and g5311 (n5424, n_172, n_2482);
  not g5312 (n_2483, n5366);
  and g5313 (n5425, n_171, n_2483);
  not g5314 (n_2484, n5424);
  and g5315 (n5426, n_2484, n5425);
  not g5316 (n_2485, n5365);
  and g5317 (n5427, n_174, n_2485);
  not g5318 (n_2486, n5426);
  and g5319 (n5428, n_2486, n5427);
  not g5320 (n_2487, n5364);
  and g5321 (n5429, n2532, n_2487);
  not g5322 (n_2488, n5428);
  and g5323 (n5430, n_2488, n5429);
  not g5324 (n_2489, n5355);
  and g5325 (n5431, n_176, n_2489);
  not g5326 (n_2490, n5430);
  and g5327 (n5432, n_2490, n5431);
  not g5328 (n_2491, n5336);
  and g5329 (n5433, n_157, n_2491);
  not g5330 (n_2492, n5432);
  and g5331 (n5434, n_2492, n5433);
  not g5332 (n_2493, n5332);
  and g5333 (n5435, n_158, n_2493);
  not g5334 (n_2494, n5434);
  and g5335 (n5436, n_2494, n5435);
  not g5336 (n_2495, n5328);
  and g5337 (n5437, n3328, n_2495);
  not g5338 (n_2496, n5436);
  and g5339 (n5438, n_2496, n5437);
  not g5340 (n_2498, pi0245);
  not g5341 (n_2499, n5313);
  and g5342 (n5439, n_2498, n_2499);
  not g5343 (n_2500, n5438);
  and g5344 (n5440, n_2500, n5439);
  and g5345 (n5441, n_909, n5312);
  and g5346 (n5442, n_824, n5441);
  and g5347 (n5443, n_997, n_2382);
  and g5348 (n5444, n_2401, n5443);
  not g5349 (n_2501, n5444);
  and g5350 (n5445, n_20, n_2501);
  not g5351 (n_2502, n5445);
  and g5352 (n5446, n_2385, n_2502);
  not g5353 (n_2503, n5446);
  and g5354 (n5447, n_26, n_2503);
  not g5355 (n_2504, n5447);
  and g5356 (n5448, n_2394, n_2504);
  not g5357 (n_2505, n5448);
  and g5358 (n5449, n_36, n_2505);
  not g5359 (n_2506, n5449);
  and g5360 (n5450, n_2396, n_2506);
  and g5361 (n5451, n3331, n5450);
  and g5362 (n5452, n_826, n5441);
  not g5363 (n_2507, n5452);
  and g5364 (n5453, pi0062, n_2507);
  not g5365 (n_2508, n5451);
  and g5366 (n5454, n_2508, n5453);
  not g5367 (n_2509, n5441);
  and g5368 (n5455, n_179, n_2509);
  not g5369 (n_2510, n5450);
  and g5370 (n5456, n2537, n_2510);
  not g5371 (n_2511, n5455);
  and g5372 (n5457, pi0056, n_2511);
  not g5373 (n_2512, n5456);
  and g5374 (n5458, n_2512, n5457);
  and g5375 (n5459, n2572, n5450);
  and g5376 (n5460, n_204, n5441);
  not g5377 (n_2513, n5460);
  and g5378 (n5461, pi0055, n_2513);
  not g5379 (n_2514, n5459);
  and g5380 (n5462, n_2514, n5461);
  and g5381 (n5463, pi0299, n_2509);
  not g5382 (n_2515, n5350);
  not g5383 (n_2516, n5463);
  and g5384 (n5464, n_2515, n_2516);
  and g5385 (n5465, n_841, n5464);
  and g5386 (n5466, n_251, n5464);
  and g5387 (n5467, pi0299, n_2510);
  not g5388 (n_2517, n5467);
  and g5389 (n5468, n_2515, n_2517);
  and g5390 (n5469, n2625, n5468);
  not g5391 (n_2518, n5466);
  not g5392 (n_2519, n5469);
  and g5393 (n5470, n_2518, n_2519);
  not g5394 (n_2520, n5470);
  and g5395 (n5471, n2533, n_2520);
  and g5396 (n5472, n_257, n5464);
  not g5397 (n_2521, n5472);
  and g5398 (n5473, pi0092, n_2521);
  not g5399 (n_2522, n5471);
  and g5400 (n5474, n_2522, n5473);
  and g5401 (n5475, pi0075, n5464);
  and g5402 (n5476, pi0087, n5470);
  and g5403 (n5477, pi0038, n5464);
  not g5404 (n_2523, n5468);
  and g5405 (n5478, pi0039, n_2523);
  and g5406 (n5479, n_266, n_938);
  and g5407 (n5480, pi0166, n3508);
  not g5408 (n_2524, n5479);
  and g5409 (n5481, n_2398, n_2524);
  not g5410 (n_2525, n5480);
  and g5411 (n5482, n_2525, n5481);
  and g5412 (n5483, n_266, n_879);
  not g5413 (n_2526, n5483);
  and g5414 (n5484, pi0875, n_2526);
  not g5415 (n_2527, n5482);
  and g5416 (n5485, n_188, n_2527);
  not g5417 (n_2528, n5484);
  and g5418 (n5486, n_2528, n5485);
  not g5419 (n_2529, n5486);
  and g5420 (n5487, n5375, n_2529);
  not g5421 (n_2530, n5487);
  and g5422 (n5488, n_2385, n_2530);
  not g5423 (n_2531, n5488);
  and g5424 (n5489, n_26, n_2531);
  not g5425 (n_2532, n5489);
  and g5426 (n5490, n_2394, n_2532);
  not g5427 (n_2533, n5490);
  and g5428 (n5491, n_36, n_2533);
  not g5429 (n_2534, n5491);
  and g5430 (n5492, n5390, n_2534);
  not g5431 (n_2535, n5492);
  and g5432 (n5493, n5395, n_2535);
  not g5433 (n_2536, n5478);
  and g5434 (n5494, n_161, n_2536);
  not g5435 (n_2537, n5493);
  and g5436 (n5495, n_2537, n5494);
  not g5437 (n_2538, n5477);
  and g5438 (n5496, n_164, n_2538);
  not g5439 (n_2539, n5495);
  and g5440 (n5497, n_2539, n5496);
  and g5441 (n5498, n_260, n5464);
  and g5442 (n5499, n_2469, n5443);
  not g5443 (n_2540, n5499);
  and g5444 (n5500, n_20, n_2540);
  not g5445 (n_2541, n5500);
  and g5446 (n5501, n_2385, n_2541);
  not g5447 (n_2542, n5501);
  and g5448 (n5502, n_26, n_2542);
  not g5449 (n_2543, n5502);
  and g5450 (n5503, n_2394, n_2543);
  not g5451 (n_2544, n5503);
  and g5452 (n5504, n_36, n_2544);
  not g5453 (n_2545, n5504);
  and g5454 (n5505, n_2396, n_2545);
  not g5455 (n_2546, n5505);
  and g5456 (n5506, pi0299, n_2546);
  and g5457 (n5507, n2530, n_2515);
  not g5458 (n_2547, n5506);
  and g5459 (n5508, n_2547, n5507);
  not g5460 (n_2548, n5498);
  and g5461 (n5509, pi0100, n_2548);
  not g5462 (n_2549, n5508);
  and g5463 (n5510, n_2549, n5509);
  not g5464 (n_2550, n5497);
  not g5465 (n_2551, n5510);
  and g5466 (n5511, n_2550, n_2551);
  not g5467 (n_2552, n5511);
  and g5468 (n5512, n_172, n_2552);
  not g5469 (n_2553, n5476);
  and g5470 (n5513, n_171, n_2553);
  not g5471 (n_2554, n5512);
  and g5472 (n5514, n_2554, n5513);
  not g5473 (n_2555, n5475);
  and g5474 (n5515, n_174, n_2555);
  not g5475 (n_2556, n5514);
  and g5476 (n5516, n_2556, n5515);
  not g5477 (n_2557, n5474);
  and g5478 (n5517, n2532, n_2557);
  not g5479 (n_2558, n5516);
  and g5480 (n5518, n_2558, n5517);
  not g5481 (n_2559, n5465);
  and g5482 (n5519, n_176, n_2559);
  not g5483 (n_2560, n5518);
  and g5484 (n5520, n_2560, n5519);
  not g5485 (n_2561, n5462);
  and g5486 (n5521, n_157, n_2561);
  not g5487 (n_2562, n5520);
  and g5488 (n5522, n_2562, n5521);
  not g5489 (n_2563, n5458);
  and g5490 (n5523, n_158, n_2563);
  not g5491 (n_2564, n5522);
  and g5492 (n5524, n_2564, n5523);
  not g5493 (n_2565, n5454);
  and g5494 (n5525, n3328, n_2565);
  not g5495 (n_2566, n5524);
  and g5496 (n5526, n_2566, n5525);
  not g5497 (n_2567, n5442);
  and g5498 (n5527, pi0245, n_2567);
  not g5499 (n_2568, n5526);
  and g5500 (n5528, n_2568, n5527);
  or g5501 (po0163, n5440, n5528);
  and g5502 (n5530, pi0215, pi1135);
  and g5503 (n5531, pi0216, pi0279);
  and g5504 (n5532, pi0879, n_145);
  not g5505 (n_2572, n5532);
  and g5506 (n5533, pi0105, n_2572);
  and g5507 (n5534, n_180, n_264);
  not g5508 (n_2573, n5533);
  not g5509 (n_2574, n5534);
  and g5510 (n5535, n_2573, n_2574);
  and g5511 (n5536, pi0228, n5535);
  and g5512 (n5537, pi0161, n_188);
  not g5513 (n_2575, n5536);
  not g5514 (n_2576, n5537);
  and g5515 (n5538, n_2575, n_2576);
  not g5516 (n_2577, n5538);
  and g5517 (n5539, n_20, n_2577);
  not g5518 (n_2578, n5531);
  not g5519 (n_2579, n5539);
  and g5520 (n5540, n_2578, n_2579);
  not g5521 (n_2580, n5540);
  and g5522 (n5541, n_26, n_2580);
  not g5523 (n_2581, pi1135);
  and g5524 (n5542, n_2581, n_29);
  not g5525 (n_2583, pi0938);
  and g5526 (n5543, n_2583, n2452);
  not g5527 (n_2584, n5542);
  and g5528 (n5544, pi0221, n_2584);
  not g5529 (n_2585, n5543);
  and g5530 (n5545, n_2585, n5544);
  not g5531 (n_2586, n5541);
  not g5532 (n_2587, n5545);
  and g5533 (n5546, n_2586, n_2587);
  not g5534 (n_2588, n5546);
  and g5535 (n5547, n_36, n_2588);
  not g5536 (n_2589, n5530);
  not g5537 (n_2590, n5547);
  and g5538 (n5548, n_2589, n_2590);
  and g5539 (n5549, n_824, n5548);
  and g5540 (n5550, n_826, n5548);
  not g5541 (n_2591, pi0879);
  and g5542 (n5551, n_2591, n2521);
  and g5543 (n5552, n_1324, n_2576);
  not g5544 (n_2592, n5551);
  not g5545 (n_2593, n5552);
  and g5546 (n5553, n_2592, n_2593);
  not g5547 (n_2594, n5553);
  and g5548 (n5554, n_2575, n_2594);
  not g5549 (n_2595, n5554);
  and g5550 (n5555, n_20, n_2595);
  not g5551 (n_2596, n5555);
  and g5552 (n5556, n_2578, n_2596);
  not g5553 (n_2597, n5556);
  and g5554 (n5557, n_26, n_2597);
  not g5555 (n_2598, n5557);
  and g5556 (n5558, n_2587, n_2598);
  not g5557 (n_2599, n5558);
  and g5558 (n5559, n_36, n_2599);
  not g5559 (n_2600, n5559);
  and g5560 (n5560, n_2589, n_2600);
  and g5561 (n5561, n3331, n5560);
  not g5562 (n_2601, n5550);
  and g5563 (n5562, pi0062, n_2601);
  not g5564 (n_2602, n5561);
  and g5565 (n5563, n_2602, n5562);
  not g5566 (n_2603, n5548);
  and g5567 (n5564, n_179, n_2603);
  not g5568 (n_2604, n5560);
  and g5569 (n5565, n2537, n_2604);
  not g5570 (n_2605, n5564);
  and g5571 (n5566, pi0056, n_2605);
  not g5572 (n_2606, n5565);
  and g5573 (n5567, n_2606, n5566);
  and g5574 (n5568, n_204, n5548);
  and g5575 (n5569, n2572, n5560);
  not g5576 (n_2607, n5568);
  and g5577 (n5570, pi0055, n_2607);
  not g5578 (n_2608, n5569);
  and g5579 (n5571, n_2608, n5570);
  and g5580 (n5572, pi0223, pi1135);
  and g5581 (n5573, n_2581, n_221);
  and g5582 (n5574, n_2583, n2591);
  not g5583 (n_2609, n5573);
  and g5584 (n5575, pi0222, n_2609);
  not g5585 (n_2610, n5574);
  and g5586 (n5576, n_2610, n5575);
  not g5587 (n_2611, pi0279);
  and g5588 (n5577, pi0224, n_2611);
  and g5589 (n5578, n_219, n_2591);
  and g5590 (n5579, n_145, n5578);
  not g5591 (n_2612, n5577);
  and g5592 (n5580, n_226, n_2612);
  not g5593 (n_2613, n5579);
  and g5594 (n5581, n_2613, n5580);
  not g5595 (n_2614, n5576);
  not g5596 (n_2615, n5581);
  and g5597 (n5582, n_2614, n_2615);
  not g5598 (n_2616, n5582);
  and g5599 (n5583, n_223, n_2616);
  not g5600 (n_2617, n5572);
  not g5601 (n_2618, n5583);
  and g5602 (n5584, n_2617, n_2618);
  not g5603 (n_2619, n5584);
  and g5604 (n5585, n_234, n_2619);
  and g5605 (n5586, n2604, n_2572);
  not g5606 (n_2620, n5586);
  and g5607 (n5587, n5585, n_2620);
  and g5608 (n5588, pi0299, n_2603);
  not g5609 (n_2621, n5587);
  not g5610 (n_2622, n5588);
  and g5611 (n5589, n_2621, n_2622);
  and g5612 (n5590, n_841, n5589);
  and g5613 (n5591, n_251, n5589);
  and g5614 (n5592, pi0299, n_2604);
  not g5615 (n_2623, n5592);
  and g5616 (n5593, n_2621, n_2623);
  and g5617 (n5594, n2625, n5593);
  not g5618 (n_2624, n5591);
  not g5619 (n_2625, n5594);
  and g5620 (n5595, n_2624, n_2625);
  not g5621 (n_2626, n5595);
  and g5622 (n5596, n2533, n_2626);
  and g5623 (n5597, n_257, n5589);
  not g5624 (n_2627, n5597);
  and g5625 (n5598, pi0092, n_2627);
  not g5626 (n_2628, n5596);
  and g5627 (n5599, n_2628, n5598);
  and g5628 (n5600, pi0075, n5589);
  and g5629 (n5601, pi0087, n5595);
  and g5630 (n5602, pi0038, n5589);
  not g5631 (n_2629, n5593);
  and g5632 (n5603, pi0039, n_2629);
  and g5633 (n5604, n_234, n_2617);
  and g5634 (n5605, n5369, n_2614);
  not g5635 (n_2630, n5605);
  and g5636 (n5606, n5583, n_2630);
  not g5637 (n_2631, n5606);
  and g5638 (n5607, n5604, n_2631);
  not g5639 (n_2632, n5535);
  and g5640 (n5608, n3498, n_2632);
  not g5641 (n_2633, n5608);
  and g5642 (n5609, n_20, n_2633);
  and g5643 (n5610, pi0161, n3499);
  and g5644 (n5611, n_264, n_1174);
  not g5645 (n_2634, n5610);
  and g5646 (n5612, pi0879, n_2634);
  not g5647 (n_2635, n5611);
  and g5648 (n5613, n_2635, n5612);
  and g5649 (n5614, pi0161, n_2591);
  and g5650 (n5615, n_879, n5614);
  not g5651 (n_2636, n5613);
  not g5652 (n_2637, n5615);
  and g5653 (n5616, n_2636, n_2637);
  not g5654 (n_2638, n5616);
  and g5655 (n5617, n_188, n_2638);
  not g5656 (n_2639, n5617);
  and g5657 (n5618, n_939, n_2639);
  not g5658 (n_2640, n5618);
  and g5659 (n5619, n5609, n_2640);
  not g5660 (n_2641, n5619);
  and g5661 (n5620, n_2578, n_2641);
  not g5662 (n_2642, n5620);
  and g5663 (n5621, n_26, n_2642);
  not g5664 (n_2643, n5621);
  and g5665 (n5622, n_2587, n_2643);
  not g5666 (n_2644, n5622);
  and g5667 (n5623, n_36, n_2644);
  and g5668 (n5624, pi0299, n_2589);
  not g5669 (n_2645, n5623);
  and g5670 (n5625, n_2645, n5624);
  not g5671 (n_2646, n5607);
  and g5672 (n5626, n_162, n_2646);
  not g5673 (n_2647, n5625);
  and g5674 (n5627, n_2647, n5626);
  not g5675 (n_2648, n5603);
  and g5676 (n5628, n_161, n_2648);
  not g5677 (n_2649, n5627);
  and g5678 (n5629, n_2649, n5628);
  not g5679 (n_2650, n5602);
  and g5680 (n5630, n_164, n_2650);
  not g5681 (n_2651, n5629);
  and g5682 (n5631, n_2651, n5630);
  and g5683 (n5632, n_260, n5589);
  and g5684 (n5633, n_2591, n3387);
  not g5685 (n_2652, n5633);
  and g5686 (n5634, pi0161, n_2652);
  and g5687 (n5635, n_263, n_266);
  and g5688 (n5636, n_855, n5635);
  not g5689 (n_2653, n5635);
  and g5690 (n5637, n_858, n_2653);
  not g5691 (n_2654, n5636);
  and g5692 (n5638, pi0879, n_2654);
  not g5693 (n_2655, n5637);
  and g5694 (n5639, n_2655, n5638);
  not g5695 (n_2656, n5634);
  not g5696 (n_2657, n5639);
  and g5697 (n5640, n_2656, n_2657);
  not g5698 (n_2658, n5640);
  and g5699 (n5641, n_188, n_2658);
  not g5700 (n_2659, n5641);
  and g5701 (n5642, n_2575, n_2659);
  not g5702 (n_2660, n5642);
  and g5703 (n5643, n_20, n_2660);
  not g5704 (n_2661, n5643);
  and g5705 (n5644, n_2578, n_2661);
  not g5706 (n_2662, n5644);
  and g5707 (n5645, n_26, n_2662);
  not g5708 (n_2663, n5645);
  and g5709 (n5646, n_2587, n_2663);
  not g5710 (n_2664, n5646);
  and g5711 (n5647, n_36, n_2664);
  not g5712 (n_2665, n5647);
  and g5713 (n5648, n_2589, n_2665);
  not g5714 (n_2666, n5648);
  and g5715 (n5649, pi0299, n_2666);
  and g5716 (n5650, n2530, n_2621);
  not g5717 (n_2667, n5649);
  and g5718 (n5651, n_2667, n5650);
  not g5719 (n_2668, n5632);
  and g5720 (n5652, pi0100, n_2668);
  not g5721 (n_2669, n5651);
  and g5722 (n5653, n_2669, n5652);
  not g5723 (n_2670, n5631);
  not g5724 (n_2671, n5653);
  and g5725 (n5654, n_2670, n_2671);
  not g5726 (n_2672, n5654);
  and g5727 (n5655, n_172, n_2672);
  not g5728 (n_2673, n5601);
  and g5729 (n5656, n_171, n_2673);
  not g5730 (n_2674, n5655);
  and g5731 (n5657, n_2674, n5656);
  not g5732 (n_2675, n5600);
  and g5733 (n5658, n_174, n_2675);
  not g5734 (n_2676, n5657);
  and g5735 (n5659, n_2676, n5658);
  not g5736 (n_2677, n5599);
  and g5737 (n5660, n2532, n_2677);
  not g5738 (n_2678, n5659);
  and g5739 (n5661, n_2678, n5660);
  not g5740 (n_2679, n5590);
  and g5741 (n5662, n_176, n_2679);
  not g5742 (n_2680, n5661);
  and g5743 (n5663, n_2680, n5662);
  not g5744 (n_2681, n5571);
  and g5745 (n5664, n_157, n_2681);
  not g5746 (n_2682, n5663);
  and g5747 (n5665, n_2682, n5664);
  not g5748 (n_2683, n5567);
  and g5749 (n5666, n_158, n_2683);
  not g5750 (n_2684, n5665);
  and g5751 (n5667, n_2684, n5666);
  not g5752 (n_2685, n5563);
  and g5753 (n5668, n3328, n_2685);
  not g5754 (n_2686, n5667);
  and g5755 (n5669, n_2686, n5668);
  not g5756 (n_2688, pi0244);
  not g5757 (n_2689, n5549);
  and g5758 (n5670, n_2688, n_2689);
  not g5759 (n_2690, n5669);
  and g5760 (n5671, n_2690, n5670);
  and g5761 (n5672, n_909, n5548);
  and g5762 (n5673, n_824, n5672);
  and g5763 (n5674, n_997, n_2575);
  and g5764 (n5675, n_2594, n5674);
  not g5765 (n_2691, n5675);
  and g5766 (n5676, n_20, n_2691);
  not g5767 (n_2692, n5676);
  and g5768 (n5677, n_2578, n_2692);
  not g5769 (n_2693, n5677);
  and g5770 (n5678, n_26, n_2693);
  not g5771 (n_2694, n5678);
  and g5772 (n5679, n_2587, n_2694);
  not g5773 (n_2695, n5679);
  and g5774 (n5680, n_36, n_2695);
  not g5775 (n_2696, n5680);
  and g5776 (n5681, n_2589, n_2696);
  and g5777 (n5682, n3331, n5681);
  and g5778 (n5683, n_826, n5672);
  not g5779 (n_2697, n5683);
  and g5780 (n5684, pi0062, n_2697);
  not g5781 (n_2698, n5682);
  and g5782 (n5685, n_2698, n5684);
  not g5783 (n_2699, n5672);
  and g5784 (n5686, n_179, n_2699);
  not g5785 (n_2700, n5681);
  and g5786 (n5687, n2537, n_2700);
  not g5787 (n_2701, n5686);
  and g5788 (n5688, pi0056, n_2701);
  not g5789 (n_2702, n5687);
  and g5790 (n5689, n_2702, n5688);
  and g5791 (n5690, n2572, n5681);
  and g5792 (n5691, n_204, n5672);
  not g5793 (n_2703, n5691);
  and g5794 (n5692, pi0055, n_2703);
  not g5795 (n_2704, n5690);
  and g5796 (n5693, n_2704, n5692);
  and g5797 (n5694, pi0299, n_2699);
  not g5798 (n_2705, n5585);
  not g5799 (n_2706, n5694);
  and g5800 (n5695, n_2705, n_2706);
  and g5801 (n5696, n_841, n5695);
  and g5802 (n5697, n_251, n5695);
  and g5803 (n5698, pi0299, n_2700);
  not g5804 (n_2707, n5698);
  and g5805 (n5699, n_2705, n_2707);
  and g5806 (n5700, n2625, n5699);
  not g5807 (n_2708, n5697);
  not g5808 (n_2709, n5700);
  and g5809 (n5701, n_2708, n_2709);
  not g5810 (n_2710, n5701);
  and g5811 (n5702, n2533, n_2710);
  and g5812 (n5703, n_257, n5695);
  not g5813 (n_2711, n5703);
  and g5814 (n5704, pi0092, n_2711);
  not g5815 (n_2712, n5702);
  and g5816 (n5705, n_2712, n5704);
  and g5817 (n5706, pi0075, n5695);
  and g5818 (n5707, pi0087, n5701);
  and g5819 (n5708, pi0038, n5695);
  not g5820 (n_2713, n5699);
  and g5821 (n5709, pi0039, n_2713);
  and g5822 (n5710, n_2437, n5582);
  not g5823 (n_2714, n5710);
  and g5824 (n5711, n_223, n_2714);
  not g5825 (n_2715, n5711);
  and g5826 (n5712, n5604, n_2715);
  and g5827 (n5713, n_264, n_938);
  and g5828 (n5714, pi0161, n3508);
  not g5829 (n_2716, n5713);
  and g5830 (n5715, n_2591, n_2716);
  not g5831 (n_2717, n5714);
  and g5832 (n5716, n_2717, n5715);
  and g5833 (n5717, n_264, n_879);
  not g5834 (n_2718, n5717);
  and g5835 (n5718, pi0879, n_2718);
  not g5836 (n_2719, n5716);
  and g5837 (n5719, n_188, n_2719);
  not g5838 (n_2720, n5718);
  and g5839 (n5720, n_2720, n5719);
  not g5840 (n_2721, n5720);
  and g5841 (n5721, n5609, n_2721);
  not g5842 (n_2722, n5721);
  and g5843 (n5722, n_2578, n_2722);
  not g5844 (n_2723, n5722);
  and g5845 (n5723, n_26, n_2723);
  not g5846 (n_2724, n5723);
  and g5847 (n5724, n_2587, n_2724);
  not g5848 (n_2725, n5724);
  and g5849 (n5725, n_36, n_2725);
  not g5850 (n_2726, n5725);
  and g5851 (n5726, n5624, n_2726);
  not g5852 (n_2727, n5712);
  and g5853 (n5727, n_162, n_2727);
  not g5854 (n_2728, n5726);
  and g5855 (n5728, n_2728, n5727);
  not g5856 (n_2729, n5709);
  and g5857 (n5729, n_161, n_2729);
  not g5858 (n_2730, n5728);
  and g5859 (n5730, n_2730, n5729);
  not g5860 (n_2731, n5708);
  and g5861 (n5731, n_164, n_2731);
  not g5862 (n_2732, n5730);
  and g5863 (n5732, n_2732, n5731);
  and g5864 (n5733, n_260, n5695);
  and g5865 (n5734, n_2659, n5674);
  not g5866 (n_2733, n5734);
  and g5867 (n5735, n_20, n_2733);
  not g5868 (n_2734, n5735);
  and g5869 (n5736, n_2578, n_2734);
  not g5870 (n_2735, n5736);
  and g5871 (n5737, n_26, n_2735);
  not g5872 (n_2736, n5737);
  and g5873 (n5738, n_2587, n_2736);
  not g5874 (n_2737, n5738);
  and g5875 (n5739, n_36, n_2737);
  not g5876 (n_2738, n5739);
  and g5877 (n5740, n_2589, n_2738);
  not g5878 (n_2739, n5740);
  and g5879 (n5741, pi0299, n_2739);
  and g5880 (n5742, n2530, n_2705);
  not g5881 (n_2740, n5741);
  and g5882 (n5743, n_2740, n5742);
  not g5883 (n_2741, n5733);
  and g5884 (n5744, pi0100, n_2741);
  not g5885 (n_2742, n5743);
  and g5886 (n5745, n_2742, n5744);
  not g5887 (n_2743, n5732);
  not g5888 (n_2744, n5745);
  and g5889 (n5746, n_2743, n_2744);
  not g5890 (n_2745, n5746);
  and g5891 (n5747, n_172, n_2745);
  not g5892 (n_2746, n5707);
  and g5893 (n5748, n_171, n_2746);
  not g5894 (n_2747, n5747);
  and g5895 (n5749, n_2747, n5748);
  not g5896 (n_2748, n5706);
  and g5897 (n5750, n_174, n_2748);
  not g5898 (n_2749, n5749);
  and g5899 (n5751, n_2749, n5750);
  not g5900 (n_2750, n5705);
  and g5901 (n5752, n2532, n_2750);
  not g5902 (n_2751, n5751);
  and g5903 (n5753, n_2751, n5752);
  not g5904 (n_2752, n5696);
  and g5905 (n5754, n_176, n_2752);
  not g5906 (n_2753, n5753);
  and g5907 (n5755, n_2753, n5754);
  not g5908 (n_2754, n5693);
  and g5909 (n5756, n_157, n_2754);
  not g5910 (n_2755, n5755);
  and g5911 (n5757, n_2755, n5756);
  not g5912 (n_2756, n5689);
  and g5913 (n5758, n_158, n_2756);
  not g5914 (n_2757, n5757);
  and g5915 (n5759, n_2757, n5758);
  not g5916 (n_2758, n5685);
  and g5917 (n5760, n3328, n_2758);
  not g5918 (n_2759, n5759);
  and g5919 (n5761, n_2759, n5760);
  not g5920 (n_2760, n5673);
  and g5921 (n5762, pi0244, n_2760);
  not g5922 (n_2761, n5761);
  and g5923 (n5763, n_2761, n5762);
  or g5924 (po0164, n5671, n5763);
  and g5925 (n5765, pi0216, pi0278);
  not g5926 (n_2763, n5765);
  and g5927 (n5766, n_26, n_2763);
  and g5928 (n5767, n_180, pi0152);
  and g5929 (n5768, pi0846, n_145);
  and g5930 (n5769, pi0105, n5768);
  not g5931 (n_2765, n5767);
  not g5932 (n_2766, n5769);
  and g5933 (n5770, n_2765, n_2766);
  not g5934 (n_2767, n5770);
  and g5935 (n5771, pi0228, n_2767);
  and g5936 (n5772, pi0152, n_188);
  not g5937 (n_2768, n5771);
  not g5938 (n_2769, n5772);
  and g5939 (n5773, n_2768, n_2769);
  not g5940 (n_2770, n5773);
  and g5941 (n5774, n_20, n_2770);
  not g5942 (n_2771, n5774);
  and g5943 (n5775, n5766, n_2771);
  not g5944 (n_2773, pi0930);
  and g5945 (n5776, pi0833, n_2773);
  and g5946 (n5777, n_20, pi0221);
  and g5947 (n5778, n5776, n5777);
  and g5948 (n5779, pi0221, n_29);
  not g5949 (n_2774, n5779);
  and g5950 (n5780, n_36, n_2774);
  not g5951 (n_2775, n5778);
  and g5952 (n5781, n_2775, n5780);
  not g5953 (n_2776, n5775);
  and g5954 (n5782, n_2776, n5781);
  not g5955 (n_2777, n5782);
  and g5956 (n5783, n_909, n_2777);
  not g5957 (n_2778, n5783);
  and g5958 (n5784, n_824, n_2778);
  and g5959 (n5785, n_826, n_2778);
  and g5960 (n5786, n_997, n_2768);
  and g5961 (n5787, n_263, n_207);
  not g5962 (n_2779, pi0846);
  and g5963 (n5788, n_2779, n2521);
  not g5964 (n_2780, n5787);
  and g5965 (n5789, n_188, n_2780);
  not g5966 (n_2781, n5788);
  and g5967 (n5790, n_2781, n5789);
  not g5968 (n_2782, n5790);
  and g5969 (n5791, n5786, n_2782);
  not g5970 (n_2783, n5791);
  and g5971 (n5792, n_20, n_2783);
  not g5972 (n_2784, n5792);
  and g5973 (n5793, n5766, n_2784);
  not g5974 (n_2785, n5793);
  and g5975 (n5794, n5781, n_2785);
  and g5976 (n5795, n3331, n5794);
  not g5977 (n_2786, n5785);
  and g5978 (n5796, pi0062, n_2786);
  not g5979 (n_2787, n5795);
  and g5980 (n5797, n_2787, n5796);
  not g5981 (n_2788, n5794);
  and g5982 (n5798, n2537, n_2788);
  and g5983 (n5799, n_179, n5783);
  not g5984 (n_2789, n5799);
  and g5985 (n5800, pi0056, n_2789);
  not g5986 (n_2790, n5798);
  and g5987 (n5801, n_2790, n5800);
  and g5988 (n5802, n_204, n_2778);
  and g5989 (n5803, n2572, n5794);
  not g5990 (n_2791, n5802);
  and g5991 (n5804, pi0055, n_2791);
  not g5992 (n_2792, n5803);
  and g5993 (n5805, n_2792, n5804);
  and g5994 (n5806, pi0224, pi0278);
  not g5995 (n_2793, n5806);
  and g5996 (n5807, n_226, n_2793);
  and g5997 (n5808, n_219, n5768);
  not g5998 (n_2794, n5808);
  and g5999 (n5809, n5807, n_2794);
  and g6000 (n5810, pi0222, n_219);
  and g6001 (n5811, n5776, n5810);
  not g6002 (n_2795, n5811);
  and g6003 (n5812, n2593, n_2795);
  not g6004 (n_2796, n5809);
  and g6005 (n5813, n_2796, n5812);
  not g6006 (n_2797, n5813);
  and g6007 (n5814, n_234, n_2797);
  and g6008 (n5815, n_1160, n5814);
  and g6009 (n5816, pi0299, n5783);
  not g6010 (n_2798, n5815);
  not g6011 (n_2799, n5816);
  and g6012 (n5817, n_2798, n_2799);
  and g6013 (n5818, n_841, n5817);
  and g6014 (n5819, n_251, n5817);
  and g6015 (n5820, pi0299, n_2788);
  not g6016 (n_2800, n5820);
  and g6017 (n5821, n_2798, n_2800);
  and g6018 (n5822, n2625, n5821);
  not g6019 (n_2801, n5819);
  not g6020 (n_2802, n5822);
  and g6021 (n5823, n_2801, n_2802);
  not g6022 (n_2803, n5823);
  and g6023 (n5824, n2533, n_2803);
  and g6024 (n5825, n_257, n5817);
  not g6025 (n_2804, n5825);
  and g6026 (n5826, pi0092, n_2804);
  not g6027 (n_2805, n5824);
  and g6028 (n5827, n_2805, n5826);
  and g6029 (n5828, pi0075, n5817);
  and g6030 (n5829, pi0087, n5823);
  and g6031 (n5830, pi0038, n5817);
  not g6032 (n_2806, n5821);
  and g6033 (n5831, pi0039, n_2806);
  and g6034 (n5832, n_2779, n3488);
  not g6035 (n_2807, n5832);
  and g6036 (n5833, n_219, n_2807);
  not g6037 (n_2808, n5833);
  and g6038 (n5834, n5807, n_2808);
  not g6039 (n_2809, n5834);
  and g6040 (n5835, n_2795, n_2809);
  and g6041 (n5836, n_224, n3470);
  and g6042 (n5837, n5835, n5836);
  and g6043 (n5838, pi0228, n_2765);
  and g6044 (n5839, pi0105, n_2807);
  not g6045 (n_2810, n5839);
  and g6046 (n5840, n5838, n_2810);
  not g6047 (n_2811, n5840);
  and g6048 (n5841, n_20, n_2811);
  and g6049 (n5842, n_263, n3499);
  and g6050 (n5843, pi0152, n_1174);
  not g6051 (n_2812, n5842);
  and g6052 (n5844, n_2779, n_2812);
  not g6053 (n_2813, n5843);
  and g6054 (n5845, n_2813, n5844);
  and g6055 (n5846, n_263, pi0846);
  and g6056 (n5847, n_879, n5846);
  not g6057 (n_2814, n5845);
  not g6058 (n_2815, n5847);
  and g6059 (n5848, n_2814, n_2815);
  not g6060 (n_2816, n5848);
  and g6061 (n5849, n_188, n_2816);
  not g6062 (n_2817, n5849);
  and g6063 (n5850, n5841, n_2817);
  not g6064 (n_2818, n5850);
  and g6065 (n5851, n5766, n_2818);
  not g6066 (n_2819, n5851);
  and g6067 (n5852, n_2775, n_2819);
  and g6068 (n5853, n_36, pi0299);
  and g6069 (n5854, n_2774, n5853);
  and g6070 (n5855, n5852, n5854);
  not g6071 (n_2820, n5837);
  and g6072 (n5856, n_162, n_2820);
  not g6073 (n_2821, n5855);
  and g6074 (n5857, n_2821, n5856);
  not g6075 (n_2822, n5831);
  and g6076 (n5858, n_161, n_2822);
  not g6077 (n_2823, n5857);
  and g6078 (n5859, n_2823, n5858);
  not g6079 (n_2824, n5830);
  and g6080 (n5860, n_164, n_2824);
  not g6081 (n_2825, n5859);
  and g6082 (n5861, n_2825, n5860);
  and g6083 (n5862, n_260, n5817);
  and g6084 (n5863, pi0846, n_863);
  not g6085 (n_2826, n5863);
  and g6086 (n5864, n_862, n_2826);
  not g6087 (n_2827, n5864);
  and g6088 (n5865, n_188, n_2827);
  not g6089 (n_2828, n5865);
  and g6090 (n5866, n5786, n_2828);
  not g6091 (n_2829, n5866);
  and g6092 (n5867, n_20, n_2829);
  not g6093 (n_2830, n5867);
  and g6094 (n5868, n5766, n_2830);
  not g6095 (n_2831, n5868);
  and g6096 (n5869, n5781, n_2831);
  not g6097 (n_2832, n5869);
  and g6098 (n5870, pi0299, n_2832);
  and g6099 (n5871, n2530, n_2798);
  not g6100 (n_2833, n5870);
  and g6101 (n5872, n_2833, n5871);
  not g6102 (n_2834, n5862);
  and g6103 (n5873, pi0100, n_2834);
  not g6104 (n_2835, n5872);
  and g6105 (n5874, n_2835, n5873);
  not g6106 (n_2836, n5861);
  not g6107 (n_2837, n5874);
  and g6108 (n5875, n_2836, n_2837);
  not g6109 (n_2838, n5875);
  and g6110 (n5876, n_172, n_2838);
  not g6111 (n_2839, n5829);
  and g6112 (n5877, n_171, n_2839);
  not g6113 (n_2840, n5876);
  and g6114 (n5878, n_2840, n5877);
  not g6115 (n_2841, n5828);
  and g6116 (n5879, n_174, n_2841);
  not g6117 (n_2842, n5878);
  and g6118 (n5880, n_2842, n5879);
  not g6119 (n_2843, n5827);
  and g6120 (n5881, n2532, n_2843);
  not g6121 (n_2844, n5880);
  and g6122 (n5882, n_2844, n5881);
  not g6123 (n_2845, n5818);
  and g6124 (n5883, n_176, n_2845);
  not g6125 (n_2846, n5882);
  and g6126 (n5884, n_2846, n5883);
  not g6127 (n_2847, n5805);
  and g6128 (n5885, n_157, n_2847);
  not g6129 (n_2848, n5884);
  and g6130 (n5886, n_2848, n5885);
  not g6131 (n_2849, n5801);
  and g6132 (n5887, n_158, n_2849);
  not g6133 (n_2850, n5886);
  and g6134 (n5888, n_2850, n5887);
  not g6135 (n_2851, n5797);
  and g6136 (n5889, n3328, n_2851);
  not g6137 (n_2852, n5888);
  and g6138 (n5890, n_2852, n5889);
  not g6139 (n_2854, n5784);
  and g6140 (n5891, pi0242, n_2854);
  not g6141 (n_2855, n5890);
  and g6142 (n5892, n_2855, n5891);
  and g6143 (n5893, n_824, n5782);
  and g6144 (n5894, n_826, n5782);
  and g6145 (n5895, n_2768, n_2782);
  not g6146 (n_2856, n5895);
  and g6147 (n5896, n_20, n_2856);
  not g6148 (n_2857, n5896);
  and g6149 (n5897, n5766, n_2857);
  not g6150 (n_2858, n5897);
  and g6151 (n5898, n5781, n_2858);
  and g6152 (n5899, n3331, n5898);
  not g6153 (n_2859, n5894);
  and g6154 (n5900, pi0062, n_2859);
  not g6155 (n_2860, n5899);
  and g6156 (n5901, n_2860, n5900);
  and g6157 (n5902, n_179, n_2777);
  not g6158 (n_2861, n5898);
  and g6159 (n5903, n2537, n_2861);
  not g6160 (n_2862, n5902);
  and g6161 (n5904, pi0056, n_2862);
  not g6162 (n_2863, n5903);
  and g6163 (n5905, n_2863, n5904);
  and g6164 (n5906, n_204, n5782);
  and g6165 (n5907, n2572, n5898);
  not g6166 (n_2864, n5906);
  and g6167 (n5908, pi0055, n_2864);
  not g6168 (n_2865, n5907);
  and g6169 (n5909, n_2865, n5908);
  and g6170 (n5910, pi0299, n_2777);
  not g6171 (n_2866, n5814);
  not g6172 (n_2867, n5910);
  and g6173 (n5911, n_2866, n_2867);
  and g6174 (n5912, n_841, n5911);
  and g6175 (n5913, n_251, n5911);
  and g6176 (n5914, pi0299, n_2861);
  not g6177 (n_2868, n5914);
  and g6178 (n5915, n_2866, n_2868);
  and g6179 (n5916, n2625, n5915);
  not g6180 (n_2869, n5913);
  not g6181 (n_2870, n5916);
  and g6182 (n5917, n_2869, n_2870);
  not g6183 (n_2871, n5917);
  and g6184 (n5918, n2533, n_2871);
  and g6185 (n5919, n_257, n5911);
  not g6186 (n_2872, n5919);
  and g6187 (n5920, pi0092, n_2872);
  not g6188 (n_2873, n5918);
  and g6189 (n5921, n_2873, n5920);
  and g6190 (n5922, pi0075, n5911);
  and g6191 (n5923, pi0087, n5917);
  and g6192 (n5924, pi0038, n5911);
  not g6193 (n_2874, n5915);
  and g6194 (n5925, pi0039, n_2874);
  and g6195 (n5926, n_929, n5808);
  not g6196 (n_2875, n5926);
  and g6197 (n5927, n5807, n_2875);
  and g6198 (n5928, n_2795, n5836);
  not g6199 (n_2876, n5927);
  and g6200 (n5929, n_2876, n5928);
  and g6201 (n5930, n_936, n5838);
  and g6202 (n5931, pi0152, n_2779);
  and g6203 (n5932, n_879, n5931);
  and g6204 (n5933, pi0152, n3499);
  and g6205 (n5934, n_263, n_1174);
  not g6206 (n_2877, n5933);
  and g6207 (n5935, pi0846, n_2877);
  not g6208 (n_2878, n5934);
  and g6209 (n5936, n_2878, n5935);
  not g6210 (n_2879, n5932);
  and g6211 (n5937, n_188, n_2879);
  not g6212 (n_2880, n5936);
  and g6213 (n5938, n_2880, n5937);
  not g6214 (n_2881, n5930);
  and g6215 (n5939, n5841, n_2881);
  not g6216 (n_2882, n5938);
  and g6217 (n5940, n_2882, n5939);
  not g6218 (n_2883, n5940);
  and g6219 (n5941, n5766, n_2883);
  not g6220 (n_2884, n5941);
  and g6221 (n5942, n_2775, n_2884);
  and g6222 (n5943, n5854, n5942);
  not g6223 (n_2885, n5929);
  and g6224 (n5944, n_162, n_2885);
  not g6225 (n_2886, n5943);
  and g6226 (n5945, n_2886, n5944);
  not g6227 (n_2887, n5925);
  and g6228 (n5946, n_161, n_2887);
  not g6229 (n_2888, n5945);
  and g6230 (n5947, n_2888, n5946);
  not g6231 (n_2889, n5924);
  and g6232 (n5948, n_164, n_2889);
  not g6233 (n_2890, n5947);
  and g6234 (n5949, n_2890, n5948);
  and g6235 (n5950, n_260, n5911);
  and g6236 (n5951, n_2768, n_2828);
  not g6237 (n_2891, n5951);
  and g6238 (n5952, n_20, n_2891);
  not g6239 (n_2892, n5952);
  and g6240 (n5953, n5766, n_2892);
  not g6241 (n_2893, n5953);
  and g6242 (n5954, n5781, n_2893);
  not g6243 (n_2894, n5954);
  and g6244 (n5955, pi0299, n_2894);
  and g6245 (n5956, n2530, n_2866);
  not g6246 (n_2895, n5955);
  and g6247 (n5957, n_2895, n5956);
  not g6248 (n_2896, n5950);
  and g6249 (n5958, pi0100, n_2896);
  not g6250 (n_2897, n5957);
  and g6251 (n5959, n_2897, n5958);
  not g6252 (n_2898, n5949);
  not g6253 (n_2899, n5959);
  and g6254 (n5960, n_2898, n_2899);
  not g6255 (n_2900, n5960);
  and g6256 (n5961, n_172, n_2900);
  not g6257 (n_2901, n5923);
  and g6258 (n5962, n_171, n_2901);
  not g6259 (n_2902, n5961);
  and g6260 (n5963, n_2902, n5962);
  not g6261 (n_2903, n5922);
  and g6262 (n5964, n_174, n_2903);
  not g6263 (n_2904, n5963);
  and g6264 (n5965, n_2904, n5964);
  not g6265 (n_2905, n5921);
  and g6266 (n5966, n2532, n_2905);
  not g6267 (n_2906, n5965);
  and g6268 (n5967, n_2906, n5966);
  not g6269 (n_2907, n5912);
  and g6270 (n5968, n_176, n_2907);
  not g6271 (n_2908, n5967);
  and g6272 (n5969, n_2908, n5968);
  not g6273 (n_2909, n5909);
  and g6274 (n5970, n_157, n_2909);
  not g6275 (n_2910, n5969);
  and g6276 (n5971, n_2910, n5970);
  not g6277 (n_2911, n5905);
  and g6278 (n5972, n_158, n_2911);
  not g6279 (n_2912, n5971);
  and g6280 (n5973, n_2912, n5972);
  not g6281 (n_2913, n5901);
  and g6282 (n5974, n3328, n_2913);
  not g6283 (n_2914, n5973);
  and g6284 (n5975, n_2914, n5974);
  not g6285 (n_2915, pi0242);
  not g6286 (n_2916, n5893);
  and g6287 (n5976, n_2915, n_2916);
  not g6288 (n_2917, n5975);
  and g6289 (n5977, n_2917, n5976);
  not g6290 (n_2918, n5892);
  not g6291 (n_2919, n5977);
  and g6292 (n5978, n_2918, n_2919);
  not g6293 (n_2921, pi1134);
  not g6294 (n_2922, n5978);
  and g6295 (n5979, n_2921, n_2922);
  and g6296 (n5980, n_2776, n_2775);
  not g6297 (n_2923, n5980);
  and g6298 (n5981, n_36, n_2923);
  and g6299 (n5982, n_824, n5981);
  and g6300 (n5983, n_826, n5981);
  and g6301 (n5984, n_2775, n_2858);
  not g6302 (n_2924, n5984);
  and g6303 (n5985, n_36, n_2924);
  and g6304 (n5986, n3331, n5985);
  not g6305 (n_2925, n5983);
  and g6306 (n5987, pi0062, n_2925);
  not g6307 (n_2926, n5986);
  and g6308 (n5988, n_2926, n5987);
  not g6309 (n_2927, n5981);
  and g6310 (n5989, n_179, n_2927);
  not g6311 (n_2928, n5985);
  and g6312 (n5990, n2537, n_2928);
  not g6313 (n_2929, n5989);
  and g6314 (n5991, pi0056, n_2929);
  not g6315 (n_2930, n5990);
  and g6316 (n5992, n_2930, n5991);
  and g6317 (n5993, n_204, n5981);
  and g6318 (n5994, n2572, n5985);
  not g6319 (n_2931, n5993);
  and g6320 (n5995, pi0055, n_2931);
  not g6321 (n_2932, n5994);
  and g6322 (n5996, n_2932, n5995);
  and g6323 (n5997, n2593, n5815);
  not g6324 (n_2933, n5997);
  and g6325 (n5998, n_234, n_2933);
  and g6326 (n5999, n_223, n5809);
  not g6327 (n_2934, n5999);
  and g6328 (n6000, n5998, n_2934);
  and g6329 (n6001, pi0299, n_2927);
  not g6330 (n_2935, n6000);
  not g6331 (n_2936, n6001);
  and g6332 (n6002, n_2935, n_2936);
  and g6333 (n6003, n_841, n6002);
  and g6334 (n6004, n_251, n6002);
  and g6335 (n6005, pi0299, n_2928);
  not g6336 (n_2937, n6005);
  and g6337 (n6006, n_2935, n_2937);
  and g6338 (n6007, n2625, n6006);
  not g6339 (n_2938, n6004);
  not g6340 (n_2939, n6007);
  and g6341 (n6008, n_2938, n_2939);
  not g6342 (n_2940, n6008);
  and g6343 (n6009, n2533, n_2940);
  and g6344 (n6010, n_257, n6002);
  not g6345 (n_2941, n6010);
  and g6346 (n6011, pi0092, n_2941);
  not g6347 (n_2942, n6009);
  and g6348 (n6012, n_2942, n6011);
  and g6349 (n6013, pi0075, n6002);
  and g6350 (n6014, pi0087, n6008);
  and g6351 (n6015, pi0038, n6002);
  not g6352 (n_2943, n6006);
  and g6353 (n6016, pi0039, n_2943);
  and g6354 (n6017, n3470, n5927);
  not g6355 (n_2944, n5942);
  and g6356 (n6018, n5853, n_2944);
  not g6357 (n_2945, n5835);
  and g6358 (n6019, n3470, n_2945);
  not g6359 (n_2946, n6019);
  and g6360 (n6020, n_162, n_2946);
  not g6361 (n_2947, n6017);
  and g6362 (n6021, n_2947, n6020);
  not g6363 (n_2948, n6018);
  and g6364 (n6022, n_2948, n6021);
  not g6365 (n_2949, n6016);
  and g6366 (n6023, n_161, n_2949);
  not g6367 (n_2950, n6022);
  and g6368 (n6024, n_2950, n6023);
  not g6369 (n_2951, n6015);
  and g6370 (n6025, n_164, n_2951);
  not g6371 (n_2952, n6024);
  and g6372 (n6026, n_2952, n6025);
  and g6373 (n6027, n_260, n6002);
  and g6374 (n6028, n_2775, n_2893);
  not g6375 (n_2953, n6028);
  and g6376 (n6029, n_36, n_2953);
  not g6377 (n_2954, n6029);
  and g6378 (n6030, pi0299, n_2954);
  and g6379 (n6031, n2530, n_2935);
  not g6380 (n_2955, n6030);
  and g6381 (n6032, n_2955, n6031);
  not g6382 (n_2956, n6027);
  and g6383 (n6033, pi0100, n_2956);
  not g6384 (n_2957, n6032);
  and g6385 (n6034, n_2957, n6033);
  not g6386 (n_2958, n6026);
  not g6387 (n_2959, n6034);
  and g6388 (n6035, n_2958, n_2959);
  not g6389 (n_2960, n6035);
  and g6390 (n6036, n_172, n_2960);
  not g6391 (n_2961, n6014);
  and g6392 (n6037, n_171, n_2961);
  not g6393 (n_2962, n6036);
  and g6394 (n6038, n_2962, n6037);
  not g6395 (n_2963, n6013);
  and g6396 (n6039, n_174, n_2963);
  not g6397 (n_2964, n6038);
  and g6398 (n6040, n_2964, n6039);
  not g6399 (n_2965, n6012);
  and g6400 (n6041, n2532, n_2965);
  not g6401 (n_2966, n6040);
  and g6402 (n6042, n_2966, n6041);
  not g6403 (n_2967, n6003);
  and g6404 (n6043, n_176, n_2967);
  not g6405 (n_2968, n6042);
  and g6406 (n6044, n_2968, n6043);
  not g6407 (n_2969, n5996);
  and g6408 (n6045, n_157, n_2969);
  not g6409 (n_2970, n6044);
  and g6410 (n6046, n_2970, n6045);
  not g6411 (n_2971, n5992);
  and g6412 (n6047, n_158, n_2971);
  not g6413 (n_2972, n6046);
  and g6414 (n6048, n_2972, n6047);
  not g6415 (n_2973, n5988);
  and g6416 (n6049, n3328, n_2973);
  not g6417 (n_2974, n6048);
  and g6418 (n6050, n_2974, n6049);
  not g6419 (n_2975, n5982);
  and g6420 (n6051, n_2915, n_2975);
  not g6421 (n_2976, n6050);
  and g6422 (n6052, n_2976, n6051);
  and g6423 (n6053, n_909, n5981);
  and g6424 (n6054, n_824, n6053);
  and g6425 (n6055, n_2775, n_2785);
  not g6426 (n_2977, n6055);
  and g6427 (n6056, n_36, n_2977);
  and g6428 (n6057, n3331, n6056);
  and g6429 (n6058, n_826, n6053);
  not g6430 (n_2978, n6058);
  and g6431 (n6059, pi0062, n_2978);
  not g6432 (n_2979, n6057);
  and g6433 (n6060, n_2979, n6059);
  not g6434 (n_2980, n6053);
  and g6435 (n6061, n_179, n_2980);
  not g6436 (n_2981, n6056);
  and g6437 (n6062, n2537, n_2981);
  not g6438 (n_2982, n6061);
  and g6439 (n6063, pi0056, n_2982);
  not g6440 (n_2983, n6062);
  and g6441 (n6064, n_2983, n6063);
  and g6442 (n6065, n2572, n6056);
  and g6443 (n6066, n_204, n6053);
  not g6444 (n_2984, n6066);
  and g6445 (n6067, pi0055, n_2984);
  not g6446 (n_2985, n6065);
  and g6447 (n6068, n_2985, n6067);
  and g6448 (n6069, pi0299, n_2980);
  not g6449 (n_2986, n5998);
  not g6450 (n_2987, n6069);
  and g6451 (n6070, n_2986, n_2987);
  and g6452 (n6071, n_841, n6070);
  and g6453 (n6072, n_251, n6070);
  and g6454 (n6073, pi0299, n_2981);
  not g6455 (n_2988, n6073);
  and g6456 (n6074, n_2986, n_2988);
  and g6457 (n6075, n2625, n6074);
  not g6458 (n_2989, n6072);
  not g6459 (n_2990, n6075);
  and g6460 (n6076, n_2989, n_2990);
  not g6461 (n_2991, n6076);
  and g6462 (n6077, n2533, n_2991);
  and g6463 (n6078, n_257, n6070);
  not g6464 (n_2992, n6078);
  and g6465 (n6079, pi0092, n_2992);
  not g6466 (n_2993, n6077);
  and g6467 (n6080, n_2993, n6079);
  and g6468 (n6081, pi0075, n6070);
  and g6469 (n6082, pi0087, n6076);
  and g6470 (n6083, pi0038, n6070);
  not g6471 (n_2994, n6074);
  and g6472 (n6084, pi0039, n_2994);
  not g6473 (n_2995, n5852);
  and g6474 (n6085, n_2995, n5853);
  not g6475 (n_2996, n6085);
  and g6476 (n6086, n6020, n_2996);
  not g6477 (n_2997, n6084);
  and g6478 (n6087, n_161, n_2997);
  not g6479 (n_2998, n6086);
  and g6480 (n6088, n_2998, n6087);
  not g6481 (n_2999, n6083);
  and g6482 (n6089, n_164, n_2999);
  not g6483 (n_3000, n6088);
  and g6484 (n6090, n_3000, n6089);
  and g6485 (n6091, n_260, n6070);
  and g6486 (n6092, n_2775, n_2831);
  not g6487 (n_3001, n6092);
  and g6488 (n6093, n_36, n_3001);
  not g6489 (n_3002, n6093);
  and g6490 (n6094, pi0299, n_3002);
  and g6491 (n6095, n2530, n_2986);
  not g6492 (n_3003, n6094);
  and g6493 (n6096, n_3003, n6095);
  not g6494 (n_3004, n6091);
  and g6495 (n6097, pi0100, n_3004);
  not g6496 (n_3005, n6096);
  and g6497 (n6098, n_3005, n6097);
  not g6498 (n_3006, n6090);
  not g6499 (n_3007, n6098);
  and g6500 (n6099, n_3006, n_3007);
  not g6501 (n_3008, n6099);
  and g6502 (n6100, n_172, n_3008);
  not g6503 (n_3009, n6082);
  and g6504 (n6101, n_171, n_3009);
  not g6505 (n_3010, n6100);
  and g6506 (n6102, n_3010, n6101);
  not g6507 (n_3011, n6081);
  and g6508 (n6103, n_174, n_3011);
  not g6509 (n_3012, n6102);
  and g6510 (n6104, n_3012, n6103);
  not g6511 (n_3013, n6080);
  and g6512 (n6105, n2532, n_3013);
  not g6513 (n_3014, n6104);
  and g6514 (n6106, n_3014, n6105);
  not g6515 (n_3015, n6071);
  and g6516 (n6107, n_176, n_3015);
  not g6517 (n_3016, n6106);
  and g6518 (n6108, n_3016, n6107);
  not g6519 (n_3017, n6068);
  and g6520 (n6109, n_157, n_3017);
  not g6521 (n_3018, n6108);
  and g6522 (n6110, n_3018, n6109);
  not g6523 (n_3019, n6064);
  and g6524 (n6111, n_158, n_3019);
  not g6525 (n_3020, n6110);
  and g6526 (n6112, n_3020, n6111);
  not g6527 (n_3021, n6060);
  and g6528 (n6113, n3328, n_3021);
  not g6529 (n_3022, n6112);
  and g6530 (n6114, n_3022, n6113);
  not g6531 (n_3023, n6054);
  and g6532 (n6115, pi0242, n_3023);
  not g6533 (n_3024, n6114);
  and g6534 (n6116, n_3024, n6115);
  not g6535 (n_3025, n6052);
  and g6536 (n6117, pi1134, n_3025);
  not g6537 (n_3026, n6116);
  and g6538 (n6118, n_3026, n6117);
  not g6539 (n_3027, n5979);
  not g6540 (n_3028, n6118);
  and g6541 (po0165, n_3027, n_3028);
  and g6542 (n6120, pi0057, pi0059);
  and g6543 (n6121, n2521, n2538);
  not g6544 (n_3029, n6121);
  and g6545 (n6122, n_824, n_3029);
  not g6546 (n_3030, n6120);
  not g6547 (n_3031, n6122);
  and g6548 (n6123, n_3030, n_3031);
  not g6549 (n_3032, n6123);
  and g6550 (n6124, pi0057, n_3032);
  and g6551 (n6125, n2512, n2625);
  and g6552 (n6126, n2536, n6125);
  not g6553 (n_3033, n6126);
  and g6554 (n6127, pi0056, n_3033);
  and g6555 (n6128, n_167, n2534);
  and g6556 (n6129, n6125, n6128);
  not g6557 (n_3034, n6129);
  and g6558 (n6130, pi0074, n_3034);
  not g6559 (n_3035, n6130);
  and g6560 (n6131, n_176, n_3035);
  not g6561 (n_3036, n6125);
  and g6562 (n6132, pi0087, n_3036);
  not g6563 (n_3037, n6132);
  and g6564 (n6133, n_171, n_3037);
  and g6565 (n6134, n_167, n_174);
  and g6566 (n6135, n_162, n2512);
  not g6567 (n_3038, n6135);
  and g6568 (n6136, pi0038, n_3038);
  not g6569 (n_3039, n6136);
  and g6570 (n6137, n_164, n_3039);
  and g6571 (n6138, pi0058, n2502);
  not g6572 (n_3040, n6138);
  and g6573 (n6139, n_43, n_3040);
  and g6574 (n6140, n2720, n2769);
  and g6575 (n6141, n2874, n6140);
  not g6576 (n_3041, n6141);
  and g6577 (n6142, n2781, n_3041);
  not g6578 (n_3042, n6142);
  and g6579 (n6143, n_453, n_3042);
  not g6580 (n_3043, n6143);
  and g6581 (n6144, n_123, n_3043);
  not g6582 (n_3044, n6144);
  and g6583 (n6145, n2775, n_3044);
  and g6584 (n6146, n_113, n2889);
  not g6585 (n_3045, n6145);
  and g6586 (n6147, n_3045, n6146);
  and g6587 (n6148, n_357, n_459);
  not g6588 (n_3046, n6147);
  and g6589 (n6149, n_3046, n6148);
  not g6590 (n_3047, n6149);
  and g6591 (n6150, n_108, n_3047);
  and g6592 (n6151, n2700, n_356);
  not g6593 (n_3048, n6150);
  and g6594 (n6152, n_3048, n6151);
  not g6595 (n_3049, n6152);
  and g6596 (n6153, n6139, n_3049);
  not g6597 (n_3050, n6153);
  and g6598 (n6154, n_466, n_3050);
  not g6599 (n_3051, n6154);
  and g6600 (n6155, n_131, n_3051);
  not g6601 (n_3052, pi0841);
  and g6602 (n6156, n_3052, n2503);
  not g6603 (n_3053, n6156);
  and g6604 (n6157, pi0093, n_3053);
  not g6605 (n_3054, n6155);
  not g6606 (n_3055, n6157);
  and g6607 (n6158, n_3054, n_3055);
  not g6608 (n_3056, n6158);
  and g6609 (n6159, n_130, n_3056);
  and g6610 (n6160, n_139, n_339);
  not g6611 (n_3057, n6159);
  and g6612 (n6161, n_3057, n6160);
  not g6613 (n_3058, n6161);
  and g6614 (n6162, n_138, n_3058);
  not g6615 (n_3059, n6162);
  and g6616 (n6163, n2748, n_3059);
  not g6617 (n_3060, n6163);
  and g6618 (n6164, n3168, n_3060);
  not g6619 (n_3061, n6164);
  and g6620 (n6165, n2746, n_3061);
  not g6621 (n_3062, n6165);
  and g6622 (n6166, n2744, n_3062);
  and g6623 (n6167, n_305, n_234);
  and g6624 (n6168, n_271, pi0299);
  not g6625 (n_3063, n6167);
  not g6626 (n_3064, n6168);
  and g6627 (n6169, n_3063, n_3064);
  and g6628 (n6170, n_130, n2508);
  and g6629 (n6171, n_143, n6170);
  and g6630 (n6172, n2915, n6171);
  not g6631 (n_3065, n6172);
  and g6632 (n6173, pi0032, n_3065);
  not g6633 (n_3066, n6169);
  not g6634 (n_3067, n6173);
  and g6635 (n6174, n_3066, n_3067);
  and g6636 (n6175, n_875, n6169);
  not g6637 (n_3068, n6174);
  not g6638 (n_3069, n6175);
  and g6639 (n6176, n_3068, n_3069);
  not g6640 (n_3070, n6166);
  not g6641 (n_3071, n6176);
  and g6642 (n6177, n_3070, n_3071);
  not g6643 (n_3072, n6177);
  and g6644 (n6178, n_144, n_3072);
  not g6645 (n_3073, n6178);
  and g6646 (n6179, n_345, n_3073);
  not g6647 (n_3074, n6179);
  and g6648 (n6180, n_162, n_3074);
  and g6649 (n6181, pi0835, pi0984);
  not g6650 (n_3078, pi1001);
  and g6651 (n6182, n_280, n_3078);
  not g6652 (n_3080, pi0979);
  not g6653 (n_3081, n6182);
  and g6654 (n6183, n_3080, n_3081);
  not g6655 (n_3082, n6181);
  and g6656 (n6184, n_3082, n6183);
  not g6657 (n_3084, pi0287);
  and g6658 (n6185, n_3084, n6184);
  and g6659 (n6186, pi0835, pi0950);
  and g6660 (n6187, n6185, n6186);
  and g6661 (n6188, n2928, n6187);
  and g6662 (n6189, pi0222, pi0224);
  not g6663 (n_3087, pi0642);
  and g6664 (n6190, pi0603, n_3087);
  not g6665 (n_3090, pi0614);
  not g6666 (n_3091, pi0616);
  and g6667 (n6191, n_3090, n_3091);
  and g6668 (n6192, n6190, n6191);
  not g6669 (n_3093, pi0662);
  and g6670 (n6193, n_3093, pi0680);
  not g6671 (n_3096, pi0661);
  and g6672 (n6194, n_3096, n6193);
  not g6673 (n_3098, pi0681);
  and g6674 (n6195, n_3098, n6194);
  or g6675 (po1101, n6192, n6195);
  not g6676 (n_3100, pi0468);
  and g6677 (n6197, n_4, n_3100);
  not g6678 (n_3102, n6197);
  and g6679 (n6198, po1101, n_3102);
  not g6680 (n_3105, pi0587);
  not g6681 (n_3106, pi0602);
  not g6695 (n_3119, n6205);
  and g6696 (n6206, n6197, n_3119);
  not g6697 (n_3120, n6198);
  not g6698 (n_3121, n6206);
  and g6699 (n6207, n_3120, n_3121);
  and g6700 (n6208, n6188, n6189);
  not g6701 (n_3122, n6207);
  and g6702 (n6209, n_3122, n6208);
  not g6703 (n_3123, n6209);
  and g6704 (n6210, n2521, n_3123);
  not g6705 (n_3124, n6210);
  and g6706 (n6211, n_223, n_3124);
  and g6707 (n6212, pi1092, n6187);
  not g6708 (n_3126, pi0824);
  not g6709 (n_3127, pi0829);
  and g6710 (n6213, n_3126, n_3127);
  not g6711 (n_3128, pi1091);
  and g6712 (n6214, pi0824, n_3128);
  and g6713 (n6215, pi1093, n_538);
  not g6714 (n_3129, n6214);
  and g6715 (n6216, n_3129, n6215);
  not g6716 (n_3130, n6213);
  not g6717 (n_3131, n6216);
  and g6718 (n6217, n_3130, n_3131);
  and g6719 (n6218, n6212, n6217);
  not g6720 (n_3132, n6218);
  and g6721 (n6219, n_3102, n_3132);
  not g6722 (n_3133, n6219);
  and g6723 (n6220, po1101, n_3133);
  not g6724 (n_3134, n6220);
  and g6725 (n6221, n2521, n_3134);
  and g6726 (n6222, n2512, n6197);
  and g6727 (n6223, po1101, n6222);
  not g6728 (n_3135, n6221);
  not g6729 (n_3136, n6223);
  and g6730 (n6224, n_3135, n_3136);
  not g6731 (n_3137, n6224);
  and g6732 (n6225, n6205, n_3137);
  not g6733 (n_3138, n6192);
  and g6734 (n6226, n_3138, n_3102);
  not g6735 (n_3139, n6195);
  and g6736 (n6227, n_3139, n6226);
  not g6737 (n_3140, n6227);
  and g6738 (n6228, n6218, n_3140);
  not g6739 (n_3141, n6228);
  and g6740 (n6229, n2521, n_3141);
  and g6741 (n6230, n_3119, n6229);
  not g6742 (n_3142, n6230);
  and g6743 (n6231, pi0223, n_3142);
  not g6744 (n_3143, n6225);
  and g6745 (n6232, n_3143, n6231);
  not g6746 (n_3144, n6211);
  and g6747 (n6233, n_234, n_3144);
  not g6748 (n_3145, n6232);
  and g6749 (n6234, n_3145, n6233);
  and g6750 (n6235, pi0216, pi0221);
  not g6751 (n_3148, pi0907);
  not g6752 (n_3149, pi0947);
  and g6753 (n6236, n_3148, n_3149);
  and g6765 (n6242, n6236, n6241);
  not g6766 (n_3162, n6242);
  and g6767 (n6243, n6197, n_3162);
  not g6768 (n_3163, n6243);
  and g6769 (n6244, n_3120, n_3163);
  and g6770 (n6245, n6188, n6235);
  not g6771 (n_3164, n6244);
  and g6772 (n6246, n_3164, n6245);
  not g6773 (n_3165, n6246);
  and g6774 (n6247, n2521, n_3165);
  not g6775 (n_3166, n6247);
  and g6776 (n6248, n_36, n_3166);
  and g6777 (n6249, n6229, n_3162);
  and g6778 (n6250, n_3137, n6242);
  not g6779 (n_3167, n6249);
  and g6780 (n6251, pi0215, n_3167);
  not g6781 (n_3168, n6250);
  and g6782 (n6252, n_3168, n6251);
  not g6783 (n_3169, n6248);
  and g6784 (n6253, pi0299, n_3169);
  not g6785 (n_3170, n6252);
  and g6786 (n6254, n_3170, n6253);
  not g6787 (n_3171, n6234);
  and g6788 (n6255, pi0039, n_3171);
  not g6789 (n_3172, n6254);
  and g6790 (n6256, n_3172, n6255);
  not g6791 (n_3173, n6180);
  not g6792 (n_3174, n6256);
  and g6793 (n6257, n_3173, n_3174);
  not g6794 (n_3175, n6257);
  and g6795 (n6258, n_161, n_3175);
  not g6796 (n_3176, n6258);
  and g6797 (n6259, n6137, n_3176);
  and g6798 (n6260, n_738, n_302);
  and g6799 (n6261, n_234, n6260);
  and g6800 (n6262, pi0299, n2640);
  not g6801 (n_3177, n6261);
  not g6802 (n_3178, n6262);
  and g6803 (n6263, n_3177, n_3178);
  and g6804 (n6264, n_855, n6263);
  not g6805 (n_3181, pi0041);
  not g6806 (n_3182, pi0099);
  and g6807 (n6265, n_3181, n_3182);
  not g6808 (n_3184, pi0101);
  and g6809 (n6266, n_3184, n6265);
  not g6810 (n_3187, pi0042);
  not g6811 (n_3188, pi0043);
  and g6812 (n6267, n_3187, n_3188);
  not g6813 (n_3190, pi0052);
  and g6814 (n6268, n_3190, n6267);
  not g6815 (n_3193, pi0113);
  not g6816 (n_3194, pi0116);
  and g6817 (n6269, n_3193, n_3194);
  not g6818 (n_3197, pi0114);
  not g6819 (n_3198, pi0115);
  and g6820 (n6270, n_3197, n_3198);
  and g6821 (n6271, n6269, n6270);
  and g6822 (n6272, n6268, n6271);
  and g6823 (n6273, n6266, n6272);
  not g6824 (n_3200, n6273);
  or g6825 (po1057, pi0044, n_3200);
  not g6826 (n_3202, pi0683);
  and g6827 (n6275, n_3202, po1057);
  and g6828 (n6276, pi0129, pi0250);
  and g6829 (n6277, n2932, n_3130);
  not g6830 (n_3206, pi1093);
  and g6831 (po0740, n_3206, n6277);
  not g6832 (n_3208, pi0250);
  not g6833 (n_3209, po0740);
  and g6834 (n6279, n_3208, n_3209);
  not g6835 (n_3210, n6276);
  not g6836 (n_3211, n6279);
  and g6837 (n6280, n_3210, n_3211);
  not g6838 (n_3212, n6275);
  not g6839 (n_3213, n6280);
  and g6840 (n6281, n_3212, n_3213);
  not g6841 (n_3214, n6263);
  and g6842 (n6282, n_3214, po1057);
  and g6843 (n6283, n6281, n6282);
  and g6844 (n6284, n_162, n2521);
  and g6845 (n6285, n_161, pi0100);
  and g6846 (n6286, n6284, n6285);
  not g6847 (n_3215, n6264);
  not g6848 (n_3216, n6283);
  and g6849 (n6287, n_3215, n_3216);
  and g6850 (n6288, n6286, n6287);
  not g6851 (n_3217, n6288);
  and g6852 (n6289, n_172, n_3217);
  not g6853 (n_3218, n6259);
  and g6854 (n6290, n_3218, n6289);
  and g6855 (n6291, n6133, n6134);
  not g6856 (n_3219, n6290);
  and g6857 (n6292, n_3219, n6291);
  not g6858 (n_3220, n6292);
  and g6859 (n6293, n_168, n_3220);
  not g6860 (n_3221, n6293);
  and g6861 (n6294, n6131, n_3221);
  not g6862 (n_3222, n6294);
  and g6863 (n6295, n_157, n_3222);
  not g6864 (n_3223, n6127);
  not g6865 (n_3224, n6295);
  and g6866 (n6296, n_3223, n_3224);
  not g6867 (n_3225, n6296);
  and g6868 (n6297, n_158, n_3225);
  and g6869 (n6298, n3330, n6125);
  not g6870 (n_3226, n6298);
  and g6871 (n6299, pi0062, n_3226);
  not g6872 (n_3227, n6299);
  and g6873 (n6300, n_792, n_3227);
  not g6874 (n_3228, n6297);
  and g6875 (n6301, n_3228, n6300);
  not g6876 (n_3229, n6301);
  and g6877 (n6302, n_796, n_3229);
  not g6878 (n_3230, n6124);
  not g6879 (n_3231, n6302);
  and g6880 (po0167, n_3230, n_3231);
  and g6881 (n6304, n_176, n2529);
  and g6882 (n6305, n_792, n6304);
  not g6883 (n_3232, n6305);
  and g6884 (n6306, n_188, n_3232);
  not g6885 (n_3233, n6306);
  and g6886 (n6307, pi0057, n_3233);
  and g6887 (n6308, n_3139, n_3102);
  and g6888 (n6309, n_3148, n6197);
  not g6889 (n_3234, n6308);
  not g6890 (n_3235, n6309);
  and g6891 (n6310, n_3234, n_3235);
  and g6892 (n6311, n_188, n_204);
  and g6893 (n6312, pi0030, pi0228);
  not g6894 (n_3237, n6312);
  and g6895 (n6313, n_1324, n_3237);
  not g6896 (n_3238, n6311);
  not g6897 (n_3239, n6313);
  and g6898 (n6314, n_3238, n_3239);
  and g6899 (n6315, n6310, n6314);
  and g6900 (n6316, n6307, n6315);
  not g6901 (n_3240, n6304);
  and g6902 (n6317, n_188, n_3240);
  not g6903 (n_3241, n6317);
  and g6904 (n6318, n6315, n_3241);
  not g6905 (n_3242, n6318);
  and g6906 (n6319, pi0059, n_3242);
  and g6907 (n6320, n6310, n6312);
  not g6908 (n_3243, n2529);
  and g6909 (n6321, n_3243, n6320);
  not g6910 (n_3244, n6315);
  and g6911 (n6322, pi0055, n_3244);
  and g6912 (n6323, n_167, n2569);
  and g6913 (n6324, pi0299, n6310);
  and g6914 (n6325, n_3106, n6197);
  not g6915 (n_3245, n6325);
  and g6916 (n6326, n_3234, n_3245);
  and g6917 (n6327, n_234, n6326);
  not g6918 (n_3246, n6324);
  not g6919 (n_3247, n6327);
  and g6920 (n6328, n_3246, n_3247);
  not g6921 (n_3248, n6328);
  and g6922 (n6329, n6312, n_3248);
  not g6923 (n_3249, n6323);
  not g6924 (n_3250, n6329);
  and g6925 (n6330, n_3249, n_3250);
  and g6926 (n6331, n_766, n6329);
  and g6927 (n6332, n_162, n_3239);
  and g6928 (n6333, n_3248, n6332);
  and g6929 (n6334, n2620, n6333);
  not g6930 (n_3251, n6331);
  not g6931 (n_3252, n6334);
  and g6932 (n6335, n_3251, n_3252);
  and g6933 (n6336, n2569, n6335);
  and g6934 (n6337, n_167, n6336);
  not g6935 (n_3253, n6330);
  and g6936 (n6338, pi0074, n_3253);
  not g6937 (n_3254, n6337);
  and g6938 (n6339, n_3254, n6338);
  not g6939 (n_3255, n2569);
  and g6940 (n6340, n_3255, n_3250);
  not g6941 (n_3256, n6336);
  not g6942 (n_3257, n6340);
  and g6943 (n6341, n_3256, n_3257);
  not g6944 (n_3258, n6341);
  and g6945 (n6342, pi0054, n_3258);
  and g6946 (n6343, n_171, n6335);
  and g6947 (n6344, pi0075, n_3250);
  not g6948 (n_3259, n6344);
  and g6949 (n6345, pi0092, n_3259);
  not g6950 (n_3260, n6343);
  and g6951 (n6346, n_3260, n6345);
  and g6952 (n6347, pi0075, n6335);
  and g6953 (n6348, pi0087, n6329);
  and g6954 (n6349, n_260, n6329);
  and g6955 (n6350, n6312, n6326);
  and g6956 (n6351, n2521, n_3213);
  and g6957 (n6352, pi0683, po1057);
  and g6958 (n6353, n6351, n6352);
  and g6959 (n6354, n_3234, n6353);
  and g6960 (n6355, n6260, n6354);
  not g6961 (n_3261, n6260);
  and g6962 (n6356, pi0252, n_3261);
  and g6963 (n6357, pi0252, n6222);
  and g6964 (n6358, n_3139, n6357);
  and g6965 (n6359, pi0252, n2521);
  and g6966 (n6360, n6195, n6359);
  not g6967 (n_3262, n6358);
  not g6968 (n_3263, n6360);
  and g6969 (n6361, n_3262, n_3263);
  not g6970 (n_3264, n6361);
  and g6971 (n6362, n6356, n_3264);
  not g6972 (n_3265, n6355);
  not g6973 (n_3266, n6362);
  and g6974 (n6363, n_3265, n_3266);
  and g6975 (n6364, n_188, n_3245);
  not g6976 (n_3267, n6363);
  and g6977 (n6365, n_3267, n6364);
  not g6978 (n_3268, n6350);
  and g6979 (n6366, n_234, n_3268);
  not g6980 (n_3269, n6365);
  and g6981 (n6367, n_3269, n6366);
  not g6982 (n_3270, n6320);
  and g6983 (n6368, pi0299, n_3270);
  not g6984 (n_3271, n6354);
  and g6985 (n6369, n2640, n_3271);
  and g6986 (n6370, n_272, n6361);
  not g6992 (n_3274, n6373);
  and g6993 (n6374, n6368, n_3274);
  not g6994 (n_3275, n6374);
  and g6995 (n6375, n2530, n_3275);
  not g6996 (n_3276, n6367);
  and g6997 (n6376, n_3276, n6375);
  not g6998 (n_3277, n6349);
  and g6999 (n6377, pi0100, n_3277);
  not g7000 (n_3278, n6376);
  and g7001 (n6378, n_3278, n6377);
  and g7002 (n6379, n_36, pi0221);
  and g7003 (n6380, n_3084, n2521);
  and g7004 (n6381, pi0835, n6184);
  and g7005 (n6382, n6380, n6381);
  and g7006 (n6383, pi0824, pi1093);
  and g7007 (n6384, n2932, n6383);
  and g7008 (n6385, n6382, n6384);
  and g7009 (n6386, n_3128, n6385);
  and g7010 (n6387, pi1091, n2923);
  not g7011 (n_3279, n6387);
  and g7012 (n6388, n6384, n_3279);
  not g7013 (n_3280, n6388);
  and g7014 (n6389, n_494, n_3280);
  not g7015 (n_3281, n6389);
  and g7016 (n6390, pi1091, n_3281);
  and g7017 (n6391, n6382, n6390);
  not g7018 (n_3282, n6386);
  not g7019 (n_3283, n6391);
  and g7020 (n6392, n_3282, n_3283);
  not g7021 (n_3284, n6392);
  and g7022 (n6393, pi0216, n_3284);
  and g7023 (n6394, n_3127, n_489);
  not g7024 (n_3285, n6394);
  and g7025 (n6395, pi1091, n_3285);
  not g7026 (n_3286, n6395);
  and g7027 (n6396, n6385, n_3286);
  and g7028 (n6397, n_20, n6396);
  not g7029 (n_3287, n6393);
  not g7030 (n_3288, n6397);
  and g7031 (n6398, n_3287, n_3288);
  not g7032 (n_3289, n6398);
  and g7033 (n6399, n_188, n_3289);
  not g7034 (n_3290, n6399);
  and g7035 (n6400, n_3237, n_3290);
  not g7036 (n_3291, n6400);
  and g7037 (n6401, n6379, n_3291);
  not g7038 (n_3292, n6401);
  and g7039 (n6402, n_3237, n_3292);
  not g7040 (n_3293, n6402);
  and g7041 (n6403, n6310, n_3293);
  not g7042 (n_3294, n6403);
  and g7043 (n6404, pi0299, n_3294);
  and g7044 (n6405, pi0222, n_223);
  not g7045 (n_3295, n6396);
  and g7046 (n6406, n_219, n_3295);
  and g7047 (n6407, pi0224, n6392);
  not g7048 (n_3296, n6406);
  and g7049 (n6408, n6405, n_3296);
  not g7050 (n_3297, n6407);
  and g7051 (n6409, n_3297, n6408);
  and g7052 (n6410, n_188, n6409);
  not g7053 (n_3298, n6410);
  and g7054 (n6411, n_3237, n_3298);
  not g7055 (n_3299, n6411);
  and g7056 (n6412, n6326, n_3299);
  not g7057 (n_3300, n6412);
  and g7058 (n6413, n_234, n_3300);
  not g7059 (n_3301, n6413);
  and g7060 (n6414, pi0039, n_3301);
  not g7061 (n_3302, n6404);
  and g7062 (n6415, n_3302, n6414);
  and g7063 (n6416, pi0158, pi0159);
  and g7064 (n6417, pi0160, pi0197);
  and g7065 (n6418, n6416, n6417);
  not g7066 (n_3307, n2755);
  and g7067 (n6419, pi0091, n_3307);
  not g7068 (n_3308, n6419);
  and g7069 (n6420, n_42, n_3308);
  not g7070 (n_3310, pi0314);
  and g7071 (n6421, n_109, n_3310);
  and g7072 (n6422, n2765, n_459);
  and g7073 (n6423, pi0067, n2483);
  and g7074 (n6424, pi0085, n2827);
  not g7075 (n_3311, n6424);
  and g7076 (n6425, n2469, n_3311);
  not g7077 (n_3312, n6425);
  and g7078 (n6426, n2831, n_3312);
  not g7079 (n_3313, n6426);
  and g7080 (n6427, n2478, n_3313);
  and g7081 (n6428, n_411, n_408);
  not g7082 (n_3314, n6427);
  and g7083 (n6429, n_3314, n6428);
  and g7084 (n6430, n2479, n6429);
  not g7085 (n_3315, n6430);
  and g7086 (n6431, n_413, n_3315);
  not g7087 (n_3316, n6431);
  and g7088 (n6432, n2804, n_3316);
  not g7089 (n_3317, n6423);
  and g7090 (n6433, n2797, n_3317);
  not g7091 (n_3318, n6432);
  and g7092 (n6434, n_3318, n6433);
  not g7093 (n_3319, n6434);
  and g7094 (n6435, n2796, n_3319);
  not g7095 (n_3320, n6435);
  and g7096 (n6436, n_57, n_3320);
  not g7097 (n_3321, n2487);
  or g7098 (po1049, pi0064, n_3321);
  not g7099 (n_3323, po1049);
  and g7100 (n6438, n2791, n_3323);
  not g7101 (n_3324, n6436);
  and g7102 (n6439, n_3324, n6438);
  not g7103 (n_3325, n6439);
  and g7104 (n6440, n_105, n_3325);
  and g7105 (n6441, n2845, n6438);
  not g7106 (n_3326, n6441);
  and g7107 (n6442, n6440, n_3326);
  and g7108 (n6443, n_53, n_368);
  and g7109 (n6444, n2463, n6443);
  not g7110 (n_3327, n6442);
  and g7111 (n6445, n_3327, n6444);
  not g7112 (n_3328, n6445);
  and g7113 (n6446, n2785, n_3328);
  not g7114 (n_3329, n6446);
  and g7115 (n6447, n2877, n_3329);
  not g7116 (n_3330, n6447);
  and g7117 (n6448, n2719, n_3330);
  not g7118 (n_3331, n6448);
  and g7119 (n6449, n_333, n_3331);
  not g7120 (n_3332, n6449);
  and g7121 (n6450, n_119, n_3332);
  and g7122 (n6451, n_127, n2496);
  and g7123 (n6452, n2783, n6451);
  not g7124 (n_3333, n6450);
  and g7125 (n6453, n_3333, n6452);
  not g7126 (n_3334, n6453);
  and g7127 (n6454, n2889, n_3334);
  not g7128 (n_3335, n6454);
  and g7129 (n6455, n6422, n_3335);
  not g7130 (n_3336, n6455);
  and g7131 (n6456, n6421, n_3336);
  and g7132 (n6457, n_109, pi0314);
  not g7133 (n_3337, n6440);
  and g7134 (n6458, n_3337, n6444);
  not g7135 (n_3338, n6458);
  and g7136 (n6459, n2785, n_3338);
  not g7137 (n_3339, n6459);
  and g7138 (n6460, n2877, n_3339);
  not g7139 (n_3340, n6460);
  and g7140 (n6461, n2719, n_3340);
  not g7141 (n_3341, n6461);
  and g7142 (n6462, n_333, n_3341);
  not g7143 (n_3342, n6462);
  and g7144 (n6463, n_119, n_3342);
  not g7145 (n_3343, n6463);
  and g7146 (n6464, n6452, n_3343);
  not g7147 (n_3344, n6464);
  and g7148 (n6465, n2889, n_3344);
  not g7149 (n_3345, n6465);
  and g7150 (n6466, n6422, n_3345);
  not g7151 (n_3346, n6466);
  and g7152 (n6467, n6457, n_3346);
  not g7153 (n_3347, n6467);
  and g7154 (n6468, n6420, n_3347);
  not g7155 (n_3348, n6456);
  and g7156 (n6469, n_3348, n6468);
  not g7157 (n_3349, n6469);
  and g7158 (n6470, n_43, n_3349);
  not g7159 (n_3350, n6470);
  and g7160 (n6471, n_466, n_3350);
  not g7161 (n_3351, n6471);
  and g7162 (n6472, n_131, n_3351);
  not g7163 (n_3352, n2914);
  and g7164 (n6473, pi0093, n_3352);
  not g7165 (n_3353, n6473);
  and g7166 (n6474, n_130, n_3353);
  not g7167 (n_3354, n6472);
  and g7168 (n6475, n_3354, n6474);
  not g7169 (n_3355, n6475);
  and g7170 (n6476, n_139, n_3355);
  not g7171 (n_3356, n6476);
  and g7172 (n6477, n3100, n_3356);
  not g7173 (n_3357, n6477);
  and g7174 (n6478, n_134, n_3357);
  and g7175 (n6479, n_144, n2510);
  and g7176 (n6480, n_348, n6479);
  not g7177 (n_3358, n6478);
  and g7178 (n6481, n_3358, n6480);
  not g7179 (n_3359, n6481);
  and g7180 (n6482, n_692, n_3359);
  and g7181 (n6483, n_3052, n2728);
  and g7182 (n6484, n2962, n6483);
  and g7183 (n6485, n2736, n6484);
  and g7184 (n6486, pi0032, n6485);
  and g7185 (n6487, n_144, n6486);
  and g7186 (n6488, n_271, n6487);
  not g7187 (n_3360, n6488);
  and g7188 (n6489, n6482, n_3360);
  not g7189 (n_3361, n6489);
  and g7190 (n6490, n_3102, n_3361);
  and g7191 (n6491, n_108, n2493);
  and g7192 (n6492, n_457, n_3334);
  not g7193 (n_3362, n6492);
  and g7194 (n6493, n6491, n_3362);
  not g7195 (n_3363, n6493);
  and g7196 (n6494, n6421, n_3363);
  and g7197 (n6495, n_457, n_3344);
  not g7198 (n_3364, n6495);
  and g7199 (n6496, n6491, n_3364);
  not g7200 (n_3365, n6496);
  and g7201 (n6497, n6457, n_3365);
  not g7202 (n_3366, n6497);
  and g7203 (n6498, n6420, n_3366);
  not g7204 (n_3367, n6494);
  and g7205 (n6499, n_3367, n6498);
  not g7206 (n_3368, n6499);
  and g7207 (n6500, n_43, n_3368);
  not g7208 (n_3369, n6500);
  and g7209 (n6501, n_466, n_3369);
  not g7210 (n_3370, n6501);
  and g7211 (n6502, n_131, n_3370);
  not g7212 (n_3371, n6502);
  and g7213 (n6503, n6474, n_3371);
  not g7214 (n_3372, n6503);
  and g7215 (n6504, n_139, n_3372);
  not g7216 (n_3373, n6504);
  and g7217 (n6505, n3100, n_3373);
  not g7218 (n_3374, n6505);
  and g7219 (n6506, n_134, n_3374);
  not g7220 (n_3375, n6506);
  and g7221 (n6507, n6480, n_3375);
  not g7222 (n_3376, n6507);
  and g7223 (n6508, n_692, n_3376);
  and g7224 (n6509, n_3360, n6508);
  not g7225 (n_3377, n6509);
  and g7226 (n6510, n6197, n_3377);
  not g7227 (n_3378, n6490);
  not g7228 (n_3379, n6510);
  and g7229 (n6511, n_3378, n_3379);
  not g7230 (n_3380, n6511);
  and g7231 (n6512, n6310, n_3380);
  not g7232 (n_3381, n6512);
  and g7233 (n6513, n6418, n_3381);
  and g7234 (n6514, n6310, n_3361);
  not g7235 (n_3382, n6418);
  not g7236 (n_3383, n6514);
  and g7237 (n6515, n_3382, n_3383);
  not g7238 (n_3384, n6515);
  and g7239 (n6516, n_188, n_3384);
  not g7240 (n_3385, n6513);
  and g7241 (n6517, n_3385, n6516);
  not g7242 (n_3386, n6517);
  and g7243 (n6518, n6368, n_3386);
  and g7244 (n6519, n_305, n6487);
  not g7245 (n_3387, n6519);
  and g7246 (n6520, n6482, n_3387);
  not g7247 (n_3388, n6520);
  and g7248 (n6521, n_188, n_3388);
  not g7249 (n_3389, n6521);
  and g7250 (n6522, n_3237, n_3389);
  not g7251 (n_3390, n6522);
  and g7252 (n6523, n6326, n_3390);
  not g7253 (n_3391, n6523);
  and g7254 (n6524, n_234, n_3391);
  and g7258 (n6528, n_234, n6527);
  not g7259 (n_3396, n6524);
  not g7260 (n_3397, n6528);
  and g7261 (n6529, n_3396, n_3397);
  and g7262 (n6530, n_3102, n_3388);
  and g7263 (n6531, n6508, n_3387);
  not g7264 (n_3398, n6531);
  and g7265 (n6532, n6197, n_3398);
  not g7266 (n_3399, n6530);
  not g7267 (n_3400, n6532);
  and g7268 (n6533, n_3399, n_3400);
  and g7269 (n6534, n_188, n6326);
  not g7270 (n_3401, n6533);
  and g7271 (n6535, n_3401, n6534);
  not g7272 (n_3402, n6535);
  and g7273 (n6536, n_3268, n_3402);
  not g7274 (n_3403, n6536);
  and g7275 (n6537, n6527, n_3403);
  not g7276 (n_3404, n6529);
  not g7277 (n_3405, n6537);
  and g7278 (n6538, n_3404, n_3405);
  not g7279 (n_3407, n6518);
  and g7280 (n6539, pi0232, n_3407);
  not g7281 (n_3408, n6538);
  and g7282 (n6540, n_3408, n6539);
  and g7283 (n6541, n_188, n6514);
  not g7284 (n_3409, n6541);
  and g7285 (n6542, n6368, n_3409);
  not g7286 (n_3410, pi0232);
  not g7287 (n_3411, n6542);
  and g7288 (n6543, n_3410, n_3411);
  and g7289 (n6544, n_3396, n6543);
  not g7290 (n_3412, n6540);
  not g7291 (n_3413, n6544);
  and g7292 (n6545, n_3412, n_3413);
  not g7293 (n_3414, n6545);
  and g7294 (n6546, n_162, n_3414);
  not g7295 (n_3415, n6415);
  and g7296 (n6547, n_161, n_3415);
  not g7297 (n_3416, n6546);
  and g7298 (n6548, n_3416, n6547);
  and g7299 (n6549, pi0038, n_3250);
  not g7300 (n_3417, n6333);
  and g7301 (n6550, n_3417, n6549);
  not g7302 (n_3418, n6548);
  not g7303 (n_3419, n6550);
  and g7304 (n6551, n_3418, n_3419);
  not g7305 (n_3420, n6551);
  and g7306 (n6552, n_164, n_3420);
  not g7307 (n_3421, n6378);
  and g7308 (n6553, n_172, n_3421);
  not g7309 (n_3422, n6552);
  and g7310 (n6554, n_3422, n6553);
  not g7311 (n_3423, n6348);
  and g7312 (n6555, n_171, n_3423);
  not g7313 (n_3424, n6554);
  and g7314 (n6556, n_3424, n6555);
  not g7315 (n_3425, n6347);
  and g7316 (n6557, n_174, n_3425);
  not g7317 (n_3426, n6556);
  and g7318 (n6558, n_3426, n6557);
  not g7319 (n_3427, n6346);
  and g7320 (n6559, n_167, n_3427);
  not g7321 (n_3428, n6558);
  and g7322 (n6560, n_3428, n6559);
  not g7323 (n_3429, n6342);
  and g7324 (n6561, n_168, n_3429);
  not g7325 (n_3430, n6560);
  and g7326 (n6562, n_3430, n6561);
  not g7327 (n_3431, n6339);
  and g7328 (n6563, n_176, n_3431);
  not g7329 (n_3432, n6562);
  and g7330 (n6564, n_3432, n6563);
  not g7331 (n_3433, n6322);
  and g7332 (n6565, n2529, n_3433);
  not g7333 (n_3434, n6564);
  and g7334 (n6566, n_3434, n6565);
  not g7335 (n_3435, n6321);
  and g7336 (n6567, n_792, n_3435);
  not g7337 (n_3436, n6566);
  and g7338 (n6568, n_3436, n6567);
  not g7339 (n_3437, n6319);
  and g7340 (n6569, n_796, n_3437);
  not g7341 (n_3438, n6568);
  and g7342 (n6570, n_3438, n6569);
  not g7343 (n_3439, n6316);
  not g7344 (n_3440, n6570);
  and g7345 (po0171, n_3439, n_3440);
  and g7346 (n6572, n_3149, n6197);
  not g7347 (n_3441, n6226);
  not g7348 (n_3442, n6572);
  and g7349 (n6573, n_3441, n_3442);
  and g7350 (n6574, n6314, n6573);
  and g7351 (n6575, n6307, n6574);
  and g7352 (n6576, n_3241, n6574);
  not g7353 (n_3443, n6576);
  and g7354 (n6577, pi0059, n_3443);
  and g7355 (n6578, n6312, n6573);
  and g7356 (n6579, n_3243, n6578);
  not g7357 (n_3444, n6574);
  and g7358 (n6580, pi0055, n_3444);
  not g7359 (n_3445, n6573);
  and g7360 (n6581, pi0299, n_3445);
  and g7361 (n6582, n_3105, n6197);
  not g7362 (n_3446, n6582);
  and g7363 (n6583, n_3441, n_3446);
  not g7364 (n_3447, n6583);
  and g7365 (n6584, n_234, n_3447);
  not g7366 (n_3448, n6581);
  not g7367 (n_3449, n6584);
  and g7368 (n6585, n_3448, n_3449);
  and g7369 (n6586, n6312, n6585);
  not g7370 (n_3450, n6586);
  and g7371 (n6587, n_3249, n_3450);
  and g7372 (n6588, n_766, n6586);
  and g7373 (n6589, n6332, n6585);
  and g7374 (n6590, n2620, n6589);
  not g7375 (n_3451, n6588);
  not g7376 (n_3452, n6590);
  and g7377 (n6591, n_3451, n_3452);
  and g7378 (n6592, n2569, n6591);
  and g7379 (n6593, n_167, n6592);
  not g7380 (n_3453, n6587);
  and g7381 (n6594, pi0074, n_3453);
  not g7382 (n_3454, n6593);
  and g7383 (n6595, n_3454, n6594);
  and g7384 (n6596, n_3255, n_3450);
  not g7385 (n_3455, n6592);
  not g7386 (n_3456, n6596);
  and g7387 (n6597, n_3455, n_3456);
  not g7388 (n_3457, n6597);
  and g7389 (n6598, pi0054, n_3457);
  and g7390 (n6599, n_171, n6591);
  and g7391 (n6600, pi0075, n_3450);
  not g7392 (n_3458, n6600);
  and g7393 (n6601, pi0092, n_3458);
  not g7394 (n_3459, n6599);
  and g7395 (n6602, n_3459, n6601);
  and g7396 (n6603, pi0075, n6591);
  and g7397 (n6604, pi0087, n6586);
  and g7398 (n6605, n_260, n6586);
  not g7399 (n_3460, n6578);
  and g7400 (n6606, pi0299, n_3460);
  and g7401 (n6607, n_3441, n6353);
  and g7402 (n6608, n2640, n_3442);
  and g7403 (n6609, n6607, n6608);
  not g7404 (n_3461, n6357);
  and g7405 (n6610, n_3138, n_3461);
  not g7406 (n_3462, n6359);
  and g7407 (n6611, n6192, n_3462);
  not g7408 (n_3463, n6610);
  not g7409 (n_3464, n6611);
  and g7410 (n6612, n_3463, n_3464);
  and g7411 (n6613, n6192, n_3102);
  not g7412 (n_3465, n6613);
  and g7413 (n6614, n_3149, n_3465);
  not g7414 (n_3466, n6614);
  and g7415 (n6615, n_272, n_3466);
  and g7416 (n6616, n6612, n6615);
  not g7417 (n_3467, n6609);
  not g7418 (n_3468, n6616);
  and g7419 (n6617, n_3467, n_3468);
  not g7420 (n_3469, n6617);
  and g7421 (n6618, n_188, n_3469);
  not g7422 (n_3470, n6618);
  and g7423 (n6619, n6606, n_3470);
  and g7424 (n6620, n_188, n2669);
  and g7425 (n6621, n_3446, n6612);
  not g7426 (n_3471, n6621);
  and g7427 (n6622, n6620, n_3471);
  and g7428 (n6623, n_3105, n_3465);
  not g7429 (n_3472, n6612);
  and g7430 (n6624, pi0142, n_3472);
  not g7431 (n_3473, n6607);
  and g7432 (n6625, n_738, n_3473);
  and g7439 (n6629, n6312, n6583);
  not g7440 (n_3477, n6620);
  not g7441 (n_3478, n6629);
  and g7442 (n6630, n_3477, n_3478);
  not g7443 (n_3479, n6628);
  and g7444 (n6631, n_3479, n6630);
  not g7445 (n_3480, n6622);
  not g7446 (n_3481, n6631);
  and g7447 (n6632, n_3480, n_3481);
  not g7448 (n_3482, n6632);
  and g7449 (n6633, n_234, n_3482);
  not g7450 (n_3483, n6619);
  and g7451 (n6634, n2530, n_3483);
  not g7452 (n_3484, n6633);
  and g7453 (n6635, n_3484, n6634);
  not g7454 (n_3485, n6605);
  and g7455 (n6636, pi0100, n_3485);
  not g7456 (n_3486, n6635);
  and g7457 (n6637, n_3486, n6636);
  and g7458 (n6638, n_3299, n6583);
  not g7459 (n_3487, n6638);
  and g7460 (n6639, n_234, n_3487);
  and g7461 (n6640, pi0299, n6379);
  not g7462 (n_3488, n6606);
  not g7463 (n_3489, n6640);
  and g7464 (n6641, n_3488, n_3489);
  and g7465 (n6642, n6401, n6573);
  not g7466 (n_3490, n6641);
  not g7467 (n_3491, n6642);
  and g7468 (n6643, n_3490, n_3491);
  not g7469 (n_3492, n6639);
  and g7470 (n6644, pi0039, n_3492);
  not g7471 (n_3493, n6643);
  and g7472 (n6645, n_3493, n6644);
  and g7473 (n6646, n_3380, n6573);
  not g7474 (n_3494, n6646);
  and g7475 (n6647, n6418, n_3494);
  and g7476 (n6648, n_3361, n6573);
  not g7477 (n_3495, n6648);
  and g7478 (n6649, n_3382, n_3495);
  not g7479 (n_3496, n6649);
  and g7480 (n6650, n_188, n_3496);
  not g7481 (n_3497, n6647);
  and g7482 (n6651, n_3497, n6650);
  not g7483 (n_3498, n6651);
  and g7484 (n6652, n6606, n_3498);
  and g7485 (n6653, n_3390, n6583);
  not g7486 (n_3499, n6527);
  and g7487 (n6654, n_3499, n6653);
  and g7488 (n6655, n_188, n6583);
  and g7489 (n6656, n_3401, n6655);
  not g7490 (n_3500, n6656);
  and g7491 (n6657, n_3478, n_3500);
  not g7492 (n_3501, n6657);
  and g7493 (n6658, n6527, n_3501);
  not g7494 (n_3502, n6654);
  and g7495 (n6659, n_234, n_3502);
  not g7496 (n_3503, n6658);
  and g7497 (n6660, n_3503, n6659);
  not g7498 (n_3504, n6652);
  and g7499 (n6661, pi0232, n_3504);
  not g7500 (n_3505, n6660);
  and g7501 (n6662, n_3505, n6661);
  and g7502 (n6663, n_188, n6648);
  not g7503 (n_3506, n6663);
  and g7504 (n6664, n6606, n_3506);
  not g7505 (n_3507, n6653);
  and g7506 (n6665, n_234, n_3507);
  not g7507 (n_3508, n6664);
  and g7508 (n6666, n_3410, n_3508);
  not g7509 (n_3509, n6665);
  and g7510 (n6667, n_3509, n6666);
  not g7511 (n_3510, n6662);
  not g7512 (n_3511, n6667);
  and g7513 (n6668, n_3510, n_3511);
  not g7514 (n_3512, n6668);
  and g7515 (n6669, n_162, n_3512);
  not g7516 (n_3513, n6645);
  and g7517 (n6670, n_161, n_3513);
  not g7518 (n_3514, n6669);
  and g7519 (n6671, n_3514, n6670);
  and g7520 (n6672, pi0038, n_3450);
  not g7521 (n_3515, n6589);
  and g7522 (n6673, n_3515, n6672);
  not g7523 (n_3516, n6671);
  not g7524 (n_3517, n6673);
  and g7525 (n6674, n_3516, n_3517);
  not g7526 (n_3518, n6674);
  and g7527 (n6675, n_164, n_3518);
  not g7528 (n_3519, n6637);
  and g7529 (n6676, n_172, n_3519);
  not g7530 (n_3520, n6675);
  and g7531 (n6677, n_3520, n6676);
  not g7532 (n_3521, n6604);
  and g7533 (n6678, n_171, n_3521);
  not g7534 (n_3522, n6677);
  and g7535 (n6679, n_3522, n6678);
  not g7536 (n_3523, n6603);
  and g7537 (n6680, n_174, n_3523);
  not g7538 (n_3524, n6679);
  and g7539 (n6681, n_3524, n6680);
  not g7540 (n_3525, n6602);
  and g7541 (n6682, n_167, n_3525);
  not g7542 (n_3526, n6681);
  and g7543 (n6683, n_3526, n6682);
  not g7544 (n_3527, n6598);
  and g7545 (n6684, n_168, n_3527);
  not g7546 (n_3528, n6683);
  and g7547 (n6685, n_3528, n6684);
  not g7548 (n_3529, n6595);
  and g7549 (n6686, n_176, n_3529);
  not g7550 (n_3530, n6685);
  and g7551 (n6687, n_3530, n6686);
  not g7552 (n_3531, n6580);
  and g7553 (n6688, n2529, n_3531);
  not g7554 (n_3532, n6687);
  and g7555 (n6689, n_3532, n6688);
  not g7556 (n_3533, n6579);
  and g7557 (n6690, n_792, n_3533);
  not g7558 (n_3534, n6689);
  and g7559 (n6691, n_3534, n6690);
  not g7560 (n_3535, n6577);
  and g7561 (n6692, n_796, n_3535);
  not g7562 (n_3536, n6691);
  and g7563 (n6693, n_3536, n6692);
  not g7564 (n_3537, n6575);
  not g7565 (n_3538, n6693);
  and g7566 (po0172, n_3537, n_3538);
  and g7567 (n6695, pi0030, n6197);
  and g7568 (n6696, pi0228, n6695);
  and g7569 (n6697, pi0970, n6696);
  and g7570 (n6698, n_188, pi0970);
  and g7571 (n6699, n6222, n6698);
  and g7572 (n6700, n2572, n6699);
  and g7573 (n6701, n6305, n6700);
  not g7574 (n_3539, n6697);
  not g7575 (n_3540, n6701);
  and g7576 (n6702, n_3539, n_3540);
  not g7577 (n_3541, n6702);
  and g7578 (n6703, pi0057, n_3541);
  and g7579 (n6704, n6304, n6700);
  and g7580 (n6705, pi0059, n_3539);
  not g7581 (n_3542, n6704);
  and g7582 (n6706, n_3542, n6705);
  and g7583 (n6707, n_3243, n6697);
  and g7584 (n6708, pi0055, n_3539);
  not g7585 (n_3543, n6700);
  and g7586 (n6709, n_3543, n6708);
  and g7587 (n6710, pi0299, pi0970);
  and g7588 (n6711, n_234, pi0967);
  not g7589 (n_3544, n6710);
  not g7590 (n_3545, n6711);
  and g7591 (n6712, n_3544, n_3545);
  not g7592 (n_3546, n6712);
  and g7593 (n6713, n6696, n_3546);
  not g7594 (n_3547, n6713);
  and g7595 (n6714, n_3249, n_3547);
  and g7596 (n6715, n_766, n6713);
  and g7597 (n6716, pi0299, n_3539);
  not g7598 (n_3548, n6699);
  and g7599 (n6717, n_3548, n6716);
  not g7600 (n_3549, n6695);
  and g7601 (n6718, pi0228, n_3549);
  not g7602 (n_3550, n6222);
  and g7603 (n6719, n_188, n_3550);
  not g7604 (n_3551, n6718);
  not g7605 (n_3552, n6719);
  and g7606 (n6720, n_3551, n_3552);
  and g7607 (n6721, pi0967, n6720);
  not g7608 (n_3553, n6721);
  and g7609 (n6722, n_234, n_3553);
  not g7610 (n_3554, n6717);
  and g7611 (n6723, n_162, n_3554);
  not g7612 (n_3555, n6722);
  and g7613 (n6724, n_3555, n6723);
  and g7614 (n6725, n2620, n6724);
  not g7615 (n_3556, n6715);
  not g7616 (n_3557, n6725);
  and g7617 (n6726, n_3556, n_3557);
  and g7618 (n6727, n2569, n6726);
  and g7619 (n6728, n_167, n6727);
  not g7620 (n_3558, n6714);
  and g7621 (n6729, pi0074, n_3558);
  not g7622 (n_3559, n6728);
  and g7623 (n6730, n_3559, n6729);
  and g7624 (n6731, n_3255, n_3547);
  not g7625 (n_3560, n6727);
  not g7626 (n_3561, n6731);
  and g7627 (n6732, n_3560, n_3561);
  not g7628 (n_3562, n6732);
  and g7629 (n6733, pi0054, n_3562);
  and g7630 (n6734, n_171, n6726);
  and g7631 (n6735, pi0075, n_3547);
  not g7632 (n_3563, n6735);
  and g7633 (n6736, pi0092, n_3563);
  not g7634 (n_3564, n6734);
  and g7635 (n6737, n_3564, n6736);
  and g7636 (n6738, pi0075, n6726);
  and g7637 (n6739, pi0087, n6713);
  and g7638 (n6740, n_260, n6713);
  and g7639 (n6741, n_272, n_3461);
  and g7640 (n6742, n6197, n6353);
  not g7641 (n_3565, n6742);
  and g7642 (n6743, n2640, n_3565);
  not g7643 (n_3566, n6741);
  and g7644 (n6744, n_188, n_3566);
  not g7645 (n_3567, n6743);
  and g7646 (n6745, n_3567, n6744);
  and g7647 (n6746, pi0970, n6745);
  not g7648 (n_3568, n6746);
  and g7649 (n6747, n6716, n_3568);
  and g7650 (n6748, n_3261, n6357);
  and g7651 (n6749, n6260, n6742);
  not g7652 (n_3569, n6748);
  and g7653 (n6750, n_188, n_3569);
  not g7654 (n_3570, n6749);
  and g7655 (n6751, n_3570, n6750);
  not g7656 (n_3571, n6751);
  and g7657 (n6752, n_3551, n_3571);
  and g7658 (n6753, pi0967, n6752);
  not g7659 (n_3572, n6753);
  and g7660 (n6754, n_234, n_3572);
  not g7661 (n_3573, n6747);
  and g7662 (n6755, n2530, n_3573);
  not g7663 (n_3574, n6754);
  and g7664 (n6756, n_3574, n6755);
  not g7665 (n_3575, n6740);
  and g7666 (n6757, pi0100, n_3575);
  not g7667 (n_3576, n6756);
  and g7668 (n6758, n_3576, n6757);
  and g7669 (n6759, n6379, n_3289);
  and g7670 (n6760, n6197, n6759);
  not g7671 (n_3577, n6760);
  and g7672 (n6761, n_188, n_3577);
  not g7673 (n_3578, n6761);
  and g7674 (n6762, n6710, n_3578);
  and g7675 (n6763, n6197, n6409);
  not g7676 (n_3579, n6763);
  and g7677 (n6764, n_188, n_3579);
  not g7678 (n_3580, n6764);
  and g7679 (n6765, n6711, n_3580);
  not g7680 (n_3581, n6762);
  not g7681 (n_3582, n6765);
  and g7682 (n6766, n_3581, n_3582);
  and g7683 (n6767, pi0039, n_3551);
  not g7684 (n_3583, n6766);
  and g7685 (n6768, n_3583, n6767);
  and g7686 (n6769, n6197, n_3390);
  not g7687 (n_3584, n6769);
  and g7688 (n6770, n_3499, n_3584);
  and g7689 (n6771, n_3388, n_3499);
  and g7690 (n6772, n_188, n6532);
  not g7691 (n_3585, n6696);
  not g7692 (n_3586, n6771);
  and g7693 (n6773, n_3585, n_3586);
  not g7694 (n_3587, n6772);
  and g7695 (n6774, n_3587, n6773);
  not g7696 (n_3588, n6770);
  not g7697 (n_3589, n6774);
  and g7698 (n6775, n_3588, n_3589);
  and g7699 (n6776, pi0967, n6775);
  not g7700 (n_3590, n6776);
  and g7701 (n6777, n_234, n_3590);
  and g7702 (n6778, n6197, n_3361);
  and g7703 (n6779, n6698, n6778);
  not g7704 (n_3591, n6779);
  and g7705 (n6780, n6716, n_3591);
  and g7706 (n6781, pi0299, n6416);
  not g7707 (n_3592, n6780);
  not g7708 (n_3593, n6781);
  and g7709 (n6782, n_3592, n_3593);
  and g7710 (n6783, n6417, n_3379);
  not g7711 (n_3594, n6417);
  and g7712 (n6784, n_3594, n6489);
  not g7713 (n_3595, n6783);
  not g7714 (n_3596, n6784);
  and g7715 (n6785, n_3595, n_3596);
  and g7716 (n6786, n6197, n6785);
  and g7717 (n6787, n6698, n6786);
  not g7718 (n_3597, n6787);
  and g7719 (n6788, n_3539, n_3597);
  not g7720 (n_3598, n6788);
  and g7721 (n6789, n6416, n_3598);
  not g7722 (n_3599, n6782);
  not g7723 (n_3600, n6789);
  and g7724 (n6790, n_3599, n_3600);
  not g7725 (n_3601, n6777);
  and g7726 (n6791, pi0232, n_3601);
  not g7727 (n_3602, n6790);
  and g7728 (n6792, n_3602, n6791);
  and g7729 (n6793, pi0967, n6769);
  not g7730 (n_3603, n6793);
  and g7731 (n6794, n_234, n_3603);
  and g7732 (n6795, n_3410, n_3592);
  not g7733 (n_3604, n6794);
  and g7734 (n6796, n_3604, n6795);
  not g7735 (n_3605, n6792);
  not g7736 (n_3606, n6796);
  and g7737 (n6797, n_3605, n_3606);
  not g7738 (n_3607, n6797);
  and g7739 (n6798, n_162, n_3607);
  not g7740 (n_3608, n6768);
  and g7741 (n6799, n_161, n_3608);
  not g7742 (n_3609, n6798);
  and g7743 (n6800, n_3609, n6799);
  and g7744 (n6801, pi0039, n6713);
  not g7745 (n_3610, n6801);
  and g7746 (n6802, pi0038, n_3610);
  not g7747 (n_3611, n6724);
  and g7748 (n6803, n_3611, n6802);
  not g7749 (n_3612, n6800);
  not g7750 (n_3613, n6803);
  and g7751 (n6804, n_3612, n_3613);
  not g7752 (n_3614, n6804);
  and g7753 (n6805, n_164, n_3614);
  not g7754 (n_3615, n6758);
  and g7755 (n6806, n_172, n_3615);
  not g7756 (n_3616, n6805);
  and g7757 (n6807, n_3616, n6806);
  not g7758 (n_3617, n6739);
  and g7759 (n6808, n_171, n_3617);
  not g7760 (n_3618, n6807);
  and g7761 (n6809, n_3618, n6808);
  not g7762 (n_3619, n6738);
  and g7763 (n6810, n_174, n_3619);
  not g7764 (n_3620, n6809);
  and g7765 (n6811, n_3620, n6810);
  not g7766 (n_3621, n6737);
  and g7767 (n6812, n_167, n_3621);
  not g7768 (n_3622, n6811);
  and g7769 (n6813, n_3622, n6812);
  not g7770 (n_3623, n6733);
  and g7771 (n6814, n_168, n_3623);
  not g7772 (n_3624, n6813);
  and g7773 (n6815, n_3624, n6814);
  not g7774 (n_3625, n6730);
  and g7775 (n6816, n_176, n_3625);
  not g7776 (n_3626, n6815);
  and g7777 (n6817, n_3626, n6816);
  not g7778 (n_3627, n6709);
  and g7779 (n6818, n2529, n_3627);
  not g7780 (n_3628, n6817);
  and g7781 (n6819, n_3628, n6818);
  not g7782 (n_3629, n6707);
  and g7783 (n6820, n_792, n_3629);
  not g7784 (n_3630, n6819);
  and g7785 (n6821, n_3630, n6820);
  not g7786 (n_3631, n6706);
  and g7787 (n6822, n_796, n_3631);
  not g7788 (n_3632, n6821);
  and g7789 (n6823, n_3632, n6822);
  not g7790 (n_3633, n6703);
  not g7791 (n_3634, n6823);
  and g7792 (po0173, n_3633, n_3634);
  and g7793 (n6825, pi0972, n6696);
  and g7794 (n6826, n_188, pi0972);
  and g7795 (n6827, n6222, n6826);
  and g7796 (n6828, n2572, n6827);
  and g7797 (n6829, n6305, n6828);
  not g7798 (n_3635, n6825);
  not g7799 (n_3636, n6829);
  and g7800 (n6830, n_3635, n_3636);
  not g7801 (n_3637, n6830);
  and g7802 (n6831, pi0057, n_3637);
  and g7803 (n6832, n6304, n6828);
  and g7804 (n6833, pi0059, n_3635);
  not g7805 (n_3638, n6832);
  and g7806 (n6834, n_3638, n6833);
  and g7807 (n6835, n_3243, n6825);
  and g7808 (n6836, pi0055, n_3635);
  not g7809 (n_3639, n6828);
  and g7810 (n6837, n_3639, n6836);
  and g7811 (n6838, n_234, pi0961);
  and g7812 (n6839, pi0299, pi0972);
  not g7813 (n_3640, n6838);
  not g7814 (n_3641, n6839);
  and g7815 (n6840, n_3640, n_3641);
  not g7816 (n_3642, n6840);
  and g7817 (n6841, n6696, n_3642);
  not g7818 (n_3643, n6841);
  and g7819 (n6842, n_3249, n_3643);
  and g7820 (n6843, n_766, n6841);
  and g7821 (n6844, pi0299, n_3635);
  not g7822 (n_3644, n6827);
  and g7823 (n6845, n_3644, n6844);
  and g7824 (n6846, pi0961, n6720);
  not g7825 (n_3645, n6846);
  and g7826 (n6847, n_234, n_3645);
  not g7827 (n_3646, n6845);
  and g7828 (n6848, n_162, n_3646);
  not g7829 (n_3647, n6847);
  and g7830 (n6849, n_3647, n6848);
  and g7831 (n6850, n2620, n6849);
  not g7832 (n_3648, n6843);
  not g7833 (n_3649, n6850);
  and g7834 (n6851, n_3648, n_3649);
  and g7835 (n6852, n2569, n6851);
  and g7836 (n6853, n_167, n6852);
  not g7837 (n_3650, n6842);
  and g7838 (n6854, pi0074, n_3650);
  not g7839 (n_3651, n6853);
  and g7840 (n6855, n_3651, n6854);
  and g7841 (n6856, n_3255, n_3643);
  not g7842 (n_3652, n6852);
  not g7843 (n_3653, n6856);
  and g7844 (n6857, n_3652, n_3653);
  not g7845 (n_3654, n6857);
  and g7846 (n6858, pi0054, n_3654);
  and g7847 (n6859, n_171, n6851);
  and g7848 (n6860, pi0075, n_3643);
  not g7849 (n_3655, n6860);
  and g7850 (n6861, pi0092, n_3655);
  not g7851 (n_3656, n6859);
  and g7852 (n6862, n_3656, n6861);
  and g7853 (n6863, pi0075, n6851);
  and g7854 (n6864, pi0087, n6841);
  and g7855 (n6865, n_260, n6841);
  and g7856 (n6866, pi0972, n6745);
  not g7857 (n_3657, n6866);
  and g7858 (n6867, n6844, n_3657);
  and g7859 (n6868, pi0961, n6752);
  not g7860 (n_3658, n6868);
  and g7861 (n6869, n_234, n_3658);
  not g7862 (n_3659, n6867);
  and g7863 (n6870, n2530, n_3659);
  not g7864 (n_3660, n6869);
  and g7865 (n6871, n_3660, n6870);
  not g7866 (n_3661, n6865);
  and g7867 (n6872, pi0100, n_3661);
  not g7868 (n_3662, n6871);
  and g7869 (n6873, n_3662, n6872);
  and g7870 (n6874, n_3580, n6838);
  and g7871 (n6875, n_3578, n6839);
  not g7872 (n_3663, n6874);
  not g7873 (n_3664, n6875);
  and g7874 (n6876, n_3663, n_3664);
  not g7875 (n_3665, n6876);
  and g7876 (n6877, n6767, n_3665);
  and g7877 (n6878, pi0961, n6775);
  not g7878 (n_3666, n6878);
  and g7879 (n6879, n_234, n_3666);
  and g7880 (n6880, n6778, n6826);
  not g7881 (n_3667, n6880);
  and g7882 (n6881, n6844, n_3667);
  not g7883 (n_3668, n6881);
  and g7884 (n6882, n_3593, n_3668);
  and g7885 (n6883, n6786, n6826);
  not g7886 (n_3669, n6883);
  and g7887 (n6884, n_3635, n_3669);
  not g7888 (n_3670, n6884);
  and g7889 (n6885, n6416, n_3670);
  not g7890 (n_3671, n6882);
  not g7891 (n_3672, n6885);
  and g7892 (n6886, n_3671, n_3672);
  not g7893 (n_3673, n6879);
  and g7894 (n6887, pi0232, n_3673);
  not g7895 (n_3674, n6886);
  and g7896 (n6888, n_3674, n6887);
  and g7897 (n6889, pi0961, n6769);
  not g7898 (n_3675, n6889);
  and g7899 (n6890, n_234, n_3675);
  and g7900 (n6891, n_3410, n_3668);
  not g7901 (n_3676, n6890);
  and g7902 (n6892, n_3676, n6891);
  not g7903 (n_3677, n6888);
  not g7904 (n_3678, n6892);
  and g7905 (n6893, n_3677, n_3678);
  not g7906 (n_3679, n6893);
  and g7907 (n6894, n_162, n_3679);
  not g7908 (n_3680, n6877);
  and g7909 (n6895, n_161, n_3680);
  not g7910 (n_3681, n6894);
  and g7911 (n6896, n_3681, n6895);
  and g7912 (n6897, pi0039, n6841);
  not g7913 (n_3682, n6897);
  and g7914 (n6898, pi0038, n_3682);
  not g7915 (n_3683, n6849);
  and g7916 (n6899, n_3683, n6898);
  not g7917 (n_3684, n6896);
  not g7918 (n_3685, n6899);
  and g7919 (n6900, n_3684, n_3685);
  not g7920 (n_3686, n6900);
  and g7921 (n6901, n_164, n_3686);
  not g7922 (n_3687, n6873);
  and g7923 (n6902, n_172, n_3687);
  not g7924 (n_3688, n6901);
  and g7925 (n6903, n_3688, n6902);
  not g7926 (n_3689, n6864);
  and g7927 (n6904, n_171, n_3689);
  not g7928 (n_3690, n6903);
  and g7929 (n6905, n_3690, n6904);
  not g7930 (n_3691, n6863);
  and g7931 (n6906, n_174, n_3691);
  not g7932 (n_3692, n6905);
  and g7933 (n6907, n_3692, n6906);
  not g7934 (n_3693, n6862);
  and g7935 (n6908, n_167, n_3693);
  not g7936 (n_3694, n6907);
  and g7937 (n6909, n_3694, n6908);
  not g7938 (n_3695, n6858);
  and g7939 (n6910, n_168, n_3695);
  not g7940 (n_3696, n6909);
  and g7941 (n6911, n_3696, n6910);
  not g7942 (n_3697, n6855);
  and g7943 (n6912, n_176, n_3697);
  not g7944 (n_3698, n6911);
  and g7945 (n6913, n_3698, n6912);
  not g7946 (n_3699, n6837);
  and g7947 (n6914, n2529, n_3699);
  not g7948 (n_3700, n6913);
  and g7949 (n6915, n_3700, n6914);
  not g7950 (n_3701, n6835);
  and g7951 (n6916, n_792, n_3701);
  not g7952 (n_3702, n6915);
  and g7953 (n6917, n_3702, n6916);
  not g7954 (n_3703, n6834);
  and g7955 (n6918, n_796, n_3703);
  not g7956 (n_3704, n6917);
  and g7957 (n6919, n_3704, n6918);
  not g7958 (n_3705, n6831);
  not g7959 (n_3706, n6919);
  and g7960 (po0174, n_3705, n_3706);
  and g7961 (n6921, pi0960, n6696);
  and g7962 (n6922, n_188, pi0960);
  and g7963 (n6923, n6222, n6922);
  and g7964 (n6924, n2572, n6923);
  and g7965 (n6925, n6305, n6924);
  not g7966 (n_3707, n6921);
  not g7967 (n_3708, n6925);
  and g7968 (n6926, n_3707, n_3708);
  not g7969 (n_3709, n6926);
  and g7970 (n6927, pi0057, n_3709);
  and g7971 (n6928, n6304, n6924);
  and g7972 (n6929, pi0059, n_3707);
  not g7973 (n_3710, n6928);
  and g7974 (n6930, n_3710, n6929);
  and g7975 (n6931, n_3243, n6921);
  and g7976 (n6932, pi0055, n_3707);
  not g7977 (n_3711, n6924);
  and g7978 (n6933, n_3711, n6932);
  and g7979 (n6934, n_234, pi0977);
  and g7980 (n6935, pi0299, pi0960);
  not g7981 (n_3712, n6934);
  not g7982 (n_3713, n6935);
  and g7983 (n6936, n_3712, n_3713);
  not g7984 (n_3714, n6936);
  and g7985 (n6937, n6696, n_3714);
  not g7986 (n_3715, n6937);
  and g7987 (n6938, n_3249, n_3715);
  and g7988 (n6939, n_766, n6937);
  and g7989 (n6940, pi0299, n_3707);
  not g7990 (n_3716, n6923);
  and g7991 (n6941, n_3716, n6940);
  and g7992 (n6942, pi0977, n6720);
  not g7993 (n_3717, n6942);
  and g7994 (n6943, n_234, n_3717);
  not g7995 (n_3718, n6941);
  and g7996 (n6944, n_162, n_3718);
  not g7997 (n_3719, n6943);
  and g7998 (n6945, n_3719, n6944);
  and g7999 (n6946, n2620, n6945);
  not g8000 (n_3720, n6939);
  not g8001 (n_3721, n6946);
  and g8002 (n6947, n_3720, n_3721);
  and g8003 (n6948, n2569, n6947);
  and g8004 (n6949, n_167, n6948);
  not g8005 (n_3722, n6938);
  and g8006 (n6950, pi0074, n_3722);
  not g8007 (n_3723, n6949);
  and g8008 (n6951, n_3723, n6950);
  and g8009 (n6952, n_3255, n_3715);
  not g8010 (n_3724, n6948);
  not g8011 (n_3725, n6952);
  and g8012 (n6953, n_3724, n_3725);
  not g8013 (n_3726, n6953);
  and g8014 (n6954, pi0054, n_3726);
  and g8015 (n6955, n_171, n6947);
  and g8016 (n6956, pi0075, n_3715);
  not g8017 (n_3727, n6956);
  and g8018 (n6957, pi0092, n_3727);
  not g8019 (n_3728, n6955);
  and g8020 (n6958, n_3728, n6957);
  and g8021 (n6959, pi0075, n6947);
  and g8022 (n6960, pi0087, n6937);
  and g8023 (n6961, n_260, n6937);
  and g8024 (n6962, pi0960, n6745);
  not g8025 (n_3729, n6962);
  and g8026 (n6963, n6940, n_3729);
  and g8027 (n6964, pi0977, n6752);
  not g8028 (n_3730, n6964);
  and g8029 (n6965, n_234, n_3730);
  not g8030 (n_3731, n6963);
  and g8031 (n6966, n2530, n_3731);
  not g8032 (n_3732, n6965);
  and g8033 (n6967, n_3732, n6966);
  not g8034 (n_3733, n6961);
  and g8035 (n6968, pi0100, n_3733);
  not g8036 (n_3734, n6967);
  and g8037 (n6969, n_3734, n6968);
  and g8038 (n6970, n_3580, n6934);
  and g8039 (n6971, n_3578, n6935);
  not g8040 (n_3735, n6970);
  not g8041 (n_3736, n6971);
  and g8042 (n6972, n_3735, n_3736);
  not g8043 (n_3737, n6972);
  and g8044 (n6973, n6767, n_3737);
  and g8045 (n6974, pi0977, n6775);
  not g8046 (n_3738, n6974);
  and g8047 (n6975, n_234, n_3738);
  and g8048 (n6976, n6778, n6922);
  not g8049 (n_3739, n6976);
  and g8050 (n6977, n6940, n_3739);
  not g8051 (n_3740, n6977);
  and g8052 (n6978, n_3593, n_3740);
  and g8053 (n6979, n6786, n6922);
  not g8054 (n_3741, n6979);
  and g8055 (n6980, n_3707, n_3741);
  not g8056 (n_3742, n6980);
  and g8057 (n6981, n6416, n_3742);
  not g8058 (n_3743, n6978);
  not g8059 (n_3744, n6981);
  and g8060 (n6982, n_3743, n_3744);
  not g8061 (n_3745, n6975);
  and g8062 (n6983, pi0232, n_3745);
  not g8063 (n_3746, n6982);
  and g8064 (n6984, n_3746, n6983);
  and g8065 (n6985, pi0977, n6769);
  not g8066 (n_3747, n6985);
  and g8067 (n6986, n_234, n_3747);
  and g8068 (n6987, n_3410, n_3740);
  not g8069 (n_3748, n6986);
  and g8070 (n6988, n_3748, n6987);
  not g8071 (n_3749, n6984);
  not g8072 (n_3750, n6988);
  and g8073 (n6989, n_3749, n_3750);
  not g8074 (n_3751, n6989);
  and g8075 (n6990, n_162, n_3751);
  not g8076 (n_3752, n6973);
  and g8077 (n6991, n_161, n_3752);
  not g8078 (n_3753, n6990);
  and g8079 (n6992, n_3753, n6991);
  and g8080 (n6993, pi0039, n6937);
  not g8081 (n_3754, n6993);
  and g8082 (n6994, pi0038, n_3754);
  not g8083 (n_3755, n6945);
  and g8084 (n6995, n_3755, n6994);
  not g8085 (n_3756, n6992);
  not g8086 (n_3757, n6995);
  and g8087 (n6996, n_3756, n_3757);
  not g8088 (n_3758, n6996);
  and g8089 (n6997, n_164, n_3758);
  not g8090 (n_3759, n6969);
  and g8091 (n6998, n_172, n_3759);
  not g8092 (n_3760, n6997);
  and g8093 (n6999, n_3760, n6998);
  not g8094 (n_3761, n6960);
  and g8095 (n7000, n_171, n_3761);
  not g8096 (n_3762, n6999);
  and g8097 (n7001, n_3762, n7000);
  not g8098 (n_3763, n6959);
  and g8099 (n7002, n_174, n_3763);
  not g8100 (n_3764, n7001);
  and g8101 (n7003, n_3764, n7002);
  not g8102 (n_3765, n6958);
  and g8103 (n7004, n_167, n_3765);
  not g8104 (n_3766, n7003);
  and g8105 (n7005, n_3766, n7004);
  not g8106 (n_3767, n6954);
  and g8107 (n7006, n_168, n_3767);
  not g8108 (n_3768, n7005);
  and g8109 (n7007, n_3768, n7006);
  not g8110 (n_3769, n6951);
  and g8111 (n7008, n_176, n_3769);
  not g8112 (n_3770, n7007);
  and g8113 (n7009, n_3770, n7008);
  not g8114 (n_3771, n6933);
  and g8115 (n7010, n2529, n_3771);
  not g8116 (n_3772, n7009);
  and g8117 (n7011, n_3772, n7010);
  not g8118 (n_3773, n6931);
  and g8119 (n7012, n_792, n_3773);
  not g8120 (n_3774, n7011);
  and g8121 (n7013, n_3774, n7012);
  not g8122 (n_3775, n6930);
  and g8123 (n7014, n_796, n_3775);
  not g8124 (n_3776, n7013);
  and g8125 (n7015, n_3776, n7014);
  not g8126 (n_3777, n6927);
  not g8127 (n_3778, n7015);
  and g8128 (po0175, n_3777, n_3778);
  and g8129 (n7017, pi0963, n6696);
  and g8130 (n7018, n_188, pi0963);
  and g8131 (n7019, n6222, n7018);
  and g8132 (n7020, n2572, n7019);
  and g8133 (n7021, n6305, n7020);
  not g8134 (n_3779, n7017);
  not g8135 (n_3780, n7021);
  and g8136 (n7022, n_3779, n_3780);
  not g8137 (n_3781, n7022);
  and g8138 (n7023, pi0057, n_3781);
  and g8139 (n7024, n6304, n7020);
  and g8140 (n7025, pi0059, n_3779);
  not g8141 (n_3782, n7024);
  and g8142 (n7026, n_3782, n7025);
  and g8143 (n7027, n_3243, n7017);
  and g8144 (n7028, pi0055, n_3779);
  not g8145 (n_3783, n7020);
  and g8146 (n7029, n_3783, n7028);
  and g8147 (n7030, n_234, pi0969);
  and g8148 (n7031, pi0299, pi0963);
  not g8149 (n_3784, n7030);
  not g8150 (n_3785, n7031);
  and g8151 (n7032, n_3784, n_3785);
  not g8152 (n_3786, n7032);
  and g8153 (n7033, n6696, n_3786);
  not g8154 (n_3787, n7033);
  and g8155 (n7034, n_3249, n_3787);
  and g8156 (n7035, n_766, n7033);
  and g8157 (n7036, pi0299, n_3779);
  not g8158 (n_3788, n7019);
  and g8159 (n7037, n_3788, n7036);
  and g8160 (n7038, pi0969, n6720);
  not g8161 (n_3789, n7038);
  and g8162 (n7039, n_234, n_3789);
  not g8163 (n_3790, n7037);
  and g8164 (n7040, n_162, n_3790);
  not g8165 (n_3791, n7039);
  and g8166 (n7041, n_3791, n7040);
  and g8167 (n7042, n2620, n7041);
  not g8168 (n_3792, n7035);
  not g8169 (n_3793, n7042);
  and g8170 (n7043, n_3792, n_3793);
  and g8171 (n7044, n2569, n7043);
  and g8172 (n7045, n_167, n7044);
  not g8173 (n_3794, n7034);
  and g8174 (n7046, pi0074, n_3794);
  not g8175 (n_3795, n7045);
  and g8176 (n7047, n_3795, n7046);
  and g8177 (n7048, n_3255, n_3787);
  not g8178 (n_3796, n7044);
  not g8179 (n_3797, n7048);
  and g8180 (n7049, n_3796, n_3797);
  not g8181 (n_3798, n7049);
  and g8182 (n7050, pi0054, n_3798);
  and g8183 (n7051, n_171, n7043);
  and g8184 (n7052, pi0075, n_3787);
  not g8185 (n_3799, n7052);
  and g8186 (n7053, pi0092, n_3799);
  not g8187 (n_3800, n7051);
  and g8188 (n7054, n_3800, n7053);
  and g8189 (n7055, pi0075, n7043);
  and g8190 (n7056, pi0087, n7033);
  and g8191 (n7057, n_260, n7033);
  and g8192 (n7058, pi0963, n6745);
  not g8193 (n_3801, n7058);
  and g8194 (n7059, n7036, n_3801);
  and g8195 (n7060, pi0969, n6752);
  not g8196 (n_3802, n7060);
  and g8197 (n7061, n_234, n_3802);
  not g8198 (n_3803, n7059);
  and g8199 (n7062, n2530, n_3803);
  not g8200 (n_3804, n7061);
  and g8201 (n7063, n_3804, n7062);
  not g8202 (n_3805, n7057);
  and g8203 (n7064, pi0100, n_3805);
  not g8204 (n_3806, n7063);
  and g8205 (n7065, n_3806, n7064);
  and g8206 (n7066, n_3580, n7030);
  and g8207 (n7067, n_3578, n7031);
  not g8208 (n_3807, n7066);
  not g8209 (n_3808, n7067);
  and g8210 (n7068, n_3807, n_3808);
  not g8211 (n_3809, n7068);
  and g8212 (n7069, n6767, n_3809);
  and g8213 (n7070, pi0969, n6775);
  not g8214 (n_3810, n7070);
  and g8215 (n7071, n_234, n_3810);
  and g8216 (n7072, n6778, n7018);
  not g8217 (n_3811, n7072);
  and g8218 (n7073, n7036, n_3811);
  not g8219 (n_3812, n7073);
  and g8220 (n7074, n_3593, n_3812);
  and g8221 (n7075, n6786, n7018);
  not g8222 (n_3813, n7075);
  and g8223 (n7076, n_3779, n_3813);
  not g8224 (n_3814, n7076);
  and g8225 (n7077, n6416, n_3814);
  not g8226 (n_3815, n7074);
  not g8227 (n_3816, n7077);
  and g8228 (n7078, n_3815, n_3816);
  not g8229 (n_3817, n7071);
  and g8230 (n7079, pi0232, n_3817);
  not g8231 (n_3818, n7078);
  and g8232 (n7080, n_3818, n7079);
  and g8233 (n7081, pi0969, n6769);
  not g8234 (n_3819, n7081);
  and g8235 (n7082, n_234, n_3819);
  and g8236 (n7083, n_3410, n_3812);
  not g8237 (n_3820, n7082);
  and g8238 (n7084, n_3820, n7083);
  not g8239 (n_3821, n7080);
  not g8240 (n_3822, n7084);
  and g8241 (n7085, n_3821, n_3822);
  not g8242 (n_3823, n7085);
  and g8243 (n7086, n_162, n_3823);
  not g8244 (n_3824, n7069);
  and g8245 (n7087, n_161, n_3824);
  not g8246 (n_3825, n7086);
  and g8247 (n7088, n_3825, n7087);
  and g8248 (n7089, pi0039, n7033);
  not g8249 (n_3826, n7089);
  and g8250 (n7090, pi0038, n_3826);
  not g8251 (n_3827, n7041);
  and g8252 (n7091, n_3827, n7090);
  not g8253 (n_3828, n7088);
  not g8254 (n_3829, n7091);
  and g8255 (n7092, n_3828, n_3829);
  not g8256 (n_3830, n7092);
  and g8257 (n7093, n_164, n_3830);
  not g8258 (n_3831, n7065);
  and g8259 (n7094, n_172, n_3831);
  not g8260 (n_3832, n7093);
  and g8261 (n7095, n_3832, n7094);
  not g8262 (n_3833, n7056);
  and g8263 (n7096, n_171, n_3833);
  not g8264 (n_3834, n7095);
  and g8265 (n7097, n_3834, n7096);
  not g8266 (n_3835, n7055);
  and g8267 (n7098, n_174, n_3835);
  not g8268 (n_3836, n7097);
  and g8269 (n7099, n_3836, n7098);
  not g8270 (n_3837, n7054);
  and g8271 (n7100, n_167, n_3837);
  not g8272 (n_3838, n7099);
  and g8273 (n7101, n_3838, n7100);
  not g8274 (n_3839, n7050);
  and g8275 (n7102, n_168, n_3839);
  not g8276 (n_3840, n7101);
  and g8277 (n7103, n_3840, n7102);
  not g8278 (n_3841, n7047);
  and g8279 (n7104, n_176, n_3841);
  not g8280 (n_3842, n7103);
  and g8281 (n7105, n_3842, n7104);
  not g8282 (n_3843, n7029);
  and g8283 (n7106, n2529, n_3843);
  not g8284 (n_3844, n7105);
  and g8285 (n7107, n_3844, n7106);
  not g8286 (n_3845, n7027);
  and g8287 (n7108, n_792, n_3845);
  not g8288 (n_3846, n7107);
  and g8289 (n7109, n_3846, n7108);
  not g8290 (n_3847, n7026);
  and g8291 (n7110, n_796, n_3847);
  not g8292 (n_3848, n7109);
  and g8293 (n7111, n_3848, n7110);
  not g8294 (n_3849, n7023);
  not g8295 (n_3850, n7111);
  and g8296 (po0176, n_3849, n_3850);
  and g8297 (n7113, pi0975, n6696);
  and g8298 (n7114, n_188, pi0975);
  and g8299 (n7115, n6222, n7114);
  and g8300 (n7116, n2572, n7115);
  and g8301 (n7117, n6305, n7116);
  not g8302 (n_3851, n7113);
  not g8303 (n_3852, n7117);
  and g8304 (n7118, n_3851, n_3852);
  not g8305 (n_3853, n7118);
  and g8306 (n7119, pi0057, n_3853);
  and g8307 (n7120, n6304, n7116);
  and g8308 (n7121, pi0059, n_3851);
  not g8309 (n_3854, n7120);
  and g8310 (n7122, n_3854, n7121);
  and g8311 (n7123, n_3243, n7113);
  and g8312 (n7124, pi0055, n_3851);
  not g8313 (n_3855, n7116);
  and g8314 (n7125, n_3855, n7124);
  and g8315 (n7126, n_234, pi0971);
  and g8316 (n7127, pi0299, pi0975);
  not g8317 (n_3856, n7126);
  not g8318 (n_3857, n7127);
  and g8319 (n7128, n_3856, n_3857);
  not g8320 (n_3858, n7128);
  and g8321 (n7129, n6696, n_3858);
  not g8322 (n_3859, n7129);
  and g8323 (n7130, n_3249, n_3859);
  and g8324 (n7131, n_766, n7129);
  and g8325 (n7132, pi0299, n_3851);
  not g8326 (n_3860, n7115);
  and g8327 (n7133, n_3860, n7132);
  and g8328 (n7134, pi0971, n6720);
  not g8329 (n_3861, n7134);
  and g8330 (n7135, n_234, n_3861);
  not g8331 (n_3862, n7133);
  and g8332 (n7136, n_162, n_3862);
  not g8333 (n_3863, n7135);
  and g8334 (n7137, n_3863, n7136);
  and g8335 (n7138, n2620, n7137);
  not g8336 (n_3864, n7131);
  not g8337 (n_3865, n7138);
  and g8338 (n7139, n_3864, n_3865);
  and g8339 (n7140, n2569, n7139);
  and g8340 (n7141, n_167, n7140);
  not g8341 (n_3866, n7130);
  and g8342 (n7142, pi0074, n_3866);
  not g8343 (n_3867, n7141);
  and g8344 (n7143, n_3867, n7142);
  and g8345 (n7144, n_3255, n_3859);
  not g8346 (n_3868, n7140);
  not g8347 (n_3869, n7144);
  and g8348 (n7145, n_3868, n_3869);
  not g8349 (n_3870, n7145);
  and g8350 (n7146, pi0054, n_3870);
  and g8351 (n7147, n_171, n7139);
  and g8352 (n7148, pi0075, n_3859);
  not g8353 (n_3871, n7148);
  and g8354 (n7149, pi0092, n_3871);
  not g8355 (n_3872, n7147);
  and g8356 (n7150, n_3872, n7149);
  and g8357 (n7151, pi0075, n7139);
  and g8358 (n7152, pi0087, n7129);
  and g8359 (n7153, n_260, n7129);
  and g8360 (n7154, pi0975, n6745);
  not g8361 (n_3873, n7154);
  and g8362 (n7155, n7132, n_3873);
  and g8363 (n7156, pi0971, n6752);
  not g8364 (n_3874, n7156);
  and g8365 (n7157, n_234, n_3874);
  not g8366 (n_3875, n7155);
  and g8367 (n7158, n2530, n_3875);
  not g8368 (n_3876, n7157);
  and g8369 (n7159, n_3876, n7158);
  not g8370 (n_3877, n7153);
  and g8371 (n7160, pi0100, n_3877);
  not g8372 (n_3878, n7159);
  and g8373 (n7161, n_3878, n7160);
  and g8374 (n7162, n_3580, n7126);
  and g8375 (n7163, n_3578, n7127);
  not g8376 (n_3879, n7162);
  not g8377 (n_3880, n7163);
  and g8378 (n7164, n_3879, n_3880);
  not g8379 (n_3881, n7164);
  and g8380 (n7165, n6767, n_3881);
  and g8381 (n7166, pi0971, n6775);
  not g8382 (n_3882, n7166);
  and g8383 (n7167, n_234, n_3882);
  and g8384 (n7168, n6778, n7114);
  not g8385 (n_3883, n7168);
  and g8386 (n7169, n7132, n_3883);
  not g8387 (n_3884, n7169);
  and g8388 (n7170, n_3593, n_3884);
  and g8389 (n7171, n6786, n7114);
  not g8390 (n_3885, n7171);
  and g8391 (n7172, n_3851, n_3885);
  not g8392 (n_3886, n7172);
  and g8393 (n7173, n6416, n_3886);
  not g8394 (n_3887, n7170);
  not g8395 (n_3888, n7173);
  and g8396 (n7174, n_3887, n_3888);
  not g8397 (n_3889, n7167);
  and g8398 (n7175, pi0232, n_3889);
  not g8399 (n_3890, n7174);
  and g8400 (n7176, n_3890, n7175);
  and g8401 (n7177, pi0971, n6769);
  not g8402 (n_3891, n7177);
  and g8403 (n7178, n_234, n_3891);
  and g8404 (n7179, n_3410, n_3884);
  not g8405 (n_3892, n7178);
  and g8406 (n7180, n_3892, n7179);
  not g8407 (n_3893, n7176);
  not g8408 (n_3894, n7180);
  and g8409 (n7181, n_3893, n_3894);
  not g8410 (n_3895, n7181);
  and g8411 (n7182, n_162, n_3895);
  not g8412 (n_3896, n7165);
  and g8413 (n7183, n_161, n_3896);
  not g8414 (n_3897, n7182);
  and g8415 (n7184, n_3897, n7183);
  and g8416 (n7185, pi0039, n7129);
  not g8417 (n_3898, n7185);
  and g8418 (n7186, pi0038, n_3898);
  not g8419 (n_3899, n7137);
  and g8420 (n7187, n_3899, n7186);
  not g8421 (n_3900, n7184);
  not g8422 (n_3901, n7187);
  and g8423 (n7188, n_3900, n_3901);
  not g8424 (n_3902, n7188);
  and g8425 (n7189, n_164, n_3902);
  not g8426 (n_3903, n7161);
  and g8427 (n7190, n_172, n_3903);
  not g8428 (n_3904, n7189);
  and g8429 (n7191, n_3904, n7190);
  not g8430 (n_3905, n7152);
  and g8431 (n7192, n_171, n_3905);
  not g8432 (n_3906, n7191);
  and g8433 (n7193, n_3906, n7192);
  not g8434 (n_3907, n7151);
  and g8435 (n7194, n_174, n_3907);
  not g8436 (n_3908, n7193);
  and g8437 (n7195, n_3908, n7194);
  not g8438 (n_3909, n7150);
  and g8439 (n7196, n_167, n_3909);
  not g8440 (n_3910, n7195);
  and g8441 (n7197, n_3910, n7196);
  not g8442 (n_3911, n7146);
  and g8443 (n7198, n_168, n_3911);
  not g8444 (n_3912, n7197);
  and g8445 (n7199, n_3912, n7198);
  not g8446 (n_3913, n7143);
  and g8447 (n7200, n_176, n_3913);
  not g8448 (n_3914, n7199);
  and g8449 (n7201, n_3914, n7200);
  not g8450 (n_3915, n7125);
  and g8451 (n7202, n2529, n_3915);
  not g8452 (n_3916, n7201);
  and g8453 (n7203, n_3916, n7202);
  not g8454 (n_3917, n7123);
  and g8455 (n7204, n_792, n_3917);
  not g8456 (n_3918, n7203);
  and g8457 (n7205, n_3918, n7204);
  not g8458 (n_3919, n7122);
  and g8459 (n7206, n_796, n_3919);
  not g8460 (n_3920, n7205);
  and g8461 (n7207, n_3920, n7206);
  not g8462 (n_3921, n7119);
  not g8463 (n_3922, n7207);
  and g8464 (po0177, n_3921, n_3922);
  and g8465 (n7209, pi0978, n6696);
  and g8466 (n7210, n_188, pi0978);
  and g8467 (n7211, n2572, n7210);
  and g8468 (n7212, n6222, n7211);
  and g8469 (n7213, n6305, n7212);
  not g8470 (n_3923, n7209);
  not g8471 (n_3924, n7213);
  and g8472 (n7214, n_3923, n_3924);
  not g8473 (n_3925, n7214);
  and g8474 (n7215, pi0057, n_3925);
  and g8475 (n7216, n6304, n7212);
  and g8476 (n7217, pi0059, n_3923);
  not g8477 (n_3926, n7216);
  and g8478 (n7218, n_3926, n7217);
  and g8479 (n7219, n_3243, n7209);
  and g8480 (n7220, pi0055, n_3923);
  not g8481 (n_3927, n7212);
  and g8482 (n7221, n_3927, n7220);
  and g8483 (n7222, n_234, pi0974);
  and g8484 (n7223, pi0299, pi0978);
  not g8485 (n_3928, n7222);
  not g8486 (n_3929, n7223);
  and g8487 (n7224, n_3928, n_3929);
  not g8488 (n_3930, n7224);
  and g8489 (n7225, n6696, n_3930);
  not g8490 (n_3931, n7225);
  and g8491 (n7226, n_3249, n_3931);
  and g8492 (n7227, n6720, n_3930);
  and g8493 (n7228, n_188, n_766);
  not g8494 (n_3932, n7228);
  and g8495 (n7229, n7227, n_3932);
  not g8496 (n_3933, n7229);
  and g8497 (n7230, n2569, n_3933);
  and g8498 (n7231, n_167, n7230);
  not g8499 (n_3934, n7226);
  and g8500 (n7232, pi0074, n_3934);
  not g8501 (n_3935, n7231);
  and g8502 (n7233, n_3935, n7232);
  and g8503 (n7234, n_3255, n_3931);
  not g8504 (n_3936, n7230);
  not g8505 (n_3937, n7234);
  and g8506 (n7235, n_3936, n_3937);
  not g8507 (n_3938, n7235);
  and g8508 (n7236, pi0054, n_3938);
  and g8509 (n7237, n_171, n_3933);
  and g8510 (n7238, pi0075, n_3931);
  not g8511 (n_3939, n7238);
  and g8512 (n7239, pi0092, n_3939);
  not g8513 (n_3940, n7237);
  and g8514 (n7240, n_3940, n7239);
  and g8515 (n7241, pi0075, n_3933);
  and g8516 (n7242, pi0087, n7225);
  and g8517 (n7243, n_260, n7225);
  and g8518 (n7244, pi0299, n_3923);
  and g8519 (n7245, pi0978, n6745);
  not g8520 (n_3941, n7245);
  and g8521 (n7246, n7244, n_3941);
  and g8522 (n7247, pi0974, n6752);
  not g8523 (n_3942, n7247);
  and g8524 (n7248, n_234, n_3942);
  not g8525 (n_3943, n7246);
  and g8526 (n7249, n2530, n_3943);
  not g8527 (n_3944, n7248);
  and g8528 (n7250, n_3944, n7249);
  not g8529 (n_3945, n7243);
  and g8530 (n7251, pi0100, n_3945);
  not g8531 (n_3946, n7250);
  and g8532 (n7252, n_3946, n7251);
  and g8533 (n7253, pi0039, n7225);
  and g8534 (n7254, n_162, n7227);
  not g8535 (n_3947, n7253);
  and g8536 (n7255, pi0038, n_3947);
  not g8537 (n_3948, n7254);
  and g8538 (n7256, n_3948, n7255);
  and g8539 (n7257, n_3580, n7222);
  and g8540 (n7258, n_3578, n7223);
  not g8541 (n_3949, n7257);
  not g8542 (n_3950, n7258);
  and g8543 (n7259, n_3949, n_3950);
  not g8544 (n_3951, n7259);
  and g8545 (n7260, n6767, n_3951);
  and g8546 (n7261, pi0974, n6775);
  not g8547 (n_3952, n7261);
  and g8548 (n7262, n_234, n_3952);
  and g8549 (n7263, n6778, n7210);
  not g8550 (n_3953, n7263);
  and g8551 (n7264, n7244, n_3953);
  not g8552 (n_3954, n7264);
  and g8553 (n7265, n_3593, n_3954);
  and g8554 (n7266, n6786, n7210);
  not g8555 (n_3955, n7266);
  and g8556 (n7267, n_3923, n_3955);
  not g8557 (n_3956, n7267);
  and g8558 (n7268, n6416, n_3956);
  not g8559 (n_3957, n7265);
  not g8560 (n_3958, n7268);
  and g8561 (n7269, n_3957, n_3958);
  not g8562 (n_3959, n7262);
  and g8563 (n7270, pi0232, n_3959);
  not g8564 (n_3960, n7269);
  and g8565 (n7271, n_3960, n7270);
  and g8566 (n7272, pi0974, n6769);
  not g8567 (n_3961, n7272);
  and g8568 (n7273, n_234, n_3961);
  and g8569 (n7274, n_3410, n_3954);
  not g8570 (n_3962, n7273);
  and g8571 (n7275, n_3962, n7274);
  not g8572 (n_3963, n7271);
  not g8573 (n_3964, n7275);
  and g8574 (n7276, n_3963, n_3964);
  not g8575 (n_3965, n7276);
  and g8576 (n7277, n_162, n_3965);
  not g8577 (n_3966, n7260);
  and g8578 (n7278, n_161, n_3966);
  not g8579 (n_3967, n7277);
  and g8580 (n7279, n_3967, n7278);
  not g8581 (n_3968, n7256);
  not g8582 (n_3969, n7279);
  and g8583 (n7280, n_3968, n_3969);
  not g8584 (n_3970, n7280);
  and g8585 (n7281, n_164, n_3970);
  not g8586 (n_3971, n7252);
  and g8587 (n7282, n_172, n_3971);
  not g8588 (n_3972, n7281);
  and g8589 (n7283, n_3972, n7282);
  not g8590 (n_3973, n7242);
  and g8591 (n7284, n_171, n_3973);
  not g8592 (n_3974, n7283);
  and g8593 (n7285, n_3974, n7284);
  not g8594 (n_3975, n7241);
  and g8595 (n7286, n_174, n_3975);
  not g8596 (n_3976, n7285);
  and g8597 (n7287, n_3976, n7286);
  not g8598 (n_3977, n7240);
  and g8599 (n7288, n_167, n_3977);
  not g8600 (n_3978, n7287);
  and g8601 (n7289, n_3978, n7288);
  not g8602 (n_3979, n7236);
  and g8603 (n7290, n_168, n_3979);
  not g8604 (n_3980, n7289);
  and g8605 (n7291, n_3980, n7290);
  not g8606 (n_3981, n7233);
  and g8607 (n7292, n_176, n_3981);
  not g8608 (n_3982, n7291);
  and g8609 (n7293, n_3982, n7292);
  not g8610 (n_3983, n7221);
  and g8611 (n7294, n2529, n_3983);
  not g8612 (n_3984, n7293);
  and g8613 (n7295, n_3984, n7294);
  not g8614 (n_3985, n7219);
  and g8615 (n7296, n_792, n_3985);
  not g8616 (n_3986, n7295);
  and g8617 (n7297, n_3986, n7296);
  not g8618 (n_3987, n7218);
  and g8619 (n7298, n_796, n_3987);
  not g8620 (n_3988, n7297);
  and g8621 (n7299, n_3988, n7298);
  not g8622 (n_3989, n7215);
  not g8623 (n_3990, n7299);
  and g8624 (po0178, n_3989, n_3990);
  and g8625 (n7301, n2620, n6284);
  not g8626 (n_3991, n7301);
  and g8627 (n7302, pi0075, n_3991);
  and g8628 (n7303, n2533, n2608);
  and g8629 (n7304, n6284, n7303);
  not g8630 (n_3992, n7304);
  and g8631 (n7305, pi0092, n_3992);
  not g8632 (n_3993, n7302);
  not g8633 (n_3994, n7305);
  and g8634 (n7306, n_3993, n_3994);
  and g8635 (n7307, pi0299, n_3164);
  and g8636 (n7308, n6759, n7307);
  and g8637 (n7309, n_234, n_3122);
  and g8638 (n7310, n6409, n7309);
  not g8639 (n_3995, n7310);
  and g8640 (n7311, pi0039, n_3995);
  not g8641 (n_3996, n7308);
  and g8642 (n7312, n_3996, n7311);
  and g8643 (n7313, pi0299, n6489);
  and g8644 (n7314, n_234, n6520);
  not g8645 (n_3997, n7313);
  and g8646 (n7315, n_3410, n_3997);
  not g8647 (n_3998, n7314);
  and g8648 (n7316, n_3998, n7315);
  and g8649 (n7317, n6527, n6532);
  not g8654 (n_4000, n6416);
  and g8655 (n7321, n_4000, n7313);
  and g8656 (n7322, n_3378, n6781);
  not g8657 (n_4001, n6785);
  and g8658 (n7323, n_4001, n7322);
  not g8665 (n_4005, n7316);
  and g8666 (n7327, n_162, n_4005);
  not g8667 (n_4006, n7326);
  and g8668 (n7328, n_4006, n7327);
  not g8669 (n_4007, n7312);
  not g8670 (n_4008, n7328);
  and g8671 (n7329, n_4007, n_4008);
  not g8672 (n_4009, n7329);
  and g8673 (n7330, n_161, n_4009);
  not g8674 (n_4010, n7330);
  and g8675 (n7331, n_3039, n_4010);
  not g8676 (n_4011, n7331);
  and g8677 (n7332, n_164, n_4011);
  and g8678 (n7333, n_161, n6284);
  not g8679 (n_4012, n7333);
  and g8680 (n7334, pi0100, n_4012);
  not g8681 (n_4013, n7334);
  and g8682 (n7335, n6289, n_4013);
  not g8683 (n_4014, n7332);
  and g8684 (n7336, n_4014, n7335);
  not g8685 (n_4015, n7336);
  and g8686 (n7337, n2569, n_4015);
  not g8687 (n_4016, n7337);
  and g8688 (n7338, n7306, n_4016);
  not g8689 (n_4017, n7338);
  and g8690 (n7339, n_167, n_4017);
  and g8691 (n7340, n_174, n7304);
  not g8692 (n_4018, n7340);
  and g8693 (n7341, pi0054, n_4018);
  not g8694 (n_4019, n7339);
  not g8695 (n_4020, n7341);
  and g8696 (n7342, n_4019, n_4020);
  not g8697 (n_4021, n7342);
  and g8698 (n7343, n_168, n_4021);
  not g8699 (n_4022, n7343);
  and g8700 (n7344, n_3035, n_4022);
  not g8701 (n_4023, n7344);
  and g8702 (n7345, n_176, n_4023);
  and g8703 (n7346, n2535, n6125);
  not g8704 (n_4024, n7346);
  and g8705 (n7347, pi0055, n_4024);
  not g8706 (n_4025, n7347);
  and g8707 (n7348, n_157, n_4025);
  and g8708 (n7349, n_158, n7348);
  not g8709 (n_4026, n7345);
  and g8710 (n7350, n_4026, n7349);
  not g8711 (n_4027, n7350);
  and g8712 (n7351, n3328, n_4027);
  not g8713 (n_4028, n7351);
  and g8714 (po0195, n6123, n_4028);
  not g8715 (po1110, pi0954);
  not g8716 (n_4032, po0195);
  and g8717 (n7353, po1110, n_4032);
  and g8718 (n7354, pi0024, pi0954);
  not g8719 (n_4034, n7353);
  not g8720 (n_4035, n7354);
  and g8721 (po0182, n_4034, n_4035);
  and g8722 (n7356, n2531, n3335);
  and g8723 (n7357, n3330, n7356);
  not g8724 (n_4036, n7357);
  and g8725 (n7358, n_19, n_4036);
  not g8726 (n_4037, n7358);
  and g8727 (n7359, pi0062, n_4037);
  and g8728 (n7360, n2537, n3335);
  and g8729 (n7361, pi0056, n_19);
  not g8730 (n_4038, n7360);
  and g8731 (n7362, n_4038, n7361);
  and g8732 (n7363, n2531, n6128);
  and g8733 (n7364, n3335, n7363);
  and g8734 (n7365, n_168, n7364);
  not g8735 (n_4039, n7365);
  and g8736 (n7366, n_19, n_4039);
  not g8737 (n_4040, n7366);
  and g8738 (n7367, pi0055, n_4040);
  and g8739 (n7368, n_19, n_841);
  and g8740 (n7369, n3335, n3373);
  not g8741 (n_4041, n7369);
  and g8742 (n7370, n_19, n_4041);
  not g8743 (n_4042, n7370);
  and g8744 (n7371, pi0092, n_4042);
  and g8745 (n7372, pi0075, n_19);
  not g8746 (n_4043, n7356);
  and g8747 (n7373, n_19, n_4043);
  not g8748 (n_4044, n7373);
  and g8749 (n7374, pi0087, n_4044);
  and g8750 (n7375, n_164, n4730);
  not g8751 (n_4045, n6356);
  and g8752 (n7376, n2521, n_4045);
  not g8753 (n_4046, n7376);
  and g8754 (n7377, n_234, n_4046);
  and g8755 (n7378, pi0299, n_1567);
  not g8756 (n_4047, n7377);
  not g8757 (n_4048, n7378);
  and g8758 (n7379, n_4047, n_4048);
  and g8759 (n7380, pi0100, n3335);
  and g8760 (n7381, n7379, n7380);
  not g8761 (n_4049, n7381);
  and g8762 (n7382, n_162, n_4049);
  not g8763 (n_4050, n7375);
  and g8764 (n7383, n_4050, n7382);
  and g8765 (n7384, n_164, n3335);
  not g8766 (n_4051, n7384);
  and g8767 (n7385, pi0039, n_4051);
  not g8768 (n_4052, n7385);
  and g8769 (n7386, n_161, n_4052);
  not g8770 (n_4053, n7383);
  and g8771 (n7387, n_4053, n7386);
  not g8772 (n_4054, n7387);
  and g8773 (n7388, n_19, n_4054);
  not g8774 (n_4055, n7388);
  and g8775 (n7389, n_172, n_4055);
  not g8776 (n_4056, n7374);
  and g8777 (n7390, n_171, n_4056);
  not g8778 (n_4057, n7389);
  and g8779 (n7391, n_4057, n7390);
  not g8780 (n_4058, n7372);
  and g8781 (n7392, n_174, n_4058);
  not g8782 (n_4059, n7391);
  and g8783 (n7393, n_4059, n7392);
  not g8784 (n_4060, n7371);
  and g8785 (n7394, n2532, n_4060);
  not g8786 (n_4061, n7393);
  and g8787 (n7395, n_4061, n7394);
  not g8788 (n_4062, n7368);
  and g8789 (n7396, n_176, n_4062);
  not g8790 (n_4063, n7395);
  and g8791 (n7397, n_4063, n7396);
  not g8792 (n_4064, n7367);
  and g8793 (n7398, n_157, n_4064);
  not g8794 (n_4065, n7397);
  and g8795 (n7399, n_4065, n7398);
  not g8796 (n_4066, n7362);
  and g8797 (n7400, n_158, n_4066);
  not g8798 (n_4067, n7399);
  and g8799 (n7401, n_4067, n7400);
  not g8800 (n_4068, n7359);
  not g8801 (n_4069, n7401);
  and g8802 (n7402, n_4068, n_4069);
  not g8803 (n_4070, n7402);
  and g8804 (n7403, n3328, n_4070);
  and g8805 (n7404, n2441, n_824);
  or g8806 (po0183, n7403, n7404);
  and g8807 (n7406, pi0119, pi1056);
  and g8808 (n7407, n_188, pi0252);
  not g8809 (n_4073, pi0119);
  not g8810 (n_4074, n7407);
  and g8811 (n7408, n_4073, n_4074);
  not g8812 (n_4075, n7408);
  and g8813 (n7409, n_3100, n_4075);
  not g8814 (n_4076, n7409);
  or g8815 (po0184, n7406, n_4076);
  and g8816 (n7411, pi0119, pi1077);
  or g8817 (po0185, n_4076, n7411);
  and g8818 (n7413, pi0119, pi1073);
  or g8819 (po0186, n_4076, n7413);
  and g8820 (n7415, pi0119, pi1041);
  or g8821 (po0187, n_4076, n7415);
  and g8822 (n7417, pi0824, n2932);
  not g8823 (n_4081, pi0122);
  and g8824 (n7418, n_4081, pi1093);
  and g8825 (n7419, n7417, n7418);
  and g8826 (n7420, n_3128, n7419);
  and g8827 (n7421, n_47, n7420);
  and g8828 (n7422, pi0567, n7421);
  not g8829 (n_4085, pi0285);
  not g8830 (n_4086, pi0286);
  and g8831 (n7423, n_4085, n_4086);
  not g8832 (n_4088, pi0289);
  and g8833 (n7424, n_4088, n7423);
  not g8834 (n_4090, pi0288);
  and g8835 (n7425, n_4090, n7424);
  or g8836 (po1038, pi0057, n_3232);
  not g8837 (n_4091, n7425);
  and g8838 (n7427, n_4091, po1038);
  and g8839 (n7428, n7422, n7427);
  and g8840 (n7429, n_168, n6134);
  and g8841 (n7430, n_4081, pi0829);
  and g8842 (n7431, n2961, n_3055);
  and g8843 (n7432, n_3052, n2703);
  and g8844 (n7433, pi0090, n7432);
  not g8845 (n_4093, n7433);
  and g8846 (n7434, n_131, n_4093);
  not g8847 (n_4094, n7434);
  and g8848 (n7435, n7431, n_4094);
  not g8849 (n_4095, n7435);
  and g8850 (n7436, n_138, n_4095);
  and g8851 (n7437, n_46, pi0098);
  and g8852 (n7438, n_51, n_49);
  and g8853 (n7439, n_125, n7438);
  and g8854 (n7440, n2767, n7439);
  and g8855 (n7441, n2495, n7437);
  and g8856 (n7442, n7440, n7441);
  not g8857 (n_4096, n7442);
  and g8858 (n7443, n_122, n_4096);
  not g8859 (n_4097, n7443);
  and g8860 (n7444, n2717, n_4097);
  and g8861 (n7445, n_130, n2704);
  and g8862 (n7446, n_139, n7445);
  and g8863 (n7447, n7444, n7446);
  not g8864 (n_4098, n7447);
  and g8865 (n7448, n7436, n_4098);
  not g8866 (n_4099, n7448);
  and g8867 (n7449, n_350, n_4099);
  and g8868 (n7450, n_135, n2519);
  and g8869 (n7451, n7449, n7450);
  and g8870 (n7452, n6277, n7451);
  not g8871 (n_4100, n7430);
  and g8872 (n7453, n_4100, n7452);
  not g8873 (n_4101, n7449);
  and g8874 (n7454, n_135, n_4101);
  not g8875 (n_4102, n6484);
  and g8876 (n7455, pi0096, n_4102);
  not g8877 (n_4103, n7455);
  and g8878 (n7456, n2519, n_4103);
  and g8879 (n7457, n2932, n7430);
  and g8880 (n7458, n7456, n7457);
  not g8881 (n_4104, n7454);
  and g8882 (n7459, n_4104, n7458);
  not g8883 (n_4105, n7453);
  not g8884 (n_4106, n7459);
  and g8885 (n7460, n_4105, n_4106);
  not g8886 (n_4107, n7460);
  and g8887 (n7461, n_3206, n_4107);
  not g8888 (n_4108, n7461);
  and g8889 (n7462, n_172, n_4108);
  and g8890 (n7463, n2521, po0740);
  not g8891 (n_4109, n7463);
  and g8892 (n7464, pi0087, n_4109);
  and g8893 (n7465, n_171, n2531);
  not g8894 (n_4110, n7464);
  and g8895 (n7466, n_4110, n7465);
  not g8896 (n_4111, n7462);
  and g8897 (n7467, n_4111, n7466);
  not g8898 (n_4112, pi0567);
  not g8899 (n_4113, n7467);
  and g8900 (n7468, n_4112, n_4113);
  not g8901 (n_4114, n7468);
  and g8902 (n7469, n7429, n_4114);
  and g8903 (n7470, n_234, n_302);
  and g8904 (n7471, pi0299, n_269);
  not g8905 (n_4115, n7470);
  not g8906 (n_4116, n7471);
  and g8907 (n7472, n_4115, n_4116);
  and g8908 (n7473, pi0232, n6197);
  and g8909 (n7474, n7472, n7473);
  not g8910 (n_4117, n7474);
  and g8911 (n7475, n2610, n_4117);
  not g8912 (n_4118, n7475);
  and g8913 (n7476, n7421, n_4118);
  not g8914 (n_4119, pi0024);
  and g8915 (n7477, n_4119, n6359);
  and g8916 (n7478, n_489, po1057);
  and g8917 (n7479, pi1093, n7457);
  and g8918 (n7480, n7478, n7479);
  and g8919 (n7481, n7477, n7480);
  not g8920 (n_4120, n7481);
  and g8921 (n7482, pi1091, n_4120);
  not g8922 (n_4121, n7482);
  and g8923 (n7483, n7475, n_4121);
  and g8924 (n7484, n_47, n7417);
  and g8925 (n7485, n7418, n7484);
  not g8926 (n_4122, n7485);
  and g8927 (n7486, n_3128, n_4122);
  not g8928 (n_4123, n7486);
  and g8929 (n7487, n7483, n_4123);
  not g8930 (n_4124, n7476);
  and g8931 (n7488, pi0075, n_4124);
  not g8932 (n_4125, n7487);
  and g8933 (n7489, n_4125, n7488);
  and g8934 (n7490, pi1093, n2923);
  not g8935 (n_4126, n7490);
  and g8936 (n7491, n6277, n_4126);
  and g8937 (n7492, n2521, n7491);
  not g8938 (n_4127, n7492);
  and g8939 (n7493, pi1091, n_4127);
  and g8940 (n7494, n_3128, n_4109);
  and g8941 (n7495, n2521, n7417);
  and g8942 (n7496, pi0122, n7495);
  and g8943 (n7497, n_4081, n7484);
  not g8944 (n_4128, n7496);
  not g8945 (n_4129, n7497);
  and g8946 (n7498, n_4128, n_4129);
  not g8947 (n_4130, n7498);
  and g8948 (n7499, pi1093, n_4130);
  not g8949 (n_4131, n7499);
  and g8950 (n7500, n7494, n_4131);
  not g8951 (n_4132, n7493);
  and g8952 (n7501, n2625, n_4132);
  not g8953 (n_4133, n7500);
  and g8954 (n7502, n_4133, n7501);
  not g8955 (n_4134, n7421);
  not g8956 (n_4135, n7502);
  and g8957 (n7503, n_4134, n_4135);
  not g8958 (n_4136, n7503);
  and g8959 (n7504, pi0087, n_4136);
  and g8960 (n7505, n_260, n7421);
  and g8961 (n7506, pi0228, n_4117);
  not g8962 (n_4137, n7506);
  and g8963 (n7507, n_4134, n_4137);
  and g8964 (n7508, n2521, n7480);
  not g8965 (n_4138, n7508);
  and g8966 (n7509, pi1091, n_4138);
  not g8967 (n_4139, n7509);
  and g8968 (n7510, n_4123, n_4139);
  not g8969 (n_4140, n7510);
  and g8970 (n7511, n7506, n_4140);
  not g8971 (n_4141, n7507);
  and g8972 (n7512, n2530, n_4141);
  not g8973 (n_4142, n7511);
  and g8974 (n7513, n_4142, n7512);
  not g8975 (n_4143, n7505);
  and g8976 (n7514, pi0100, n_4143);
  not g8977 (n_4144, n7513);
  and g8978 (n7515, n_4144, n7514);
  and g8979 (n7516, pi0038, n7421);
  and g8980 (n7517, pi1093, n_489);
  and g8981 (n7518, n_350, n7450);
  not g8982 (n_4145, n7436);
  and g8983 (n7519, n_4145, n7518);
  and g8984 (n7520, n7417, n7519);
  and g8985 (n7521, n_3127, n7520);
  and g8986 (n7522, n_4119, n2756);
  and g8991 (n7527, n_109, n7526);
  not g8992 (n_4146, n7522);
  not g8993 (n_4147, n7527);
  and g8994 (n7528, n_4146, n_4147);
  and g8995 (n7529, n2461, n7431);
  not g8996 (n_4148, n7528);
  and g8997 (n7530, n_4148, n7529);
  not g8998 (n_4149, n7530);
  and g8999 (n7531, n7436, n_4149);
  not g9000 (n_4150, n7531);
  and g9001 (n7532, n_350, n_4150);
  not g9002 (n_4151, n7532);
  and g9003 (n7533, n_135, n_4151);
  and g9004 (n7534, n2933, n7456);
  not g9005 (n_4152, n7533);
  and g9006 (n7535, n_4152, n7534);
  not g9007 (n_4153, n7521);
  not g9008 (n_4154, n7535);
  and g9009 (n7536, n_4153, n_4154);
  not g9010 (n_4155, n7536);
  and g9011 (n7537, n_4081, n_4155);
  and g9012 (n7538, pi0122, n6277);
  and g9013 (n7539, n7519, n7538);
  not g9014 (n_4156, n7537);
  not g9015 (n_4157, n7539);
  and g9016 (n7540, n_4156, n_4157);
  not g9017 (n_4158, n7540);
  and g9018 (n7541, n7517, n_4158);
  not g9019 (n_4159, n7541);
  and g9020 (n7542, pi1091, n_4159);
  and g9021 (n7543, n_4108, n7542);
  not g9022 (n_4160, n7543);
  and g9023 (n7544, n_162, n_4160);
  and g9024 (n7545, n_3128, n_4108);
  and g9025 (n7546, pi0122, n7520);
  not g9026 (n_4161, n7546);
  and g9027 (n7547, n_4129, n_4161);
  not g9028 (n_4162, n7547);
  and g9029 (n7548, pi1093, n_4162);
  not g9030 (n_4163, n7548);
  and g9031 (n7549, n7545, n_4163);
  not g9032 (n_4164, n7549);
  and g9033 (n7550, n7544, n_4164);
  and g9034 (n7551, n_223, n5810);
  not g9035 (n_4165, n7551);
  and g9036 (n7552, n7421, n_4165);
  and g9037 (n7553, n_489, n2925);
  and g9038 (n7554, n6382, n7553);
  and g9039 (n7555, n2926, n7554);
  not g9040 (n_4166, n7555);
  and g9041 (n7556, pi1091, n_4166);
  not g9042 (n_4167, n7556);
  and g9043 (n7557, n_4123, n_4167);
  and g9044 (n7558, n6198, n7557);
  and g9045 (n7559, n_3120, n7421);
  not g9046 (n_4168, n7558);
  not g9047 (n_4169, n7559);
  and g9048 (n7560, n_4168, n_4169);
  and g9049 (n7561, n6205, n7560);
  and g9050 (n7562, n_3140, n7557);
  and g9051 (n7563, n6227, n7421);
  not g9052 (n_4170, n7562);
  not g9053 (n_4171, n7563);
  and g9054 (n7564, n_4170, n_4171);
  and g9055 (n7565, n_3119, n7564);
  not g9056 (n_4172, n7561);
  and g9057 (n7566, n7551, n_4172);
  not g9058 (n_4173, n7565);
  and g9059 (n7567, n_4173, n7566);
  not g9060 (n_4174, n7552);
  and g9061 (n7568, n_234, n_4174);
  not g9062 (n_4175, n7567);
  and g9063 (n7569, n_4175, n7568);
  and g9064 (n7570, n_20, n6379);
  not g9065 (n_4176, n7570);
  and g9066 (n7571, n7421, n_4176);
  and g9067 (n7572, n6242, n7560);
  and g9068 (n7573, n_3162, n7564);
  not g9069 (n_4177, n7572);
  and g9070 (n7574, n7570, n_4177);
  not g9071 (n_4178, n7573);
  and g9072 (n7575, n_4178, n7574);
  not g9073 (n_4179, n7571);
  and g9074 (n7576, pi0299, n_4179);
  not g9075 (n_4180, n7575);
  and g9076 (n7577, n_4180, n7576);
  not g9077 (n_4181, n7569);
  and g9078 (n7578, pi0039, n_4181);
  not g9079 (n_4182, n7577);
  and g9080 (n7579, n_4182, n7578);
  not g9081 (n_4183, n7550);
  not g9082 (n_4184, n7579);
  and g9083 (n7580, n_4183, n_4184);
  not g9084 (n_4185, n7580);
  and g9085 (n7581, n_161, n_4185);
  not g9086 (n_4186, n7516);
  and g9087 (n7582, n_164, n_4186);
  not g9088 (n_4187, n7581);
  and g9089 (n7583, n_4187, n7582);
  not g9090 (n_4188, n7515);
  and g9091 (n7584, n_172, n_4188);
  not g9092 (n_4189, n7583);
  and g9093 (n7585, n_4189, n7584);
  not g9094 (n_4190, n7504);
  and g9095 (n7586, n_171, n_4190);
  not g9096 (n_4191, n7585);
  and g9097 (n7587, n_4191, n7586);
  not g9098 (n_4192, n7489);
  not g9099 (n_4193, n7587);
  and g9100 (n7588, n_4192, n_4193);
  not g9101 (n_4194, n7588);
  and g9102 (n7589, pi0567, n_4194);
  not g9103 (n_4195, n7589);
  and g9104 (n7590, n7469, n_4195);
  not g9105 (n_4196, n7429);
  and g9106 (n7591, n7422, n_4196);
  not g9107 (n_4197, n7590);
  not g9108 (n_4198, n7591);
  and g9109 (n7592, n_4197, n_4198);
  and g9110 (n7593, n_4091, n7592);
  and g9111 (n7594, pi1091, n7478);
  and g9112 (n7595, n7457, n7594);
  and g9113 (n7596, n7477, n7595);
  and g9114 (n7597, pi1093, n7596);
  and g9115 (n7598, n7475, n7597);
  not g9116 (n_4199, n7598);
  and g9117 (n7599, pi0075, n_4199);
  not g9118 (n_4200, n7545);
  and g9119 (n7600, n_4160, n_4200);
  not g9120 (n_4201, n7600);
  and g9121 (n7601, n_162, n_4201);
  and g9122 (n7602, pi1091, n7555);
  and g9123 (n7603, n_3164, n7602);
  and g9124 (n7604, n_20, n6640);
  and g9125 (n7605, n7603, n7604);
  and g9126 (n7606, n_3122, n7602);
  and g9127 (n7607, n_234, n6405);
  and g9128 (n7608, n_219, n7607);
  and g9129 (n7609, n7606, n7608);
  not g9130 (n_4202, n7605);
  and g9131 (n7610, pi0039, n_4202);
  not g9132 (n_4203, n7609);
  and g9133 (n7611, n_4203, n7610);
  not g9134 (n_4204, n7611);
  and g9135 (n7612, n_161, n_4204);
  not g9136 (n_4205, n7601);
  and g9137 (n7613, n_4205, n7612);
  not g9138 (n_4206, n7613);
  and g9139 (n7614, n_164, n_4206);
  not g9144 (n_4208, n7617);
  and g9145 (n7618, n7614, n_4208);
  and g9146 (n7619, pi1091, n7508);
  and g9147 (n7620, pi0228, n7619);
  and g9148 (n7621, n2530, n_4117);
  and g9149 (n7622, n7620, n7621);
  not g9150 (n_4209, n7622);
  and g9151 (n7623, pi0100, n_4209);
  not g9152 (n_4210, n7618);
  not g9153 (n_4211, n7623);
  and g9154 (n7624, n_4210, n_4211);
  not g9155 (n_4212, n7624);
  and g9156 (n7625, n_172, n_4212);
  and g9157 (n7626, n_3128, pi1093);
  not g9158 (n_4213, n7495);
  and g9159 (n7627, n_4213, n7626);
  not g9160 (n_4214, n7626);
  and g9161 (n7628, n_4127, n_4214);
  not g9162 (n_4215, n7628);
  and g9163 (n7629, n2625, n_4215);
  not g9164 (n_4216, n7627);
  and g9165 (n7630, n_4216, n7629);
  not g9166 (n_4217, n7630);
  and g9167 (n7631, pi0087, n_4217);
  not g9168 (n_4218, n7625);
  not g9169 (n_4219, n7631);
  and g9170 (n7632, n_4218, n_4219);
  not g9171 (n_4220, n7632);
  and g9172 (n7633, n_171, n_4220);
  not g9173 (n_4221, n7599);
  not g9174 (n_4222, n7633);
  and g9175 (n7634, n_4221, n_4222);
  not g9176 (n_4223, n7634);
  and g9177 (n7635, pi0567, n_4223);
  not g9178 (n_4224, n7635);
  and g9179 (n7636, n7469, n_4224);
  not g9180 (n_4225, n7636);
  and g9181 (n7637, n7425, n_4225);
  not g9182 (n_4226, po1038);
  not g9183 (n_4227, n7593);
  and g9184 (n7638, n_4226, n_4227);
  not g9185 (n_4228, n7637);
  and g9186 (n7639, n_4228, n7638);
  not g9187 (n_4230, n7428);
  and g9188 (n7640, pi0217, n_4230);
  not g9189 (n_4231, n7639);
  and g9190 (n7641, n_4231, n7640);
  not g9191 (n_4234, pi1161);
  not g9192 (n_4235, pi1162);
  and g9193 (n7642, n_4234, n_4235);
  not g9194 (n_4237, pi1163);
  and g9195 (n7643, n_4237, n7642);
  not g9196 (n_4239, pi0592);
  and g9197 (n7644, n_4239, n7422);
  and g9198 (n7645, pi0592, n7422);
  not g9199 (n_4242, pi0363);
  not g9200 (n_4243, pi0372);
  and g9201 (n7646, n_4242, n_4243);
  and g9202 (n7647, pi0363, pi0372);
  not g9203 (n_4244, n7646);
  not g9204 (n_4245, n7647);
  and g9205 (n7648, n_4244, n_4245);
  not g9206 (n_4247, n7648);
  and g9207 (n7649, pi0386, n_4247);
  not g9208 (n_4248, pi0386);
  and g9209 (n7650, n_4248, n7648);
  not g9210 (n_4249, n7649);
  not g9211 (n_4250, n7650);
  and g9212 (n7651, n_4249, n_4250);
  not g9213 (n_4253, pi0388);
  and g9214 (n7652, pi0338, n_4253);
  not g9215 (n_4254, pi0338);
  and g9216 (n7653, n_4254, pi0388);
  not g9217 (n_4255, n7652);
  not g9218 (n_4256, n7653);
  and g9219 (n7654, n_4255, n_4256);
  not g9220 (n_4259, pi0339);
  and g9221 (n7655, pi0337, n_4259);
  not g9222 (n_4260, pi0337);
  and g9223 (n7656, n_4260, pi0339);
  not g9224 (n_4261, n7655);
  not g9225 (n_4262, n7656);
  and g9226 (n7657, n_4261, n_4262);
  and g9227 (n7658, pi0387, n7657);
  not g9228 (n_4264, pi0387);
  not g9229 (n_4265, n7657);
  and g9230 (n7659, n_4264, n_4265);
  not g9231 (n_4266, n7658);
  not g9232 (n_4267, n7659);
  and g9233 (n7660, n_4266, n_4267);
  not g9234 (n_4269, n7660);
  and g9235 (n7661, pi0380, n_4269);
  not g9236 (n_4270, pi0380);
  and g9237 (n7662, n_4270, n7660);
  not g9238 (n_4271, n7661);
  not g9239 (n_4272, n7662);
  and g9240 (n7663, n_4271, n_4272);
  not g9241 (n_4273, n7663);
  and g9242 (n7664, n7654, n_4273);
  not g9243 (n_4274, n7654);
  and g9244 (n7665, n_4274, n7663);
  not g9245 (n_4275, n7664);
  not g9246 (n_4276, n7665);
  and g9247 (n7666, n_4275, n_4276);
  and g9248 (n7667, n7651, n7666);
  not g9249 (n_4277, n7651);
  not g9250 (n_4278, n7666);
  and g9251 (n7668, n_4277, n_4278);
  not g9252 (n_4279, n7667);
  not g9253 (n_4280, n7668);
  and g9254 (n7669, n_4279, n_4280);
  not g9255 (n_4282, n7669);
  and g9256 (n7670, pi1196, n_4282);
  not g9257 (n_4285, pi0368);
  not g9258 (n_4286, pi0389);
  and g9259 (n7671, n_4285, n_4286);
  and g9260 (n7672, pi0368, pi0389);
  not g9261 (n_4287, n7671);
  not g9262 (n_4288, n7672);
  and g9263 (n7673, n_4287, n_4288);
  not g9264 (n_4291, pi0447);
  and g9265 (n7674, pi0365, n_4291);
  not g9266 (n_4292, pi0365);
  and g9267 (n7675, n_4292, pi0447);
  not g9268 (n_4293, n7674);
  not g9269 (n_4294, n7675);
  and g9270 (n7676, n_4293, n_4294);
  not g9271 (n_4297, pi0383);
  and g9272 (n7677, pi0336, n_4297);
  not g9273 (n_4298, pi0336);
  and g9274 (n7678, n_4298, pi0383);
  not g9275 (n_4299, n7677);
  not g9276 (n_4300, n7678);
  and g9277 (n7679, n_4299, n_4300);
  not g9278 (n_4303, pi0366);
  and g9279 (n7680, pi0364, n_4303);
  not g9280 (n_4304, pi0364);
  and g9281 (n7681, n_4304, pi0366);
  not g9282 (n_4305, n7680);
  not g9283 (n_4306, n7681);
  and g9284 (n7682, n_4305, n_4306);
  and g9285 (n7683, n7679, n7682);
  not g9286 (n_4307, n7679);
  not g9287 (n_4308, n7682);
  and g9288 (n7684, n_4307, n_4308);
  not g9289 (n_4309, n7683);
  not g9290 (n_4310, n7684);
  and g9291 (n7685, n_4309, n_4310);
  and g9292 (n7686, n7676, n7685);
  not g9293 (n_4311, n7676);
  not g9294 (n_4312, n7685);
  and g9295 (n7687, n_4311, n_4312);
  not g9296 (n_4313, n7686);
  not g9297 (n_4314, n7687);
  and g9298 (n7688, n_4313, n_4314);
  not g9299 (n_4316, n7688);
  and g9300 (n7689, pi0367, n_4316);
  not g9301 (n_4317, pi0367);
  and g9302 (n7690, n_4317, n7688);
  not g9303 (n_4318, n7689);
  not g9304 (n_4319, n7690);
  and g9305 (n7691, n_4318, n_4319);
  and g9306 (n7692, n7673, n7691);
  not g9307 (n_4320, n7673);
  not g9308 (n_4321, n7691);
  and g9309 (n7693, n_4320, n_4321);
  not g9310 (n_4323, n7692);
  and g9311 (n7694, pi1197, n_4323);
  not g9312 (n_4324, n7693);
  and g9313 (n7695, n_4324, n7694);
  not g9314 (n_4325, n7670);
  not g9315 (n_4326, n7695);
  and g9316 (n7696, n_4325, n_4326);
  not g9317 (n_4327, n7696);
  and g9318 (n7697, pi0592, n_4327);
  not g9319 (n_4330, pi0382);
  and g9320 (n7698, pi0379, n_4330);
  not g9321 (n_4331, pi0379);
  and g9322 (n7699, n_4331, pi0382);
  not g9323 (n_4332, n7698);
  not g9324 (n_4333, n7699);
  and g9325 (n7700, n_4332, n_4333);
  not g9326 (n_4336, pi0439);
  and g9327 (n7701, pi0376, n_4336);
  not g9328 (n_4337, pi0376);
  and g9329 (n7702, n_4337, pi0439);
  not g9330 (n_4338, n7701);
  not g9331 (n_4339, n7702);
  and g9332 (n7703, n_4338, n_4339);
  and g9333 (n7704, pi0381, n7703);
  not g9334 (n_4341, pi0381);
  not g9335 (n_4342, n7703);
  and g9336 (n7705, n_4341, n_4342);
  not g9337 (n_4343, n7704);
  not g9338 (n_4344, n7705);
  and g9339 (n7706, n_4343, n_4344);
  not g9340 (n_4347, pi0385);
  and g9341 (n7707, pi0317, n_4347);
  not g9342 (n_4348, pi0317);
  and g9343 (n7708, n_4348, pi0385);
  not g9344 (n_4349, n7707);
  not g9345 (n_4350, n7708);
  and g9346 (n7709, n_4349, n_4350);
  and g9347 (n7710, pi0378, n7709);
  not g9348 (n_4352, pi0378);
  not g9349 (n_4353, n7709);
  and g9350 (n7711, n_4352, n_4353);
  not g9351 (n_4354, n7710);
  not g9352 (n_4355, n7711);
  and g9353 (n7712, n_4354, n_4355);
  not g9354 (n_4356, n7712);
  and g9355 (n7713, n7706, n_4356);
  not g9356 (n_4357, n7706);
  and g9357 (n7714, n_4357, n7712);
  not g9358 (n_4358, n7713);
  not g9359 (n_4359, n7714);
  and g9360 (n7715, n_4358, n_4359);
  and g9361 (n7716, n7700, n7715);
  not g9362 (n_4360, n7700);
  not g9363 (n_4361, n7715);
  and g9364 (n7717, n_4360, n_4361);
  not g9365 (n_4362, n7716);
  not g9366 (n_4363, n7717);
  and g9367 (n7718, n_4362, n_4363);
  not g9368 (n_4365, pi0377);
  not g9369 (n_4366, n7718);
  and g9370 (n7719, n_4365, n_4366);
  and g9371 (n7720, pi0377, n7718);
  not g9372 (n_4367, n7719);
  not g9373 (n_4368, n7720);
  and g9374 (n7721, n_4367, n_4368);
  not g9375 (n_4369, n7721);
  and g9376 (n7722, n7696, n_4369);
  not g9377 (n_4370, n7722);
  and g9378 (n7723, pi0592, n_4370);
  not g9379 (n_4371, n7723);
  and g9380 (n7724, n7422, n_4371);
  not g9381 (n_4373, n7724);
  and g9382 (n7725, pi1199, n_4373);
  not g9383 (n_4374, n7697);
  not g9384 (n_4375, n7725);
  and g9385 (n7726, n_4374, n_4375);
  and g9386 (n7727, n7645, n7726);
  not g9387 (n_4377, pi1198);
  and g9388 (n7728, n_4377, n7727);
  not g9389 (n_4380, pi0442);
  and g9390 (n7729, pi0384, n_4380);
  not g9391 (n_4381, pi0384);
  and g9392 (n7730, n_4381, pi0442);
  not g9393 (n_4382, n7729);
  not g9394 (n_4383, n7730);
  and g9395 (n7731, n_4382, n_4383);
  not g9396 (n_4385, n7731);
  and g9397 (n7732, pi0440, n_4385);
  not g9398 (n_4386, pi0440);
  and g9399 (n7733, n_4386, n7731);
  not g9400 (n_4387, n7732);
  not g9401 (n_4388, n7733);
  and g9402 (n7734, n_4387, n_4388);
  not g9403 (n_4391, pi0369);
  not g9404 (n_4392, pi0374);
  and g9405 (n7735, n_4391, n_4392);
  and g9406 (n7736, pi0369, pi0374);
  not g9407 (n_4393, n7735);
  not g9408 (n_4394, n7736);
  and g9409 (n7737, n_4393, n_4394);
  not g9410 (n_4396, pi0370);
  not g9411 (n_4397, n7737);
  and g9412 (n7738, n_4396, n_4397);
  and g9413 (n7739, pi0370, n7737);
  not g9414 (n_4398, n7738);
  not g9415 (n_4399, n7739);
  and g9416 (n7740, n_4398, n_4399);
  not g9417 (n_4401, pi0371);
  not g9418 (n_4402, n7740);
  and g9419 (n7741, n_4401, n_4402);
  and g9420 (n7742, pi0371, n7740);
  not g9421 (n_4403, n7741);
  not g9422 (n_4404, n7742);
  and g9423 (n7743, n_4403, n_4404);
  not g9424 (n_4406, pi0373);
  not g9425 (n_4407, n7743);
  and g9426 (n7744, n_4406, n_4407);
  and g9427 (n7745, pi0373, n7743);
  not g9428 (n_4408, n7744);
  not g9429 (n_4409, n7745);
  and g9430 (n7746, n_4408, n_4409);
  not g9431 (n_4411, n7746);
  and g9432 (n7747, pi0375, n_4411);
  not g9433 (n_4412, pi0375);
  and g9434 (n7748, n_4412, n7746);
  not g9435 (n_4413, n7747);
  not g9436 (n_4414, n7748);
  and g9437 (n7749, n_4413, n_4414);
  not g9438 (n_4415, n7734);
  not g9439 (n_4416, n7749);
  and g9440 (n7750, n_4415, n_4416);
  and g9441 (n7751, n7734, n7749);
  not g9442 (n_4417, n7750);
  not g9443 (n_4418, n7751);
  and g9444 (n7752, n_4417, n_4418);
  and g9445 (n7753, n7727, n7752);
  not g9446 (n_4419, n7644);
  not g9447 (n_4420, n7728);
  and g9448 (n7754, n_4419, n_4420);
  not g9449 (n_4421, n7753);
  and g9450 (n7755, n_4421, n7754);
  not g9451 (n_4423, pi0590);
  not g9452 (n_4424, n7755);
  and g9453 (n7756, n_4423, n_4424);
  and g9454 (n7757, pi0351, pi1199);
  not g9455 (n_4428, pi0346);
  and g9456 (n7758, pi0345, n_4428);
  not g9457 (n_4429, pi0345);
  and g9458 (n7759, n_4429, pi0346);
  not g9459 (n_4430, n7758);
  not g9460 (n_4431, n7759);
  and g9461 (n7760, n_4430, n_4431);
  not g9462 (n_4433, n7760);
  and g9463 (n7761, pi0323, n_4433);
  not g9464 (n_4434, pi0323);
  and g9465 (n7762, n_4434, n7760);
  not g9466 (n_4435, n7761);
  not g9467 (n_4436, n7762);
  and g9468 (n7763, n_4435, n_4436);
  not g9469 (n_4439, pi0450);
  and g9470 (n7764, pi0358, n_4439);
  not g9471 (n_4440, pi0358);
  and g9472 (n7765, n_4440, pi0450);
  not g9473 (n_4441, n7764);
  not g9474 (n_4442, n7765);
  and g9475 (n7766, n_4441, n_4442);
  not g9476 (n_4443, n7766);
  and g9477 (n7767, n7763, n_4443);
  not g9478 (n_4444, n7763);
  and g9479 (n7768, n_4444, n7766);
  not g9480 (n_4445, n7767);
  not g9481 (n_4446, n7768);
  and g9482 (n7769, n_4445, n_4446);
  not g9483 (n_4449, pi0327);
  not g9484 (n_4450, pi0362);
  and g9485 (n7770, n_4449, n_4450);
  and g9486 (n7771, pi0327, pi0362);
  not g9487 (n_4451, n7770);
  not g9488 (n_4452, n7771);
  and g9489 (n7772, n_4451, n_4452);
  not g9490 (n_4455, pi0344);
  and g9491 (n7773, pi0343, n_4455);
  not g9492 (n_4456, pi0343);
  and g9493 (n7774, n_4456, pi0344);
  not g9494 (n_4457, n7773);
  not g9495 (n_4458, n7774);
  and g9496 (n7775, n_4457, n_4458);
  not g9497 (n_4459, n7775);
  and g9498 (n7776, n7772, n_4459);
  not g9499 (n_4460, n7772);
  and g9500 (n7777, n_4460, n7775);
  not g9501 (n_4461, n7776);
  not g9502 (n_4462, n7777);
  and g9503 (n7778, n_4461, n_4462);
  and g9504 (n7779, n7769, n7778);
  not g9505 (n_4463, n7769);
  not g9506 (n_4464, n7778);
  and g9507 (n7780, n_4463, n_4464);
  not g9508 (n_4465, n7779);
  and g9509 (n7781, pi1197, n_4465);
  not g9510 (n_4466, n7780);
  and g9511 (n7782, n_4466, n7781);
  not g9512 (n_4469, pi0460);
  and g9513 (n7783, pi0320, n_4469);
  not g9514 (n_4470, pi0320);
  and g9515 (n7784, n_4470, pi0460);
  not g9516 (n_4471, n7783);
  not g9517 (n_4472, n7784);
  and g9518 (n7785, n_4471, n_4472);
  not g9519 (n_4474, n7785);
  and g9520 (n7786, pi0342, n_4474);
  not g9521 (n_4475, pi0342);
  and g9522 (n7787, n_4475, n7785);
  not g9523 (n_4476, n7786);
  not g9524 (n_4477, n7787);
  and g9525 (n7788, n_4476, n_4477);
  not g9526 (n_4480, pi0455);
  and g9527 (n7789, pi0452, n_4480);
  not g9528 (n_4481, pi0452);
  and g9529 (n7790, n_4481, pi0455);
  not g9530 (n_4482, n7789);
  not g9531 (n_4483, n7790);
  and g9532 (n7791, n_4482, n_4483);
  and g9533 (n7792, pi0355, n7791);
  not g9534 (n_4485, pi0355);
  not g9535 (n_4486, n7791);
  and g9536 (n7793, n_4485, n_4486);
  not g9537 (n_4487, n7792);
  not g9538 (n_4488, n7793);
  and g9539 (n7794, n_4487, n_4488);
  not g9540 (n_4491, pi0458);
  and g9541 (n7795, pi0361, n_4491);
  not g9542 (n_4492, pi0361);
  and g9543 (n7796, n_4492, pi0458);
  not g9544 (n_4493, n7795);
  not g9545 (n_4494, n7796);
  and g9546 (n7797, n_4493, n_4494);
  and g9547 (n7798, n7794, n7797);
  not g9548 (n_4495, n7794);
  not g9549 (n_4496, n7797);
  and g9550 (n7799, n_4495, n_4496);
  not g9551 (n_4497, n7798);
  not g9552 (n_4498, n7799);
  and g9553 (n7800, n_4497, n_4498);
  not g9554 (n_4500, pi0441);
  and g9555 (n7801, n_4500, n7800);
  not g9556 (n_4501, n7800);
  and g9557 (n7802, pi0441, n_4501);
  not g9558 (n_4502, n7801);
  and g9559 (n7803, n_4239, n_4502);
  not g9560 (n_4503, n7802);
  and g9561 (n7804, n_4503, n7803);
  and g9562 (n7805, n7422, n7788);
  not g9563 (n_4504, n7804);
  and g9564 (n7806, n_4504, n7805);
  and g9565 (n7807, pi0361, n_4500);
  and g9566 (n7808, n_4492, pi0441);
  not g9567 (n_4505, n7807);
  not g9568 (n_4506, n7808);
  and g9569 (n7809, n_4505, n_4506);
  and g9570 (n7810, n7788, n7809);
  not g9571 (n_4507, n7788);
  not g9572 (n_4508, n7809);
  and g9573 (n7811, n_4507, n_4508);
  not g9574 (n_4509, n7810);
  not g9575 (n_4510, n7811);
  and g9576 (n7812, n_4509, n_4510);
  and g9577 (n7813, pi0458, n7812);
  not g9578 (n_4511, n7812);
  and g9579 (n7814, n_4491, n_4511);
  not g9580 (n_4512, n7813);
  not g9581 (n_4513, n7814);
  and g9582 (n7815, n_4512, n_4513);
  and g9583 (n7816, n7794, n7815);
  not g9584 (n_4514, n7815);
  and g9585 (n7817, n_4495, n_4514);
  not g9586 (n_4515, n7816);
  not g9587 (n_4516, n7817);
  and g9588 (n7818, n_4515, n_4516);
  and g9589 (n7819, n_4239, n7818);
  and g9590 (n7820, n7422, n_4507);
  not g9591 (n_4517, n7819);
  and g9592 (n7821, n_4517, n7820);
  not g9593 (n_4518, n7806);
  and g9594 (n7822, pi1196, n_4518);
  not g9595 (n_4519, n7821);
  and g9596 (n7823, n_4519, n7822);
  not g9597 (n_4520, n7823);
  and g9598 (n7824, n_4377, n_4520);
  and g9599 (n7825, pi1196, n7818);
  not g9600 (n_4523, pi0347);
  and g9601 (n7826, pi0321, n_4523);
  not g9602 (n_4524, pi0321);
  and g9603 (n7827, n_4524, pi0347);
  not g9604 (n_4525, n7826);
  not g9605 (n_4526, n7827);
  and g9606 (n7828, n_4525, n_4526);
  not g9607 (n_4529, pi0349);
  and g9608 (n7829, pi0316, n_4529);
  not g9609 (n_4530, pi0316);
  and g9610 (n7830, n_4530, pi0349);
  not g9611 (n_4531, n7829);
  not g9612 (n_4532, n7830);
  and g9613 (n7831, n_4531, n_4532);
  and g9614 (n7832, pi0348, n7831);
  not g9615 (n_4534, pi0348);
  not g9616 (n_4535, n7831);
  and g9617 (n7833, n_4534, n_4535);
  not g9618 (n_4536, n7832);
  not g9619 (n_4537, n7833);
  and g9620 (n7834, n_4536, n_4537);
  not g9621 (n_4540, pi0359);
  and g9622 (n7835, pi0315, n_4540);
  not g9623 (n_4541, pi0315);
  and g9624 (n7836, n_4541, pi0359);
  not g9625 (n_4542, n7835);
  not g9626 (n_4543, n7836);
  and g9627 (n7837, n_4542, n_4543);
  and g9628 (n7838, pi0322, n7837);
  not g9629 (n_4545, pi0322);
  not g9630 (n_4546, n7837);
  and g9631 (n7839, n_4545, n_4546);
  not g9632 (n_4547, n7838);
  not g9633 (n_4548, n7839);
  and g9634 (n7840, n_4547, n_4548);
  not g9635 (n_4549, n7840);
  and g9636 (n7841, n7834, n_4549);
  not g9637 (n_4550, n7834);
  and g9638 (n7842, n_4550, n7840);
  not g9639 (n_4551, n7841);
  not g9640 (n_4552, n7842);
  and g9641 (n7843, n_4551, n_4552);
  and g9642 (n7844, n7828, n7843);
  not g9643 (n_4553, n7828);
  not g9644 (n_4554, n7843);
  and g9645 (n7845, n_4553, n_4554);
  not g9646 (n_4555, n7844);
  not g9647 (n_4556, n7845);
  and g9648 (n7846, n_4555, n_4556);
  not g9649 (n_4558, n7846);
  and g9650 (n7847, pi0350, n_4558);
  not g9651 (n_4559, pi0350);
  and g9652 (n7848, n_4559, n7846);
  not g9653 (n_4560, n7847);
  not g9654 (n_4561, n7848);
  and g9655 (n7849, n_4560, n_4561);
  not g9656 (n_4562, n7825);
  and g9657 (n7850, n_4562, n7849);
  and g9658 (n7851, pi1198, n7644);
  and g9659 (n7852, n7850, n7851);
  not g9660 (n_4563, n7824);
  not g9661 (n_4564, n7852);
  and g9662 (n7853, n_4563, n_4564);
  not g9663 (n_4565, n7782);
  not g9664 (n_4566, n7853);
  and g9665 (n7854, n_4565, n_4566);
  not g9666 (n_4567, n7854);
  and g9667 (n7855, n_4239, n_4567);
  not g9668 (n_4568, n7855);
  and g9669 (n7856, n7422, n_4568);
  not g9670 (n_4569, n7757);
  not g9671 (n_4570, n7856);
  and g9672 (n7857, n_4569, n_4570);
  not g9673 (n_4571, n7645);
  and g9674 (n7858, pi1199, n_4571);
  and g9675 (n7859, pi0351, n7858);
  not g9676 (n_4572, n7857);
  not g9677 (n_4573, n7859);
  and g9678 (n7860, n_4572, n_4573);
  not g9679 (n_4575, pi0461);
  not g9680 (n_4576, n7860);
  and g9681 (n7861, n_4575, n_4576);
  not g9682 (n_4577, pi0351);
  and g9683 (n7862, n_4577, pi1199);
  not g9684 (n_4578, n7862);
  and g9685 (n7863, n_4570, n_4578);
  and g9686 (n7864, n_4577, n7858);
  not g9687 (n_4579, n7863);
  not g9688 (n_4580, n7864);
  and g9689 (n7865, n_4579, n_4580);
  not g9690 (n_4581, n7865);
  and g9691 (n7866, pi0461, n_4581);
  not g9692 (n_4582, n7861);
  not g9693 (n_4583, n7866);
  and g9694 (n7867, n_4582, n_4583);
  not g9695 (n_4585, pi0357);
  not g9696 (n_4586, n7867);
  and g9697 (n7868, n_4585, n_4586);
  and g9698 (n7869, n_4575, n_4581);
  and g9699 (n7870, pi0461, n_4576);
  not g9700 (n_4587, n7869);
  not g9701 (n_4588, n7870);
  and g9702 (n7871, n_4587, n_4588);
  not g9703 (n_4589, n7871);
  and g9704 (n7872, pi0357, n_4589);
  not g9705 (n_4590, n7868);
  not g9706 (n_4591, n7872);
  and g9707 (n7873, n_4590, n_4591);
  not g9708 (n_4593, pi0356);
  not g9709 (n_4594, n7873);
  and g9710 (n7874, n_4593, n_4594);
  and g9711 (n7875, n_4585, n_4589);
  and g9712 (n7876, pi0357, n_4586);
  not g9713 (n_4595, n7875);
  not g9714 (n_4596, n7876);
  and g9715 (n7877, n_4595, n_4596);
  not g9716 (n_4597, n7877);
  and g9717 (n7878, pi0356, n_4597);
  not g9718 (n_4600, pi0462);
  and g9719 (n7879, pi0360, n_4600);
  not g9720 (n_4601, pi0360);
  and g9721 (n7880, n_4601, pi0462);
  not g9722 (n_4602, n7879);
  not g9723 (n_4603, n7880);
  and g9724 (n7881, n_4602, n_4603);
  not g9725 (n_4606, pi0353);
  and g9726 (n7882, pi0352, n_4606);
  not g9727 (n_4607, pi0352);
  and g9728 (n7883, n_4607, pi0353);
  not g9729 (n_4608, n7882);
  not g9730 (n_4609, n7883);
  and g9731 (n7884, n_4608, n_4609);
  and g9732 (n7885, n7881, n7884);
  not g9733 (n_4610, n7881);
  not g9734 (n_4611, n7884);
  and g9735 (n7886, n_4610, n_4611);
  not g9736 (n_4612, n7885);
  not g9737 (n_4613, n7886);
  and g9738 (n7887, n_4612, n_4613);
  not g9739 (n_4615, n7887);
  and g9740 (n7888, pi0354, n_4615);
  not g9741 (n_4616, pi0354);
  and g9742 (n7889, n_4616, n7887);
  not g9743 (n_4617, n7888);
  not g9744 (n_4618, n7889);
  and g9745 (n7890, n_4617, n_4618);
  not g9746 (n_4619, n7874);
  and g9747 (n7891, n_4619, n7890);
  not g9748 (n_4620, n7878);
  and g9749 (n7892, n_4620, n7891);
  and g9750 (n7893, n_4593, n_4597);
  and g9751 (n7894, pi0356, n_4594);
  not g9752 (n_4621, n7890);
  not g9753 (n_4622, n7893);
  and g9754 (n7895, n_4621, n_4622);
  not g9755 (n_4623, n7894);
  and g9756 (n7896, n_4623, n7895);
  not g9757 (n_4624, n7892);
  not g9758 (n_4625, n7896);
  and g9759 (n7897, n_4624, n_4625);
  not g9760 (n_4626, n7897);
  and g9761 (n7898, pi0590, n_4626);
  not g9762 (n_4628, pi0591);
  not g9763 (n_4629, n7756);
  and g9764 (n7899, n_4628, n_4629);
  not g9765 (n_4630, n7898);
  and g9766 (n7900, n_4630, n7899);
  and g9767 (n7901, pi0590, n7422);
  and g9768 (n7902, pi1197, n_4571);
  not g9769 (n_4633, pi0409);
  and g9770 (n7903, pi0318, n_4633);
  not g9771 (n_4634, pi0318);
  and g9772 (n7904, n_4634, pi0409);
  not g9773 (n_4635, n7903);
  not g9774 (n_4636, n7904);
  and g9775 (n7905, n_4635, n_4636);
  not g9776 (n_4639, pi0402);
  and g9777 (n7906, pi0401, n_4639);
  not g9778 (n_4640, pi0401);
  and g9779 (n7907, n_4640, pi0402);
  not g9780 (n_4641, n7906);
  not g9781 (n_4642, n7907);
  and g9782 (n7908, n_4641, n_4642);
  and g9783 (n7909, pi0406, n7908);
  not g9784 (n_4644, pi0406);
  not g9785 (n_4645, n7908);
  and g9786 (n7910, n_4644, n_4645);
  not g9787 (n_4646, n7909);
  not g9788 (n_4647, n7910);
  and g9789 (n7911, n_4646, n_4647);
  not g9790 (n_4650, pi0403);
  not g9791 (n_4651, pi0405);
  and g9792 (n7912, n_4650, n_4651);
  and g9793 (n7913, pi0403, pi0405);
  not g9794 (n_4652, n7912);
  not g9795 (n_4653, n7913);
  and g9796 (n7914, n_4652, n_4653);
  not g9797 (n_4656, pi0326);
  and g9798 (n7915, pi0325, n_4656);
  not g9799 (n_4657, pi0325);
  and g9800 (n7916, n_4657, pi0326);
  not g9801 (n_4658, n7915);
  not g9802 (n_4659, n7916);
  and g9803 (n7917, n_4658, n_4659);
  and g9804 (n7918, n7914, n7917);
  not g9805 (n_4660, n7914);
  not g9806 (n_4661, n7917);
  and g9807 (n7919, n_4660, n_4661);
  not g9808 (n_4662, n7918);
  not g9809 (n_4663, n7919);
  and g9810 (n7920, n_4662, n_4663);
  not g9811 (n_4664, n7920);
  and g9812 (n7921, n7911, n_4664);
  not g9813 (n_4665, n7911);
  and g9814 (n7922, n_4665, n7920);
  not g9815 (n_4666, n7921);
  not g9816 (n_4667, n7922);
  and g9817 (n7923, n_4666, n_4667);
  and g9818 (n7924, n7905, n7923);
  not g9819 (n_4668, n7905);
  not g9820 (n_4669, n7923);
  and g9821 (n7925, n_4668, n_4669);
  not g9822 (n_4670, n7924);
  not g9823 (n_4671, n7925);
  and g9824 (n7926, n_4670, n_4671);
  not g9825 (n_4672, n7926);
  and g9826 (n7927, n7485, n_4672);
  and g9827 (n7928, n_3128, n7927);
  and g9828 (n7929, pi0567, n7928);
  not g9829 (n_4675, pi0410);
  and g9830 (n7930, pi0390, n_4675);
  not g9831 (n_4676, pi0390);
  and g9832 (n7931, n_4676, pi0410);
  not g9833 (n_4677, n7930);
  not g9834 (n_4678, n7931);
  and g9835 (n7932, n_4677, n_4678);
  not g9836 (n_4681, pi0412);
  and g9837 (n7933, pi0397, n_4681);
  not g9838 (n_4682, pi0397);
  and g9839 (n7934, n_4682, pi0412);
  not g9840 (n_4683, n7933);
  not g9841 (n_4684, n7934);
  and g9842 (n7935, n_4683, n_4684);
  and g9843 (n7936, pi0404, n7935);
  not g9844 (n_4686, pi0404);
  not g9845 (n_4687, n7935);
  and g9846 (n7937, n_4686, n_4687);
  not g9847 (n_4688, n7936);
  not g9848 (n_4689, n7937);
  and g9849 (n7938, n_4688, n_4689);
  not g9850 (n_4692, pi0324);
  and g9851 (n7939, pi0319, n_4692);
  not g9852 (n_4693, pi0319);
  and g9853 (n7940, n_4693, pi0324);
  not g9854 (n_4694, n7939);
  not g9855 (n_4695, n7940);
  and g9856 (n7941, n_4694, n_4695);
  not g9857 (n_4697, n7941);
  and g9858 (n7942, pi0456, n_4697);
  not g9859 (n_4698, pi0456);
  and g9860 (n7943, n_4698, n7941);
  not g9861 (n_4699, n7942);
  not g9862 (n_4700, n7943);
  and g9863 (n7944, n_4699, n_4700);
  not g9864 (n_4701, n7944);
  and g9865 (n7945, n7938, n_4701);
  not g9866 (n_4702, n7938);
  and g9867 (n7946, n_4702, n7944);
  not g9868 (n_4703, n7945);
  not g9869 (n_4704, n7946);
  and g9870 (n7947, n_4703, n_4704);
  and g9871 (n7948, n7932, n7947);
  not g9872 (n_4705, n7932);
  not g9873 (n_4706, n7947);
  and g9874 (n7949, n_4705, n_4706);
  not g9875 (n_4707, n7948);
  not g9876 (n_4708, n7949);
  and g9877 (n7950, n_4707, n_4708);
  and g9878 (n7951, pi0411, n7950);
  not g9879 (n_4710, pi0411);
  not g9880 (n_4711, n7950);
  and g9881 (n7952, n_4710, n_4711);
  not g9882 (n_4712, n7951);
  not g9883 (n_4713, n7952);
  and g9884 (n7953, n_4712, n_4713);
  not g9885 (n_4714, n7953);
  and g9886 (n7954, pi1196, n_4714);
  and g9887 (n7955, n_4239, n7929);
  not g9888 (n_4715, n7954);
  and g9889 (n7956, n_4715, n7955);
  not g9890 (n_4716, n7956);
  and g9891 (n7957, n7858, n_4716);
  and g9892 (n7958, n_4239, pi1196);
  not g9893 (n_4717, n7958);
  and g9894 (n7959, n7422, n_4717);
  and g9895 (n7960, n7485, n7953);
  and g9896 (n7961, n_3128, n7960);
  and g9897 (n7962, pi0567, n7961);
  and g9898 (n7963, n7958, n7962);
  not g9899 (n_4718, pi1199);
  not g9900 (n_4719, n7959);
  and g9901 (n7964, n_4718, n_4719);
  not g9902 (n_4720, n7963);
  and g9903 (n7965, n_4720, n7964);
  not g9904 (n_4721, n7957);
  not g9905 (n_4722, n7965);
  and g9906 (n7966, n_4721, n_4722);
  not g9907 (n_4723, pi1197);
  not g9908 (n_4724, n7966);
  and g9909 (n7967, n_4723, n_4724);
  not g9910 (n_4725, n7902);
  not g9911 (n_4726, n7967);
  and g9912 (n7968, n_4725, n_4726);
  not g9913 (n_4728, n7968);
  and g9914 (n7969, pi0333, n_4728);
  and g9915 (n7970, pi1198, n_4571);
  not g9916 (n_4729, n7970);
  and g9917 (n7971, n7966, n_4729);
  not g9918 (n_4732, pi0408);
  and g9919 (n7972, pi0328, n_4732);
  not g9920 (n_4733, pi0328);
  and g9921 (n7973, n_4733, pi0408);
  not g9922 (n_4734, n7972);
  not g9923 (n_4735, n7973);
  and g9924 (n7974, n_4734, n_4735);
  not g9925 (n_4738, pi0394);
  not g9926 (n_4739, pi0396);
  and g9927 (n7975, n_4738, n_4739);
  and g9928 (n7976, pi0394, pi0396);
  not g9929 (n_4740, n7975);
  not g9930 (n_4741, n7976);
  and g9931 (n7977, n_4740, n_4741);
  not g9932 (n_4742, n7977);
  and g9933 (n7978, n7974, n_4742);
  not g9934 (n_4743, n7974);
  and g9935 (n7979, n_4743, n7977);
  not g9936 (n_4744, n7978);
  not g9937 (n_4745, n7979);
  and g9938 (n7980, n_4744, n_4745);
  not g9939 (n_4748, pi0399);
  and g9940 (n7981, pi0398, n_4748);
  not g9941 (n_4749, pi0398);
  and g9942 (n7982, n_4749, pi0399);
  not g9943 (n_4750, n7981);
  not g9944 (n_4751, n7982);
  and g9945 (n7983, n_4750, n_4751);
  and g9946 (n7984, pi0395, n7983);
  not g9947 (n_4753, pi0395);
  not g9948 (n_4754, n7983);
  and g9949 (n7985, n_4753, n_4754);
  not g9950 (n_4755, n7984);
  not g9951 (n_4756, n7985);
  and g9952 (n7986, n_4755, n_4756);
  not g9953 (n_4758, n7986);
  and g9954 (n7987, pi0329, n_4758);
  not g9955 (n_4759, pi0329);
  and g9956 (n7988, n_4759, n7986);
  not g9957 (n_4760, n7987);
  not g9958 (n_4761, n7988);
  and g9959 (n7989, n_4760, n_4761);
  not g9960 (n_4763, n7989);
  and g9961 (n7990, pi0400, n_4763);
  not g9962 (n_4764, pi0400);
  and g9963 (n7991, n_4764, n7989);
  not g9964 (n_4765, n7990);
  not g9965 (n_4766, n7991);
  and g9966 (n7992, n_4765, n_4766);
  and g9967 (n7993, n7980, n7992);
  not g9968 (n_4767, n7980);
  not g9969 (n_4768, n7992);
  and g9970 (n7994, n_4767, n_4768);
  not g9971 (n_4769, n7993);
  not g9972 (n_4770, n7994);
  and g9973 (n7995, n_4769, n_4770);
  not g9974 (n_4771, n7971);
  not g9975 (n_4772, n7995);
  and g9976 (n7996, n_4771, n_4772);
  not g9977 (n_4773, pi0333);
  and g9978 (n7997, n_4773, n_4724);
  not g9979 (n_4774, n7996);
  not g9980 (n_4775, n7997);
  and g9981 (n7998, n_4774, n_4775);
  not g9982 (n_4776, n7969);
  and g9983 (n7999, n_4776, n7998);
  not g9984 (n_4778, pi0391);
  not g9985 (n_4779, n7999);
  and g9986 (n8000, n_4778, n_4779);
  and g9987 (n8001, n_4773, n_4728);
  and g9988 (n8002, n7966, n_4774);
  not g9989 (n_4780, n8001);
  and g9990 (n8003, n_4780, n8002);
  not g9991 (n_4781, n8003);
  and g9992 (n8004, pi0391, n_4781);
  not g9993 (n_4782, n8000);
  not g9994 (n_4783, n8004);
  and g9995 (n8005, n_4782, n_4783);
  not g9996 (n_4785, pi0392);
  not g9997 (n_4786, n8005);
  and g9998 (n8006, n_4785, n_4786);
  and g9999 (n8007, n_4778, n_4781);
  and g10000 (n8008, pi0391, n_4779);
  not g10001 (n_4787, n8007);
  not g10002 (n_4788, n8008);
  and g10003 (n8009, n_4787, n_4788);
  not g10004 (n_4789, n8009);
  and g10005 (n8010, pi0392, n_4789);
  not g10006 (n_4790, n8006);
  not g10007 (n_4791, n8010);
  and g10008 (n8011, n_4790, n_4791);
  not g10009 (n_4793, pi0393);
  not g10010 (n_4794, n8011);
  and g10011 (n8012, n_4793, n_4794);
  and g10012 (n8013, n_4785, n_4789);
  and g10013 (n8014, pi0392, n_4786);
  not g10014 (n_4795, n8013);
  not g10015 (n_4796, n8014);
  and g10016 (n8015, n_4795, n_4796);
  not g10017 (n_4797, n8015);
  and g10018 (n8016, pi0393, n_4797);
  not g10019 (n_4800, pi0463);
  and g10020 (n8017, pi0407, n_4800);
  not g10021 (n_4801, pi0407);
  and g10022 (n8018, n_4801, pi0463);
  not g10023 (n_4802, n8017);
  not g10024 (n_4803, n8018);
  and g10025 (n8019, n_4802, n_4803);
  not g10026 (n_4806, pi0413);
  and g10027 (n8020, pi0335, n_4806);
  not g10028 (n_4807, pi0335);
  and g10029 (n8021, n_4807, pi0413);
  not g10030 (n_4808, n8020);
  not g10031 (n_4809, n8021);
  and g10032 (n8022, n_4808, n_4809);
  and g10033 (n8023, n8019, n8022);
  not g10034 (n_4810, n8019);
  not g10035 (n_4811, n8022);
  and g10036 (n8024, n_4810, n_4811);
  not g10037 (n_4812, n8023);
  not g10038 (n_4813, n8024);
  and g10039 (n8025, n_4812, n_4813);
  not g10040 (n_4815, n8025);
  and g10041 (n8026, pi0334, n_4815);
  not g10042 (n_4816, pi0334);
  and g10043 (n8027, n_4816, n8025);
  not g10044 (n_4817, n8026);
  not g10045 (n_4818, n8027);
  and g10046 (n8028, n_4817, n_4818);
  not g10047 (n_4819, n8012);
  and g10048 (n8029, n_4819, n8028);
  not g10049 (n_4820, n8016);
  and g10050 (n8030, n_4820, n8029);
  and g10051 (n8031, n_4793, n_4797);
  and g10052 (n8032, pi0393, n_4794);
  not g10053 (n_4821, n8028);
  not g10054 (n_4822, n8031);
  and g10055 (n8033, n_4821, n_4822);
  not g10056 (n_4823, n8032);
  and g10057 (n8034, n_4823, n8033);
  not g10058 (n_4824, n8030);
  not g10059 (n_4825, n8034);
  and g10060 (n8035, n_4824, n_4825);
  not g10061 (n_4826, n8035);
  and g10062 (n8036, n_4423, n_4826);
  not g10063 (n_4827, n7901);
  and g10064 (n8037, pi0591, n_4827);
  not g10065 (n_4828, n8036);
  and g10066 (n8038, n_4828, n8037);
  not g10067 (n_4829, n7900);
  not g10068 (n_4830, n8038);
  and g10069 (n8039, n_4829, n_4830);
  not g10070 (n_4832, pi0588);
  not g10071 (n_4833, n8039);
  and g10072 (n8040, n_4832, n_4833);
  and g10073 (n8041, n_4423, n_4628);
  not g10074 (n_4834, n8041);
  and g10075 (n8042, n7422, n_4834);
  not g10076 (n_4837, pi0417);
  not g10077 (n_4838, pi0418);
  and g10078 (n8043, n_4837, n_4838);
  and g10079 (n8044, pi0417, pi0418);
  not g10080 (n_4839, n8043);
  not g10081 (n_4840, n8044);
  and g10082 (n8045, n_4839, n_4840);
  and g10083 (n8046, pi0437, n8045);
  not g10084 (n_4842, pi0437);
  not g10085 (n_4843, n8045);
  and g10086 (n8047, n_4842, n_4843);
  not g10087 (n_4844, n8046);
  not g10088 (n_4845, n8047);
  and g10089 (n8048, n_4844, n_4845);
  not g10090 (n_4848, pi0464);
  and g10091 (n8049, pi0453, n_4848);
  not g10092 (n_4849, pi0453);
  and g10093 (n8050, n_4849, pi0464);
  not g10094 (n_4850, n8049);
  not g10095 (n_4851, n8050);
  and g10096 (n8051, n_4850, n_4851);
  and g10097 (n8052, n8048, n8051);
  not g10098 (n_4852, n8048);
  not g10099 (n_4853, n8051);
  and g10100 (n8053, n_4852, n_4853);
  not g10101 (n_4854, n8052);
  not g10102 (n_4855, n8053);
  and g10103 (n8054, n_4854, n_4855);
  not g10104 (n_4858, pi0431);
  and g10105 (n8055, pi0415, n_4858);
  not g10106 (n_4859, pi0415);
  and g10107 (n8056, n_4859, pi0431);
  not g10108 (n_4860, n8055);
  not g10109 (n_4861, n8056);
  and g10110 (n8057, n_4860, n_4861);
  not g10111 (n_4864, pi0438);
  and g10112 (n8058, pi0416, n_4864);
  not g10113 (n_4865, pi0416);
  and g10114 (n8059, n_4865, pi0438);
  not g10115 (n_4866, n8058);
  not g10116 (n_4867, n8059);
  and g10117 (n8060, n_4866, n_4867);
  and g10118 (n8061, n8057, n8060);
  not g10119 (n_4868, n8057);
  not g10120 (n_4869, n8060);
  and g10121 (n8062, n_4868, n_4869);
  not g10122 (n_4870, n8061);
  not g10123 (n_4871, n8062);
  and g10124 (n8063, n_4870, n_4871);
  not g10125 (n_4872, n8063);
  and g10126 (n8064, n8054, n_4872);
  not g10127 (n_4873, n8054);
  and g10128 (n8065, n_4873, n8063);
  not g10129 (n_4874, n8064);
  and g10130 (n8066, pi1197, n_4874);
  not g10131 (n_4875, n8065);
  and g10132 (n8067, n_4875, n8066);
  not g10133 (n_4878, pi0454);
  and g10134 (n8068, pi0421, n_4878);
  not g10135 (n_4879, pi0421);
  and g10136 (n8069, n_4879, pi0454);
  not g10137 (n_4880, n8068);
  not g10138 (n_4881, n8069);
  and g10139 (n8070, n_4880, n_4881);
  not g10140 (n_4884, pi0459);
  and g10141 (n8071, pi0432, n_4884);
  not g10142 (n_4885, pi0432);
  and g10143 (n8072, n_4885, pi0459);
  not g10144 (n_4886, n8071);
  not g10145 (n_4887, n8072);
  and g10146 (n8073, n_4886, n_4887);
  not g10147 (n_4888, n8073);
  and g10148 (n8074, n8070, n_4888);
  not g10149 (n_4889, n8070);
  and g10150 (n8075, n_4889, n8073);
  not g10151 (n_4890, n8074);
  not g10152 (n_4891, n8075);
  and g10153 (n8076, n_4890, n_4891);
  not g10154 (n_4894, pi0419);
  not g10155 (n_4895, pi0420);
  and g10156 (n8077, n_4894, n_4895);
  and g10157 (n8078, pi0419, pi0420);
  not g10158 (n_4896, n8077);
  not g10159 (n_4897, n8078);
  and g10160 (n8079, n_4896, n_4897);
  not g10161 (n_4900, pi0424);
  and g10162 (n8080, pi0423, n_4900);
  not g10163 (n_4901, pi0423);
  and g10164 (n8081, n_4901, pi0424);
  not g10165 (n_4902, n8080);
  not g10166 (n_4903, n8081);
  and g10167 (n8082, n_4902, n_4903);
  not g10168 (n_4904, n8082);
  and g10169 (n8083, n8079, n_4904);
  not g10170 (n_4905, n8079);
  and g10171 (n8084, n_4905, n8082);
  not g10172 (n_4906, n8083);
  not g10173 (n_4907, n8084);
  and g10174 (n8085, n_4906, n_4907);
  and g10175 (n8086, n8076, n8085);
  not g10176 (n_4908, n8076);
  not g10177 (n_4909, n8085);
  and g10178 (n8087, n_4908, n_4909);
  not g10179 (n_4910, n8086);
  not g10180 (n_4911, n8087);
  and g10181 (n8088, n_4910, n_4911);
  not g10182 (n_4913, n8088);
  and g10183 (n8089, pi0425, n_4913);
  not g10184 (n_4914, pi0425);
  and g10185 (n8090, n_4914, n8088);
  not g10186 (n_4915, n8089);
  and g10187 (n8091, pi1198, n_4915);
  not g10188 (n_4916, n8090);
  and g10189 (n8092, n_4916, n8091);
  not g10190 (n_4917, n8067);
  not g10191 (n_4918, n8092);
  and g10192 (n8093, n_4917, n_4918);
  not g10193 (n_4921, pi0429);
  not g10194 (n_4922, pi0435);
  and g10195 (n8094, n_4921, n_4922);
  and g10196 (n8095, pi0429, pi0435);
  not g10197 (n_4923, n8094);
  not g10198 (n_4924, n8095);
  and g10199 (n8096, n_4923, n_4924);
  not g10200 (n_4927, pi0446);
  and g10201 (n8097, pi0434, n_4927);
  not g10202 (n_4928, pi0434);
  and g10203 (n8098, n_4928, pi0446);
  not g10204 (n_4929, n8097);
  not g10205 (n_4930, n8098);
  and g10206 (n8099, n_4929, n_4930);
  not g10207 (n_4933, pi0422);
  and g10208 (n8100, pi0414, n_4933);
  not g10209 (n_4934, pi0414);
  and g10210 (n8101, n_4934, pi0422);
  not g10211 (n_4935, n8100);
  not g10212 (n_4936, n8101);
  and g10213 (n8102, n_4935, n_4936);
  and g10214 (n8103, n8099, n8102);
  not g10215 (n_4937, n8099);
  not g10216 (n_4938, n8102);
  and g10217 (n8104, n_4937, n_4938);
  not g10218 (n_4939, n8103);
  not g10219 (n_4940, n8104);
  and g10220 (n8105, n_4939, n_4940);
  and g10221 (n8106, n8096, n8105);
  not g10222 (n_4941, n8096);
  not g10223 (n_4942, n8105);
  and g10224 (n8107, n_4941, n_4942);
  not g10225 (n_4943, n8106);
  not g10226 (n_4944, n8107);
  and g10227 (n8108, n_4943, n_4944);
  not g10228 (n_4947, pi0443);
  and g10229 (n8109, pi0436, n_4947);
  not g10230 (n_4948, pi0436);
  and g10231 (n8110, n_4948, pi0443);
  not g10232 (n_4949, n8109);
  not g10233 (n_4950, n8110);
  and g10234 (n8111, n_4949, n_4950);
  not g10235 (n_4952, pi0444);
  and g10236 (n8112, n_4952, n8111);
  not g10237 (n_4953, n8111);
  and g10238 (n8113, pi0444, n_4953);
  not g10239 (n_4954, n8112);
  not g10240 (n_4955, n8113);
  and g10241 (n8114, n_4954, n_4955);
  not g10242 (n_4956, n8108);
  not g10243 (n_4957, n8114);
  and g10244 (n8115, n_4956, n_4957);
  and g10245 (n8116, n8108, n8114);
  not g10246 (n_4958, n8115);
  and g10247 (n8117, n7958, n_4958);
  not g10248 (n_4959, n8116);
  and g10249 (n8118, n_4959, n8117);
  not g10250 (n_4960, n8118);
  and g10251 (n8119, n8093, n_4960);
  and g10252 (n8120, n7644, n8119);
  and g10253 (n8121, n_4718, n_4571);
  not g10254 (n_4961, n8120);
  and g10255 (n8122, n_4961, n8121);
  not g10256 (n_4964, pi0451);
  and g10257 (n8123, pi0433, n_4964);
  not g10258 (n_4965, pi0433);
  and g10259 (n8124, n_4965, pi0451);
  not g10260 (n_4966, n8123);
  not g10261 (n_4967, n8124);
  and g10262 (n8125, n_4966, n_4967);
  and g10263 (n8126, pi0449, n8125);
  not g10264 (n_4969, pi0449);
  not g10265 (n_4970, n8125);
  and g10266 (n8127, n_4969, n_4970);
  not g10267 (n_4971, n8126);
  not g10268 (n_4972, n8127);
  and g10269 (n8128, n_4971, n_4972);
  not g10270 (n_4974, pi0427);
  and g10271 (n8129, n_4974, pi0428);
  not g10272 (n_4976, pi0428);
  and g10273 (n8130, pi0427, n_4976);
  not g10274 (n_4977, n8129);
  not g10275 (n_4978, n8130);
  and g10276 (n8131, n_4977, n_4978);
  not g10277 (n_4980, n8131);
  and g10278 (n8132, pi0430, n_4980);
  not g10279 (n_4981, pi0430);
  and g10280 (n8133, n_4981, n8131);
  not g10281 (n_4982, n8132);
  not g10282 (n_4983, n8133);
  and g10283 (n8134, n_4982, n_4983);
  not g10284 (n_4985, pi0426);
  not g10285 (n_4986, n8134);
  and g10286 (n8135, n_4985, n_4986);
  and g10287 (n8136, pi0426, n8134);
  not g10288 (n_4987, n8135);
  not g10289 (n_4988, n8136);
  and g10290 (n8137, n_4987, n_4988);
  not g10291 (n_4990, pi0445);
  not g10292 (n_4991, n8137);
  and g10293 (n8138, n_4990, n_4991);
  and g10294 (n8139, pi0445, n8137);
  not g10295 (n_4992, n8138);
  not g10296 (n_4993, n8139);
  and g10297 (n8140, n_4992, n_4993);
  not g10298 (n_4995, pi0448);
  not g10299 (n_4996, n8140);
  and g10300 (n8141, n_4995, n_4996);
  and g10301 (n8142, pi0448, n8140);
  not g10302 (n_4997, n8141);
  not g10303 (n_4998, n8142);
  and g10304 (n8143, n_4997, n_4998);
  not g10305 (n_4999, n8143);
  and g10306 (n8144, n8120, n_4999);
  not g10307 (n_5000, n8144);
  and g10308 (n8145, n_4571, n_5000);
  not g10309 (n_5001, n8145);
  and g10310 (n8146, n8128, n_5001);
  and g10311 (n8147, n8120, n8143);
  not g10312 (n_5002, n8147);
  and g10313 (n8148, n_4571, n_5002);
  not g10314 (n_5003, n8128);
  not g10315 (n_5004, n8148);
  and g10316 (n8149, n_5003, n_5004);
  not g10317 (n_5005, n8146);
  and g10318 (n8150, pi1199, n_5005);
  not g10319 (n_5006, n8149);
  and g10320 (n8151, n_5006, n8150);
  not g10321 (n_5007, n8122);
  and g10322 (n8152, n8041, n_5007);
  not g10323 (n_5008, n8151);
  and g10324 (n8153, n_5008, n8152);
  not g10325 (n_5009, n8042);
  and g10326 (n8154, pi0588, n_5009);
  not g10327 (n_5010, n8153);
  and g10328 (n8155, n_5010, n8154);
  not g10329 (n_5011, n8155);
  and g10330 (n8156, n7427, n_5011);
  not g10331 (n_5012, n8040);
  and g10332 (n8157, n_5012, n8156);
  and g10333 (n8158, n7636, n_4834);
  and g10334 (n8159, n_172, n_4211);
  not g10335 (n_5013, n7614);
  and g10336 (n8160, n_5013, n8159);
  and g10337 (n8161, pi0087, n_164);
  and g10338 (n8162, n2530, n8161);
  and g10339 (n8163, n_4132, n8162);
  not g10340 (n_5014, n7494);
  and g10341 (n8164, n_5014, n8163);
  not g10342 (n_5015, n8164);
  and g10343 (n8165, n_171, n_5015);
  not g10344 (n_5016, n8160);
  and g10345 (n8166, n_5016, n8165);
  not g10346 (n_5017, n8166);
  and g10347 (n8167, n_4221, n_5017);
  not g10348 (n_5018, n8167);
  and g10349 (n8168, pi0567, n_5018);
  not g10350 (n_5019, n8168);
  and g10351 (n8169, n7469, n_5019);
  not g10352 (n_5020, n8169);
  and g10353 (n8170, n_4239, n_5020);
  and g10354 (n8171, pi0592, n_4225);
  not g10355 (n_5021, n8170);
  not g10356 (n_5022, n8171);
  and g10357 (n8172, n_5021, n_5022);
  not g10358 (n_5023, n8093);
  and g10359 (n8173, n_5023, n8172);
  not g10360 (n_5024, pi1196);
  and g10361 (n8174, n_5024, n_4225);
  and g10362 (n8175, n_4947, n_4239);
  not g10363 (n_5025, n8175);
  and g10364 (n8176, n_4225, n_5025);
  and g10365 (n8177, n_5020, n8175);
  not g10366 (n_5026, n8176);
  not g10367 (n_5027, n8177);
  and g10368 (n8178, n_5026, n_5027);
  not g10369 (n_5028, n8178);
  and g10370 (n8179, n_4952, n_5028);
  and g10371 (n8180, pi0443, n_4239);
  not g10372 (n_5029, n8180);
  and g10373 (n8181, n_4225, n_5029);
  and g10374 (n8182, n_5020, n8180);
  not g10375 (n_5030, n8181);
  not g10376 (n_5031, n8182);
  and g10377 (n8183, n_5030, n_5031);
  not g10378 (n_5032, n8183);
  and g10379 (n8184, pi0444, n_5032);
  not g10380 (n_5033, n8179);
  not g10381 (n_5034, n8184);
  and g10382 (n8185, n_5033, n_5034);
  not g10383 (n_5035, n8185);
  and g10384 (n8186, n_4948, n_5035);
  and g10385 (n8187, n_4952, n_5032);
  and g10386 (n8188, pi0444, n_5028);
  not g10387 (n_5036, n8187);
  not g10388 (n_5037, n8188);
  and g10389 (n8189, n_5036, n_5037);
  not g10390 (n_5038, n8189);
  and g10391 (n8190, pi0436, n_5038);
  not g10392 (n_5039, n8186);
  and g10393 (n8191, n8108, n_5039);
  not g10394 (n_5040, n8190);
  and g10395 (n8192, n_5040, n8191);
  and g10396 (n8193, n_4948, n_5038);
  and g10397 (n8194, pi0436, n_5035);
  not g10398 (n_5041, n8193);
  and g10399 (n8195, n_4956, n_5041);
  not g10400 (n_5042, n8194);
  and g10401 (n8196, n_5042, n8195);
  not g10402 (n_5043, n8192);
  and g10403 (n8197, pi1196, n_5043);
  not g10404 (n_5044, n8196);
  and g10405 (n8198, n_5044, n8197);
  not g10406 (n_5045, n8174);
  and g10407 (n8199, n8093, n_5045);
  not g10408 (n_5046, n8198);
  and g10409 (n8200, n_5046, n8199);
  not g10410 (n_5047, n8173);
  not g10411 (n_5048, n8200);
  and g10412 (n8201, n_5047, n_5048);
  and g10413 (n8202, n_4718, n8201);
  not g10414 (n_5049, n8201);
  and g10415 (n8203, pi0428, n_5049);
  and g10416 (n8204, n_4976, n8172);
  not g10417 (n_5050, n8203);
  not g10418 (n_5051, n8204);
  and g10419 (n8205, n_5050, n_5051);
  not g10420 (n_5052, n8205);
  and g10421 (n8206, n_4974, n_5052);
  and g10422 (n8207, n_4976, n_5049);
  and g10423 (n8208, pi0428, n8172);
  not g10424 (n_5053, n8207);
  not g10425 (n_5054, n8208);
  and g10426 (n8209, n_5053, n_5054);
  not g10427 (n_5055, n8209);
  and g10428 (n8210, pi0427, n_5055);
  not g10429 (n_5056, n8206);
  not g10430 (n_5057, n8210);
  and g10431 (n8211, n_5056, n_5057);
  not g10432 (n_5058, n8211);
  and g10433 (n8212, pi0430, n_5058);
  and g10434 (n8213, n_4974, n_5055);
  and g10435 (n8214, pi0427, n_5052);
  not g10436 (n_5059, n8213);
  not g10437 (n_5060, n8214);
  and g10438 (n8215, n_5059, n_5060);
  not g10439 (n_5061, n8215);
  and g10440 (n8216, n_4981, n_5061);
  not g10441 (n_5062, n8212);
  not g10442 (n_5063, n8216);
  and g10443 (n8217, n_5062, n_5063);
  not g10444 (n_5064, n8217);
  and g10445 (n8218, pi0426, n_5064);
  and g10446 (n8219, pi0430, n_5061);
  and g10447 (n8220, n_4981, n_5058);
  not g10448 (n_5065, n8219);
  not g10449 (n_5066, n8220);
  and g10450 (n8221, n_5065, n_5066);
  not g10451 (n_5067, n8221);
  and g10452 (n8222, n_4985, n_5067);
  not g10453 (n_5068, n8218);
  not g10454 (n_5069, n8222);
  and g10455 (n8223, n_5068, n_5069);
  not g10456 (n_5070, n8223);
  and g10457 (n8224, pi0445, n_5070);
  and g10458 (n8225, pi0426, n_5067);
  and g10459 (n8226, n_4985, n_5064);
  not g10460 (n_5071, n8225);
  not g10461 (n_5072, n8226);
  and g10462 (n8227, n_5071, n_5072);
  not g10463 (n_5073, n8227);
  and g10464 (n8228, n_4990, n_5073);
  not g10465 (n_5074, n8224);
  not g10466 (n_5075, n8228);
  and g10467 (n8229, n_5074, n_5075);
  and g10468 (n8230, pi0448, n_5003);
  and g10469 (n8231, n_4995, n8128);
  not g10470 (n_5076, n8230);
  not g10471 (n_5077, n8231);
  and g10472 (n8232, n_5076, n_5077);
  not g10473 (n_5078, n8229);
  not g10474 (n_5079, n8232);
  and g10475 (n8233, n_5078, n_5079);
  and g10476 (n8234, pi0445, n_5073);
  and g10477 (n8235, n_4990, n_5070);
  not g10478 (n_5080, n8234);
  not g10479 (n_5081, n8235);
  and g10480 (n8236, n_5080, n_5081);
  not g10481 (n_5082, n8236);
  and g10482 (n8237, n8232, n_5082);
  not g10483 (n_5083, n8233);
  and g10484 (n8238, pi1199, n_5083);
  not g10485 (n_5084, n8237);
  and g10486 (n8239, n_5084, n8238);
  not g10487 (n_5085, n8202);
  and g10488 (n8240, n8041, n_5085);
  not g10489 (n_5086, n8239);
  and g10490 (n8241, n_5086, n8240);
  not g10491 (n_5087, n8158);
  and g10492 (n8242, n7425, n_5087);
  not g10493 (n_5088, n8241);
  and g10494 (n8243, n_5088, n8242);
  not g10495 (n_5089, n7592);
  and g10496 (n8244, n_5089, n_4834);
  and g10497 (n8245, n_5024, n7592);
  and g10498 (n8246, n7592, n_5025);
  and g10499 (n8247, n_4948, pi0444);
  and g10500 (n8248, pi0436, n_4952);
  not g10501 (n_5090, n8247);
  not g10502 (n_5091, n8248);
  and g10503 (n8249, n_5090, n_5091);
  not g10504 (n_5092, n8249);
  and g10505 (n8250, n8108, n_5092);
  and g10506 (n8251, n_4956, n8249);
  not g10507 (n_5093, n8250);
  not g10508 (n_5094, n8251);
  and g10509 (n8252, n_5093, n_5094);
  and g10510 (n8253, n_5027, n8252);
  not g10511 (n_5095, n8246);
  and g10512 (n8254, n_5095, n8253);
  and g10513 (n8255, n7592, n_5029);
  not g10514 (n_5096, n8252);
  and g10515 (n8256, n_5031, n_5096);
  not g10516 (n_5097, n8255);
  and g10517 (n8257, n_5097, n8256);
  not g10518 (n_5098, n8254);
  and g10519 (n8258, pi1196, n_5098);
  not g10520 (n_5099, n8257);
  and g10521 (n8259, n_5099, n8258);
  not g10522 (n_5100, n8245);
  not g10523 (n_5101, n8259);
  and g10524 (n8260, n_5100, n_5101);
  not g10525 (n_5102, n8260);
  and g10526 (n8261, n8093, n_5102);
  and g10527 (n8262, pi0592, n7592);
  not g10528 (n_5103, n8262);
  and g10529 (n8263, n_5021, n_5103);
  not g10530 (n_5104, n8263);
  and g10531 (n8264, n_5023, n_5104);
  not g10532 (n_5105, n8261);
  not g10533 (n_5106, n8264);
  and g10534 (n8265, n_5105, n_5106);
  not g10535 (n_5107, n8265);
  and g10536 (n8266, n_4718, n_5107);
  and g10537 (n8267, n_4976, n8263);
  and g10538 (n8268, pi0428, n8265);
  not g10539 (n_5108, n8267);
  and g10540 (n8269, pi0427, n_5108);
  not g10541 (n_5109, n8268);
  and g10542 (n8270, n_5109, n8269);
  and g10543 (n8271, n_4976, n8265);
  and g10544 (n8272, pi0428, n8263);
  not g10545 (n_5110, n8272);
  and g10546 (n8273, n_4974, n_5110);
  not g10547 (n_5111, n8271);
  and g10548 (n8274, n_5111, n8273);
  not g10549 (n_5112, n8270);
  not g10550 (n_5113, n8274);
  and g10551 (n8275, n_5112, n_5113);
  not g10552 (n_5114, n8275);
  and g10553 (n8276, n_4981, n_5114);
  and g10554 (n8277, n8131, n8263);
  and g10555 (n8278, n_4980, n8265);
  not g10556 (n_5115, n8277);
  not g10557 (n_5116, n8278);
  and g10558 (n8279, n_5115, n_5116);
  and g10559 (n8280, pi0430, n8279);
  not g10560 (n_5117, n8276);
  not g10561 (n_5118, n8280);
  and g10562 (n8281, n_5117, n_5118);
  not g10563 (n_5119, n8281);
  and g10564 (n8282, n_4985, n_5119);
  and g10565 (n8283, pi0430, n_5114);
  and g10566 (n8284, n_4981, n8279);
  not g10567 (n_5120, n8283);
  not g10568 (n_5121, n8284);
  and g10569 (n8285, n_5120, n_5121);
  not g10570 (n_5122, n8285);
  and g10571 (n8286, pi0426, n_5122);
  not g10572 (n_5123, n8282);
  not g10573 (n_5124, n8286);
  and g10574 (n8287, n_5123, n_5124);
  not g10575 (n_5125, n8287);
  and g10576 (n8288, n_4990, n_5125);
  and g10577 (n8289, n_4985, n_5122);
  and g10578 (n8290, pi0426, n_5119);
  not g10579 (n_5126, n8289);
  not g10580 (n_5127, n8290);
  and g10581 (n8291, n_5126, n_5127);
  not g10582 (n_5128, n8291);
  and g10583 (n8292, pi0445, n_5128);
  not g10584 (n_5129, n8288);
  not g10585 (n_5130, n8292);
  and g10586 (n8293, n_5129, n_5130);
  and g10587 (n8294, pi0448, n8293);
  and g10588 (n8295, n_4990, n_5128);
  and g10589 (n8296, pi0445, n_5125);
  not g10590 (n_5131, n8295);
  not g10591 (n_5132, n8296);
  and g10592 (n8297, n_5131, n_5132);
  and g10593 (n8298, n_4995, n8297);
  not g10594 (n_5133, n8294);
  and g10595 (n8299, n_5003, n_5133);
  not g10596 (n_5134, n8298);
  and g10597 (n8300, n_5134, n8299);
  and g10598 (n8301, n_4995, n8293);
  and g10599 (n8302, pi0448, n8297);
  not g10600 (n_5135, n8301);
  and g10601 (n8303, n8128, n_5135);
  not g10602 (n_5136, n8302);
  and g10603 (n8304, n_5136, n8303);
  not g10604 (n_5137, n8300);
  not g10605 (n_5138, n8304);
  and g10606 (n8305, n_5137, n_5138);
  not g10607 (n_5139, n8305);
  and g10608 (n8306, pi1199, n_5139);
  not g10609 (n_5140, n8266);
  and g10610 (n8307, n8041, n_5140);
  not g10611 (n_5141, n8306);
  and g10612 (n8308, n_5141, n8307);
  not g10613 (n_5142, n8244);
  and g10614 (n8309, n_4091, n_5142);
  not g10615 (n_5143, n8308);
  and g10616 (n8310, n_5143, n8309);
  not g10617 (n_5144, n8243);
  not g10618 (n_5145, n8310);
  and g10619 (n8311, n_5144, n_5145);
  not g10620 (n_5146, n8311);
  and g10621 (n8312, pi0588, n_5146);
  and g10622 (n8313, pi0591, n7636);
  not g10623 (n_5147, n8172);
  and g10624 (n8314, n7825, n_5147);
  and g10625 (n8315, n_4559, n_4239);
  not g10626 (n_5148, n8315);
  and g10627 (n8316, n_4225, n_5148);
  and g10628 (n8317, n_5020, n8315);
  not g10629 (n_5149, n8317);
  and g10630 (n8318, n7846, n_5149);
  not g10631 (n_5150, n8316);
  and g10632 (n8319, n_5150, n8318);
  and g10633 (n8320, pi0350, n_4239);
  not g10634 (n_5151, n8320);
  and g10635 (n8321, n_4225, n_5151);
  and g10636 (n8322, n_5020, n8320);
  not g10637 (n_5152, n8322);
  and g10638 (n8323, n_4558, n_5152);
  not g10639 (n_5153, n8321);
  and g10640 (n8324, n_5153, n8323);
  not g10641 (n_5154, n8319);
  and g10642 (n8325, n_4562, n_5154);
  not g10643 (n_5155, n8324);
  and g10644 (n8326, n_5155, n8325);
  not g10645 (n_5156, n8314);
  and g10646 (n8327, pi1198, n_5156);
  not g10647 (n_5157, n8326);
  and g10648 (n8328, n_5157, n8327);
  and g10649 (n8329, n_4480, n_5147);
  and g10650 (n8330, pi0455, n_4225);
  not g10651 (n_5158, n8329);
  not g10652 (n_5159, n8330);
  and g10653 (n8331, n_5158, n_5159);
  not g10654 (n_5160, n8331);
  and g10655 (n8332, n_4481, n_5160);
  and g10656 (n8333, pi0455, n_5147);
  and g10657 (n8334, n_4480, n_4225);
  not g10658 (n_5161, n8333);
  not g10659 (n_5162, n8334);
  and g10660 (n8335, n_5161, n_5162);
  not g10661 (n_5163, n8335);
  and g10662 (n8336, pi0452, n_5163);
  not g10663 (n_5164, n8332);
  not g10664 (n_5165, n8336);
  and g10665 (n8337, n_5164, n_5165);
  not g10666 (n_5166, n8337);
  and g10667 (n8338, n_4485, n_5166);
  and g10668 (n8339, n_4481, n_5163);
  and g10669 (n8340, pi0452, n_5160);
  not g10670 (n_5167, n8339);
  not g10671 (n_5168, n8340);
  and g10672 (n8341, n_5167, n_5168);
  not g10673 (n_5169, n8341);
  and g10674 (n8342, pi0355, n_5169);
  not g10675 (n_5170, n8338);
  not g10676 (n_5171, n8342);
  and g10677 (n8343, n_5170, n_5171);
  not g10678 (n_5172, n8343);
  and g10679 (n8344, pi0458, n_5172);
  and g10680 (n8345, n_4485, n_5169);
  and g10681 (n8346, pi0355, n_5166);
  not g10682 (n_5173, n8345);
  not g10683 (n_5174, n8346);
  and g10684 (n8347, n_5173, n_5174);
  not g10685 (n_5175, n8347);
  and g10686 (n8348, n_4491, n_5175);
  not g10687 (n_5176, n8344);
  and g10688 (n8349, n7812, n_5176);
  not g10689 (n_5177, n8348);
  and g10690 (n8350, n_5177, n8349);
  and g10691 (n8351, pi0458, n_5175);
  and g10692 (n8352, n_4491, n_5172);
  not g10693 (n_5178, n8351);
  and g10694 (n8353, n_4511, n_5178);
  not g10695 (n_5179, n8352);
  and g10696 (n8354, n_5179, n8353);
  not g10697 (n_5180, n8350);
  and g10698 (n8355, pi1196, n_5180);
  not g10699 (n_5181, n8354);
  and g10700 (n8356, n_5181, n8355);
  and g10701 (n8357, n_4377, n_5045);
  not g10702 (n_5182, n8356);
  and g10703 (n8358, n_5182, n8357);
  not g10704 (n_5183, n8328);
  not g10705 (n_5184, n8358);
  and g10706 (n8359, n_5183, n_5184);
  not g10707 (n_5185, n8359);
  and g10708 (n8360, n_4565, n_5185);
  and g10709 (n8361, n7782, n8172);
  not g10710 (n_5186, n8360);
  not g10711 (n_5187, n8361);
  and g10712 (n8362, n_5186, n_5187);
  and g10713 (n8363, n_4578, n8362);
  and g10714 (n8364, pi1199, n_5147);
  and g10715 (n8365, n_4577, n8364);
  not g10716 (n_5188, n8363);
  not g10717 (n_5189, n8365);
  and g10718 (n8366, n_5188, n_5189);
  not g10719 (n_5190, n8366);
  and g10720 (n8367, n_4575, n_5190);
  and g10721 (n8368, n_4569, n8362);
  and g10722 (n8369, pi0351, n8364);
  not g10723 (n_5191, n8368);
  not g10724 (n_5192, n8369);
  and g10725 (n8370, n_5191, n_5192);
  not g10726 (n_5193, n8370);
  and g10727 (n8371, pi0461, n_5193);
  not g10728 (n_5194, n8367);
  not g10729 (n_5195, n8371);
  and g10730 (n8372, n_5194, n_5195);
  not g10731 (n_5196, n8372);
  and g10732 (n8373, n_4585, n_5196);
  and g10733 (n8374, n_4575, n_5193);
  and g10734 (n8375, pi0461, n_5190);
  not g10735 (n_5197, n8374);
  not g10736 (n_5198, n8375);
  and g10737 (n8376, n_5197, n_5198);
  not g10738 (n_5199, n8376);
  and g10739 (n8377, pi0357, n_5199);
  not g10740 (n_5200, n8373);
  not g10741 (n_5201, n8377);
  and g10742 (n8378, n_5200, n_5201);
  not g10743 (n_5202, n8378);
  and g10744 (n8379, n_4593, n_5202);
  and g10745 (n8380, n_4585, n_5199);
  and g10746 (n8381, pi0357, n_5196);
  not g10747 (n_5203, n8380);
  not g10748 (n_5204, n8381);
  and g10749 (n8382, n_5203, n_5204);
  not g10750 (n_5205, n8382);
  and g10751 (n8383, pi0356, n_5205);
  not g10752 (n_5206, n8379);
  not g10753 (n_5207, n8383);
  and g10754 (n8384, n_5206, n_5207);
  not g10755 (n_5208, n8384);
  and g10756 (n8385, n_4621, n_5208);
  and g10757 (n8386, n_4593, n_5205);
  and g10758 (n8387, pi0356, n_5202);
  not g10759 (n_5209, n8386);
  not g10760 (n_5210, n8387);
  and g10761 (n8388, n_5209, n_5210);
  not g10762 (n_5211, n8388);
  and g10763 (n8389, n7890, n_5211);
  not g10764 (n_5212, n8385);
  and g10765 (n8390, n_4628, n_5212);
  not g10766 (n_5213, n8389);
  and g10767 (n8391, n_5213, n8390);
  not g10768 (n_5214, n8313);
  and g10769 (n8392, pi0590, n_5214);
  not g10770 (n_5215, n8391);
  and g10771 (n8393, n_5215, n8392);
  and g10772 (n8394, pi1197, n_5147);
  and g10773 (n8395, pi1198, n_4772);
  and g10774 (n8396, n8172, n8395);
  and g10775 (n8397, n_171, n7954);
  not g10776 (n_5216, n8397);
  and g10777 (n8398, n_4672, n_5216);
  and g10778 (n8399, n7617, n8398);
  not g10779 (n_5217, n8399);
  and g10780 (n8400, n7614, n_5217);
  not g10781 (n_5218, n8400);
  and g10782 (n8401, n8159, n_5218);
  and g10783 (n8402, n_4215, n8162);
  and g10784 (n8403, n7495, n_4672);
  not g10785 (n_5219, n8403);
  and g10786 (n8404, n7626, n_5219);
  not g10787 (n_5220, n8404);
  and g10788 (n8405, n8402, n_5220);
  and g10789 (n8406, n_5024, n8405);
  and g10790 (n8407, n7495, n7953);
  not g10791 (n_5221, n8407);
  and g10792 (n8408, n7626, n_5221);
  not g10793 (n_5222, n8408);
  and g10794 (n8409, n8405, n_5222);
  and g10795 (n8410, n_171, n_4239);
  not g10803 (n_5226, n8410);
  and g10804 (n8415, n_4223, n_5226);
  and g10805 (n8416, n8402, n_5222);
  and g10806 (n8417, n7617, n7953);
  not g10807 (n_5227, n8417);
  and g10808 (n8418, n7614, n_5227);
  not g10809 (n_5228, n8418);
  and g10810 (n8419, n8159, n_5228);
  and g10816 (n8423, n_5024, n7633);
  not g10817 (n_5231, n8422);
  not g10818 (n_5232, n8423);
  and g10819 (n8424, n_5231, n_5232);
  not g10820 (n_5233, n8424);
  and g10821 (n8425, n_4718, n_5233);
  not g10822 (n_5234, n8414);
  not g10823 (n_5235, n8415);
  and g10824 (n8426, n_5234, n_5235);
  not g10825 (n_5236, n8425);
  and g10826 (n8427, n_5236, n8426);
  not g10827 (n_5237, n8427);
  and g10828 (n8428, pi0567, n_5237);
  not g10829 (n_5238, n8395);
  and g10830 (n8429, n7469, n_5238);
  not g10831 (n_5239, n8428);
  and g10832 (n8430, n_5239, n8429);
  not g10833 (n_5240, n8396);
  not g10834 (n_5241, n8430);
  and g10835 (n8431, n_5240, n_5241);
  and g10836 (n8432, n_4723, n8431);
  not g10837 (n_5242, n8394);
  not g10838 (n_5243, n8432);
  and g10839 (n8433, n_5242, n_5243);
  not g10840 (n_5244, n8433);
  and g10841 (n8434, pi0333, n_5244);
  and g10842 (n8435, n_4773, n8431);
  not g10843 (n_5245, n8434);
  not g10844 (n_5246, n8435);
  and g10845 (n8436, n_5245, n_5246);
  not g10846 (n_5247, n8436);
  and g10847 (n8437, pi0391, n_5247);
  not g10848 (n_5248, n8431);
  and g10849 (n8438, pi0333, n_5248);
  and g10850 (n8439, n_4773, n8433);
  not g10851 (n_5249, n8438);
  not g10852 (n_5250, n8439);
  and g10853 (n8440, n_5249, n_5250);
  and g10854 (n8441, n_4778, n8440);
  not g10855 (n_5251, n8437);
  not g10856 (n_5252, n8441);
  and g10857 (n8442, n_5251, n_5252);
  not g10858 (n_5253, n8442);
  and g10859 (n8443, n_4785, n_5253);
  and g10860 (n8444, n_4778, n_5247);
  and g10861 (n8445, pi0391, n8440);
  not g10862 (n_5254, n8444);
  not g10863 (n_5255, n8445);
  and g10864 (n8446, n_5254, n_5255);
  not g10865 (n_5256, n8446);
  and g10866 (n8447, pi0392, n_5256);
  not g10867 (n_5257, n8443);
  not g10868 (n_5258, n8447);
  and g10869 (n8448, n_5257, n_5258);
  not g10870 (n_5259, n8448);
  and g10871 (n8449, n_4793, n_5259);
  and g10872 (n8450, n_4785, n_5256);
  and g10873 (n8451, pi0392, n_5253);
  not g10874 (n_5260, n8450);
  not g10875 (n_5261, n8451);
  and g10876 (n8452, n_5260, n_5261);
  not g10877 (n_5262, n8452);
  and g10878 (n8453, pi0393, n_5262);
  not g10879 (n_5263, n8449);
  not g10880 (n_5264, n8453);
  and g10881 (n8454, n_5263, n_5264);
  and g10882 (n8455, n_4816, n8454);
  and g10883 (n8456, n_4793, n_5262);
  and g10884 (n8457, pi0393, n_5259);
  not g10885 (n_5265, n8456);
  not g10886 (n_5266, n8457);
  and g10887 (n8458, n_5265, n_5266);
  and g10888 (n8459, pi0334, n8458);
  not g10889 (n_5267, n8455);
  and g10890 (n8460, n8025, n_5267);
  not g10891 (n_5268, n8459);
  and g10892 (n8461, n_5268, n8460);
  and g10893 (n8462, n_4816, n8458);
  and g10894 (n8463, pi0334, n8454);
  not g10895 (n_5269, n8462);
  and g10896 (n8464, n_4815, n_5269);
  not g10897 (n_5270, n8463);
  and g10898 (n8465, n_5270, n8464);
  not g10899 (n_5271, n8461);
  and g10900 (n8466, pi0591, n_5271);
  not g10901 (n_5272, n8465);
  and g10902 (n8467, n_5272, n8466);
  and g10903 (n8468, pi0377, pi0592);
  not g10904 (n_5273, n8468);
  and g10905 (n8469, n_4225, n_5273);
  and g10906 (n8470, n_5020, n8468);
  not g10907 (n_5274, n8470);
  and g10908 (n8471, n_4366, n_5274);
  not g10909 (n_5275, n8469);
  and g10910 (n8472, n_5275, n8471);
  and g10911 (n8473, n_4365, pi0592);
  not g10912 (n_5276, n8473);
  and g10913 (n8474, n_4225, n_5276);
  and g10914 (n8475, n_5020, n8473);
  not g10915 (n_5277, n8475);
  and g10916 (n8476, n7718, n_5277);
  not g10917 (n_5278, n8474);
  and g10918 (n8477, n_5278, n8476);
  not g10919 (n_5279, n8472);
  not g10920 (n_5280, n8477);
  and g10921 (n8478, n_5279, n_5280);
  not g10922 (n_5281, n8478);
  and g10923 (n8479, n7696, n_5281);
  and g10924 (n8480, pi0592, n_5020);
  and g10925 (n8481, n_4239, n_4225);
  not g10926 (n_5282, n8480);
  not g10927 (n_5283, n8481);
  and g10928 (n8482, n_5282, n_5283);
  and g10929 (n8483, n_4327, n8482);
  not g10930 (n_5284, n8479);
  not g10931 (n_5285, n8483);
  and g10932 (n8484, n_5284, n_5285);
  and g10933 (n8485, pi1199, n8484);
  and g10934 (n8486, n7636, n_4326);
  and g10935 (n8487, n7695, n8482);
  not g10936 (n_5286, n8486);
  not g10937 (n_5287, n8487);
  and g10938 (n8488, n_5286, n_5287);
  not g10939 (n_5288, n8488);
  and g10940 (n8489, n7669, n_5288);
  and g10941 (n8490, n_5024, n_4326);
  not g10942 (n_5289, n8490);
  and g10943 (n8491, n8482, n_5289);
  and g10944 (n8492, n_5024, n8486);
  not g10945 (n_5290, n8491);
  not g10946 (n_5291, n8492);
  and g10947 (n8493, n_5290, n_5291);
  not g10948 (n_5292, n8493);
  and g10949 (n8494, n_4282, n_5292);
  not g10950 (n_5293, n8489);
  and g10951 (n8495, n_4718, n_5293);
  not g10952 (n_5294, n8494);
  and g10953 (n8496, n_5294, n8495);
  not g10954 (n_5295, n8485);
  not g10955 (n_5296, n8496);
  and g10956 (n8497, n_5295, n_5296);
  not g10957 (n_5297, n8497);
  and g10958 (n8498, n_4392, n_5297);
  and g10959 (n8499, n_4377, pi1199);
  and g10960 (n8500, n8484, n8499);
  and g10961 (n8501, n_4377, n8496);
  not g10962 (n_5298, n8482);
  and g10963 (n8502, pi1198, n_5298);
  not g10964 (n_5299, n8500);
  not g10965 (n_5300, n8502);
  and g10966 (n8503, n_5299, n_5300);
  not g10967 (n_5301, n8501);
  and g10968 (n8504, n_5301, n8503);
  not g10969 (n_5302, n8504);
  and g10970 (n8505, pi0374, n_5302);
  not g10971 (n_5303, n8498);
  not g10972 (n_5304, n8505);
  and g10973 (n8506, n_5303, n_5304);
  not g10974 (n_5305, n8506);
  and g10975 (n8507, pi0369, n_5305);
  and g10976 (n8508, n_4392, n_5302);
  and g10977 (n8509, pi0374, n_5297);
  not g10978 (n_5306, n8508);
  not g10979 (n_5307, n8509);
  and g10980 (n8510, n_5306, n_5307);
  not g10981 (n_5308, n8510);
  and g10982 (n8511, n_4391, n_5308);
  not g10983 (n_5309, n8507);
  not g10984 (n_5310, n8511);
  and g10985 (n8512, n_5309, n_5310);
  not g10986 (n_5311, n8512);
  and g10987 (n8513, n_4396, n_5311);
  and g10988 (n8514, n_4391, n_5305);
  and g10989 (n8515, pi0369, n_5308);
  not g10990 (n_5312, n8514);
  not g10991 (n_5313, n8515);
  and g10992 (n8516, n_5312, n_5313);
  not g10993 (n_5314, n8516);
  and g10994 (n8517, pi0370, n_5314);
  not g10995 (n_5315, n8513);
  not g10996 (n_5316, n8517);
  and g10997 (n8518, n_5315, n_5316);
  not g10998 (n_5317, n8518);
  and g10999 (n8519, n_4401, n_5317);
  and g11000 (n8520, n_4396, n_5314);
  and g11001 (n8521, pi0370, n_5311);
  not g11002 (n_5318, n8520);
  not g11003 (n_5319, n8521);
  and g11004 (n8522, n_5318, n_5319);
  not g11005 (n_5320, n8522);
  and g11006 (n8523, pi0371, n_5320);
  not g11007 (n_5321, n8519);
  not g11008 (n_5322, n8523);
  and g11009 (n8524, n_5321, n_5322);
  not g11010 (n_5323, n8524);
  and g11011 (n8525, n_4406, n_5323);
  and g11012 (n8526, n_4401, n_5320);
  and g11013 (n8527, pi0371, n_5317);
  not g11014 (n_5324, n8526);
  not g11015 (n_5325, n8527);
  and g11016 (n8528, n_5324, n_5325);
  not g11017 (n_5326, n8528);
  and g11018 (n8529, pi0373, n_5326);
  not g11019 (n_5327, n8525);
  not g11020 (n_5328, n8529);
  and g11021 (n8530, n_5327, n_5328);
  and g11022 (n8531, n_4412, n8530);
  and g11023 (n8532, n_4406, n_5326);
  and g11024 (n8533, pi0373, n_5323);
  not g11025 (n_5329, n8532);
  not g11026 (n_5330, n8533);
  and g11027 (n8534, n_5329, n_5330);
  and g11028 (n8535, pi0375, n8534);
  not g11029 (n_5331, n8531);
  and g11030 (n8536, n7734, n_5331);
  not g11031 (n_5332, n8535);
  and g11032 (n8537, n_5332, n8536);
  and g11033 (n8538, pi0375, n8530);
  and g11034 (n8539, n_4412, n8534);
  not g11035 (n_5333, n8538);
  and g11036 (n8540, n_4415, n_5333);
  not g11037 (n_5334, n8539);
  and g11038 (n8541, n_5334, n8540);
  not g11039 (n_5335, n8537);
  and g11040 (n8542, n_4628, n_5335);
  not g11041 (n_5336, n8541);
  and g11042 (n8543, n_5336, n8542);
  not g11043 (n_5337, n8467);
  and g11044 (n8544, n_4423, n_5337);
  not g11045 (n_5338, n8543);
  and g11046 (n8545, n_5338, n8544);
  not g11047 (n_5339, n8545);
  and g11048 (n8546, n7425, n_5339);
  not g11049 (n_5340, n8393);
  and g11050 (n8547, n_5340, n8546);
  and g11051 (n8548, pi0591, n_5089);
  and g11052 (n8549, n7782, n_5104);
  and g11053 (n8550, n7825, n_5104);
  and g11054 (n8551, n7592, n_5151);
  not g11055 (n_5341, n8551);
  and g11056 (n8552, n8323, n_5341);
  and g11057 (n8553, n7592, n_5148);
  not g11058 (n_5342, n8553);
  and g11059 (n8554, n8318, n_5342);
  not g11060 (n_5343, n8552);
  and g11061 (n8555, n_4562, n_5343);
  not g11062 (n_5344, n8554);
  and g11063 (n8556, n_5344, n8555);
  not g11064 (n_5345, n8550);
  and g11065 (n8557, pi1198, n_5345);
  not g11066 (n_5346, n8556);
  and g11067 (n8558, n_5346, n8557);
  and g11068 (n8559, pi0455, n_5104);
  and g11069 (n8560, n_4480, n7592);
  not g11070 (n_5347, n8559);
  not g11071 (n_5348, n8560);
  and g11072 (n8561, n_5347, n_5348);
  not g11073 (n_5349, n8561);
  and g11074 (n8562, n_4481, n_5349);
  and g11075 (n8563, n_4480, n_5104);
  and g11076 (n8564, pi0455, n7592);
  not g11077 (n_5350, n8563);
  not g11078 (n_5351, n8564);
  and g11079 (n8565, n_5350, n_5351);
  not g11080 (n_5352, n8565);
  and g11081 (n8566, pi0452, n_5352);
  and g11082 (n8567, pi0355, n_4514);
  and g11083 (n8568, n_4485, n7815);
  not g11084 (n_5353, n8567);
  not g11085 (n_5354, n8568);
  and g11086 (n8569, n_5353, n_5354);
  not g11087 (n_5355, n8562);
  not g11088 (n_5356, n8569);
  and g11089 (n8570, n_5355, n_5356);
  not g11090 (n_5357, n8566);
  and g11091 (n8571, n_5357, n8570);
  and g11092 (n8572, n_4481, n_5352);
  and g11093 (n8573, pi0452, n_5349);
  not g11094 (n_5358, n8572);
  and g11095 (n8574, n8569, n_5358);
  not g11096 (n_5359, n8573);
  and g11097 (n8575, n_5359, n8574);
  not g11098 (n_5360, n8571);
  and g11099 (n8576, pi1196, n_5360);
  not g11100 (n_5361, n8575);
  and g11101 (n8577, n_5361, n8576);
  and g11102 (n8578, n_4377, n_5100);
  not g11103 (n_5362, n8577);
  and g11104 (n8579, n_5362, n8578);
  not g11105 (n_5363, n8558);
  and g11106 (n8580, n_4565, n_5363);
  not g11107 (n_5364, n8579);
  and g11108 (n8581, n_5364, n8580);
  not g11109 (n_5365, n8549);
  not g11110 (n_5366, n8581);
  and g11111 (n8582, n_5365, n_5366);
  not g11112 (n_5367, n8582);
  and g11113 (n8583, n_4578, n_5367);
  and g11114 (n8584, pi1199, n_5104);
  and g11115 (n8585, n_4577, n8584);
  not g11116 (n_5368, n8583);
  not g11117 (n_5369, n8585);
  and g11118 (n8586, n_5368, n_5369);
  not g11119 (n_5370, n8586);
  and g11120 (n8587, n_4575, n_5370);
  and g11121 (n8588, n_4569, n_5367);
  and g11122 (n8589, pi0351, n8584);
  not g11123 (n_5371, n8588);
  not g11124 (n_5372, n8589);
  and g11125 (n8590, n_5371, n_5372);
  not g11126 (n_5373, n8590);
  and g11127 (n8591, pi0461, n_5373);
  not g11128 (n_5374, n8587);
  not g11129 (n_5375, n8591);
  and g11130 (n8592, n_5374, n_5375);
  not g11131 (n_5376, n8592);
  and g11132 (n8593, n_4585, n_5376);
  and g11133 (n8594, n_4575, n_5373);
  and g11134 (n8595, pi0461, n_5370);
  not g11135 (n_5377, n8594);
  not g11136 (n_5378, n8595);
  and g11137 (n8596, n_5377, n_5378);
  not g11138 (n_5379, n8596);
  and g11139 (n8597, pi0357, n_5379);
  not g11140 (n_5380, n8593);
  not g11141 (n_5381, n8597);
  and g11142 (n8598, n_5380, n_5381);
  not g11143 (n_5382, n8598);
  and g11144 (n8599, n_4593, n_5382);
  and g11145 (n8600, n_4585, n_5379);
  and g11146 (n8601, pi0357, n_5376);
  not g11147 (n_5383, n8600);
  not g11148 (n_5384, n8601);
  and g11149 (n8602, n_5383, n_5384);
  not g11150 (n_5385, n8602);
  and g11151 (n8603, pi0356, n_5385);
  not g11152 (n_5386, n8599);
  not g11153 (n_5387, n8603);
  and g11154 (n8604, n_5386, n_5387);
  not g11155 (n_5388, n8604);
  and g11156 (n8605, n_4621, n_5388);
  and g11157 (n8606, n_4593, n_5385);
  and g11158 (n8607, pi0356, n_5382);
  not g11159 (n_5389, n8606);
  not g11160 (n_5390, n8607);
  and g11161 (n8608, n_5389, n_5390);
  not g11162 (n_5391, n8608);
  and g11163 (n8609, n7890, n_5391);
  not g11164 (n_5392, n8605);
  and g11165 (n8610, n_4628, n_5392);
  not g11166 (n_5393, n8609);
  and g11167 (n8611, n_5393, n8610);
  not g11168 (n_5394, n8548);
  and g11169 (n8612, pi0590, n_5394);
  not g11170 (n_5395, n8611);
  and g11171 (n8613, n_5395, n8612);
  and g11172 (n8614, n_4196, n7962);
  and g11173 (n8615, pi0038, n7961);
  not g11174 (n_5396, n8615);
  and g11175 (n8616, n_164, n_5396);
  and g11176 (n8617, n7545, n_4714);
  not g11177 (n_5397, n8617);
  and g11178 (n8618, n7550, n_5397);
  and g11179 (n8619, n_4176, n7961);
  not g11180 (n_5398, n8619);
  and g11181 (n8620, pi0299, n_5398);
  and g11182 (n8621, n_3140, n7602);
  not g11183 (n_5399, n7961);
  not g11184 (n_5400, n8621);
  and g11185 (n8622, n_5399, n_5400);
  and g11186 (n8623, n_3162, n8622);
  and g11187 (n8624, n6198, n7602);
  not g11188 (n_5401, n8624);
  and g11189 (n8625, n_5399, n_5401);
  and g11190 (n8626, n6242, n8625);
  not g11191 (n_5402, n8623);
  and g11192 (n8627, n7570, n_5402);
  not g11193 (n_5403, n8626);
  and g11194 (n8628, n_5403, n8627);
  not g11195 (n_5404, n8628);
  and g11196 (n8629, n8620, n_5404);
  and g11197 (n8630, n_4165, n7961);
  not g11198 (n_5405, n8630);
  and g11199 (n8631, n_234, n_5405);
  and g11200 (n8632, n_3119, n8622);
  and g11201 (n8633, n6205, n8625);
  not g11202 (n_5406, n8632);
  and g11203 (n8634, n7551, n_5406);
  not g11204 (n_5407, n8633);
  and g11205 (n8635, n_5407, n8634);
  not g11206 (n_5408, n8635);
  and g11207 (n8636, n8631, n_5408);
  not g11208 (n_5409, n8629);
  and g11209 (n8637, pi0039, n_5409);
  not g11210 (n_5410, n8636);
  and g11211 (n8638, n_5410, n8637);
  not g11212 (n_5411, n8618);
  not g11213 (n_5412, n8638);
  and g11214 (n8639, n_5411, n_5412);
  not g11215 (n_5413, n8639);
  and g11216 (n8640, n_161, n_5413);
  not g11217 (n_5414, n8640);
  and g11218 (n8641, n8616, n_5414);
  and g11219 (n8642, n7623, n_5399);
  not g11220 (n_5415, n8641);
  not g11221 (n_5416, n8642);
  and g11222 (n8643, n_5415, n_5416);
  not g11223 (n_5417, n8643);
  and g11224 (n8644, n_172, n_5417);
  and g11225 (n8645, n_251, n7961);
  not g11226 (n_5418, n8645);
  and g11227 (n8646, pi0087, n_5418);
  and g11228 (n8647, n7494, n_4714);
  not g11229 (n_5419, n8647);
  and g11230 (n8648, n7502, n_5419);
  not g11231 (n_5420, n8648);
  and g11232 (n8649, n8646, n_5420);
  not g11233 (n_5421, n8644);
  not g11234 (n_5422, n8649);
  and g11235 (n8650, n_5421, n_5422);
  not g11236 (n_5423, n8650);
  and g11237 (n8651, n_171, n_5423);
  and g11238 (n8652, n_4118, n7961);
  not g11239 (n_5424, n8652);
  and g11240 (n8653, pi0075, n_5424);
  not g11241 (n_5425, n7960);
  and g11242 (n8654, n_3128, n_5425);
  not g11243 (n_5426, n8654);
  and g11244 (n8655, n7483, n_5426);
  not g11245 (n_5427, n8655);
  and g11246 (n8656, n8653, n_5427);
  not g11247 (n_5428, n8651);
  not g11248 (n_5429, n8656);
  and g11249 (n8657, n_5428, n_5429);
  not g11250 (n_5430, n8657);
  and g11251 (n8658, pi0567, n_5430);
  not g11252 (n_5431, n8658);
  and g11253 (n8659, n7469, n_5431);
  not g11254 (n_5432, n8614);
  and g11255 (n8660, n7958, n_5432);
  not g11256 (n_5433, n8659);
  and g11257 (n8661, n_5433, n8660);
  and g11258 (n8662, n_4718, n_5100);
  not g11259 (n_5434, n8661);
  and g11260 (n8663, n_5434, n8662);
  and g11261 (n8664, n7484, n_4672);
  and g11262 (n8665, n8614, n8664);
  not g11263 (n_5435, n8665);
  and g11264 (n8666, n7958, n_5435);
  and g11265 (n8667, n_4196, n7929);
  and g11266 (n8668, n_4239, n_5024);
  not g11267 (n_5436, n8667);
  and g11268 (n8669, n_5436, n8668);
  not g11269 (n_5437, n8666);
  not g11270 (n_5438, n8669);
  and g11271 (n8670, n_5437, n_5438);
  not g11272 (n_5439, n7469);
  not g11273 (n_5440, n8670);
  and g11274 (n8671, n_5439, n_5440);
  and g11275 (n8672, n_4176, n7928);
  not g11276 (n_5441, n8672);
  and g11277 (n8673, pi0299, n_5441);
  not g11278 (n_5442, n8620);
  not g11279 (n_5443, n8673);
  and g11280 (n8674, n_5442, n_5443);
  and g11281 (n8675, n_4672, n7961);
  not g11282 (n_5444, n8675);
  and g11283 (n8676, n_5401, n_5444);
  and g11284 (n8677, n6242, n8676);
  and g11285 (n8678, n_5400, n_5444);
  and g11286 (n8679, n_3162, n8678);
  not g11287 (n_5445, n8677);
  and g11288 (n8680, n7570, n_5445);
  not g11289 (n_5446, n8679);
  and g11290 (n8681, n_5446, n8680);
  not g11291 (n_5447, n8674);
  not g11292 (n_5448, n8681);
  and g11293 (n8682, n_5447, n_5448);
  and g11294 (n8683, n_4165, n7928);
  not g11295 (n_5449, n8683);
  and g11296 (n8684, n_234, n_5449);
  not g11297 (n_5450, n8631);
  not g11298 (n_5451, n8684);
  and g11299 (n8685, n_5450, n_5451);
  and g11300 (n8686, n6205, n8676);
  and g11301 (n8687, n_3119, n8678);
  not g11302 (n_5452, n8686);
  and g11303 (n8688, n7551, n_5452);
  not g11304 (n_5453, n8687);
  and g11305 (n8689, n_5453, n8688);
  not g11306 (n_5454, n8685);
  not g11307 (n_5455, n8689);
  and g11308 (n8690, n_5454, n_5455);
  not g11309 (n_5456, n8682);
  and g11310 (n8691, pi0039, n_5456);
  not g11311 (n_5457, n8690);
  and g11312 (n8692, n_5457, n8691);
  and g11313 (n8693, n7520, n_4672);
  not g11314 (n_5458, n8693);
  and g11315 (n8694, pi0122, n_5458);
  not g11316 (n_5459, n8664);
  and g11317 (n8695, n_4081, n_5459);
  not g11318 (n_5460, n8695);
  and g11319 (n8696, pi1093, n_5460);
  not g11320 (n_5461, n8694);
  and g11321 (n8697, n_5461, n8696);
  not g11322 (n_5462, n8697);
  and g11323 (n8698, n7545, n_5462);
  not g11324 (n_5463, n8698);
  and g11325 (n8699, n8618, n_5463);
  not g11326 (n_5464, n8692);
  not g11327 (n_5465, n8699);
  and g11328 (n8700, n_5464, n_5465);
  not g11329 (n_5466, n8700);
  and g11330 (n8701, n_161, n_5466);
  and g11331 (n8702, pi0038, n7928);
  not g11332 (n_5467, n8702);
  and g11333 (n8703, n_164, n_5467);
  not g11334 (n_5468, n8616);
  not g11335 (n_5469, n8703);
  and g11336 (n8704, n_5468, n_5469);
  not g11337 (n_5470, n8701);
  not g11338 (n_5471, n8704);
  and g11339 (n8705, n_5470, n_5471);
  and g11340 (n8706, n_260, n8675);
  and g11341 (n8707, n_3410, n_5444);
  not g11342 (n_5472, n7620);
  and g11343 (n8708, n_5472, n8707);
  and g11344 (n8709, n6197, n_4116);
  not g11345 (n_5473, n8709);
  and g11346 (n8710, n_4115, n_5473);
  and g11347 (n8711, pi0228, n8710);
  not g11348 (n_5474, n8711);
  and g11349 (n8712, n8675, n_5474);
  and g11350 (n8713, n7470, n7619);
  and g11351 (n8714, n_3128, n_5444);
  not g11352 (n_5475, n8714);
  and g11353 (n8715, n8710, n_5475);
  and g11354 (n8716, n_4139, n8715);
  not g11355 (n_5476, n8713);
  not g11356 (n_5477, n8716);
  and g11357 (n8717, n_5476, n_5477);
  not g11358 (n_5478, n8717);
  and g11359 (n8718, pi0228, n_5478);
  not g11360 (n_5479, n8712);
  and g11361 (n8719, pi0232, n_5479);
  not g11362 (n_5480, n8718);
  and g11363 (n8720, n_5480, n8719);
  not g11364 (n_5481, n8708);
  and g11365 (n8721, n2530, n_5481);
  not g11366 (n_5482, n8720);
  and g11367 (n8722, n_5482, n8721);
  not g11368 (n_5483, n8706);
  and g11369 (n8723, pi0100, n_5483);
  not g11370 (n_5484, n8722);
  and g11371 (n8724, n_5484, n8723);
  not g11372 (n_5485, n8705);
  not g11373 (n_5486, n8724);
  and g11374 (n8725, n_5485, n_5486);
  not g11375 (n_5487, n8725);
  and g11376 (n8726, n_172, n_5487);
  and g11377 (n8727, n_251, n7928);
  not g11378 (n_5488, n8727);
  and g11379 (n8728, pi0087, n_5488);
  not g11380 (n_5489, n8646);
  not g11381 (n_5490, n8728);
  and g11382 (n8729, n_5489, n_5490);
  and g11383 (n8730, n7494, n7926);
  not g11384 (n_5491, n8730);
  and g11385 (n8731, n7502, n_5491);
  and g11386 (n8732, n_5419, n8731);
  not g11387 (n_5492, n8729);
  not g11388 (n_5493, n8732);
  and g11389 (n8733, n_5492, n_5493);
  not g11390 (n_5494, n8726);
  not g11391 (n_5495, n8733);
  and g11392 (n8734, n_5494, n_5495);
  not g11393 (n_5496, n8734);
  and g11394 (n8735, n_171, n_5496);
  and g11395 (n8736, n_4118, n7928);
  not g11396 (n_5497, n8736);
  and g11397 (n8737, pi0075, n_5497);
  not g11398 (n_5498, n8653);
  not g11399 (n_5499, n8737);
  and g11400 (n8738, n_5498, n_5499);
  and g11401 (n8739, n7483, n_5475);
  not g11402 (n_5500, n8738);
  not g11403 (n_5501, n8739);
  and g11404 (n8740, n_5500, n_5501);
  not g11405 (n_5502, n8735);
  not g11406 (n_5503, n8740);
  and g11407 (n8741, n_5502, n_5503);
  not g11408 (n_5504, n8741);
  and g11409 (n8742, n8666, n_5504);
  not g11410 (n_5505, n8731);
  and g11411 (n8743, n8728, n_5505);
  not g11412 (n_5506, n7928);
  and g11413 (n8744, n7623, n_5506);
  and g11414 (n8745, n7544, n_5463);
  and g11415 (n8746, n_5506, n_5400);
  and g11416 (n8747, n_3162, n8746);
  and g11417 (n8748, n_5506, n_5401);
  and g11418 (n8749, n6242, n8748);
  not g11419 (n_5507, n8747);
  and g11420 (n8750, n7570, n_5507);
  not g11421 (n_5508, n8749);
  and g11422 (n8751, n_5508, n8750);
  not g11423 (n_5509, n8751);
  and g11424 (n8752, n8673, n_5509);
  and g11425 (n8753, n_3119, n8746);
  and g11426 (n8754, n6205, n8748);
  not g11427 (n_5510, n8753);
  and g11428 (n8755, n7551, n_5510);
  not g11429 (n_5511, n8754);
  and g11430 (n8756, n_5511, n8755);
  not g11431 (n_5512, n8756);
  and g11432 (n8757, n8684, n_5512);
  not g11433 (n_5513, n8752);
  and g11434 (n8758, pi0039, n_5513);
  not g11435 (n_5514, n8757);
  and g11436 (n8759, n_5514, n8758);
  not g11437 (n_5515, n8745);
  not g11438 (n_5516, n8759);
  and g11439 (n8760, n_5515, n_5516);
  not g11440 (n_5517, n8760);
  and g11441 (n8761, n_161, n_5517);
  not g11442 (n_5518, n8761);
  and g11443 (n8762, n8703, n_5518);
  not g11444 (n_5519, n8744);
  not g11445 (n_5520, n8762);
  and g11446 (n8763, n_5519, n_5520);
  not g11447 (n_5521, n8763);
  and g11448 (n8764, n_172, n_5521);
  not g11449 (n_5522, n8743);
  not g11450 (n_5523, n8764);
  and g11451 (n8765, n_5522, n_5523);
  not g11452 (n_5524, n8765);
  and g11453 (n8766, n_171, n_5524);
  not g11454 (n_5525, n7927);
  and g11455 (n8767, n_3128, n_5525);
  not g11456 (n_5526, n8767);
  and g11457 (n8768, n7483, n_5526);
  not g11458 (n_5527, n8768);
  and g11459 (n8769, n8737, n_5527);
  not g11460 (n_5528, n8766);
  not g11461 (n_5529, n8769);
  and g11462 (n8770, n_5528, n_5529);
  not g11463 (n_5530, n8770);
  and g11464 (n8771, n8669, n_5530);
  not g11465 (n_5531, n8742);
  not g11466 (n_5532, n8771);
  and g11467 (n8772, n_5531, n_5532);
  not g11468 (n_5533, n8772);
  and g11469 (n8773, pi0567, n_5533);
  not g11470 (n_5534, n8671);
  and g11471 (n8774, pi1199, n_5534);
  not g11472 (n_5535, n8773);
  and g11473 (n8775, n_5535, n8774);
  not g11474 (n_5536, n8663);
  and g11475 (n8776, n_5238, n_5536);
  not g11476 (n_5537, n8775);
  and g11477 (n8777, n_5537, n8776);
  and g11478 (n8778, n8170, n8395);
  not g11479 (n_5538, n8778);
  and g11480 (n8779, n_5103, n_5538);
  not g11481 (n_5539, n8777);
  and g11482 (n8780, n_5539, n8779);
  not g11483 (n_5540, n8780);
  and g11484 (n8781, n_4723, n_5540);
  and g11485 (n8782, pi1197, n_5104);
  not g11486 (n_5541, n8781);
  not g11487 (n_5542, n8782);
  and g11488 (n8783, n_5541, n_5542);
  not g11489 (n_5543, n8783);
  and g11490 (n8784, n_4773, n_5543);
  and g11491 (n8785, pi0333, n_5540);
  not g11492 (n_5544, n8784);
  not g11493 (n_5545, n8785);
  and g11494 (n8786, n_5544, n_5545);
  not g11495 (n_5546, n8786);
  and g11496 (n8787, n_4778, n_5546);
  and g11497 (n8788, n_4773, n_5540);
  and g11498 (n8789, pi0333, n_5543);
  not g11499 (n_5547, n8788);
  not g11500 (n_5548, n8789);
  and g11501 (n8790, n_5547, n_5548);
  not g11502 (n_5549, n8790);
  and g11503 (n8791, pi0391, n_5549);
  not g11504 (n_5550, n8787);
  not g11505 (n_5551, n8791);
  and g11506 (n8792, n_5550, n_5551);
  not g11507 (n_5552, n8792);
  and g11508 (n8793, n_4785, n_5552);
  and g11509 (n8794, n_4778, n_5549);
  and g11510 (n8795, pi0391, n_5546);
  not g11511 (n_5553, n8794);
  not g11512 (n_5554, n8795);
  and g11513 (n8796, n_5553, n_5554);
  not g11514 (n_5555, n8796);
  and g11515 (n8797, pi0392, n_5555);
  not g11516 (n_5556, n8793);
  not g11517 (n_5557, n8797);
  and g11518 (n8798, n_5556, n_5557);
  and g11519 (n8799, pi0393, n8028);
  and g11520 (n8800, n_4793, n_4821);
  not g11521 (n_5558, n8799);
  not g11522 (n_5559, n8800);
  and g11523 (n8801, n_5558, n_5559);
  not g11524 (n_5560, n8798);
  not g11525 (n_5561, n8801);
  and g11526 (n8802, n_5560, n_5561);
  and g11527 (n8803, n_4785, n_5555);
  and g11528 (n8804, pi0392, n_5552);
  not g11529 (n_5562, n8803);
  not g11530 (n_5563, n8804);
  and g11531 (n8805, n_5562, n_5563);
  not g11532 (n_5564, n8805);
  and g11533 (n8806, n8801, n_5564);
  not g11534 (n_5565, n8802);
  and g11535 (n8807, pi0591, n_5565);
  not g11536 (n_5566, n8806);
  and g11537 (n8808, n_5566, n8807);
  and g11538 (n8809, n_4239, n7592);
  not g11539 (n_5567, n8809);
  and g11540 (n8810, n_5282, n_5567);
  and g11541 (n8811, n_4327, n8810);
  and g11542 (n8812, n_5089, n7696);
  not g11543 (n_5568, n8812);
  and g11544 (n8813, n_4718, n_5568);
  not g11545 (n_5569, n8811);
  and g11546 (n8814, n_5569, n8813);
  and g11547 (n8815, n7592, n_5276);
  not g11548 (n_5570, n8815);
  and g11549 (n8816, n8476, n_5570);
  and g11550 (n8817, n7592, n_5273);
  not g11551 (n_5571, n8817);
  and g11552 (n8818, n8471, n_5571);
  not g11553 (n_5572, n8816);
  not g11554 (n_5573, n8818);
  and g11555 (n8819, n_5572, n_5573);
  not g11556 (n_5574, n8819);
  and g11557 (n8820, n7696, n_5574);
  and g11558 (n8821, pi1199, n_5569);
  not g11559 (n_5575, n8820);
  and g11560 (n8822, n_5575, n8821);
  not g11561 (n_5576, n8814);
  not g11562 (n_5577, n8822);
  and g11563 (n8823, n_5576, n_5577);
  not g11564 (n_5578, n8823);
  and g11565 (n8824, n_4392, n_5578);
  and g11566 (n8825, n_4377, n_5578);
  not g11567 (n_5579, n8810);
  and g11568 (n8826, pi1198, n_5579);
  not g11569 (n_5580, n8825);
  not g11570 (n_5581, n8826);
  and g11571 (n8827, n_5580, n_5581);
  not g11572 (n_5582, n8827);
  and g11573 (n8828, pi0374, n_5582);
  not g11574 (n_5583, n8824);
  not g11575 (n_5584, n8828);
  and g11576 (n8829, n_5583, n_5584);
  not g11577 (n_5585, n8829);
  and g11578 (n8830, pi0369, n_5585);
  and g11579 (n8831, n_4392, n_5582);
  and g11580 (n8832, pi0374, n_5578);
  not g11581 (n_5586, n8831);
  not g11582 (n_5587, n8832);
  and g11583 (n8833, n_5586, n_5587);
  not g11584 (n_5588, n8833);
  and g11585 (n8834, n_4391, n_5588);
  not g11586 (n_5589, n8830);
  not g11587 (n_5590, n8834);
  and g11588 (n8835, n_5589, n_5590);
  not g11589 (n_5591, n8835);
  and g11590 (n8836, n_4396, n_5591);
  and g11591 (n8837, n_4391, n_5585);
  and g11592 (n8838, pi0369, n_5588);
  not g11593 (n_5592, n8837);
  not g11594 (n_5593, n8838);
  and g11595 (n8839, n_5592, n_5593);
  not g11596 (n_5594, n8839);
  and g11597 (n8840, pi0370, n_5594);
  not g11598 (n_5595, n8836);
  not g11599 (n_5596, n8840);
  and g11600 (n8841, n_5595, n_5596);
  not g11601 (n_5597, n8841);
  and g11602 (n8842, n_4401, n_5597);
  and g11603 (n8843, n_4396, n_5594);
  and g11604 (n8844, pi0370, n_5591);
  not g11605 (n_5598, n8843);
  not g11606 (n_5599, n8844);
  and g11607 (n8845, n_5598, n_5599);
  not g11608 (n_5600, n8845);
  and g11609 (n8846, pi0371, n_5600);
  not g11610 (n_5601, n8842);
  not g11611 (n_5602, n8846);
  and g11612 (n8847, n_5601, n_5602);
  and g11613 (n8848, pi0375, n7734);
  and g11614 (n8849, n_4412, n_4415);
  not g11615 (n_5603, n8848);
  not g11616 (n_5604, n8849);
  and g11617 (n8850, n_5603, n_5604);
  not g11618 (n_5605, n8850);
  and g11619 (n8851, pi0373, n_5605);
  and g11620 (n8852, n_4406, n8850);
  not g11621 (n_5606, n8851);
  not g11622 (n_5607, n8852);
  and g11623 (n8853, n_5606, n_5607);
  not g11624 (n_5608, n8847);
  not g11625 (n_5609, n8853);
  and g11626 (n8854, n_5608, n_5609);
  and g11627 (n8855, n_4401, n_5600);
  and g11628 (n8856, pi0371, n_5597);
  not g11629 (n_5610, n8855);
  not g11630 (n_5611, n8856);
  and g11631 (n8857, n_5610, n_5611);
  not g11632 (n_5612, n8857);
  and g11633 (n8858, n8853, n_5612);
  not g11634 (n_5613, n8854);
  and g11635 (n8859, n_4628, n_5613);
  not g11636 (n_5614, n8858);
  and g11637 (n8860, n_5614, n8859);
  not g11638 (n_5615, n8808);
  and g11639 (n8861, n_4423, n_5615);
  not g11640 (n_5616, n8860);
  and g11641 (n8862, n_5616, n8861);
  not g11642 (n_5617, n8862);
  and g11643 (n8863, n_4091, n_5617);
  not g11644 (n_5618, n8613);
  and g11645 (n8864, n_5618, n8863);
  not g11646 (n_5619, n8864);
  and g11647 (n8865, n_4832, n_5619);
  not g11648 (n_5620, n8547);
  and g11649 (n8866, n_5620, n8865);
  not g11650 (n_5621, n8312);
  and g11651 (n8867, n_4226, n_5621);
  not g11652 (n_5622, n8866);
  and g11653 (n8868, n_5622, n8867);
  not g11654 (n_5623, pi0217);
  not g11655 (n_5624, n8157);
  and g11656 (n8869, n_5623, n_5624);
  not g11657 (n_5625, n8868);
  and g11658 (n8870, n_5625, n8869);
  not g11659 (n_5626, n7641);
  and g11660 (n8871, n_5626, n7643);
  not g11661 (n_5627, n8870);
  and g11662 (n8872, n_5627, n8871);
  and g11663 (n8873, pi1161, n_4237);
  and g11664 (n8874, n2926, n8873);
  not g11665 (n_5629, pi0031);
  and g11666 (n8875, n_5629, pi1162);
  and g11667 (n8876, n8874, n8875);
  or g11668 (po0189, n8872, n8876);
  and g11669 (n8878, n2529, n3328);
  and g11670 (n8879, n_176, n_168);
  and g11671 (n8880, n8878, n8879);
  and g11672 (n8881, n6134, n8880);
  and g11673 (n8882, pi0100, n2530);
  not g11674 (n_5630, po1057);
  and g11675 (n8883, n_3214, n_5630);
  and g11676 (n8884, n6351, n8883);
  and g11677 (n8885, n_186, n8884);
  and g11678 (n8886, n_186, pi0252);
  and g11679 (n8887, pi0129, n2521);
  and g11680 (n8888, po1057, n_4117);
  not g11681 (n_5631, n8888);
  and g11682 (n8889, n6263, n_5631);
  and g11683 (n8890, n8886, n8889);
  and g11684 (n8891, n8887, n8890);
  not g11685 (n_5632, n8885);
  not g11686 (n_5633, n8891);
  and g11687 (n8892, n_5632, n_5633);
  not g11688 (n_5634, n8892);
  and g11689 (n8893, n8882, n_5634);
  and g11690 (n8894, n_4119, n_43);
  and g11691 (n8895, n6171, n8894);
  and g11692 (n8896, n2497, n2714);
  and g11693 (n8897, n2701, n8896);
  and g11694 (n8898, pi0050, n2777);
  and g11695 (n8899, n2495, n8898);
  and g11696 (n8900, n_131, n8897);
  and g11697 (n8901, n8899, n8900);
  and g11698 (n8902, n8895, n8901);
  and g11699 (n8903, pi0829, n_3206);
  and g11700 (n8904, n2932, n8903);
  or g11701 (po0840, n2928, n8904);
  not g11702 (n_5636, po0840);
  and g11703 (n8906, n_4091, n_5636);
  not g11704 (n_5637, n8906);
  and g11705 (n8907, n_186, n_5637);
  not g11706 (n_5638, n8907);
  and g11707 (n8908, n8902, n_5638);
  and g11708 (n8909, n_90, n_69);
  and g11709 (n8910, n2462, n2804);
  and g11710 (n8911, n_61, n2471);
  and g11711 (n8912, n8910, n8911);
  and g11712 (n8913, n_81, n_53);
  and g11713 (n8914, n7438, n8913);
  and g11714 (n8915, n_87, n_79);
  and g11715 (n8916, n2466, n2797);
  and g11719 (n8920, n_83, n_68);
  and g11720 (n8921, n_103, n_105);
  and g11721 (n8922, n2487, n8921);
  and g11730 (n8931, n2495, n8930);
  and g11731 (n8932, n8897, n8931);
  not g11732 (n_5639, n8932);
  and g11733 (n8933, pi0024, n_5639);
  not g11734 (n_5640, n8898);
  not g11735 (n_5641, n8930);
  and g11736 (n8934, n_5640, n_5641);
  and g11737 (n8935, n2499, n2702);
  not g11738 (n_5642, n8934);
  and g11739 (n8936, n_5642, n8935);
  not g11740 (n_5643, n8936);
  and g11741 (n8937, n_4119, n_5643);
  and g11742 (n8938, n2507, n2736);
  not g11750 (n_5646, n8908);
  not g11751 (n_5647, n8943);
  and g11752 (n8944, n_5646, n_5647);
  not g11753 (n_5648, n8944);
  and g11754 (n8945, n_142, n_5648);
  and g11755 (n8946, n_4119, n_3052);
  not g11756 (n_5649, n8946);
  and g11757 (n8947, pi0032, n_5649);
  and g11758 (n8948, n2710, n8947);
  not g11759 (n_5650, n8945);
  not g11760 (n_5651, n8948);
  and g11761 (n8949, n_5650, n_5651);
  not g11762 (n_5652, n8949);
  and g11763 (n8950, n_3066, n_5652);
  not g11764 (n_5653, n8902);
  and g11765 (n8951, n_142, n_5653);
  and g11766 (n8952, n6169, n_3067);
  not g11767 (n_5654, n8951);
  and g11768 (n8953, n_5654, n8952);
  not g11769 (n_5655, n8950);
  not g11770 (n_5656, n8953);
  and g11771 (n8954, n_5655, n_5656);
  and g11772 (n8955, n_144, n2531);
  not g11773 (n_5657, n8954);
  and g11774 (n8956, n_5657, n8955);
  not g11775 (n_5658, n8893);
  not g11776 (n_5659, n8956);
  and g11777 (n8957, n_5658, n_5659);
  not g11778 (n_5660, n8957);
  and g11779 (n8958, n2533, n_5660);
  and g11780 (n8959, n_4119, n2505);
  and g11781 (n8960, n2519, n2705);
  and g11782 (n8961, n_138, n8960);
  and g11783 (n8962, n8959, n8961);
  and g11784 (n8963, n_5636, n8962);
  and g11785 (n8964, pi0252, n_5631);
  and g11786 (n8965, n_172, n2530);
  and g11787 (n8966, pi0075, n_164);
  and g11788 (n8967, n8965, n8966);
  not g11790 (n_5661, n6282);
  not g11792 (n_5662, n8964);
  not g11795 (n_5663, n8958);
  not g11796 (n_5664, n8971);
  and g11797 (n8972, n_5663, n_5664);
  not g11798 (n_5665, n8972);
  and g11799 (po0190, n8881, n_5665);
  not g11800 (n_5668, pi0195);
  not g11801 (n_5669, pi0196);
  and g11802 (n8974, n_5668, n_5669);
  not g11803 (n_5671, pi0138);
  and g11804 (n8975, n_5671, n8974);
  not g11805 (n_5673, pi0139);
  and g11806 (n8976, n_5673, n8975);
  not g11807 (n_5675, pi0118);
  and g11808 (n8977, n_5675, n8976);
  not g11809 (n_5677, pi0079);
  and g11810 (n8978, n_5677, n8977);
  not g11811 (n_5679, pi0034);
  and g11812 (n8979, n_5679, n8978);
  not g11813 (n_5681, pi0033);
  not g11814 (n_5682, n8979);
  and g11815 (n8980, n_5681, n_5682);
  and g11816 (n8981, pi0149, pi0157);
  not g11817 (n_5685, pi0149);
  not g11818 (n_5686, pi0157);
  and g11819 (n8982, n_5685, n_5686);
  not g11820 (n_5687, n8982);
  and g11821 (n8983, n6197, n_5687);
  not g11822 (n_5688, n8981);
  and g11823 (n8984, n_5688, n8983);
  and g11824 (n8985, pi0232, n8984);
  not g11825 (n_5689, n8985);
  and g11826 (n8986, pi0075, n_5689);
  and g11827 (n8987, pi0100, n_5689);
  not g11828 (n_5690, n8986);
  not g11829 (n_5691, n8987);
  and g11830 (n8988, n_5690, n_5691);
  and g11831 (n8989, n_171, n_164);
  and g11832 (n8990, n7473, n8989);
  and g11833 (n8991, pi0164, n8990);
  not g11834 (n_5693, n8991);
  and g11835 (n8992, n8988, n_5693);
  not g11836 (n_5694, n8992);
  and g11837 (n8993, n_168, n_5694);
  and g11838 (n8994, pi0169, n8990);
  not g11839 (n_5695, n8994);
  and g11840 (n8995, n8988, n_5695);
  not g11841 (n_5696, n8995);
  and g11842 (n8996, pi0074, n_5696);
  not g11843 (n_5697, n8993);
  and g11844 (n8997, n_824, n_5697);
  not g11845 (n_5698, n8996);
  and g11846 (n8998, n_5698, n8997);
  and g11847 (n8999, pi0054, n_5694);
  and g11848 (n9000, pi0164, n7473);
  and g11849 (n9001, pi0038, n9000);
  and g11850 (n9002, n8989, n9001);
  not g11851 (n_5699, n9002);
  and g11852 (n9003, n8988, n_5699);
  not g11853 (n_5700, n8999);
  and g11854 (n9004, n_5700, n9003);
  not g11855 (n_5701, n9004);
  and g11856 (n9005, n_168, n_5701);
  not g11857 (n_5702, n9005);
  and g11858 (n9006, n_5698, n_5702);
  not g11859 (n_5703, n9006);
  and g11860 (n9007, n_3243, n_5703);
  not g11861 (n_5704, n9007);
  and g11862 (n9008, n3328, n_5704);
  not g11863 (n_5705, n8984);
  and g11864 (n9009, pi0299, n_5705);
  and g11865 (n9010, pi0178, pi0183);
  not g11866 (n_5708, pi0178);
  not g11867 (n_5709, pi0183);
  and g11868 (n9011, n_5708, n_5709);
  not g11869 (n_5710, n9011);
  and g11870 (n9012, n6197, n_5710);
  not g11871 (n_5711, n9010);
  and g11872 (n9013, n_5711, n9012);
  not g11873 (n_5712, n9013);
  and g11874 (n9014, n_234, n_5712);
  not g11875 (n_5713, n9009);
  and g11876 (n9015, pi0232, n_5713);
  not g11877 (n_5714, n9014);
  and g11878 (n9016, n_5714, n9015);
  not g11879 (n_5715, n9016);
  and g11880 (n9017, pi0100, n_5715);
  and g11881 (n9018, pi0075, n_5715);
  not g11882 (n_5716, n9017);
  not g11883 (n_5717, n9018);
  and g11884 (n9019, n_5716, n_5717);
  and g11885 (n9020, pi0191, n_234);
  and g11886 (n9021, pi0169, pi0299);
  not g11887 (n_5719, n9020);
  not g11888 (n_5720, n9021);
  and g11889 (n9022, n_5719, n_5720);
  not g11890 (n_5721, n9022);
  and g11891 (n9023, n8990, n_5721);
  not g11892 (n_5722, n9023);
  and g11893 (n9024, n9019, n_5722);
  not g11894 (n_5723, n9024);
  and g11895 (n9025, pi0074, n_5723);
  not g11896 (n_5724, n9025);
  and g11897 (n9026, n_176, n_5724);
  not g11898 (n_5726, pi0186);
  and g11899 (n9027, n_5726, n_234);
  not g11900 (n_5727, pi0164);
  and g11901 (n9028, n_5727, pi0299);
  not g11902 (n_5728, n9027);
  not g11903 (n_5729, n9028);
  and g11904 (n9029, n_5728, n_5729);
  and g11905 (n9030, n7473, n9029);
  and g11906 (n9031, n8989, n9030);
  not g11907 (n_5730, n9031);
  and g11908 (n9032, n9019, n_5730);
  not g11909 (n_5731, n9032);
  and g11910 (n9033, pi0054, n_5731);
  and g11911 (n9034, pi0038, n9030);
  not g11912 (n_5732, n9034);
  and g11913 (n9035, pi0087, n_5732);
  and g11914 (n9036, pi0216, n6379);
  and g11915 (n9037, n6243, n_3284);
  not g11916 (n_5733, n9037);
  and g11917 (n9038, pi0154, n_5733);
  and g11918 (n9039, n6243, n6396);
  not g11919 (n_5734, n9039);
  and g11920 (n9040, n_820, n_5734);
  not g11921 (n_5735, n9040);
  and g11922 (n9041, n_263, n_5735);
  not g11923 (n_5736, n9038);
  and g11924 (n9042, n_5736, n9041);
  and g11925 (n9043, n6197, n7602);
  and g11926 (n9044, n_3162, n9043);
  and g11927 (n9045, pi0152, pi0154);
  and g11928 (n9046, n9044, n9045);
  not g11929 (n_5737, n9042);
  not g11930 (n_5738, n9046);
  and g11931 (n9047, n_5737, n_5738);
  not g11932 (n_5739, n9047);
  and g11933 (n9048, n9036, n_5739);
  not g11934 (n_5740, n9048);
  and g11935 (n9049, pi0299, n_5740);
  not g11936 (n_5742, pi0176);
  and g11937 (n9050, n_5742, pi0232);
  and g11938 (n9051, pi0224, n6405);
  and g11939 (n9052, n6206, n6396);
  and g11940 (n9053, n9051, n9052);
  and g11941 (n9054, n_299, n9053);
  not g11942 (n_5743, n9054);
  and g11943 (n9055, n_234, n_5743);
  not g11944 (n_5744, n9055);
  and g11945 (n9056, n9050, n_5744);
  and g11946 (n9057, pi0176, pi0232);
  and g11947 (n9058, n6206, n9051);
  and g11948 (n9059, n7602, n9058);
  and g11949 (n9060, pi0174, n9059);
  and g11950 (n9061, n_3284, n9051);
  and g11951 (n9062, n6206, n9061);
  and g11952 (n9063, n_299, n9062);
  not g11953 (n_5745, n9060);
  and g11954 (n9064, n_234, n_5745);
  not g11955 (n_5746, n9063);
  and g11956 (n9065, n_5746, n9064);
  not g11957 (n_5747, n9065);
  and g11958 (n9066, n9057, n_5747);
  not g11959 (n_5748, n9056);
  not g11960 (n_5749, n9066);
  and g11961 (n9067, n_5748, n_5749);
  not g11962 (n_5750, n9049);
  and g11963 (n9068, pi0039, n_5750);
  not g11964 (n_5751, n9067);
  and g11965 (n9069, n_5751, n9068);
  and g11966 (n9070, n3181, n6197);
  and g11967 (n9071, pi0180, n9070);
  not g11968 (n_5752, n7432);
  and g11969 (n9072, pi0090, n_5752);
  and g11970 (n9073, n_134, n_131);
  and g11971 (n9074, n2707, n9073);
  not g11972 (n_5753, n9072);
  and g11973 (n9075, n_5753, n9074);
  and g11974 (n9076, n_68, n_91);
  and g11975 (n9077, n_90, n2468);
  and g11976 (n9078, n_95, n2467);
  and g11977 (n9079, n_97, n9077);
  and g11978 (n9080, n9078, n9079);
  and g11979 (n9081, n_53, n8921);
  and g11980 (n9082, n2466, n9081);
  and g11981 (n9083, n2464, n9082);
  and g11987 (n9089, n8935, n9088);
  and g11988 (n9090, n2487, n9089);
  not g11989 (n_5754, n9090);
  and g11990 (n9091, n6139, n_5754);
  not g11991 (n_5755, n9091);
  and g11992 (n9092, n9075, n_5755);
  and g11993 (n9093, n2518, n6197);
  and g11994 (n9094, n_143, n9093);
  and g11995 (n9095, n9092, n9094);
  and g11996 (n9096, n_5709, n9095);
  and g11997 (n9097, pi0183, n6197);
  not g11998 (n_5756, n6139);
  and g11999 (n9098, n2504, n_5756);
  and g12000 (n9099, n_5753, n9098);
  and g12001 (n9100, n2485, n9083);
  and g12002 (n9101, n_117, n9100);
  not g12003 (n_5757, n9101);
  and g12004 (n9102, pi0053, n_5757);
  and g12005 (n9103, n_117, n8898);
  not g12006 (n_5758, n9103);
  and g12007 (n9104, n2719, n_5758);
  not g12008 (n_5759, n9102);
  not g12009 (n_5760, n9104);
  and g12010 (n9105, n_5759, n_5760);
  and g12011 (n9106, n2494, n9088);
  not g12012 (n_5761, n9106);
  and g12013 (n9107, n2487, n_5761);
  not g12014 (n_5762, n9105);
  and g12015 (n9108, n_5762, n9107);
  not g12016 (n_5763, n9108);
  and g12017 (n9109, n2720, n_5763);
  and g12018 (n9110, n_43, n2717);
  and g12019 (n9111, n2504, n9110);
  and g12020 (n9112, n2723, n9111);
  and g12021 (n9113, n2487, n9112);
  and g12022 (n9114, n9109, n9113);
  not g12023 (n_5764, n9114);
  and g12024 (n9115, n_139, n_5764);
  not g12025 (n_5765, n9099);
  and g12026 (n9116, n_5765, n9115);
  and g12027 (n9117, n2519, n3100);
  not g12028 (n_5766, n9116);
  and g12029 (n9118, n_5766, n9117);
  not g12030 (n_5767, n9115);
  and g12031 (n9119, n_5767, n9117);
  not g12032 (n_5768, n6487);
  not g12033 (n_5769, n9119);
  and g12034 (n9120, n_5768, n_5769);
  not g12035 (n_5770, n9120);
  and g12036 (n9121, n_305, n_5770);
  not g12037 (n_5771, n9118);
  not g12038 (n_5772, n9121);
  and g12039 (n9122, n_5771, n_5772);
  not g12040 (n_5773, n9122);
  and g12041 (n9123, n9097, n_5773);
  not g12042 (n_5774, n9096);
  and g12043 (n9124, n_299, n_5774);
  not g12044 (n_5775, n9123);
  and g12045 (n9125, n_5775, n9124);
  and g12046 (n9126, n_5760, n9112);
  not g12047 (n_5776, n9126);
  and g12048 (n9127, n_139, n_5776);
  and g12049 (n9128, n_5765, n9127);
  not g12050 (n_5777, n9128);
  and g12051 (n9129, n9117, n_5777);
  not g12052 (n_5778, n9129);
  and g12053 (n9130, n_3387, n_5778);
  not g12054 (n_5779, n9130);
  and g12055 (n9131, n6197, n_5779);
  and g12056 (n9132, pi0183, n9131);
  and g12057 (n9133, n_5756, n9075);
  and g12058 (n9134, n9094, n9133);
  and g12059 (n9135, n_5709, n9134);
  not g12060 (n_5780, n9135);
  and g12061 (n9136, pi0174, n_5780);
  not g12062 (n_5781, n9132);
  and g12063 (n9137, n_5781, n9136);
  not g12064 (n_5782, n9125);
  not g12065 (n_5783, n9137);
  and g12066 (n9138, n_5782, n_5783);
  not g12067 (n_5785, n9138);
  and g12068 (n9139, pi0193, n_5785);
  and g12069 (n9140, n_143, n6197);
  and g12070 (n9141, n_43, n9074);
  and g12071 (n9142, n9090, n9141);
  and g12072 (n9143, n2518, n9142);
  and g12073 (n9144, n9140, n9143);
  and g12074 (n9145, n_299, n_5709);
  and g12075 (n9146, n9144, n9145);
  and g12076 (n9147, n_3387, n_5769);
  and g12077 (n9148, n_299, n9147);
  not g12078 (n_5786, n9127);
  and g12079 (n9149, n9117, n_5786);
  not g12080 (n_5787, n9149);
  and g12081 (n9150, n_3387, n_5787);
  and g12082 (n9151, pi0174, n9150);
  not g12083 (n_5788, n9151);
  and g12084 (n9152, n9097, n_5788);
  not g12085 (n_5789, n9148);
  and g12086 (n9153, n_5789, n9152);
  not g12087 (n_5790, pi0193);
  not g12088 (n_5791, n9146);
  and g12089 (n9154, n_5790, n_5791);
  not g12090 (n_5792, n9153);
  and g12091 (n9155, n_5792, n9154);
  not g12092 (n_5793, n9139);
  not g12093 (n_5794, n9155);
  and g12094 (n9156, n_5793, n_5794);
  not g12095 (n_5795, n9071);
  and g12096 (n9157, n_234, n_5795);
  not g12097 (n_5796, n9156);
  and g12098 (n9158, n_5796, n9157);
  and g12099 (n9159, n_162, pi0232);
  and g12100 (n9160, pi0158, n9070);
  and g12101 (n9161, pi0172, n9118);
  and g12102 (n9162, n_3360, n_5769);
  and g12103 (n9163, n_263, n9162);
  not g12104 (n_5797, n9161);
  and g12105 (n9164, n_5797, n9163);
  and g12106 (n9165, pi0172, n9129);
  and g12107 (n9166, n_3360, n_5787);
  not g12108 (n_5798, n9165);
  and g12109 (n9167, pi0152, n_5798);
  and g12110 (n9168, n9166, n9167);
  and g12116 (n9172, n_263, n9095);
  not g12117 (n_5801, n9134);
  not g12118 (n_5802, n9172);
  and g12119 (n9173, n_5801, n_5802);
  not g12120 (n_5803, n9173);
  and g12121 (n9174, pi0172, n_5803);
  and g12122 (n9175, n_263, n_1362);
  and g12123 (n9176, n9144, n9175);
  not g12124 (n_5804, n9174);
  not g12125 (n_5805, n9176);
  and g12126 (n9177, n_5804, n_5805);
  not g12127 (n_5806, n9177);
  and g12128 (n9178, n_5685, n_5806);
  not g12135 (n_5810, n9181);
  and g12136 (n9182, n9159, n_5810);
  not g12137 (n_5811, n9158);
  and g12138 (n9183, n_5811, n9182);
  not g12139 (n_5812, n9069);
  not g12140 (n_5813, n9183);
  and g12141 (n9184, n_5812, n_5813);
  not g12142 (n_5814, n9184);
  and g12143 (n9185, n_161, n_5814);
  and g12144 (n9186, pi0299, n7473);
  and g12145 (n9187, n_3038, n9186);
  not g12146 (n_5815, n9187);
  and g12147 (n9188, n_5726, n_5815);
  not g12148 (n_5816, n6284);
  and g12149 (n9189, n_5816, n7473);
  not g12150 (n_5817, n9189);
  and g12151 (n9190, pi0186, n_5817);
  not g12152 (n_5818, n9190);
  and g12153 (n9191, pi0164, n_5818);
  not g12154 (n_5819, n9188);
  and g12155 (n9192, n_5819, n9191);
  and g12156 (n9193, n_234, n7473);
  and g12157 (n9194, n_3038, n9193);
  and g12158 (n9195, n_5727, pi0186);
  and g12159 (n9196, n9194, n9195);
  not g12160 (n_5820, n9192);
  not g12161 (n_5821, n9196);
  and g12162 (n9197, n_5820, n_5821);
  not g12163 (n_5822, n9197);
  and g12164 (n9198, pi0038, n_5822);
  not g12165 (n_5823, n9198);
  and g12166 (n9199, n_172, n_5823);
  not g12167 (n_5824, n9185);
  and g12168 (n9200, n_5824, n9199);
  not g12169 (n_5825, n9035);
  and g12170 (n9201, n_164, n_5825);
  not g12171 (n_5826, n9200);
  and g12172 (n9202, n_5826, n9201);
  not g12173 (n_5827, n9202);
  and g12174 (n9203, n_5716, n_5827);
  not g12175 (n_5828, n9203);
  and g12176 (n9204, n2569, n_5828);
  and g12177 (n9205, n_171, pi0092);
  and g12178 (n9206, n_164, n9034);
  not g12179 (n_5829, n9206);
  and g12180 (n9207, n_5716, n_5829);
  and g12181 (n9208, n_161, n_172);
  not g12182 (n_5830, n3383);
  and g12183 (n9209, pi0232, n_5830);
  and g12184 (n9210, n_5742, n_234);
  not g12185 (n_5831, n9210);
  and g12186 (n9211, n6197, n_5831);
  and g12187 (n9212, n9209, n9211);
  not g12191 (n_5832, n9215);
  and g12192 (n9216, n9207, n_5832);
  not g12193 (n_5833, n9216);
  and g12194 (n9217, n9205, n_5833);
  not g12195 (n_5834, n9217);
  and g12196 (n9218, n_5717, n_5834);
  not g12197 (n_5835, n9204);
  and g12198 (n9219, n_5835, n9218);
  not g12199 (n_5836, n9219);
  and g12200 (n9220, n_167, n_5836);
  not g12201 (n_5837, n9033);
  not g12202 (n_5838, n9220);
  and g12203 (n9221, n_5837, n_5838);
  not g12204 (n_5839, n9221);
  and g12205 (n9222, n_168, n_5839);
  not g12206 (n_5840, n9222);
  and g12207 (n9223, n9026, n_5840);
  and g12208 (n9224, pi0055, n_5698);
  and g12209 (n9225, n_174, n_5690);
  not g12210 (n_5841, n9000);
  and g12211 (n9226, pi0038, n_5841);
  not g12212 (n_5842, n9226);
  and g12213 (n9227, n2568, n_5842);
  and g12214 (n9228, pi0149, n7473);
  and g12215 (n9229, n6135, n9228);
  not g12216 (n_5843, n9229);
  and g12217 (n9230, n_161, n_5843);
  not g12218 (n_5844, n9230);
  and g12219 (n9231, n9227, n_5844);
  and g12220 (n9232, n8161, n9001);
  not g12221 (n_5845, n9232);
  and g12222 (n9233, n_5691, n_5845);
  not g12223 (n_5846, n9231);
  and g12224 (n9234, n_5846, n9233);
  not g12225 (n_5847, n9234);
  and g12226 (n9235, n_171, n_5847);
  not g12227 (n_5848, n9235);
  and g12228 (n9236, n9225, n_5848);
  and g12229 (n9237, pi0092, n9003);
  not g12230 (n_5849, n9237);
  and g12231 (n9238, n_167, n_5849);
  not g12232 (n_5850, n9236);
  and g12233 (n9239, n_5850, n9238);
  not g12234 (n_5851, n9239);
  and g12235 (n9240, n_5700, n_5851);
  not g12236 (n_5852, n9240);
  and g12237 (n9241, n_168, n_5852);
  not g12238 (n_5853, n9241);
  and g12239 (n9242, n9224, n_5853);
  not g12240 (n_5854, n9242);
  and g12241 (n9243, n2529, n_5854);
  not g12242 (n_5855, n9223);
  and g12243 (n9244, n_5855, n9243);
  not g12244 (n_5856, n9244);
  and g12245 (n9245, n9008, n_5856);
  not g12246 (n_5857, n8998);
  not g12247 (n_5858, n9245);
  and g12248 (n9246, n_5857, n_5858);
  not g12249 (n_5859, n9246);
  and g12250 (n9247, n8980, n_5859);
  and g12251 (n9248, n_143, n2487);
  and g12252 (n9249, n_161, n9248);
  and g12253 (n9250, n8989, n9249);
  and g12254 (n9251, n2532, n9250);
  and g12255 (n9252, n_3243, n9251);
  and g12256 (n9253, n2716, n2720);
  and g12257 (n9254, n_116, n9253);
  and g12258 (n9255, n9101, n9254);
  and g12259 (n9256, n_42, n9255);
  and g12260 (n9257, n7445, n9256);
  and g12261 (n9258, n_142, n2508);
  and g12262 (n9259, n9257, n9258);
  and g12263 (n9260, n_144, n9259);
  not g12264 (n_5860, n9228);
  and g12265 (n9261, n_162, n_5860);
  and g12266 (n9262, n9260, n9261);
  not g12267 (n_5861, n9262);
  and g12268 (n9263, n9248, n_5861);
  not g12269 (n_5862, n9263);
  and g12270 (n9264, n_161, n_5862);
  not g12271 (n_5863, n9264);
  and g12272 (n9265, n9227, n_5863);
  not g12273 (n_5864, n9248);
  and g12274 (n9266, n_161, n_5864);
  not g12275 (n_5865, n9266);
  and g12276 (n9267, n_164, n_5865);
  and g12277 (n9268, n_5842, n9267);
  and g12278 (n9269, pi0087, n9268);
  not g12279 (n_5866, n9269);
  and g12280 (n9270, n_5691, n_5866);
  not g12281 (n_5867, n9265);
  and g12282 (n9271, n_5867, n9270);
  not g12283 (n_5868, n9271);
  and g12284 (n9272, n_171, n_5868);
  not g12285 (n_5869, n9272);
  and g12286 (n9273, n9225, n_5869);
  and g12287 (n9274, n_171, n9268);
  and g12288 (n9275, pi0092, n8988);
  not g12289 (n_5870, n9274);
  and g12290 (n9276, n_5870, n9275);
  not g12291 (n_5871, n9276);
  and g12292 (n9277, n_167, n_5871);
  not g12293 (n_5872, n9273);
  and g12294 (n9278, n_5872, n9277);
  not g12295 (n_5873, n9278);
  and g12296 (n9279, n_5700, n_5873);
  not g12297 (n_5874, n9279);
  and g12298 (n9280, n_168, n_5874);
  not g12299 (n_5875, n9280);
  and g12300 (n9281, n9224, n_5875);
  and g12301 (n9282, n2609, n9260);
  not g12302 (n_5876, n9212);
  and g12303 (n9283, n_5876, n9282);
  and g12304 (n9284, n2608, n9248);
  not g12305 (n_5877, n9283);
  and g12306 (n9285, n_5877, n9284);
  not g12307 (n_5878, n9285);
  and g12308 (n9286, n9207, n_5878);
  not g12309 (n_5879, n9286);
  and g12310 (n9287, n9205, n_5879);
  not g12311 (n_5880, n9284);
  and g12312 (n9288, pi0087, n_5880);
  and g12313 (n9289, n9207, n9288);
  not g12314 (n_5881, n9036);
  and g12315 (n9290, n_5881, n9248);
  not g12316 (n_5882, n9290);
  and g12317 (n9291, pi0299, n_5882);
  and g12318 (n9292, n6383, n_3286);
  and g12319 (n9293, n6212, n9292);
  not g12320 (n_5883, n6188);
  not g12321 (n_5884, n9293);
  and g12322 (n9294, n_5883, n_5884);
  not g12323 (n_5885, n9294);
  and g12324 (n9295, n9260, n_5885);
  and g12325 (n9296, n6198, n9295);
  not g12326 (n_5886, n9296);
  and g12327 (n9297, n9248, n_5886);
  and g12328 (n9298, n6197, n9295);
  not g12329 (n_5887, n9298);
  and g12330 (n9299, n9248, n_5887);
  not g12331 (n_5888, n9299);
  and g12332 (n9300, n_3162, n_5888);
  not g12333 (n_5889, n9300);
  and g12334 (n9301, n9297, n_5889);
  not g12335 (n_5890, n9301);
  and g12336 (n9302, n9291, n_5890);
  not g12337 (n_5891, n9051);
  and g12338 (n9303, n_5891, n9248);
  not g12339 (n_5892, n9297);
  not g12340 (n_5893, n9303);
  and g12341 (n9304, n_5892, n_5893);
  and g12342 (n9305, n_3119, n_5888);
  and g12343 (n9306, n_5893, n9305);
  not g12344 (n_5894, n9304);
  not g12345 (n_5895, n9306);
  and g12346 (n9307, n_5894, n_5895);
  not g12347 (n_5896, n9307);
  and g12348 (n9308, n_234, n_5896);
  not g12349 (n_5897, n9302);
  not g12350 (n_5898, n9308);
  and g12351 (n9309, n_5897, n_5898);
  not g12352 (n_5899, n9309);
  and g12353 (n9310, n_3410, n_5899);
  and g12354 (n9311, n9260, n9293);
  and g12355 (n9312, n6197, n9311);
  not g12356 (n_5900, n9312);
  and g12357 (n9313, n9248, n_5900);
  not g12358 (n_5901, n9313);
  and g12359 (n9314, n_3119, n_5901);
  and g12360 (n9315, n_5893, n9314);
  and g12361 (n9316, pi0174, n9315);
  not g12362 (n_5902, n9316);
  and g12363 (n9317, n_5894, n_5902);
  not g12364 (n_5903, n9317);
  and g12365 (n9318, n_234, n_5903);
  not g12366 (n_5904, n9311);
  and g12367 (n9319, n9248, n_5904);
  not g12368 (n_5905, n9319);
  and g12369 (n9320, n6243, n_5905);
  and g12370 (n9321, pi0152, n9320);
  not g12371 (n_5906, n9321);
  and g12372 (n9322, n9297, n_5906);
  not g12373 (n_5907, n9322);
  and g12374 (n9323, pi0154, n_5907);
  and g12375 (n9324, n6188, n9260);
  and g12376 (n9325, n_3140, n9324);
  not g12377 (n_5908, n9325);
  and g12378 (n9326, n9248, n_5908);
  and g12379 (n9327, n6197, n9326);
  and g12380 (n9328, n_263, n9327);
  and g12381 (n9329, n_820, n_5890);
  not g12382 (n_5909, n9328);
  and g12383 (n9330, n_5909, n9329);
  not g12384 (n_5910, n9323);
  and g12385 (n9331, n9036, n_5910);
  not g12386 (n_5911, n9330);
  and g12387 (n9332, n_5911, n9331);
  not g12388 (n_5912, n9332);
  and g12389 (n9333, n9291, n_5912);
  not g12390 (n_5913, n9318);
  not g12391 (n_5914, n9333);
  and g12392 (n9334, n_5913, n_5914);
  and g12393 (n9335, n6206, n9324);
  and g12394 (n9336, n9051, n9248);
  not g12395 (n_5915, n9335);
  and g12396 (n9337, n_5915, n9336);
  not g12397 (n_5916, n9337);
  and g12398 (n9338, n_5893, n_5916);
  and g12399 (n9339, n_234, n9338);
  not g12400 (n_5917, n9339);
  and g12401 (n9340, n9334, n_5917);
  not g12402 (n_5918, n9340);
  and g12403 (n9341, n9050, n_5918);
  not g12404 (n_5919, n9334);
  and g12405 (n9342, n9057, n_5919);
  not g12406 (n_5920, n9310);
  and g12412 (n9346, pi0095, n_5864);
  not g12413 (n_5923, n9346);
  and g12414 (n9347, n_145, n_5923);
  and g12415 (n9348, n_143, n_15);
  not g12416 (n_5924, n9259);
  and g12417 (n9349, n2487, n_5924);
  and g12418 (n9350, n9348, n9349);
  not g12419 (n_5925, n9347);
  not g12420 (n_5926, n9350);
  and g12421 (n9351, n_5925, n_5926);
  and g12422 (n9352, pi0032, n_5864);
  not g12423 (n_5927, n2506);
  and g12424 (n9353, n2487, n_5927);
  not g12425 (n_5928, n9257);
  and g12426 (n9354, n2487, n_5928);
  not g12427 (n_5929, n9354);
  and g12428 (n9355, pi0070, n_5929);
  not g12429 (n_5930, n9255);
  and g12430 (n9356, n2487, n_5930);
  not g12431 (n_5931, n9356);
  and g12432 (n9357, pi0058, n_5931);
  not g12433 (n_5932, n2716);
  and g12434 (n9358, n2487, n_5932);
  not g12435 (n_5933, n2720);
  and g12436 (n9359, n_3321, n_5933);
  not g12437 (n_5934, n9359);
  and g12438 (n9360, n2716, n_5934);
  not g12439 (n_5935, n9109);
  and g12440 (n9361, n_5935, n9360);
  not g12441 (n_5936, n9358);
  and g12442 (n9362, n_42, n_5936);
  not g12443 (n_5937, n9361);
  and g12444 (n9363, n_5937, n9362);
  not g12445 (n_5938, n9357);
  not g12446 (n_5939, n9363);
  and g12447 (n9364, n_5938, n_5939);
  not g12448 (n_5940, n9364);
  and g12449 (n9365, n_43, n_5940);
  and g12450 (n9366, n_3052, n9256);
  not g12451 (n_5941, n9366);
  and g12452 (n9367, n2487, n_5941);
  not g12453 (n_5942, n9367);
  and g12454 (n9368, pi0090, n_5942);
  not g12455 (n_5943, n9368);
  and g12456 (n9369, n2504, n_5943);
  not g12457 (n_5944, n9365);
  and g12458 (n9370, n_5944, n9369);
  not g12459 (n_5945, n2504);
  and g12460 (n9371, n2487, n_5945);
  not g12461 (n_5946, n9371);
  and g12462 (n9372, n_139, n_5946);
  not g12463 (n_5947, n9370);
  and g12464 (n9373, n_5947, n9372);
  not g12465 (n_5948, n9355);
  not g12466 (n_5949, n9373);
  and g12467 (n9374, n_5948, n_5949);
  not g12468 (n_5950, n9374);
  and g12469 (n9375, n_138, n_5950);
  and g12470 (n9376, pi0051, n_3321);
  not g12471 (n_5951, n9376);
  and g12472 (n9377, n2506, n_5951);
  not g12473 (n_5952, n9375);
  and g12474 (n9378, n_5952, n9377);
  not g12475 (n_5953, n9353);
  not g12476 (n_5954, n9378);
  and g12477 (n9379, n_5953, n_5954);
  not g12478 (n_5955, n9379);
  and g12479 (n9380, n_143, n_5955);
  not g12480 (n_5956, n9380);
  and g12481 (n9381, n_142, n_5956);
  not g12482 (n_5957, n9352);
  not g12483 (n_5958, n9381);
  and g12484 (n9382, n_5957, n_5958);
  not g12485 (n_5959, n9382);
  and g12486 (n9383, n_144, n_5959);
  not g12487 (n_5960, n9351);
  not g12488 (n_5961, n9383);
  and g12489 (n9384, n_5960, n_5961);
  and g12490 (n9385, n9141, n9366);
  not g12491 (n_5962, n9385);
  and g12492 (n9386, n9248, n_5962);
  not g12493 (n_5963, n9386);
  and g12494 (n9387, pi0032, n_5963);
  not g12495 (n_5964, n9387);
  and g12496 (n9388, n_5958, n_5964);
  not g12497 (n_5965, n9388);
  and g12498 (n9389, n_144, n_5965);
  and g12499 (n9390, n_305, n9389);
  not g12500 (n_5966, n9390);
  and g12501 (n9391, n9384, n_5966);
  and g12502 (n9392, n_3102, n9391);
  and g12503 (n9393, n9105, n9253);
  not g12504 (n_5967, n9393);
  and g12505 (n9394, n2487, n_5967);
  not g12506 (n_5968, n9394);
  and g12507 (n9395, n_42, n_5968);
  not g12508 (n_5969, n9395);
  and g12509 (n9396, n_5938, n_5969);
  not g12510 (n_5970, n9396);
  and g12511 (n9397, n_43, n_5970);
  not g12512 (n_5971, n9397);
  and g12513 (n9398, n9369, n_5971);
  not g12514 (n_5972, n9398);
  and g12515 (n9399, n9372, n_5972);
  not g12516 (n_5973, n9399);
  and g12517 (n9400, n_5948, n_5973);
  not g12518 (n_5974, n9400);
  and g12519 (n9401, n_138, n_5974);
  not g12520 (n_5975, n9401);
  and g12521 (n9402, n9377, n_5975);
  not g12522 (n_5976, n9402);
  and g12523 (n9403, n_5953, n_5976);
  not g12524 (n_5977, n9403);
  and g12525 (n9404, n_143, n_5977);
  not g12526 (n_5978, n9404);
  and g12527 (n9405, n_142, n_5978);
  not g12528 (n_5979, n9405);
  and g12529 (n9406, n_5964, n_5979);
  not g12530 (n_5980, n9406);
  and g12531 (n9407, n_144, n_5980);
  and g12532 (n9408, n_305, n9407);
  and g12533 (n9409, n6197, n_5923);
  and g12534 (n9410, n_5957, n_5979);
  not g12535 (n_5981, n9410);
  and g12536 (n9411, n_144, n_5981);
  not g12537 (n_5982, n9411);
  and g12538 (n9412, n9409, n_5982);
  not g12539 (n_5983, n9408);
  and g12540 (n9413, n_5983, n9412);
  not g12541 (n_5984, n9392);
  not g12542 (n_5985, n9413);
  and g12543 (n9414, n_5984, n_5985);
  not g12544 (n_5986, n9414);
  and g12545 (n9415, n_5709, n_5986);
  and g12546 (n9416, n_143, n_5957);
  not g12547 (n_5987, n6170);
  and g12548 (n9417, n2487, n_5987);
  not g12549 (n_5988, n9417);
  and g12550 (n9418, n_142, n_5988);
  and g12551 (n9419, pi0093, n_3321);
  not g12552 (n_5989, n9419);
  and g12553 (n9420, n6170, n_5989);
  and g12554 (n9421, n2487, n_5938);
  not g12555 (n_5990, n9421);
  and g12556 (n9422, n_43, n_5990);
  not g12557 (n_5991, n9422);
  and g12558 (n9423, n_5943, n_5991);
  not g12559 (n_5992, n9423);
  and g12560 (n9424, n_131, n_5992);
  not g12561 (n_5993, n9424);
  and g12562 (n9425, n9420, n_5993);
  not g12563 (n_5994, n9425);
  and g12564 (n9426, n9418, n_5994);
  not g12565 (n_5995, n9426);
  and g12566 (n9427, n9416, n_5995);
  not g12567 (n_5996, n9427);
  and g12568 (n9428, n_144, n_5996);
  not g12569 (n_5997, n9428);
  and g12570 (n9429, n9409, n_5997);
  not g12571 (n_5998, n9429);
  and g12572 (n9430, n_5984, n_5998);
  not g12573 (n_5999, n9430);
  and g12574 (n9431, pi0183, n_5999);
  not g12575 (n_6000, n9415);
  not g12576 (n_6001, n9431);
  and g12577 (n9432, n_6000, n_6001);
  and g12578 (n9433, n_144, n9432);
  and g12579 (n9434, n_299, n_5960);
  not g12580 (n_6002, n9433);
  and g12581 (n9435, n_6002, n9434);
  not g12582 (n_6003, n9097);
  not g12583 (n_6004, n9391);
  and g12584 (n9436, n_6003, n_6004);
  and g12585 (n9437, n_43, n9089);
  not g12586 (n_6005, n9437);
  and g12587 (n9438, n9423, n_6005);
  not g12588 (n_6006, n9438);
  and g12589 (n9439, n_131, n_6006);
  not g12590 (n_6007, n9439);
  and g12591 (n9440, n9420, n_6007);
  not g12592 (n_6008, n9440);
  and g12593 (n9441, n9418, n_6008);
  not g12594 (n_6009, n9441);
  and g12595 (n9442, n9416, n_6009);
  not g12596 (n_6010, n9442);
  and g12597 (n9443, n_144, n_6010);
  not g12598 (n_6011, n9443);
  and g12599 (n9444, n_5960, n_6011);
  not g12600 (n_6012, n9444);
  and g12601 (n9445, n6197, n_6012);
  and g12602 (n9446, pi0183, n9445);
  not g12603 (n_6013, n9446);
  and g12604 (n9447, pi0174, n_6013);
  not g12605 (n_6014, n9436);
  and g12606 (n9448, n_6014, n9447);
  not g12607 (n_6015, pi0180);
  not g12608 (n_6016, n9448);
  and g12609 (n9449, n_6015, n_6016);
  not g12610 (n_6017, n9435);
  and g12611 (n9450, n_6017, n9449);
  not g12612 (n_6018, n9432);
  and g12613 (n9451, n_299, n_6018);
  and g12614 (n9452, n9409, n_6011);
  not g12615 (n_6019, n9452);
  and g12616 (n9453, n_5984, n_6019);
  not g12617 (n_6020, n9453);
  and g12618 (n9454, pi0183, n_6020);
  and g12619 (n9455, n_5923, n_5961);
  and g12620 (n9456, n_5966, n9455);
  and g12621 (n9457, n9140, n9456);
  not g12622 (n_6021, n9457);
  and g12623 (n9458, n_5984, n_6021);
  not g12624 (n_6022, n9458);
  and g12625 (n9459, n_5709, n_6022);
  not g12626 (n_6023, n9454);
  not g12627 (n_6024, n9459);
  and g12628 (n9460, n_6023, n_6024);
  not g12629 (n_6025, n9460);
  and g12630 (n9461, pi0174, n_6025);
  not g12631 (n_6026, n9451);
  and g12632 (n9462, pi0180, n_6026);
  not g12633 (n_6027, n9461);
  and g12634 (n9463, n_6027, n9462);
  not g12635 (n_6028, n9450);
  not g12636 (n_6029, n9463);
  and g12637 (n9464, n_6028, n_6029);
  not g12638 (n_6030, n9464);
  and g12639 (n9465, n_5790, n_6030);
  and g12640 (n9466, n_143, n_3321);
  not g12641 (n_6031, n9466);
  and g12642 (n9467, pi0032, n_6031);
  and g12643 (n9468, n2461, n2504);
  not g12644 (n_6032, n9468);
  and g12645 (n9469, n_3321, n_6032);
  and g12646 (n9470, n7445, n9363);
  not g12647 (n_6033, n9469);
  not g12648 (n_6034, n9470);
  and g12649 (n9471, n_6033, n_6034);
  not g12650 (n_6035, n9471);
  and g12651 (n9472, n_139, n_6035);
  not g12652 (n_6036, n9472);
  and g12653 (n9473, n_5948, n_6036);
  not g12654 (n_6037, n9473);
  and g12655 (n9474, n_138, n_6037);
  not g12656 (n_6038, n9474);
  and g12657 (n9475, n9377, n_6038);
  and g12658 (n9476, n_143, n_5953);
  not g12659 (n_6039, n9475);
  and g12660 (n9477, n_6039, n9476);
  not g12661 (n_6040, n9477);
  and g12662 (n9478, n_142, n_6040);
  not g12663 (n_6041, n9467);
  not g12664 (n_6042, n9478);
  and g12665 (n9479, n_6041, n_6042);
  not g12666 (n_6043, n2736);
  and g12667 (n9480, n_6043, n_5864);
  not g12668 (n_6044, n9479);
  not g12669 (n_6045, n9480);
  and g12670 (n9481, n_6044, n_6045);
  not g12671 (n_6046, n9481);
  and g12672 (n9482, n_144, n_6046);
  not g12673 (n_6047, n9482);
  and g12674 (n9483, n_5960, n_6047);
  and g12675 (n9484, n_5923, n_6047);
  and g12676 (n9485, pi0095, n_6031);
  and g12677 (n9486, n_143, n_5963);
  not g12678 (n_6048, n9486);
  and g12679 (n9487, pi0032, n_6048);
  not g12680 (n_6049, n9487);
  and g12681 (n9488, n_6042, n_6049);
  not g12682 (n_6050, n9488);
  and g12683 (n9489, n_144, n_6050);
  not g12684 (n_6051, n9485);
  not g12685 (n_6052, n9489);
  and g12686 (n9490, n_6051, n_6052);
  not g12687 (n_6053, n9490);
  and g12688 (n9491, n9484, n_6053);
  not g12689 (n_6054, n9491);
  and g12690 (n9492, n_305, n_6054);
  not g12691 (n_6055, n9492);
  and g12692 (n9493, n6197, n_6055);
  and g12693 (n9494, n6197, n_5864);
  not g12694 (n_6056, n9493);
  not g12695 (n_6057, n9494);
  and g12696 (n9495, n_6056, n_6057);
  not g12697 (n_6058, n9495);
  and g12698 (n9496, n9483, n_6058);
  not g12699 (n_6059, n9496);
  and g12700 (n9497, n_5984, n_6059);
  not g12701 (n_6060, n9497);
  and g12702 (n9498, n_5709, n_6060);
  and g12703 (n9499, n2704, n6170);
  and g12704 (n9500, n8935, n9499);
  and g12705 (n9501, n_142, n9500);
  and g12706 (n9502, n9088, n9501);
  not g12707 (n_6061, n9502);
  and g12708 (n9503, n9248, n_6061);
  not g12709 (n_6062, n9503);
  and g12710 (n9504, n_144, n_6062);
  not g12711 (n_6063, n9504);
  and g12712 (n9505, n6197, n_6063);
  and g12713 (n9506, n_5960, n9505);
  not g12714 (n_6064, n9506);
  and g12715 (n9507, n_5984, n_6064);
  not g12716 (n_6065, n9507);
  and g12717 (n9508, pi0183, n_6065);
  not g12718 (n_6066, n9508);
  and g12719 (n9509, pi0174, n_6066);
  not g12720 (n_6067, n9498);
  and g12721 (n9510, n_6067, n9509);
  and g12722 (n9511, n_3102, n_6004);
  and g12723 (n9512, n7445, n9395);
  not g12724 (n_6068, n9512);
  and g12725 (n9513, n_6033, n_6068);
  not g12726 (n_6069, n9513);
  and g12727 (n9514, n_139, n_6069);
  not g12728 (n_6070, n9514);
  and g12729 (n9515, n_5948, n_6070);
  not g12730 (n_6071, n9515);
  and g12731 (n9516, n_138, n_6071);
  not g12732 (n_6072, n9516);
  and g12733 (n9517, n9377, n_6072);
  not g12734 (n_6073, n9517);
  and g12735 (n9518, n_5953, n_6073);
  not g12736 (n_6074, n9518);
  and g12737 (n9519, n_143, n_6074);
  not g12738 (n_6075, n9519);
  and g12739 (n9520, n_142, n_6075);
  not g12740 (n_6076, n9520);
  and g12741 (n9521, n_5957, n_6076);
  not g12742 (n_6077, n9521);
  and g12743 (n9522, n_144, n_6077);
  not g12744 (n_6078, n9522);
  and g12745 (n9523, n_5960, n_6078);
  and g12746 (n9524, n_5964, n_6076);
  not g12747 (n_6079, n9524);
  and g12748 (n9525, n_144, n_6079);
  and g12749 (n9526, n_305, n9525);
  not g12750 (n_6080, n9526);
  and g12751 (n9527, n9523, n_6080);
  not g12752 (n_6081, n9527);
  and g12753 (n9528, n6197, n_6081);
  not g12754 (n_6082, n9511);
  not g12755 (n_6083, n9528);
  and g12756 (n9529, n_6082, n_6083);
  and g12757 (n9530, n_5709, n9529);
  and g12758 (n9531, n_144, n_5864);
  not g12759 (n_6084, n9531);
  and g12760 (n9532, n_5960, n_6084);
  and g12761 (n9533, n6197, n9532);
  not g12762 (n_6085, n9533);
  and g12763 (n9534, n_5984, n_6085);
  not g12764 (n_6086, n9534);
  and g12765 (n9535, pi0183, n_6086);
  not g12766 (n_6087, n9530);
  and g12767 (n9536, n_299, n_6087);
  not g12768 (n_6088, n9535);
  and g12769 (n9537, n_6088, n9536);
  not g12770 (n_6089, n9537);
  and g12771 (n9538, n_6015, n_6089);
  not g12772 (n_6090, n9510);
  and g12773 (n9539, n_6090, n9538);
  and g12774 (n9540, n9409, n_6063);
  not g12775 (n_6091, n9540);
  and g12776 (n9541, n_5984, n_6091);
  not g12777 (n_6092, n9541);
  and g12778 (n9542, pi0183, n_6092);
  and g12779 (n9543, n9484, n9493);
  not g12780 (n_6093, n9543);
  and g12781 (n9544, n_5984, n_6093);
  not g12782 (n_6094, n9544);
  and g12783 (n9545, n_5709, n_6094);
  not g12784 (n_6095, n9542);
  and g12785 (n9546, pi0174, n_6095);
  not g12786 (n_6096, n9545);
  and g12787 (n9547, n_6096, n9546);
  and g12788 (n9548, n_6057, n_6082);
  and g12789 (n9549, pi0183, n9548);
  and g12790 (n9550, n_143, n9518);
  not g12791 (n_6097, n9550);
  and g12792 (n9551, n_142, n_6097);
  not g12793 (n_6098, n9551);
  and g12794 (n9552, n_6041, n_6098);
  not g12795 (n_6099, n9552);
  and g12796 (n9553, n_144, n_6099);
  not g12797 (n_6100, n9553);
  and g12798 (n9554, n_6051, n_6100);
  not g12799 (n_6101, n9554);
  and g12800 (n9555, pi0198, n_6101);
  and g12801 (n9556, n_6049, n_6098);
  not g12802 (n_6102, n9556);
  and g12803 (n9557, n_144, n_6102);
  not g12804 (n_6103, n9557);
  and g12805 (n9558, n_6051, n_6103);
  not g12806 (n_6104, n9558);
  and g12807 (n9559, n_305, n_6104);
  not g12808 (n_6105, n9555);
  not g12809 (n_6106, n9559);
  and g12810 (n9560, n_6105, n_6106);
  not g12811 (n_6107, n9560);
  and g12812 (n9561, n9140, n_6107);
  not g12813 (n_6108, n9561);
  and g12814 (n9562, n_5984, n_6108);
  not g12815 (n_6109, n9562);
  and g12816 (n9563, n_5709, n_6109);
  not g12817 (n_6110, n9549);
  and g12818 (n9564, n_299, n_6110);
  not g12819 (n_6111, n9563);
  and g12820 (n9565, n_6111, n9564);
  not g12821 (n_6112, n9547);
  and g12822 (n9566, pi0180, n_6112);
  not g12823 (n_6113, n9565);
  and g12824 (n9567, n_6113, n9566);
  not g12825 (n_6114, n9539);
  and g12826 (n9568, pi0193, n_6114);
  not g12827 (n_6115, n9567);
  and g12828 (n9569, n_6115, n9568);
  not g12829 (n_6116, n9465);
  not g12830 (n_6117, n9569);
  and g12831 (n9570, n_6116, n_6117);
  not g12832 (n_6118, n9570);
  and g12833 (n9571, n_234, n_6118);
  and g12834 (n9572, pi0158, pi0299);
  and g12835 (n9573, n_271, n9389);
  not g12836 (n_6119, n9573);
  and g12837 (n9574, n9384, n_6119);
  and g12838 (n9575, n_3102, n9574);
  and g12839 (n9576, n_271, n9407);
  not g12840 (n_6120, n9576);
  and g12841 (n9577, n9412, n_6120);
  not g12842 (n_6121, n9575);
  not g12843 (n_6122, n9577);
  and g12844 (n9578, n_6121, n_6122);
  not g12845 (n_6123, n9578);
  and g12846 (n9579, n_263, n_6123);
  not g12847 (n_6124, n9574);
  and g12848 (n9580, n_3102, n_6124);
  and g12849 (n9581, n9455, n_6119);
  not g12850 (n_6125, n9581);
  and g12851 (n9582, n6197, n_6125);
  not g12852 (n_6126, n9580);
  not g12853 (n_6127, n9582);
  and g12854 (n9583, n_6126, n_6127);
  and g12855 (n9584, pi0152, n9583);
  not g12856 (n_6128, n9579);
  and g12857 (n9585, n_1362, n_6128);
  not g12858 (n_6129, n9584);
  and g12859 (n9586, n_6129, n9585);
  not g12860 (n_6130, n9525);
  and g12861 (n9587, n_5923, n_6130);
  not g12862 (n_6131, n9587);
  and g12863 (n9588, n_271, n_6131);
  not g12864 (n_6132, n9588);
  and g12865 (n9589, n6197, n_6132);
  and g12866 (n9590, n_5923, n_6078);
  and g12867 (n9591, n9589, n9590);
  not g12868 (n_6133, n9591);
  and g12869 (n9592, n_6121, n_6133);
  not g12870 (n_6134, n9592);
  and g12871 (n9593, n_263, n_6134);
  and g12872 (n9594, n_271, n_6054);
  not g12873 (n_6135, n9594);
  and g12874 (n9595, n6197, n_6135);
  and g12875 (n9596, n9484, n9595);
  not g12876 (n_6136, n9596);
  and g12877 (n9597, n_6121, n_6136);
  not g12878 (n_6137, n9597);
  and g12879 (n9598, pi0152, n_6137);
  not g12880 (n_6138, n9593);
  and g12881 (n9599, pi0172, n_6138);
  not g12882 (n_6139, n9598);
  and g12883 (n9600, n_6139, n9599);
  not g12884 (n_6140, n9586);
  not g12885 (n_6141, n9600);
  and g12886 (n9601, n_6140, n_6141);
  not g12887 (n_6142, n9601);
  and g12888 (n9602, n9572, n_6142);
  not g12889 (n_6143, pi0158);
  and g12890 (n9603, n_6143, pi0299);
  and g12891 (n9604, n_5960, n_5982);
  and g12892 (n9605, n_6120, n9604);
  and g12893 (n9606, n6197, n9605);
  not g12894 (n_6144, n9606);
  and g12895 (n9607, n_263, n_6144);
  and g12896 (n9608, pi0152, n_6124);
  not g12897 (n_6145, n9607);
  and g12898 (n9609, n_1362, n_6145);
  not g12899 (n_6146, n9608);
  and g12900 (n9610, n_6146, n9609);
  not g12901 (n_6147, n9595);
  and g12902 (n9611, n_6057, n_6147);
  not g12903 (n_6148, n9611);
  and g12904 (n9612, n9483, n_6148);
  not g12905 (n_6149, n9612);
  and g12906 (n9613, pi0152, n_6149);
  not g12907 (n_6150, n9589);
  and g12908 (n9614, n_6057, n_6150);
  not g12909 (n_6151, n9614);
  and g12910 (n9615, n9523, n_6151);
  not g12911 (n_6152, n9615);
  and g12912 (n9616, n_263, n_6152);
  not g12913 (n_6153, n9616);
  and g12914 (n9617, pi0172, n_6153);
  not g12915 (n_6154, n9613);
  and g12916 (n9618, n_6154, n9617);
  not g12922 (n_6157, n9621);
  and g12923 (n9622, n_5685, n_6157);
  not g12924 (n_6158, n9602);
  and g12925 (n9623, n_6158, n9622);
  and g12926 (n9624, n_6019, n_6121);
  not g12927 (n_6159, n9624);
  and g12928 (n9625, pi0152, n_6159);
  and g12929 (n9626, n_5998, n_6121);
  not g12930 (n_6160, n9626);
  and g12931 (n9627, n_263, n_6160);
  not g12932 (n_6161, n9625);
  and g12933 (n9628, n_1362, n_6161);
  not g12934 (n_6162, n9627);
  and g12935 (n9629, n_6162, n9628);
  and g12936 (n9630, n_6091, n_6121);
  not g12937 (n_6163, n9630);
  and g12938 (n9631, pi0152, n_6163);
  and g12939 (n9632, n_6057, n_6126);
  and g12940 (n9633, n_263, n9632);
  not g12941 (n_6164, n9631);
  and g12942 (n9634, pi0172, n_6164);
  not g12943 (n_6165, n9633);
  and g12944 (n9635, n_6165, n9634);
  not g12945 (n_6166, n9629);
  not g12946 (n_6167, n9635);
  and g12947 (n9636, n_6166, n_6167);
  not g12948 (n_6168, n9636);
  and g12949 (n9637, n9572, n_6168);
  and g12950 (n9638, n_6064, n_6121);
  not g12951 (n_6169, n9638);
  and g12952 (n9639, pi0152, n_6169);
  and g12953 (n9640, n_6085, n_6121);
  not g12954 (n_6170, n9640);
  and g12955 (n9641, n_263, n_6170);
  not g12956 (n_6171, n9639);
  and g12957 (n9642, pi0172, n_6171);
  not g12958 (n_6172, n9641);
  and g12959 (n9643, n_6172, n9642);
  and g12960 (n9644, n_5960, n_5997);
  not g12961 (n_6173, n9644);
  and g12962 (n9645, n6197, n_6173);
  not g12963 (n_6174, n9645);
  and g12964 (n9646, n_6126, n_6174);
  and g12965 (n9647, n_263, n9646);
  not g12966 (n_6175, n9445);
  and g12967 (n9648, n_6175, n_6126);
  and g12968 (n9649, pi0152, n9648);
  not g12969 (n_6176, n9647);
  and g12970 (n9650, n_1362, n_6176);
  not g12971 (n_6177, n9649);
  and g12972 (n9651, n_6177, n9650);
  not g12973 (n_6178, n9643);
  not g12974 (n_6179, n9651);
  and g12975 (n9652, n_6178, n_6179);
  not g12976 (n_6180, n9652);
  and g12977 (n9653, n9603, n_6180);
  not g12978 (n_6181, n9637);
  and g12979 (n9654, pi0149, n_6181);
  not g12980 (n_6182, n9653);
  and g12981 (n9655, n_6182, n9654);
  not g12982 (n_6183, n9623);
  not g12983 (n_6184, n9655);
  and g12984 (n9656, n_6183, n_6184);
  not g12985 (n_6185, n9571);
  not g12986 (n_6186, n9656);
  and g12987 (n9657, n_6185, n_6186);
  not g12988 (n_6187, n9657);
  and g12989 (n9658, pi0232, n_6187);
  and g12990 (n9659, n_3066, n9389);
  not g12991 (n_6188, n9659);
  and g12992 (n9660, n9384, n_6188);
  not g12993 (n_6189, n9660);
  and g12994 (n9661, n_3410, n_6189);
  not g12995 (n_6190, n9661);
  and g12996 (n9662, n_162, n_6190);
  not g12997 (n_6191, n9658);
  and g12998 (n9663, n_6191, n9662);
  not g12999 (n_6192, n9345);
  not g13000 (n_6193, n9663);
  and g13001 (n9664, n_6192, n_6193);
  not g13002 (n_6194, n9664);
  and g13003 (n9665, n_161, n_6194);
  not g13004 (n_6195, n9665);
  and g13005 (n9666, n_5823, n_6195);
  not g13006 (n_6196, n9666);
  and g13007 (n9667, n_164, n_6196);
  and g13008 (n9668, n_172, n_5716);
  not g13009 (n_6197, n9667);
  and g13010 (n9669, n_6197, n9668);
  not g13011 (n_6198, n9289);
  and g13012 (n9670, n2569, n_6198);
  not g13013 (n_6199, n9669);
  and g13014 (n9671, n_6199, n9670);
  not g13015 (n_6200, n9287);
  and g13016 (n9672, n_5717, n_6200);
  not g13017 (n_6201, n9671);
  and g13018 (n9673, n_6201, n9672);
  not g13019 (n_6202, n9673);
  and g13020 (n9674, n_167, n_6202);
  not g13021 (n_6203, n9674);
  and g13022 (n9675, n_5837, n_6203);
  not g13023 (n_6204, n9675);
  and g13024 (n9676, n_168, n_6204);
  not g13025 (n_6205, n9676);
  and g13026 (n9677, n9026, n_6205);
  not g13027 (n_6206, n9281);
  and g13028 (n9678, n2529, n_6206);
  not g13029 (n_6207, n9677);
  and g13030 (n9679, n_6207, n9678);
  not g13031 (n_6208, n9252);
  and g13032 (n9680, n9008, n_6208);
  not g13033 (n_6209, n9679);
  and g13034 (n9681, n_6209, n9680);
  not g13035 (n_6210, n9681);
  and g13036 (n9682, n_5857, n_6210);
  not g13037 (n_6211, n8980);
  not g13038 (n_6212, n9682);
  and g13039 (n9683, n_6211, n_6212);
  not g13040 (n_6213, n9247);
  and g13041 (n9684, po1110, n_6213);
  not g13042 (n_6214, n9683);
  and g13043 (n9685, n_6214, n9684);
  and g13044 (n9686, pi0033, n_5859);
  and g13045 (n9687, n_5681, n_6212);
  not g13046 (n_6215, n9686);
  and g13047 (n9688, pi0954, n_6215);
  not g13048 (n_6216, n9687);
  and g13049 (n9689, n_6216, n9688);
  not g13050 (n_6217, n9685);
  not g13051 (n_6218, n9689);
  and g13052 (po0191, n_6217, n_6218);
  and g13053 (n9691, pi0197, n8982);
  not g13054 (n_6219, pi0197);
  and g13055 (n9692, n_6219, n_5687);
  not g13056 (n_6220, n9691);
  not g13057 (n_6221, n9692);
  and g13058 (n9693, n_6220, n_6221);
  and g13059 (n9694, pi0162, n6197);
  not g13060 (n_6223, n9694);
  and g13061 (n9695, n9693, n_6223);
  and g13062 (n9696, n9691, n9694);
  not g13063 (n_6224, pi0162);
  and g13064 (n9697, n_6224, n_6219);
  not g13065 (n_6225, n9697);
  and g13066 (n9698, n8983, n_6225);
  not g13067 (n_6226, n9698);
  and g13068 (n9699, n6197, n_6226);
  not g13069 (n_6227, n9696);
  and g13070 (n9700, n_6227, n9699);
  not g13071 (n_6228, n9693);
  not g13072 (n_6229, n9700);
  and g13073 (n9701, n_6228, n_6229);
  not g13074 (n_6230, n9695);
  not g13075 (n_6231, n9701);
  and g13076 (n9702, n_6230, n_6231);
  and g13077 (n9703, pi0232, n9702);
  not g13078 (n_6232, n8989);
  and g13079 (n9704, n_6232, n9703);
  and g13080 (n9705, pi0167, n7473);
  and g13081 (n9706, n8989, n9705);
  not g13082 (n_6234, n9704);
  not g13083 (n_6235, n9706);
  and g13084 (n9707, n_6234, n_6235);
  and g13085 (n9708, n_168, n9707);
  and g13086 (n9709, pi0148, n8990);
  not g13087 (n_6236, n9709);
  and g13088 (n9710, pi0074, n_6236);
  and g13089 (n9711, n_6234, n9710);
  not g13090 (n_6237, n9708);
  not g13091 (n_6238, n9711);
  and g13092 (n9712, n_6237, n_6238);
  and g13093 (n9713, n_824, n9712);
  and g13094 (n9714, n_167, n_6234);
  and g13095 (n9715, pi0038, n9706);
  not g13096 (n_6239, n9715);
  and g13097 (n9716, n9714, n_6239);
  and g13098 (n9717, n_168, n9716);
  not g13099 (n_6240, n9717);
  and g13100 (n9718, n9712, n_6240);
  not g13101 (n_6241, n9718);
  and g13102 (n9719, n_3243, n_6241);
  not g13103 (n_6242, n9719);
  and g13104 (n9720, n3328, n_6242);
  and g13105 (n9721, pi0140, pi0145);
  not g13106 (n_6244, n9721);
  and g13107 (n9722, n9011, n_6244);
  not g13108 (n_6245, pi0140);
  not g13109 (n_6246, pi0145);
  and g13110 (n9723, n_6245, n_6246);
  not g13111 (n_6247, n9723);
  and g13112 (n9724, n6197, n_6247);
  and g13113 (n9725, n9722, n9724);
  and g13114 (n9726, n_6244, n_6247);
  not g13115 (n_6248, n9726);
  and g13116 (n9727, n9012, n_6248);
  not g13117 (n_6249, n9725);
  and g13118 (n9728, n_234, n_6249);
  not g13119 (n_6250, n9727);
  and g13120 (n9729, n_6250, n9728);
  not g13121 (n_6251, n9702);
  and g13122 (n9730, pi0299, n_6251);
  not g13123 (n_6252, n9729);
  and g13124 (n9731, pi0232, n_6252);
  not g13125 (n_6253, n9730);
  and g13126 (n9732, n_6253, n9731);
  not g13127 (n_6254, n9732);
  and g13128 (n9733, pi0100, n_6254);
  and g13129 (n9734, pi0075, n_6254);
  not g13130 (n_6255, n9733);
  not g13131 (n_6256, n9734);
  and g13132 (n9735, n_6255, n_6256);
  and g13133 (n9736, pi0141, n_234);
  and g13134 (n9737, pi0148, pi0299);
  not g13135 (n_6258, n9736);
  not g13136 (n_6259, n9737);
  and g13137 (n9738, n_6258, n_6259);
  not g13138 (n_6260, n9738);
  and g13139 (n9739, n7473, n_6260);
  not g13140 (n_6261, n9739);
  and g13141 (n9740, n8989, n_6261);
  not g13142 (n_6262, n9740);
  and g13143 (n9741, n9735, n_6262);
  not g13144 (n_6263, n9741);
  and g13145 (n9742, pi0074, n_6263);
  not g13146 (n_6264, n9742);
  and g13147 (n9743, n_176, n_6264);
  and g13148 (n9744, pi0188, n_234);
  and g13149 (n9745, pi0167, pi0299);
  not g13150 (n_6266, n9744);
  not g13151 (n_6267, n9745);
  and g13152 (n9746, n_6266, n_6267);
  not g13153 (n_6268, n9746);
  and g13154 (n9747, n7473, n_6268);
  not g13155 (n_6269, n9747);
  and g13156 (n9748, n_164, n_6269);
  and g13157 (n9749, n_171, n9748);
  not g13158 (n_6270, n9749);
  and g13159 (n9750, n9735, n_6270);
  not g13160 (n_6271, n9750);
  and g13161 (n9751, pi0054, n_6271);
  not g13162 (n_6272, pi0188);
  and g13163 (n9752, n_6272, n_5815);
  and g13164 (n9753, pi0188, n9194);
  not g13165 (n_6273, pi0167);
  not g13166 (n_6274, n9753);
  and g13167 (n9754, n_6273, n_6274);
  and g13168 (n9755, pi0167, pi0188);
  and g13169 (n9756, n_5817, n9755);
  not g13170 (n_6275, n9752);
  not g13171 (n_6276, n9756);
  and g13172 (n9757, n_6275, n_6276);
  not g13173 (n_6277, n9754);
  and g13174 (n9758, n_6277, n9757);
  not g13175 (n_6278, n9758);
  and g13176 (n9759, pi0038, n_6278);
  and g13177 (n9760, n_161, pi0155);
  not g13178 (n_6280, n9044);
  and g13179 (n9761, pi0161, n_6280);
  and g13180 (n9762, n_264, n_5733);
  not g13181 (n_6281, n9762);
  and g13182 (n9763, n9036, n_6281);
  not g13183 (n_6282, n9761);
  and g13184 (n9764, n_6282, n9763);
  not g13185 (n_6283, n9764);
  and g13186 (n9765, n9760, n_6283);
  not g13187 (n_6284, pi0155);
  and g13188 (n9766, n_161, n_6284);
  and g13189 (n9767, n_264, n9036);
  and g13190 (n9768, n9039, n9767);
  not g13191 (n_6285, n9768);
  and g13192 (n9769, n9766, n_6285);
  not g13193 (n_6286, n9765);
  not g13194 (n_6287, n9769);
  and g13195 (n9770, n_6286, n_6287);
  not g13196 (n_6288, n9770);
  and g13197 (n9771, pi0299, n_6288);
  not g13198 (n_6290, pi0177);
  and g13199 (n9772, n_6290, n_234);
  and g13200 (n9773, n_298, n9053);
  not g13201 (n_6291, n9773);
  and g13202 (n9774, n9772, n_6291);
  and g13203 (n9775, n_298, n9062);
  and g13204 (n9776, pi0177, n_234);
  and g13205 (n9777, pi0144, n9059);
  not g13206 (n_6292, n9777);
  and g13207 (n9778, n9776, n_6292);
  not g13208 (n_6293, n9775);
  and g13209 (n9779, n_6293, n9778);
  not g13210 (n_6294, n9774);
  and g13211 (n9780, pi0232, n_6294);
  not g13212 (n_6295, n9779);
  and g13213 (n9781, n_6295, n9780);
  not g13214 (n_6296, n9781);
  and g13215 (n9782, n_161, n_6296);
  not g13216 (n_6297, n9771);
  not g13217 (n_6298, n9782);
  and g13218 (n9783, n_6297, n_6298);
  not g13219 (n_6299, n9783);
  and g13220 (n9784, pi0039, n_6299);
  not g13221 (n_6300, n9095);
  and g13222 (n9785, n_268, n_6300);
  not g13223 (n_6301, n9144);
  and g13224 (n9786, pi0146, n_6301);
  not g13225 (n_6302, n9786);
  and g13226 (n9787, n_264, n_6302);
  not g13227 (n_6303, n9785);
  and g13228 (n9788, n_6303, n9787);
  and g13229 (n9789, n_268, pi0161);
  and g13230 (n9790, n9134, n9789);
  not g13231 (n_6304, n9788);
  not g13232 (n_6305, n9790);
  and g13233 (n9791, n_6304, n_6305);
  not g13234 (n_6306, n9791);
  and g13235 (n9792, n_6224, n_6306);
  not g13236 (n_6307, pi0159);
  and g13237 (n9793, n_6307, pi0299);
  and g13238 (n9794, pi0159, pi0299);
  and g13239 (n9795, n_6224, n9070);
  not g13240 (n_6308, n9795);
  and g13241 (n9796, n9794, n_6308);
  not g13242 (n_6309, n9793);
  not g13243 (n_6310, n9796);
  and g13244 (n9797, n_6309, n_6310);
  not g13245 (n_6311, n9797);
  and g13246 (n9798, n_6223, n_6311);
  and g13247 (n9799, pi0159, n3181);
  and g13248 (n9800, n_268, n9129);
  not g13249 (n_6312, n9800);
  and g13250 (n9801, n9166, n_6312);
  not g13251 (n_6313, n9801);
  and g13252 (n9802, pi0161, n_6313);
  and g13253 (n9803, n_268, n9118);
  not g13254 (n_6314, n9803);
  and g13255 (n9804, n9162, n_6314);
  not g13256 (n_6315, n9804);
  and g13257 (n9805, n_264, n_6315);
  not g13264 (n_6319, n9798);
  not g13265 (n_6320, n9808);
  and g13266 (n9809, n_6319, n_6320);
  not g13267 (n_6321, n9792);
  not g13268 (n_6322, n9809);
  and g13269 (n9810, n_6321, n_6322);
  and g13270 (n9811, pi0181, n9070);
  and g13271 (n9812, pi0140, n_3102);
  and g13272 (n9813, n_738, n9134);
  not g13273 (n_6323, n9813);
  and g13274 (n9814, n_6245, n_6323);
  and g13275 (n9815, n_738, n9129);
  not g13276 (n_6324, n9815);
  and g13277 (n9816, pi0140, n_6324);
  and g13278 (n9817, n9150, n9816);
  not g13279 (n_6325, n9814);
  not g13280 (n_6326, n9817);
  and g13281 (n9818, n_6325, n_6326);
  not g13282 (n_6327, n9818);
  and g13283 (n9819, pi0144, n_6327);
  and g13284 (n9820, n_738, n9095);
  and g13285 (n9821, pi0142, n9144);
  not g13286 (n_6328, n9821);
  and g13287 (n9822, n_6245, n_6328);
  not g13288 (n_6329, n9820);
  and g13289 (n9823, n_6329, n9822);
  and g13290 (n9824, n_738, n9118);
  and g13291 (n9825, pi0140, n9147);
  not g13292 (n_6330, n9824);
  and g13293 (n9826, n_6330, n9825);
  not g13294 (n_6331, n9823);
  not g13295 (n_6332, n9826);
  and g13296 (n9827, n_6331, n_6332);
  not g13297 (n_6333, n9827);
  and g13298 (n9828, n_298, n_6333);
  not g13299 (n_6334, n9812);
  not g13300 (n_6335, n9819);
  and g13301 (n9829, n_6334, n_6335);
  not g13302 (n_6336, n9828);
  and g13303 (n9830, n_6336, n9829);
  not g13304 (n_6337, n9811);
  and g13305 (n9831, n_234, n_6337);
  not g13306 (n_6338, n9830);
  and g13307 (n9832, n_6338, n9831);
  not g13308 (n_6339, n9810);
  and g13309 (n9833, pi0232, n_6339);
  not g13310 (n_6340, n9832);
  and g13311 (n9834, n_6340, n9833);
  not g13312 (n_6341, n9834);
  and g13313 (n9835, n2530, n_6341);
  not g13314 (n_6342, n9759);
  not g13315 (n_6343, n9784);
  and g13316 (n9836, n_6342, n_6343);
  not g13317 (n_6344, n9835);
  and g13318 (n9837, n_6344, n9836);
  not g13319 (n_6345, n9837);
  and g13320 (n9838, n_164, n_6345);
  not g13321 (n_6346, n9838);
  and g13322 (n9839, n_6255, n_6346);
  not g13323 (n_6347, n9839);
  and g13324 (n9840, n_172, n_6347);
  not g13325 (n_6348, n9748);
  and g13326 (n9841, n_958, n_6348);
  and g13327 (n9842, n_6255, n9841);
  not g13328 (n_6349, n9842);
  and g13329 (n9843, pi0087, n_6349);
  not g13330 (n_6350, n9840);
  not g13331 (n_6351, n9843);
  and g13332 (n9844, n_6350, n_6351);
  not g13333 (n_6352, n9844);
  and g13334 (n9845, n2569, n_6352);
  and g13335 (n9846, pi0038, n_6268);
  and g13336 (n9847, pi0155, pi0299);
  not g13337 (n_6353, n9776);
  not g13338 (n_6354, n9847);
  and g13339 (n9848, n_6353, n_6354);
  not g13340 (n_6355, n9848);
  and g13341 (n9849, n2530, n_6355);
  and g13342 (n9850, n2512, n9849);
  not g13343 (n_6356, n9846);
  not g13344 (n_6357, n9850);
  and g13345 (n9851, n_6356, n_6357);
  not g13346 (n_6358, n9851);
  and g13347 (n9852, n7473, n_6358);
  not g13348 (n_6359, n9852);
  and g13349 (n9853, n_164, n_6359);
  not g13350 (n_6360, n9853);
  and g13351 (n9854, n_6255, n_6360);
  not g13352 (n_6361, n9854);
  and g13353 (n9855, n_172, n_6361);
  not g13354 (n_6362, n9855);
  and g13355 (n9856, n_6351, n_6362);
  not g13356 (n_6363, n9856);
  and g13357 (n9857, n9205, n_6363);
  not g13358 (n_6364, n9857);
  and g13359 (n9858, n_6256, n_6364);
  not g13360 (n_6365, n9845);
  and g13361 (n9859, n_6365, n9858);
  not g13362 (n_6366, n9859);
  and g13363 (n9860, n_167, n_6366);
  not g13364 (n_6367, n9751);
  not g13365 (n_6368, n9860);
  and g13366 (n9861, n_6367, n_6368);
  not g13367 (n_6369, n9861);
  and g13368 (n9862, n_168, n_6369);
  not g13369 (n_6370, n9862);
  and g13370 (n9863, n9743, n_6370);
  and g13371 (n9864, pi0055, n_6238);
  and g13372 (n9865, pi0054, n9707);
  and g13373 (n9866, pi0038, n9705);
  not g13378 (n_6371, n9866);
  not g13379 (n_6372, n9870);
  and g13380 (n9871, n_6371, n_6372);
  not g13381 (n_6373, n9871);
  and g13382 (n9872, n8989, n_6373);
  not g13383 (n_6374, n9872);
  and g13384 (n9873, n9714, n_6374);
  not g13385 (n_6375, n9865);
  not g13386 (n_6376, n9873);
  and g13387 (n9874, n_6375, n_6376);
  not g13388 (n_6377, n9874);
  and g13389 (n9875, n_168, n_6377);
  not g13390 (n_6378, n9875);
  and g13391 (n9876, n9864, n_6378);
  not g13392 (n_6379, n9876);
  and g13393 (n9877, n2529, n_6379);
  not g13394 (n_6380, n9863);
  and g13395 (n9878, n_6380, n9877);
  not g13396 (n_6381, n9878);
  and g13397 (n9879, n9720, n_6381);
  not g13398 (n_6382, n9713);
  not g13399 (n_6383, n9879);
  and g13400 (n9880, n_6382, n_6383);
  and g13401 (n9881, pi0034, n9880);
  not g13402 (n_6384, n9251);
  and g13403 (n9882, n_3243, n_6384);
  not g13404 (n_6385, n9882);
  and g13405 (n9883, n3328, n_6385);
  not g13406 (n_6386, n9720);
  not g13407 (n_6387, n9883);
  and g13408 (n9884, n_6386, n_6387);
  not g13409 (n_6388, n9250);
  and g13410 (n9885, n_6388, n9716);
  not g13411 (n_6389, n6134);
  not g13412 (n_6390, n9885);
  and g13413 (n9886, n_6389, n_6390);
  not g13414 (n_6391, n9703);
  and g13415 (n9887, pi0075, n_6391);
  and g13416 (n9888, pi0100, n_6391);
  and g13417 (n9889, n9282, n_6223);
  not g13418 (n_6392, n9889);
  and g13419 (n9890, n9249, n_6392);
  not g13420 (n_6393, n9890);
  and g13421 (n9891, n_164, n_6393);
  and g13422 (n9892, n_3410, n9282);
  not g13423 (n_6394, n9891);
  not g13424 (n_6395, n9892);
  and g13425 (n9893, n_6394, n_6395);
  not g13426 (n_6396, n9893);
  and g13427 (n9894, n_6371, n_6396);
  not g13428 (n_6397, n9888);
  not g13429 (n_6398, n9894);
  and g13430 (n9895, n_6397, n_6398);
  not g13431 (n_6399, n9895);
  and g13432 (n9896, n_171, n_6399);
  not g13433 (n_6400, n9887);
  and g13434 (n9897, n_174, n_6400);
  not g13435 (n_6401, n9896);
  and g13436 (n9898, n_6401, n9897);
  not g13437 (n_6402, n9886);
  not g13438 (n_6403, n9898);
  and g13439 (n9899, n_6402, n_6403);
  not g13440 (n_6404, n9899);
  and g13441 (n9900, n_6375, n_6404);
  not g13442 (n_6405, n9900);
  and g13443 (n9901, n_168, n_6405);
  not g13444 (n_6406, n9901);
  and g13445 (n9902, n9864, n_6406);
  and g13446 (n9903, pi0146, n9646);
  and g13447 (n9904, n_268, n_6170);
  not g13448 (n_6407, n9903);
  and g13449 (n9905, n_264, n_6407);
  not g13450 (n_6408, n9904);
  and g13451 (n9906, n_6408, n9905);
  and g13452 (n9907, pi0146, n9648);
  and g13453 (n9908, n_268, n_6169);
  not g13454 (n_6409, n9907);
  and g13455 (n9909, pi0161, n_6409);
  not g13456 (n_6410, n9908);
  and g13457 (n9910, n_6410, n9909);
  not g13458 (n_6411, n9906);
  not g13459 (n_6412, n9910);
  and g13460 (n9911, n_6411, n_6412);
  not g13461 (n_6413, n9911);
  and g13462 (n9912, pi0162, n_6413);
  and g13463 (n9913, n_264, n_6144);
  and g13464 (n9914, pi0161, n_6124);
  not g13465 (n_6414, n9913);
  and g13466 (n9915, pi0146, n_6414);
  not g13467 (n_6415, n9914);
  and g13468 (n9916, n_6415, n9915);
  and g13469 (n9917, n_264, n_6152);
  and g13470 (n9918, pi0161, n_6149);
  not g13471 (n_6416, n9917);
  and g13472 (n9919, n_268, n_6416);
  not g13473 (n_6417, n9918);
  and g13474 (n9920, n_6417, n9919);
  not g13480 (n_6420, n9912);
  not g13481 (n_6421, n9923);
  and g13482 (n9924, n_6420, n_6421);
  not g13483 (n_6422, n9924);
  and g13484 (n9925, n9793, n_6422);
  and g13485 (n9926, pi0142, n9391);
  and g13486 (n9927, n_738, n_6060);
  not g13487 (n_6423, n9926);
  and g13488 (n9928, n_6245, n_6423);
  not g13489 (n_6424, n9927);
  and g13490 (n9929, n_6424, n9928);
  and g13491 (n9930, pi0142, n_6175);
  and g13492 (n9931, n_6082, n9930);
  and g13493 (n9932, n_738, n_6065);
  not g13494 (n_6425, n9931);
  and g13495 (n9933, pi0140, n_6425);
  not g13496 (n_6426, n9932);
  and g13497 (n9934, n_6426, n9933);
  not g13498 (n_6427, n9929);
  not g13499 (n_6428, n9934);
  and g13500 (n9935, n_6427, n_6428);
  not g13501 (n_6429, pi0181);
  not g13502 (n_6430, n9935);
  and g13503 (n9936, n_6429, n_6430);
  and g13504 (n9937, n_738, n_6094);
  and g13505 (n9938, pi0142, n_6022);
  not g13506 (n_6431, n9938);
  and g13507 (n9939, n_6245, n_6431);
  not g13508 (n_6432, n9937);
  and g13509 (n9940, n_6432, n9939);
  and g13510 (n9941, pi0142, n_6020);
  and g13511 (n9942, n_738, n_6092);
  not g13512 (n_6433, n9941);
  and g13513 (n9943, pi0140, n_6433);
  not g13514 (n_6434, n9942);
  and g13515 (n9944, n_6434, n9943);
  not g13516 (n_6435, n9940);
  not g13517 (n_6436, n9944);
  and g13518 (n9945, n_6435, n_6436);
  not g13519 (n_6437, n9945);
  and g13520 (n9946, pi0181, n_6437);
  not g13521 (n_6438, n9946);
  and g13522 (n9947, pi0144, n_6438);
  not g13523 (n_6439, n9936);
  and g13524 (n9948, n_6439, n9947);
  and g13525 (n9949, n_5983, n9604);
  not g13526 (n_6440, n9949);
  and g13527 (n9950, n6197, n_6440);
  not g13528 (n_6441, n9950);
  and g13529 (n9951, pi0142, n_6441);
  and g13530 (n9952, n_6082, n9951);
  and g13531 (n9953, n_738, n9529);
  not g13532 (n_6442, n9952);
  and g13533 (n9954, n_6245, n_6442);
  not g13534 (n_6443, n9953);
  and g13535 (n9955, n_6443, n9954);
  and g13536 (n9956, pi0142, n_6174);
  and g13537 (n9957, n_6082, n9956);
  and g13538 (n9958, n_738, n_6086);
  not g13539 (n_6444, n9957);
  and g13540 (n9959, pi0140, n_6444);
  not g13541 (n_6445, n9958);
  and g13542 (n9960, n_6445, n9959);
  not g13543 (n_6446, n9955);
  not g13544 (n_6447, n9960);
  and g13545 (n9961, n_6446, n_6447);
  not g13546 (n_6448, n9961);
  and g13547 (n9962, n_6429, n_6448);
  and g13548 (n9963, pi0142, n_5986);
  and g13549 (n9964, n_738, n_6109);
  not g13550 (n_6449, n9963);
  and g13551 (n9965, n_6245, n_6449);
  not g13552 (n_6450, n9964);
  and g13553 (n9966, n_6450, n9965);
  and g13554 (n9967, n_738, n9548);
  and g13555 (n9968, pi0142, n_5999);
  not g13556 (n_6451, n9967);
  and g13557 (n9969, pi0140, n_6451);
  not g13558 (n_6452, n9968);
  and g13559 (n9970, n_6452, n9969);
  not g13560 (n_6453, n9966);
  not g13561 (n_6454, n9970);
  and g13562 (n9971, n_6453, n_6454);
  not g13563 (n_6455, n9971);
  and g13564 (n9972, pi0181, n_6455);
  not g13565 (n_6456, n9962);
  and g13566 (n9973, n_298, n_6456);
  not g13567 (n_6457, n9972);
  and g13568 (n9974, n_6457, n9973);
  not g13569 (n_6458, n9974);
  and g13570 (n9975, n_234, n_6458);
  not g13571 (n_6459, n9948);
  and g13572 (n9976, n_6459, n9975);
  and g13573 (n9977, pi0146, n9583);
  and g13574 (n9978, n_268, n_6137);
  not g13575 (n_6460, n9977);
  and g13576 (n9979, pi0161, n_6460);
  not g13577 (n_6461, n9978);
  and g13578 (n9980, n_6461, n9979);
  and g13579 (n9981, pi0146, n_6123);
  and g13580 (n9982, n_268, n_6134);
  not g13581 (n_6462, n9981);
  and g13582 (n9983, n_264, n_6462);
  not g13583 (n_6463, n9982);
  and g13584 (n9984, n_6463, n9983);
  not g13585 (n_6464, n9980);
  and g13586 (n9985, n_6224, n_6464);
  not g13587 (n_6465, n9984);
  and g13588 (n9986, n_6465, n9985);
  and g13589 (n9987, n_268, n9632);
  and g13590 (n9988, pi0146, n_6160);
  not g13591 (n_6466, n9987);
  and g13592 (n9989, n_264, n_6466);
  not g13593 (n_6467, n9988);
  and g13594 (n9990, n_6467, n9989);
  and g13595 (n9991, pi0146, n_6159);
  and g13596 (n9992, n_268, n_6163);
  not g13597 (n_6468, n9991);
  and g13598 (n9993, pi0161, n_6468);
  not g13599 (n_6469, n9992);
  and g13600 (n9994, n_6469, n9993);
  not g13601 (n_6470, n9990);
  and g13602 (n9995, pi0162, n_6470);
  not g13603 (n_6471, n9994);
  and g13604 (n9996, n_6471, n9995);
  not g13605 (n_6472, n9986);
  and g13606 (n9997, n9794, n_6472);
  not g13607 (n_6473, n9996);
  and g13608 (n9998, n_6473, n9997);
  not g13609 (n_6474, n9925);
  not g13610 (n_6475, n9998);
  and g13611 (n9999, n_6474, n_6475);
  not g13612 (n_6476, n9976);
  and g13613 (n10000, n_6476, n9999);
  not g13614 (n_6477, n10000);
  and g13615 (n10001, pi0232, n_6477);
  not g13616 (n_6478, n10001);
  and g13617 (n10002, n_6190, n_6478);
  not g13618 (n_6479, n10002);
  and g13619 (n10003, n2530, n_6479);
  and g13620 (n10004, pi0144, n9307);
  and g13621 (n10005, n_298, n_5894);
  not g13622 (n_6480, n9338);
  and g13623 (n10006, n_6480, n10005);
  not g13624 (n_6481, n10006);
  and g13625 (n10007, n9772, n_6481);
  not g13626 (n_6482, n10004);
  and g13627 (n10008, n_6482, n10007);
  not g13628 (n_6483, n9315);
  and g13629 (n10009, n_5894, n_6483);
  not g13630 (n_6484, n10005);
  and g13631 (n10010, n9776, n_6484);
  not g13632 (n_6485, n10009);
  and g13633 (n10011, n_6485, n10010);
  not g13634 (n_6486, n10008);
  not g13635 (n_6487, n10011);
  and g13636 (n10012, n_6486, n_6487);
  not g13637 (n_6488, n10012);
  and g13638 (n10013, pi0232, n_6488);
  not g13639 (n_6489, n10013);
  and g13640 (n10014, n_5920, n_6489);
  not g13641 (n_6490, n10014);
  and g13642 (n10015, n_161, n_6490);
  and g13643 (n10016, n_264, n9327);
  not g13644 (n_6491, n10016);
  and g13645 (n10017, n_5890, n_6491);
  not g13646 (n_6492, n10017);
  and g13647 (n10018, n9036, n_6492);
  and g13648 (n10019, n9291, n9766);
  not g13649 (n_6493, n10018);
  and g13650 (n10020, n_6493, n10019);
  and g13651 (n10021, pi0161, n9320);
  and g13652 (n10022, n9036, n9297);
  not g13653 (n_6494, n10021);
  and g13654 (n10023, n_6494, n10022);
  and g13655 (n10024, n9291, n9760);
  not g13656 (n_6495, n10023);
  and g13657 (n10025, n_6495, n10024);
  not g13658 (n_6496, n10020);
  not g13659 (n_6497, n10025);
  and g13660 (n10026, n_6496, n_6497);
  not g13661 (n_6498, n10026);
  and g13662 (n10027, pi0232, n_6498);
  not g13663 (n_6499, n10015);
  not g13664 (n_6500, n10027);
  and g13665 (n10028, n_6499, n_6500);
  not g13666 (n_6501, n10028);
  and g13667 (n10029, pi0039, n_6501);
  and g13673 (n10033, pi0038, n_6269);
  not g13674 (n_6504, n10033);
  and g13675 (n10034, n_5865, n_6504);
  and g13676 (n10035, pi0087, n10034);
  not g13677 (n_6505, n10035);
  and g13678 (n10036, n_164, n_6505);
  not g13679 (n_6506, n10032);
  and g13680 (n10037, n_6506, n10036);
  not g13681 (n_6507, n10037);
  and g13682 (n10038, n_6255, n_6507);
  not g13683 (n_6508, n10038);
  and g13684 (n10039, n2569, n_6508);
  and g13685 (n10040, n_161, n9848);
  not g13686 (n_6509, n10040);
  and g13687 (n10041, n7473, n_6509);
  not g13688 (n_6510, n10041);
  and g13689 (n10042, n9282, n_6510);
  not g13690 (n_6511, n10042);
  and g13691 (n10043, n10034, n_6511);
  not g13692 (n_6512, n10043);
  and g13693 (n10044, n_164, n_6512);
  not g13694 (n_6513, n10044);
  and g13695 (n10045, n_6255, n_6513);
  not g13696 (n_6514, n10045);
  and g13697 (n10046, n9205, n_6514);
  not g13698 (n_6515, n10046);
  and g13699 (n10047, n_6256, n_6515);
  not g13700 (n_6516, n10039);
  and g13701 (n10048, n_6516, n10047);
  not g13702 (n_6517, n10048);
  and g13703 (n10049, n_167, n_6517);
  not g13704 (n_6518, n10049);
  and g13705 (n10050, n_6367, n_6518);
  not g13706 (n_6519, n10050);
  and g13707 (n10051, n_168, n_6519);
  not g13708 (n_6520, n10051);
  and g13709 (n10052, n9743, n_6520);
  not g13710 (n_6521, n9902);
  and g13711 (n10053, n2529, n_6521);
  not g13712 (n_6522, n10052);
  and g13713 (n10054, n_6522, n10053);
  not g13714 (n_6523, n9884);
  not g13715 (n_6524, n10054);
  and g13716 (n10055, n_6523, n_6524);
  not g13717 (n_6525, n10055);
  and g13718 (n10056, n_6382, n_6525);
  and g13719 (n10057, n_5679, n10056);
  and g13720 (n10058, n_5681, po1110);
  not g13721 (n_6526, n9881);
  not g13722 (n_6527, n10058);
  and g13723 (n10059, n_6526, n_6527);
  not g13724 (n_6528, n10057);
  and g13725 (n10060, n_6528, n10059);
  not g13726 (n_6529, n8978);
  and g13727 (n10061, n_5679, n_6529);
  and g13728 (n10062, n9880, n10061);
  not g13729 (n_6530, n10061);
  and g13730 (n10063, n10056, n_6530);
  not g13731 (n_6531, n10062);
  and g13732 (n10064, n10058, n_6531);
  not g13733 (n_6532, n10063);
  and g13734 (n10065, n_6532, n10064);
  not g13735 (n_6533, n10060);
  not g13736 (n_6534, n10065);
  and g13737 (po0192, n_6533, n_6534);
  and g13738 (n10067, n2529, n2572);
  and g13739 (n10068, n8962, n10067);
  and g13740 (n10069, n_176, n10068);
  not g13741 (n_6535, n10069);
  and g13742 (n10070, pi0059, n_6535);
  and g13743 (n10071, n_4119, n7340);
  not g13744 (n_6536, n10071);
  and g13745 (n10072, pi0054, n_6536);
  and g13746 (n10073, pi0137, n8884);
  and g13747 (n10074, n2923, n2930);
  not g13748 (n_6537, n10074);
  and g13749 (n10075, n7417, n_6537);
  and g13750 (n10076, pi0683, n10075);
  and g13751 (n10077, pi0252, po1057);
  not g13752 (n_6538, n10076);
  and g13753 (n10078, n_6538, n10077);
  and g13754 (n10079, pi0146, n7471);
  and g13755 (n10080, pi0142, n7470);
  not g13756 (n_6539, n10079);
  not g13757 (n_6540, n10080);
  and g13758 (n10081, n_6539, n_6540);
  not g13759 (n_6541, n7472);
  and g13760 (n10082, n_6541, n10081);
  not g13761 (n_6542, n10078);
  not g13762 (n_6543, n10082);
  and g13763 (n10083, n_6542, n_6543);
  not g13764 (n_6544, n10083);
  and g13765 (n10084, n_4117, n_6544);
  not g13766 (n_6545, n8886);
  not g13767 (n_6546, n10084);
  and g13768 (n10085, n_6545, n_6546);
  not g13769 (n_6547, n8889);
  and g13770 (n10086, n6263, n_6547);
  and g13771 (n10087, n_6542, n10086);
  not g13772 (n_6548, n10085);
  not g13773 (n_6549, n10087);
  and g13774 (n10088, n_6548, n_6549);
  not g13775 (n_6550, n10088);
  and g13776 (n10089, n8887, n_6550);
  not g13777 (n_6551, n10073);
  not g13778 (n_6552, n10089);
  and g13779 (n10090, n_6551, n_6552);
  not g13780 (n_6553, n10090);
  and g13781 (n10091, n8882, n_6553);
  and g13782 (n10092, n_43, n6138);
  not g13783 (n_6554, n10092);
  and g13784 (n10093, n_131, n_6554);
  not g13785 (n_6555, n10093);
  and g13786 (n10094, n_3055, n_6555);
  not g13787 (n_6556, n10094);
  and g13788 (n10095, n_130, n_6556);
  not g13789 (n_6557, n2915);
  and g13790 (n10096, pi0035, n_6557);
  not g13791 (n_6558, n10096);
  and g13792 (n10097, n8938, n_6558);
  not g13793 (n_6559, n10095);
  and g13794 (n10098, n_6559, n10097);
  and g13795 (n10099, n_142, n10098);
  not g13799 (n_6560, n10099);
  not g13800 (n_6561, n10102);
  and g13801 (n10103, n_6560, n_6561);
  and g13802 (n10104, n_144, n_3066);
  not g13803 (n_6562, n10103);
  and g13804 (n10105, n_6562, n10104);
  and g13805 (n10106, n6169, n_6559);
  and g13806 (n10107, n_186, n_3066);
  and g13807 (n10108, n2924, n7479);
  not g13808 (n_6563, n10107);
  and g13809 (n10109, n_4091, n_6563);
  and g13810 (n10110, n10108, n10109);
  and g13811 (n10111, n_4081, n_3209);
  and g13812 (n10112, n7425, n_6563);
  and g13813 (n10113, n10111, n10112);
  not g13814 (n_6564, n10110);
  not g13815 (n_6565, n10113);
  and g13816 (n10114, n_6564, n_6565);
  not g13817 (n_6566, n10106);
  and g13818 (n10115, n_6566, n10114);
  and g13819 (n10116, n2704, n8932);
  not g13820 (n_6567, n10116);
  and g13821 (n10117, n10095, n_6567);
  not g13827 (n_6570, n10098);
  and g13828 (n10121, n_346, n_6570);
  and g13829 (n10122, pi1082, n2518);
  not g13830 (n_6572, n10121);
  and g13831 (n10123, n_6572, n10122);
  not g13838 (n_6576, n8962);
  and g13839 (n10127, pi0038, n_6576);
  not g13845 (n_6579, n10091);
  not g13846 (n_6580, n10130);
  and g13847 (n10131, n_6579, n_6580);
  not g13848 (n_6581, n10131);
  and g13849 (n10132, n2533, n_6581);
  and g13850 (n10133, pi0137, n_5636);
  and g13851 (n10134, n_5661, n10133);
  not g13852 (n_6582, n10134);
  and g13853 (n10135, n_5662, n_6582);
  not g13854 (n_6583, n10135);
  and g13855 (n10136, n8967, n_6583);
  and g13856 (n10137, n8962, n10136);
  not g13857 (n_6584, n10132);
  not g13858 (n_6585, n10137);
  and g13859 (n10138, n_6584, n_6585);
  not g13860 (n_6586, n10138);
  and g13861 (n10139, n_174, n_6586);
  not g13862 (n_6587, n10139);
  and g13863 (n10140, n_167, n_6587);
  not g13869 (n_6590, n10143);
  and g13870 (n10144, n_792, n_6590);
  not g13871 (n_6591, n10070);
  and g13872 (n10145, n_796, n_6591);
  not g13873 (n_6592, n10144);
  and g13874 (po0193, n_6592, n10145);
  and g13875 (n10147, n2717, n2771);
  and g13879 (n10151, n_65, n10150);
  and g13880 (n10152, n_64, n_57);
  and g13881 (n10153, n_60, n2802);
  and g13886 (n10158, n10147, n10157);
  and g13887 (n10159, n_42, n7522);
  not g13888 (n_6593, n10158);
  not g13889 (n_6594, n10159);
  and g13890 (n10160, n_6593, n_6594);
  and g13891 (n10161, n2704, n6479);
  and g13892 (n10162, n6170, n10161);
  and g13893 (n10163, n2532, n_4226);
  and g13894 (n10164, n3373, n10163);
  and g13895 (n10165, n_174, n10164);
  and g13896 (n10166, n10162, n10165);
  and g13897 (n10167, po0740, n10166);
  not g13898 (n_6595, n10160);
  and g13899 (po0194, n_6595, n10167);
  and g13900 (n10169, n_105, n_429);
  and g13901 (n10170, n_87, n_69);
  and g13902 (n10171, n8920, n10170);
  and g13903 (n10172, n_57, n2487);
  and g13904 (n10173, n_85, n2472);
  and g13905 (n10174, n10172, n10173);
  and g13913 (n10182, pi0332, n10181);
  not g13914 (n_6596, n10182);
  and g13915 (n10183, n_103, n_6596);
  and g13916 (n10184, n6479, n9468);
  and g13917 (n10185, n2501, n10184);
  and g13918 (n10186, n2508, n10185);
  not g13925 (n_6598, n10191);
  and g13926 (n10192, n_161, n_6598);
  and g13927 (n10193, n_162, n2519);
  and g13928 (n10194, pi0024, n10193);
  and g13929 (n10195, n2709, n10194);
  not g13930 (n_6599, n10195);
  and g13931 (n10196, pi0038, n_6599);
  and g13932 (n10197, n2571, n_4226);
  not g13933 (n_6600, n10192);
  and g13934 (n10198, n_6600, n10197);
  not g13935 (n_6601, n10196);
  and g13936 (po0196, n_6601, n10198);
  and g13937 (n10200, n_161, n10197);
  not g13938 (n_6603, pi1082);
  and g13939 (n10201, pi0786, n_6603);
  not g13940 (n_6604, pi0984);
  not g13941 (n_6605, n2932);
  and g13942 (n10202, n_6604, n_6605);
  not g13943 (n_6606, n10202);
  and g13944 (n10203, pi0835, n_6606);
  not g13945 (n_6607, n10203);
  and g13946 (n10204, n6183, n_6607);
  not g13947 (n_6608, n10204);
  and g13948 (n10205, n6217, n_6608);
  and g13949 (n10206, pi1093, n10205);
  and g13950 (n10207, n6184, n6380);
  not g13951 (n_6609, n10206);
  and g13952 (n10208, n_6609, n10207);
  and g13953 (n10209, n_223, n10208);
  and g13954 (n10210, n6198, n10205);
  not g13955 (n_6610, n10210);
  and g13956 (n10211, n10207, n_6610);
  and g13957 (n10212, n6205, n10211);
  and g13958 (n10213, n_3140, n10205);
  not g13959 (n_6611, n10213);
  and g13960 (n10214, n10207, n_6611);
  and g13961 (n10215, n_3119, n10214);
  not g13962 (n_6612, n10212);
  and g13963 (n10216, n_234, n_6612);
  not g13964 (n_6613, n10215);
  and g13965 (n10217, n_6613, n10216);
  not g13966 (n_6614, n10209);
  and g13967 (n10218, n_6614, n10217);
  and g13968 (n10219, n_36, n10208);
  and g13969 (n10220, n6242, n10211);
  and g13970 (n10221, n_3162, n10214);
  not g13971 (n_6615, n10220);
  and g13972 (n10222, pi0299, n_6615);
  not g13973 (n_6616, n10221);
  and g13974 (n10223, n_6616, n10222);
  not g13975 (n_6617, n10219);
  and g13976 (n10224, n_6617, n10223);
  not g13977 (n_6618, n10201);
  not g13978 (n_6619, n10218);
  and g13979 (n10225, n_6618, n_6619);
  not g13980 (n_6620, n10224);
  and g13981 (n10226, n_6620, n10225);
  and g13982 (n10227, n5853, n_3164);
  and g13983 (n10228, n3470, n_3122);
  not g13984 (n_6621, n10227);
  not g13985 (n_6622, n10228);
  and g13986 (n10229, n_6621, n_6622);
  not g13991 (n_6624, n10226);
  not g13992 (n_6625, n10232);
  and g13993 (n10233, n_6624, n_6625);
  not g13994 (n_6626, n10233);
  and g13995 (n10234, pi0039, n_6626);
  and g13996 (n10235, n_162, n_144);
  and g13997 (n10236, n6169, n6486);
  not g13998 (n_6628, pi0986);
  and g13999 (n10237, n_6628, n_3209);
  not g14000 (n_6629, n10237);
  and g14001 (n10238, pi0252, n_6629);
  not g14002 (n_6630, n10238);
  and g14003 (n10239, pi0314, n_6630);
  and g14004 (n10240, pi0108, n2714);
  and g14005 (n10241, n2773, n10240);
  and g14006 (n10242, n_3052, n2494);
  and g14007 (n10243, n2720, n10242);
  and g14008 (n10244, n2714, n_360);
  and g14009 (n10245, n8921, n9076);
  and g14010 (n10246, n_56, n_65);
  and g14011 (n10247, n10245, n10246);
  not g14024 (n_6631, n10241);
  and g14025 (n10260, n_108, n_6631);
  not g14026 (n_6632, n10259);
  and g14027 (n10261, n_6632, n10260);
  and g14028 (n10262, n6151, n10239);
  not g14029 (n_6633, n10261);
  and g14030 (n10263, n_6633, n10262);
  and g14031 (n10264, n_108, n_3052);
  and g14032 (n10265, n10256, n10264);
  not g14033 (n_6634, n2760);
  not g14034 (n_6635, n10265);
  and g14035 (n10266, n_6634, n_6635);
  not g14041 (n_6638, n10263);
  not g14042 (n_6639, n10269);
  and g14043 (n10270, n_6638, n_6639);
  not g14044 (n_6640, n10270);
  and g14045 (n10271, n2704, n_6640);
  not g14046 (n_6641, n10271);
  and g14047 (n10272, n_130, n_6641);
  not g14048 (n_6642, n6483);
  and g14049 (n10273, pi0035, n_6642);
  not g14050 (n_6643, n10273);
  and g14051 (n10274, n2508, n_6643);
  and g14052 (n10275, n2510, n10274);
  not g14053 (n_6644, n10272);
  and g14054 (n10276, n_6644, n10275);
  not g14055 (n_6645, n10236);
  not g14056 (n_6646, n10276);
  and g14057 (n10277, n_6645, n_6646);
  not g14058 (n_6647, n10277);
  and g14059 (n10278, n10235, n_6647);
  not g14060 (n_6648, n10234);
  not g14061 (n_6649, n10278);
  and g14062 (n10279, n_6648, n_6649);
  not g14063 (n_6650, n10279);
  and g14064 (po0197, n10200, n_6650);
  and g14071 (n10287, n6479, n10286);
  not g14072 (n_6651, n10287);
  and g14073 (n10288, pi1082, n_6651);
  and g14074 (n10289, n2518, n_874);
  not g14075 (n_6652, n10286);
  and g14076 (n10290, n_143, n_6652);
  not g14077 (n_6653, n10290);
  and g14078 (n10291, n10289, n_6653);
  not g14079 (n_6654, n10291);
  and g14080 (n10292, n_6603, n_6654);
  not g14081 (n_6655, n10288);
  and g14082 (n10293, n10165, n_6655);
  not g14083 (n_6656, n10292);
  and g14084 (po0198, n_6656, n10293);
  and g14085 (n10295, n_301, n6197);
  and g14086 (n10296, pi0144, n10295);
  and g14087 (n10297, n_299, n10296);
  not g14088 (n_6657, n10297);
  and g14089 (n10298, n_234, n_6657);
  and g14090 (n10299, n_266, n6197);
  and g14091 (n10300, pi0161, n10299);
  and g14092 (n10301, n_263, n10300);
  not g14093 (n_6658, n10301);
  and g14094 (n10302, n_4115, n_6658);
  not g14095 (n_6659, n10298);
  and g14096 (n10303, pi0232, n_6659);
  not g14097 (n_6660, n10302);
  and g14098 (n10304, n_6660, n10303);
  not g14099 (n_6661, n10304);
  and g14100 (n10305, n_134, n_6661);
  not g14101 (n_6662, n10305);
  and g14102 (n10306, pi0039, n_6662);
  and g14103 (n10307, n_3181, n_134);
  not g14104 (n_6663, n10307);
  and g14105 (n10308, n_162, n_6663);
  not g14106 (n_6664, n10306);
  not g14107 (n_6665, n10308);
  and g14108 (n10309, n_6664, n_6665);
  not g14109 (n_6666, n2620);
  and g14110 (n10310, n_6666, n10309);
  and g14111 (n10311, n_4137, n_6663);
  and g14112 (n10312, n_538, n10307);
  not g14113 (n_6667, n10312);
  and g14114 (n10313, n7506, n_6667);
  and g14115 (n10314, n_3181, pi0072);
  not g14116 (n_6668, n10314);
  and g14117 (n10315, n2924, n_6668);
  not g14118 (n_6669, pi0044);
  and g14119 (n10316, n_6669, n2521);
  and g14120 (n10317, n_3184, n10316);
  and g14121 (n10318, n7479, n10317);
  and g14122 (n10319, n7477, n10318);
  not g14123 (n_6670, n10319);
  and g14124 (n10320, pi0041, n_6670);
  and g14125 (n10321, n_3182, n6272);
  and g14126 (n10322, n_134, pi0101);
  not g14127 (n_6671, n10322);
  and g14128 (n10323, n_3181, n_6671);
  and g14129 (n10324, pi0252, n6479);
  and g14130 (n10325, n_4119, n2709);
  and g14131 (n10326, n7479, n10324);
  and g14132 (n10327, n10325, n10326);
  and g14133 (n10328, n_6669, n10327);
  and g14134 (n10329, n10323, n10328);
  not g14135 (n_6672, n10321);
  and g14136 (n10330, n_6672, n10329);
  not g14137 (n_6673, n10330);
  and g14138 (n10331, n10315, n_6673);
  not g14139 (n_6674, n10320);
  and g14140 (n10332, n_6674, n10331);
  not g14141 (n_6675, n10332);
  and g14142 (n10333, n10313, n_6675);
  not g14143 (n_6676, n10311);
  not g14144 (n_6677, n10333);
  and g14145 (n10334, n_6676, n_6677);
  not g14146 (n_6678, n10334);
  and g14147 (n10335, n_162, n_6678);
  and g14148 (n10336, n2620, n_6664);
  not g14149 (n_6679, n10335);
  and g14150 (n10337, n_6679, n10336);
  not g14151 (n_6680, n10310);
  and g14152 (n10338, pi0075, n_6680);
  not g14153 (n_6681, n10337);
  and g14154 (n10339, n_6681, n10338);
  and g14155 (n10340, n_958, n10308);
  and g14156 (n10341, n_188, n10307);
  and g14157 (n10342, n2709, n6479);
  and g14158 (n10343, n_6669, n10342);
  and g14159 (n10344, n10323, n10343);
  not g14160 (n_6682, n10344);
  and g14161 (n10345, n_6668, n_6682);
  not g14162 (n_6683, n10317);
  and g14163 (n10346, pi0041, n_6683);
  and g14164 (n10347, pi0228, n10345);
  not g14165 (n_6684, n10346);
  and g14166 (n10348, n_6684, n10347);
  not g14167 (n_6685, n10341);
  and g14168 (n10349, n2625, n_6685);
  not g14169 (n_6686, n10348);
  and g14170 (n10350, n_6686, n10349);
  not g14176 (n_6689, n10309);
  and g14177 (n10354, pi0038, n_6689);
  not g14178 (n_6690, n10318);
  and g14179 (n10355, pi0041, n_6690);
  and g14180 (n10356, n2924, n_6672);
  not g14181 (n_6691, n10315);
  not g14182 (n_6692, n10356);
  and g14183 (n10357, n_6691, n_6692);
  not g14184 (n_6693, n7479);
  and g14185 (n10358, n_134, n_6693);
  not g14186 (n_6694, n10345);
  not g14187 (n_6695, n10358);
  and g14188 (n10359, n_6694, n_6695);
  and g14189 (n10360, n_6672, n10359);
  not g14190 (n_6696, n10355);
  not g14191 (n_6697, n10357);
  and g14192 (n10361, n_6696, n_6697);
  not g14193 (n_6698, n10360);
  and g14194 (n10362, n_6698, n10361);
  not g14195 (n_6699, n10362);
  and g14196 (n10363, n10313, n_6699);
  not g14197 (n_6700, n10363);
  and g14198 (n10364, n_6676, n_6700);
  not g14199 (n_6701, n10364);
  and g14200 (n10365, n_162, n_6701);
  not g14201 (n_6702, n10365);
  and g14202 (n10366, n_6664, n_6702);
  not g14203 (n_6703, n10366);
  and g14204 (n10367, n6285, n_6703);
  and g14205 (n10368, pi0287, n2521);
  and g14206 (n10369, n10304, n10368);
  not g14207 (n_6704, n10369);
  and g14208 (n10370, n_6662, n_6704);
  not g14209 (n_6705, n10370);
  and g14210 (n10371, pi0039, n_6705);
  not g14211 (n_6708, pi0959);
  and g14212 (n10372, pi0901, n_6708);
  not g14213 (n_6710, pi0480);
  and g14214 (n10373, n_6710, pi0949);
  and g14215 (n10374, n2717, n2780);
  and g14216 (n10375, n2708, n10374);
  not g14217 (n_6712, n10373);
  and g14218 (n10376, n_6712, n10375);
  and g14219 (n10377, n2708, n10373);
  and g14220 (n10378, n2700, n_357);
  and g14221 (n10379, n_112, n6451);
  and g14222 (n10380, n2780, n10379);
  not g14223 (n_6713, n10380);
  and g14224 (n10381, n_113, n_6713);
  not g14229 (n_6715, n10376);
  and g14230 (n10385, n10372, n_6715);
  not g14231 (n_6716, n10384);
  and g14232 (n10386, n_6716, n10385);
  and g14233 (n10387, n2701, n2758);
  and g14234 (n10388, pi0110, n10387);
  and g14235 (n10389, n10377, n10388);
  not g14236 (n_6717, n10372);
  not g14237 (n_6718, n10389);
  and g14238 (n10390, n_6717, n_6718);
  and g14239 (n10391, n_3208, pi0252);
  and g14245 (n10395, n_134, n10394);
  and g14246 (n10396, n10162, n10388);
  not g14247 (n_6721, n10391);
  and g14248 (n10397, n10373, n_6721);
  and g14249 (n10398, n10396, n10397);
  not g14250 (n_6722, n10395);
  not g14251 (n_6723, n10398);
  and g14252 (n10399, n_6722, n_6723);
  not g14253 (n_6724, n10399);
  and g14254 (n10400, n_6669, n_6724);
  and g14255 (n10401, n_3184, n10400);
  not g14256 (n_6725, n10401);
  and g14257 (n10402, pi0041, n_6725);
  and g14258 (n10403, pi0044, pi0072);
  and g14259 (n10404, n6479, n_6721);
  and g14260 (n10405, n10389, n10404);
  not g14261 (n_6726, n10405);
  and g14262 (n10406, n_134, n_6726);
  not g14263 (n_6727, n10394);
  and g14264 (n10407, n_6727, n10406);
  not g14265 (n_6728, n10407);
  and g14266 (n10408, n_6669, n_6728);
  not g14267 (n_6729, n10403);
  not g14268 (n_6730, n10408);
  and g14269 (n10409, n_6729, n_6730);
  and g14270 (n10410, n_3184, n10409);
  not g14271 (n_6731, n10410);
  and g14272 (n10411, n10323, n_6731);
  not g14273 (n_6732, n10402);
  not g14274 (n_6733, n10411);
  and g14275 (n10412, n_6732, n_6733);
  not g14276 (n_6734, n10412);
  and g14277 (n10413, n_188, n_6734);
  not g14278 (n_6735, n7451);
  and g14279 (n10414, n_134, n_6735);
  not g14280 (n_6736, n7457);
  and g14281 (n10415, n_6736, n10414);
  and g14282 (n10416, n6479, n_4103);
  and g14283 (n10417, n_4104, n10416);
  and g14284 (n10418, n_134, n7457);
  not g14285 (n_6737, n10417);
  and g14286 (n10419, n_6737, n10418);
  not g14287 (n_6738, n10415);
  and g14288 (n10420, n_3206, n_6738);
  not g14289 (n_6739, n10419);
  and g14290 (n10421, n_6739, n10420);
  not g14291 (n_6740, n10421);
  and g14292 (n10422, n10414, n_6740);
  not g14293 (n_6741, n10422);
  and g14294 (n10423, n_6669, n_6741);
  not g14295 (n_6742, n10423);
  and g14296 (n10424, n_6729, n_6742);
  and g14297 (n10425, n_3184, n10424);
  not g14298 (n_6743, n10425);
  and g14299 (n10426, n10323, n_6743);
  and g14300 (n10427, n7451, n_6736);
  and g14301 (n10428, n_3206, n_4106);
  not g14302 (n_6744, n10427);
  and g14303 (n10429, n_6744, n10428);
  not g14304 (n_6745, n10429);
  and g14305 (n10430, n_6669, n_6745);
  and g14306 (n10431, pi1093, n_6735);
  not g14307 (n_6746, n10431);
  and g14308 (n10432, n10430, n_6746);
  and g14309 (n10433, n_3184, n10432);
  not g14310 (n_6747, n10433);
  and g14311 (n10434, pi0041, n_6747);
  not g14312 (n_6748, n10434);
  and g14313 (n10435, n_538, n_6748);
  not g14314 (n_6749, n10426);
  and g14315 (n10436, n_6749, n10435);
  and g14316 (n10437, n2935, n_4097);
  and g14317 (n10438, n2937, n10437);
  not g14318 (n_6750, n10438);
  and g14319 (n10439, n_4146, n_6750);
  not g14320 (n_6751, n10439);
  and g14321 (n10440, n2461, n_6751);
  not g14322 (n_6752, n10440);
  and g14323 (n10441, n7434, n_6752);
  not g14324 (n_6753, n10441);
  and g14325 (n10442, n7431, n_6753);
  not g14326 (n_6754, n10442);
  and g14327 (n10443, n_138, n_6754);
  not g14328 (n_6755, n10443);
  and g14329 (n10444, n_350, n_6755);
  not g14330 (n_6756, n10444);
  and g14331 (n10445, n_135, n_6756);
  and g14332 (n10446, n10416, n10418);
  not g14333 (n_6757, n10445);
  and g14334 (n10447, n_6757, n10446);
  not g14335 (n_6758, n10447);
  and g14336 (n10448, n_6744, n_6758);
  and g14337 (n10449, pi1093, n10448);
  not g14338 (n_6759, n10449);
  and g14339 (n10450, n10430, n_6759);
  and g14340 (n10451, n_3184, n10450);
  not g14341 (n_6760, n10451);
  and g14342 (n10452, pi0041, n_6760);
  and g14343 (n10453, n_134, n10448);
  not g14344 (n_6761, n10453);
  and g14345 (n10454, pi1093, n_6761);
  not g14346 (n_6762, n10454);
  and g14347 (n10455, n_6740, n_6762);
  not g14348 (n_6763, n10455);
  and g14349 (n10456, n_6669, n_6763);
  not g14350 (n_6764, n10456);
  and g14351 (n10457, n_6729, n_6764);
  and g14352 (n10458, n_3184, n10457);
  not g14353 (n_6765, n10458);
  and g14354 (n10459, n10323, n_6765);
  not g14355 (n_6766, n10459);
  and g14356 (n10460, n2924, n_6766);
  not g14357 (n_6767, n10452);
  and g14358 (n10461, n_6767, n10460);
  not g14359 (n_6768, n10436);
  and g14360 (n10462, pi0228, n_6768);
  not g14361 (n_6769, n10461);
  and g14362 (n10463, n_6769, n10462);
  not g14363 (n_6770, n10413);
  and g14364 (n10464, n_162, n_6770);
  not g14365 (n_6771, n10463);
  and g14366 (n10465, n_6771, n10464);
  not g14367 (n_6772, n10371);
  and g14368 (n10466, n2608, n_6772);
  not g14369 (n_6773, n10465);
  and g14370 (n10467, n_6773, n10466);
  not g14377 (n_6777, n10353);
  and g14378 (n10471, n_171, n_6777);
  not g14379 (n_6778, n10470);
  and g14380 (n10472, n_6778, n10471);
  not g14381 (n_6779, n10339);
  not g14382 (n_6780, n10472);
  and g14383 (n10473, n_6779, n_6780);
  not g14384 (n_6781, n10473);
  and g14385 (n10474, n7429, n_6781);
  and g14386 (n10475, n_4196, n_6689);
  not g14387 (n_6782, n10475);
  and g14388 (n10476, n_4226, n_6782);
  not g14389 (n_6783, n10474);
  and g14390 (n10477, n_6783, n10476);
  and g14391 (n10478, pi0039, pi0232);
  and g14392 (n10479, n10301, n10478);
  not g14397 (n_6785, n10477);
  not g14398 (n_6786, n10482);
  and g14399 (po0199, n_6785, n_6786);
  and g14400 (n10484, pi0211, pi0214);
  and g14401 (n10485, pi0212, n10484);
  not g14402 (n_6791, pi0219);
  not g14403 (n_6792, n10485);
  and g14404 (n10486, n_6791, n_6792);
  and g14405 (n10487, pi0207, pi0208);
  and g14406 (n10488, pi0042, n_134);
  and g14407 (n10489, n_6666, n10488);
  not g14408 (n_6795, n10488);
  and g14409 (n10490, n_4137, n_6795);
  and g14410 (n10491, n_3198, n2924);
  not g14411 (n_6796, n10491);
  and g14412 (n10492, n10488, n_6796);
  not g14413 (n_6797, n10492);
  and g14414 (n10493, n7506, n_6797);
  and g14415 (n10494, pi0114, n_6795);
  not g14416 (n_6798, n10494);
  and g14417 (n10495, n10491, n_6798);
  and g14418 (n10496, n6266, n10328);
  and g14419 (n10497, n_3193, n10496);
  and g14420 (n10498, n_3194, n10497);
  not g14421 (n_6799, n10498);
  and g14422 (n10499, n10488, n_6799);
  and g14423 (n10500, n6265, n10317);
  and g14424 (n10501, n6269, n10500);
  and g14425 (n10502, n7479, n10501);
  not g14426 (n_6800, n6268);
  and g14427 (n10503, n_3197, n_6800);
  and g14428 (n10504, n10502, n10503);
  and g14429 (n10505, n7477, n10504);
  and g14430 (n10506, n_3187, n10505);
  not g14431 (n_6801, n10499);
  and g14432 (n10507, n_3197, n_6801);
  not g14433 (n_6802, n10506);
  and g14434 (n10508, n_6802, n10507);
  not g14435 (n_6803, n10508);
  and g14436 (n10509, n10495, n_6803);
  not g14437 (n_6804, n10509);
  and g14438 (n10510, n10493, n_6804);
  not g14439 (n_6805, n10490);
  and g14440 (n10511, n2620, n_6805);
  not g14441 (n_6806, n10510);
  and g14442 (n10512, n_6806, n10511);
  not g14443 (n_6807, n10489);
  and g14444 (n10513, n_162, n_6807);
  not g14445 (n_6808, n10512);
  and g14446 (n10514, n_6808, n10513);
  and g14447 (n10515, n_134, pi0199);
  not g14448 (n_6810, n10515);
  and g14449 (n10516, n_3410, n_6810);
  not g14450 (n_6811, n10516);
  and g14451 (n10517, n_234, n_6811);
  not g14452 (n_6812, n10295);
  and g14453 (n10518, n_134, n_6812);
  and g14454 (n10519, pi0199, n10518);
  not g14455 (n_6813, n10519);
  and g14456 (n10520, pi0232, n_6813);
  not g14457 (n_6814, n10520);
  and g14458 (n10521, n10517, n_6814);
  and g14459 (n10522, n_266, n7473);
  not g14460 (n_6815, n10522);
  and g14461 (n10523, n_134, n_6815);
  and g14462 (n10524, pi0299, n10523);
  not g14463 (n_6816, n10524);
  and g14464 (n10525, pi0039, n_6816);
  not g14465 (n_6817, n10521);
  and g14466 (n10526, n_6817, n10525);
  not g14467 (n_6818, n10514);
  not g14468 (n_6819, n10526);
  and g14469 (n10527, n_6818, n_6819);
  not g14470 (n_6820, n10527);
  and g14471 (n10528, pi0075, n_6820);
  and g14472 (n10529, n_162, n_6795);
  and g14473 (n10530, n_958, n10529);
  and g14474 (n10531, n6266, n10343);
  and g14475 (n10532, pi0228, n10531);
  and g14476 (n10533, n6271, n10532);
  not g14477 (n_6821, n10533);
  and g14478 (n10534, n10488, n_6821);
  and g14479 (n10535, pi0228, n10501);
  and g14480 (n10536, n_3198, n10535);
  and g14481 (n10537, n_3197, n10536);
  and g14482 (n10538, n_3187, n10537);
  not g14483 (n_6822, n10534);
  and g14484 (n10539, n2625, n_6822);
  not g14485 (n_6823, n10538);
  and g14486 (n10540, n_6823, n10539);
  not g14487 (n_6824, n10530);
  and g14488 (n10541, pi0087, n_6824);
  not g14489 (n_6825, n10540);
  and g14490 (n10542, n_6825, n10541);
  and g14491 (n10543, n_6819, n10542);
  and g14492 (n10544, pi0115, n_6795);
  and g14493 (n10545, pi0042, n_3197);
  and g14494 (n10546, pi0072, pi0116);
  and g14495 (n10547, pi0072, pi0113);
  not g14496 (n_6826, n6265);
  and g14497 (n10548, pi0072, n_6826);
  and g14498 (n10549, n_3182, n10411);
  not g14499 (n_6827, n10548);
  not g14500 (n_6828, n10549);
  and g14501 (n10550, n_6827, n_6828);
  not g14502 (n_6829, n10550);
  and g14503 (n10551, n_3193, n_6829);
  not g14504 (n_6830, n10547);
  not g14505 (n_6831, n10551);
  and g14506 (n10552, n_6830, n_6831);
  not g14507 (n_6832, n10552);
  and g14508 (n10553, n_3194, n_6832);
  not g14509 (n_6833, n10546);
  not g14510 (n_6834, n10553);
  and g14511 (n10554, n_6833, n_6834);
  not g14512 (n_6835, n10554);
  and g14513 (n10555, n10545, n_6835);
  and g14514 (n10556, n6265, n10401);
  and g14515 (n10557, n_3193, n10556);
  and g14516 (n10558, n_3194, n10557);
  not g14517 (n_6836, n10558);
  and g14518 (n10559, n_3187, n_6836);
  not g14519 (n_6837, n10559);
  and g14520 (n10560, n_6798, n_6837);
  not g14521 (n_6838, n10555);
  and g14522 (n10561, n_6838, n10560);
  not g14523 (n_6839, n10561);
  and g14524 (n10562, n_3198, n_6839);
  not g14525 (n_6840, n10544);
  and g14526 (n10563, n_188, n_6840);
  not g14527 (n_6841, n10562);
  and g14528 (n10564, n_6841, n10563);
  and g14529 (n10565, n_3182, n10459);
  not g14530 (n_6842, n10565);
  and g14531 (n10566, n_6827, n_6842);
  not g14532 (n_6843, n10566);
  and g14533 (n10567, n_3193, n_6843);
  not g14534 (n_6844, n10567);
  and g14535 (n10568, n_6830, n_6844);
  not g14536 (n_6845, n10568);
  and g14537 (n10569, n_3194, n_6845);
  not g14538 (n_6846, n10569);
  and g14539 (n10570, n_6833, n_6846);
  not g14540 (n_6847, n10570);
  and g14541 (n10571, n10545, n_6847);
  and g14542 (n10572, n6265, n10451);
  and g14543 (n10573, n6269, n10572);
  not g14544 (n_6848, n10573);
  and g14545 (n10574, n_3187, n_6848);
  not g14546 (n_6849, n10574);
  and g14547 (n10575, n_6798, n_6849);
  not g14548 (n_6850, n10571);
  and g14549 (n10576, n_6850, n10575);
  not g14550 (n_6851, n10576);
  and g14551 (n10577, n10491, n_6851);
  and g14552 (n10578, n_3198, n_538);
  and g14553 (n10579, n6265, n10433);
  and g14554 (n10580, n6269, n10579);
  and g14555 (n10581, n_3187, n10580);
  and g14556 (n10582, n_3182, n10426);
  not g14557 (n_6852, n10582);
  and g14558 (n10583, n_6827, n_6852);
  not g14559 (n_6853, n10583);
  and g14560 (n10584, n_3193, n_6853);
  not g14561 (n_6854, n10584);
  and g14562 (n10585, n_6830, n_6854);
  not g14563 (n_6855, n10585);
  and g14564 (n10586, n_3194, n_6855);
  not g14565 (n_6856, n10586);
  and g14566 (n10587, n_6833, n_6856);
  and g14567 (n10588, pi0042, n10587);
  not g14568 (n_6857, n10581);
  and g14569 (n10589, n_3197, n_6857);
  not g14570 (n_6858, n10588);
  and g14571 (n10590, n_6858, n10589);
  not g14572 (n_6859, n10590);
  and g14573 (n10591, n_6798, n_6859);
  not g14574 (n_6860, n10591);
  and g14575 (n10592, n10578, n_6860);
  not g14581 (n_6863, n10564);
  and g14582 (n10596, n_162, n_6863);
  not g14583 (n_6864, n10595);
  and g14584 (n10597, n_6864, n10596);
  and g14585 (n10598, pi0232, pi0299);
  and g14586 (n10599, n10299, n10368);
  not g14587 (n_6865, n10523);
  and g14588 (n10600, n_6865, n10598);
  not g14589 (n_6866, n10599);
  and g14590 (n10601, n_6866, n10600);
  and g14591 (n10602, pi0232, n_234);
  and g14592 (n10603, n6197, n10368);
  and g14593 (n10604, n_301, n10603);
  not g14594 (n_6867, n10518);
  not g14595 (n_6868, n10604);
  and g14596 (n10605, n_6867, n_6868);
  not g14597 (n_6869, n10605);
  and g14598 (n10606, pi0199, n_6869);
  not g14599 (n_6870, n10606);
  and g14600 (n10607, n10602, n_6870);
  and g14601 (n10608, pi0072, n_3410);
  not g14602 (n_6871, n10608);
  and g14603 (n10609, pi0299, n_6871);
  not g14604 (n_6872, n10609);
  and g14605 (n10610, n10516, n_6872);
  not g14606 (n_6873, n10601);
  not g14607 (n_6874, n10610);
  and g14608 (n10611, n_6873, n_6874);
  not g14609 (n_6875, n10607);
  and g14610 (n10612, n_6875, n10611);
  not g14611 (n_6876, n10612);
  and g14612 (n10613, pi0039, n_6876);
  not g14613 (n_6877, n10597);
  not g14614 (n_6878, n10613);
  and g14615 (n10614, n_6877, n_6878);
  not g14616 (n_6879, n10614);
  and g14617 (n10615, n2608, n_6879);
  and g14618 (n10616, n6269, n10531);
  not g14619 (n_6880, n10616);
  and g14620 (n10617, n_134, n_6880);
  not g14621 (n_6881, n10617);
  and g14622 (n10618, n_6695, n_6881);
  not g14623 (n_6882, n10618);
  and g14624 (n10619, pi0042, n_6882);
  and g14625 (n10620, n_3187, n10504);
  not g14626 (n_6883, n10619);
  and g14627 (n10621, n_3197, n_6883);
  not g14628 (n_6884, n10620);
  and g14629 (n10622, n_6884, n10621);
  not g14630 (n_6885, n10622);
  and g14631 (n10623, n10495, n_6885);
  not g14632 (n_6886, n10623);
  and g14633 (n10624, n10493, n_6886);
  not g14634 (n_6887, n10624);
  and g14635 (n10625, n_6805, n_6887);
  not g14636 (n_6888, n10625);
  and g14637 (n10626, n_162, n_6888);
  not g14638 (n_6889, n10626);
  and g14639 (n10627, n_6819, n_6889);
  not g14640 (n_6890, n10627);
  and g14641 (n10628, n6285, n_6890);
  not g14642 (n_6891, n10529);
  and g14643 (n10629, n_6819, n_6891);
  not g14644 (n_6892, n10629);
  and g14645 (n10630, pi0038, n_6892);
  not g14646 (n_6893, n10630);
  and g14647 (n10631, n_172, n_6893);
  not g14648 (n_6894, n10628);
  and g14649 (n10632, n_6894, n10631);
  not g14650 (n_6895, n10615);
  and g14651 (n10633, n_6895, n10632);
  not g14652 (n_6896, n10543);
  and g14653 (n10634, n_171, n_6896);
  not g14654 (n_6897, n10633);
  and g14655 (n10635, n_6897, n10634);
  not g14656 (n_6898, n10528);
  and g14657 (n10636, n7429, n_6898);
  not g14658 (n_6899, n10635);
  and g14659 (n10637, n_6899, n10636);
  not g14660 (n_6900, n10487);
  not g14661 (n_6901, n10637);
  and g14662 (n10638, n_6900, n_6901);
  and g14663 (n10639, n_134, pi0200);
  not g14664 (n_6903, n10639);
  and g14665 (n10640, n_3410, n_6903);
  not g14666 (n_6904, n10640);
  and g14667 (n10641, n_234, n_6904);
  and g14668 (n10642, pi0200, n10518);
  not g14669 (n_6905, n10642);
  and g14670 (n10643, pi0232, n_6905);
  not g14671 (n_6906, n10643);
  and g14672 (n10644, n10641, n_6906);
  not g14673 (n_6907, n10644);
  and g14674 (n10645, pi0039, n_6907);
  and g14675 (n10646, n_6817, n10645);
  not g14676 (n_6908, n10646);
  and g14677 (n10647, n_6891, n_6908);
  and g14678 (n10648, n_4196, n10647);
  not g14679 (n_6909, n10648);
  and g14680 (n10649, n10487, n_6909);
  and g14681 (n10650, n10526, n10645);
  not g14682 (n_6910, n10650);
  and g14683 (n10651, n_6818, n_6910);
  not g14684 (n_6911, n10651);
  and g14685 (n10652, pi0075, n_6911);
  and g14686 (n10653, n_6889, n_6910);
  not g14687 (n_6912, n10653);
  and g14688 (n10654, n6285, n_6912);
  not g14689 (n_6913, n10647);
  and g14690 (n10655, pi0038, n_6913);
  not g14691 (n_6914, n10655);
  and g14692 (n10656, n_172, n_6914);
  not g14693 (n_6915, n10631);
  not g14694 (n_6916, n10656);
  and g14695 (n10657, n_6915, n_6916);
  and g14696 (n10658, pi0232, n_6870);
  and g14697 (n10659, pi0200, n_6869);
  not g14698 (n_6917, n10659);
  and g14699 (n10660, n10658, n_6917);
  and g14700 (n10661, n_234, n10660);
  and g14701 (n10662, n10610, n_6903);
  not g14702 (n_6918, n10662);
  and g14703 (n10663, n_6873, n_6918);
  not g14704 (n_6919, n10661);
  and g14705 (n10664, n_6919, n10663);
  not g14706 (n_6920, n10664);
  and g14707 (n10665, pi0039, n_6920);
  not g14708 (n_6921, n10665);
  and g14709 (n10666, n_6877, n_6921);
  not g14710 (n_6922, n10666);
  and g14711 (n10667, n2608, n_6922);
  not g14712 (n_6923, n10654);
  not g14713 (n_6924, n10657);
  and g14714 (n10668, n_6923, n_6924);
  not g14715 (n_6925, n10667);
  and g14716 (n10669, n_6925, n10668);
  and g14717 (n10670, n10541, n_6910);
  and g14718 (n10671, n_6825, n10670);
  not g14719 (n_6926, n10671);
  and g14720 (n10672, n_171, n_6926);
  not g14721 (n_6927, n10669);
  and g14722 (n10673, n_6927, n10672);
  not g14723 (n_6928, n10652);
  and g14724 (n10674, n7429, n_6928);
  not g14725 (n_6929, n10673);
  and g14726 (n10675, n_6929, n10674);
  not g14727 (n_6930, n10675);
  and g14728 (n10676, n10649, n_6930);
  not g14729 (n_6931, n10638);
  not g14730 (n_6932, n10676);
  and g14731 (n10677, n_6931, n_6932);
  and g14732 (n10678, n_4196, n10629);
  not g14733 (n_6933, n10486);
  not g14734 (n_6934, n10678);
  and g14735 (n10679, n_6933, n_6934);
  not g14736 (n_6935, n10677);
  and g14737 (n10680, n_6935, n10679);
  and g14738 (n10681, pi0039, n_6817);
  not g14739 (n_6936, n10681);
  and g14740 (n10682, n_6818, n_6936);
  not g14741 (n_6937, n10682);
  and g14742 (n10683, pi0075, n_6937);
  and g14743 (n10684, n10542, n_6936);
  and g14744 (n10685, n_6889, n_6936);
  not g14745 (n_6938, n10685);
  and g14746 (n10686, n6285, n_6938);
  and g14747 (n10687, n_6891, n_6936);
  not g14748 (n_6939, n10687);
  and g14749 (n10688, pi0038, n_6939);
  not g14750 (n_6940, n10658);
  and g14751 (n10689, n10517, n_6940);
  not g14752 (n_6941, n10689);
  and g14753 (n10690, pi0039, n_6941);
  not g14754 (n_6942, n10690);
  and g14755 (n10691, n_6877, n_6942);
  not g14756 (n_6943, n10691);
  and g14757 (n10692, n2608, n_6943);
  not g14764 (n_6947, n10684);
  and g14765 (n10696, n_171, n_6947);
  not g14766 (n_6948, n10695);
  and g14767 (n10697, n_6948, n10696);
  not g14768 (n_6949, n10683);
  and g14769 (n10698, n7429, n_6949);
  not g14770 (n_6950, n10697);
  and g14771 (n10699, n_6950, n10698);
  and g14772 (n10700, n_4196, n10687);
  not g14773 (n_6951, n10700);
  and g14774 (n10701, n_6900, n_6951);
  not g14775 (n_6952, n10699);
  and g14776 (n10702, n_6952, n10701);
  and g14777 (n10703, n_6818, n_6908);
  not g14778 (n_6953, n10703);
  and g14779 (n10704, pi0075, n_6953);
  and g14780 (n10705, n10542, n_6908);
  not g14781 (n_6954, n10517);
  not g14782 (n_6955, n10641);
  and g14783 (n10706, n_6954, n_6955);
  not g14784 (n_6956, n10660);
  not g14785 (n_6957, n10706);
  and g14786 (n10707, n_6956, n_6957);
  not g14787 (n_6958, n10707);
  and g14788 (n10708, pi0039, n_6958);
  not g14789 (n_6959, n10708);
  and g14790 (n10709, n_6877, n_6959);
  not g14791 (n_6960, n10709);
  and g14792 (n10710, n2608, n_6960);
  and g14793 (n10711, n_6889, n_6908);
  not g14794 (n_6961, n10711);
  and g14795 (n10712, n6285, n_6961);
  not g14796 (n_6962, n10712);
  and g14797 (n10713, n10656, n_6962);
  not g14798 (n_6963, n10710);
  and g14799 (n10714, n_6963, n10713);
  not g14800 (n_6964, n10705);
  and g14801 (n10715, n_171, n_6964);
  not g14802 (n_6965, n10714);
  and g14803 (n10716, n_6965, n10715);
  not g14804 (n_6966, n10704);
  and g14805 (n10717, n7429, n_6966);
  not g14806 (n_6967, n10716);
  and g14807 (n10718, n_6967, n10717);
  not g14808 (n_6968, n10718);
  and g14809 (n10719, n10649, n_6968);
  not g14810 (n_6969, n10702);
  not g14811 (n_6970, n10719);
  and g14812 (n10720, n_6969, n_6970);
  not g14813 (n_6971, n10720);
  and g14814 (n10721, n10486, n_6971);
  not g14815 (n_6972, n10680);
  and g14816 (n10722, n_4226, n_6972);
  not g14817 (n_6973, n10721);
  and g14818 (n10723, n_6973, n10722);
  and g14819 (n10724, n_6933, n10523);
  not g14820 (n_6974, n10724);
  and g14821 (n10725, pi0039, n_6974);
  and g14822 (n10726, po1038, n_6891);
  not g14823 (n_6975, n10725);
  and g14824 (n10727, n_6975, n10726);
  or g14825 (po0200, n10723, n10727);
  and g14826 (n10729, pi0043, n_134);
  not g14827 (n_6976, n10729);
  and g14828 (n10730, n_4137, n_6976);
  and g14829 (n10731, n_3187, n6270);
  and g14830 (n10732, n2924, n10731);
  not g14831 (n_6977, n10732);
  and g14832 (n10733, n10729, n_6977);
  not g14833 (n_6978, n10733);
  and g14834 (n10734, n7506, n_6978);
  and g14835 (n10735, n_134, n_6799);
  and g14836 (n10736, pi0043, n10735);
  and g14837 (n10737, n_3188, pi0052);
  and g14838 (n10738, n7477, n10502);
  and g14839 (n10739, n10737, n10738);
  not g14840 (n_6979, n10736);
  not g14841 (n_6980, n10739);
  and g14842 (n10740, n_6979, n_6980);
  not g14843 (n_6981, n10740);
  and g14844 (n10741, n10732, n_6981);
  not g14845 (n_6982, n10741);
  and g14846 (n10742, n10734, n_6982);
  not g14847 (n_6983, n10730);
  not g14848 (n_6984, n10742);
  and g14849 (n10743, n_6983, n_6984);
  not g14850 (n_6985, n10743);
  and g14851 (n10744, n_162, n_6985);
  not g14852 (n_6986, n10744);
  and g14853 (n10745, n2620, n_6986);
  and g14854 (n10746, n_162, n_6976);
  not g14855 (n_6987, n10746);
  and g14856 (n10747, n_6666, n_6987);
  not g14857 (n_6988, n10745);
  not g14858 (n_6989, n10747);
  and g14859 (n10748, n_6988, n_6989);
  not g14860 (n_6990, n10645);
  not g14861 (n_6991, n10748);
  and g14862 (n10749, n_6990, n_6991);
  not g14863 (n_6992, n10749);
  and g14864 (n10750, pi0075, n_6992);
  and g14865 (n10751, n_958, n10746);
  not g14866 (n_6993, n10501);
  and g14867 (n10752, n_3188, n_6993);
  and g14868 (n10753, pi0043, n_6881);
  and g14869 (n10754, pi0228, n10731);
  not g14870 (n_6994, n10753);
  and g14871 (n10755, n_6994, n10754);
  not g14872 (n_6995, n10752);
  and g14873 (n10756, n_6995, n10755);
  not g14874 (n_6996, n10754);
  and g14875 (n10757, n10729, n_6996);
  not g14876 (n_6997, n10757);
  and g14877 (n10758, n2625, n_6997);
  not g14878 (n_6998, n10756);
  and g14879 (n10759, n_6998, n10758);
  not g14880 (n_6999, n10751);
  and g14881 (n10760, pi0087, n_6999);
  not g14882 (n_7000, n10759);
  and g14883 (n10761, n_7000, n10760);
  and g14884 (n10762, n_6990, n10761);
  and g14885 (n10763, n10502, n10737);
  and g14886 (n10764, pi0043, n_6882);
  not g14887 (n_7001, n10763);
  not g14888 (n_7002, n10764);
  and g14889 (n10765, n_7001, n_7002);
  not g14890 (n_7003, n10765);
  and g14891 (n10766, n10732, n_7003);
  not g14892 (n_7004, n10766);
  and g14893 (n10767, n10734, n_7004);
  not g14894 (n_7005, n10767);
  and g14895 (n10768, n_6983, n_7005);
  not g14896 (n_7006, n10768);
  and g14897 (n10769, n_162, n_7006);
  not g14898 (n_7007, n10769);
  and g14899 (n10770, n_6990, n_7007);
  not g14900 (n_7008, n10770);
  and g14901 (n10771, n6285, n_7008);
  and g14902 (n10772, n_6990, n_6987);
  not g14903 (n_7009, n10772);
  and g14904 (n10773, pi0038, n_7009);
  and g14905 (n10774, pi0232, n_6917);
  not g14906 (n_7010, n10774);
  and g14907 (n10775, n10641, n_7010);
  not g14908 (n_7011, n10775);
  and g14909 (n10776, pi0039, n_7011);
  and g14910 (n10777, n_188, n_6836);
  not g14911 (n_7012, n10579);
  and g14912 (n10778, n_538, n_7012);
  not g14913 (n_7013, n10572);
  and g14914 (n10779, n2924, n_7013);
  not g14915 (n_7014, n10778);
  not g14916 (n_7015, n10779);
  and g14917 (n10780, n_7014, n_7015);
  and g14918 (n10781, n6269, n10780);
  not g14919 (n_7016, n10781);
  and g14920 (n10782, pi0228, n_7016);
  not g14921 (n_7017, n10777);
  not g14922 (n_7018, n10782);
  and g14923 (n10783, n_7017, n_7018);
  not g14924 (n_7019, n10783);
  and g14925 (n10784, n_3188, n_7019);
  not g14926 (n_7020, n10731);
  and g14927 (n10785, n_6976, n_7020);
  not g14928 (n_7021, n10587);
  and g14929 (n10786, n_538, n_7021);
  and g14930 (n10787, n2924, n_6847);
  not g14931 (n_7022, n10786);
  not g14932 (n_7023, n10787);
  and g14933 (n10788, n_7022, n_7023);
  not g14934 (n_7024, n10788);
  and g14935 (n10789, pi0228, n_7024);
  and g14936 (n10790, n_188, n_6835);
  not g14937 (n_7025, n10789);
  not g14938 (n_7026, n10790);
  and g14939 (n10791, n_7025, n_7026);
  and g14940 (n10792, pi0043, n10731);
  not g14941 (n_7027, n10791);
  and g14942 (n10793, n_7027, n10792);
  not g14943 (n_7028, n10784);
  not g14944 (n_7029, n10785);
  and g14945 (n10794, n_7028, n_7029);
  not g14946 (n_7030, n10793);
  and g14947 (n10795, n_7030, n10794);
  not g14948 (n_7031, n10795);
  and g14949 (n10796, n_162, n_7031);
  not g14950 (n_7032, n10776);
  not g14951 (n_7033, n10796);
  and g14952 (n10797, n_7032, n_7033);
  not g14953 (n_7034, n10797);
  and g14954 (n10798, n2608, n_7034);
  not g14961 (n_7038, n10762);
  and g14962 (n10802, n_171, n_7038);
  not g14963 (n_7039, n10801);
  and g14964 (n10803, n_7039, n10802);
  not g14965 (n_7040, n10750);
  and g14966 (n10804, n7429, n_7040);
  not g14967 (n_7041, n10803);
  and g14968 (n10805, n_7041, n10804);
  and g14969 (n10806, n_4196, n10772);
  not g14970 (n_7042, n10806);
  and g14971 (n10807, n_6900, n_7042);
  not g14972 (n_7043, n10805);
  and g14973 (n10808, n_7043, n10807);
  not g14974 (n_7044, pi0199);
  not g14975 (n_7045, pi0200);
  and g14976 (n10809, n_7044, n_7045);
  not g14977 (n_7046, n10809);
  and g14978 (n10810, n_234, n_7046);
  not g14979 (n_7047, n10810);
  and g14980 (n10811, n_134, n_7047);
  not g14981 (n_7048, n10811);
  and g14982 (n10812, n_3410, n_7048);
  not g14983 (n_7049, n10812);
  and g14984 (n10813, n_234, n_7049);
  and g14985 (n10814, n10518, n10809);
  not g14986 (n_7050, n10814);
  and g14987 (n10815, pi0232, n_7050);
  not g14988 (n_7051, n10815);
  and g14989 (n10816, n10813, n_7051);
  not g14990 (n_7052, n10816);
  and g14991 (n10817, pi0039, n_7052);
  not g14992 (n_7053, n10817);
  and g14993 (n10818, n_6987, n_7053);
  and g14994 (n10819, n_4196, n10818);
  and g14995 (n10820, n_6991, n_7053);
  not g14996 (n_7054, n10820);
  and g14997 (n10821, pi0075, n_7054);
  and g14998 (n10822, n_7007, n_7053);
  not g14999 (n_7055, n10822);
  and g15000 (n10823, n6285, n_7055);
  not g15001 (n_7056, n10818);
  and g15002 (n10824, pi0038, n_7056);
  and g15003 (n10825, n_6869, n10809);
  not g15004 (n_7057, n10825);
  and g15005 (n10826, pi0232, n_7057);
  not g15006 (n_7058, n10826);
  and g15007 (n10827, n10813, n_7058);
  not g15008 (n_7059, n10827);
  and g15009 (n10828, pi0039, n_7059);
  not g15010 (n_7060, n10828);
  and g15011 (n10829, n_7033, n_7060);
  not g15012 (n_7061, n10829);
  and g15013 (n10830, n2608, n_7061);
  not g15020 (n_7065, n2531);
  and g15021 (n10834, n_7065, n_7056);
  not g15022 (n_7066, n10834);
  and g15023 (n10835, n10761, n_7066);
  not g15024 (n_7067, n10835);
  and g15025 (n10836, n_171, n_7067);
  not g15026 (n_7068, n10833);
  and g15027 (n10837, n_7068, n10836);
  not g15028 (n_7069, n10821);
  and g15029 (n10838, n7429, n_7069);
  not g15030 (n_7070, n10837);
  and g15031 (n10839, n_7070, n10838);
  not g15032 (n_7071, n10819);
  and g15033 (n10840, n10487, n_7071);
  not g15034 (n_7072, n10839);
  and g15035 (n10841, n_7072, n10840);
  not g15036 (n_7073, n10808);
  not g15037 (n_7074, n10841);
  and g15038 (n10842, n_7073, n_7074);
  and g15039 (n10843, pi0212, pi0214);
  not g15040 (n_7075, pi0211);
  and g15041 (n10844, n_7075, n_6791);
  not g15042 (n_7076, n10844);
  and g15043 (n10845, n10843, n_7076);
  not g15044 (n_7077, n10843);
  and g15045 (n10846, n_7075, n_7077);
  not g15046 (n_7078, n10845);
  not g15047 (n_7079, n10846);
  and g15048 (n10847, n_7078, n_7079);
  not g15049 (n_7080, n10842);
  not g15050 (n_7081, n10847);
  and g15051 (n10848, n_7080, n_7081);
  and g15052 (n10849, n10525, n_6907);
  not g15053 (n_7082, n10849);
  and g15054 (n10850, n_6991, n_7082);
  not g15055 (n_7083, n10850);
  and g15056 (n10851, pi0075, n_7083);
  and g15057 (n10852, n10761, n_7082);
  and g15058 (n10853, n_7007, n_7082);
  not g15059 (n_7084, n10853);
  and g15060 (n10854, n6285, n_7084);
  and g15061 (n10855, n_6987, n_7082);
  not g15062 (n_7085, n10855);
  and g15063 (n10856, pi0038, n_7085);
  and g15064 (n10857, n10602, n_6917);
  and g15065 (n10858, n_6872, n10640);
  not g15066 (n_7086, n10858);
  and g15067 (n10859, n_6873, n_7086);
  not g15068 (n_7087, n10857);
  and g15069 (n10860, n_7087, n10859);
  not g15070 (n_7088, n10860);
  and g15071 (n10861, pi0039, n_7088);
  not g15072 (n_7089, n10861);
  and g15073 (n10862, n_7033, n_7089);
  not g15074 (n_7090, n10862);
  and g15075 (n10863, n2608, n_7090);
  not g15082 (n_7094, n10852);
  and g15083 (n10867, n_171, n_7094);
  not g15084 (n_7095, n10866);
  and g15085 (n10868, n_7095, n10867);
  not g15086 (n_7096, n10851);
  and g15087 (n10869, n7429, n_7096);
  not g15088 (n_7097, n10868);
  and g15089 (n10870, n_7097, n10869);
  and g15090 (n10871, n_4196, n10855);
  not g15091 (n_7098, n10871);
  and g15092 (n10872, n_6900, n_7098);
  not g15093 (n_7099, n10870);
  and g15094 (n10873, n_7099, n10872);
  and g15095 (n10874, n_6816, n10817);
  not g15096 (n_7100, n10874);
  and g15097 (n10875, n_6987, n_7100);
  and g15098 (n10876, n_4196, n10875);
  and g15099 (n10877, n_6991, n_7100);
  not g15100 (n_7101, n10877);
  and g15101 (n10878, pi0075, n_7101);
  and g15102 (n10879, n10761, n_7100);
  and g15103 (n10880, n_7007, n_7100);
  not g15104 (n_7102, n10880);
  and g15105 (n10881, n6285, n_7102);
  not g15106 (n_7103, n10875);
  and g15107 (n10882, pi0038, n_7103);
  and g15108 (n10883, n10602, n_7057);
  and g15109 (n10884, n_6873, n_7049);
  not g15110 (n_7104, n10883);
  and g15111 (n10885, n_7104, n10884);
  not g15112 (n_7105, n10885);
  and g15113 (n10886, pi0039, n_7105);
  not g15114 (n_7106, n10886);
  and g15115 (n10887, n_7033, n_7106);
  not g15116 (n_7107, n10887);
  and g15117 (n10888, n2608, n_7107);
  not g15124 (n_7111, n10879);
  and g15125 (n10892, n_171, n_7111);
  not g15126 (n_7112, n10891);
  and g15127 (n10893, n_7112, n10892);
  not g15128 (n_7113, n10878);
  and g15129 (n10894, n7429, n_7113);
  not g15130 (n_7114, n10893);
  and g15131 (n10895, n_7114, n10894);
  not g15132 (n_7115, n10876);
  and g15133 (n10896, n10487, n_7115);
  not g15134 (n_7116, n10895);
  and g15135 (n10897, n_7116, n10896);
  not g15136 (n_7117, n10873);
  not g15137 (n_7118, n10897);
  and g15138 (n10898, n_7117, n_7118);
  not g15139 (n_7119, n10898);
  and g15140 (n10899, n10847, n_7119);
  not g15141 (n_7120, n10848);
  and g15142 (n10900, n_4226, n_7120);
  not g15143 (n_7121, n10899);
  and g15144 (n10901, n_7121, n10900);
  and g15145 (n10902, n10523, n10847);
  not g15146 (n_7122, n10902);
  and g15147 (n10903, pi0039, n_7122);
  and g15148 (n10904, po1038, n_6987);
  not g15149 (n_7123, n10903);
  and g15150 (n10905, n_7123, n10904);
  or g15151 (po0201, n10901, n10905);
  and g15152 (n10907, n_134, n7474);
  not g15153 (n_7124, n10907);
  and g15154 (n10908, pi0039, n_7124);
  and g15155 (n10909, pi0044, n_134);
  not g15156 (n_7125, n10909);
  and g15157 (n10910, n_162, n_7125);
  not g15158 (n_7126, n10908);
  not g15159 (n_7127, n10910);
  and g15160 (n10911, n_7126, n_7127);
  and g15161 (n10912, n_6666, n10911);
  and g15162 (n10913, n_4137, n_7125);
  not g15163 (n_7128, n10913);
  and g15164 (n10914, n_162, n_7128);
  and g15165 (n10915, n_538, n10909);
  not g15166 (n_7129, n10915);
  and g15167 (n10916, n7506, n_7129);
  and g15168 (n10917, n7594, n_6729);
  and g15169 (n10918, n7479, n10316);
  and g15170 (n10919, n7477, n10918);
  not g15171 (n_7130, n10327);
  and g15172 (n10920, pi0044, n_7130);
  not g15173 (n_7131, n10919);
  not g15174 (n_7132, n10920);
  and g15175 (n10921, n_7131, n_7132);
  not g15176 (n_7133, n10921);
  and g15177 (n10922, n10917, n_7133);
  not g15178 (n_7134, n10922);
  and g15179 (n10923, n10916, n_7134);
  not g15180 (n_7135, n10923);
  and g15181 (n10924, n10914, n_7135);
  and g15182 (n10925, pi0039, n7474);
  and g15183 (n10926, n_134, n10925);
  not g15184 (n_7136, n10924);
  not g15185 (n_7137, n10926);
  and g15186 (n10927, n_7136, n_7137);
  not g15187 (n_7138, n10927);
  and g15188 (n10928, n2620, n_7138);
  not g15189 (n_7139, n10912);
  and g15190 (n10929, pi0075, n_7139);
  not g15191 (n_7140, n10928);
  and g15192 (n10930, n_7140, n10929);
  and g15193 (n10931, pi0228, n2608);
  and g15194 (n10932, n10316, n10931);
  and g15195 (n10933, n10342, n10931);
  not g15196 (n_7141, n10933);
  and g15197 (n10934, n10909, n_7141);
  not g15198 (n_7142, n10934);
  and g15199 (n10935, n_162, n_7142);
  not g15200 (n_7143, n10932);
  and g15201 (n10936, n_7143, n10935);
  and g15202 (n10937, pi0087, n_7126);
  not g15203 (n_7144, n10936);
  and g15204 (n10938, n_7144, n10937);
  not g15205 (n_7145, n10911);
  and g15206 (n10939, pi0038, n_7145);
  and g15207 (n10940, n7479, n10342);
  not g15208 (n_7146, n10940);
  and g15209 (n10941, pi0044, n_7146);
  not g15210 (n_7147, n10918);
  not g15211 (n_7148, n10941);
  and g15212 (n10942, n_7147, n_7148);
  not g15213 (n_7149, n10942);
  and g15214 (n10943, n10917, n_7149);
  not g15215 (n_7150, n10943);
  and g15216 (n10944, n10916, n_7150);
  not g15217 (n_7151, n10944);
  and g15218 (n10945, n10914, n_7151);
  and g15219 (n10946, n6285, n_7137);
  not g15220 (n_7152, n10945);
  and g15221 (n10947, n_7152, n10946);
  and g15222 (n10948, pi0287, n10342);
  not g15223 (n_7153, n10948);
  and g15224 (n10949, n_134, n_7153);
  and g15225 (n10950, n10925, n10949);
  and g15226 (n10951, pi0044, n10407);
  not g15227 (n_7154, n10951);
  and g15228 (n10952, n_188, n_7154);
  not g15229 (n_7155, n10400);
  and g15230 (n10953, n_7155, n10952);
  and g15231 (n10954, pi0044, n10455);
  not g15232 (n_7156, n10450);
  and g15233 (n10955, n2924, n_7156);
  not g15234 (n_7157, n10954);
  and g15235 (n10956, n_7157, n10955);
  and g15236 (n10957, pi0044, n10422);
  not g15237 (n_7158, n10432);
  and g15238 (n10958, n_538, n_7158);
  not g15239 (n_7159, n10957);
  and g15240 (n10959, n_7159, n10958);
  not g15241 (n_7160, n10956);
  not g15242 (n_7161, n10959);
  and g15243 (n10960, n_7160, n_7161);
  not g15244 (n_7162, n10960);
  and g15245 (n10961, pi0228, n_7162);
  not g15246 (n_7163, n10953);
  and g15247 (n10962, n_162, n_7163);
  not g15248 (n_7164, n10961);
  and g15249 (n10963, n_7164, n10962);
  not g15250 (n_7165, n10950);
  and g15251 (n10964, n2608, n_7165);
  not g15252 (n_7166, n10963);
  and g15253 (n10965, n_7166, n10964);
  not g15260 (n_7170, n10938);
  and g15261 (n10969, n_171, n_7170);
  not g15262 (n_7171, n10968);
  and g15263 (n10970, n_7171, n10969);
  not g15264 (n_7172, n10930);
  not g15265 (n_7173, n10970);
  and g15266 (n10971, n_7172, n_7173);
  not g15267 (n_7174, n10971);
  and g15268 (n10972, n7429, n_7174);
  and g15269 (n10973, n_4196, n_7145);
  not g15270 (n_7175, n10973);
  and g15271 (n10974, n_4226, n_7175);
  not g15272 (n_7176, n10972);
  and g15273 (n10975, n_7176, n10974);
  and g15274 (n10976, n2639, n7473);
  and g15275 (n10977, n_134, n10976);
  not g15276 (n_7177, n10977);
  and g15277 (n10978, pi0039, n_7177);
  and g15278 (n10979, po1038, n_7127);
  not g15279 (n_7178, n10978);
  and g15280 (n10980, n_7178, n10979);
  or g15281 (po0202, n10975, n10980);
  and g15282 (n10982, n_161, pi0039);
  and g15283 (n10983, n10197, n10982);
  and g15284 (n10984, pi0979, n10983);
  and g15285 (po0203, n6380, n10984);
  and g15286 (n10986, n_53, n_85);
  and g15287 (n10987, n_95, n10986);
  and g15288 (n10988, n_83, n_73);
  and g15289 (n10989, n8909, n10988);
  and g15301 (n11001, n_3052, n11000);
  and g15302 (n11002, n2702, n2888);
  and g15303 (n11003, pi0024, n11002);
  not g15304 (n_7179, n11001);
  not g15305 (n_7180, n11003);
  and g15306 (n11004, n_7179, n_7180);
  not g15307 (n_7181, n11004);
  and g15308 (po0204, n10166, n_7181);
  and g15309 (n11006, n_94, n2474);
  not g15314 (n_7182, n11010);
  and g15315 (n11011, n_97, n_7182);
  and g15316 (n11012, n8916, n9081);
  and g15317 (n11013, n_64, n_61);
  and g15318 (n11014, n2487, n11013);
  and g15323 (n11018, n_416, n11017);
  not g15324 (n_7184, n11018);
  and g15325 (n11019, n_46, n_7184);
  and g15326 (n11020, n_442, n7438);
  not g15327 (n_7185, n11019);
  and g15328 (n11021, n2754, n_7185);
  and g15329 (n11022, n11020, n11021);
  and g15330 (n11023, n2700, n11022);
  not g15331 (n_7186, n11023);
  and g15332 (n11024, n_6594, n_7186);
  not g15333 (n_7187, n11024);
  and g15334 (n11025, n10162, n_7187);
  not g15335 (n_7188, n11025);
  and g15336 (n11026, n7490, n_7188);
  and g15337 (n11027, n_97, n11017);
  not g15338 (n_7189, n11027);
  and g15339 (n11028, n_46, n_7189);
  not g15340 (n_7190, n11028);
  and g15341 (n11029, n11020, n_7190);
  and g15342 (n11030, n10186, n11029);
  and g15343 (n11031, n_3126, n2932);
  and g15344 (n11032, n11030, n11031);
  and g15345 (n11033, n_6605, n11025);
  not g15346 (n_7191, n11032);
  and g15347 (n11034, pi0829, n_7191);
  not g15348 (n_7192, n11033);
  and g15349 (n11035, n_7192, n11034);
  and g15350 (n11036, n_489, n11035);
  not g15351 (n_7193, n11026);
  not g15352 (n_7194, n11036);
  and g15353 (n11037, n_7193, n_7194);
  not g15354 (n_7195, n11037);
  and g15355 (n11038, pi1091, n_7195);
  not g15356 (n_7196, n7417);
  and g15357 (n11039, n_7196, n11025);
  not g15358 (n_7197, n11039);
  and g15359 (n11040, n_3127, n_7197);
  not g15360 (n_7198, n11035);
  not g15361 (n_7199, n11040);
  and g15362 (n11041, n_7198, n_7199);
  not g15363 (n_7200, n11041);
  and g15364 (n11042, n_3206, n_7200);
  and g15365 (n11043, n7417, n10162);
  and g15366 (n11044, n_6595, n11043);
  and g15367 (n11045, n_3285, n_4214);
  not g15368 (n_7201, n11044);
  not g15369 (n_7202, n11045);
  and g15370 (n11046, n_7201, n_7202);
  and g15371 (n11047, n_7197, n11046);
  and g15378 (n11051, n_134, pi0841);
  and g15379 (n11052, n2705, n11051);
  and g15384 (n11057, n2464, n2487);
  and g15385 (n11058, n_61, n2804);
  and g15386 (n11059, n10245, n11058);
  and g15387 (n11060, n8909, n8916);
  and g15388 (n11061, n11059, n11060);
  and g15394 (n11067, n2706, n8935);
  and g15395 (n11068, n11066, n11067);
  and g15396 (n11069, n10161, n11052);
  and g15397 (n11070, n11068, n11069);
  not g15398 (n_7206, n11070);
  and g15399 (n11071, n_168, n_7206);
  and g15400 (n11072, pi0074, n_6576);
  and g15406 (n11076, pi0024, n8897);
  not g15407 (n_7209, n10374);
  not g15408 (n_7210, n11076);
  and g15409 (n11077, n_7209, n_7210);
  and g15410 (n11078, n_280, n_5631);
  and g15411 (n11079, pi0252, n_5636);
  not g15412 (n_7211, n11078);
  not g15413 (n_7212, n11079);
  and g15414 (n11080, n_7211, n_7212);
  and g15415 (n11081, pi0024, n_125);
  not g15416 (n_7213, n8899);
  and g15417 (n11082, n_7213, n11081);
  and g15423 (n11086, n2962, n7450);
  not g15429 (n_7217, n11085);
  not g15430 (n_7218, n11090);
  and g15431 (n11091, n_7217, n_7218);
  not g15432 (n_7219, n11091);
  and g15433 (n11092, n_164, n_7219);
  and g15434 (n11093, pi0100, n_3214);
  and g15435 (n11094, n6353, n11093);
  not g15436 (n_7220, n11092);
  not g15437 (n_7221, n11094);
  and g15438 (n11095, n_7220, n_7221);
  and g15439 (n11096, n2530, n2533);
  not g15440 (n_7222, n11095);
  and g15441 (n11097, n_7222, n11096);
  and g15442 (n11098, n6282, n8967);
  and g15443 (n11099, n8963, n11098);
  not g15444 (n_7223, n11097);
  not g15445 (n_7224, n11099);
  and g15446 (n11100, n_7223, n_7224);
  not g15447 (n_7225, n11100);
  and g15448 (po0208, n8881, n_7225);
  and g15449 (n11102, n9082, n11057);
  and g15450 (n11103, n2467, n11102);
  and g15451 (n11104, n_65, n11103);
  and g15452 (n11105, n2804, n11104);
  and g15453 (n11106, n2700, n10166);
  and g15454 (n11107, n2754, n11106);
  and g15455 (n11108, n2807, n11105);
  and g15456 (po0209, n11107, n11108);
  and g15457 (n11110, n_6791, n10846);
  and g15458 (n11111, pi0052, n_134);
  not g15459 (n_7226, n11111);
  and g15460 (n11112, n_162, n_7226);
  not g15461 (n_7227, n10525);
  not g15462 (n_7228, n11112);
  and g15463 (n11113, n_7227, n_7228);
  not g15464 (n_7229, n11113);
  and g15465 (n11114, n_4196, n_7229);
  and g15466 (n11115, n_6873, n10609);
  not g15467 (n_7230, n11115);
  and g15468 (n11116, pi0039, n_7230);
  and g15469 (n11117, n6267, n6270);
  not g15470 (n_7231, n11117);
  and g15471 (n11118, n_7226, n_7231);
  and g15472 (n11119, n_3190, n10558);
  and g15473 (n11120, pi0052, n10554);
  not g15474 (n_7232, n11119);
  and g15475 (n11121, n11117, n_7232);
  not g15476 (n_7233, n11120);
  and g15477 (n11122, n_7233, n11121);
  not g15478 (n_7234, n11118);
  and g15479 (n11123, n_188, n_7234);
  not g15480 (n_7235, n11122);
  and g15481 (n11124, n_7235, n11123);
  and g15482 (n11125, n_3197, n6267);
  and g15483 (n11126, n_3190, n10573);
  and g15484 (n11127, pi0052, n10570);
  not g15485 (n_7236, n11126);
  and g15486 (n11128, n10491, n_7236);
  not g15487 (n_7237, n11127);
  and g15488 (n11129, n_7237, n11128);
  and g15489 (n11130, n_3190, n10580);
  and g15490 (n11131, pi0052, n10587);
  not g15491 (n_7238, n11130);
  and g15492 (n11132, n10578, n_7238);
  not g15493 (n_7239, n11131);
  and g15494 (n11133, n_7239, n11132);
  not g15495 (n_7240, n11129);
  not g15496 (n_7241, n11133);
  and g15497 (n11134, n_7240, n_7241);
  not g15498 (n_7242, n11134);
  and g15499 (n11135, n11125, n_7242);
  and g15500 (n11136, pi0228, n_7234);
  not g15501 (n_7243, n11135);
  and g15502 (n11137, n_7243, n11136);
  not g15503 (n_7244, n11124);
  and g15504 (n11138, n_162, n_7244);
  not g15505 (n_7245, n11137);
  and g15506 (n11139, n_7245, n11138);
  not g15507 (n_7246, n11116);
  not g15508 (n_7247, n11139);
  and g15509 (n11140, n_7246, n_7247);
  not g15510 (n_7248, n11140);
  and g15511 (n11141, n2608, n_7248);
  and g15512 (n11142, pi0038, n_7229);
  and g15513 (n11143, n7506, n10491);
  and g15514 (n11144, n11125, n11143);
  and g15515 (n11145, n7479, n11144);
  and g15516 (n11146, n10616, n11145);
  not g15517 (n_7249, n11146);
  and g15518 (n11147, n11111, n_7249);
  not g15519 (n_7250, n11147);
  and g15520 (n11148, n_162, n_7250);
  not g15521 (n_7251, n11148);
  and g15522 (n11149, n_7227, n_7251);
  not g15523 (n_7252, n11149);
  and g15524 (n11150, n6285, n_7252);
  not g15525 (n_7253, n11142);
  not g15526 (n_7254, n11150);
  and g15527 (n11151, n_7253, n_7254);
  not g15528 (n_7255, n11141);
  and g15529 (n11152, n_7255, n11151);
  not g15530 (n_7256, n11152);
  and g15531 (n11153, n_172, n_7256);
  and g15532 (n11154, n_958, n11113);
  not g15533 (n_7257, n11154);
  and g15534 (n11155, pi0087, n_7257);
  and g15535 (n11156, pi0228, n11117);
  and g15536 (n11157, n_3190, n10501);
  and g15537 (n11158, pi0052, n10617);
  not g15538 (n_7258, n11157);
  not g15539 (n_7259, n11158);
  and g15540 (n11159, n_7258, n_7259);
  not g15541 (n_7260, n11159);
  and g15542 (n11160, n11156, n_7260);
  not g15543 (n_7261, n11156);
  and g15544 (n11161, n11111, n_7261);
  not g15545 (n_7262, n11160);
  not g15546 (n_7263, n11161);
  and g15547 (n11162, n_7262, n_7263);
  and g15548 (n11163, n_162, n11162);
  and g15549 (n11164, n2608, n_7227);
  not g15550 (n_7264, n11163);
  and g15551 (n11165, n_7264, n11164);
  not g15552 (n_7265, n11165);
  and g15553 (n11166, n11155, n_7265);
  not g15554 (n_7266, n11166);
  and g15555 (n11167, n10487, n_7266);
  not g15556 (n_7267, n11153);
  and g15557 (n11168, n_7267, n11167);
  and g15558 (n11169, n_7053, n_7228);
  and g15559 (n11170, n_958, n11169);
  and g15560 (n11171, n2608, n_7100);
  and g15561 (n11172, n_7264, n11171);
  not g15562 (n_7268, n11170);
  and g15563 (n11173, n11155, n_7268);
  not g15564 (n_7269, n11172);
  and g15565 (n11174, n_7269, n11173);
  and g15566 (n11175, n_7106, n_7247);
  not g15567 (n_7270, n11175);
  and g15568 (n11176, n2608, n_7270);
  and g15569 (n11177, n_7100, n_7251);
  not g15570 (n_7271, n11177);
  and g15571 (n11178, n6285, n_7271);
  not g15572 (n_7272, n11169);
  and g15573 (n11179, pi0038, n_7272);
  and g15574 (n11180, n_7229, n11179);
  not g15575 (n_7273, n11178);
  not g15576 (n_7274, n11180);
  and g15577 (n11181, n_7273, n_7274);
  not g15578 (n_7275, n11176);
  and g15579 (n11182, n_7275, n11181);
  not g15580 (n_7276, n11182);
  and g15581 (n11183, n_172, n_7276);
  not g15582 (n_7277, n11174);
  and g15583 (n11184, n_6900, n_7277);
  not g15584 (n_7278, n11183);
  and g15585 (n11185, n_7278, n11184);
  not g15586 (n_7279, n11168);
  not g15587 (n_7280, n11185);
  and g15588 (n11186, n_7279, n_7280);
  not g15589 (n_7281, n11186);
  and g15590 (n11187, n_171, n_7281);
  and g15591 (n11188, n10498, n11144);
  and g15592 (n11189, n2620, n11188);
  and g15593 (n11190, n_162, n11111);
  not g15594 (n_7282, n11189);
  and g15595 (n11191, n_7282, n11190);
  not g15596 (n_7283, n11191);
  and g15597 (n11192, n_162, n_7283);
  and g15598 (n11193, n_6900, n10874);
  and g15599 (n11194, n10487, n10525);
  not g15606 (n_7287, n11197);
  and g15607 (n11198, n7429, n_7287);
  not g15608 (n_7288, n11187);
  and g15609 (n11199, n_7288, n11198);
  not g15610 (n_7289, n11114);
  and g15611 (n11200, n11110, n_7289);
  not g15612 (n_7290, n11199);
  and g15613 (n11201, n_7290, n11200);
  and g15614 (n11202, n_4196, n_6900);
  and g15615 (n11203, n11169, n11202);
  not g15616 (n_7291, n11190);
  and g15617 (n11204, n_4196, n_7291);
  and g15618 (n11205, pi0075, n11191);
  and g15619 (n11206, pi0100, n_7291);
  and g15620 (n11207, pi0038, n_7291);
  and g15621 (n11208, n_161, n11162);
  not g15622 (n_7292, n11207);
  not g15623 (n_7293, n11208);
  and g15624 (n11209, n_7292, n_7293);
  not g15625 (n_7294, n11209);
  and g15626 (n11210, n_164, n_7294);
  and g15627 (n11211, n_164, n10982);
  not g15628 (n_7295, n11211);
  and g15629 (n11212, pi0087, n_7295);
  not g15630 (n_7296, n11206);
  and g15631 (n11213, n_7296, n11212);
  not g15632 (n_7297, n11210);
  and g15633 (n11214, n_7297, n11213);
  and g15634 (n11215, pi0100, n_7250);
  and g15635 (n11216, n_164, n11139);
  not g15636 (n_7298, n11215);
  and g15637 (n11217, n_162, n_7298);
  not g15638 (n_7299, n11216);
  and g15639 (n11218, n_7299, n11217);
  not g15640 (n_7300, n11218);
  and g15641 (n11219, n_161, n_7300);
  and g15642 (n11220, n_172, n_7292);
  not g15643 (n_7301, n11219);
  and g15644 (n11221, n_7301, n11220);
  not g15645 (n_7302, n11214);
  not g15646 (n_7303, n11221);
  and g15647 (n11222, n_7302, n_7303);
  not g15648 (n_7304, n11222);
  and g15649 (n11223, n_171, n_7304);
  not g15650 (n_7305, n11205);
  and g15651 (n11224, n7429, n_7305);
  not g15652 (n_7306, n11223);
  and g15653 (n11225, n_7306, n11224);
  not g15654 (n_7307, n11204);
  and g15655 (n11226, n10487, n_7307);
  not g15656 (n_7308, n11225);
  and g15657 (n11227, n_7308, n11226);
  and g15658 (n11228, n2608, n_7053);
  and g15659 (n11229, n_7264, n11228);
  not g15660 (n_7309, n11229);
  and g15661 (n11230, n_7268, n_7309);
  not g15662 (n_7310, n11230);
  and g15663 (n11231, pi0087, n_7310);
  and g15664 (n11232, n_7060, n_7247);
  not g15665 (n_7311, n11232);
  and g15666 (n11233, n2608, n_7311);
  and g15667 (n11234, n_7053, n_7251);
  not g15668 (n_7312, n11234);
  and g15669 (n11235, n6285, n_7312);
  not g15676 (n_7316, n11231);
  and g15677 (n11239, n_171, n_7316);
  not g15678 (n_7317, n11238);
  and g15679 (n11240, n_7317, n11239);
  and g15680 (n11241, n_6666, n11169);
  not g15681 (n_7318, n11188);
  and g15682 (n11242, n11111, n_7318);
  not g15683 (n_7319, n11242);
  and g15684 (n11243, n_162, n_7319);
  and g15685 (n11244, n2620, n_7053);
  not g15686 (n_7320, n11243);
  and g15687 (n11245, n_7320, n11244);
  not g15688 (n_7321, n11241);
  and g15689 (n11246, pi0075, n_7321);
  not g15690 (n_7322, n11245);
  and g15691 (n11247, n_7322, n11246);
  not g15697 (n_7325, n11227);
  not g15698 (n_7326, n11250);
  and g15699 (n11251, n_7325, n_7326);
  not g15700 (n_7327, n11110);
  not g15701 (n_7328, n11251);
  and g15702 (n11252, n_7327, n_7328);
  and g15709 (n11256, pi0039, n11110);
  and g15710 (n11257, n10523, n11256);
  and g15711 (n11258, po1038, n_7291);
  not g15712 (n_7332, n11257);
  and g15713 (n11259, n_7332, n11258);
  not g15714 (n_7333, n11255);
  not g15715 (n_7334, n11259);
  and g15716 (po0210, n_7333, n_7334);
  and g15717 (n11261, n_3084, n_3080);
  and g15718 (n11262, n6181, n11261);
  not g15719 (n_7335, n11262);
  and g15720 (n11263, pi0039, n_7335);
  and g15721 (n11264, pi0024, n10162);
  and g15725 (n11268, n11264, n11267);
  not g15726 (n_7336, n11268);
  and g15727 (n11269, n_162, n_7336);
  not g15728 (n_7337, n11263);
  and g15733 (n11273, n8897, n9254);
  and g15742 (n11282, n11273, n11281);
  and g15743 (n11283, n_3052, n2704);
  and g15744 (n11284, n8960, n11283);
  not g15748 (n_7339, n11287);
  and g15749 (n11288, n_167, n_7339);
  and g15750 (n11289, n2621, n10195);
  not g15751 (n_7340, n11289);
  and g15752 (n11290, pi0054, n_7340);
  not g15753 (n_7341, n11288);
  and g15754 (n11291, n8880, n_7341);
  not g15755 (n_7342, n11290);
  and g15756 (po0212, n_7342, n11291);
  and g15757 (n11293, n_167, n11289);
  and g15758 (n11294, n_168, n11293);
  not g15759 (n_7343, n11294);
  and g15760 (n11295, pi0055, n_7343);
  and g15765 (n11300, n6479, n9500);
  and g15766 (n11301, n2465, n2572);
  and g15767 (n11302, n11300, n11301);
  and g15768 (n11303, n11299, n11302);
  not g15769 (n_7344, n11303);
  and g15770 (n11304, n_176, n_7344);
  not g15771 (n_7345, n11304);
  and g15772 (n11305, n8878, n_7345);
  not g15773 (n_7346, n11295);
  and g15774 (po0213, n_7346, n11305);
  and g15775 (n11307, n2518, n2537);
  and g15776 (n11308, n6172, n11307);
  not g15777 (n_7347, n11308);
  and g15778 (n11309, pi0056, n_7347);
  and g15779 (n11310, pi0056, n_158);
  and g15780 (n11311, pi0055, n10068);
  not g15781 (n_7348, n11310);
  not g15782 (n_7349, n11311);
  and g15783 (n11312, n_7348, n_7349);
  not g15784 (n_7350, n11309);
  and g15785 (n11313, n3328, n_7350);
  not g15786 (n_7351, n11312);
  and g15787 (po0214, n_7351, n11313);
  and g15788 (n11315, n6304, n11294);
  not g15789 (n_7352, n11315);
  and g15790 (n11316, pi0057, n_7352);
  and g15791 (n11317, n6485, n11307);
  and g15792 (n11318, n_157, pi0062);
  not g15793 (n_7354, pi0924);
  and g15794 (n11319, n_7354, n11318);
  not g15795 (n_7355, n11319);
  and g15796 (n11320, n_7348, n_7355);
  not g15797 (n_7356, n11320);
  and g15798 (n11321, n11317, n_7356);
  not g15799 (n_7357, n11321);
  and g15800 (n11322, n_796, n_7357);
  not g15801 (n_7358, n11316);
  and g15802 (n11323, n_792, n_7358);
  not g15803 (n_7359, n11322);
  and g15804 (po0215, n_7359, n11323);
  and g15805 (n11325, n_131, n11086);
  and g15806 (n11326, n10165, n11325);
  and g15807 (po0216, n7433, n11326);
  and g15808 (n11328, pi0059, n_7352);
  and g15809 (n11329, pi0924, n11318);
  and g15810 (n11330, n11317, n11329);
  not g15811 (n_7360, n11330);
  and g15812 (n11331, n_792, n_7360);
  not g15813 (n_7361, n11328);
  and g15814 (n11332, n_796, n_7361);
  not g15815 (n_7362, n11331);
  and g15816 (po0217, n_7362, n11332);
  not g15824 (n_7363, n11337);
  not g15825 (n_7364, n11340);
  and g15826 (n11341, n_7363, n_7364);
  not g15827 (n_7365, n11341);
  and g15828 (po0218, n10200, n_7365);
  and g15829 (n11343, pi0841, n11000);
  and g15830 (n11344, n_4119, n11273);
  and g15831 (n11345, n2718, n11344);
  not g15832 (n_7366, n11343);
  not g15833 (n_7367, n11345);
  and g15834 (n11346, n_7366, n_7367);
  not g15835 (n_7368, n11346);
  and g15836 (po0219, n10166, n_7368);
  and g15837 (n11348, pi0057, n_6535);
  and g15838 (n11349, n11308, n11318);
  not g15839 (n_7369, n11349);
  and g15840 (n11350, n_796, n_7369);
  not g15841 (n_7370, n11348);
  and g15842 (n11351, n_792, n_7370);
  not g15843 (n_7371, n11350);
  and g15844 (po0220, n_7371, n11351);
  and g15845 (n11353, n2861, n8935);
  and g15846 (n11354, n9100, n11353);
  and g15847 (n11355, pi0999, n11354);
  and g15848 (n11356, n_4119, n11002);
  not g15849 (n_7373, n11355);
  not g15850 (n_7374, n11356);
  and g15851 (n11357, n_7373, n_7374);
  not g15852 (n_7375, n11357);
  and g15853 (po0221, n10166, n_7375);
  and g15854 (n11359, n_100, pi0107);
  and g15855 (n11360, n9100, n11359);
  not g15856 (n_7376, n11360);
  and g15857 (n11361, n_3052, n_7376);
  and g15858 (n11362, n2486, n11359);
  not g15859 (n_7377, n11362);
  and g15860 (n11363, n_103, n_7377);
  not g15861 (n_7378, n11363);
  and g15862 (n11364, n2465, n_7378);
  and g15863 (n11365, n10169, n11364);
  not g15864 (n_7379, n11365);
  and g15865 (n11366, pi0841, n_7379);
  not g15866 (n_7380, n11361);
  and g15867 (n11367, n11107, n_7380);
  not g15868 (n_7381, n11366);
  and g15869 (po0222, n_7381, n11367);
  and g15870 (n11369, pi0039, n10201);
  and g15876 (n11373, pi0199, n_234);
  and g15877 (n11374, n2570, n2608);
  and g15878 (n11375, pi0314, n2464);
  and g15879 (n11376, n11300, n11375);
  not g15886 (n_7384, n11382);
  and g15887 (n11383, n_6791, n_7384);
  and g15888 (n11384, n_7044, n_234);
  and g15889 (n11385, n2572, n11379);
  not g15890 (n_7385, n11384);
  and g15891 (n11386, n_7385, n11385);
  not g15892 (n_7386, n11386);
  and g15893 (n11387, pi0219, n_7386);
  not g15894 (n_7387, n11383);
  and g15895 (n11388, n_4226, n_7387);
  not g15896 (n_7388, n11387);
  and g15897 (po0224, n_7388, n11388);
  and g15903 (n11395, n_3164, n6396);
  and g15904 (n11396, n3310, n5853);
  and g15905 (n11397, n11395, n11396);
  and g15906 (n11398, n_3122, n6396);
  and g15907 (n11399, n3351, n3470);
  and g15908 (n11400, n11398, n11399);
  not g15909 (n_7389, n11397);
  not g15910 (n_7390, n11400);
  and g15911 (n11401, n_7389, n_7390);
  not g15912 (n_7391, n11401);
  and g15913 (po0226, n10983, n_7391);
  and g15914 (n11403, pi0069, n11058);
  and g15915 (n11404, n10153, n11403);
  not g15916 (n_7392, n11404);
  and g15917 (n11405, n_57, n_7392);
  not g15927 (n_7394, n11409);
  not g15928 (n_7395, n11413);
  and g15929 (n11414, n_7394, n_7395);
  not g15930 (n_7396, n11414);
  and g15931 (po0227, n11107, n_7396);
  and g15932 (n11416, n2505, n2749);
  and g15933 (n11417, n_135, n11416);
  and g15934 (n11418, n10194, n11417);
  and g15935 (n11419, pi0198, pi0589);
  and g15936 (n11420, n3471, n_3122);
  and g15937 (n11421, n11419, n11420);
  and g15938 (n11422, pi0210, pi0589);
  and g15939 (n11423, n_26, n5853);
  and g15940 (n11424, n_20, n11423);
  and g15941 (n11425, n_3164, n11424);
  and g15942 (n11426, n11422, n11425);
  not g15943 (n_7398, n11421);
  not g15944 (n_7399, n11426);
  and g15945 (n11427, n_7398, n_7399);
  not g15949 (n_7402, n11427);
  not g15951 (n_7403, n11430);
  and g15952 (n11431, n_3084, n_7403);
  not g15953 (n_7404, n11431);
  and g15954 (n11432, pi0039, n_7404);
  and g15955 (n11433, n2521, n11432);
  not g15956 (n_7405, n11418);
  not g15957 (n_7406, n11433);
  and g15958 (n11434, n_7405, n_7406);
  not g15959 (n_7407, n11434);
  and g15960 (po0228, n10200, n_7407);
  and g15961 (n11436, n2469, n2481);
  and g15962 (n11437, n6424, n11436);
  and g15963 (n11438, n11014, n11437);
  and g15964 (n11439, n_103, n8916);
  and g15965 (n11440, n11438, n11439);
  not g15966 (n_7408, n11440);
  and g15967 (n11441, n_105, n_7408);
  and g15968 (n11442, n_51, n8935);
  and g15969 (n11443, n6444, n11442);
  and g15970 (n11444, n_7044, pi0200);
  and g15971 (n11445, n_234, n11444);
  and g15972 (n11446, pi0211, n_6791);
  and g15973 (n11447, pi0299, n11446);
  not g15974 (n_7409, n11445);
  not g15975 (n_7410, n11447);
  and g15976 (n11448, n_7409, n_7410);
  not g15977 (n_7411, n11448);
  not g15986 (n_7413, n11452);
  not g15987 (n_7414, n11455);
  and g15988 (n11456, n_7413, n_7414);
  not g15989 (n_7415, n11456);
  and g15990 (po0229, n10165, n_7415);
  and g15991 (n11458, pi0024, n2709);
  and g15992 (n11459, pi0072, n11458);
  and g15993 (n11460, pi0088, n10147);
  not g15997 (n_7416, n11459);
  not g15998 (n_7417, n11463);
  and g15999 (n11464, n_7416, n_7417);
  not g16000 (n_7418, n11464);
  and g16001 (n11465, n6479, n_7418);
  not g16002 (n_7419, n11465);
  and g16003 (n11466, n_162, n_7419);
  and g16004 (n11467, n7604, n11395);
  and g16005 (n11468, n7608, n11398);
  not g16006 (n_7420, n11467);
  and g16007 (n11469, pi0039, n_7420);
  not g16008 (n_7421, n11468);
  and g16009 (n11470, n_7421, n11469);
  not g16010 (n_7422, n11470);
  and g16011 (n11471, n10200, n_7422);
  not g16012 (n_7423, n11466);
  and g16013 (po0230, n_7423, n11471);
  and g16014 (n11473, n_3310, pi1050);
  and g16015 (n11474, n9090, n10162);
  and g16016 (n11475, n11473, n11474);
  not g16017 (n_7425, n11475);
  and g16018 (n11476, n_162, n_7425);
  and g16019 (n11477, n9051, n11398);
  not g16020 (n_7426, n11477);
  and g16021 (n11478, n_234, n_7426);
  and g16022 (n11479, n9036, n11395);
  not g16023 (n_7427, n11479);
  and g16024 (n11480, pi0299, n_7427);
  not g16025 (n_7428, n11478);
  not g16026 (n_7429, n11480);
  and g16027 (n11481, n_7428, n_7429);
  not g16028 (n_7430, n11481);
  and g16029 (n11482, pi0039, n_7430);
  not g16030 (n_7431, n11476);
  and g16031 (n11483, n10200, n_7431);
  not g16032 (n_7432, n11482);
  and g16033 (po0231, n_7432, n11483);
  and g16034 (n11485, pi0074, n11293);
  and g16035 (n11486, n2964, n7526);
  not g16036 (n_7433, n11486);
  and g16037 (n11487, n_135, n_7433);
  and g16038 (n11488, n_135, n_3206);
  and g16039 (n11489, n7417, n11488);
  and g16040 (n11490, n_135, n_3066);
  not g16041 (n_7434, n11490);
  and g16042 (n11491, pi0479, n_7434);
  not g16049 (n_7437, n11487);
  not g16052 (n_7438, n11485);
  not g16053 (n_7439, n11497);
  and g16054 (n11498, n_7438, n_7439);
  not g16055 (n_7440, n11498);
  and g16056 (po0232, n_4226, n_7440);
  and g16057 (n11500, n2620, n10195);
  not g16058 (n_7441, n11500);
  and g16059 (n11501, pi0075, n_7441);
  and g16060 (n11502, pi0096, n_3206);
  and g16061 (n11503, n2931, n_7437);
  not g16062 (n_7442, n11502);
  not g16063 (n_7443, n11503);
  and g16064 (n11504, n_7442, n_7443);
  not g16065 (n_7444, n11504);
  and g16066 (n11505, n2610, n_7444);
  and g16067 (n11506, n7534, n11505);
  not g16068 (n_7445, n11506);
  and g16069 (n11507, n_171, n_7445);
  not g16070 (n_7446, n11501);
  and g16071 (n11508, n8881, n_7446);
  not g16072 (n_7447, n11507);
  and g16073 (po0233, n_7447, n11508);
  and g16074 (n11510, n8930, n10186);
  not g16075 (n_7448, n10111);
  and g16076 (n11511, n_7448, n11510);
  not g16077 (n_7449, n11511);
  and g16078 (n11512, po1057, n_7449);
  and g16079 (n11513, n2519, n10375);
  and g16080 (n11514, pi0252, n2933);
  not g16081 (n_7450, n11514);
  and g16082 (n11515, n11513, n_7450);
  and g16083 (n11516, n_186, n11515);
  and g16084 (n11517, n_186, n2924);
  not g16085 (n_7451, n8931);
  and g16086 (n11518, n_125, n_7451);
  not g16087 (n_7452, n8897);
  and g16088 (n11519, n_7452, n_7209);
  not g16089 (n_7453, n11518);
  and g16090 (n11520, n10162, n_7453);
  not g16091 (n_7454, n11519);
  and g16092 (n11521, n_7454, n11520);
  not g16093 (n_7455, n2933);
  not g16094 (n_7456, n11521);
  and g16095 (n11522, n_7455, n_7456);
  and g16096 (n11523, n_280, n11521);
  and g16097 (n11524, pi0252, n11510);
  not g16098 (n_7457, n11524);
  and g16099 (n11525, n2933, n_7457);
  not g16100 (n_7458, n11523);
  and g16101 (n11526, n_7458, n11525);
  not g16102 (n_7459, n11522);
  not g16103 (n_7460, n11526);
  and g16104 (n11527, n_7459, n_7460);
  not g16105 (n_7461, n11527);
  and g16106 (n11528, pi0122, n_7461);
  and g16107 (n11529, n7417, n11522);
  not g16108 (n_7462, n6277);
  not g16109 (n_7463, n11513);
  and g16110 (n11530, n_7462, n_7463);
  not g16111 (n_7464, n11530);
  and g16112 (n11531, n_7460, n_7464);
  not g16113 (n_7465, n11529);
  and g16114 (n11532, n_7465, n11531);
  not g16115 (n_7466, n11532);
  and g16116 (n11533, n_4081, n_7466);
  not g16117 (n_7467, n11528);
  not g16118 (n_7468, n11533);
  and g16119 (n11534, n_7467, n_7468);
  not g16120 (n_7469, n11534);
  and g16121 (n11535, n_3206, n_7469);
  not g16122 (n_7470, n11515);
  and g16123 (n11536, n_4081, n_7470);
  not g16124 (n_7471, n11536);
  and g16125 (n11537, n_7467, n_7471);
  not g16126 (n_7472, n11537);
  and g16127 (n11538, pi1093, n_7472);
  not g16128 (n_7473, n11535);
  not g16129 (n_7474, n11538);
  and g16130 (n11539, n_7473, n_7474);
  not g16131 (n_7475, n11539);
  and g16132 (n11540, n2924, n_7475);
  not g16133 (n_7476, n11517);
  not g16134 (n_7477, n11540);
  and g16135 (n11541, n_7476, n_7477);
  not g16136 (n_7478, n11516);
  not g16137 (n_7479, n11541);
  and g16138 (n11542, n_7478, n_7479);
  and g16139 (n11543, n_4081, n11513);
  and g16140 (n11544, pi1093, n_7456);
  not g16141 (n_7480, n7418);
  not g16142 (n_7481, n11544);
  and g16143 (n11545, n_7480, n_7481);
  not g16144 (n_7482, n11543);
  not g16145 (n_7483, n11545);
  and g16146 (n11546, n_7482, n_7483);
  not g16147 (n_7484, n11546);
  and g16148 (n11547, n_7473, n_7484);
  not g16149 (n_7485, n11547);
  and g16150 (n11548, n_538, n_7485);
  and g16151 (n11549, n_186, n_538);
  not g16152 (n_7486, n11548);
  not g16153 (n_7487, n11549);
  and g16154 (n11550, n_7486, n_7487);
  and g16155 (n11551, pi0252, pi1092);
  and g16156 (n11552, n_3206, n11551);
  and g16157 (n11553, n2925, n11552);
  not g16158 (n_7488, n11553);
  and g16159 (n11554, n_186, n_7488);
  and g16160 (n11555, n11513, n11554);
  not g16161 (n_7489, n11550);
  not g16162 (n_7490, n11555);
  and g16163 (n11556, n_7489, n_7490);
  not g16164 (n_7491, n11542);
  not g16165 (n_7492, n11556);
  and g16166 (n11557, n_7491, n_7492);
  not g16167 (n_7493, n11557);
  and g16168 (n11558, n_5630, n_7493);
  and g16169 (n11559, n_186, po1057);
  not g16170 (n_7494, n11512);
  not g16171 (n_7495, n11559);
  and g16172 (n11560, n_7494, n_7495);
  not g16173 (n_7496, n11558);
  and g16174 (n11561, n_7496, n11560);
  not g16175 (n_7497, n11561);
  and g16176 (n11562, n_271, n_7497);
  and g16177 (n11563, n_7477, n_7486);
  not g16178 (n_7498, n11563);
  and g16179 (n11564, n_5630, n_7498);
  not g16180 (n_7499, n11564);
  and g16181 (n11565, n_7494, n_7499);
  not g16182 (n_7500, n11565);
  and g16183 (n11566, pi0210, n_7500);
  not g16184 (n_7501, n11562);
  not g16185 (n_7502, n11566);
  and g16186 (n11567, n_7501, n_7502);
  and g16187 (n11568, n2638, n10299);
  not g16188 (n_7503, n11567);
  not g16189 (n_7504, n11568);
  and g16190 (n11569, n_7503, n_7504);
  and g16191 (n11570, n_271, n_7493);
  and g16192 (n11571, pi0210, n_7498);
  not g16193 (n_7505, n11570);
  not g16194 (n_7506, n11571);
  and g16195 (n11572, n_7505, n_7506);
  not g16196 (n_7507, n11572);
  and g16197 (n11573, n11568, n_7507);
  not g16198 (n_7508, n11573);
  and g16199 (n11574, pi0299, n_7508);
  not g16200 (n_7509, n11569);
  and g16201 (n11575, n_7509, n11574);
  and g16202 (n11576, n_305, n_7497);
  and g16203 (n11577, pi0198, n_7500);
  not g16204 (n_7510, n11576);
  not g16205 (n_7511, n11577);
  and g16206 (n11578, n_7510, n_7511);
  and g16207 (n11579, n2669, n6197);
  not g16208 (n_7512, n11578);
  not g16209 (n_7513, n11579);
  and g16210 (n11580, n_7512, n_7513);
  and g16211 (n11581, pi0198, n_7498);
  and g16212 (n11582, n_305, n_7493);
  not g16213 (n_7514, n11581);
  not g16214 (n_7515, n11582);
  and g16215 (n11583, n_7514, n_7515);
  not g16216 (n_7516, n11583);
  and g16217 (n11584, n11579, n_7516);
  not g16218 (n_7517, n11584);
  and g16219 (n11585, n_234, n_7517);
  not g16220 (n_7518, n11580);
  and g16221 (n11586, n_7518, n11585);
  not g16222 (n_7519, n11575);
  not g16223 (n_7520, n11586);
  and g16224 (n11587, n_7519, n_7520);
  not g16225 (n_7521, n11587);
  and g16226 (n11588, pi0232, n_7521);
  and g16227 (n11589, pi0299, n_7503);
  and g16228 (n11590, n_234, n_7512);
  not g16229 (n_7522, n11589);
  and g16230 (n11591, n_3410, n_7522);
  not g16231 (n_7523, n11590);
  and g16232 (n11592, n_7523, n11591);
  not g16233 (n_7524, n11588);
  not g16234 (n_7525, n11592);
  and g16235 (n11593, n_7524, n_7525);
  not g16236 (n_7526, n11593);
  and g16237 (n11594, n7425, n_7526);
  and g16238 (n11595, n_538, n11544);
  and g16239 (n11596, n2933, n_7463);
  and g16240 (n11597, n_7450, n_7459);
  not g16241 (n_7527, n11596);
  and g16242 (n11598, n_7527, n11597);
  not g16243 (n_7528, n11598);
  and g16244 (n11599, n7418, n_7528);
  not g16245 (n_7529, n11599);
  and g16246 (n11600, n_7467, n_7529);
  not g16247 (n_7530, n11600);
  and g16248 (n11601, n2924, n_7530);
  and g16249 (n11602, n_3206, n_7461);
  not g16250 (n_7531, n11595);
  not g16251 (n_7532, n11602);
  and g16252 (n11603, n_7531, n_7532);
  not g16253 (n_7533, n11601);
  and g16254 (n11604, n_7533, n11603);
  and g16255 (n11605, n_5630, n11604);
  and g16256 (n11606, po1057, n11510);
  not g16257 (n_7534, n10108);
  and g16258 (n11607, n_7534, n11606);
  not g16259 (n_7535, n11605);
  not g16260 (n_7536, n11607);
  and g16261 (n11608, n_7535, n_7536);
  not g16262 (n_7537, n11608);
  and g16263 (n11609, pi0210, n_7537);
  and g16264 (n11610, n8904, n11559);
  and g16265 (n11611, pi0137, n11602);
  and g16266 (n11612, n_186, n_7528);
  and g16267 (n11613, n_3206, n11612);
  not g16268 (n_7538, n11611);
  and g16269 (n11614, n_7481, n_7538);
  not g16270 (n_7539, n11613);
  and g16271 (n11615, n_7539, n11614);
  and g16272 (n11616, n_5630, n11615);
  not g16273 (n_7540, n11606);
  not g16274 (n_7541, n11616);
  and g16275 (n11617, n_7540, n_7541);
  not g16276 (n_7542, n11610);
  and g16277 (n11618, n_538, n_7542);
  not g16278 (n_7543, n11617);
  and g16279 (n11619, n_7543, n11618);
  and g16280 (n11620, pi0137, n_7480);
  not g16281 (n_7544, n11620);
  and g16282 (n11621, n2933, n_7544);
  not g16283 (n_7545, n11621);
  and g16284 (n11622, n11510, n_7545);
  not g16285 (n_7546, n11622);
  and g16286 (n11623, po1057, n_7546);
  and g16287 (n11624, pi0137, n_7530);
  not g16288 (n_7547, n11612);
  and g16289 (n11625, n_7538, n_7547);
  not g16290 (n_7548, n11624);
  and g16291 (n11626, n_7548, n11625);
  not g16292 (n_7549, n11626);
  and g16293 (n11627, n_5630, n_7549);
  not g16294 (n_7550, n11623);
  and g16295 (n11628, n2924, n_7550);
  not g16296 (n_7551, n11627);
  and g16297 (n11629, n_7551, n11628);
  not g16298 (n_7552, n11619);
  not g16299 (n_7553, n11629);
  and g16300 (n11630, n_7552, n_7553);
  not g16301 (n_7554, n11630);
  and g16302 (n11631, n_271, n_7554);
  not g16303 (n_7555, n11609);
  not g16304 (n_7556, n11631);
  and g16305 (n11632, n_7555, n_7556);
  not g16306 (n_7557, n11632);
  and g16307 (n11633, n_7504, n_7557);
  and g16308 (n11634, n_538, n11615);
  and g16309 (n11635, n2924, n11626);
  not g16310 (n_7558, n11634);
  not g16311 (n_7559, n11635);
  and g16312 (n11636, n_7558, n_7559);
  and g16313 (n11637, n_271, n11636);
  not g16314 (n_7560, n11604);
  and g16315 (n11638, pi0210, n_7560);
  not g16316 (n_7561, n11638);
  and g16317 (n11639, n11568, n_7561);
  not g16318 (n_7562, n11637);
  and g16319 (n11640, n_7562, n11639);
  not g16320 (n_7563, n11640);
  and g16321 (n11641, pi0299, n_7563);
  not g16322 (n_7564, n11633);
  and g16323 (n11642, n_7564, n11641);
  and g16324 (n11643, pi0198, n_7537);
  and g16325 (n11644, n_305, n_7554);
  not g16326 (n_7565, n11643);
  not g16327 (n_7566, n11644);
  and g16328 (n11645, n_7565, n_7566);
  not g16329 (n_7567, n11645);
  and g16330 (n11646, n_7513, n_7567);
  not g16331 (n_7568, n11636);
  and g16332 (n11647, n_305, n_7568);
  and g16333 (n11648, pi0198, n11604);
  not g16334 (n_7569, n11647);
  not g16335 (n_7570, n11648);
  and g16336 (n11649, n_7569, n_7570);
  not g16337 (n_7571, n11649);
  and g16338 (n11650, n11579, n_7571);
  not g16339 (n_7572, n11650);
  and g16340 (n11651, n_234, n_7572);
  not g16341 (n_7573, n11646);
  and g16342 (n11652, n_7573, n11651);
  not g16343 (n_7574, n11642);
  not g16344 (n_7575, n11652);
  and g16345 (n11653, n_7574, n_7575);
  not g16346 (n_7576, n11653);
  and g16347 (n11654, pi0232, n_7576);
  and g16348 (n11655, n_234, n_7567);
  and g16349 (n11656, pi0299, n_7557);
  not g16350 (n_7577, n11655);
  and g16351 (n11657, n_3410, n_7577);
  not g16352 (n_7578, n11656);
  and g16353 (n11658, n_7578, n11657);
  not g16354 (n_7579, n11658);
  and g16355 (n11659, n_4091, n_7579);
  not g16356 (n_7580, n11654);
  and g16357 (n11660, n_7580, n11659);
  not g16358 (n_7581, n11594);
  not g16359 (n_7582, n11660);
  and g16360 (n11661, n_7581, n_7582);
  not g16361 (n_7583, n11661);
  and g16362 (po0234, n10165, n_7583);
  and g16363 (n11663, pi0086, n8897);
  and g16364 (n11664, n2778, n11663);
  not g16365 (n_7584, n11664);
  and g16366 (n11665, pi0314, n_7584);
  and g16367 (n11666, n2769, n2784);
  not g16368 (n_7585, n11666);
  and g16369 (n11667, n_119, n_7585);
  not g16370 (n_7586, n11667);
  and g16371 (n11668, n6452, n_7586);
  and g16372 (n11669, n2702, n11668);
  not g16373 (n_7587, n11669);
  and g16374 (n11670, n_3310, n_7587);
  not g16375 (n_7588, n11665);
  and g16376 (n11671, n10166, n_7588);
  not g16377 (n_7589, n11670);
  and g16378 (po0235, n_7589, n11671);
  and g16379 (n11673, pi0119, pi0232);
  and g16380 (po0236, n_3100, n11673);
  and g16381 (n11675, pi0163, n_6229);
  not g16382 (n_7591, pi0163);
  and g16383 (n11676, n_7591, n_6227);
  and g16384 (n11677, n_6226, n11676);
  not g16385 (n_7592, n11675);
  not g16386 (n_7593, n11677);
  and g16387 (n11678, n_7592, n_7593);
  and g16388 (n11679, pi0232, n11678);
  and g16389 (n11680, n_6232, n11679);
  not g16390 (n_7594, n11680);
  and g16391 (n11681, pi0074, n_7594);
  not g16392 (n_7595, n11679);
  and g16393 (n11682, pi0075, n_7595);
  and g16394 (n11683, pi0100, n_7595);
  not g16395 (n_7596, n11682);
  not g16396 (n_7597, n11683);
  and g16397 (n11684, n_7596, n_7597);
  and g16398 (n11685, pi0147, n7473);
  and g16399 (n11686, n8989, n11685);
  not g16400 (n_7599, n11686);
  and g16401 (n11687, n11684, n_7599);
  not g16402 (n_7600, n11681);
  and g16403 (n11688, n_824, n_7600);
  and g16404 (n11689, n11687, n11688);
  not g16405 (n_7601, n11687);
  and g16406 (n11690, pi0054, n_7601);
  and g16407 (n11691, n_161, n_143);
  not g16408 (n_7602, n11685);
  and g16409 (n11692, pi0038, n_7602);
  not g16410 (n_7603, n11692);
  and g16411 (n11693, n_164, n_7603);
  not g16412 (n_7604, n11691);
  and g16413 (n11694, n_7604, n11693);
  not g16414 (n_7605, n11694);
  and g16415 (n11695, n_7597, n_7605);
  not g16416 (n_7606, n11695);
  and g16417 (n11696, n_171, n_7606);
  not g16418 (n_7607, n11696);
  and g16419 (n11697, n_7596, n_7607);
  not g16420 (n_7608, n11697);
  and g16421 (n11698, n_167, n_7608);
  not g16422 (n_7609, n11690);
  not g16423 (n_7610, n11698);
  and g16424 (n11699, n_7609, n_7610);
  not g16425 (n_7611, n11699);
  and g16426 (n11700, n_168, n_7611);
  not g16427 (n_7612, n11700);
  and g16428 (n11701, n_7600, n_7612);
  not g16429 (n_7613, n11701);
  and g16430 (n11702, n_3243, n_7613);
  not g16431 (n_7614, n11702);
  and g16432 (n11703, n3328, n_7614);
  not g16433 (n_7615, n9722);
  and g16434 (n11704, n_7615, n9724);
  not g16435 (n_7617, pi0184);
  and g16436 (n11705, n_7617, n11704);
  and g16437 (n11706, pi0184, n6197);
  not g16438 (n_7618, n11704);
  and g16439 (n11707, n_7618, n11706);
  not g16440 (n_7619, n11705);
  and g16441 (n11708, n_234, n_7619);
  not g16442 (n_7620, n11707);
  and g16443 (n11709, n_7620, n11708);
  not g16444 (n_7621, n11678);
  and g16445 (n11710, pi0299, n_7621);
  not g16446 (n_7622, n11709);
  and g16447 (n11711, pi0232, n_7622);
  not g16448 (n_7623, n11710);
  and g16449 (n11712, n_7623, n11711);
  and g16450 (n11713, n_6232, n11712);
  not g16451 (n_7624, n11713);
  and g16452 (n11714, pi0074, n_7624);
  not g16453 (n_7625, n11714);
  and g16454 (n11715, n_176, n_7625);
  not g16455 (n_7627, pi0187);
  and g16456 (n11716, n_7627, n_234);
  not g16457 (n_7628, pi0147);
  and g16458 (n11717, n_7628, pi0299);
  not g16459 (n_7629, n11716);
  not g16460 (n_7630, n11717);
  and g16461 (n11718, n_7629, n_7630);
  and g16462 (n11719, n7473, n11718);
  not g16463 (n_7631, n11719);
  and g16464 (n11720, n8989, n_7631);
  not g16465 (n_7632, n11720);
  and g16466 (n11721, pi0054, n_7632);
  and g16467 (n11722, n_7624, n11721);
  not g16468 (n_7633, n11712);
  and g16469 (n11723, pi0075, n_7633);
  and g16470 (n11724, pi0100, n_7633);
  and g16471 (n11725, pi0038, n_7631);
  not g16472 (n_7634, n11725);
  and g16473 (n11726, n_164, n_7634);
  not g16474 (n_7636, pi0179);
  and g16475 (n11727, n_7636, n_234);
  not g16476 (n_7638, pi0156);
  and g16477 (n11728, n_7638, pi0299);
  not g16478 (n_7639, n11727);
  not g16479 (n_7640, n11728);
  and g16480 (n11729, n_7639, n_7640);
  and g16481 (n11730, n7473, n11729);
  not g16485 (n_7641, n11733);
  and g16486 (n11734, n11691, n_7641);
  not g16487 (n_7642, n11734);
  and g16488 (n11735, n11726, n_7642);
  not g16489 (n_7643, n11724);
  not g16490 (n_7644, n11735);
  and g16491 (n11736, n_7643, n_7644);
  not g16492 (n_7645, n11736);
  and g16493 (n11737, n9205, n_7645);
  and g16494 (n11738, n_7627, n_5815);
  and g16495 (n11739, pi0187, n_5817);
  not g16496 (n_7646, n11739);
  and g16497 (n11740, pi0147, n_7646);
  not g16498 (n_7647, n11738);
  and g16499 (n11741, n_7647, n11740);
  and g16500 (n11742, n_7628, pi0187);
  and g16501 (n11743, n9194, n11742);
  not g16502 (n_7648, n11741);
  not g16503 (n_7649, n11743);
  and g16504 (n11744, n_7648, n_7649);
  not g16505 (n_7650, n11744);
  and g16506 (n11745, pi0038, n_7650);
  and g16507 (n11746, n2509, n9093);
  and g16508 (n11747, n_3162, n9036);
  and g16509 (n11748, pi0156, n6188);
  and g16510 (n11749, n_266, n9293);
  not g16511 (n_7651, n11748);
  not g16512 (n_7652, n11749);
  and g16513 (n11750, n_7651, n_7652);
  not g16514 (n_7653, n11750);
  and g16515 (n11751, n11747, n_7653);
  and g16516 (n11752, n11746, n11751);
  and g16517 (n11753, n_143, pi0299);
  not g16518 (n_7654, n11752);
  and g16519 (n11754, n_7654, n11753);
  and g16520 (n11755, n_301, n9293);
  and g16521 (n11756, pi0179, n6188);
  not g16522 (n_7655, n11755);
  not g16523 (n_7656, n11756);
  and g16524 (n11757, n_7655, n_7656);
  and g16529 (n11761, n_143, n_234);
  not g16530 (n_7658, n11760);
  and g16531 (n11762, n_7658, n11761);
  not g16532 (n_7659, n11754);
  and g16533 (n11763, pi0039, n_7659);
  not g16534 (n_7660, n11762);
  and g16535 (n11764, n_7660, n11763);
  not g16536 (n_7662, pi0175);
  and g16537 (n11765, n_7662, n_234);
  and g16538 (n11766, pi0184, n9147);
  not g16539 (n_7663, n9143);
  and g16540 (n11767, n_7617, n_7663);
  not g16541 (n_7664, n11767);
  and g16542 (n11768, n_301, n_7664);
  not g16543 (n_7665, n11766);
  and g16544 (n11769, n_7665, n11768);
  and g16545 (n11770, n_142, pi0095);
  and g16546 (n11771, n_15, n11770);
  and g16547 (n11772, n2509, n11771);
  and g16548 (n11773, pi0182, n11772);
  and g16549 (n11774, pi0184, pi0189);
  not g16550 (n_7666, n9150);
  and g16551 (n11775, n_7666, n11774);
  not g16552 (n_7667, n11773);
  not g16553 (n_7668, n11775);
  and g16554 (n11776, n_7667, n_7668);
  not g16555 (n_7669, n11769);
  and g16556 (n11777, n_7669, n11776);
  not g16557 (n_7670, n11777);
  and g16558 (n11778, n6197, n_7670);
  not g16559 (n_7671, n11778);
  and g16560 (n11779, n_143, n_7671);
  not g16561 (n_7672, n11779);
  and g16562 (n11780, n11765, n_7672);
  and g16563 (n11781, n6197, n11772);
  and g16564 (n11782, pi0153, n9093);
  and g16565 (n11783, n9133, n11782);
  and g16566 (n11784, n9143, n10299);
  not g16572 (n_7675, n11781);
  and g16573 (n11788, n_7675, n11787);
  and g16574 (n11789, pi0040, n_3102);
  and g16575 (n11790, pi0166, n6197);
  not g16576 (n_7676, n11772);
  and g16577 (n11791, n_143, n_7676);
  and g16578 (n11792, n9166, n11791);
  not g16579 (n_7677, n11792);
  and g16580 (n11793, n11790, n_7677);
  and g16581 (n11794, n9162, n11791);
  not g16582 (n_7678, n11794);
  and g16583 (n11795, n10299, n_7678);
  not g16584 (n_7679, n11793);
  and g16585 (n11796, n_187, n_7679);
  not g16586 (n_7680, n11795);
  and g16587 (n11797, n_7680, n11796);
  and g16588 (n11798, n_271, n_5770);
  and g16589 (n11799, n_5771, n11791);
  not g16590 (n_7681, n11798);
  and g16591 (n11800, n_7681, n11799);
  not g16592 (n_7682, n11800);
  and g16593 (n11801, n10299, n_7682);
  and g16594 (n11802, n_5778, n11792);
  not g16595 (n_7683, n11802);
  and g16596 (n11803, n11790, n_7683);
  not g16597 (n_7684, n11803);
  and g16598 (n11804, pi0153, n_7684);
  not g16599 (n_7685, n11801);
  and g16600 (n11805, n_7685, n11804);
  not g16601 (n_7686, n11797);
  not g16602 (n_7687, n11805);
  and g16603 (n11806, n_7686, n_7687);
  not g16604 (n_7688, n11789);
  and g16605 (n11807, pi0163, n_7688);
  not g16606 (n_7689, n11806);
  and g16607 (n11808, n_7689, n11807);
  not g16608 (n_7690, n11808);
  and g16609 (n11809, pi0160, n_7690);
  and g16610 (n11810, pi0153, n9118);
  not g16611 (n_7691, n11810);
  and g16612 (n11811, n9162, n_7691);
  not g16613 (n_7692, n11811);
  and g16614 (n11812, n10299, n_7692);
  and g16615 (n11813, pi0153, n9129);
  not g16616 (n_7693, n11813);
  and g16617 (n11814, n9166, n_7693);
  not g16618 (n_7694, n11814);
  and g16619 (n11815, n11790, n_7694);
  not g16625 (n_7697, pi0160);
  not g16626 (n_7698, n11787);
  and g16627 (n11819, n_7697, n_7698);
  not g16628 (n_7699, n11818);
  and g16629 (n11820, n_7699, n11819);
  not g16630 (n_7700, n11809);
  not g16631 (n_7701, n11820);
  and g16632 (n11821, n_7700, n_7701);
  not g16633 (n_7702, n11788);
  and g16634 (n11822, pi0299, n_7702);
  not g16635 (n_7703, n11821);
  and g16636 (n11823, n_7703, n11822);
  and g16637 (n11824, n_5772, n11799);
  not g16638 (n_7704, n11824);
  and g16639 (n11825, n10295, n_7704);
  and g16640 (n11826, pi0189, n6197);
  and g16641 (n11827, n9130, n11791);
  not g16642 (n_7705, n11827);
  and g16643 (n11828, n11826, n_7705);
  and g16650 (n11833, pi0175, n_234);
  not g16651 (n_7708, n9133);
  and g16652 (n11834, pi0189, n_7708);
  not g16653 (n_7709, n9092);
  and g16654 (n11835, n_301, n_7709);
  not g16655 (n_7710, n11834);
  and g16656 (n11836, n2518, n_7710);
  not g16657 (n_7711, n11835);
  and g16658 (n11837, n_7711, n11836);
  not g16659 (n_7712, n11837);
  and g16660 (n11838, n_7667, n_7712);
  not g16661 (n_7713, n11838);
  and g16662 (n11839, n6197, n_7713);
  not g16663 (n_7714, n11839);
  and g16664 (n11840, n_7617, n_7714);
  and g16665 (n11841, pi0189, n9131);
  and g16666 (n11842, n_5773, n10295);
  not g16667 (n_7715, pi0182);
  not g16673 (n_7718, n11840);
  not g16674 (n_7719, n11845);
  and g16675 (n11846, n_7718, n_7719);
  not g16676 (n_7720, n11846);
  and g16677 (n11847, n_143, n_7720);
  not g16678 (n_7721, n11832);
  and g16679 (n11848, n_7721, n11833);
  not g16680 (n_7722, n11847);
  and g16681 (n11849, n_7722, n11848);
  not g16682 (n_7723, n11780);
  not g16683 (n_7724, n11849);
  and g16684 (n11850, n_7723, n_7724);
  not g16685 (n_7725, n11823);
  and g16686 (n11851, n_7725, n11850);
  not g16687 (n_7726, n11851);
  and g16688 (n11852, n_162, n_7726);
  not g16689 (n_7727, n11764);
  and g16690 (n11853, pi0232, n_7727);
  not g16691 (n_7728, n11852);
  and g16692 (n11854, n_7728, n11853);
  and g16693 (n11855, n_143, n_3410);
  not g16694 (n_7729, n11855);
  and g16695 (n11856, n_161, n_7729);
  not g16696 (n_7730, n11854);
  and g16697 (n11857, n_7730, n11856);
  not g16698 (n_7731, n11745);
  not g16699 (n_7732, n11857);
  and g16700 (n11858, n_7731, n_7732);
  not g16701 (n_7733, n11858);
  and g16702 (n11859, n2568, n_7733);
  and g16703 (n11860, pi0087, n_7604);
  and g16704 (n11861, n11726, n11860);
  not g16705 (n_7734, n11861);
  and g16706 (n11862, n_7643, n_7734);
  not g16707 (n_7735, n11859);
  and g16708 (n11863, n_7735, n11862);
  not g16709 (n_7736, n11863);
  and g16710 (n11864, n2569, n_7736);
  not g16711 (n_7737, n11723);
  not g16712 (n_7738, n11737);
  and g16713 (n11865, n_7737, n_7738);
  not g16714 (n_7739, n11864);
  and g16715 (n11866, n_7739, n11865);
  not g16716 (n_7740, n11866);
  and g16717 (n11867, n_167, n_7740);
  not g16718 (n_7741, n11722);
  not g16719 (n_7742, n11867);
  and g16720 (n11868, n_7741, n_7742);
  not g16721 (n_7743, n11868);
  and g16722 (n11869, n_168, n_7743);
  not g16723 (n_7744, n11869);
  and g16724 (n11870, n11715, n_7744);
  and g16725 (n11871, pi0055, n_7600);
  and g16726 (n11872, pi0163, pi0232);
  not g16730 (n_7745, n11875);
  and g16731 (n11876, n11691, n_7745);
  and g16732 (n11877, n_171, n11693);
  not g16733 (n_7746, n11876);
  and g16734 (n11878, n_7746, n11877);
  not g16735 (n_7747, n11878);
  and g16736 (n11879, n11684, n_7747);
  not g16737 (n_7748, n11879);
  and g16738 (n11880, n_167, n_7748);
  not g16739 (n_7749, n11880);
  and g16740 (n11881, n_7609, n_7749);
  not g16741 (n_7750, n11881);
  and g16742 (n11882, n_168, n_7750);
  not g16743 (n_7751, n11882);
  and g16744 (n11883, n11871, n_7751);
  not g16745 (n_7752, n11883);
  and g16746 (n11884, n2529, n_7752);
  not g16747 (n_7753, n11870);
  and g16748 (n11885, n_7753, n11884);
  not g16749 (n_7754, n11885);
  and g16750 (n11886, n11703, n_7754);
  not g16751 (n_7755, n11689);
  not g16752 (n_7756, n11886);
  and g16753 (n11887, n_7755, n_7756);
  and g16754 (n11888, pi0079, n11887);
  not g16755 (n_7757, n9260);
  and g16756 (n11889, n2487, n_7757);
  not g16757 (n_7758, n11889);
  and g16758 (n11890, n_143, n_7758);
  and g16759 (n11891, n_3102, n9260);
  not g16760 (n_7759, n11891);
  and g16761 (n11892, n9248, n_7759);
  and g16762 (n11893, n11872, n11892);
  not g16763 (n_7760, n11893);
  and g16764 (n11894, n11890, n_7760);
  not g16765 (n_7761, n11894);
  and g16766 (n11895, n_162, n_7761);
  and g16767 (n11896, pi0039, n_6031);
  not g16768 (n_7762, n11896);
  and g16769 (n11897, n9208, n_7762);
  not g16770 (n_7763, n11895);
  and g16771 (n11898, n_7763, n11897);
  and g16772 (n11899, pi0087, n_3321);
  and g16773 (n11900, n11691, n11899);
  not g16774 (n_7764, n11900);
  and g16775 (n11901, n11693, n_7764);
  not g16776 (n_7765, n11898);
  and g16777 (n11902, n_7765, n11901);
  not g16778 (n_7766, n11902);
  and g16779 (n11903, n_7597, n_7766);
  not g16780 (n_7767, n11903);
  and g16781 (n11904, n2569, n_7767);
  and g16782 (n11905, n_5880, n11695);
  not g16783 (n_7768, n11905);
  and g16784 (n11906, n9205, n_7768);
  not g16785 (n_7769, n11906);
  and g16786 (n11907, n_7596, n_7769);
  not g16787 (n_7770, n11904);
  and g16788 (n11908, n_7770, n11907);
  not g16789 (n_7771, n11908);
  and g16790 (n11909, n_167, n_7771);
  not g16791 (n_7772, n11909);
  and g16792 (n11910, n_7609, n_7772);
  not g16793 (n_7773, n11910);
  and g16794 (n11911, n_168, n_7773);
  not g16795 (n_7774, n11911);
  and g16796 (n11912, n11871, n_7774);
  and g16797 (n11913, n11726, n_7764);
  and g16798 (n11914, n2487, n11730);
  not g16799 (n_7775, n11914);
  and g16800 (n11915, n11890, n_7775);
  not g16801 (n_7776, n11915);
  and g16802 (n11916, n_162, n_7776);
  not g16803 (n_7777, n11916);
  and g16804 (n11917, n11897, n_7777);
  not g16805 (n_7778, n11917);
  and g16806 (n11918, n11913, n_7778);
  not g16807 (n_7779, n11918);
  and g16808 (n11919, n_7643, n_7779);
  not g16809 (n_7780, n11919);
  and g16810 (n11920, n9205, n_7780);
  and g16811 (n11921, pi0087, n11913);
  and g16812 (n11922, n_143, n_5892);
  not g16813 (n_7781, n11922);
  and g16814 (n11923, n6242, n_7781);
  and g16815 (n11924, n6227, n9466);
  not g16816 (n_7782, n9295);
  and g16817 (n11925, n2487, n_7782);
  not g16818 (n_7783, n11925);
  and g16819 (n11926, n_143, n_7783);
  and g16820 (n11927, n_3140, n11926);
  not g16821 (n_7784, n11924);
  not g16822 (n_7785, n11927);
  and g16823 (n11928, n_7784, n_7785);
  and g16824 (n11929, n_3162, n11928);
  not g16825 (n_7786, n11923);
  not g16826 (n_7787, n11929);
  and g16827 (n11930, n_7786, n_7787);
  and g16828 (n11931, n9291, n11930);
  and g16829 (n11932, n6205, n_7781);
  and g16830 (n11933, n_3119, n11928);
  not g16831 (n_7788, n11932);
  not g16832 (n_7789, n11933);
  and g16833 (n11934, n_7788, n_7789);
  not g16834 (n_7790, n11934);
  and g16835 (n11935, n9051, n_7790);
  and g16836 (n11936, n_5891, n_6031);
  not g16837 (n_7791, n11936);
  and g16838 (n11937, n_234, n_7791);
  not g16839 (n_7792, n11935);
  and g16840 (n11938, n_7792, n11937);
  not g16841 (n_7793, n11931);
  and g16842 (n11939, n_3410, n_7793);
  not g16843 (n_7794, n11938);
  and g16844 (n11940, n_7794, n11939);
  and g16845 (n11941, n_301, n_7781);
  and g16846 (n11942, n2487, n_5904);
  not g16847 (n_7795, n11942);
  and g16848 (n11943, n9140, n_7795);
  and g16849 (n11944, n6198, n11926);
  not g16850 (n_7796, n11944);
  and g16851 (n11945, n_7784, n_7796);
  not g16852 (n_7797, n11943);
  and g16853 (n11946, n_7797, n11945);
  and g16854 (n11947, pi0189, n_3119);
  and g16855 (n11948, n11946, n11947);
  not g16856 (n_7798, n11941);
  not g16857 (n_7799, n11948);
  and g16858 (n11949, n_7798, n_7799);
  not g16859 (n_7800, n11949);
  and g16860 (n11950, pi0179, n_7800);
  not g16861 (n_7801, n11928);
  and g16862 (n11951, pi0189, n_7801);
  and g16863 (n11952, n9140, n9324);
  and g16864 (n11953, n_3321, n9140);
  not g16865 (n_7802, n11952);
  not g16866 (n_7803, n11953);
  and g16867 (n11954, n_7802, n_7803);
  and g16868 (n11955, n11945, n11954);
  not g16869 (n_7804, n11955);
  and g16870 (n11956, n_301, n_7804);
  not g16876 (n_7807, n11959);
  and g16877 (n11960, n_7788, n_7807);
  not g16878 (n_7808, n11950);
  and g16879 (n11961, n_7808, n11960);
  not g16880 (n_7809, n11961);
  and g16881 (n11962, n9051, n_7809);
  not g16882 (n_7810, n11962);
  and g16883 (n11963, n_7791, n_7810);
  not g16884 (n_7811, n11963);
  and g16885 (n11964, n_234, n_7811);
  and g16886 (n11965, n_5881, n9466);
  not g16887 (n_7812, n11965);
  and g16888 (n11966, pi0299, n_7812);
  and g16889 (n11967, n_266, n_3162);
  not g16890 (n_7813, n11930);
  not g16891 (n_7814, n11967);
  and g16892 (n11968, n_7813, n_7814);
  and g16893 (n11969, n11955, n11967);
  not g16894 (n_7815, n11969);
  and g16895 (n11970, n9036, n_7815);
  not g16896 (n_7816, n11968);
  and g16897 (n11971, n_7816, n11970);
  not g16898 (n_7817, n11971);
  and g16899 (n11972, n11966, n_7817);
  not g16900 (n_7818, n11964);
  not g16901 (n_7819, n11972);
  and g16902 (n11973, n_7818, n_7819);
  and g16903 (n11974, n_7638, pi0232);
  not g16904 (n_7820, n11973);
  and g16905 (n11975, n_7820, n11974);
  and g16906 (n11976, pi0166, n_3162);
  and g16907 (n11977, n11946, n11976);
  not g16908 (n_7821, n11976);
  and g16909 (n11978, n_7781, n_7821);
  not g16910 (n_7822, n11978);
  and g16911 (n11979, n9036, n_7822);
  not g16912 (n_7823, n11977);
  and g16913 (n11980, n_7823, n11979);
  not g16914 (n_7824, n11980);
  and g16915 (n11981, n11966, n_7824);
  not g16916 (n_7825, n11981);
  and g16917 (n11982, n_7818, n_7825);
  and g16918 (n11983, pi0156, pi0232);
  not g16919 (n_7826, n11982);
  and g16920 (n11984, n_7826, n11983);
  and g16927 (n11988, n_145, n_6051);
  not g16928 (n_7830, n9349);
  and g16929 (n11989, n9348, n_7830);
  not g16930 (n_7831, n11988);
  not g16931 (n_7832, n11989);
  and g16932 (n11990, n_7831, n_7832);
  not g16933 (n_7833, n9456);
  and g16934 (n11991, n_143, n_7833);
  not g16935 (n_7834, n11991);
  and g16936 (n11992, n_144, n_7834);
  not g16937 (n_7835, n11990);
  not g16938 (n_7836, n11992);
  and g16939 (n11993, n_7835, n_7836);
  and g16940 (n11994, n_234, n11993);
  and g16941 (n11995, n_143, n_6125);
  not g16942 (n_7837, n11995);
  and g16943 (n11996, n_144, n_7837);
  not g16944 (n_7838, n11996);
  and g16945 (n11997, n_7835, n_7838);
  and g16946 (n11998, pi0299, n11997);
  not g16947 (n_7839, n11994);
  and g16948 (n11999, n_3410, n_7839);
  not g16949 (n_7840, n11998);
  and g16950 (n12000, n_7840, n11999);
  and g16951 (n12001, n_3102, n11993);
  and g16952 (n12002, n_143, n_5996);
  not g16953 (n_7841, n12002);
  and g16954 (n12003, n_144, n_7841);
  and g16955 (n12004, n_143, n_6010);
  and g16956 (n12005, pi0189, n12004);
  not g16957 (n_7842, n12005);
  and g16958 (n12006, n12003, n_7842);
  and g16959 (n12007, n_7715, n11990);
  and g16960 (n12008, pi0182, n9485);
  not g16963 (n_7844, n12007);
  not g16967 (n_7846, n12011);
  and g16968 (n12012, pi0184, n_7846);
  and g16969 (n12013, n_143, n9403);
  not g16970 (n_7847, n12013);
  and g16971 (n12014, n_142, n_7847);
  not g16972 (n_7848, n12014);
  and g16973 (n12015, n_6049, n_7848);
  not g16974 (n_7849, n12015);
  and g16975 (n12016, n_144, n_7849);
  not g16976 (n_7850, n12016);
  and g16977 (n12017, n_6051, n_7850);
  not g16978 (n_7851, n12017);
  and g16979 (n12018, n_305, n_7851);
  and g16980 (n12019, n_6041, n_7848);
  not g16981 (n_7852, n12019);
  and g16982 (n12020, n_144, n_7852);
  not g16983 (n_7853, n12020);
  and g16984 (n12021, n_6051, n_7853);
  not g16985 (n_7854, n12021);
  and g16986 (n12022, pi0198, n_7854);
  not g16987 (n_7855, n12018);
  and g16988 (n12023, n10295, n_7855);
  not g16989 (n_7856, n12022);
  and g16990 (n12024, n_7856, n12023);
  and g16991 (n12025, n11826, n11991);
  not g16997 (n_7859, n12012);
  not g16998 (n_7860, n12028);
  and g16999 (n12029, n_7859, n_7860);
  not g17000 (n_7861, n12029);
  and g17001 (n12030, n11765, n_7861);
  and g17002 (n12031, pi0095, n_7715);
  and g17003 (n12032, n_143, n_6062);
  and g17004 (n12033, n_144, pi0189);
  not g17005 (n_7862, n12033);
  and g17006 (n12034, n2487, n_7862);
  not g17007 (n_7863, n12034);
  and g17008 (n12035, n12032, n_7863);
  not g17009 (n_7864, n12031);
  not g17010 (n_7865, n12035);
  and g17011 (n12036, n_7864, n_7865);
  not g17012 (n_7866, n12036);
  and g17013 (n12037, n11706, n_7866);
  and g17014 (n12038, n_7844, n12037);
  and g17015 (n12039, n9560, n10295);
  and g17016 (n12040, n_305, n_6053);
  and g17017 (n12041, n_144, n_6044);
  not g17018 (n_7867, n12041);
  and g17019 (n12042, n_6051, n_7867);
  not g17020 (n_7868, n12042);
  and g17021 (n12043, pi0198, n_7868);
  not g17022 (n_7869, n12040);
  and g17023 (n12044, n11826, n_7869);
  not g17024 (n_7870, n12043);
  and g17025 (n12045, n_7870, n12044);
  not g17026 (n_7871, n12039);
  and g17027 (n12046, pi0182, n_7871);
  not g17028 (n_7872, n12045);
  and g17029 (n12047, n_7872, n12046);
  and g17030 (n12048, n_6052, n_7835);
  not g17031 (n_7873, n12048);
  and g17032 (n12049, n_305, n_7873);
  and g17033 (n12050, n_7835, n_7867);
  not g17034 (n_7874, n12050);
  and g17035 (n12051, pi0198, n_7874);
  not g17036 (n_7875, n12049);
  and g17037 (n12052, n11826, n_7875);
  not g17038 (n_7876, n12051);
  and g17039 (n12053, n_7876, n12052);
  not g17040 (n_7877, n12053);
  and g17041 (n12054, n_7715, n_7877);
  not g17042 (n_7878, n12047);
  not g17043 (n_7879, n12054);
  and g17044 (n12055, n_7878, n_7879);
  and g17045 (n12056, n_6107, n_7864);
  and g17046 (n12057, n10295, n_7835);
  not g17047 (n_7880, n12056);
  and g17048 (n12058, n_7880, n12057);
  not g17049 (n_7881, n12055);
  not g17050 (n_7882, n12058);
  and g17051 (n12059, n_7881, n_7882);
  not g17052 (n_7883, n12059);
  and g17053 (n12060, n_7617, n_7883);
  not g17054 (n_7884, n12038);
  and g17055 (n12061, n11833, n_7884);
  not g17056 (n_7885, n12060);
  and g17057 (n12062, n_7885, n12061);
  not g17058 (n_7886, n12030);
  not g17059 (n_7887, n12062);
  and g17060 (n12063, n_7886, n_7887);
  not g17061 (n_7888, n12001);
  not g17062 (n_7889, n12063);
  and g17063 (n12064, n_7888, n_7889);
  and g17064 (n12065, n_3102, n11997);
  not g17065 (n_7890, n12032);
  and g17066 (n12066, n_144, n_7890);
  not g17067 (n_7891, n12066);
  and g17068 (n12067, pi0166, n_7891);
  not g17069 (n_7892, n11474);
  and g17070 (n12068, n_7892, n_7891);
  not g17071 (n_7893, n12067);
  and g17072 (n12069, pi0153, n_7893);
  not g17073 (n_7894, n12068);
  and g17074 (n12070, n_7894, n12069);
  and g17075 (n12071, pi0166, n12004);
  not g17076 (n_7895, n12071);
  and g17077 (n12072, n12003, n_7895);
  and g17078 (n12073, n_187, n12072);
  and g17085 (n12078, n6197, n_6051);
  and g17086 (n12079, n12067, n12078);
  and g17087 (n12080, n9466, n10299);
  not g17088 (n_7898, n12080);
  and g17089 (n12081, pi0153, n_7898);
  not g17090 (n_7899, n12079);
  and g17091 (n12082, n_7899, n12081);
  not g17092 (n_7900, n12072);
  and g17093 (n12083, n_7900, n12078);
  not g17094 (n_7901, n12083);
  and g17095 (n12084, n_187, n_7901);
  not g17096 (n_7902, n12082);
  and g17097 (n12085, pi0160, n_7902);
  not g17098 (n_7903, n12084);
  and g17099 (n12086, n_7903, n12085);
  not g17100 (n_7904, n12077);
  and g17101 (n12087, pi0163, n_7904);
  not g17102 (n_7905, n12086);
  and g17103 (n12088, n_7905, n12087);
  and g17104 (n12089, pi0210, n_7874);
  and g17105 (n12090, n_271, n_7873);
  not g17106 (n_7906, n12089);
  and g17107 (n12091, n11790, n_7906);
  not g17108 (n_7907, n12090);
  and g17109 (n12092, n_7907, n12091);
  and g17110 (n12093, n_6103, n_7835);
  not g17111 (n_7908, n12093);
  and g17112 (n12094, n_271, n_7908);
  and g17113 (n12095, n_6100, n_7835);
  not g17114 (n_7909, n12095);
  and g17115 (n12096, pi0210, n_7909);
  not g17116 (n_7910, n12094);
  and g17117 (n12097, n10299, n_7910);
  not g17118 (n_7911, n12096);
  and g17119 (n12098, n_7911, n12097);
  not g17120 (n_7912, n12092);
  and g17121 (n12099, pi0153, n_7912);
  not g17122 (n_7913, n12098);
  and g17123 (n12100, n_7913, n12099);
  and g17124 (n12101, pi0166, n11997);
  and g17125 (n12102, n_7835, n_7853);
  not g17126 (n_7914, n12102);
  and g17127 (n12103, pi0210, n_7914);
  and g17128 (n12104, n_7835, n_7850);
  not g17129 (n_7915, n12104);
  and g17130 (n12105, n_271, n_7915);
  not g17131 (n_7916, n12103);
  and g17132 (n12106, n10299, n_7916);
  not g17133 (n_7917, n12105);
  and g17134 (n12107, n_7917, n12106);
  not g17135 (n_7918, n12107);
  and g17136 (n12108, n_187, n_7918);
  not g17137 (n_7919, n12101);
  and g17138 (n12109, n_7919, n12108);
  not g17139 (n_7920, n12100);
  and g17140 (n12110, n_7697, n_7920);
  not g17141 (n_7921, n12109);
  and g17142 (n12111, n_7921, n12110);
  and g17143 (n12112, pi0210, n_6101);
  and g17144 (n12113, n_271, n_6104);
  not g17145 (n_7922, n12112);
  and g17146 (n12114, n10299, n_7922);
  not g17147 (n_7923, n12113);
  and g17148 (n12115, n_7923, n12114);
  and g17149 (n12116, n_271, n_6053);
  and g17150 (n12117, pi0210, n_7868);
  not g17151 (n_7924, n12116);
  and g17152 (n12118, n11790, n_7924);
  not g17153 (n_7925, n12117);
  and g17154 (n12119, n_7925, n12118);
  not g17155 (n_7926, n12115);
  and g17156 (n12120, pi0153, n_7926);
  not g17157 (n_7927, n12119);
  and g17158 (n12121, n_7927, n12120);
  and g17159 (n12122, n11790, n11995);
  and g17160 (n12123, n_271, n_7851);
  and g17161 (n12124, pi0210, n_7854);
  not g17162 (n_7928, n12123);
  and g17163 (n12125, n10299, n_7928);
  not g17164 (n_7929, n12124);
  and g17165 (n12126, n_7929, n12125);
  not g17166 (n_7930, n12126);
  and g17167 (n12127, n_187, n_7930);
  not g17168 (n_7931, n12122);
  and g17169 (n12128, n_7931, n12127);
  not g17170 (n_7932, n12121);
  and g17171 (n12129, pi0160, n_7932);
  not g17172 (n_7933, n12128);
  and g17173 (n12130, n_7933, n12129);
  not g17174 (n_7934, n12130);
  and g17175 (n12131, n_7591, n_7934);
  not g17176 (n_7935, n12111);
  and g17177 (n12132, n_7935, n12131);
  not g17178 (n_7936, n12088);
  not g17179 (n_7937, n12132);
  and g17180 (n12133, n_7936, n_7937);
  not g17181 (n_7938, n12065);
  and g17182 (n12134, pi0299, n_7938);
  not g17183 (n_7939, n12133);
  and g17184 (n12135, n_7939, n12134);
  and g17185 (n12136, n_6812, n11993);
  and g17186 (n12137, pi0198, n_7914);
  and g17187 (n12138, n_305, n_7915);
  not g17188 (n_7940, n12137);
  and g17189 (n12139, n10295, n_7940);
  not g17190 (n_7941, n12138);
  and g17191 (n12140, n_7941, n12139);
  not g17198 (n_7944, n12064);
  not g17199 (n_7945, n12144);
  and g17200 (n12145, n_7944, n_7945);
  not g17201 (n_7946, n12135);
  and g17202 (n12146, n_7946, n12145);
  not g17203 (n_7947, n12146);
  and g17204 (n12147, pi0232, n_7947);
  not g17205 (n_7948, n12000);
  and g17206 (n12148, n_162, n_7948);
  not g17207 (n_7949, n12147);
  and g17208 (n12149, n_7949, n12148);
  not g17209 (n_7950, n11987);
  and g17210 (n12150, n_161, n_7950);
  not g17211 (n_7951, n12149);
  and g17212 (n12151, n_7951, n12150);
  not g17213 (n_7952, n12151);
  and g17214 (n12152, n_7731, n_7952);
  not g17215 (n_7953, n12152);
  and g17216 (n12153, n2568, n_7953);
  not g17217 (n_7954, n11921);
  and g17218 (n12154, n_7643, n_7954);
  not g17219 (n_7955, n12153);
  and g17220 (n12155, n_7955, n12154);
  not g17221 (n_7956, n12155);
  and g17222 (n12156, n2569, n_7956);
  not g17223 (n_7957, n11920);
  and g17224 (n12157, n_7737, n_7957);
  not g17225 (n_7958, n12156);
  and g17226 (n12158, n_7958, n12157);
  not g17227 (n_7959, n12158);
  and g17228 (n12159, n_167, n_7959);
  not g17229 (n_7960, n12159);
  and g17230 (n12160, n_7741, n_7960);
  not g17231 (n_7961, n12160);
  and g17232 (n12161, n_168, n_7961);
  not g17233 (n_7962, n12161);
  and g17234 (n12162, n11715, n_7962);
  not g17235 (n_7963, n11912);
  and g17236 (n12163, n2529, n_7963);
  not g17237 (n_7964, n12162);
  and g17238 (n12164, n_7964, n12163);
  and g17239 (n12165, n_6208, n11703);
  not g17240 (n_7965, n12164);
  and g17241 (n12166, n_7965, n12165);
  not g17242 (n_7966, n12166);
  and g17243 (n12167, n_7755, n_7966);
  and g17244 (n12168, n_5677, n12167);
  and g17245 (n12169, n_5679, n10058);
  not g17246 (n_7967, n11888);
  not g17247 (n_7968, n12169);
  and g17248 (n12170, n_7967, n_7968);
  not g17249 (n_7969, n12168);
  and g17250 (n12171, n_7969, n12170);
  not g17251 (n_7970, n8977);
  and g17252 (n12172, n_5677, n_7970);
  and g17253 (n12173, n11887, n12172);
  not g17254 (n_7971, n12172);
  and g17255 (n12174, n12167, n_7971);
  not g17256 (n_7972, n12173);
  and g17257 (n12175, n12169, n_7972);
  not g17258 (n_7973, n12174);
  and g17259 (n12176, n_7973, n12175);
  or g17260 (po0237, n12171, n12176);
  and g17261 (n12178, pi0098, pi1092);
  and g17262 (n12179, pi1093, n12178);
  and g17263 (n12180, n_4112, n2926);
  not g17264 (n_7974, n12179);
  not g17265 (n_7975, n12180);
  and g17266 (n12181, n_7974, n_7975);
  not g17267 (n_7977, pi0080);
  not g17268 (n_7978, n12181);
  and g17269 (n12182, n_7977, n_7978);
  not g17270 (n_7979, n12182);
  and g17271 (n12183, pi0217, n_7979);
  and g17272 (n12184, n7425, n12181);
  and g17273 (n12185, n_4834, n12181);
  not g17274 (n_7980, n12185);
  and g17275 (n12186, pi0588, n_7980);
  and g17276 (n12187, pi0592, n_5023);
  not g17277 (n_7981, n8119);
  and g17278 (n12188, n7422, n_7981);
  not g17279 (n_7982, n12187);
  and g17280 (n12189, n_7982, n12188);
  not g17281 (n_7983, n12189);
  and g17282 (n12190, n12181, n_7983);
  not g17283 (n_7984, n12190);
  and g17284 (n12191, n_4718, n_7984);
  and g17285 (n12192, pi0428, n_7984);
  and g17286 (n12193, n_4419, n12181);
  not g17287 (n_7985, n12193);
  and g17288 (n12194, n_4976, n_7985);
  not g17289 (n_7986, n12192);
  not g17290 (n_7987, n12194);
  and g17291 (n12195, n_7986, n_7987);
  not g17292 (n_7988, n12195);
  and g17293 (n12196, n_4974, n_7988);
  and g17294 (n12197, n_4976, n_7984);
  and g17295 (n12198, pi0428, n_7985);
  not g17296 (n_7989, n12197);
  not g17297 (n_7990, n12198);
  and g17298 (n12199, n_7989, n_7990);
  not g17299 (n_7991, n12199);
  and g17300 (n12200, pi0427, n_7991);
  not g17301 (n_7992, n12196);
  not g17302 (n_7993, n12200);
  and g17303 (n12201, n_7992, n_7993);
  not g17304 (n_7994, n12201);
  and g17305 (n12202, n_4981, n_7994);
  and g17306 (n12203, n_4974, n_7991);
  and g17307 (n12204, pi0427, n_7988);
  not g17308 (n_7995, n12203);
  not g17309 (n_7996, n12204);
  and g17310 (n12205, n_7995, n_7996);
  not g17311 (n_7997, n12205);
  and g17312 (n12206, pi0430, n_7997);
  not g17313 (n_7998, n12202);
  not g17314 (n_7999, n12206);
  and g17315 (n12207, n_7998, n_7999);
  not g17316 (n_8000, n12207);
  and g17317 (n12208, n_4985, n_8000);
  and g17318 (n12209, n_4981, n_7997);
  and g17319 (n12210, pi0430, n_7994);
  not g17320 (n_8001, n12209);
  not g17321 (n_8002, n12210);
  and g17322 (n12211, n_8001, n_8002);
  not g17323 (n_8003, n12211);
  and g17324 (n12212, pi0426, n_8003);
  not g17325 (n_8004, n12208);
  not g17326 (n_8005, n12212);
  and g17327 (n12213, n_8004, n_8005);
  not g17328 (n_8006, n12213);
  and g17329 (n12214, n_4990, n_8006);
  and g17330 (n12215, n_4985, n_8003);
  and g17331 (n12216, pi0426, n_8000);
  not g17332 (n_8007, n12215);
  not g17333 (n_8008, n12216);
  and g17334 (n12217, n_8007, n_8008);
  not g17335 (n_8009, n12217);
  and g17336 (n12218, pi0445, n_8009);
  not g17337 (n_8010, n12214);
  not g17338 (n_8011, n12218);
  and g17339 (n12219, n_8010, n_8011);
  not g17340 (n_8012, n12219);
  and g17341 (n12220, pi0448, n_8012);
  and g17342 (n12221, n_4990, n_8009);
  and g17343 (n12222, pi0445, n_8006);
  not g17344 (n_8013, n12221);
  not g17345 (n_8014, n12222);
  and g17346 (n12223, n_8013, n_8014);
  not g17347 (n_8015, n12223);
  and g17348 (n12224, n_4995, n_8015);
  not g17349 (n_8016, n12220);
  and g17350 (n12225, n8128, n_8016);
  not g17351 (n_8017, n12224);
  and g17352 (n12226, n_8017, n12225);
  and g17353 (n12227, n_4995, n_8012);
  and g17354 (n12228, pi0448, n_8015);
  not g17355 (n_8018, n12227);
  and g17356 (n12229, n_5003, n_8018);
  not g17357 (n_8019, n12228);
  and g17358 (n12230, n_8019, n12229);
  not g17359 (n_8020, n12226);
  and g17360 (n12231, pi1199, n_8020);
  not g17361 (n_8021, n12230);
  and g17362 (n12232, n_8021, n12231);
  not g17363 (n_8022, n12191);
  and g17364 (n12233, n8041, n_8022);
  not g17365 (n_8023, n12232);
  and g17366 (n12234, n_8023, n12233);
  not g17367 (n_8024, n12234);
  and g17368 (n12235, n12186, n_8024);
  and g17369 (n12236, pi0591, n_7978);
  not g17370 (n_8025, n12236);
  and g17371 (n12237, pi0590, n_8025);
  and g17372 (n12238, n_4571, n12181);
  and g17373 (n12239, n7854, n12238);
  and g17374 (n12240, n_4569, n12239);
  not g17375 (n_8026, n12240);
  and g17376 (n12241, n_7985, n_8026);
  not g17377 (n_8027, n12241);
  and g17378 (n12242, pi0461, n_8027);
  and g17379 (n12243, n_4578, n12239);
  not g17380 (n_8028, n12243);
  and g17381 (n12244, n_7985, n_8028);
  not g17382 (n_8029, n12244);
  and g17383 (n12245, n_4575, n_8029);
  not g17384 (n_8030, n12242);
  not g17385 (n_8031, n12245);
  and g17386 (n12246, n_8030, n_8031);
  not g17387 (n_8032, n12246);
  and g17388 (n12247, pi0357, n_8032);
  and g17389 (n12248, pi0461, n_8029);
  and g17390 (n12249, n_4575, n_8027);
  not g17391 (n_8033, n12248);
  not g17392 (n_8034, n12249);
  and g17393 (n12250, n_8033, n_8034);
  not g17394 (n_8035, n12250);
  and g17395 (n12251, n_4585, n_8035);
  not g17396 (n_8036, n12247);
  not g17397 (n_8037, n12251);
  and g17398 (n12252, n_8036, n_8037);
  not g17399 (n_8038, n12252);
  and g17400 (n12253, pi0356, n_8038);
  and g17401 (n12254, pi0357, n_8035);
  and g17402 (n12255, n_4585, n_8032);
  not g17403 (n_8039, n12254);
  not g17404 (n_8040, n12255);
  and g17405 (n12256, n_8039, n_8040);
  not g17406 (n_8041, n12256);
  and g17407 (n12257, n_4593, n_8041);
  not g17408 (n_8042, n12253);
  not g17409 (n_8043, n12257);
  and g17410 (n12258, n_8042, n_8043);
  and g17411 (n12259, pi0354, n12258);
  and g17412 (n12260, pi0356, n_8041);
  and g17413 (n12261, n_4593, n_8038);
  not g17414 (n_8044, n12260);
  not g17415 (n_8045, n12261);
  and g17416 (n12262, n_8044, n_8045);
  and g17417 (n12263, n_4616, n12262);
  not g17418 (n_8046, n12259);
  and g17419 (n12264, n_4615, n_8046);
  not g17420 (n_8047, n12263);
  and g17421 (n12265, n_8047, n12264);
  and g17422 (n12266, pi0354, n12262);
  and g17423 (n12267, n_4616, n12258);
  not g17424 (n_8048, n12266);
  and g17425 (n12268, n7887, n_8048);
  not g17426 (n_8049, n12267);
  and g17427 (n12269, n_8049, n12268);
  not g17428 (n_8050, n12265);
  and g17429 (n12270, n_4628, n_8050);
  not g17430 (n_8051, n12269);
  and g17431 (n12271, n_8051, n12270);
  not g17432 (n_8052, n12271);
  and g17433 (n12272, n12237, n_8052);
  and g17434 (n12273, n_4723, n_5238);
  not g17435 (n_8053, n12273);
  and g17436 (n12274, n_7985, n_8053);
  and g17437 (n12275, pi0592, n_7978);
  and g17438 (n12276, n_5024, n_7978);
  not g17439 (n_8054, n12275);
  not g17440 (n_8055, n12276);
  and g17441 (n12277, n_8054, n_8055);
  and g17442 (n12278, pi0397, n_4686);
  and g17443 (n12279, n_4682, pi0404);
  not g17444 (n_8056, n12278);
  not g17445 (n_8057, n12279);
  and g17446 (n12280, n_8056, n_8057);
  not g17447 (n_8058, n12280);
  and g17448 (n12281, pi0411, n_8058);
  and g17449 (n12282, n_4710, n12280);
  not g17450 (n_8059, n12281);
  not g17451 (n_8060, n12282);
  and g17452 (n12283, n_8059, n_8060);
  and g17453 (n12284, n_4705, n12283);
  not g17454 (n_8061, n12283);
  and g17455 (n12285, n7932, n_8061);
  not g17456 (n_8062, n12284);
  not g17457 (n_8063, n12285);
  and g17458 (n12286, n_8062, n_8063);
  not g17459 (n_8064, n12286);
  and g17460 (n12287, n7417, n_8064);
  not g17461 (n_8065, n12178);
  not g17462 (n_8066, n12287);
  and g17463 (n12288, n_8065, n_8066);
  not g17464 (n_8067, n12288);
  and g17465 (n12289, n_4681, n_8067);
  and g17466 (n12290, n7417, n12286);
  not g17467 (n_8068, n12290);
  and g17468 (n12291, n_8065, n_8068);
  not g17469 (n_8069, n12291);
  and g17470 (n12292, pi0412, n_8069);
  not g17471 (n_8070, n12289);
  and g17472 (n12293, n7944, n_8070);
  not g17473 (n_8071, n12292);
  and g17474 (n12294, n_8071, n12293);
  and g17475 (n12295, pi0412, n_8067);
  and g17476 (n12296, n_4681, n_8069);
  not g17477 (n_8072, n12295);
  and g17478 (n12297, n_4701, n_8072);
  not g17479 (n_8073, n12296);
  and g17480 (n12298, n_8073, n12297);
  not g17481 (n_8074, n12294);
  and g17482 (n12299, n_4081, n_8074);
  not g17483 (n_8075, n12298);
  and g17484 (n12300, n_8075, n12299);
  not g17485 (n_8076, n12300);
  and g17486 (n12301, n_8065, n_8076);
  not g17487 (n_8077, n12301);
  and g17488 (n12302, n7626, n_8077);
  and g17489 (n12303, pi1091, n12179);
  not g17490 (n_8078, n12302);
  not g17491 (n_8079, n12303);
  and g17492 (n12304, n_8078, n_8079);
  not g17493 (n_8080, n12304);
  and g17494 (n12305, pi0567, n_8080);
  not g17495 (n_8081, n12305);
  and g17496 (n12306, n_7975, n_8081);
  not g17497 (n_8082, n12306);
  and g17498 (n12307, n7958, n_8082);
  not g17499 (n_8083, n12307);
  and g17500 (n12308, n12277, n_8083);
  not g17501 (n_8084, n12308);
  and g17502 (n12309, n_4718, n_8084);
  and g17503 (n12310, n_4081, n7417);
  not g17504 (n_8085, n12310);
  and g17505 (n12311, n_8065, n_8085);
  and g17506 (n12312, n_4214, n_8079);
  and g17507 (n12313, n7417, n7926);
  and g17508 (n12314, n_4081, n_8065);
  not g17509 (n_8086, n12313);
  and g17510 (n12315, n_8086, n12314);
  not g17511 (n_8087, n12312);
  not g17512 (n_8088, n12315);
  and g17513 (n12316, n_8087, n_8088);
  not g17514 (n_8089, n12311);
  and g17515 (n12317, n_8089, n12316);
  and g17516 (n12318, pi0567, n12317);
  not g17517 (n_8090, n12318);
  and g17518 (n12319, n_7975, n_8090);
  and g17519 (n12320, n_8081, n12319);
  not g17520 (n_8091, n12320);
  and g17521 (n12321, n7958, n_8091);
  not g17522 (n_8092, n12319);
  and g17523 (n12322, n8668, n_8092);
  not g17524 (n_8093, n12322);
  and g17525 (n12323, n_8054, n_8093);
  not g17526 (n_8094, n12321);
  and g17527 (n12324, n_8094, n12323);
  not g17528 (n_8095, n12324);
  and g17529 (n12325, pi1199, n_8095);
  not g17530 (n_8096, n12309);
  not g17531 (n_8097, n12325);
  and g17532 (n12326, n_8096, n_8097);
  not g17533 (n_8098, n12326);
  and g17534 (n12327, n12273, n_8098);
  not g17535 (n_8099, n12274);
  not g17536 (n_8100, n12327);
  and g17537 (n12328, n_8099, n_8100);
  not g17538 (n_8101, n12328);
  and g17539 (n12329, pi0333, n_8101);
  and g17540 (n12330, n8395, n_7985);
  and g17541 (n12331, n_5238, n_8098);
  not g17542 (n_8102, n12330);
  not g17543 (n_8103, n12331);
  and g17544 (n12332, n_8102, n_8103);
  not g17545 (n_8104, n12332);
  and g17546 (n12333, n_4773, n_8104);
  not g17547 (n_8105, n12329);
  not g17548 (n_8106, n12333);
  and g17549 (n12334, n_8105, n_8106);
  not g17550 (n_8107, n12334);
  and g17551 (n12335, pi0391, n_8107);
  and g17552 (n12336, n_4773, n_8101);
  and g17553 (n12337, pi0333, n_8104);
  not g17554 (n_8108, n12336);
  not g17555 (n_8109, n12337);
  and g17556 (n12338, n_8108, n_8109);
  not g17557 (n_8110, n12338);
  and g17558 (n12339, n_4778, n_8110);
  and g17559 (n12340, pi0392, n8801);
  and g17560 (n12341, n_4785, n_5561);
  not g17561 (n_8111, n12340);
  not g17562 (n_8112, n12341);
  and g17563 (n12342, n_8111, n_8112);
  not g17564 (n_8113, n12335);
  not g17565 (n_8114, n12342);
  and g17566 (n12343, n_8113, n_8114);
  not g17567 (n_8115, n12339);
  and g17568 (n12344, n_8115, n12343);
  and g17569 (n12345, pi0391, n_8110);
  and g17570 (n12346, n_4778, n_8107);
  not g17571 (n_8116, n12345);
  and g17572 (n12347, n12342, n_8116);
  not g17573 (n_8117, n12346);
  and g17574 (n12348, n_8117, n12347);
  not g17575 (n_8118, n12344);
  and g17576 (n12349, pi0591, n_8118);
  not g17577 (n_8119, n12348);
  and g17578 (n12350, n_8119, n12349);
  and g17579 (n12351, n_4419, n_4424);
  not g17580 (n_8120, n7726);
  and g17581 (n12352, n7422, n_8120);
  not g17582 (n_8121, n12352);
  and g17583 (n12353, n_4377, n_8121);
  not g17584 (n_8122, n12353);
  and g17585 (n12354, n_4729, n_8122);
  not g17586 (n_8123, n12351);
  and g17587 (n12355, n_8123, n12354);
  not g17588 (n_8124, n12355);
  and g17589 (n12356, n12181, n_8124);
  not g17590 (n_8125, n12356);
  and g17591 (n12357, n_4628, n_8125);
  not g17592 (n_8126, n12357);
  and g17593 (n12358, n_4423, n_8126);
  not g17594 (n_8127, n12350);
  and g17595 (n12359, n_8127, n12358);
  not g17596 (n_8128, n12272);
  and g17597 (n12360, n_4832, n_8128);
  not g17598 (n_8129, n12359);
  and g17599 (n12361, n_8129, n12360);
  not g17600 (n_8130, n12235);
  and g17601 (n12362, n_4091, n_8130);
  not g17602 (n_8131, n12361);
  and g17603 (n12363, n_8131, n12362);
  and g17609 (n12367, pi0567, n7429);
  not g17610 (n_8134, n7420);
  and g17611 (n12368, n_8134, n_7974);
  and g17612 (n12369, n_4081, n12368);
  not g17613 (n_8135, n12369);
  and g17614 (n12370, n7626, n_8135);
  and g17615 (n12371, n2625, n_8079);
  not g17616 (n_8136, n12370);
  and g17617 (n12372, n_8136, n12371);
  and g17618 (n12373, pi0824, pi0950);
  and g17619 (n12374, n_113, n2701);
  and g17620 (n12375, n_46, n2495);
  and g17621 (n12376, n10379, n12375);
  and g17622 (n12377, n12374, n12376);
  and g17623 (n12378, n7440, n12377);
  and g17624 (n12379, n7446, n12378);
  and g17625 (n12380, pi0051, n12379);
  and g17626 (n12381, pi0090, pi0093);
  not g17633 (n_8139, n12380);
  not g17634 (n_8140, n12385);
  and g17635 (n12386, n_8139, n_8140);
  and g17636 (n12387, n7450, n12373);
  not g17637 (n_8141, n12386);
  and g17638 (n12388, n_8141, n12387);
  not g17639 (n_8142, n12388);
  and g17640 (n12389, n_47, n_8142);
  not g17641 (n_8143, n12389);
  and g17642 (n12390, pi1092, n_8143);
  and g17643 (n12391, n_172, n12371);
  not g17644 (n_8144, n12390);
  and g17645 (n12392, n_8144, n12391);
  and g17646 (n12393, n2520, n12373);
  and g17647 (n12394, n12379, n12393);
  not g17648 (n_8145, n12394);
  and g17649 (n12395, n_47, n_8145);
  not g17650 (n_8146, n12395);
  and g17651 (n12396, pi1092, n_8146);
  and g17652 (n12397, pi0087, n12371);
  not g17653 (n_8147, n12396);
  and g17654 (n12398, n_8147, n12397);
  not g17655 (n_8148, n12392);
  not g17656 (n_8149, n12398);
  and g17657 (n12399, n_8148, n_8149);
  not g17658 (n_8150, n12399);
  and g17659 (n12400, pi0122, n_8150);
  not g17660 (n_8151, n12372);
  not g17661 (n_8152, n12400);
  and g17662 (n12401, n_8151, n_8152);
  not g17663 (n_8153, n12401);
  and g17664 (n12402, n_171, n_8153);
  not g17665 (n_8154, n7465);
  and g17666 (n12403, n_8154, n12368);
  not g17667 (n_8155, n12403);
  and g17668 (n12404, n12367, n_8155);
  not g17669 (n_8156, n12402);
  and g17670 (n12405, n_8156, n12404);
  not g17671 (n_8157, n12368);
  and g17672 (n12406, n_4196, n_8157);
  not g17673 (n_8158, n12406);
  and g17674 (n12407, n_7975, n_8158);
  not g17675 (n_8159, n12405);
  and g17676 (n12408, n_8159, n12407);
  not g17677 (n_8160, n12408);
  and g17678 (n12409, n_4239, n_8160);
  not g17679 (n_8161, n12409);
  and g17680 (n12410, n_8054, n_8161);
  and g17681 (n12411, n_5023, n12410);
  and g17682 (n12412, n8093, n_8055);
  and g17683 (n12413, n_4947, n_7978);
  not g17684 (n_8162, n12410);
  and g17685 (n12414, pi0443, n_8162);
  not g17686 (n_8163, n12413);
  not g17687 (n_8164, n12414);
  and g17688 (n12415, n_8163, n_8164);
  and g17689 (n12416, n8249, n12415);
  and g17690 (n12417, pi0443, n_7978);
  and g17691 (n12418, n_4947, n_8162);
  not g17692 (n_8165, n12417);
  not g17693 (n_8166, n12418);
  and g17694 (n12419, n_8165, n_8166);
  and g17695 (n12420, n_5092, n12419);
  not g17696 (n_8167, n12416);
  not g17697 (n_8168, n12420);
  and g17698 (n12421, n_8167, n_8168);
  not g17699 (n_8169, n12421);
  and g17700 (n12422, pi0435, n_8169);
  and g17701 (n12423, n_4952, n12419);
  and g17702 (n12424, pi0444, n12415);
  not g17703 (n_8170, n12423);
  and g17704 (n12425, n_4948, n_8170);
  not g17705 (n_8171, n12424);
  and g17706 (n12426, n_8171, n12425);
  and g17707 (n12427, n_4952, n12415);
  and g17708 (n12428, pi0444, n12419);
  not g17709 (n_8172, n12427);
  and g17710 (n12429, pi0436, n_8172);
  not g17711 (n_8173, n12428);
  and g17712 (n12430, n_8173, n12429);
  not g17713 (n_8174, n12426);
  not g17714 (n_8175, n12430);
  and g17715 (n12431, n_8174, n_8175);
  and g17716 (n12432, n_4922, n12431);
  not g17717 (n_8176, n12422);
  not g17718 (n_8177, n12432);
  and g17719 (n12433, n_8176, n_8177);
  and g17720 (n12434, n_4921, n12433);
  and g17721 (n12435, n_4922, n_8169);
  and g17722 (n12436, pi0435, n12431);
  not g17723 (n_8178, n12435);
  not g17724 (n_8179, n12436);
  and g17725 (n12437, n_8178, n_8179);
  and g17726 (n12438, pi0429, n12437);
  not g17727 (n_8180, n12434);
  and g17728 (n12439, n8105, n_8180);
  not g17729 (n_8181, n12438);
  and g17730 (n12440, n_8181, n12439);
  and g17731 (n12441, n_4921, n12437);
  and g17732 (n12442, pi0429, n12433);
  not g17733 (n_8182, n12441);
  and g17734 (n12443, n_4942, n_8182);
  not g17735 (n_8183, n12442);
  and g17736 (n12444, n_8183, n12443);
  not g17737 (n_8184, n12440);
  and g17738 (n12445, pi1196, n_8184);
  not g17739 (n_8185, n12444);
  and g17740 (n12446, n_8185, n12445);
  not g17741 (n_8186, n12446);
  and g17742 (n12447, n12412, n_8186);
  not g17743 (n_8187, n12411);
  not g17744 (n_8188, n12447);
  and g17745 (n12448, n_8187, n_8188);
  and g17746 (n12449, n_4718, n12448);
  not g17747 (n_8189, n12448);
  and g17748 (n12450, pi0428, n_8189);
  and g17749 (n12451, n_4976, n12410);
  not g17750 (n_8190, n12450);
  not g17751 (n_8191, n12451);
  and g17752 (n12452, n_8190, n_8191);
  not g17753 (n_8192, n12452);
  and g17754 (n12453, n_4974, n_8192);
  and g17755 (n12454, n_4976, n_8189);
  and g17756 (n12455, pi0428, n12410);
  not g17757 (n_8193, n12454);
  not g17758 (n_8194, n12455);
  and g17759 (n12456, n_8193, n_8194);
  not g17760 (n_8195, n12456);
  and g17761 (n12457, pi0427, n_8195);
  not g17762 (n_8196, n12453);
  not g17763 (n_8197, n12457);
  and g17764 (n12458, n_8196, n_8197);
  not g17765 (n_8198, n12458);
  and g17766 (n12459, pi0430, n_8198);
  and g17767 (n12460, n_4974, n_8195);
  and g17768 (n12461, pi0427, n_8192);
  not g17769 (n_8199, n12460);
  not g17770 (n_8200, n12461);
  and g17771 (n12462, n_8199, n_8200);
  not g17772 (n_8201, n12462);
  and g17773 (n12463, n_4981, n_8201);
  not g17774 (n_8202, n12459);
  not g17775 (n_8203, n12463);
  and g17776 (n12464, n_8202, n_8203);
  not g17777 (n_8204, n12464);
  and g17778 (n12465, pi0426, n_8204);
  and g17779 (n12466, pi0430, n_8201);
  and g17780 (n12467, n_4981, n_8198);
  not g17781 (n_8205, n12466);
  not g17782 (n_8206, n12467);
  and g17783 (n12468, n_8205, n_8206);
  not g17784 (n_8207, n12468);
  and g17785 (n12469, n_4985, n_8207);
  not g17786 (n_8208, n12465);
  not g17787 (n_8209, n12469);
  and g17788 (n12470, n_8208, n_8209);
  not g17789 (n_8210, n12470);
  and g17790 (n12471, pi0445, n_8210);
  and g17791 (n12472, pi0426, n_8207);
  and g17792 (n12473, n_4985, n_8204);
  not g17793 (n_8211, n12472);
  not g17794 (n_8212, n12473);
  and g17795 (n12474, n_8211, n_8212);
  not g17796 (n_8213, n12474);
  and g17797 (n12475, n_4990, n_8213);
  not g17798 (n_8214, n12471);
  not g17799 (n_8215, n12475);
  and g17800 (n12476, n_8214, n_8215);
  and g17801 (n12477, pi0448, n12476);
  and g17802 (n12478, pi0445, n_8213);
  and g17803 (n12479, n_4990, n_8210);
  not g17804 (n_8216, n12478);
  not g17805 (n_8217, n12479);
  and g17806 (n12480, n_8216, n_8217);
  and g17807 (n12481, n_4995, n12480);
  not g17808 (n_8218, n12477);
  and g17809 (n12482, n_5003, n_8218);
  not g17810 (n_8219, n12481);
  and g17811 (n12483, n_8219, n12482);
  and g17812 (n12484, n_4995, n12476);
  and g17813 (n12485, pi0448, n12480);
  not g17814 (n_8220, n12484);
  and g17815 (n12486, n8128, n_8220);
  not g17816 (n_8221, n12485);
  and g17817 (n12487, n_8221, n12486);
  not g17818 (n_8222, n12483);
  and g17819 (n12488, pi1199, n_8222);
  not g17820 (n_8223, n12487);
  and g17821 (n12489, n_8223, n12488);
  not g17822 (n_8224, n12449);
  and g17823 (n12490, n8041, n_8224);
  not g17824 (n_8225, n12489);
  and g17825 (n12491, n_8225, n12490);
  not g17826 (n_8226, n12491);
  and g17827 (n12492, n12186, n_8226);
  and g17828 (n12493, n7850, n12181);
  not g17829 (n_8227, n7850);
  and g17830 (n12494, n_8227, n12410);
  not g17831 (n_8228, n12493);
  not g17832 (n_8229, n12494);
  and g17833 (n12495, n_8228, n_8229);
  not g17834 (n_8230, n12495);
  and g17835 (n12496, pi1198, n_8230);
  and g17836 (n12497, n_4377, n_8055);
  and g17837 (n12498, n7791, n12181);
  and g17838 (n12499, n_4486, n12410);
  not g17839 (n_8231, n12498);
  not g17840 (n_8232, n12499);
  and g17841 (n12500, n_8231, n_8232);
  not g17842 (n_8233, n12500);
  and g17843 (n12501, n_4485, n_8233);
  and g17844 (n12502, pi0455, n_7978);
  and g17845 (n12503, n_4480, n_8162);
  not g17846 (n_8234, n12502);
  not g17847 (n_8235, n12503);
  and g17848 (n12504, n_8234, n_8235);
  not g17849 (n_8236, n12504);
  and g17850 (n12505, n_4481, n_8236);
  and g17851 (n12506, n_4480, n_7978);
  and g17852 (n12507, pi0455, n_8162);
  not g17853 (n_8237, n12506);
  not g17854 (n_8238, n12507);
  and g17855 (n12508, n_8237, n_8238);
  not g17856 (n_8239, n12508);
  and g17857 (n12509, pi0452, n_8239);
  not g17858 (n_8240, n12505);
  not g17859 (n_8241, n12509);
  and g17860 (n12510, n_8240, n_8241);
  and g17861 (n12511, pi0355, n12510);
  not g17862 (n_8242, n12501);
  not g17863 (n_8243, n12511);
  and g17864 (n12512, n_8242, n_8243);
  and g17865 (n12513, n_4491, n12512);
  and g17866 (n12514, pi0355, n_8233);
  and g17867 (n12515, n_4485, n12510);
  not g17868 (n_8244, n12514);
  not g17869 (n_8245, n12515);
  and g17870 (n12516, n_8244, n_8245);
  and g17871 (n12517, pi0458, n12516);
  not g17872 (n_8246, n12513);
  and g17873 (n12518, n7812, n_8246);
  not g17874 (n_8247, n12517);
  and g17875 (n12519, n_8247, n12518);
  and g17876 (n12520, n_4491, n12516);
  and g17877 (n12521, pi0458, n12512);
  not g17878 (n_8248, n12520);
  and g17879 (n12522, n_4511, n_8248);
  not g17880 (n_8249, n12521);
  and g17881 (n12523, n_8249, n12522);
  not g17882 (n_8250, n12519);
  and g17883 (n12524, pi1196, n_8250);
  not g17884 (n_8251, n12523);
  and g17885 (n12525, n_8251, n12524);
  not g17886 (n_8252, n12525);
  and g17887 (n12526, n12497, n_8252);
  not g17888 (n_8253, n12496);
  not g17889 (n_8254, n12526);
  and g17890 (n12527, n_8253, n_8254);
  not g17891 (n_8255, n12527);
  and g17892 (n12528, n_4565, n_8255);
  and g17893 (n12529, n7782, n12410);
  not g17894 (n_8256, n12528);
  not g17895 (n_8257, n12529);
  and g17896 (n12530, n_8256, n_8257);
  and g17897 (n12531, n_4569, n12530);
  and g17898 (n12532, pi1199, n_8162);
  and g17899 (n12533, pi0351, n12532);
  not g17900 (n_8258, n12531);
  not g17901 (n_8259, n12533);
  and g17902 (n12534, n_8258, n_8259);
  not g17903 (n_8260, n12534);
  and g17904 (n12535, n_4575, n_8260);
  and g17905 (n12536, n_4578, n12530);
  and g17906 (n12537, n_4577, n12532);
  not g17907 (n_8261, n12536);
  not g17908 (n_8262, n12537);
  and g17909 (n12538, n_8261, n_8262);
  not g17910 (n_8263, n12538);
  and g17911 (n12539, pi0461, n_8263);
  not g17912 (n_8264, n12535);
  not g17913 (n_8265, n12539);
  and g17914 (n12540, n_8264, n_8265);
  not g17915 (n_8266, n12540);
  and g17916 (n12541, n_4585, n_8266);
  and g17917 (n12542, n_4575, n_8263);
  and g17918 (n12543, pi0461, n_8260);
  not g17919 (n_8267, n12542);
  not g17920 (n_8268, n12543);
  and g17921 (n12544, n_8267, n_8268);
  not g17922 (n_8269, n12544);
  and g17923 (n12545, pi0357, n_8269);
  not g17924 (n_8270, n12541);
  not g17925 (n_8271, n12545);
  and g17926 (n12546, n_8270, n_8271);
  not g17927 (n_8272, n12546);
  and g17928 (n12547, n_4593, n_8272);
  and g17929 (n12548, n_4585, n_8269);
  and g17930 (n12549, pi0357, n_8266);
  not g17931 (n_8273, n12548);
  not g17932 (n_8274, n12549);
  and g17933 (n12550, n_8273, n_8274);
  not g17934 (n_8275, n12550);
  and g17935 (n12551, pi0356, n_8275);
  not g17936 (n_8276, n12547);
  not g17937 (n_8277, n12551);
  and g17938 (n12552, n_8276, n_8277);
  not g17939 (n_8278, n12552);
  and g17940 (n12553, n_4616, n_8278);
  and g17941 (n12554, n_4593, n_8275);
  and g17942 (n12555, pi0356, n_8272);
  not g17943 (n_8279, n12554);
  not g17944 (n_8280, n12555);
  and g17945 (n12556, n_8279, n_8280);
  not g17946 (n_8281, n12556);
  and g17947 (n12557, pi0354, n_8281);
  not g17948 (n_8282, n12553);
  and g17949 (n12558, n_4615, n_8282);
  not g17950 (n_8283, n12557);
  and g17951 (n12559, n_8283, n12558);
  and g17952 (n12560, n_4616, n_8281);
  and g17953 (n12561, pi0354, n_8278);
  not g17954 (n_8284, n12560);
  and g17955 (n12562, n7887, n_8284);
  not g17956 (n_8285, n12561);
  and g17957 (n12563, n_8285, n12562);
  not g17958 (n_8286, n12559);
  and g17959 (n12564, n_4628, n_8286);
  not g17960 (n_8287, n12563);
  and g17961 (n12565, n_8287, n12564);
  not g17962 (n_8288, n12565);
  and g17963 (n12566, n12237, n_8288);
  and g17964 (n12567, n_8053, n12410);
  and g17965 (n12568, n7429, n_7975);
  not g17966 (n_8289, n12568);
  and g17967 (n12569, n_8082, n_8289);
  and g17968 (n12570, pi0075, n12304);
  and g17969 (n12571, n_4710, n12178);
  not g17970 (n_8290, n12571);
  and g17971 (n12572, n7950, n_8290);
  and g17972 (n12573, pi0411, n12396);
  not g17973 (n_8291, n12573);
  and g17974 (n12574, n12572, n_8291);
  and g17975 (n12575, n_4710, n12396);
  and g17976 (n12576, n_4711, n_8065);
  not g17977 (n_8292, n12576);
  and g17978 (n12577, n_4713, n_8292);
  not g17979 (n_8293, n12575);
  not g17980 (n_8294, n12577);
  and g17981 (n12578, n_8293, n_8294);
  not g17982 (n_8295, n12574);
  not g17983 (n_8296, n12578);
  and g17984 (n12579, n_8295, n_8296);
  and g17985 (n12580, pi0122, n12579);
  not g17986 (n_8297, n12580);
  and g17987 (n12581, n_8076, n_8297);
  not g17988 (n_8298, n12581);
  and g17989 (n12582, n7626, n_8298);
  not g17990 (n_8299, n12582);
  and g17991 (n12583, n12397, n_8299);
  and g17992 (n12584, pi0411, n12390);
  not g17993 (n_8300, n12584);
  and g17994 (n12585, n12572, n_8300);
  and g17995 (n12586, n_4710, n12390);
  not g17996 (n_8301, n12586);
  and g17997 (n12587, n_8294, n_8301);
  not g17998 (n_8302, n12585);
  not g17999 (n_8303, n12587);
  and g18000 (n12588, n_8302, n_8303);
  and g18001 (n12589, pi0122, n12588);
  not g18002 (n_8304, n12589);
  and g18003 (n12590, n_8076, n_8304);
  not g18004 (n_8305, n12590);
  and g18005 (n12591, n7626, n_8305);
  not g18006 (n_8306, n12591);
  and g18007 (n12592, n12391, n_8306);
  and g18008 (n12593, n_251, n12304);
  not g18009 (n_8307, n12583);
  not g18010 (n_8308, n12593);
  and g18011 (n12594, n_8307, n_8308);
  not g18012 (n_8309, n12592);
  and g18013 (n12595, n_8309, n12594);
  not g18014 (n_8310, n12595);
  and g18015 (n12596, n_171, n_8310);
  not g18016 (n_8311, n12570);
  and g18017 (n12597, n12367, n_8311);
  not g18018 (n_8312, n12596);
  and g18019 (n12598, n_8312, n12597);
  not g18020 (n_8313, n12569);
  not g18021 (n_8314, n12598);
  and g18022 (n12599, n_8313, n_8314);
  not g18023 (n_8315, n12599);
  and g18024 (n12600, n7958, n_8315);
  not g18025 (n_8316, n12600);
  and g18026 (n12601, n_8055, n_8316);
  not g18027 (n_8317, n12601);
  and g18028 (n12602, n_4718, n_8317);
  and g18029 (n12603, n_8091, n_8289);
  not g18030 (n_8318, n12317);
  and g18031 (n12604, n_8154, n_8318);
  and g18032 (n12605, n_8078, n12604);
  not g18033 (n_8319, n12316);
  and g18034 (n12606, n2625, n_8319);
  and g18035 (n12607, n_8078, n12606);
  and g18036 (n12608, n_4081, n12313);
  and g18037 (n12609, n7926, n12390);
  and g18038 (n12610, n_4672, n12178);
  not g18039 (n_8320, n12609);
  not g18040 (n_8321, n12610);
  and g18041 (n12611, n_8320, n_8321);
  and g18042 (n12612, n12391, n12611);
  and g18043 (n12613, n_4711, n_8301);
  not g18044 (n_8322, n12613);
  and g18045 (n12614, n_8302, n_8322);
  not g18046 (n_8323, n12614);
  and g18047 (n12615, n12612, n_8323);
  and g18048 (n12616, n7926, n12396);
  not g18049 (n_8324, n12616);
  and g18050 (n12617, n12397, n_8324);
  not g18051 (n_8325, n12579);
  and g18052 (n12618, n_8325, n12617);
  not g18053 (n_8326, n12615);
  not g18054 (n_8327, n12618);
  and g18055 (n12619, n_8326, n_8327);
  not g18056 (n_8328, n12608);
  and g18057 (n12620, n_8076, n_8328);
  not g18058 (n_8329, n12619);
  and g18059 (n12621, n_8329, n12620);
  not g18060 (n_8330, n12607);
  not g18061 (n_8331, n12621);
  and g18062 (n12622, n_8330, n_8331);
  not g18063 (n_8332, n12622);
  and g18064 (n12623, n_171, n_8332);
  not g18065 (n_8333, n12605);
  and g18066 (n12624, n12367, n_8333);
  not g18067 (n_8334, n12623);
  and g18068 (n12625, n_8334, n12624);
  not g18069 (n_8335, n12603);
  not g18070 (n_8336, n12625);
  and g18071 (n12626, n_8335, n_8336);
  not g18072 (n_8337, n12626);
  and g18073 (n12627, n7958, n_8337);
  and g18074 (n12628, n_8092, n_8289);
  and g18075 (n12629, n_8321, n_8324);
  and g18076 (n12630, n12397, n12629);
  not g18077 (n_8338, n12612);
  not g18078 (n_8339, n12630);
  and g18079 (n12631, n_8338, n_8339);
  not g18080 (n_8340, n12631);
  and g18081 (n12632, pi0122, n_8340);
  not g18082 (n_8341, n12606);
  not g18083 (n_8342, n12632);
  and g18084 (n12633, n_8341, n_8342);
  not g18085 (n_8343, n12633);
  and g18086 (n12634, n_171, n_8343);
  not g18087 (n_8344, n12604);
  and g18088 (n12635, n12367, n_8344);
  not g18089 (n_8345, n12634);
  and g18090 (n12636, n_8345, n12635);
  not g18091 (n_8346, n12628);
  not g18092 (n_8347, n12636);
  and g18093 (n12637, n_8346, n_8347);
  not g18094 (n_8348, n12637);
  and g18095 (n12638, n8668, n_8348);
  not g18096 (n_8349, n12627);
  not g18097 (n_8350, n12638);
  and g18098 (n12639, n_8349, n_8350);
  not g18099 (n_8351, n12639);
  and g18100 (n12640, pi1199, n_8351);
  not g18101 (n_8352, n12640);
  and g18102 (n12641, n_8054, n_8352);
  not g18103 (n_8353, n12602);
  and g18104 (n12642, n_8353, n12641);
  and g18105 (n12643, n12273, n12642);
  not g18106 (n_8354, n12567);
  not g18107 (n_8355, n12643);
  and g18108 (n12644, n_8354, n_8355);
  not g18109 (n_8356, n12644);
  and g18110 (n12645, pi0333, n_8356);
  and g18111 (n12646, n8395, n_8162);
  not g18112 (n_8357, n12642);
  and g18113 (n12647, n_5238, n_8357);
  not g18114 (n_8358, n12646);
  not g18115 (n_8359, n12647);
  and g18116 (n12648, n_8358, n_8359);
  and g18117 (n12649, n_4773, n12648);
  not g18118 (n_8360, n12645);
  not g18119 (n_8361, n12649);
  and g18120 (n12650, n_8360, n_8361);
  not g18121 (n_8362, n12650);
  and g18122 (n12651, pi0391, n_8362);
  not g18123 (n_8363, n12648);
  and g18124 (n12652, pi0333, n_8363);
  and g18125 (n12653, n_4773, n12644);
  not g18126 (n_8364, n12652);
  not g18127 (n_8365, n12653);
  and g18128 (n12654, n_8364, n_8365);
  and g18129 (n12655, n_4778, n12654);
  not g18130 (n_8366, n12651);
  not g18131 (n_8367, n12655);
  and g18132 (n12656, n_8366, n_8367);
  not g18133 (n_8368, n12656);
  and g18134 (n12657, pi0392, n_8368);
  and g18135 (n12658, n_4778, n12650);
  not g18136 (n_8369, n12654);
  and g18137 (n12659, pi0391, n_8369);
  not g18138 (n_8370, n12658);
  not g18139 (n_8371, n12659);
  and g18140 (n12660, n_8370, n_8371);
  and g18141 (n12661, n_4785, n12660);
  not g18142 (n_8372, n12657);
  not g18143 (n_8373, n12661);
  and g18144 (n12662, n_8372, n_8373);
  not g18145 (n_8374, n12662);
  and g18146 (n12663, pi0393, n_8374);
  and g18147 (n12664, n_4785, n_8368);
  and g18148 (n12665, pi0392, n12660);
  not g18149 (n_8375, n12664);
  not g18150 (n_8376, n12665);
  and g18151 (n12666, n_8375, n_8376);
  not g18152 (n_8377, n12666);
  and g18153 (n12667, n_4793, n_8377);
  not g18154 (n_8378, n12663);
  not g18155 (n_8379, n12667);
  and g18156 (n12668, n_8378, n_8379);
  not g18157 (n_8380, n12668);
  and g18158 (n12669, n_4821, n_8380);
  and g18159 (n12670, pi0393, n_8377);
  and g18160 (n12671, n_4793, n_8374);
  not g18161 (n_8381, n12670);
  not g18162 (n_8382, n12671);
  and g18163 (n12672, n_8381, n_8382);
  not g18164 (n_8383, n12672);
  and g18165 (n12673, n8028, n_8383);
  not g18166 (n_8384, n12669);
  and g18167 (n12674, pi0591, n_8384);
  not g18168 (n_8385, n12673);
  and g18169 (n12675, n_8385, n12674);
  and g18170 (n12676, n_4239, n_7978);
  and g18171 (n12677, pi0592, n_8160);
  not g18172 (n_8386, n12676);
  not g18173 (n_8387, n12677);
  and g18174 (n12678, n_8386, n_8387);
  and g18175 (n12679, n_4370, n12678);
  and g18176 (n12680, n7722, n12181);
  not g18177 (n_8388, n12679);
  not g18178 (n_8389, n12680);
  and g18179 (n12681, n_8388, n_8389);
  and g18180 (n12682, pi1199, n12681);
  and g18181 (n12683, n7670, n12678);
  and g18182 (n12684, n_4723, n_7978);
  not g18183 (n_8390, n12684);
  and g18184 (n12685, n_4325, n_8390);
  and g18185 (n12686, pi0367, n_7978);
  not g18186 (n_8391, n12678);
  and g18187 (n12687, n_4317, n_8391);
  not g18188 (n_8392, n12686);
  not g18189 (n_8393, n12687);
  and g18190 (n12688, n_8392, n_8393);
  not g18191 (n_8394, n12688);
  and g18192 (n12689, n7673, n_8394);
  and g18193 (n12690, n_4317, n_7978);
  and g18194 (n12691, pi0367, n_8391);
  not g18195 (n_8395, n12690);
  not g18196 (n_8396, n12691);
  and g18197 (n12692, n_8395, n_8396);
  not g18198 (n_8397, n12692);
  and g18199 (n12693, n_4320, n_8397);
  not g18200 (n_8398, n12689);
  not g18201 (n_8399, n12693);
  and g18202 (n12694, n_8398, n_8399);
  not g18203 (n_8400, n12694);
  and g18204 (n12695, n7676, n_8400);
  and g18205 (n12696, n_4320, n12688);
  and g18206 (n12697, n7673, n12692);
  not g18207 (n_8401, n12696);
  not g18208 (n_8402, n12697);
  and g18209 (n12698, n_8401, n_8402);
  and g18210 (n12699, n_4311, n12698);
  not g18211 (n_8403, n12695);
  and g18212 (n12700, n_4312, n_8403);
  not g18213 (n_8404, n12699);
  and g18214 (n12701, n_8404, n12700);
  and g18215 (n12702, n_4311, n_8400);
  and g18216 (n12703, n7676, n12698);
  not g18217 (n_8405, n12702);
  and g18218 (n12704, n7685, n_8405);
  not g18219 (n_8406, n12703);
  and g18220 (n12705, n_8406, n12704);
  not g18221 (n_8407, n12701);
  and g18222 (n12706, pi1197, n_8407);
  not g18223 (n_8408, n12705);
  and g18224 (n12707, n_8408, n12706);
  not g18225 (n_8409, n12707);
  and g18226 (n12708, n12685, n_8409);
  not g18227 (n_8410, n12683);
  and g18228 (n12709, n_4718, n_8410);
  not g18229 (n_8411, n12708);
  and g18230 (n12710, n_8411, n12709);
  not g18231 (n_8412, n12682);
  not g18232 (n_8413, n12710);
  and g18233 (n12711, n_8412, n_8413);
  not g18234 (n_8414, n12711);
  and g18235 (n12712, n_4392, n_8414);
  and g18236 (n12713, n8499, n12681);
  and g18237 (n12714, n_4377, n12710);
  and g18238 (n12715, pi1198, n_8391);
  not g18239 (n_8415, n12713);
  not g18240 (n_8416, n12715);
  and g18241 (n12716, n_8415, n_8416);
  not g18242 (n_8417, n12714);
  and g18243 (n12717, n_8417, n12716);
  not g18244 (n_8418, n12717);
  and g18245 (n12718, pi0374, n_8418);
  not g18246 (n_8419, n12712);
  not g18247 (n_8420, n12718);
  and g18248 (n12719, n_8419, n_8420);
  not g18249 (n_8421, n12719);
  and g18250 (n12720, pi0369, n_8421);
  and g18251 (n12721, n_4392, n_8418);
  and g18252 (n12722, pi0374, n_8414);
  not g18253 (n_8422, n12721);
  not g18254 (n_8423, n12722);
  and g18255 (n12723, n_8422, n_8423);
  not g18256 (n_8424, n12723);
  and g18257 (n12724, n_4391, n_8424);
  and g18258 (n12725, pi0371, n8853);
  and g18259 (n12726, n_4401, n_5609);
  not g18260 (n_8425, n12725);
  not g18261 (n_8426, n12726);
  and g18262 (n12727, n_8425, n_8426);
  not g18263 (n_8427, n12727);
  and g18264 (n12728, pi0370, n_8427);
  and g18265 (n12729, n_4396, n12727);
  not g18266 (n_8428, n12728);
  not g18267 (n_8429, n12729);
  and g18268 (n12730, n_8428, n_8429);
  not g18269 (n_8430, n12720);
  and g18270 (n12731, n_8430, n12730);
  not g18271 (n_8431, n12724);
  and g18272 (n12732, n_8431, n12731);
  and g18273 (n12733, n_4391, n_8421);
  and g18274 (n12734, pi0369, n_8424);
  not g18275 (n_8432, n12730);
  not g18276 (n_8433, n12733);
  and g18277 (n12735, n_8432, n_8433);
  not g18278 (n_8434, n12734);
  and g18279 (n12736, n_8434, n12735);
  not g18280 (n_8435, n12732);
  and g18281 (n12737, n_4628, n_8435);
  not g18282 (n_8436, n12736);
  and g18283 (n12738, n_8436, n12737);
  not g18284 (n_8437, n12675);
  and g18285 (n12739, n_4423, n_8437);
  not g18286 (n_8438, n12738);
  and g18287 (n12740, n_8438, n12739);
  not g18288 (n_8439, n12740);
  and g18289 (n12741, n_4832, n_8439);
  not g18290 (n_8440, n12566);
  and g18291 (n12742, n_8440, n12741);
  not g18292 (n_8441, n12742);
  and g18293 (n12743, n_4091, n_8441);
  not g18294 (n_8442, n12492);
  and g18295 (n12744, n_8442, n12743);
  and g18296 (n12745, n_4196, n12181);
  and g18297 (n12746, pi0075, n12179);
  and g18298 (n12747, n_8079, n_8147);
  and g18299 (n12748, n8162, n_8087);
  not g18300 (n_8443, n12747);
  and g18301 (n12749, n_8443, n12748);
  and g18302 (n12750, n_8079, n_8144);
  and g18303 (n12751, n2610, n_8087);
  not g18304 (n_8444, n12750);
  and g18305 (n12752, n_8444, n12751);
  and g18306 (n12753, n_251, n12179);
  not g18307 (n_8445, n12749);
  not g18308 (n_8446, n12753);
  and g18309 (n12754, n_8445, n_8446);
  not g18310 (n_8447, n12752);
  and g18311 (n12755, n_8447, n12754);
  not g18312 (n_8448, n12755);
  and g18313 (n12756, n_171, n_8448);
  not g18314 (n_8449, n12746);
  not g18315 (n_8450, n12756);
  and g18316 (n12757, n_8449, n_8450);
  not g18317 (n_8451, n12757);
  and g18318 (n12758, pi0567, n_8451);
  not g18319 (n_8452, n12758);
  and g18320 (n12759, n12568, n_8452);
  not g18321 (n_8453, n12745);
  not g18322 (n_8454, n12759);
  and g18323 (n12760, n_8453, n_8454);
  and g18324 (n12761, n_4239, n12760);
  not g18325 (n_8455, n12761);
  and g18326 (n12762, n_8054, n_8455);
  and g18327 (n12763, n_5023, n12762);
  not g18328 (n_8456, n12762);
  and g18329 (n12764, pi0443, n_8456);
  not g18330 (n_8457, n12764);
  and g18331 (n12765, n_8163, n_8457);
  and g18332 (n12766, n8249, n12765);
  and g18333 (n12767, n_4947, n_8456);
  not g18334 (n_8458, n12767);
  and g18335 (n12768, n_8165, n_8458);
  and g18336 (n12769, n_5092, n12768);
  not g18337 (n_8459, n12766);
  not g18338 (n_8460, n12769);
  and g18339 (n12770, n_8459, n_8460);
  not g18340 (n_8461, n12770);
  and g18341 (n12771, pi0435, n_8461);
  and g18342 (n12772, n_4952, n12768);
  and g18343 (n12773, pi0444, n12765);
  not g18344 (n_8462, n12772);
  and g18345 (n12774, n_4948, n_8462);
  not g18346 (n_8463, n12773);
  and g18347 (n12775, n_8463, n12774);
  and g18348 (n12776, n_4952, n12765);
  and g18349 (n12777, pi0444, n12768);
  not g18350 (n_8464, n12776);
  and g18351 (n12778, pi0436, n_8464);
  not g18352 (n_8465, n12777);
  and g18353 (n12779, n_8465, n12778);
  not g18354 (n_8466, n12775);
  not g18355 (n_8467, n12779);
  and g18356 (n12780, n_8466, n_8467);
  and g18357 (n12781, n_4922, n12780);
  not g18358 (n_8468, n12771);
  not g18359 (n_8469, n12781);
  and g18360 (n12782, n_8468, n_8469);
  and g18361 (n12783, n_4921, n12782);
  and g18362 (n12784, n_4922, n_8461);
  and g18363 (n12785, pi0435, n12780);
  not g18364 (n_8470, n12784);
  not g18365 (n_8471, n12785);
  and g18366 (n12786, n_8470, n_8471);
  and g18367 (n12787, pi0429, n12786);
  not g18368 (n_8472, n12783);
  and g18369 (n12788, n8105, n_8472);
  not g18370 (n_8473, n12787);
  and g18371 (n12789, n_8473, n12788);
  and g18372 (n12790, n_4921, n12786);
  and g18373 (n12791, pi0429, n12782);
  not g18374 (n_8474, n12790);
  and g18375 (n12792, n_4942, n_8474);
  not g18376 (n_8475, n12791);
  and g18377 (n12793, n_8475, n12792);
  not g18378 (n_8476, n12789);
  and g18379 (n12794, pi1196, n_8476);
  not g18380 (n_8477, n12793);
  and g18381 (n12795, n_8477, n12794);
  not g18382 (n_8478, n12795);
  and g18383 (n12796, n12412, n_8478);
  not g18384 (n_8479, n12763);
  not g18385 (n_8480, n12796);
  and g18386 (n12797, n_8479, n_8480);
  and g18387 (n12798, n_4718, n12797);
  not g18388 (n_8481, n12797);
  and g18389 (n12799, n_4976, n_8481);
  and g18390 (n12800, pi0428, n12762);
  not g18391 (n_8482, n12799);
  not g18392 (n_8483, n12800);
  and g18393 (n12801, n_8482, n_8483);
  not g18394 (n_8484, n12801);
  and g18395 (n12802, n_4974, n_8484);
  and g18396 (n12803, pi0428, n_8481);
  and g18397 (n12804, n_4976, n12762);
  not g18398 (n_8485, n12803);
  not g18399 (n_8486, n12804);
  and g18400 (n12805, n_8485, n_8486);
  not g18401 (n_8487, n12805);
  and g18402 (n12806, pi0427, n_8487);
  not g18403 (n_8488, n12802);
  not g18404 (n_8489, n12806);
  and g18405 (n12807, n_8488, n_8489);
  not g18406 (n_8490, n12807);
  and g18407 (n12808, pi0430, n_8490);
  and g18408 (n12809, n_4974, n_8487);
  and g18409 (n12810, pi0427, n_8484);
  not g18410 (n_8491, n12809);
  not g18411 (n_8492, n12810);
  and g18412 (n12811, n_8491, n_8492);
  not g18413 (n_8493, n12811);
  and g18414 (n12812, n_4981, n_8493);
  not g18415 (n_8494, n12808);
  not g18416 (n_8495, n12812);
  and g18417 (n12813, n_8494, n_8495);
  not g18418 (n_8496, n12813);
  and g18419 (n12814, pi0426, n_8496);
  and g18420 (n12815, pi0430, n_8493);
  and g18421 (n12816, n_4981, n_8490);
  not g18422 (n_8497, n12815);
  not g18423 (n_8498, n12816);
  and g18424 (n12817, n_8497, n_8498);
  not g18425 (n_8499, n12817);
  and g18426 (n12818, n_4985, n_8499);
  not g18427 (n_8500, n12814);
  not g18428 (n_8501, n12818);
  and g18429 (n12819, n_8500, n_8501);
  not g18430 (n_8502, n12819);
  and g18431 (n12820, pi0445, n_8502);
  and g18432 (n12821, pi0426, n_8499);
  and g18433 (n12822, n_4985, n_8496);
  not g18434 (n_8503, n12821);
  not g18435 (n_8504, n12822);
  and g18436 (n12823, n_8503, n_8504);
  not g18437 (n_8505, n12823);
  and g18438 (n12824, n_4990, n_8505);
  not g18439 (n_8506, n12820);
  not g18440 (n_8507, n12824);
  and g18441 (n12825, n_8506, n_8507);
  and g18442 (n12826, pi0448, n12825);
  and g18443 (n12827, pi0445, n_8505);
  and g18444 (n12828, n_4990, n_8502);
  not g18445 (n_8508, n12827);
  not g18446 (n_8509, n12828);
  and g18447 (n12829, n_8508, n_8509);
  and g18448 (n12830, n_4995, n12829);
  not g18449 (n_8510, n12826);
  and g18450 (n12831, n8128, n_8510);
  not g18451 (n_8511, n12830);
  and g18452 (n12832, n_8511, n12831);
  and g18453 (n12833, pi0448, n12829);
  and g18454 (n12834, n_4995, n12825);
  not g18455 (n_8512, n12833);
  and g18456 (n12835, n_5003, n_8512);
  not g18457 (n_8513, n12834);
  and g18458 (n12836, n_8513, n12835);
  not g18459 (n_8514, n12832);
  and g18460 (n12837, pi1199, n_8514);
  not g18461 (n_8515, n12836);
  and g18462 (n12838, n_8515, n12837);
  not g18463 (n_8516, n12798);
  and g18464 (n12839, n8041, n_8516);
  not g18465 (n_8517, n12838);
  and g18466 (n12840, n_8517, n12839);
  not g18467 (n_8518, n12840);
  and g18468 (n12841, n12186, n_8518);
  and g18469 (n12842, n_8053, n_8456);
  and g18470 (n12843, n8410, n12568);
  not g18471 (n_8519, n12843);
  and g18472 (n12844, n_7978, n_8519);
  and g18473 (n12845, n7958, n_8453);
  and g18474 (n12846, n_8079, n_8325);
  not g18475 (n_8520, n12846);
  and g18476 (n12847, n12748, n_8520);
  not g18477 (n_8521, n12588);
  and g18478 (n12848, n_8079, n_8521);
  not g18479 (n_8522, n12848);
  and g18480 (n12849, n12751, n_8522);
  not g18481 (n_8523, n12847);
  and g18482 (n12850, n_8446, n_8523);
  not g18483 (n_8524, n12849);
  and g18484 (n12851, n_8524, n12850);
  and g18485 (n12852, n7926, n12749);
  not g18486 (n_8525, n12611);
  and g18487 (n12853, n_8525, n12752);
  not g18488 (n_8526, n12852);
  not g18489 (n_8527, n12853);
  and g18490 (n12854, n_8526, n_8527);
  and g18491 (n12855, n12851, n12854);
  not g18492 (n_8528, n12855);
  and g18493 (n12856, n12845, n_8528);
  not g18494 (n_8529, n12629);
  and g18495 (n12857, n_8529, n12749);
  not g18496 (n_8530, n12857);
  and g18497 (n12858, n_8446, n_8530);
  and g18498 (n12859, n_8527, n12858);
  and g18499 (n12860, n8668, n_8453);
  not g18500 (n_8531, n12859);
  and g18501 (n12861, n_8531, n12860);
  not g18502 (n_8532, n12856);
  not g18503 (n_8533, n12861);
  and g18504 (n12862, n_8532, n_8533);
  and g18505 (n12863, n_171, pi0567);
  not g18506 (n_8534, n12862);
  and g18507 (n12864, n_8534, n12863);
  not g18508 (n_8535, n12844);
  and g18509 (n12865, pi1199, n_8535);
  not g18510 (n_8536, n12864);
  and g18511 (n12866, n_8536, n12865);
  not g18512 (n_8537, n12851);
  and g18513 (n12867, n_171, n_8537);
  not g18514 (n_8538, n12867);
  and g18515 (n12868, n_8449, n_8538);
  not g18516 (n_8539, n12868);
  and g18517 (n12869, pi0567, n_8539);
  not g18518 (n_8540, n12869);
  and g18519 (n12870, n12568, n_8540);
  not g18520 (n_8541, n12870);
  and g18521 (n12871, n12845, n_8541);
  and g18522 (n12872, n_4718, n12277);
  not g18523 (n_8542, n12871);
  and g18524 (n12873, n_8542, n12872);
  not g18525 (n_8543, n12866);
  and g18526 (n12874, n_5238, n_8543);
  not g18527 (n_8544, n12873);
  and g18528 (n12875, n_8544, n12874);
  and g18529 (n12876, n_4723, n12875);
  not g18530 (n_8545, n12842);
  not g18531 (n_8546, n12876);
  and g18532 (n12877, n_8545, n_8546);
  not g18533 (n_8547, n12877);
  and g18534 (n12878, n_4773, n_8547);
  and g18535 (n12879, n8395, n_8456);
  not g18536 (n_8548, n12875);
  not g18537 (n_8549, n12879);
  and g18538 (n12880, n_8548, n_8549);
  not g18539 (n_8550, n12880);
  and g18540 (n12881, pi0333, n_8550);
  not g18541 (n_8551, n12878);
  not g18542 (n_8552, n12881);
  and g18543 (n12882, n_8551, n_8552);
  not g18544 (n_8553, n12882);
  and g18545 (n12883, n_4778, n_8553);
  and g18546 (n12884, pi0333, n_8547);
  and g18547 (n12885, n_4773, n_8550);
  not g18548 (n_8554, n12884);
  not g18549 (n_8555, n12885);
  and g18550 (n12886, n_8554, n_8555);
  not g18551 (n_8556, n12886);
  and g18552 (n12887, pi0391, n_8556);
  not g18553 (n_8557, n12883);
  not g18554 (n_8558, n12887);
  and g18555 (n12888, n_8557, n_8558);
  not g18556 (n_8559, n12888);
  and g18557 (n12889, n_4785, n_8559);
  and g18558 (n12890, n_4778, n_8556);
  and g18559 (n12891, pi0391, n_8553);
  not g18560 (n_8560, n12890);
  not g18561 (n_8561, n12891);
  and g18562 (n12892, n_8560, n_8561);
  not g18563 (n_8562, n12892);
  and g18564 (n12893, pi0392, n_8562);
  not g18565 (n_8563, n12889);
  not g18566 (n_8564, n12893);
  and g18567 (n12894, n_8563, n_8564);
  not g18568 (n_8565, n12894);
  and g18569 (n12895, n_4793, n_8565);
  and g18570 (n12896, n_4785, n_8562);
  and g18571 (n12897, pi0392, n_8559);
  not g18572 (n_8566, n12896);
  not g18573 (n_8567, n12897);
  and g18574 (n12898, n_8566, n_8567);
  not g18575 (n_8568, n12898);
  and g18576 (n12899, pi0393, n_8568);
  not g18577 (n_8569, n12895);
  and g18578 (n12900, n_4821, n_8569);
  not g18579 (n_8570, n12899);
  and g18580 (n12901, n_8570, n12900);
  and g18581 (n12902, n_4793, n_8568);
  and g18582 (n12903, pi0393, n_8565);
  not g18583 (n_8571, n12902);
  and g18584 (n12904, n8028, n_8571);
  not g18585 (n_8572, n12903);
  and g18586 (n12905, n_8572, n12904);
  not g18587 (n_8573, n12901);
  and g18588 (n12906, pi0591, n_8573);
  not g18589 (n_8574, n12905);
  and g18590 (n12907, n_8574, n12906);
  and g18591 (n12908, pi0592, n12760);
  not g18592 (n_8575, n12908);
  and g18593 (n12909, n_8386, n_8575);
  and g18594 (n12910, n_4370, n12909);
  and g18595 (n12911, pi1199, n_8389);
  not g18596 (n_8576, n12910);
  and g18597 (n12912, n_8576, n12911);
  and g18598 (n12913, n7673, n7688);
  and g18599 (n12914, n_4320, n_4316);
  not g18600 (n_8577, n12913);
  not g18601 (n_8578, n12914);
  and g18602 (n12915, n_8577, n_8578);
  not g18603 (n_8579, n12915);
  and g18604 (n12916, pi0367, n_8579);
  and g18605 (n12917, n_4317, n12915);
  not g18606 (n_8580, n12916);
  not g18607 (n_8581, n12917);
  and g18608 (n12918, n_8580, n_8581);
  not g18609 (n_8582, n12918);
  and g18610 (n12919, n12181, n_8582);
  and g18611 (n12920, n12909, n12918);
  not g18612 (n_8583, n12919);
  and g18613 (n12921, pi1197, n_8583);
  not g18614 (n_8584, n12920);
  and g18615 (n12922, n_8584, n12921);
  not g18616 (n_8585, n12922);
  and g18617 (n12923, n12685, n_8585);
  and g18618 (n12924, n7670, n12909);
  not g18619 (n_8586, n12924);
  and g18620 (n12925, n_4718, n_8586);
  not g18621 (n_8587, n12923);
  and g18622 (n12926, n_8587, n12925);
  not g18623 (n_8588, n12912);
  not g18624 (n_8589, n12926);
  and g18625 (n12927, n_8588, n_8589);
  not g18626 (n_8590, n12927);
  and g18627 (n12928, n_4392, n_8590);
  and g18628 (n12929, n_4377, n_8590);
  not g18629 (n_8591, n12909);
  and g18630 (n12930, pi1198, n_8591);
  not g18631 (n_8592, n12929);
  not g18632 (n_8593, n12930);
  and g18633 (n12931, n_8592, n_8593);
  not g18634 (n_8594, n12931);
  and g18635 (n12932, pi0374, n_8594);
  not g18636 (n_8595, n12928);
  not g18637 (n_8596, n12932);
  and g18638 (n12933, n_8595, n_8596);
  not g18639 (n_8597, n12933);
  and g18640 (n12934, n_4391, n_8597);
  and g18641 (n12935, n_4392, n_8594);
  and g18642 (n12936, pi0374, n_8590);
  not g18643 (n_8598, n12935);
  not g18644 (n_8599, n12936);
  and g18645 (n12937, n_8598, n_8599);
  not g18646 (n_8600, n12937);
  and g18647 (n12938, pi0369, n_8600);
  not g18648 (n_8601, n12934);
  and g18649 (n12939, n_8432, n_8601);
  not g18650 (n_8602, n12938);
  and g18651 (n12940, n_8602, n12939);
  and g18652 (n12941, pi0369, n_8597);
  and g18653 (n12942, n_4391, n_8600);
  not g18654 (n_8603, n12941);
  and g18655 (n12943, n12730, n_8603);
  not g18656 (n_8604, n12942);
  and g18657 (n12944, n_8604, n12943);
  not g18658 (n_8605, n12940);
  and g18659 (n12945, n_4628, n_8605);
  not g18660 (n_8606, n12944);
  and g18661 (n12946, n_8606, n12945);
  not g18662 (n_8607, n12946);
  and g18663 (n12947, n_4423, n_8607);
  not g18664 (n_8608, n12907);
  and g18665 (n12948, n_8608, n12947);
  and g18666 (n12949, n_8227, n12762);
  not g18667 (n_8609, n12949);
  and g18668 (n12950, n_8228, n_8609);
  not g18669 (n_8610, n12950);
  and g18670 (n12951, pi1198, n_8610);
  and g18671 (n12952, n_4486, n12762);
  not g18672 (n_8611, n12952);
  and g18673 (n12953, n_8231, n_8611);
  not g18674 (n_8612, n12953);
  and g18675 (n12954, pi0355, n_8612);
  and g18676 (n12955, n_4480, n_8456);
  not g18677 (n_8613, n12955);
  and g18678 (n12956, n_8234, n_8613);
  not g18679 (n_8614, n12956);
  and g18680 (n12957, n_4481, n_8614);
  and g18681 (n12958, pi0455, n_8456);
  not g18682 (n_8615, n12958);
  and g18683 (n12959, n_8237, n_8615);
  not g18684 (n_8616, n12959);
  and g18685 (n12960, pi0452, n_8616);
  not g18686 (n_8617, n12957);
  not g18687 (n_8618, n12960);
  and g18688 (n12961, n_8617, n_8618);
  and g18689 (n12962, n_4485, n12961);
  not g18690 (n_8619, n12954);
  not g18691 (n_8620, n12962);
  and g18692 (n12963, n_8619, n_8620);
  and g18693 (n12964, n_4491, n12963);
  and g18694 (n12965, n_4485, n_8612);
  and g18695 (n12966, pi0355, n12961);
  not g18696 (n_8621, n12965);
  not g18697 (n_8622, n12966);
  and g18698 (n12967, n_8621, n_8622);
  and g18699 (n12968, pi0458, n12967);
  not g18700 (n_8623, n12964);
  and g18701 (n12969, n_4511, n_8623);
  not g18702 (n_8624, n12968);
  and g18703 (n12970, n_8624, n12969);
  and g18704 (n12971, n_4491, n12967);
  and g18705 (n12972, pi0458, n12963);
  not g18706 (n_8625, n12971);
  and g18707 (n12973, n7812, n_8625);
  not g18708 (n_8626, n12972);
  and g18709 (n12974, n_8626, n12973);
  not g18710 (n_8627, n12970);
  and g18711 (n12975, pi1196, n_8627);
  not g18712 (n_8628, n12974);
  and g18713 (n12976, n_8628, n12975);
  not g18714 (n_8629, n12976);
  and g18715 (n12977, n12497, n_8629);
  not g18716 (n_8630, n12951);
  not g18717 (n_8631, n12977);
  and g18718 (n12978, n_8630, n_8631);
  not g18719 (n_8632, n12978);
  and g18720 (n12979, n_4565, n_8632);
  and g18721 (n12980, n7782, n12762);
  not g18722 (n_8633, n12979);
  not g18723 (n_8634, n12980);
  and g18724 (n12981, n_8633, n_8634);
  and g18725 (n12982, n_4569, n12981);
  and g18726 (n12983, pi1199, n_8456);
  and g18727 (n12984, pi0351, n12983);
  not g18728 (n_8635, n12982);
  not g18729 (n_8636, n12984);
  and g18730 (n12985, n_8635, n_8636);
  not g18731 (n_8637, n12985);
  and g18732 (n12986, n_4575, n_8637);
  and g18733 (n12987, n_4578, n12981);
  and g18734 (n12988, n_4577, n12983);
  not g18735 (n_8638, n12987);
  not g18736 (n_8639, n12988);
  and g18737 (n12989, n_8638, n_8639);
  not g18738 (n_8640, n12989);
  and g18739 (n12990, pi0461, n_8640);
  not g18740 (n_8641, n12986);
  not g18741 (n_8642, n12990);
  and g18742 (n12991, n_8641, n_8642);
  not g18743 (n_8643, n12991);
  and g18744 (n12992, n_4585, n_8643);
  and g18745 (n12993, n_4575, n_8640);
  and g18746 (n12994, pi0461, n_8637);
  not g18747 (n_8644, n12993);
  not g18748 (n_8645, n12994);
  and g18749 (n12995, n_8644, n_8645);
  not g18750 (n_8646, n12995);
  and g18751 (n12996, pi0357, n_8646);
  not g18752 (n_8647, n12992);
  not g18753 (n_8648, n12996);
  and g18754 (n12997, n_8647, n_8648);
  not g18755 (n_8649, n12997);
  and g18756 (n12998, n_4593, n_8649);
  and g18757 (n12999, n_4585, n_8646);
  and g18758 (n13000, pi0357, n_8643);
  not g18759 (n_8650, n12999);
  not g18760 (n_8651, n13000);
  and g18761 (n13001, n_8650, n_8651);
  not g18762 (n_8652, n13001);
  and g18763 (n13002, pi0356, n_8652);
  not g18764 (n_8653, n12998);
  not g18765 (n_8654, n13002);
  and g18766 (n13003, n_8653, n_8654);
  not g18767 (n_8655, n13003);
  and g18768 (n13004, n_4616, n_8655);
  and g18769 (n13005, n_4593, n_8652);
  and g18770 (n13006, pi0356, n_8649);
  not g18771 (n_8656, n13005);
  not g18772 (n_8657, n13006);
  and g18773 (n13007, n_8656, n_8657);
  not g18774 (n_8658, n13007);
  and g18775 (n13008, pi0354, n_8658);
  not g18776 (n_8659, n13004);
  and g18777 (n13009, n_4615, n_8659);
  not g18778 (n_8660, n13008);
  and g18779 (n13010, n_8660, n13009);
  and g18780 (n13011, n_4616, n_8658);
  and g18781 (n13012, pi0354, n_8655);
  not g18782 (n_8661, n13011);
  and g18783 (n13013, n7887, n_8661);
  not g18784 (n_8662, n13012);
  and g18785 (n13014, n_8662, n13013);
  not g18786 (n_8663, n13010);
  and g18787 (n13015, n_4628, n_8663);
  not g18788 (n_8664, n13014);
  and g18789 (n13016, n_8664, n13015);
  not g18790 (n_8665, n13016);
  and g18791 (n13017, n12237, n_8665);
  not g18792 (n_8666, n12948);
  and g18793 (n13018, n_4832, n_8666);
  not g18794 (n_8667, n13017);
  and g18795 (n13019, n_8667, n13018);
  not g18796 (n_8668, n13019);
  and g18797 (n13020, n7425, n_8668);
  not g18798 (n_8669, n12841);
  and g18799 (n13021, n_8669, n13020);
  not g18805 (n_8672, n12366);
  and g18806 (n13025, n_5623, n_8672);
  not g18807 (n_8673, n13024);
  and g18808 (n13026, n_8673, n13025);
  not g18809 (n_8674, n12183);
  and g18810 (n13027, n7643, n_8674);
  not g18811 (n_8675, n13026);
  and g18812 (po0238, n_8675, n13027);
  and g18813 (n13029, n_4226, n11302);
  and g18814 (n13030, pi0081, n_3310);
  and g18815 (n13031, n2489, n13030);
  not g18821 (n_8676, n13031);
  not g18822 (n_8677, n13036);
  and g18823 (n13037, n_8676, n_8677);
  not g18824 (n_8678, n13037);
  and g18825 (po0239, n13029, n_8678);
  and g18826 (n13039, pi0069, pi0314);
  and g18827 (n13040, n2792, n13039);
  not g18831 (n_8679, n13040);
  not g18832 (n_8680, n13043);
  and g18833 (n13044, n_8679, n_8680);
  and g18834 (n13045, n11103, n11107);
  not g18835 (n_8681, n13044);
  and g18836 (po0240, n_8681, n13045);
  and g18837 (n13047, n2480, n2799);
  and g18838 (n13048, pi0084, n9077);
  and g18839 (n13049, n13047, n13048);
  and g18840 (n13050, n2467, n13049);
  and g18841 (n13051, n2499, n11102);
  and g18842 (n13052, n2702, n13051);
  and g18843 (n13053, n13050, n13052);
  not g18844 (n_8682, n13053);
  and g18845 (n13054, pi0314, n_8682);
  not g18846 (n_8683, n13049);
  and g18847 (n13055, n_60, n_8683);
  not g18848 (n_8684, n13055);
  and g18849 (n13056, n13052, n_8684);
  and g18850 (n13057, n2795, n13056);
  not g18851 (n_8685, n13057);
  and g18852 (n13058, n_3310, n_8685);
  not g18853 (n_8686, n13054);
  and g18854 (n13059, n10166, n_8686);
  not g18855 (n_8687, n13058);
  and g18856 (po0241, n_8687, n13059);
  and g18857 (n13061, pi0211, pi0299);
  and g18858 (n13062, pi0219, pi0299);
  not g18859 (n_8688, n13061);
  not g18860 (n_8689, n13062);
  and g18861 (n13063, n_8688, n_8689);
  and g18862 (n13064, n_7047, n13063);
  and g18863 (n13065, n_4226, n13064);
  and g18864 (po0242, n11385, n13065);
  and g18865 (n13067, n6423, n11104);
  and g18866 (n13068, n_3310, n11105);
  and g18867 (n13069, n11437, n13068);
  not g18868 (n_8690, n13067);
  not g18869 (n_8691, n13069);
  and g18870 (n13070, n_8690, n_8691);
  not g18871 (n_8692, n13070);
  and g18872 (po0243, n11107, n_8692);
  and g18873 (n13072, n7603, n11396);
  and g18874 (n13073, n7606, n11399);
  not g18875 (n_8693, n13072);
  not g18876 (n_8694, n13073);
  and g18877 (n13074, n_8693, n_8694);
  not g18878 (n_8695, n13074);
  and g18879 (po0244, n10983, n_8695);
  and g18880 (n13076, n2845, n13051);
  and g18881 (n13077, pi0314, n10166);
  and g18882 (n13078, n2702, n13077);
  and g18883 (po0245, n13076, n13078);
  and g18884 (n13080, n2708, n7417);
  not g18890 (n_8696, n13085);
  and g18891 (n13086, n_4091, n_8696);
  and g18892 (n13087, n7417, n11030);
  not g18893 (n_8697, n13087);
  and g18894 (n13088, n_3206, n_8697);
  and g18895 (n13089, n7439, n12376);
  and g18896 (n13090, n11027, n13089);
  and g18897 (n13091, n11043, n12374);
  and g18898 (n13092, n13090, n13091);
  not g18899 (n_8698, n13092);
  and g18900 (n13093, pi1093, n_8698);
  not g18906 (n_8701, n13096);
  and g18907 (n13097, n7425, n_8701);
  not g18908 (n_8702, n13086);
  and g18909 (n13098, n_4226, n_8702);
  not g18910 (n_8703, n13097);
  and g18911 (po0246, n_8703, n13098);
  and g18915 (n13103, pi0841, n7445);
  and g18916 (n13104, n13102, n13103);
  not g18917 (n_8704, n13104);
  and g18918 (n13105, n_139, n_8704);
  not g18919 (n_8705, n8959);
  and g18920 (n13106, pi0070, n_8705);
  not g18926 (n_8708, pi1050);
  and g18927 (n13110, n_8708, n9090);
  not g18928 (n_8709, n13110);
  and g18929 (n13111, n_43, n_8709);
  and g18934 (n13115, n_42, n2756);
  not g18935 (n_8711, n13115);
  and g18936 (n13116, n_6593, n_8711);
  and g18937 (n13117, n2928, n10162);
  not g18938 (n_8712, n13116);
  and g18939 (n13118, n_8712, n13117);
  not g18944 (n_8713, n13122);
  and g18945 (n13123, n_162, n_8713);
  not g18946 (n_8714, n13118);
  and g18947 (n13124, n_8714, n13123);
  not g18948 (n_8715, n13124);
  and g18949 (n13125, n10197, n_8715);
  and g18950 (po0249, n7612, n13125);
  and g18951 (n13127, pi0092, n2521);
  and g18952 (n13128, n3373, n11473);
  and g18953 (n13129, n13127, n13128);
  and g18954 (n13130, n5853, n6235);
  and g18955 (n13131, n7603, n13130);
  and g18956 (n13132, n3470, n6189);
  and g18957 (n13133, n7606, n13132);
  not g18958 (n_8716, n13131);
  not g18959 (n_8717, n13133);
  and g18960 (n13134, n_8716, n_8717);
  and g18961 (n13135, n2534, n11211);
  not g18962 (n_8718, n13134);
  and g18963 (n13136, n_8718, n13135);
  not g18964 (n_8719, n13129);
  not g18965 (n_8720, n13136);
  and g18966 (n13137, n_8719, n_8720);
  not g18967 (n_8721, n13137);
  and g18968 (po0250, n10163, n_8721);
  and g18969 (n13139, pi0093, n11086);
  and g18970 (n13140, n2914, n13139);
  not g18971 (n_8722, n13140);
  and g18972 (n13141, n_174, n_8722);
  and g18973 (n13142, n_8708, n2521);
  not g18974 (n_8723, n13142);
  and g18975 (n13143, pi0092, n_8723);
  not g18976 (n_8724, n13141);
  and g18977 (n13144, n10164, n_8724);
  not g18978 (n_8725, n13143);
  and g18979 (po0251, n_8725, n13144);
  and g18980 (n13146, n11068, n11284);
  not g18981 (n_8726, n13146);
  and g18982 (n13147, n_5631, n_8726);
  and g18983 (n13148, n2924, n13146);
  not g18984 (n_8727, n13148);
  and g18985 (n13149, pi1093, n_8727);
  not g18986 (n_8728, n13149);
  and g18987 (n13150, n2933, n_8728);
  and g18988 (n13151, n10243, n11066);
  not g18989 (n_8729, n13151);
  and g18990 (n13152, n_362, n_8729);
  and g18991 (n13153, n2717, n10162);
  and g18992 (n13154, pi0252, n13153);
  not g18993 (n_8730, n13152);
  and g18994 (n13155, n_8730, n13154);
  not g18995 (n_8731, n13150);
  not g18996 (n_8732, n13155);
  and g18997 (n13156, n_8731, n_8732);
  not g18998 (n_8733, n13156);
  and g18999 (n13157, n_5636, n_8733);
  not g19000 (n_8734, n13157);
  and g19001 (n13158, n_8726, n_8734);
  and g19002 (n13159, pi0252, n13156);
  not g19003 (n_8735, n13158);
  not g19004 (n_8736, n13159);
  and g19005 (n13160, n_8735, n_8736);
  not g19006 (n_8737, n13160);
  and g19007 (n13161, n8888, n_8737);
  not g19008 (n_8738, n13147);
  and g19009 (n13162, n10165, n_8738);
  not g19010 (n_8739, n13161);
  and g19011 (po0252, n_8739, n13162);
  and g19012 (n13164, n2517, n11770);
  and g19013 (n13165, n11458, n13164);
  and g19014 (n13166, n_4, n10162);
  and g19015 (n13167, n11283, n13166);
  and g19016 (n13168, n13102, n13167);
  not g19017 (n_8740, n13168);
  and g19018 (n13169, n_162, n_8740);
  not g19019 (n_8741, n13165);
  and g19020 (n13170, n_8741, n13169);
  not g19021 (n_8742, n11422);
  and g19022 (n13171, n_8742, n11425);
  and g19023 (n13172, n_3284, n13171);
  and g19024 (n13173, n_3122, n_3284);
  not g19025 (n_8743, n11419);
  and g19026 (n13174, n3471, n_8743);
  and g19027 (n13175, n13173, n13174);
  not g19028 (n_8744, n13172);
  and g19029 (n13176, pi0039, n_8744);
  not g19030 (n_8745, n13175);
  and g19031 (n13177, n_8745, n13176);
  not g19032 (n_8746, n13170);
  and g19033 (n13178, n10200, n_8746);
  not g19034 (n_8747, n13177);
  and g19035 (po0253, n_8747, n13178);
  and g19036 (n13180, n10325, n13164);
  and g19037 (n13181, pi0479, n_5636);
  and g19038 (n13182, n3183, n13181);
  not g19044 (n_8749, n13182);
  not g19045 (n_8750, n13186);
  and g19046 (n13187, n_8749, n_8750);
  not g19047 (n_8751, n13187);
  and g19048 (n13188, n_144, n_8751);
  not g19049 (n_8752, n13180);
  not g19050 (n_8753, n13188);
  and g19051 (n13189, n_8752, n_8753);
  not g19052 (n_8754, n13189);
  and g19053 (po0254, n10165, n_8754);
  and g19057 (n13194, n6169, n13181);
  not g19058 (n_8755, n13194);
  and g19059 (n13195, n_3209, n_8755);
  not g19064 (n_8757, n13193);
  not g19065 (n_8758, n13198);
  and g19066 (n13199, n_8757, n_8758);
  not g19067 (n_8759, n13199);
  and g19068 (po0255, n10200, n_8759);
  and g19069 (n13201, n_174, n11474);
  not g19070 (n_8760, n13127);
  not g19071 (n_8761, n13201);
  and g19072 (n13202, n_8760, n_8761);
  and g19077 (n13206, n_134, pi0152);
  and g19078 (n13207, n10300, n13206);
  and g19079 (n13208, pi0299, n13207);
  not g19083 (n_8763, n13208);
  not g19084 (n_8764, n13211);
  and g19085 (n13212, n_8763, n_8764);
  not g19086 (n_8765, n13212);
  and g19087 (n13213, pi0232, n_8765);
  not g19088 (n_8766, n13213);
  and g19089 (n13214, pi0039, n_8766);
  and g19090 (n13215, n_134, pi0099);
  not g19091 (n_8767, n13215);
  and g19092 (n13216, n_162, n_8767);
  not g19093 (n_8768, n13214);
  not g19094 (n_8769, n13216);
  and g19095 (n13217, n_8768, n_8769);
  and g19096 (n13218, n_6666, n13217);
  and g19097 (n13219, n_4137, n_8767);
  and g19098 (n13220, n_538, n13215);
  not g19099 (n_8770, n13220);
  and g19100 (n13221, n7506, n_8770);
  not g19101 (n_8771, n10329);
  and g19102 (n13222, n_8771, n13215);
  and g19103 (n13223, n6266, n10919);
  not g19104 (n_8772, n13222);
  not g19105 (n_8773, n13223);
  and g19106 (n13224, n_8772, n_8773);
  not g19107 (n_8774, n13224);
  and g19108 (n13225, n10356, n_8774);
  not g19109 (n_8775, n13225);
  and g19110 (n13226, n13221, n_8775);
  not g19111 (n_8776, n13219);
  not g19112 (n_8777, n13226);
  and g19113 (n13227, n_8776, n_8777);
  not g19114 (n_8778, n13227);
  and g19115 (n13228, n_162, n_8778);
  and g19116 (n13229, n2620, n_8768);
  not g19117 (n_8779, n13228);
  and g19118 (n13230, n_8779, n13229);
  not g19119 (n_8780, n13218);
  and g19120 (n13231, pi0075, n_8780);
  not g19121 (n_8781, n13230);
  and g19122 (n13232, n_8781, n13231);
  and g19123 (n13233, pi0228, n10500);
  and g19124 (n13234, pi0228, n10344);
  not g19125 (n_8782, n13234);
  and g19126 (n13235, n13215, n_8782);
  not g19127 (n_8783, n13235);
  and g19128 (n13236, n2531, n_8783);
  not g19129 (n_8784, n13233);
  and g19130 (n13237, n_8784, n13236);
  not g19131 (n_8785, n13217);
  and g19132 (n13238, n_7065, n_8785);
  not g19133 (n_8786, n13238);
  and g19134 (n13239, pi0087, n_8786);
  not g19135 (n_8787, n13237);
  and g19136 (n13240, n_8787, n13239);
  and g19137 (n13241, pi0038, n_8785);
  and g19138 (n13242, n10478, n_8765);
  and g19139 (n13243, n_7153, n13242);
  and g19140 (n13244, pi0041, pi0072);
  not g19141 (n_8788, n13244);
  and g19142 (n13245, pi0099, n_8788);
  and g19143 (n13246, n_6733, n13245);
  not g19144 (n_8789, n10556);
  and g19145 (n13247, n_188, n_8789);
  not g19146 (n_8790, n13246);
  and g19147 (n13248, n_8790, n13247);
  and g19148 (n13249, n_6766, n13245);
  not g19149 (n_8791, n13249);
  and g19150 (n13250, n10779, n_8791);
  and g19151 (n13251, n_6749, n13245);
  not g19152 (n_8792, n13251);
  and g19153 (n13252, n10778, n_8792);
  not g19154 (n_8793, n13250);
  not g19155 (n_8794, n13252);
  and g19156 (n13253, n_8793, n_8794);
  not g19157 (n_8795, n13253);
  and g19158 (n13254, pi0228, n_8795);
  not g19159 (n_8796, n13248);
  and g19160 (n13255, n_162, n_8796);
  not g19161 (n_8797, n13254);
  and g19162 (n13256, n_8797, n13255);
  not g19163 (n_8798, n13243);
  and g19164 (n13257, n2608, n_8798);
  not g19165 (n_8799, n13256);
  and g19166 (n13258, n_8799, n13257);
  not g19167 (n_8800, n10359);
  and g19168 (n13259, n_8800, n13215);
  and g19169 (n13260, n6265, n10318);
  not g19170 (n_8801, n13259);
  not g19171 (n_8802, n13260);
  and g19172 (n13261, n_8801, n_8802);
  not g19173 (n_8803, n13261);
  and g19174 (n13262, n10356, n_8803);
  not g19175 (n_8804, n13262);
  and g19176 (n13263, n13221, n_8804);
  not g19177 (n_8805, n13263);
  and g19178 (n13264, n_8776, n_8805);
  not g19179 (n_8806, n13264);
  and g19180 (n13265, n_162, n_8806);
  not g19181 (n_8807, n13265);
  and g19182 (n13266, n_8768, n_8807);
  not g19183 (n_8808, n13266);
  and g19184 (n13267, n6285, n_8808);
  not g19191 (n_8812, n13240);
  and g19192 (n13271, n_171, n_8812);
  not g19193 (n_8813, n13270);
  and g19194 (n13272, n_8813, n13271);
  not g19195 (n_8814, n13232);
  not g19196 (n_8815, n13272);
  and g19197 (n13273, n_8814, n_8815);
  not g19198 (n_8816, n13273);
  and g19199 (n13274, n7429, n_8816);
  and g19200 (n13275, n_4196, n_8785);
  not g19201 (n_8817, n13275);
  and g19202 (n13276, n_4226, n_8817);
  not g19203 (n_8818, n13274);
  and g19204 (n13277, n_8818, n13276);
  and g19205 (n13278, pi0232, n13207);
  not g19206 (n_8819, n13278);
  and g19207 (n13279, pi0039, n_8819);
  and g19208 (n13280, po1038, n_8769);
  not g19209 (n_8820, n13279);
  and g19210 (n13281, n_8820, n13280);
  or g19211 (po0257, n13277, n13281);
  not g19212 (n_8821, n6281);
  and g19213 (n13283, n_3214, n_8821);
  not g19214 (n_8822, n7473);
  and g19215 (n13284, n_8822, n10078);
  not g19216 (n_8823, n13284);
  and g19217 (n13285, pi0129, n_8823);
  not g19218 (n_8824, n13285);
  and g19219 (n13286, n7472, n_8824);
  and g19220 (n13287, pi0129, n_6542);
  not g19221 (n_8825, n10081);
  not g19222 (n_8826, n13287);
  and g19223 (n13288, n_8825, n_8826);
  not g19224 (n_8827, n13283);
  not g19225 (n_8828, n13288);
  and g19226 (n13289, n_8827, n_8828);
  not g19227 (n_8829, n13286);
  and g19228 (n13290, n_8829, n13289);
  not g19236 (n_8831, n13293);
  not g19237 (n_8832, n13296);
  and g19238 (n13297, n_8831, n_8832);
  not g19239 (n_8833, n13297);
  and g19240 (n13298, n8881, n_8833);
  and g19241 (po0258, n2521, n13298);
  and g19242 (n13300, n_162, n_6671);
  and g19243 (n13301, pi0152, n3389);
  and g19244 (n13302, n6197, n13301);
  and g19245 (n13303, n_134, n13302);
  not g19246 (n_8834, n13303);
  and g19247 (n13304, pi0299, n_8834);
  and g19248 (n13305, n_298, pi0174);
  and g19249 (n13306, n10295, n13305);
  and g19250 (n13307, n_134, n13306);
  not g19251 (n_8835, n13307);
  and g19252 (n13308, n_234, n_8835);
  not g19253 (n_8836, n13304);
  and g19254 (n13309, pi0232, n_8836);
  not g19255 (n_8837, n13308);
  and g19256 (n13310, n_8837, n13309);
  not g19257 (n_8838, n13310);
  and g19258 (n13311, pi0039, n_8838);
  not g19259 (n_8839, n13300);
  not g19260 (n_8840, n13311);
  and g19261 (n13312, n_8839, n_8840);
  and g19262 (n13313, n_6666, n13312);
  and g19263 (n13314, n_4137, n_6671);
  and g19264 (n13315, n_538, n10322);
  not g19265 (n_8841, n13315);
  and g19266 (n13316, n7506, n_8841);
  and g19267 (n13317, n2924, n_3200);
  not g19268 (n_8842, n10328);
  and g19269 (n13318, n10322, n_8842);
  not g19270 (n_8843, n13318);
  and g19271 (n13319, n_6670, n_8843);
  not g19272 (n_8844, n13319);
  and g19273 (n13320, n13317, n_8844);
  not g19274 (n_8845, n13320);
  and g19275 (n13321, n13316, n_8845);
  not g19276 (n_8846, n13314);
  not g19277 (n_8847, n13321);
  and g19278 (n13322, n_8846, n_8847);
  not g19279 (n_8848, n13322);
  and g19280 (n13323, n_162, n_8848);
  and g19281 (n13324, n2620, n_8840);
  not g19282 (n_8849, n13323);
  and g19283 (n13325, n_8849, n13324);
  not g19284 (n_8850, n13313);
  and g19285 (n13326, pi0075, n_8850);
  not g19286 (n_8851, n13325);
  and g19287 (n13327, n_8851, n13326);
  and g19288 (n13328, n10343, n10931);
  not g19289 (n_8852, n13328);
  and g19290 (n13329, n10322, n_8852);
  and g19291 (n13330, n_3184, n10932);
  not g19292 (n_8853, n13329);
  and g19293 (n13331, n_162, n_8853);
  not g19294 (n_8854, n13330);
  and g19295 (n13332, n_8854, n13331);
  and g19296 (n13333, pi0087, n_8840);
  not g19297 (n_8855, n13332);
  and g19298 (n13334, n_8855, n13333);
  not g19299 (n_8856, n13312);
  and g19300 (n13335, pi0038, n_8856);
  and g19301 (n13336, n10949, n13302);
  not g19302 (n_8857, n13336);
  and g19303 (n13337, pi0299, n_8857);
  and g19304 (n13338, n10949, n13306);
  not g19305 (n_8858, n13338);
  and g19306 (n13339, n_234, n_8858);
  not g19307 (n_8859, n13337);
  and g19308 (n13340, n10478, n_8859);
  not g19309 (n_8860, n13339);
  and g19310 (n13341, n_8860, n13340);
  and g19311 (n13342, pi0101, n10409);
  and g19312 (n13343, n_188, n_6725);
  not g19313 (n_8861, n13342);
  and g19314 (n13344, n_8861, n13343);
  and g19315 (n13345, pi0101, n10457);
  and g19316 (n13346, n2924, n_6760);
  not g19317 (n_8862, n13345);
  and g19318 (n13347, n_8862, n13346);
  and g19319 (n13348, pi0101, n10424);
  and g19320 (n13349, n_538, n_6747);
  not g19321 (n_8863, n13348);
  and g19322 (n13350, n_8863, n13349);
  not g19323 (n_8864, n13347);
  not g19324 (n_8865, n13350);
  and g19325 (n13351, n_8864, n_8865);
  not g19326 (n_8866, n13351);
  and g19327 (n13352, pi0228, n_8866);
  not g19328 (n_8867, n13344);
  and g19329 (n13353, n_162, n_8867);
  not g19330 (n_8868, n13352);
  and g19331 (n13354, n_8868, n13353);
  not g19332 (n_8869, n13341);
  and g19333 (n13355, n2608, n_8869);
  not g19334 (n_8870, n13354);
  and g19335 (n13356, n_8870, n13355);
  and g19336 (n13357, n_6669, n10940);
  not g19337 (n_8871, n13357);
  and g19338 (n13358, n10322, n_8871);
  not g19339 (n_8872, n13358);
  and g19340 (n13359, n_6690, n_8872);
  not g19341 (n_8873, n13359);
  and g19342 (n13360, n13317, n_8873);
  not g19343 (n_8874, n13360);
  and g19344 (n13361, n13316, n_8874);
  not g19345 (n_8875, n13361);
  and g19346 (n13362, n_8846, n_8875);
  not g19347 (n_8876, n13362);
  and g19348 (n13363, n_162, n_8876);
  not g19349 (n_8877, n13363);
  and g19350 (n13364, n_8840, n_8877);
  not g19351 (n_8878, n13364);
  and g19352 (n13365, n6285, n_8878);
  not g19359 (n_8882, n13334);
  and g19360 (n13369, n_171, n_8882);
  not g19361 (n_8883, n13368);
  and g19362 (n13370, n_8883, n13369);
  not g19363 (n_8884, n13327);
  not g19364 (n_8885, n13370);
  and g19365 (n13371, n_8884, n_8885);
  not g19366 (n_8886, n13371);
  and g19367 (n13372, n7429, n_8886);
  and g19368 (n13373, n_4196, n_8856);
  not g19369 (n_8887, n13373);
  and g19370 (n13374, n_4226, n_8887);
  not g19371 (n_8888, n13372);
  and g19372 (n13375, n_8888, n13374);
  and g19373 (n13376, pi0232, n13303);
  not g19374 (n_8889, n13376);
  and g19375 (n13377, pi0039, n_8889);
  and g19376 (n13378, po1038, n_8839);
  not g19377 (n_8890, n13377);
  and g19378 (n13379, n_8890, n13378);
  or g19379 (po0259, n13375, n13379);
  and g19380 (n13381, n2851, n8922);
  and g19381 (po0260, n13029, n13381);
  and g19382 (n13383, pi0109, n2765);
  and g19383 (n13384, n2699, n13383);
  not g19384 (n_8891, n13384);
  and g19385 (n13385, pi0314, n_8891);
  not g19386 (n_8892, n13076);
  and g19387 (n13386, n_112, n_8892);
  not g19388 (n_8893, n13386);
  and g19389 (n13387, n6422, n_8893);
  not g19390 (n_8894, n13387);
  and g19391 (n13388, n_3310, n_8894);
  not g19392 (n_8895, n13385);
  and g19393 (n13389, n11106, n_8895);
  not g19394 (n_8896, n13388);
  and g19395 (po0261, n_8896, n13389);
  and g19396 (n13391, n7425, n_5631);
  not g19397 (n_8897, n13391);
  and g19398 (n13392, n10075, n_8897);
  not g19399 (n_8898, n13392);
  and g19400 (n13393, n10396, n_8898);
  and g19401 (n13394, po1057, n_8698);
  not g19402 (n_8899, n13090);
  and g19403 (n13395, n_113, n_8899);
  not g19408 (n_8901, n13398);
  and g19409 (n13399, n_5630, n_8901);
  and g19415 (n13403, n7474, n_6537);
  and g19416 (n13404, n13398, n13403);
  not g19417 (n_8904, n13402);
  not g19418 (n_8905, n13404);
  and g19419 (n13405, n_8904, n_8905);
  not g19420 (n_8906, n13405);
  and g19421 (n13406, n_4091, n_8906);
  not g19422 (n_8907, n13393);
  not g19423 (n_8908, n13406);
  and g19424 (n13407, n_8907, n_8908);
  not g19425 (n_8909, n13407);
  and g19426 (po0262, n10165, n_8909);
  and g19427 (n13409, pi0024, n11282);
  not g19428 (n_8910, n11281);
  and g19429 (n13410, n_116, n_8910);
  not g19430 (n_8911, n13410);
  and g19431 (n13411, n2723, n_8911);
  and g19432 (n13412, n_4119, n2717);
  and g19433 (n13413, n13411, n13412);
  not g19434 (n_8912, n13409);
  not g19435 (n_8913, n13413);
  and g19436 (n13414, n_8912, n_8913);
  not g19437 (n_8914, n13414);
  and g19438 (n13415, pi0841, n_8914);
  and g19439 (n13416, n8946, n11267);
  not g19440 (n_8915, n13415);
  not g19441 (n_8916, n13416);
  and g19442 (n13417, n_8915, n_8916);
  not g19443 (n_8917, n13417);
  and g19444 (po0264, n10166, n_8917);
  not g19445 (n_8918, pi0999);
  and g19446 (n13419, n_8918, n10166);
  and g19447 (po0265, n11354, n13419);
  and g19448 (n13421, n_122, n7442);
  not g19449 (n_8919, n13421);
  and g19450 (n13422, n_123, n_8919);
  not g19451 (n_8920, n13422);
  and g19452 (n13423, n2701, n_8920);
  and g19453 (n13424, n10244, n13423);
  not g19454 (n_8921, n13424);
  and g19455 (n13425, n_3310, n_8921);
  not g19456 (n_8922, n7444);
  and g19457 (n13426, pi0314, n_8922);
  and g19463 (n13430, n7446, n10238);
  and g19464 (n13431, n13424, n13430);
  not g19465 (n_8925, n13431);
  and g19466 (n13432, n_138, n_8925);
  not g19467 (n_8926, n13429);
  and g19468 (n13433, n_8926, n13432);
  and g19469 (n13434, n2625, n7518);
  not g19470 (n_8927, n13433);
  and g19471 (n13435, n_8927, n13434);
  not g19472 (n_8928, n13435);
  and g19473 (n13436, n_172, n_8928);
  and g19474 (n13437, n6133, n8881);
  not g19475 (n_8929, n13436);
  and g19476 (po0266, n_8929, n13437);
  and g19477 (n13439, n2784, n11442);
  and g19478 (po0267, n13077, n13439);
  and g19485 (n13447, pi0314, n13446);
  and g19486 (n13448, n8888, n10075);
  and g19487 (n13449, n10388, n13448);
  not g19488 (n_8930, n13447);
  not g19489 (n_8931, n13449);
  and g19490 (n13450, n_8930, n_8931);
  not g19491 (n_8932, n13450);
  and g19492 (po0268, n10166, n_8932);
  and g19493 (n13452, pi0072, n10325);
  and g19494 (n13453, n_3310, n13446);
  and g19495 (n13454, n9141, n13453);
  not g19496 (n_8933, n13452);
  not g19497 (n_8934, n13454);
  and g19498 (n13455, n_8933, n_8934);
  and g19499 (n13456, n6479, n10165);
  not g19500 (n_8935, n13455);
  and g19501 (po0269, n_8935, n13456);
  not g19502 (n_8937, pi0124);
  or g19503 (po0270, n_8937, pi0468);
  and g19504 (n13459, n_134, pi0113);
  and g19505 (n13460, n_162, n13459);
  not g19506 (n_8938, n13460);
  and g19507 (n13461, pi0038, n_8938);
  and g19508 (n13462, n2924, n7506);
  and g19509 (n13463, n7479, n10531);
  not g19510 (n_8939, n6272);
  not g19511 (n_8940, n13463);
  and g19512 (n13464, n_8939, n_8940);
  not g19513 (n_8941, n13464);
  and g19514 (n13465, n13462, n_8941);
  not g19515 (n_8942, n13465);
  and g19516 (n13466, n13459, n_8942);
  and g19517 (n13467, n_8939, n13462);
  and g19518 (n13468, n_3193, n13467);
  and g19519 (n13469, n13260, n13468);
  not g19520 (n_8943, n13466);
  not g19521 (n_8944, n13469);
  and g19522 (n13470, n_8943, n_8944);
  not g19523 (n_8945, n13470);
  and g19524 (n13471, n_162, n_8945);
  not g19525 (n_8946, n13471);
  and g19526 (n13472, n6285, n_8946);
  and g19527 (n13473, pi0113, n10550);
  not g19528 (n_8947, n10557);
  and g19529 (n13474, n_188, n_8947);
  not g19530 (n_8948, n13473);
  and g19531 (n13475, n_8948, n13474);
  and g19532 (n13476, n_3193, n10780);
  and g19533 (n13477, n_538, n_6749);
  not g19534 (n_8949, n13477);
  and g19535 (n13478, n_3182, n_8949);
  not g19536 (n_8950, n10460);
  and g19537 (n13479, n_8950, n13478);
  and g19538 (n13480, pi0113, n_6827);
  not g19539 (n_8951, n13479);
  and g19540 (n13481, n_8951, n13480);
  not g19541 (n_8952, n13476);
  and g19542 (n13482, pi0228, n_8952);
  not g19543 (n_8953, n13481);
  and g19544 (n13483, n_8953, n13482);
  not g19545 (n_8954, n13475);
  and g19546 (n13484, n_162, n_8954);
  not g19547 (n_8955, n13483);
  and g19548 (n13485, n_8955, n13484);
  not g19549 (n_8956, n13485);
  and g19550 (n13486, n2608, n_8956);
  not g19551 (n_8957, n13461);
  not g19552 (n_8958, n13472);
  and g19553 (n13487, n_8957, n_8958);
  not g19554 (n_8959, n13486);
  and g19555 (n13488, n_8959, n13487);
  not g19556 (n_8960, n13488);
  and g19557 (n13489, n_172, n_8960);
  and g19558 (n13490, n_958, n13460);
  not g19559 (n_8961, n10532);
  and g19560 (n13491, n_8961, n13459);
  and g19561 (n13492, n_3193, n13233);
  not g19562 (n_8962, n13491);
  not g19563 (n_8963, n13492);
  and g19564 (n13493, n_8962, n_8963);
  not g19565 (n_8964, n13493);
  and g19566 (n13494, n2531, n_8964);
  not g19567 (n_8965, n13490);
  and g19568 (n13495, pi0087, n_8965);
  not g19569 (n_8966, n13494);
  and g19570 (n13496, n_8966, n13495);
  not g19571 (n_8967, n13489);
  not g19572 (n_8968, n13496);
  and g19573 (n13497, n_8967, n_8968);
  not g19574 (n_8969, n13497);
  and g19575 (n13498, n_171, n_8969);
  and g19576 (n13499, n7477, n13469);
  not g19577 (n_8970, n10496);
  and g19578 (n13500, n_8939, n_8970);
  not g19579 (n_8971, n13500);
  and g19580 (n13501, n13462, n_8971);
  not g19581 (n_8972, n13501);
  and g19582 (n13502, n13459, n_8972);
  not g19583 (n_8973, n13499);
  not g19584 (n_8974, n13502);
  and g19585 (n13503, n_8973, n_8974);
  not g19586 (n_8975, n13503);
  and g19587 (n13504, n2610, n_8975);
  and g19588 (n13505, n_6666, n13460);
  not g19589 (n_8976, n13505);
  and g19590 (n13506, pi0075, n_8976);
  not g19591 (n_8977, n13504);
  and g19592 (n13507, n_8977, n13506);
  not g19593 (n_8978, n13498);
  not g19594 (n_8979, n13507);
  and g19595 (n13508, n_8978, n_8979);
  not g19596 (n_8980, n13508);
  and g19597 (n13509, n8881, n_8980);
  not g19598 (n_8981, n8881);
  and g19599 (n13510, n_8981, n_8938);
  not g19600 (n_8982, n13509);
  not g19601 (n_8983, n13510);
  and g19602 (po0271, n_8982, n_8983);
  and g19603 (n13512, n_134, pi0114);
  and g19604 (n13513, n_162, n13512);
  and g19605 (n13514, n_6666, n13513);
  not g19606 (n_8984, n11143);
  not g19607 (n_8985, n13512);
  and g19608 (n13515, n_8984, n_8985);
  and g19609 (n13516, pi0114, n10735);
  not g19610 (n_8986, n13516);
  and g19611 (n13517, n11143, n_8986);
  not g19612 (n_8987, n10505);
  and g19613 (n13518, n_8987, n13517);
  not g19614 (n_8988, n13515);
  and g19615 (n13519, n2610, n_8988);
  not g19616 (n_8989, n13518);
  and g19617 (n13520, n_8989, n13519);
  not g19618 (n_8990, n13514);
  and g19619 (n13521, pi0075, n_8990);
  not g19620 (n_8991, n13520);
  and g19621 (n13522, n_8991, n13521);
  not g19622 (n_8992, n13513);
  and g19623 (n13523, n_958, n_8992);
  and g19624 (n13524, pi0228, n10616);
  and g19625 (n13525, n_3198, n13524);
  not g19626 (n_8993, n13525);
  and g19627 (n13526, n13512, n_8993);
  not g19628 (n_8994, n13526);
  and g19629 (n13527, n2608, n_8994);
  not g19630 (n_8995, n10537);
  and g19631 (n13528, n_8995, n13527);
  not g19632 (n_8996, n13523);
  and g19633 (n13529, n11212, n_8996);
  not g19634 (n_8997, n13528);
  and g19635 (n13530, n_8997, n13529);
  and g19636 (n13531, pi0038, n_8992);
  and g19637 (n13532, pi0114, n_6882);
  not g19638 (n_8998, n13532);
  and g19639 (n13533, n11143, n_8998);
  not g19640 (n_8999, n10504);
  and g19641 (n13534, n_8999, n13533);
  and g19642 (n13535, n_162, n_8988);
  not g19643 (n_9000, n13534);
  and g19644 (n13536, n_9000, n13535);
  not g19645 (n_9001, n13536);
  and g19646 (n13537, n6285, n_9001);
  and g19647 (n13538, n_3197, n_7019);
  and g19648 (n13539, pi0114, n_7027);
  not g19649 (n_9002, n13538);
  not g19650 (n_9003, n13539);
  and g19651 (n13540, n_9002, n_9003);
  not g19652 (n_9004, n13540);
  and g19653 (n13541, n_3198, n_9004);
  and g19654 (n13542, pi0115, n_8985);
  not g19655 (n_9005, n13542);
  and g19656 (n13543, n_162, n_9005);
  not g19657 (n_9006, n13541);
  and g19658 (n13544, n_9006, n13543);
  not g19659 (n_9007, n13544);
  and g19660 (n13545, n2608, n_9007);
  not g19667 (n_9011, n13530);
  and g19668 (n13549, n_171, n_9011);
  not g19669 (n_9012, n13548);
  and g19670 (n13550, n_9012, n13549);
  not g19671 (n_9013, n13522);
  not g19672 (n_9014, n13550);
  and g19673 (n13551, n_9013, n_9014);
  not g19674 (n_9015, n13551);
  and g19675 (n13552, n8881, n_9015);
  and g19676 (n13553, n_8981, n_8992);
  not g19677 (n_9016, n13552);
  not g19678 (n_9017, n13553);
  and g19679 (po0272, n_9016, n_9017);
  and g19680 (n13555, n_134, pi0115);
  and g19681 (n13556, n_162, n13555);
  and g19682 (n13557, n_6666, n13556);
  not g19683 (n_9018, n13462);
  not g19684 (n_9019, n13555);
  and g19685 (n13558, n_9018, n_9019);
  and g19686 (n13559, pi0115, n10735);
  and g19687 (n13560, n_3190, n11125);
  not g19688 (n_9020, n13560);
  and g19689 (n13561, n_3198, n_9020);
  and g19690 (n13562, n10502, n13561);
  and g19691 (n13563, n7477, n13562);
  not g19692 (n_9021, n13559);
  and g19693 (n13564, n13462, n_9021);
  not g19694 (n_9022, n13563);
  and g19695 (n13565, n_9022, n13564);
  not g19696 (n_9023, n13558);
  and g19697 (n13566, n2610, n_9023);
  not g19698 (n_9024, n13565);
  and g19699 (n13567, n_9024, n13566);
  not g19700 (n_9025, n13557);
  and g19701 (n13568, pi0075, n_9025);
  not g19702 (n_9026, n13567);
  and g19703 (n13569, n_9026, n13568);
  not g19704 (n_9027, n13556);
  and g19705 (n13570, n_958, n_9027);
  not g19706 (n_9028, n13524);
  and g19707 (n13571, n_9028, n13555);
  not g19708 (n_9029, n13571);
  and g19709 (n13572, n2608, n_9029);
  not g19710 (n_9030, n10536);
  and g19711 (n13573, n_9030, n13572);
  not g19712 (n_9031, n13570);
  and g19713 (n13574, n11212, n_9031);
  not g19714 (n_9032, n13573);
  and g19715 (n13575, n_9032, n13574);
  and g19716 (n13576, pi0038, n_9027);
  and g19717 (n13577, pi0115, n_6882);
  not g19718 (n_9033, n13577);
  and g19719 (n13578, n13462, n_9033);
  not g19720 (n_9034, n13562);
  and g19721 (n13579, n_9034, n13578);
  and g19722 (n13580, n_162, n_9023);
  not g19723 (n_9035, n13579);
  and g19724 (n13581, n_9035, n13580);
  not g19725 (n_9036, n13581);
  and g19726 (n13582, n6285, n_9036);
  and g19727 (n13583, n_3198, n_7019);
  and g19728 (n13584, pi0115, n_7027);
  not g19729 (n_9037, n13583);
  and g19730 (n13585, n_162, n_9037);
  not g19731 (n_9038, n13584);
  and g19732 (n13586, n_9038, n13585);
  not g19733 (n_9039, n13586);
  and g19734 (n13587, n2608, n_9039);
  not g19741 (n_9043, n13575);
  and g19742 (n13591, n_171, n_9043);
  not g19743 (n_9044, n13590);
  and g19744 (n13592, n_9044, n13591);
  not g19745 (n_9045, n13569);
  not g19746 (n_9046, n13592);
  and g19747 (n13593, n_9045, n_9046);
  not g19748 (n_9047, n13593);
  and g19749 (n13594, n8881, n_9047);
  and g19750 (n13595, n_8981, n_9027);
  not g19751 (n_9048, n13594);
  not g19752 (n_9049, n13595);
  and g19753 (po0273, n_9048, n_9049);
  and g19754 (n13597, n_134, pi0116);
  and g19755 (n13598, n_162, n13597);
  not g19756 (n_9050, n13598);
  and g19757 (n13599, pi0038, n_9050);
  and g19758 (n13600, n_3193, n10532);
  not g19759 (n_9051, n13600);
  and g19760 (n13601, n13597, n_9051);
  not g19761 (n_9052, n13601);
  and g19762 (n13602, n_161, n_9052);
  not g19763 (n_9053, n10535);
  and g19764 (n13603, n_9053, n13602);
  not g19765 (n_9054, n13599);
  not g19766 (n_9055, n13603);
  and g19767 (n13604, n_9054, n_9055);
  not g19768 (n_9056, n13604);
  and g19769 (n13605, n_164, n_9056);
  and g19770 (n13606, pi0100, n_9050);
  not g19771 (n_9057, n13606);
  and g19772 (n13607, n11212, n_9057);
  not g19773 (n_9058, n13605);
  and g19774 (n13608, n_9058, n13607);
  and g19775 (n13609, n_538, n10580);
  and g19776 (n13610, pi0116, n10585);
  not g19777 (n_9059, n13610);
  and g19778 (n13611, n_538, n_9059);
  and g19779 (n13612, n2924, n_6845);
  not g19780 (n_9060, n13612);
  and g19781 (n13613, pi0116, n_9060);
  not g19782 (n_9061, n13613);
  and g19783 (n13614, n_6848, n_9061);
  not g19784 (n_9062, n13611);
  not g19785 (n_9063, n13614);
  and g19786 (n13615, n_9062, n_9063);
  not g19787 (n_9064, n13609);
  and g19788 (n13616, pi0228, n_9064);
  not g19789 (n_9065, n13615);
  and g19790 (n13617, n_9065, n13616);
  and g19791 (n13618, pi0116, n10552);
  not g19792 (n_9066, n13618);
  and g19793 (n13619, n10777, n_9066);
  not g19794 (n_9067, n13619);
  and g19795 (n13620, n_162, n_9067);
  not g19796 (n_9068, n13617);
  and g19797 (n13621, n_9068, n13620);
  not g19798 (n_9069, n13621);
  and g19799 (n13622, n2608, n_9069);
  and g19800 (n13623, n_9018, n13597);
  and g19801 (n13624, n_3193, n13463);
  not g19802 (n_9070, n13624);
  and g19803 (n13625, n13597, n_9070);
  not g19804 (n_9071, n10502);
  not g19805 (n_9072, n13625);
  and g19806 (n13626, n_9071, n_9072);
  not g19807 (n_9073, n13626);
  and g19808 (n13627, n13467, n_9073);
  not g19809 (n_9074, n13623);
  not g19810 (n_9075, n13627);
  and g19811 (n13628, n_9074, n_9075);
  not g19812 (n_9076, n13628);
  and g19813 (n13629, n_162, n_9076);
  not g19814 (n_9077, n13629);
  and g19815 (n13630, n6285, n_9077);
  not g19821 (n_9080, n13608);
  and g19822 (n13634, n_171, n_9080);
  not g19823 (n_9081, n13633);
  and g19824 (n13635, n_9081, n13634);
  not g19825 (n_9082, n10497);
  and g19826 (n13636, n_9082, n13597);
  not g19827 (n_9083, n10738);
  not g19828 (n_9084, n13636);
  and g19829 (n13637, n_9083, n_9084);
  not g19830 (n_9085, n13637);
  and g19831 (n13638, n13467, n_9085);
  not g19832 (n_9086, n13638);
  and g19833 (n13639, n_9074, n_9086);
  not g19834 (n_9087, n13639);
  and g19835 (n13640, n2610, n_9087);
  and g19836 (n13641, n_6666, n13598);
  not g19837 (n_9088, n13641);
  and g19838 (n13642, pi0075, n_9088);
  not g19839 (n_9089, n13640);
  and g19840 (n13643, n_9089, n13642);
  not g19841 (n_9090, n13635);
  not g19842 (n_9091, n13643);
  and g19843 (n13644, n_9090, n_9091);
  not g19844 (n_9092, n13644);
  and g19845 (n13645, n8881, n_9092);
  and g19846 (n13646, n_8981, n_9050);
  not g19847 (n_9093, n13645);
  not g19848 (n_9094, n13646);
  and g19849 (po0274, n_9093, n_9094);
  and g19850 (n13648, n3686, n7379);
  not g19851 (n_9095, n13648);
  and g19852 (n13649, n_1088, n_9095);
  not g19853 (n_9096, n13649);
  and g19854 (n13650, n_161, n_9096);
  not g19855 (n_9097, n13650);
  and g19856 (n13651, n_172, n_9097);
  not g19857 (n_9098, n13651);
  and g19858 (n13652, n6133, n_9098);
  not g19859 (n_9099, n13652);
  and g19860 (n13653, n_174, n_9099);
  and g19861 (n13654, n_167, n_3994);
  and g19862 (n13655, n_168, n13654);
  not g19863 (n_9100, n13653);
  and g19864 (n13656, n_9100, n13655);
  not g19865 (n_9101, n13656);
  and g19866 (n13657, n_176, n_9101);
  not g19867 (n_9102, n13657);
  and g19868 (n13658, n_4025, n_9102);
  not g19869 (n_9103, n13658);
  and g19870 (n13659, n_157, n_9103);
  not g19871 (n_9104, n13659);
  and g19872 (n13660, n_3223, n_9104);
  not g19873 (n_9105, n13660);
  and g19874 (n13661, n_158, n_9105);
  and g19875 (n13662, n_796, n6300);
  not g19876 (n_9106, n13661);
  and g19877 (po0275, n_9106, n13662);
  and g19878 (n13664, n_5677, n12169);
  and g19879 (n13665, pi0163, n6197);
  not g19880 (n_9107, n13665);
  and g19881 (n13666, n_7621, n_9107);
  not g19882 (n_9109, pi0150);
  not g19883 (n_9110, n13666);
  and g19884 (n13667, n_9109, n_9110);
  and g19885 (n13668, pi0150, n9699);
  and g19886 (n13669, n11676, n13668);
  not g19887 (n_9111, n13667);
  not g19888 (n_9112, n13669);
  and g19889 (n13670, n_9111, n_9112);
  not g19890 (n_9113, n13670);
  and g19891 (n13671, pi0232, n_9113);
  and g19892 (n13672, n_6232, n13671);
  not g19893 (n_9114, n13672);
  and g19894 (n13673, pi0074, n_9114);
  and g19895 (n13674, pi0165, n7473);
  and g19896 (n13675, n_161, n_167);
  not g19897 (n_9116, n13674);
  not g19898 (n_9117, n13675);
  and g19899 (n13676, n_9116, n_9117);
  and g19900 (n13677, n8989, n13676);
  and g19901 (n13678, n_168, n_9114);
  not g19902 (n_9118, n13677);
  and g19903 (n13679, n_9118, n13678);
  not g19904 (n_9119, n13673);
  not g19905 (n_9120, n13679);
  and g19906 (n13680, n_9119, n_9120);
  not g19907 (n_9121, n13680);
  and g19908 (n13681, n_3243, n_9121);
  not g19909 (n_9122, n13681);
  and g19910 (n13682, n3328, n_9122);
  not g19911 (n_9123, n13682);
  and g19912 (n13683, n_6387, n_9123);
  and g19913 (n13684, pi0055, n_9119);
  and g19914 (n13685, pi0150, n7473);
  and g19915 (n13686, n_174, n9282);
  and g19916 (n13687, n13685, n13686);
  and g19917 (n13688, n9248, n13675);
  not g19918 (n_9124, n13687);
  and g19919 (n13689, n_9124, n13688);
  not g19920 (n_9125, n13676);
  not g19921 (n_9126, n13689);
  and g19922 (n13690, n_9125, n_9126);
  not g19923 (n_9127, n13690);
  and g19924 (n13691, n8989, n_9127);
  not g19925 (n_9128, n13691);
  and g19926 (n13692, n13678, n_9128);
  not g19927 (n_9129, n13692);
  and g19928 (n13693, n13684, n_9129);
  and g19929 (n13694, n_7617, n_7618);
  not g19930 (n_9131, n13694);
  and g19931 (n13695, pi0185, n_9131);
  not g19932 (n_9132, pi0185);
  and g19933 (n13696, n_9132, n13694);
  not g19934 (n_9133, n13695);
  and g19935 (n13697, n6197, n_9133);
  not g19936 (n_9134, n13696);
  and g19937 (n13698, n_9134, n13697);
  not g19938 (n_9135, n13698);
  and g19939 (n13699, n_234, n_9135);
  and g19940 (n13700, pi0299, n13670);
  not g19941 (n_9136, n13699);
  and g19942 (n13701, pi0232, n_9136);
  not g19943 (n_9137, n13700);
  and g19944 (n13702, n_9137, n13701);
  and g19945 (n13703, n_6232, n13702);
  not g19946 (n_9138, n13703);
  and g19947 (n13704, pi0074, n_9138);
  not g19948 (n_9139, n13704);
  and g19949 (n13705, n_176, n_9139);
  not g19950 (n_9141, pi0143);
  and g19951 (n13706, n_9141, n_234);
  not g19952 (n_9142, pi0165);
  and g19953 (n13707, n_9142, pi0299);
  not g19954 (n_9143, n13706);
  not g19955 (n_9144, n13707);
  and g19956 (n13708, n_9143, n_9144);
  and g19957 (n13709, n7473, n13708);
  not g19958 (n_9145, n13709);
  and g19959 (n13710, n8989, n_9145);
  not g19960 (n_9146, n13710);
  and g19961 (n13711, pi0054, n_9146);
  and g19962 (n13712, n_9138, n13711);
  not g19963 (n_9147, n13702);
  and g19964 (n13713, pi0075, n_9147);
  and g19965 (n13714, pi0100, n_9147);
  and g19966 (n13715, pi0038, n_9145);
  not g19967 (n_9148, n13715);
  and g19968 (n13716, n_164, n_9148);
  and g19969 (n13717, n_5686, pi0299);
  and g19970 (n13718, n_5708, n_234);
  not g19971 (n_9149, n13717);
  not g19972 (n_9150, n13718);
  and g19973 (n13719, n_9149, n_9150);
  and g19974 (n13720, n7473, n13719);
  and g19975 (n13721, n9282, n13720);
  not g19976 (n_9151, n13721);
  and g19977 (n13722, n9249, n_9151);
  not g19978 (n_9152, n13722);
  and g19979 (n13723, n13716, n_9152);
  not g19980 (n_9153, n13714);
  not g19981 (n_9154, n13723);
  and g19982 (n13724, n_9153, n_9154);
  not g19983 (n_9155, n13724);
  and g19984 (n13725, n9205, n_9155);
  and g19985 (n13726, n_9141, n_5815);
  and g19986 (n13727, pi0143, n_5817);
  not g19987 (n_9156, n13727);
  and g19988 (n13728, pi0165, n_9156);
  not g19989 (n_9157, n13726);
  and g19990 (n13729, n_9157, n13728);
  and g19991 (n13730, pi0143, n_9142);
  and g19992 (n13731, n9194, n13730);
  not g19993 (n_9158, n13731);
  and g19994 (n13732, pi0038, n_9158);
  not g19995 (n_9159, n13729);
  and g19996 (n13733, n_9159, n13732);
  not g19997 (n_9160, n13733);
  and g19998 (n13734, n2568, n_9160);
  and g19999 (n13735, n_3410, n9532);
  not g20000 (n_9161, n9532);
  and g20001 (n13736, n_3102, n_9161);
  and g20002 (n13737, n6197, n_6124);
  not g20003 (n_9162, n13736);
  not g20004 (n_9163, n13737);
  and g20005 (n13738, n_9162, n_9163);
  and g20006 (n13739, pi0151, pi0168);
  not g20007 (n_9164, n13738);
  and g20008 (n13740, n_9164, n13739);
  and g20009 (n13741, n_3102, n9532);
  and g20010 (n13742, pi0151, n_2206);
  and g20011 (n13743, n_6144, n13742);
  and g20012 (n13744, n_2206, n9615);
  and g20013 (n13745, pi0168, n9612);
  not g20014 (n_9165, n13744);
  and g20015 (n13746, n_983, n_9165);
  not g20016 (n_9166, n13745);
  and g20017 (n13747, n_9166, n13746);
  not g20018 (n_9167, n13743);
  not g20019 (n_9168, n13747);
  and g20020 (n13748, n_9167, n_9168);
  not g20021 (n_9169, n13741);
  not g20022 (n_9170, n13748);
  and g20023 (n13749, n_9169, n_9170);
  not g20024 (n_9171, n13740);
  and g20025 (n13750, pi0150, n_9171);
  not g20026 (n_9172, n13749);
  and g20027 (n13751, n_9172, n13750);
  and g20028 (n13752, pi0168, n6197);
  not g20029 (n_9173, n13752);
  and g20030 (n13753, n9532, n_9173);
  and g20031 (n13754, pi0168, n9506);
  not g20032 (n_9174, n13753);
  and g20033 (n13755, n_983, n_9174);
  not g20034 (n_9175, n13754);
  and g20035 (n13756, n_9175, n13755);
  and g20036 (n13757, n_6174, n_9162);
  and g20037 (n13758, n_2206, n13757);
  and g20038 (n13759, n_6175, n_9162);
  and g20039 (n13760, pi0168, n13759);
  not g20040 (n_9176, n13758);
  and g20041 (n13761, pi0151, n_9176);
  not g20042 (n_9177, n13760);
  and g20043 (n13762, n_9177, n13761);
  not g20044 (n_9178, n13756);
  and g20045 (n13763, n_9109, n_9178);
  not g20046 (n_9179, n13762);
  and g20047 (n13764, n_9179, n13763);
  not g20048 (n_9180, n13764);
  and g20049 (n13765, pi0299, n_9180);
  not g20050 (n_9181, n13751);
  and g20051 (n13766, n_9181, n13765);
  and g20052 (n13767, n_6064, n_9169);
  not g20053 (n_9183, pi0173);
  not g20054 (n_9184, n13767);
  and g20055 (n13768, n_9183, n_9184);
  and g20056 (n13769, pi0173, n13759);
  not g20057 (n_9185, n13768);
  and g20058 (n13770, n_9132, n_9185);
  not g20059 (n_9186, n13769);
  and g20060 (n13771, n_9186, n13770);
  and g20061 (n13772, n6197, n_6004);
  and g20062 (n13773, pi0173, n_9162);
  not g20063 (n_9187, n13772);
  and g20064 (n13774, n_9187, n13773);
  and g20065 (n13775, n_6059, n_9169);
  not g20066 (n_9188, n13775);
  and g20067 (n13776, n_9183, n_9188);
  not g20068 (n_9189, n13774);
  and g20069 (n13777, pi0185, n_9189);
  not g20070 (n_9190, n13776);
  and g20071 (n13778, n_9190, n13777);
  not g20072 (n_9192, n13771);
  and g20073 (n13779, pi0190, n_9192);
  not g20074 (n_9193, n13778);
  and g20075 (n13780, n_9193, n13779);
  and g20076 (n13781, n_9183, n_6081);
  and g20077 (n13782, pi0173, n_6440);
  not g20078 (n_9194, n13781);
  and g20079 (n13783, n6197, n_9194);
  not g20080 (n_9195, n13782);
  and g20081 (n13784, n_9195, n13783);
  and g20082 (n13785, pi0185, n_9169);
  not g20083 (n_9196, n13784);
  and g20084 (n13786, n_9196, n13785);
  and g20085 (n13787, pi0173, n13757);
  and g20086 (n13788, n_9183, n9532);
  not g20087 (n_9197, n13788);
  and g20088 (n13789, n_9132, n_9197);
  not g20089 (n_9198, n13787);
  and g20090 (n13790, n_9198, n13789);
  not g20091 (n_9199, pi0190);
  not g20092 (n_9200, n13790);
  and g20093 (n13791, n_9199, n_9200);
  not g20094 (n_9201, n13786);
  and g20095 (n13792, n_9201, n13791);
  not g20096 (n_9202, n13792);
  and g20097 (n13793, n_234, n_9202);
  not g20098 (n_9203, n13780);
  and g20099 (n13794, n_9203, n13793);
  not g20100 (n_9204, n13794);
  and g20101 (n13795, pi0232, n_9204);
  not g20102 (n_9205, n13766);
  and g20103 (n13796, n_9205, n13795);
  not g20104 (n_9206, n13735);
  and g20105 (n13797, n_162, n_9206);
  not g20106 (n_9207, n13796);
  and g20107 (n13798, n_9207, n13797);
  and g20108 (n13799, pi0168, n9311);
  and g20109 (n13800, pi0157, n9324);
  not g20110 (n_9208, n13799);
  not g20111 (n_9209, n13800);
  and g20112 (n13801, n_9208, n_9209);
  and g20113 (n13802, n6197, n11747);
  not g20114 (n_9210, n13801);
  and g20115 (n13803, n_9210, n13802);
  not g20116 (n_9211, n13803);
  and g20117 (n13804, pi0299, n_9211);
  not g20118 (n_9212, n13804);
  and g20119 (n13805, n_9150, n_9212);
  not g20120 (n_9213, n13805);
  and g20121 (n13806, n9248, n_9213);
  and g20122 (n13807, pi0178, n_6480);
  not g20123 (n_9214, n13807);
  and g20124 (n13808, n_9199, n_9214);
  not g20125 (n_9215, n13808);
  and g20126 (n13809, n_234, n_9215);
  not g20127 (n_9216, n13806);
  not g20128 (n_9217, n13809);
  and g20129 (n13810, n_9216, n_9217);
  and g20130 (n13811, n6205, n_5864);
  not g20131 (n_9218, n13811);
  and g20132 (n13812, n9051, n_9218);
  and g20133 (n13813, n_5708, n13812);
  not g20134 (n_9219, n9314);
  and g20135 (n13814, n_9219, n13813);
  and g20136 (n13815, n_234, n_5893);
  and g20137 (n13816, pi0178, n13812);
  not g20138 (n_9220, n9305);
  and g20139 (n13817, n_9220, n13816);
  not g20145 (n_9223, n13820);
  and g20146 (n13821, pi0232, n_9223);
  not g20147 (n_9224, n13810);
  and g20148 (n13822, n_9224, n13821);
  and g20149 (n13823, n_3410, n9248);
  not g20150 (n_9225, n13823);
  and g20151 (n13824, pi0039, n_9225);
  not g20152 (n_9226, n13822);
  and g20153 (n13825, n_9226, n13824);
  not g20154 (n_9227, n13825);
  and g20155 (n13826, n_161, n_9227);
  not g20156 (n_9228, n13798);
  and g20157 (n13827, n_9228, n13826);
  not g20158 (n_9229, n13827);
  and g20159 (n13828, n13734, n_9229);
  and g20160 (n13829, n8161, n_9148);
  not g20161 (n_9230, n9249);
  and g20162 (n13830, n_9230, n13829);
  not g20163 (n_9231, n13830);
  and g20164 (n13831, n_9153, n_9231);
  not g20165 (n_9232, n13828);
  and g20166 (n13832, n_9232, n13831);
  not g20167 (n_9233, n13832);
  and g20168 (n13833, n2569, n_9233);
  not g20169 (n_9234, n13713);
  not g20170 (n_9235, n13725);
  and g20171 (n13834, n_9234, n_9235);
  not g20172 (n_9236, n13833);
  and g20173 (n13835, n_9236, n13834);
  not g20174 (n_9237, n13835);
  and g20175 (n13836, n_167, n_9237);
  not g20176 (n_9238, n13712);
  not g20177 (n_9239, n13836);
  and g20178 (n13837, n_9238, n_9239);
  not g20179 (n_9240, n13837);
  and g20180 (n13838, n_168, n_9240);
  not g20181 (n_9241, n13838);
  and g20182 (n13839, n13705, n_9241);
  not g20183 (n_9242, n13693);
  and g20184 (n13840, n2529, n_9242);
  not g20185 (n_9243, n13839);
  and g20186 (n13841, n_9243, n13840);
  not g20187 (n_9244, n13683);
  not g20188 (n_9245, n13841);
  and g20189 (n13842, n_9244, n_9245);
  and g20190 (n13843, n8989, n13674);
  not g20191 (n_9246, n13671);
  and g20192 (n13844, n_6232, n_9246);
  not g20198 (n_9249, n13842);
  not g20199 (n_9250, n13847);
  and g20200 (n13848, n_9249, n_9250);
  and g20201 (n13849, pi0118, n13848);
  not g20202 (n_9251, n13720);
  and g20203 (n13850, n8965, n_9251);
  and g20204 (n13851, n2521, n13850);
  not g20205 (n_9252, n13851);
  and g20206 (n13852, n13716, n_9252);
  not g20207 (n_9253, n13852);
  and g20208 (n13853, n_9153, n_9253);
  not g20209 (n_9254, n13853);
  and g20210 (n13854, n9205, n_9254);
  and g20211 (n13855, n7309, n9061);
  and g20212 (n13856, n_3164, n13130);
  and g20213 (n13857, n_3284, n13856);
  not g20214 (n_9255, n13857);
  and g20215 (n13858, n_3410, n_9255);
  not g20216 (n_9256, n13855);
  and g20217 (n13859, n_9256, n13858);
  and g20218 (n13860, n6198, n_3284);
  and g20219 (n13861, pi0157, n_5734);
  and g20220 (n13862, n_5686, n9044);
  not g20221 (n_9257, n13862);
  and g20222 (n13863, pi0168, n_9257);
  and g20223 (n13864, n_5686, n_2206);
  and g20224 (n13865, n_5733, n13864);
  not g20225 (n_9258, n13861);
  not g20226 (n_9259, n13865);
  and g20227 (n13866, n_9258, n_9259);
  not g20228 (n_9260, n13863);
  and g20229 (n13867, n_9260, n13866);
  not g20230 (n_9261, n13860);
  not g20231 (n_9262, n13867);
  and g20232 (n13868, n_9261, n_9262);
  not g20233 (n_9263, n13868);
  and g20234 (n13869, n13130, n_9263);
  and g20235 (n13870, n_5708, n_3119);
  and g20236 (n13871, n9043, n13870);
  not g20237 (n_9264, n13871);
  and g20238 (n13872, n_9261, n_9264);
  not g20239 (n_9265, n13872);
  and g20240 (n13873, pi0190, n_9265);
  not g20241 (n_9266, n9052);
  and g20242 (n13874, pi0178, n_9266);
  and g20243 (n13875, n_9261, n13874);
  not g20244 (n_9267, n13173);
  and g20245 (n13876, n_5708, n_9267);
  not g20246 (n_9268, n13875);
  and g20247 (n13877, n_9199, n_9268);
  not g20248 (n_9269, n13876);
  and g20249 (n13878, n_9269, n13877);
  not g20250 (n_9270, n13873);
  not g20251 (n_9271, n13878);
  and g20252 (n13879, n_9270, n_9271);
  not g20253 (n_9272, n13879);
  and g20254 (n13880, n13132, n_9272);
  not g20255 (n_9273, n13880);
  and g20256 (n13881, pi0232, n_9273);
  not g20257 (n_9274, n13869);
  and g20258 (n13882, n_9274, n13881);
  not g20259 (n_9275, n13859);
  and g20260 (n13883, pi0039, n_9275);
  not g20261 (n_9276, n13882);
  and g20262 (n13884, n_9276, n13883);
  and g20263 (n13885, n_3066, n_5770);
  and g20264 (n13886, n_3410, n_5771);
  not g20265 (n_9277, n13885);
  and g20266 (n13887, n_9277, n13886);
  and g20267 (n13888, n_5771, n_7681);
  not g20268 (n_9278, n13888);
  and g20269 (n13889, n_3102, n_9278);
  and g20270 (n13890, n9142, n13742);
  and g20271 (n13891, pi0168, n_7708);
  and g20272 (n13892, n_2206, n_7709);
  not g20273 (n_9279, n13891);
  and g20274 (n13893, n_983, n_9279);
  not g20275 (n_9280, n13892);
  and g20276 (n13894, n_9280, n13893);
  not g20277 (n_9281, n13890);
  not g20278 (n_9282, n13894);
  and g20279 (n13895, n_9281, n_9282);
  not g20280 (n_9283, n13895);
  and g20281 (n13896, n9094, n_9283);
  not g20282 (n_9284, n13896);
  and g20283 (n13897, pi0150, n_9284);
  and g20284 (n13898, n_983, n9129);
  not g20285 (n_9285, n13898);
  and g20286 (n13899, n9166, n_9285);
  not g20287 (n_9286, n13899);
  and g20288 (n13900, n13752, n_9286);
  and g20289 (n13901, n_983, n9118);
  not g20290 (n_9287, n13901);
  and g20291 (n13902, n9162, n_9287);
  not g20292 (n_9288, n13902);
  and g20293 (n13903, n_2206, n_9288);
  not g20294 (n_9289, n13900);
  and g20295 (n13904, n_9109, n_9289);
  not g20296 (n_9290, n13903);
  and g20297 (n13905, n_9290, n13904);
  not g20298 (n_9291, n13897);
  not g20299 (n_9292, n13905);
  and g20300 (n13906, n_9291, n_9292);
  not g20301 (n_9293, n13889);
  and g20302 (n13907, pi0299, n_9293);
  not g20303 (n_9294, n13906);
  and g20304 (n13908, n_9294, n13907);
  and g20305 (n13909, n_3102, n_5773);
  and g20306 (n13910, n6479, n9142);
  and g20307 (n13911, pi0173, n13910);
  and g20308 (n13912, n_9183, n6479);
  and g20309 (n13913, n9092, n13912);
  not g20310 (n_9295, n13911);
  not g20311 (n_9296, n13913);
  and g20312 (n13914, n_9295, n_9296);
  and g20313 (n13915, n_9199, n6197);
  not g20314 (n_9297, n13914);
  and g20315 (n13916, n_9297, n13915);
  and g20316 (n13917, n_9183, pi0190);
  and g20317 (n13918, n9134, n13917);
  not g20318 (n_9298, n13918);
  and g20319 (n13919, pi0185, n_9298);
  not g20320 (n_9299, n13916);
  and g20321 (n13920, n_9299, n13919);
  and g20322 (n13921, pi0173, n9150);
  and g20323 (n13922, pi0190, n9131);
  not g20324 (n_9300, n13921);
  and g20325 (n13923, n_9300, n13922);
  and g20326 (n13924, n_9183, n9118);
  not g20327 (n_9301, n13924);
  and g20328 (n13925, n9147, n_9301);
  not g20329 (n_9302, n13925);
  and g20330 (n13926, n_9199, n_9302);
  not g20331 (n_9303, n13923);
  and g20332 (n13927, n_9132, n_9303);
  not g20333 (n_9304, n13926);
  and g20334 (n13928, n_9304, n13927);
  not g20335 (n_9305, n13920);
  not g20336 (n_9306, n13928);
  and g20337 (n13929, n_9305, n_9306);
  not g20338 (n_9307, n13909);
  and g20339 (n13930, n_234, n_9307);
  not g20340 (n_9308, n13929);
  and g20341 (n13931, n_9308, n13930);
  not g20342 (n_9309, n13908);
  not g20343 (n_9310, n13931);
  and g20344 (n13932, n_9309, n_9310);
  not g20345 (n_9311, n13932);
  and g20346 (n13933, pi0232, n_9311);
  not g20347 (n_9312, n13887);
  and g20348 (n13934, n_162, n_9312);
  not g20349 (n_9313, n13933);
  and g20350 (n13935, n_9313, n13934);
  not g20351 (n_9314, n13884);
  not g20352 (n_9315, n13935);
  and g20353 (n13936, n_9314, n_9315);
  not g20354 (n_9316, n13936);
  and g20355 (n13937, n_161, n_9316);
  not g20356 (n_9317, n13937);
  and g20357 (n13938, n13734, n_9317);
  not g20358 (n_9318, n13829);
  and g20359 (n13939, n_9153, n_9318);
  not g20360 (n_9319, n13938);
  and g20361 (n13940, n_9319, n13939);
  not g20362 (n_9320, n13940);
  and g20363 (n13941, n2569, n_9320);
  not g20364 (n_9321, n13854);
  and g20365 (n13942, n_9234, n_9321);
  not g20366 (n_9322, n13941);
  and g20367 (n13943, n_9322, n13942);
  not g20368 (n_9323, n13943);
  and g20369 (n13944, n_167, n_9323);
  not g20370 (n_9324, n13944);
  and g20371 (n13945, n_9238, n_9324);
  not g20372 (n_9325, n13945);
  and g20373 (n13946, n_168, n_9325);
  not g20374 (n_9326, n13946);
  and g20375 (n13947, n13705, n_9326);
  and g20376 (n13948, pi0054, n13674);
  not g20379 (n_9327, n13685);
  not g20384 (n_9329, n13953);
  and g20385 (n13954, n13679, n_9329);
  not g20386 (n_9330, n13954);
  and g20387 (n13955, n13684, n_9330);
  not g20388 (n_9331, n13955);
  and g20389 (n13956, n2529, n_9331);
  not g20390 (n_9332, n13947);
  and g20391 (n13957, n_9332, n13956);
  not g20392 (n_9333, n13957);
  and g20393 (n13958, n13682, n_9333);
  not g20394 (n_9334, n13958);
  and g20395 (n13959, n_9250, n_9334);
  and g20396 (n13960, n_5675, n13959);
  not g20397 (n_9335, n13664);
  not g20398 (n_9336, n13960);
  and g20399 (n13961, n_9335, n_9336);
  not g20400 (n_9337, n13849);
  and g20401 (n13962, n_9337, n13961);
  not g20402 (n_9338, n8976);
  and g20403 (n13963, n_5675, n_9338);
  not g20404 (n_9339, n13963);
  and g20405 (n13964, n13959, n_9339);
  and g20406 (n13965, n13848, n13963);
  not g20407 (n_9340, n13964);
  and g20408 (n13966, n13664, n_9340);
  not g20409 (n_9341, n13965);
  and g20410 (n13967, n_9341, n13966);
  or g20411 (po0276, n13962, n13967);
  and g20412 (n13969, pi0128, pi0228);
  not g20413 (n_9343, n10163);
  and g20414 (n13970, n_9343, n13969);
  and g20415 (n13971, n7384, n8965);
  not g20416 (n_9344, n13969);
  not g20417 (n_9345, n13971);
  and g20418 (n13972, n_9344, n_9345);
  not g20419 (n_9346, n13972);
  and g20420 (n13973, pi0075, n_9346);
  and g20421 (n13974, pi0087, n_9344);
  and g20422 (n13975, n2530, n3335);
  not g20423 (n_9347, n13975);
  and g20424 (n13976, n_9344, n_9347);
  not g20425 (n_9348, n13976);
  and g20426 (n13977, pi0100, n_9348);
  not g20427 (n_9349, n2603);
  and g20428 (n13978, n_9349, n3470);
  and g20429 (n13979, n7606, n13978);
  not g20430 (n_9350, n3448);
  and g20431 (n13980, n_9350, n5853);
  and g20432 (n13981, n7603, n13980);
  not g20433 (n_9351, n13979);
  not g20434 (n_9352, n13981);
  and g20435 (n13982, n_9351, n_9352);
  not g20436 (n_9353, n13982);
  and g20437 (n13983, pi0039, n_9353);
  and g20438 (n13984, pi0299, n6418);
  not g20439 (n_9354, n13984);
  and g20440 (n13985, n_3397, n_9354);
  not g20441 (n_9355, n13985);
  and g20442 (n13986, n7473, n_9355);
  not g20443 (n_9356, n13986);
  and g20444 (n13987, pi0109, n_9356);
  and g20445 (n13988, n_494, n11668);
  and g20446 (n13989, n2770, n10157);
  not g20447 (n_9357, n13989);
  and g20448 (n13990, n11667, n_9357);
  not g20449 (n_9358, n13990);
  and g20450 (n13991, n2783, n_9358);
  not g20451 (n_9359, n13991);
  and g20452 (n13992, n_122, n_9359);
  not g20457 (n_9361, n13987);
  not g20458 (n_9362, n13988);
  and g20459 (n13996, n_9361, n_9362);
  not g20460 (n_9363, n13995);
  and g20461 (n13997, n_9363, n13996);
  not g20462 (n_9364, n6422);
  and g20463 (n13998, n_9364, n_9356);
  not g20464 (n_9365, n6491);
  and g20465 (n13999, n_9365, n13986);
  not g20466 (n_9366, n13998);
  not g20467 (n_9367, n13999);
  and g20468 (n14000, n_9366, n_9367);
  not g20469 (n_9368, n13997);
  and g20470 (n14001, n_9368, n14000);
  not g20471 (n_9369, n14001);
  and g20472 (n14002, n_109, n_9369);
  and g20473 (n14003, n2938, n_3308);
  not g20474 (n_9370, n14002);
  and g20475 (n14004, n_9370, n14003);
  not g20476 (n_9371, n14004);
  and g20477 (n14005, n_352, n_9371);
  and g20478 (n14006, n_162, n11086);
  not g20479 (n_9372, n14005);
  and g20480 (n14007, n_9372, n14006);
  not g20481 (n_9373, n13983);
  not g20482 (n_9374, n14007);
  and g20483 (n14008, n_9373, n_9374);
  not g20484 (n_9375, n14008);
  and g20485 (n14009, n_161, n_9375);
  and g20486 (n14010, n_188, n14009);
  not g20487 (n_9376, n14010);
  and g20488 (n14011, n_9344, n_9376);
  not g20489 (n_9377, n14011);
  and g20490 (n14012, n_164, n_9377);
  not g20491 (n_9378, n13977);
  and g20492 (n14013, n_172, n_9378);
  not g20493 (n_9379, n14012);
  and g20494 (n14014, n_9379, n14013);
  not g20495 (n_9380, n13974);
  and g20496 (n14015, n_171, n_9380);
  not g20497 (n_9381, n14014);
  and g20498 (n14016, n_9381, n14015);
  not g20499 (n_9382, n13973);
  and g20500 (n14017, n_174, n_9382);
  not g20501 (n_9383, n14016);
  and g20502 (n14018, n_9383, n14017);
  and g20503 (n14019, pi0092, n_9344);
  and g20504 (n14020, n_4041, n14019);
  not g20505 (n_9384, n14020);
  and g20506 (n14021, n10163, n_9384);
  not g20507 (n_9385, n14018);
  and g20508 (n14022, n_9385, n14021);
  or g20509 (po0277, n13970, n14022);
  and g20510 (n14024, n_5629, n_7977);
  and g20511 (n14025, pi0818, n14024);
  and g20512 (n14026, n7420, n_4196);
  not g20513 (n_9387, n14026);
  and g20514 (n14027, n_4091, n_9387);
  not g20515 (n_9389, pi0120);
  and g20516 (n14028, n_9389, n_4196);
  and g20517 (n14029, n_3206, n14028);
  not g20518 (n_9390, n14029);
  and g20519 (n14030, n14027, n_9390);
  and g20520 (n14031, pi0120, n_8134);
  and g20521 (n14032, n_9389, pi1093);
  and g20522 (n14033, n_3128, n12310);
  not g20523 (n_9391, n14033);
  and g20524 (n14034, n14032, n_9391);
  not g20525 (n_9392, n14031);
  not g20526 (n_9393, n14034);
  and g20527 (n14035, n_9392, n_9393);
  and g20528 (n14036, n2521, n7595);
  not g20529 (n_9394, n7619);
  and g20530 (n14037, n_9394, n14031);
  not g20531 (n_9395, n14037);
  and g20532 (n14038, n14036, n_9395);
  not g20533 (n_9396, n14032);
  and g20534 (n14039, n7619, n_9396);
  not g20535 (n_9397, n14038);
  not g20536 (n_9398, n14039);
  and g20537 (n14040, n_9397, n_9398);
  and g20538 (n14041, n2530, n7506);
  not g20539 (n_9399, n14040);
  and g20540 (n14042, n_9399, n14041);
  not g20541 (n_9400, n14035);
  and g20542 (n14043, pi0100, n_9400);
  not g20543 (n_9401, n14042);
  and g20544 (n14044, n_9401, n14043);
  and g20545 (n14045, pi0038, n7420);
  and g20546 (n14046, n_3206, n7460);
  and g20547 (n14047, pi0120, n14046);
  not g20548 (n_9402, n14047);
  and g20549 (n14048, n_162, n_9402);
  not g20550 (n_9403, n7452);
  and g20551 (n14049, pi0122, n_9403);
  and g20552 (n14050, n7534, n_6757);
  and g20553 (n14051, n7417, n7451);
  and g20554 (n14052, n_3127, n14051);
  not g20555 (n_9404, n14052);
  and g20556 (n14053, n_4081, n_9404);
  not g20557 (n_9405, n14050);
  and g20558 (n14054, n_9405, n14053);
  not g20559 (n_9406, n14049);
  and g20560 (n14055, n_489, n_9406);
  not g20561 (n_9407, n14054);
  and g20562 (n14056, n_9407, n14055);
  not g20563 (n_9408, n14056);
  and g20564 (n14057, n2930, n_9408);
  not g20565 (n_9409, n14051);
  and g20566 (n14058, n7626, n_9409);
  and g20567 (n14059, n_8085, n14058);
  not g20568 (n_9410, n14057);
  not g20569 (n_9411, n14059);
  and g20570 (n14060, n_9410, n_9411);
  and g20571 (n14061, n14048, n14060);
  and g20572 (n14062, n_4176, n14035);
  and g20573 (n14063, n_3120, n14035);
  not g20574 (n_9412, n7602);
  and g20575 (n14064, n_9412, n14031);
  and g20576 (n14065, pi1091, pi1092);
  and g20577 (n14066, n7554, n14065);
  not g20578 (n_9413, n14066);
  and g20579 (n14067, n14034, n_9413);
  not g20580 (n_9414, n14064);
  not g20581 (n_9415, n14067);
  and g20582 (n14068, n_9414, n_9415);
  and g20583 (n14069, n6198, n14068);
  not g20584 (n_9416, n14063);
  not g20585 (n_9417, n14069);
  and g20586 (n14070, n_9416, n_9417);
  and g20587 (n14071, n6242, n14070);
  and g20588 (n14072, n6227, n_9400);
  not g20589 (n_9418, n14068);
  and g20590 (n14073, n_3140, n_9418);
  not g20591 (n_9419, n14072);
  not g20592 (n_9420, n14073);
  and g20593 (n14074, n_9419, n_9420);
  not g20594 (n_9421, n14074);
  and g20595 (n14075, n_3162, n_9421);
  not g20596 (n_9422, n14071);
  and g20597 (n14076, n7570, n_9422);
  not g20598 (n_9423, n14075);
  and g20599 (n14077, n_9423, n14076);
  not g20600 (n_9424, n14062);
  and g20601 (n14078, pi0299, n_9424);
  not g20602 (n_9425, n14077);
  and g20603 (n14079, n_9425, n14078);
  and g20604 (n14080, n6205, n14070);
  and g20605 (n14081, n_3119, n_9421);
  not g20606 (n_9426, n14080);
  and g20607 (n14082, n7551, n_9426);
  not g20608 (n_9427, n14081);
  and g20609 (n14083, n_9427, n14082);
  and g20610 (n14084, n_4165, n14035);
  not g20611 (n_9428, n14084);
  and g20612 (n14085, n_234, n_9428);
  not g20613 (n_9429, n14083);
  and g20614 (n14086, n_9429, n14085);
  not g20615 (n_9430, n14079);
  and g20616 (n14087, pi0039, n_9430);
  not g20617 (n_9431, n14086);
  and g20618 (n14088, n_9431, n14087);
  not g20619 (n_9432, n14061);
  not g20620 (n_9433, n14088);
  and g20621 (n14089, n_9432, n_9433);
  not g20622 (n_9434, n14089);
  and g20623 (n14090, n_161, n_9434);
  and g20624 (n14091, n_9389, n_3206);
  and g20625 (n14092, pi0038, n14091);
  not g20626 (n_9435, n14092);
  and g20627 (n14093, n_164, n_9435);
  not g20628 (n_9436, n14045);
  and g20629 (n14094, n_9436, n14093);
  not g20630 (n_9437, n14090);
  and g20631 (n14095, n_9437, n14094);
  not g20632 (n_9438, n14044);
  not g20633 (n_9439, n14095);
  and g20634 (n14096, n_9438, n_9439);
  not g20635 (n_9440, n14096);
  and g20636 (n14097, n_172, n_9440);
  not g20637 (n_9441, n14091);
  and g20638 (n14098, n7631, n_9441);
  and g20639 (n14099, n_251, n7420);
  and g20640 (n14100, n7626, n_8085);
  and g20641 (n14101, n_4128, n14100);
  not g20642 (n_9442, n14101);
  and g20643 (n14102, n7629, n_9442);
  not g20644 (n_9443, n14099);
  and g20645 (n14103, pi0087, n_9443);
  not g20646 (n_9444, n14102);
  and g20647 (n14104, n_9444, n14103);
  and g20648 (n14105, n14098, n14104);
  not g20649 (n_9445, n14097);
  not g20650 (n_9446, n14105);
  and g20651 (n14106, n_9445, n_9446);
  not g20652 (n_9447, n14106);
  and g20653 (n14107, n_171, n_9447);
  and g20654 (n14108, n7474, n14035);
  not g20655 (n_9448, n7596);
  and g20656 (n14109, n_9448, n14034);
  not g20657 (n_9449, n7419);
  and g20658 (n14110, n_3128, n_9449);
  not g20659 (n_9450, n14110);
  and g20660 (n14111, n_4121, n_9450);
  not g20661 (n_9451, n14111);
  and g20662 (n14112, pi0120, n_9451);
  not g20663 (n_9452, n14112);
  and g20664 (n14113, n_4117, n_9452);
  not g20665 (n_9453, n14109);
  and g20666 (n14114, n_9453, n14113);
  not g20667 (n_9454, n14108);
  not g20668 (n_9455, n14114);
  and g20669 (n14115, n_9454, n_9455);
  not g20670 (n_9456, n14115);
  and g20671 (n14116, n2610, n_9456);
  and g20672 (n14117, n_766, n14035);
  not g20673 (n_9457, n14117);
  and g20674 (n14118, pi0075, n_9457);
  not g20675 (n_9458, n14116);
  and g20676 (n14119, n_9458, n14118);
  not g20677 (n_9459, n14119);
  and g20678 (n14120, n7429, n_9459);
  not g20679 (n_9460, n14107);
  and g20680 (n14121, n_9460, n14120);
  not g20681 (n_9461, n14121);
  and g20682 (n14122, n14030, n_9461);
  and g20683 (n14123, n7599, n_9441);
  not g20684 (n_9462, n14058);
  and g20685 (n14124, n_9410, n_9462);
  and g20686 (n14125, n14048, n14124);
  and g20687 (n14126, pi1093, n_3120);
  and g20688 (n14127, n6242, n14126);
  and g20689 (n14128, n6227, n_3162);
  and g20695 (n14132, pi0299, n_9441);
  not g20696 (n_9465, n14131);
  and g20697 (n14133, n_9465, n14132);
  and g20698 (n14134, n6205, n14126);
  and g20699 (n14135, n_3119, n6227);
  and g20705 (n14139, n_234, n_9441);
  not g20706 (n_9468, n14138);
  and g20707 (n14140, n_9468, n14139);
  not g20708 (n_9469, n14133);
  and g20709 (n14141, pi0039, n_9469);
  not g20710 (n_9470, n14140);
  and g20711 (n14142, n_9470, n14141);
  not g20712 (n_9471, n14125);
  not g20713 (n_9472, n14142);
  and g20714 (n14143, n_9471, n_9472);
  not g20715 (n_9473, n14143);
  and g20716 (n14144, n_161, n_9473);
  not g20717 (n_9474, n14144);
  and g20718 (n14145, n14093, n_9474);
  and g20719 (n14146, pi0120, n7619);
  and g20720 (n14147, n_9389, n14036);
  not g20721 (n_9475, n14146);
  not g20722 (n_9476, n14147);
  and g20723 (n14148, n_9475, n_9476);
  not g20724 (n_9477, n14148);
  and g20725 (n14149, n14041, n_9477);
  and g20726 (n14150, pi0100, n_9441);
  not g20727 (n_9478, n14149);
  and g20728 (n14151, n_9478, n14150);
  not g20729 (n_9479, n14145);
  not g20730 (n_9480, n14151);
  and g20731 (n14152, n_9479, n_9480);
  not g20732 (n_9481, n14152);
  and g20733 (n14153, n_172, n_9481);
  not g20734 (n_9482, n14098);
  not g20735 (n_9483, n14153);
  and g20736 (n14154, n_9482, n_9483);
  not g20737 (n_9484, n14154);
  and g20738 (n14155, n_171, n_9484);
  not g20739 (n_9485, n14123);
  and g20740 (n14156, n7429, n_9485);
  not g20741 (n_9486, n14155);
  and g20742 (n14157, n_9486, n14156);
  and g20743 (n14158, n7425, n_9390);
  not g20744 (n_9487, n14157);
  and g20745 (n14159, n_9487, n14158);
  not g20746 (n_9488, n14122);
  not g20747 (n_9489, n14159);
  and g20748 (n14160, n_9488, n_9489);
  not g20749 (n_9490, n14160);
  and g20750 (n14161, n14025, n_9490);
  not g20751 (n_9491, n14161);
  and g20752 (n14162, n_4226, n_9491);
  and g20753 (n14163, n_4091, n14035);
  not g20754 (n_9492, n14163);
  and g20755 (n14164, pi0120, n_9492);
  and g20756 (n14165, n14025, n_9441);
  and g20757 (n14166, n_9492, n14165);
  not g20758 (n_9493, n14166);
  and g20759 (n14167, po1038, n_9493);
  not g20760 (n_9494, n14164);
  and g20761 (n14168, n_9494, n14167);
  not g20762 (n_9495, n7643);
  not g20763 (n_9496, n14168);
  and g20764 (n14169, n_9495, n_9496);
  and g20765 (n14170, pi0951, pi0982);
  and g20766 (n14171, pi1092, n14170);
  and g20767 (n14172, pi1093, n14171);
  not g20768 (n_9499, n14172);
  and g20769 (n14173, n_9389, n_9499);
  not g20770 (n_9500, n14173);
  and g20771 (n14174, n_9492, n_9500);
  not g20772 (n_9501, n14174);
  and g20773 (n14175, n14167, n_9501);
  not g20774 (n_9502, n14175);
  and g20775 (n14176, n7643, n_9502);
  not g20776 (n_9503, n14169);
  not g20777 (n_9504, n14176);
  and g20778 (n14177, n_9503, n_9504);
  not g20779 (n_9505, n14162);
  not g20780 (n_9506, n14177);
  and g20781 (n14178, n_9505, n_9506);
  and g20782 (n14179, n14028, n_9499);
  and g20783 (n14180, n_766, n_9500);
  and g20784 (n14181, pi0120, n7597);
  and g20785 (n14182, n_3128, n14172);
  not g20786 (n_9507, n14182);
  and g20787 (n14183, n_9389, n_9507);
  and g20788 (n14184, n2930, n14171);
  not g20797 (n_9508, n14192);
  and g20798 (n14193, n14184, n_9508);
  not g20799 (n_9509, n14193);
  and g20800 (n14194, n14183, n_9509);
  not g20801 (n_9510, n14181);
  not g20802 (n_9511, n14194);
  and g20803 (n14195, n_9510, n_9511);
  not g20804 (n_9512, n14195);
  and g20805 (n14196, n_4117, n_9512);
  and g20806 (n14197, n7474, n14173);
  not g20807 (n_9513, n14197);
  and g20808 (n14198, n2610, n_9513);
  not g20809 (n_9514, n14196);
  and g20810 (n14199, n_9514, n14198);
  not g20811 (n_9515, n14180);
  and g20812 (n14200, pi0075, n_9515);
  not g20813 (n_9516, n14199);
  and g20814 (n14201, n_9516, n14200);
  and g20815 (n14202, n_251, n14173);
  not g20816 (n_9517, n14202);
  and g20817 (n14203, pi0087, n_9517);
  and g20818 (n14204, pi0950, n2521);
  and g20819 (n14205, n_489, n_3130);
  and g20820 (n14206, n14204, n14205);
  not g20821 (n_9518, n14206);
  and g20822 (n14207, n14184, n_9518);
  and g20823 (n14208, pi0824, n14204);
  not g20824 (n_9519, n14208);
  and g20825 (n14209, n14182, n_9519);
  not g20826 (n_9520, n14207);
  not g20827 (n_9521, n14209);
  and g20828 (n14210, n_9520, n_9521);
  not g20829 (n_9522, n14210);
  and g20830 (n14211, n_9389, n_9522);
  and g20831 (n14212, n_4216, n_4215);
  not g20832 (n_9523, n14212);
  and g20833 (n14213, pi0120, n_9523);
  not g20834 (n_9524, n14213);
  and g20835 (n14214, n2625, n_9524);
  not g20836 (n_9525, n14211);
  and g20837 (n14215, n_9525, n14214);
  not g20838 (n_9526, n14215);
  and g20839 (n14216, n14203, n_9526);
  and g20840 (n14217, n7430, n7478);
  and g20841 (n14218, n14204, n14217);
  not g20842 (n_9527, n14218);
  and g20843 (n14219, n14184, n_9527);
  not g20844 (n_9528, n14219);
  and g20845 (n14220, n14183, n_9528);
  not g20846 (n_9529, n14220);
  and g20847 (n14221, n_9475, n_9529);
  and g20848 (n14222, n_162, n7506);
  not g20849 (n_9530, n14221);
  and g20850 (n14223, n_9530, n14222);
  not g20851 (n_9531, n14223);
  and g20852 (n14224, pi0100, n_9531);
  not g20853 (n_9532, n14224);
  and g20854 (n14225, n_161, n_9532);
  not g20855 (n_9533, n14041);
  and g20856 (n14226, n_9533, n14173);
  not g20857 (n_9534, n14225);
  not g20858 (n_9535, n14226);
  and g20859 (n14227, n_9534, n_9535);
  and g20860 (n14228, n_4165, n14173);
  not g20861 (n_9536, n14228);
  and g20862 (n14229, n_234, n_9536);
  and g20863 (n14230, n_5400, n_9500);
  and g20864 (n14231, n_3119, n14230);
  and g20865 (n14232, n_5401, n_9500);
  and g20866 (n14233, n6205, n14232);
  not g20867 (n_9537, n14231);
  and g20868 (n14234, n7551, n_9537);
  not g20869 (n_9538, n14233);
  and g20870 (n14235, n_9538, n14234);
  not g20871 (n_9539, n14235);
  and g20872 (n14236, n14229, n_9539);
  and g20873 (n14237, n_4176, n14173);
  not g20874 (n_9540, n14237);
  and g20875 (n14238, pi0299, n_9540);
  and g20876 (n14239, n_3162, n14230);
  and g20877 (n14240, n6242, n14232);
  not g20878 (n_9541, n14239);
  and g20879 (n14241, n7570, n_9541);
  not g20880 (n_9542, n14240);
  and g20881 (n14242, n_9542, n14241);
  not g20882 (n_9543, n14242);
  and g20883 (n14243, n14238, n_9543);
  not g20884 (n_9544, n14236);
  not g20885 (n_9545, n14243);
  and g20886 (n14244, n_9544, n_9545);
  not g20887 (n_9546, n14244);
  and g20888 (n14245, pi0039, n_9546);
  and g20889 (n14246, n2771, n7437);
  and g20890 (n14247, n2767, n14246);
  and g20891 (n14248, n9110, n14247);
  and g20892 (n14249, n7431, n14248);
  not g20893 (n_9547, n14249);
  and g20894 (n14250, n7436, n_9547);
  and g20895 (n14251, pi0950, n7518);
  not g20896 (n_9548, n14250);
  and g20897 (n14252, n_9548, n14251);
  and g20898 (n14253, pi0824, n14252);
  not g20899 (n_9549, n14253);
  and g20900 (n14254, n14171, n_9549);
  and g20901 (n14255, n_3127, n14254);
  not g20902 (n_9550, n14247);
  and g20903 (n14256, n_122, n_9550);
  not g20904 (n_9551, n14256);
  and g20905 (n14257, n2935, n_9551);
  and g20906 (n14258, n2937, n14257);
  not g20907 (n_9552, n14258);
  and g20908 (n14259, n_4146, n_9552);
  not g20909 (n_9553, n14259);
  and g20910 (n14260, n2461, n_9553);
  not g20911 (n_9554, n14260);
  and g20912 (n14261, n7434, n_9554);
  not g20913 (n_9555, n14261);
  and g20914 (n14262, n7431, n_9555);
  not g20915 (n_9556, n14262);
  and g20916 (n14263, n_138, n_9556);
  not g20917 (n_9557, n14263);
  and g20918 (n14264, n_350, n_9557);
  not g20919 (n_9558, n14264);
  and g20920 (n14265, n_135, n_9558);
  and g20925 (n14269, n7430, n14171);
  not g20926 (n_9560, n14268);
  and g20927 (n14270, n_9560, n14269);
  and g20928 (n14271, pi0829, pi1092);
  not g20933 (n_9562, n14255);
  not g20934 (n_9563, n14274);
  and g20935 (n14275, n_9562, n_9563);
  not g20936 (n_9564, n14270);
  and g20937 (n14276, n_9564, n14275);
  not g20938 (n_9565, n14276);
  and g20939 (n14277, n7517, n_9565);
  and g20940 (n14278, n2923, n14172);
  not g20941 (n_9566, n14277);
  not g20942 (n_9567, n14278);
  and g20943 (n14279, n_9566, n_9567);
  not g20944 (n_9568, n14279);
  and g20945 (n14280, pi1091, n_9568);
  and g20946 (n14281, n14182, n_9549);
  not g20947 (n_9569, n14281);
  and g20948 (n14282, n_9389, n_9569);
  not g20949 (n_9570, n14280);
  and g20950 (n14283, n_9570, n14282);
  not g20951 (n_9571, n14046);
  and g20952 (n14284, n_9571, n14124);
  and g20953 (n14285, pi0120, n14284);
  not g20954 (n_9572, n14283);
  and g20955 (n14286, n_162, n_9572);
  not g20956 (n_9573, n14285);
  and g20957 (n14287, n_9573, n14286);
  not g20958 (n_9574, n14245);
  not g20959 (n_9575, n14287);
  and g20960 (n14288, n_9574, n_9575);
  not g20961 (n_9576, n14288);
  and g20962 (n14289, n2608, n_9576);
  not g20963 (n_9577, n14227);
  not g20964 (n_9578, n14289);
  and g20965 (n14290, n_9577, n_9578);
  not g20966 (n_9579, n14290);
  and g20967 (n14291, n_172, n_9579);
  not g20968 (n_9580, n14216);
  and g20969 (n14292, n_171, n_9580);
  not g20970 (n_9581, n14291);
  and g20971 (n14293, n_9581, n14292);
  not g20972 (n_9582, n14201);
  not g20973 (n_9583, n14293);
  and g20974 (n14294, n_9582, n_9583);
  not g20975 (n_9584, n14294);
  and g20976 (n14295, n7429, n_9584);
  not g20977 (n_9585, n14295);
  and g20978 (n14296, n7425, n_9585);
  and g20979 (n14297, n_9400, n_9500);
  not g20980 (n_9586, n14297);
  and g20981 (n14298, n_260, n_9586);
  and g20982 (n14299, n_4137, n14297);
  and g20983 (n14300, n_8085, n14182);
  not g20984 (n_9587, n14300);
  and g20985 (n14301, n_9528, n_9587);
  not g20986 (n_9588, n14301);
  and g20987 (n14302, n_9389, n_9588);
  not g20988 (n_9589, n14302);
  and g20989 (n14303, n_9395, n_9589);
  not g20990 (n_9590, n14303);
  and g20991 (n14304, n7506, n_9590);
  not g20992 (n_9591, n14299);
  and g20993 (n14305, n2530, n_9591);
  not g20994 (n_9592, n14304);
  and g20995 (n14306, n_9592, n14305);
  not g20996 (n_9593, n14298);
  and g20997 (n14307, pi0100, n_9593);
  not g20998 (n_9594, n14306);
  and g20999 (n14308, n_9594, n14307);
  and g21000 (n14309, pi0038, n_9586);
  and g21001 (n14310, n_9571, n14060);
  and g21002 (n14311, pi0120, n14310);
  and g21003 (n14312, n14100, n14254);
  not g21004 (n_9595, n14312);
  and g21005 (n14313, n_9389, n_9595);
  and g21006 (n14314, n_9570, n14313);
  not g21007 (n_9596, n14311);
  not g21008 (n_9597, n14314);
  and g21009 (n14315, n_9596, n_9597);
  not g21010 (n_9598, n14315);
  and g21011 (n14316, n_162, n_9598);
  not g21012 (n_9599, n7554);
  and g21013 (n14317, n_9599, n14184);
  not g21014 (n_9600, n14317);
  and g21015 (n14318, n_9587, n_9600);
  not g21016 (n_9601, n14318);
  and g21017 (n14319, n_9389, n_9601);
  not g21018 (n_9602, n14319);
  and g21019 (n14320, n_9414, n_9602);
  not g21020 (n_9603, n14320);
  and g21021 (n14321, n6198, n_9603);
  and g21022 (n14322, n_3120, n14297);
  not g21023 (n_9604, n14321);
  not g21024 (n_9605, n14322);
  and g21025 (n14323, n_9604, n_9605);
  not g21026 (n_9606, n14323);
  and g21027 (n14324, n6205, n_9606);
  and g21028 (n14325, n_3140, n_9603);
  and g21029 (n14326, n6227, n14297);
  not g21030 (n_9607, n14325);
  not g21031 (n_9608, n14326);
  and g21032 (n14327, n_9607, n_9608);
  not g21033 (n_9609, n14327);
  and g21034 (n14328, n_3119, n_9609);
  not g21035 (n_9610, n14324);
  and g21036 (n14329, n7551, n_9610);
  not g21037 (n_9611, n14328);
  and g21038 (n14330, n_9611, n14329);
  and g21039 (n14331, n_9428, n14229);
  not g21040 (n_9612, n14330);
  and g21041 (n14332, n_9612, n14331);
  and g21042 (n14333, n6242, n_9606);
  and g21043 (n14334, n_3162, n_9609);
  not g21044 (n_9613, n14333);
  and g21045 (n14335, n7570, n_9613);
  not g21046 (n_9614, n14334);
  and g21047 (n14336, n_9614, n14335);
  and g21048 (n14337, n7420, n_4176);
  not g21049 (n_9615, n14337);
  and g21050 (n14338, n14238, n_9615);
  not g21051 (n_9616, n14336);
  and g21052 (n14339, n_9616, n14338);
  not g21053 (n_9617, n14332);
  and g21054 (n14340, pi0039, n_9617);
  not g21055 (n_9618, n14339);
  and g21056 (n14341, n_9618, n14340);
  not g21057 (n_9619, n14316);
  not g21058 (n_9620, n14341);
  and g21059 (n14342, n_9619, n_9620);
  not g21060 (n_9621, n14342);
  and g21061 (n14343, n_161, n_9621);
  not g21062 (n_9622, n14309);
  and g21063 (n14344, n_164, n_9622);
  not g21064 (n_9623, n14343);
  and g21065 (n14345, n_9623, n14344);
  not g21066 (n_9624, n14308);
  not g21067 (n_9625, n14345);
  and g21068 (n14346, n_9624, n_9625);
  not g21069 (n_9626, n14346);
  and g21070 (n14347, n_172, n_9626);
  not g21071 (n_9627, n14214);
  and g21072 (n14348, n_9444, n_9627);
  and g21073 (n14349, n_9520, n_9587);
  not g21074 (n_9628, n14349);
  and g21075 (n14350, n14211, n_9628);
  not g21076 (n_9629, n14348);
  not g21077 (n_9630, n14350);
  and g21078 (n14351, n_9629, n_9630);
  and g21079 (n14352, n_9443, n14203);
  not g21080 (n_9631, n14351);
  and g21081 (n14353, n_9631, n14352);
  not g21082 (n_9632, n14347);
  not g21083 (n_9633, n14353);
  and g21084 (n14354, n_9632, n_9633);
  not g21085 (n_9634, n14354);
  and g21086 (n14355, n_171, n_9634);
  and g21087 (n14356, n7474, n_9586);
  and g21088 (n14357, n_9509, n_9587);
  not g21089 (n_9635, n14357);
  and g21090 (n14358, n_9389, n_9635);
  not g21091 (n_9636, n14358);
  and g21092 (n14359, n14113, n_9636);
  not g21093 (n_9637, n14356);
  not g21094 (n_9638, n14359);
  and g21095 (n14360, n_9637, n_9638);
  not g21096 (n_9639, n14360);
  and g21097 (n14361, n2610, n_9639);
  and g21098 (n14362, n_766, n_9586);
  not g21099 (n_9640, n14362);
  and g21100 (n14363, pi0075, n_9640);
  not g21101 (n_9641, n14361);
  and g21102 (n14364, n_9641, n14363);
  not g21103 (n_9642, n14364);
  and g21104 (n14365, n7429, n_9642);
  not g21105 (n_9643, n14355);
  and g21106 (n14366, n_9643, n14365);
  not g21107 (n_9644, n14366);
  and g21108 (n14367, n14030, n_9644);
  not g21109 (n_9645, n14296);
  not g21110 (n_9646, n14367);
  and g21111 (n14368, n_9645, n_9646);
  not g21112 (n_9647, n14179);
  and g21113 (n14369, n14176, n_9647);
  not g21114 (n_9648, n14368);
  and g21115 (n14370, n_9648, n14369);
  and g21116 (n14371, n_8134, n7623);
  not g21117 (n_9649, n14310);
  and g21118 (n14372, n_162, n_9649);
  and g21119 (n14373, n7420, n_4165);
  and g21120 (n14374, n_4167, n_9450);
  not g21121 (n_9650, n14374);
  and g21122 (n14375, n6198, n_9650);
  and g21123 (n14376, n_3120, n_8134);
  not g21124 (n_9651, n14375);
  not g21125 (n_9652, n14376);
  and g21126 (n14377, n_9651, n_9652);
  not g21127 (n_9653, n14377);
  and g21128 (n14378, n6205, n_9653);
  and g21129 (n14379, n_3140, n_9650);
  and g21130 (n14380, n6227, n_8134);
  not g21131 (n_9654, n14379);
  not g21132 (n_9655, n14380);
  and g21133 (n14381, n_9654, n_9655);
  not g21134 (n_9656, n14381);
  and g21135 (n14382, n_3119, n_9656);
  not g21136 (n_9657, n14378);
  and g21137 (n14383, n7551, n_9657);
  not g21138 (n_9658, n14382);
  and g21139 (n14384, n_9658, n14383);
  not g21140 (n_9659, n14373);
  and g21141 (n14385, n_234, n_9659);
  not g21142 (n_9660, n14384);
  and g21143 (n14386, n_9660, n14385);
  and g21144 (n14387, n6242, n_9653);
  and g21145 (n14388, n_3162, n_9656);
  not g21146 (n_9661, n14387);
  and g21147 (n14389, n7570, n_9661);
  not g21148 (n_9662, n14388);
  and g21149 (n14390, n_9662, n14389);
  and g21150 (n14391, pi0299, n_9615);
  not g21151 (n_9663, n14390);
  and g21152 (n14392, n_9663, n14391);
  not g21153 (n_9664, n14386);
  not g21154 (n_9665, n14392);
  and g21155 (n14393, n_9664, n_9665);
  not g21156 (n_9666, n14393);
  and g21157 (n14394, pi0039, n_9666);
  not g21158 (n_9667, n14394);
  and g21159 (n14395, n_161, n_9667);
  not g21160 (n_9668, n14372);
  and g21161 (n14396, n_9668, n14395);
  and g21162 (n14397, n_164, n_9436);
  not g21163 (n_9669, n14396);
  and g21164 (n14398, n_9669, n14397);
  not g21165 (n_9670, n14371);
  not g21166 (n_9671, n14398);
  and g21167 (n14399, n_9670, n_9671);
  not g21168 (n_9672, n14399);
  and g21169 (n14400, n_172, n_9672);
  not g21170 (n_9673, n14104);
  not g21171 (n_9674, n14400);
  and g21172 (n14401, n_9673, n_9674);
  not g21173 (n_9675, n14401);
  and g21174 (n14402, n_171, n_9675);
  and g21175 (n14403, n7420, n_4118);
  and g21176 (n14404, n7475, n14111);
  not g21177 (n_9676, n14403);
  and g21178 (n14405, pi0075, n_9676);
  not g21179 (n_9677, n14404);
  and g21180 (n14406, n_9677, n14405);
  not g21181 (n_9678, n14402);
  not g21182 (n_9679, n14406);
  and g21183 (n14407, n_9678, n_9679);
  not g21184 (n_9680, n14407);
  and g21185 (n14408, n14027, n_9680);
  and g21186 (n14409, n_4196, n_9492);
  not g21187 (n_9681, n14284);
  and g21188 (n14410, n_162, n_9681);
  not g21189 (n_9682, n14410);
  and g21190 (n14411, n7612, n_9682);
  not g21191 (n_9683, n14411);
  and g21192 (n14412, n_164, n_9683);
  not g21193 (n_9684, n14412);
  and g21194 (n14413, n_4211, n_9684);
  not g21195 (n_9685, n14413);
  and g21196 (n14414, n_172, n_9685);
  not g21197 (n_9686, n14414);
  and g21198 (n14415, n_4219, n_9686);
  not g21199 (n_9687, n14415);
  and g21200 (n14416, n_171, n_9687);
  not g21201 (n_9688, n14416);
  and g21202 (n14417, n_4221, n_9688);
  not g21203 (n_9689, n14028);
  and g21204 (n14418, n7425, n_9689);
  not g21205 (n_9690, n14417);
  and g21206 (n14419, n_9690, n14418);
  not g21207 (n_9691, n14408);
  not g21208 (n_9692, n14409);
  and g21209 (n14420, n_9691, n_9692);
  not g21210 (n_9693, n14419);
  and g21211 (n14421, n_9693, n14420);
  and g21212 (n14422, pi0120, n14169);
  not g21213 (n_9694, n14421);
  and g21214 (n14423, n_9694, n14422);
  not g21215 (n_9695, n14370);
  not g21216 (n_9696, n14423);
  and g21217 (n14424, n_9695, n_9696);
  not g21218 (n_9697, n14025);
  not g21219 (n_9698, n14424);
  and g21220 (n14425, n_9697, n_9698);
  or g21221 (po0278, n14178, n14425);
  not g21222 (n_9701, pi0134);
  not g21223 (n_9702, pi0135);
  and g21224 (n14427, n_9701, n_9702);
  not g21225 (n_9704, pi0136);
  and g21226 (n14428, n_9704, n14427);
  not g21227 (n_9706, pi0130);
  and g21228 (n14429, n_9706, n14428);
  not g21229 (n_9708, pi0132);
  and g21230 (n14430, n_9708, n14429);
  not g21231 (n_9710, pi0126);
  and g21232 (n14431, n_9710, n14430);
  not g21233 (n_9712, pi0121);
  and g21234 (n14432, n_9712, n14431);
  not g21235 (n_9715, pi0125);
  not g21236 (n_9716, pi0133);
  and g21237 (n14433, n_9715, n_9716);
  not g21238 (n_9717, n14433);
  and g21239 (n14434, pi0121, n_9717);
  and g21240 (n14435, n_9712, n14433);
  not g21241 (n_9718, n14434);
  not g21242 (n_9719, n14435);
  and g21243 (n14436, n_9718, n_9719);
  not g21244 (n_9720, n14432);
  not g21245 (n_9721, n14436);
  and g21246 (n14437, n_9720, n_9721);
  and g21247 (n14438, n2478, n10152);
  and g21248 (n14439, n_138, n14438);
  and g21249 (n14440, n_172, n14439);
  not g21250 (n_9722, n14437);
  and g21251 (n14441, n_9722, n14440);
  and g21252 (n14442, pi0051, pi0146);
  and g21253 (n14443, pi0051, n6197);
  and g21254 (n14444, n_268, n14443);
  not g21255 (n_9723, n14444);
  and g21256 (n14445, pi0161, n_9723);
  not g21257 (n_9724, n14439);
  and g21258 (n14446, n6197, n_9724);
  not g21259 (n_9725, n14442);
  not g21260 (n_9726, n14445);
  and g21261 (n14447, n_9725, n_9726);
  and g21262 (n14448, n14446, n14447);
  not g21263 (n_9727, n14448);
  and g21264 (n14449, n_172, n_9727);
  and g21265 (n14450, pi0087, n_9107);
  not g21266 (n_9728, n14450);
  and g21267 (n14451, pi0232, n_9728);
  not g21268 (n_9729, n14449);
  and g21269 (n14452, n_9729, n14451);
  not g21270 (n_9730, n14441);
  and g21271 (n14453, po1038, n_9730);
  not g21272 (n_9731, n14452);
  and g21273 (n14454, n_9731, n14453);
  not g21274 (n_9732, n2570);
  and g21275 (n14455, n_172, n_9732);
  and g21276 (n14456, n_9724, n14455);
  and g21277 (n14457, n_738, n14443);
  not g21278 (n_9733, n14457);
  and g21279 (n14458, pi0144, n_9733);
  and g21280 (n14459, pi0051, pi0142);
  not g21281 (n_9734, n14459);
  and g21282 (n14460, n14446, n_9734);
  not g21283 (n_9735, n14458);
  and g21284 (n14461, n_9735, n14460);
  not g21285 (n_9736, n14461);
  and g21286 (n14462, n_234, n_9736);
  and g21287 (n14463, pi0299, n_9727);
  not g21288 (n_9737, n14462);
  and g21289 (n14464, pi0232, n_9737);
  not g21290 (n_9738, n14463);
  and g21291 (n14465, n_9738, n14464);
  not g21292 (n_9739, n14465);
  and g21293 (n14466, n14456, n_9739);
  and g21294 (n14467, pi0100, n14439);
  not g21295 (n_9740, n14467);
  and g21296 (n14468, n2535, n_9740);
  and g21297 (n14469, pi0100, n14465);
  and g21298 (n14470, pi0038, n_9739);
  not g21299 (n_9741, n14470);
  and g21300 (n14471, n_164, n_9741);
  and g21301 (n14472, pi0038, n_9724);
  not g21302 (n_9742, n14472);
  and g21303 (n14473, n_164, n_9742);
  not g21304 (n_9743, n14471);
  not g21305 (n_9744, n14473);
  and g21306 (n14474, n_9743, n_9744);
  and g21307 (n14475, n_264, n_9723);
  and g21308 (n14476, n2705, n7445);
  and g21309 (n14477, n_4119, pi0314);
  and g21310 (n14478, n14476, n14477);
  and g21311 (n14479, n2467, n10151);
  and g21312 (n14480, n13047, n14479);
  and g21316 (n14484, n8897, n14478);
  and g21317 (n14485, n14483, n14484);
  and g21318 (n14486, n2519, n14485);
  and g21319 (n14487, n2770, n14480);
  and g21323 (n14491, pi0072, n6479);
  and g21324 (n14492, n14490, n14491);
  not g21325 (n_9745, n14476);
  and g21326 (n14493, n14438, n_9745);
  not g21327 (n_9746, n14493);
  and g21328 (n14494, n_138, n_9746);
  and g21329 (n14495, n_4119, n11663);
  and g21330 (n14496, n14487, n14495);
  and g21331 (n14497, pi0086, n14487);
  not g21332 (n_9747, n14483);
  not g21333 (n_9748, n14497);
  and g21334 (n14498, n_9747, n_9748);
  not g21335 (n_9749, n14498);
  and g21336 (n14499, n11076, n_9749);
  not g21337 (n_9750, n14496);
  and g21338 (n14500, n14438, n_9750);
  not g21339 (n_9751, n14499);
  and g21340 (n14501, n_9751, n14500);
  not g21341 (n_9752, n14501);
  and g21342 (n14502, n14494, n_9752);
  and g21343 (n14503, n2519, n14502);
  not g21344 (n_9753, n14503);
  and g21345 (n14504, n14439, n_9753);
  not g21346 (n_9754, n14492);
  and g21347 (n14505, n_9754, n14504);
  not g21348 (n_9755, n14486);
  and g21349 (n14506, n_9755, n14505);
  not g21350 (n_9756, n14506);
  and g21351 (n14507, n_3102, n_9756);
  and g21352 (n14508, pi0072, n10342);
  not g21353 (n_9757, n14443);
  not g21354 (n_9758, n14508);
  and g21355 (n14509, n_9757, n_9758);
  not g21356 (n_9759, n14509);
  and g21357 (n14510, n6197, n_9759);
  not g21358 (n_9760, n14507);
  not g21359 (n_9761, n14510);
  and g21360 (n14511, n_9760, n_9761);
  not g21361 (n_9762, n14511);
  and g21362 (n14512, n14475, n_9762);
  and g21363 (n14513, n14439, n_9755);
  and g21364 (n14514, n_9753, n14513);
  not g21365 (n_9763, n14514);
  and g21366 (n14515, n_3102, n_9763);
  not g21367 (n_9764, n14446);
  not g21368 (n_9765, n14515);
  and g21369 (n14516, n_9764, n_9765);
  and g21370 (n14517, n_9754, n14516);
  and g21371 (n14518, pi0146, n14517);
  and g21372 (n14519, n_138, n6197);
  and g21373 (n14520, n14438, n_9754);
  not g21374 (n_9766, n14520);
  and g21375 (n14521, n14519, n_9766);
  not g21376 (n_9767, n14521);
  and g21377 (n14522, n_268, n_9767);
  and g21378 (n14523, n_9760, n14522);
  not g21379 (n_9768, n14518);
  and g21380 (n14524, pi0161, n_9768);
  not g21381 (n_9769, n14523);
  and g21382 (n14525, n_9769, n14524);
  not g21383 (n_9770, n14512);
  not g21384 (n_9771, n14525);
  and g21385 (n14526, n_9770, n_9771);
  not g21386 (n_9772, n14526);
  and g21387 (n14527, n9572, n_9772);
  and g21388 (n14528, n_3102, n14506);
  and g21389 (n14529, n_138, n14478);
  and g21390 (n14530, n13439, n14529);
  not g21391 (n_9773, n14530);
  and g21392 (n14531, n_134, n_9773);
  not g21393 (n_9774, n14531);
  and g21394 (n14532, n6480, n_9774);
  not g21395 (n_9775, n14532);
  and g21396 (n14533, n6197, n_9775);
  not g21397 (n_9776, n14528);
  not g21398 (n_9777, n14533);
  and g21399 (n14534, n_9776, n_9777);
  not g21400 (n_9778, n14534);
  and g21401 (n14535, n_268, n_9778);
  and g21402 (n14536, n2519, n6197);
  and g21403 (n14537, n14530, n14536);
  not g21404 (n_9779, n14537);
  and g21405 (n14538, n14511, n_9779);
  and g21406 (n14539, pi0146, n14538);
  not g21407 (n_9780, n14535);
  and g21408 (n14540, n_264, n_9780);
  not g21409 (n_9781, n14539);
  and g21410 (n14541, n_9781, n14540);
  and g21411 (n14542, n14519, n14520);
  and g21412 (n14543, n_9755, n14542);
  not g21413 (n_9782, n14543);
  and g21414 (n14544, n_9757, n_9782);
  and g21415 (n14545, pi0146, n_9724);
  not g21416 (n_9783, n14544);
  not g21417 (n_9784, n14545);
  and g21418 (n14546, n_9783, n_9784);
  not g21419 (n_9785, n14546);
  and g21420 (n14547, pi0161, n_9785);
  and g21421 (n14548, n_9776, n14547);
  not g21422 (n_9786, n14541);
  not g21423 (n_9787, n14548);
  and g21424 (n14549, n_9786, n_9787);
  not g21425 (n_9788, n14549);
  and g21426 (n14550, n9603, n_9788);
  not g21427 (n_9789, n14527);
  not g21428 (n_9790, n14550);
  and g21429 (n14551, n_9789, n_9790);
  not g21430 (n_9791, n14551);
  and g21431 (n14552, pi0156, n_9791);
  not g21432 (n_9792, n14517);
  and g21433 (n14553, pi0144, n_9792);
  and g21434 (n14554, n_298, n_9762);
  not g21435 (n_9793, n14553);
  not g21436 (n_9794, n14554);
  and g21437 (n14555, n_9793, n_9794);
  not g21438 (n_9795, n14555);
  and g21439 (n14556, n_9733, n_9795);
  not g21440 (n_9796, n14556);
  and g21441 (n14557, pi0180, n_9796);
  and g21442 (n14558, n_738, n_9778);
  and g21443 (n14559, pi0142, n14538);
  not g21444 (n_9797, n14558);
  and g21445 (n14560, n_298, n_9797);
  not g21446 (n_9798, n14559);
  and g21447 (n14561, n_9798, n14560);
  and g21448 (n14562, n_9755, n14517);
  not g21449 (n_9799, n14562);
  and g21450 (n14563, n14458, n_9799);
  not g21451 (n_9800, n14563);
  and g21452 (n14564, n_6015, n_9800);
  not g21453 (n_9801, n14561);
  and g21454 (n14565, n_9801, n14564);
  not g21455 (n_9802, n14557);
  and g21456 (n14566, pi0179, n_9802);
  not g21457 (n_9803, n14565);
  and g21458 (n14567, n_9803, n14566);
  and g21459 (n14568, n14458, n_9756);
  and g21460 (n14569, n_4119, n_7584);
  and g21461 (n14570, pi0024, n_7587);
  not g21462 (n_9804, n14569);
  not g21463 (n_9805, n14570);
  and g21464 (n14571, n_9804, n_9805);
  not g21465 (n_9806, n14571);
  and g21466 (n14572, n_3310, n_9806);
  and g21467 (n14573, pi0314, n_7587);
  not g21468 (n_9807, n14572);
  not g21469 (n_9808, n14573);
  and g21470 (n14574, n_9807, n_9808);
  and g21471 (n14575, n7445, n8960);
  and g21472 (n14576, n14574, n14575);
  not g21473 (n_9809, n14576);
  and g21474 (n14577, n_138, n_9809);
  and g21475 (n14578, n_9758, n14577);
  not g21476 (n_9810, n14578);
  and g21477 (n14579, n6197, n_9810);
  not g21478 (n_9811, n14579);
  and g21479 (n14580, n_9760, n_9811);
  and g21480 (n14581, pi0142, n14580);
  and g21481 (n14582, n2708, n14574);
  not g21482 (n_9812, n14582);
  and g21483 (n14583, n_134, n_9812);
  not g21484 (n_9813, n14583);
  and g21485 (n14584, n6480, n_9813);
  not g21486 (n_9814, n14584);
  and g21487 (n14585, n6197, n_9814);
  not g21488 (n_9815, n14585);
  and g21489 (n14586, n_9776, n_9815);
  not g21490 (n_9816, n14586);
  and g21491 (n14587, n_738, n_9816);
  not g21492 (n_9817, n14581);
  and g21493 (n14588, n_298, n_9817);
  not g21494 (n_9818, n14587);
  and g21495 (n14589, n_9818, n14588);
  not g21496 (n_9819, n14568);
  and g21497 (n14590, n_6015, n_9819);
  not g21498 (n_9820, n14589);
  and g21499 (n14591, n_9820, n14590);
  not g21500 (n_9821, n14505);
  and g21501 (n14592, n_9821, n14519);
  not g21502 (n_9822, n14592);
  and g21503 (n14593, n_9760, n_9822);
  not g21504 (n_9823, n14504);
  and g21505 (n14594, n6197, n_9823);
  not g21506 (n_9824, n14594);
  and g21507 (n14595, n_738, n_9824);
  not g21508 (n_9825, n14438);
  and g21509 (n14596, n_138, n_9825);
  and g21510 (n14597, n6197, n14596);
  not g21511 (n_9826, n14536);
  not g21512 (n_9827, n14597);
  and g21513 (n14598, n_9826, n_9827);
  not g21514 (n_9828, n14502);
  and g21515 (n14599, n2519, n_9828);
  not g21516 (n_9829, n14598);
  not g21517 (n_9830, n14599);
  and g21518 (n14600, n_9829, n_9830);
  not g21519 (n_9831, n14600);
  and g21520 (n14601, pi0142, n_9831);
  not g21521 (n_9832, n14595);
  not g21522 (n_9833, n14601);
  and g21523 (n14602, n_9832, n_9833);
  not g21524 (n_9834, n14516);
  not g21525 (n_9835, n14602);
  and g21526 (n14603, n_9834, n_9835);
  not g21527 (n_9836, n14603);
  and g21528 (n14604, n14593, n_9836);
  not g21529 (n_9837, n14604);
  and g21530 (n14605, pi0144, n_9837);
  and g21531 (n14606, n2708, n14571);
  not g21532 (n_9838, n14606);
  and g21533 (n14607, n_134, n_9838);
  not g21534 (n_9839, n14607);
  and g21535 (n14608, n6480, n_9839);
  not g21536 (n_9840, n14608);
  and g21537 (n14609, n6197, n_9840);
  not g21538 (n_9841, n14609);
  and g21539 (n14610, n_9776, n_9841);
  not g21540 (n_9842, n14610);
  and g21541 (n14611, n_738, n_9842);
  and g21542 (n14612, n14536, n14606);
  not g21543 (n_9843, n14612);
  and g21544 (n14613, n_9761, n_9843);
  and g21545 (n14614, n_9760, n14613);
  and g21546 (n14615, pi0142, n14614);
  not g21547 (n_9844, n14615);
  and g21548 (n14616, n_298, n_9844);
  not g21549 (n_9845, n14611);
  and g21550 (n14617, n_9845, n14616);
  not g21551 (n_9846, n14605);
  and g21552 (n14618, pi0180, n_9846);
  not g21553 (n_9847, n14617);
  and g21554 (n14619, n_9847, n14618);
  not g21555 (n_9848, n14619);
  and g21556 (n14620, n_7636, n_9848);
  not g21557 (n_9849, n14591);
  and g21558 (n14621, n_9849, n14620);
  not g21559 (n_9850, n14567);
  not g21560 (n_9851, n14621);
  and g21561 (n14622, n_9850, n_9851);
  not g21562 (n_9852, n14622);
  and g21563 (n14623, n_234, n_9852);
  and g21564 (n14624, pi0146, n14614);
  and g21565 (n14625, n_268, n_9842);
  not g21566 (n_9853, n14624);
  and g21567 (n14626, n9572, n_9853);
  not g21568 (n_9854, n14625);
  and g21569 (n14627, n_9854, n14626);
  and g21570 (n14628, n_268, n_9816);
  and g21571 (n14629, pi0146, n14580);
  not g21572 (n_9855, n14628);
  and g21573 (n14630, n9603, n_9855);
  not g21574 (n_9856, n14629);
  and g21575 (n14631, n_9856, n14630);
  not g21576 (n_9857, n14627);
  and g21577 (n14632, n_264, n_9857);
  not g21578 (n_9858, n14631);
  and g21579 (n14633, n_9858, n14632);
  and g21580 (n14634, n_268, n_9824);
  and g21581 (n14635, pi0146, n_9831);
  not g21582 (n_9859, n14634);
  not g21583 (n_9860, n14635);
  and g21584 (n14636, n_9859, n_9860);
  not g21585 (n_9861, n14636);
  and g21586 (n14637, n_9834, n_9861);
  not g21587 (n_9862, n14637);
  and g21588 (n14638, n14593, n_9862);
  not g21589 (n_9863, n14638);
  and g21590 (n14639, n9572, n_9863);
  and g21591 (n14640, n9603, n_9723);
  and g21592 (n14641, n_9756, n14640);
  not g21593 (n_9864, n14641);
  and g21594 (n14642, pi0161, n_9864);
  not g21595 (n_9865, n14639);
  and g21596 (n14643, n_9865, n14642);
  not g21597 (n_9866, n14643);
  and g21598 (n14644, n_7638, n_9866);
  not g21599 (n_9867, n14633);
  and g21600 (n14645, n_9867, n14644);
  not g21601 (n_9868, n14552);
  not g21602 (n_9869, n14645);
  and g21603 (n14646, n_9868, n_9869);
  not g21604 (n_9870, n14623);
  and g21605 (n14647, n_9870, n14646);
  not g21606 (n_9871, n14647);
  and g21607 (n14648, n9159, n_9871);
  and g21608 (n14649, n2519, n14490);
  not g21609 (n_9872, n7607);
  and g21610 (n14650, n_3489, n_9872);
  not g21611 (n_9873, n14650);
  and g21612 (n14651, n14649, n_9873);
  and g21613 (n14652, n_3410, n14439);
  not g21614 (n_9874, n14651);
  and g21615 (n14653, n_9874, n14652);
  not g21616 (n_9875, n14649);
  and g21617 (n14654, n14439, n_9875);
  not g21618 (n_9876, n14654);
  and g21619 (n14655, n_138, n_9876);
  not g21620 (n_9877, n14655);
  and g21621 (n14656, n_3084, n_9877);
  and g21622 (n14657, n_3084, n6197);
  not g21623 (n_9878, n14657);
  and g21624 (n14658, n_9827, n_9878);
  not g21625 (n_9879, n14656);
  not g21626 (n_9880, n14658);
  and g21627 (n14659, n_9879, n_9880);
  not g21628 (n_9881, n14460);
  not g21629 (n_9882, n14659);
  and g21630 (n14660, n_9881, n_9882);
  not g21631 (n_9883, n14660);
  and g21632 (n14661, n9051, n_9883);
  and g21633 (n14662, n14438, n14661);
  and g21634 (n14663, n_9724, n_9733);
  not g21635 (n_9884, n6405);
  not g21636 (n_9885, n14663);
  and g21637 (n14664, n_9884, n_9885);
  not g21638 (n_9886, n14664);
  and g21639 (n14665, pi0144, n_9886);
  and g21640 (n14666, pi0051, n_3102);
  not g21641 (n_9887, n14666);
  and g21642 (n14667, n_9877, n_9887);
  and g21643 (n14668, n6405, n_9734);
  and g21644 (n14669, n14667, n14668);
  not g21645 (n_9888, n14669);
  and g21646 (n14670, n14665, n_9888);
  not g21647 (n_9889, n14662);
  and g21648 (n14671, n_9889, n14670);
  and g21649 (n14672, n_3102, n_9876);
  not g21650 (n_9890, n14672);
  and g21651 (n14673, n_3550, n_9890);
  not g21652 (n_9891, n14673);
  and g21653 (n14674, n_738, n_9891);
  and g21654 (n14675, n2515, n7450);
  not g21655 (n_9892, n14675);
  and g21656 (n14676, n_138, n_9892);
  not g21657 (n_9893, n14676);
  and g21658 (n14677, n6197, n_9893);
  not g21659 (n_9894, n14677);
  and g21660 (n14678, n_9890, n_9894);
  not g21661 (n_9895, n14678);
  and g21662 (n14679, pi0142, n_9895);
  not g21663 (n_9896, n14674);
  and g21664 (n14680, n6405, n_9896);
  not g21665 (n_9897, n14679);
  and g21666 (n14681, n_9897, n14680);
  not g21667 (n_9898, n14681);
  and g21668 (n14682, n_5891, n_9898);
  and g21669 (n14683, n_138, n14657);
  not g21670 (n_9899, n14683);
  and g21671 (n14684, n_9895, n_9899);
  and g21672 (n14685, pi0224, n_9733);
  and g21673 (n14686, n14684, n14685);
  not g21674 (n_9900, n14682);
  not g21675 (n_9901, n14686);
  and g21676 (n14687, n_9900, n_9901);
  and g21677 (n14688, n_9884, n14597);
  not g21678 (n_9902, n14688);
  and g21679 (n14689, n_9886, n_9902);
  not g21680 (n_9903, n14665);
  and g21681 (n14690, n_9903, n14689);
  not g21682 (n_9904, n14687);
  and g21683 (n14691, n_9904, n14690);
  not g21684 (n_9905, n14671);
  and g21685 (n14692, pi0181, n_9905);
  not g21686 (n_9906, n14691);
  and g21687 (n14693, n_9906, n14692);
  and g21688 (n14694, n_9898, n14690);
  not g21689 (n_9907, n14670);
  and g21690 (n14695, n_6429, n_9907);
  not g21691 (n_9908, n14694);
  and g21692 (n14696, n_9908, n14695);
  not g21693 (n_9909, n14696);
  and g21694 (n14697, n_234, n_9909);
  not g21695 (n_9910, n14693);
  and g21696 (n14698, n_9910, n14697);
  and g21697 (n14699, n_9723, n_9876);
  not g21698 (n_9911, n14699);
  and g21699 (n14700, pi0161, n_9911);
  and g21700 (n14701, n_268, n_9891);
  and g21701 (n14702, pi0146, n_9895);
  not g21702 (n_9912, n14701);
  and g21703 (n14703, n_264, n_9912);
  not g21704 (n_9913, n14702);
  and g21705 (n14704, n_9913, n14703);
  not g21706 (n_9914, n14700);
  not g21707 (n_9915, n14704);
  and g21708 (n14705, n_9914, n_9915);
  not g21709 (n_9916, n14705);
  and g21710 (n14706, n6379, n_9916);
  and g21711 (n14707, n_9724, n_9727);
  not g21712 (n_9917, n6379);
  not g21713 (n_9918, n14707);
  and g21714 (n14708, n_9917, n_9918);
  not g21715 (n_9919, n14708);
  and g21716 (n14709, n9793, n_9919);
  not g21717 (n_9920, n14706);
  and g21718 (n14710, n_9920, n14709);
  and g21719 (n14711, n_5881, n_9920);
  and g21720 (n14712, n14475, n14684);
  and g21721 (n14713, n14649, n_9878);
  not g21722 (n_9921, n14713);
  and g21723 (n14714, n14439, n_9921);
  not g21724 (n_9922, n14714);
  and g21725 (n14715, n14445, n_9922);
  not g21726 (n_9923, n14712);
  not g21727 (n_9924, n14715);
  and g21728 (n14716, n_9923, n_9924);
  not g21729 (n_9925, n14716);
  and g21730 (n14717, pi0216, n_9925);
  not g21731 (n_9926, n14711);
  not g21732 (n_9927, n14717);
  and g21733 (n14718, n_9926, n_9927);
  and g21734 (n14719, n9794, n_9919);
  not g21735 (n_9928, n14718);
  and g21736 (n14720, n_9928, n14719);
  not g21743 (n_9932, n14653);
  and g21744 (n14724, pi0039, n_9932);
  not g21745 (n_9933, n14723);
  and g21746 (n14725, n_9933, n14724);
  and g21747 (n14726, n_162, n_3410);
  and g21748 (n14727, n_9756, n14726);
  not g21749 (n_9934, n14725);
  not g21750 (n_9935, n14727);
  and g21751 (n14728, n_9934, n_9935);
  not g21752 (n_9936, n14648);
  and g21753 (n14729, n_9936, n14728);
  not g21754 (n_9937, n14729);
  and g21755 (n14730, n_161, n_9937);
  not g21756 (n_9938, n14474);
  not g21757 (n_9939, n14730);
  and g21758 (n14731, n_9938, n_9939);
  not g21759 (n_9940, n14469);
  and g21760 (n14732, n14468, n_9940);
  not g21761 (n_9941, n14731);
  and g21762 (n14733, n_9941, n14732);
  and g21763 (n14734, n_7617, n_234);
  and g21764 (n14735, n_7591, pi0299);
  not g21765 (n_9942, n14734);
  not g21766 (n_9943, n14735);
  and g21767 (n14736, n_9942, n_9943);
  and g21768 (n14737, n7473, n14736);
  not g21769 (n_9944, n14737);
  and g21770 (n14738, pi0087, n_9944);
  not g21771 (n_9945, n14738);
  and g21777 (n14742, n14455, n_9739);
  and g21778 (n14743, n_6143, n14463);
  and g21779 (n14744, n14445, n_9779);
  not g21780 (n_9948, n14513);
  and g21781 (n14745, n6197, n_9948);
  and g21782 (n14746, n_268, n14745);
  not g21783 (n_9949, n14485);
  and g21784 (n14747, n14438, n_9949);
  not g21785 (n_9950, n14747);
  and g21786 (n14748, n_138, n_9950);
  not g21787 (n_9951, n14748);
  and g21788 (n14749, n2519, n_9951);
  not g21789 (n_9952, n14749);
  and g21790 (n14750, n_9829, n_9952);
  and g21791 (n14751, pi0146, n14750);
  not g21792 (n_9953, n14746);
  and g21793 (n14752, n_264, n_9953);
  not g21794 (n_9954, n14751);
  and g21795 (n14753, n_9954, n14752);
  not g21796 (n_9955, n14744);
  not g21797 (n_9956, n14753);
  and g21798 (n14754, n_9955, n_9956);
  not g21799 (n_9957, n14754);
  and g21800 (n14755, n9572, n_9957);
  not g21801 (n_9958, n14743);
  and g21802 (n14756, pi0232, n_9958);
  not g21803 (n_9959, n14755);
  and g21804 (n14757, n_9959, n14756);
  and g21805 (n14758, n_7638, n2530);
  not g21806 (n_9960, n14757);
  and g21807 (n14759, n_9960, n14758);
  and g21808 (n14760, n_6307, n14463);
  and g21809 (n14761, n_6429, n14461);
  and g21810 (n14762, n_298, n_9881);
  not g21811 (n_9961, n14661);
  and g21812 (n14763, n_9961, n14762);
  and g21813 (n14764, n9051, n14657);
  and g21814 (n14765, pi0142, n_207);
  and g21815 (n14766, n_738, n_9892);
  not g21816 (n_9962, n14765);
  and g21817 (n14767, n14764, n_9962);
  not g21818 (n_9963, n14766);
  and g21819 (n14768, n_9963, n14767);
  not g21820 (n_9964, n14768);
  and g21821 (n14769, n14458, n_9964);
  not g21822 (n_9965, n14763);
  and g21823 (n14770, pi0181, n_9965);
  not g21824 (n_9966, n14769);
  and g21825 (n14771, n_9966, n14770);
  not g21826 (n_9967, n14761);
  and g21827 (n14772, n_234, n_9967);
  not g21828 (n_9968, n14771);
  and g21829 (n14773, n_9968, n14772);
  and g21830 (n14774, n_5881, n14448);
  and g21831 (n14775, n14475, n_9882);
  and g21832 (n14776, n6197, n6380);
  not g21833 (n_9969, n14776);
  and g21834 (n14777, n14445, n_9969);
  not g21835 (n_9970, n14775);
  and g21836 (n14778, n9036, n_9970);
  not g21837 (n_9971, n14777);
  and g21838 (n14779, n_9971, n14778);
  not g21839 (n_9972, n14774);
  and g21840 (n14780, n9794, n_9972);
  not g21841 (n_9973, n14779);
  and g21842 (n14781, n_9973, n14780);
  not g21849 (n_9977, n14577);
  and g21850 (n14785, n6197, n_9977);
  and g21851 (n14786, n_9725, n14785);
  not g21852 (n_9978, n14786);
  and g21853 (n14787, pi0161, n_9978);
  and g21854 (n14788, n6197, n_9763);
  and g21855 (n14789, n_268, n14788);
  and g21856 (n14790, n14476, n14747);
  and g21857 (n14791, n14501, n14790);
  not g21858 (n_9979, n14791);
  and g21859 (n14792, n14494, n_9979);
  not g21860 (n_9980, n14792);
  and g21861 (n14793, n2519, n_9980);
  not g21862 (n_9981, n14793);
  and g21863 (n14794, n_9829, n_9981);
  and g21864 (n14795, pi0146, n14794);
  not g21865 (n_9982, n14789);
  and g21866 (n14796, n_264, n_9982);
  not g21867 (n_9983, n14795);
  and g21868 (n14797, n_9983, n14796);
  not g21869 (n_9984, n14787);
  not g21870 (n_9985, n14797);
  and g21871 (n14798, n_9984, n_9985);
  not g21872 (n_9986, n14798);
  and g21873 (n14799, n9572, n_9986);
  and g21874 (n14800, n14445, n_9843);
  and g21875 (n14801, n_264, n_9861);
  not g21876 (n_9987, n14800);
  not g21877 (n_9988, n14801);
  and g21878 (n14802, n_9987, n_9988);
  not g21879 (n_9989, n14802);
  and g21880 (n14803, n9603, n_9989);
  not g21881 (n_9990, n14803);
  and g21882 (n14804, pi0232, n_9990);
  not g21883 (n_9991, n14799);
  and g21884 (n14805, n_9991, n14804);
  not g21885 (n_9992, n14805);
  and g21886 (n14806, pi0156, n_9992);
  and g21887 (n14807, n_738, n14788);
  and g21888 (n14808, pi0142, n14794);
  not g21889 (n_9993, n14807);
  and g21890 (n14809, n_298, n_9993);
  not g21891 (n_9994, n14808);
  and g21892 (n14810, n_9994, n14809);
  and g21893 (n14811, n_9734, n14785);
  not g21894 (n_9995, n14811);
  and g21895 (n14812, pi0144, n_9995);
  not g21896 (n_9996, n14810);
  and g21897 (n14813, pi0180, n_9996);
  not g21898 (n_9997, n14812);
  and g21899 (n14814, n_9997, n14813);
  and g21900 (n14815, n14458, n_9843);
  and g21901 (n14816, n_298, n_9835);
  not g21902 (n_9998, n14816);
  and g21903 (n14817, n_6015, n_9998);
  not g21904 (n_9999, n14815);
  and g21905 (n14818, n_9999, n14817);
  not g21906 (n_10000, n14818);
  and g21907 (n14819, pi0179, n_10000);
  not g21908 (n_10001, n14814);
  and g21909 (n14820, n_10001, n14819);
  and g21910 (n14821, n_6015, n14461);
  and g21911 (n14822, n_738, n14745);
  and g21912 (n14823, pi0142, n14750);
  not g21913 (n_10002, n14822);
  and g21914 (n14824, n_298, n_10002);
  not g21915 (n_10003, n14823);
  and g21916 (n14825, n_10003, n14824);
  and g21917 (n14826, n14458, n_9779);
  not g21918 (n_10004, n14825);
  and g21919 (n14827, pi0180, n_10004);
  not g21920 (n_10005, n14826);
  and g21921 (n14828, n_10005, n14827);
  not g21922 (n_10006, n14821);
  and g21923 (n14829, n_7636, n_10006);
  not g21924 (n_10007, n14828);
  and g21925 (n14830, n_10007, n14829);
  not g21926 (n_10008, n14820);
  not g21927 (n_10009, n14830);
  and g21928 (n14831, n_10008, n_10009);
  not g21929 (n_10010, n14831);
  and g21930 (n14832, n_234, n_10010);
  not g21931 (n_10011, n14806);
  and g21932 (n14833, n_162, n_10011);
  not g21933 (n_10012, n14832);
  and g21934 (n14834, n_10012, n14833);
  not g21935 (n_10013, n14784);
  and g21936 (n14835, n_161, n_10013);
  not g21937 (n_10014, n14834);
  and g21938 (n14836, n_10014, n14835);
  not g21939 (n_10015, n14759);
  and g21940 (n14837, n14471, n_10015);
  not g21941 (n_10016, n14836);
  and g21942 (n14838, n_10016, n14837);
  and g21943 (n14839, n2535, n_9940);
  not g21944 (n_10017, n14838);
  and g21945 (n14840, n_10017, n14839);
  not g21951 (n_10020, n14843);
  and g21952 (n14844, n_4226, n_10020);
  not g21953 (n_10021, n14741);
  and g21954 (n14845, n_10021, n14844);
  or g21955 (po0279, n14454, n14845);
  and g21956 (n14847, n7420, n7427);
  and g21957 (n14848, n7429, n14407);
  not g21958 (n_10022, n14848);
  and g21959 (n14849, n14027, n_10022);
  and g21960 (n14850, n7429, n14417);
  not g21961 (n_10023, n14850);
  and g21962 (n14851, n7425, n_10023);
  not g21963 (n_10024, n14849);
  and g21964 (n14852, n_4226, n_10024);
  not g21965 (n_10025, n14851);
  and g21966 (n14853, n_10025, n14852);
  or g21967 (po0280, n14847, n14853);
  not g21972 (n_10027, n14857);
  and g21973 (n14858, n_162, n_10027);
  and g21974 (n14859, n_113, n9293);
  and g21975 (n14860, n_3164, n6379);
  and g21976 (n14861, n14859, n14860);
  not g21977 (n_10028, n14861);
  and g21978 (n14862, pi0039, n_10028);
  not g21979 (n_10029, n14858);
  and g21980 (n14863, po1038, n_10029);
  not g21981 (n_10030, n14862);
  and g21982 (n14864, n_10030, n14863);
  and g21983 (n14865, pi0110, n13448);
  not g21984 (n_10031, n14865);
  and g21985 (n14866, n_162, n_10031);
  and g21986 (n14867, n_3122, n7607);
  and g21987 (n14868, n14859, n14867);
  and g21988 (n14869, pi0299, n14861);
  not g21989 (n_10032, n14868);
  and g21990 (n14870, pi0039, n_10032);
  not g21991 (n_10033, n14869);
  and g21992 (n14871, n_10033, n14870);
  not g21993 (n_10034, n14866);
  not g21994 (n_10035, n14871);
  and g21995 (n14872, n_10034, n_10035);
  and g21996 (n14873, n_161, n2571);
  not g21997 (n_10036, n14872);
  not g21998 (n_10037, n14873);
  and g21999 (n14874, n_10036, n_10037);
  not g22000 (n_10038, n10387);
  and g22001 (n14875, pi0090, n_10038);
  not g22002 (n_10039, n6429);
  and g22003 (n14876, n_95, n_10039);
  and g22004 (n14877, n_97, n2809);
  not g22005 (n_10040, n14876);
  and g22006 (n14878, n_10040, n14877);
  not g22007 (n_10041, n14878);
  and g22008 (n14879, n2468, n_10041);
  and g22009 (n14880, n_376, n_415);
  not g22010 (n_10042, n14879);
  and g22011 (n14881, n_10042, n14880);
  not g22012 (n_10043, n14881);
  and g22013 (n14882, n_60, n_10043);
  not g22014 (n_10044, n14882);
  and g22015 (n14883, n2795, n_10044);
  not g22016 (n_10045, n14883);
  and g22017 (n14884, n_57, n_10045);
  not g22018 (n_10046, n14884);
  and g22019 (n14885, n6438, n_10046);
  not g22020 (n_10047, n14885);
  and g22021 (n14886, n_105, n_10047);
  not g22022 (n_10048, n14886);
  and g22023 (n14887, n11443, n_10048);
  not g22024 (n_10049, n14887);
  and g22025 (n14888, n_43, n_10049);
  not g22026 (n_10050, n14888);
  and g22027 (n14889, n2707, n_10050);
  not g22028 (n_10051, n14875);
  and g22029 (n14890, n9073, n_10051);
  and g22030 (n14891, n14889, n14890);
  and g22031 (n14892, pi0072, n2708);
  and g22032 (n14893, n10387, n14892);
  not g22033 (n_10052, n14891);
  not g22034 (n_10053, n14893);
  and g22035 (n14894, n_10052, n_10053);
  not g22036 (n_10054, n14894);
  and g22037 (n14895, n6479, n_10054);
  not g22038 (n_10055, n14895);
  and g22039 (n14896, n_113, n_10055);
  not g22040 (n_10056, n14896);
  and g22041 (n14897, n13448, n_10056);
  and g22042 (n14898, n2897, n14889);
  not g22043 (n_10057, n14898);
  and g22044 (n14899, n_134, n_10057);
  not g22045 (n_10058, n13448);
  and g22046 (n14900, n6480, n_10058);
  not g22047 (n_10059, n14899);
  and g22048 (n14901, n_10059, n14900);
  not g22049 (n_10060, n14901);
  and g22050 (n14902, n_162, n_10060);
  not g22051 (n_10061, n14897);
  and g22052 (n14903, n_10061, n14902);
  not g22053 (n_10062, n14903);
  and g22054 (n14904, n_10035, n_10062);
  not g22055 (n_10063, n14904);
  and g22056 (n14905, n14873, n_10063);
  not g22057 (n_10064, n14874);
  and g22058 (n14906, n_4226, n_10064);
  not g22059 (n_10065, n14905);
  and g22060 (n14907, n_10065, n14906);
  not g22061 (n_10066, n14864);
  not g22062 (n_10067, n14907);
  and g22063 (po0281, n_10066, n_10067);
  and g22064 (n14909, n_9715, n14432);
  and g22065 (n14910, pi0125, pi0133);
  not g22066 (n_10068, n14910);
  and g22067 (n14911, n_9717, n_10068);
  not g22068 (n_10069, n14909);
  not g22069 (n_10070, n14911);
  and g22070 (n14912, n_10069, n_10070);
  not g22071 (n_10071, n14912);
  and g22072 (n14913, n14439, n_10071);
  and g22073 (n14914, pi0172, n14443);
  and g22074 (n14915, n_263, n14597);
  not g22075 (n_10072, n14914);
  not g22076 (n_10073, n14915);
  and g22077 (n14916, n_10072, n_10073);
  not g22078 (n_10074, n14916);
  and g22079 (n14917, pi0232, n_10074);
  not g22080 (n_10075, n14913);
  not g22081 (n_10076, n14917);
  and g22082 (n14918, n_10075, n_10076);
  not g22083 (n_10077, n14918);
  and g22084 (n14919, n_172, n_10077);
  and g22085 (n14920, pi0087, n7473);
  and g22086 (n14921, pi0162, n14920);
  not g22087 (n_10078, n14921);
  and g22088 (n14922, po1038, n_10078);
  not g22089 (n_10079, n14919);
  and g22090 (n14923, n_10079, n14922);
  and g22091 (n14924, pi0193, n14443);
  and g22092 (n14925, n_299, n14597);
  not g22093 (n_10080, n14924);
  and g22094 (n14926, n_234, n_10080);
  not g22095 (n_10081, n14925);
  and g22096 (n14927, n_10081, n14926);
  and g22097 (n14928, pi0299, n14916);
  not g22098 (n_10082, n14927);
  and g22099 (n14929, pi0232, n_10082);
  not g22100 (n_10083, n14928);
  and g22101 (n14930, n_10083, n14929);
  not g22102 (n_10084, n14930);
  and g22103 (n14931, n14455, n_10084);
  and g22104 (n14932, pi0140, n_234);
  and g22105 (n14933, pi0162, pi0299);
  not g22106 (n_10085, n14932);
  not g22107 (n_10086, n14933);
  and g22108 (n14934, n_10085, n_10086);
  not g22109 (n_10087, n14934);
  and g22110 (n14935, n7473, n_10087);
  not g22111 (n_10088, n14935);
  and g22112 (n14936, pi0087, n_10088);
  and g22113 (n14937, pi0100, n14930);
  and g22114 (n14938, n_3410, n_9758);
  not g22115 (n_10089, n14938);
  and g22116 (n14939, n_162, n_10089);
  and g22117 (n14940, n_234, n_4165);
  and g22118 (n14941, pi0299, n_4176);
  not g22119 (n_10090, n14940);
  not g22120 (n_10091, n14941);
  and g22121 (n14942, n_10090, n_10091);
  and g22122 (n14943, n2521, n14942);
  not g22123 (n_10092, n14943);
  and g22124 (n14944, n_3410, n_10092);
  not g22125 (n_10093, n14944);
  and g22126 (n14945, pi0039, n_10093);
  and g22127 (n14946, n_4176, n14916);
  and g22128 (n14947, n2521, n_3102);
  and g22129 (n14948, n6197, n_9876);
  not g22130 (n_10094, n14947);
  not g22131 (n_10095, n14948);
  and g22132 (n14949, n_10094, n_10095);
  not g22133 (n_10096, n14949);
  and g22134 (n14950, n_263, n_10096);
  and g22135 (n14951, n_9894, n_10094);
  not g22136 (n_10097, n14951);
  and g22137 (n14952, pi0152, n_10097);
  not g22138 (n_10098, n14950);
  not g22139 (n_10099, n14952);
  and g22140 (n14953, n_10098, n_10099);
  and g22141 (n14954, pi0051, n_1362);
  not g22142 (n_10100, n14953);
  not g22143 (n_10101, n14954);
  and g22144 (n14955, n_10100, n_10101);
  not g22145 (n_10102, n14955);
  and g22146 (n14956, n_20, n_10102);
  and g22147 (n14957, n6379, n14956);
  not g22148 (n_10103, n14946);
  not g22149 (n_10104, n14957);
  and g22150 (n14958, n_10103, n_10104);
  not g22151 (n_10105, n14958);
  and g22152 (n14959, n9603, n_10105);
  and g22153 (n14960, n_9917, n_10074);
  and g22154 (n14961, n14649, n14657);
  not g22155 (n_10106, n14961);
  and g22156 (n14962, n_9764, n_10106);
  and g22157 (n14963, n_263, n14962);
  and g22158 (n14964, n14657, n14675);
  not g22159 (n_10107, n14964);
  and g22160 (n14965, n_9757, n_10107);
  and g22161 (n14966, pi0152, n14965);
  not g22162 (n_10108, n14963);
  and g22163 (n14967, pi0172, n_10108);
  not g22164 (n_10109, n14966);
  and g22165 (n14968, n_10109, n14967);
  and g22166 (n14969, n_263, n_9882);
  and g22167 (n14970, pi0152, n_9969);
  not g22168 (n_10110, n14969);
  and g22169 (n14971, n_1362, n_10110);
  not g22170 (n_10111, n14970);
  and g22171 (n14972, n_10111, n14971);
  not g22172 (n_10112, n14968);
  and g22173 (n14973, pi0216, n_10112);
  not g22174 (n_10113, n14972);
  and g22175 (n14974, n_10113, n14973);
  not g22176 (n_10114, n14974);
  and g22177 (n14975, n6379, n_10114);
  not g22178 (n_10115, n14956);
  and g22179 (n14976, n_10115, n14975);
  not g22180 (n_10116, n14960);
  and g22181 (n14977, n9572, n_10116);
  not g22182 (n_10117, n14976);
  and g22183 (n14978, n_10117, n14977);
  and g22184 (n14979, n_4165, n_9764);
  and g22185 (n14980, n6197, n14655);
  not g22186 (n_10118, n14980);
  and g22187 (n14981, n_10094, n_10118);
  not g22188 (n_10119, n14979);
  not g22189 (n_10120, n14981);
  and g22190 (n14982, n_10119, n_10120);
  and g22191 (n14983, n_299, n14982);
  and g22192 (n14984, n2521, n7551);
  and g22193 (n14985, pi0174, n14984);
  not g22194 (n_10121, n14985);
  and g22195 (n14986, n_10080, n_10121);
  not g22196 (n_10122, n14983);
  and g22197 (n14987, n_10122, n14986);
  not g22198 (n_10123, n14987);
  and g22199 (n14988, n_6015, n_10123);
  and g22200 (n14989, n7551, n14949);
  and g22201 (n14990, pi0224, n_10106);
  not g22202 (n_10124, n14990);
  and g22203 (n14991, n6405, n_10124);
  not g22204 (n_10125, n14991);
  and g22205 (n14992, n_9764, n_10125);
  not g22206 (n_10126, n14989);
  not g22207 (n_10127, n14992);
  and g22208 (n14993, n_10126, n_10127);
  and g22209 (n14994, n_299, n14993);
  and g22210 (n14995, pi0224, n14965);
  not g22211 (n_10128, n14995);
  and g22212 (n14996, n6405, n_10128);
  and g22213 (n14997, n7551, n14951);
  not g22214 (n_10129, n14997);
  and g22215 (n14998, n14996, n_10129);
  not g22216 (n_10130, n14998);
  and g22217 (n14999, n_9757, n_10130);
  not g22218 (n_10131, n14999);
  and g22219 (n15000, pi0174, n_10131);
  not g22220 (n_10132, n14994);
  and g22221 (n15001, pi0193, n_10132);
  not g22222 (n_10133, n15000);
  and g22223 (n15002, n_10133, n15001);
  not g22224 (n_10134, n14764);
  and g22225 (n15003, n_4165, n_10134);
  not g22226 (n_10135, n15003);
  and g22227 (n15004, n2521, n_10135);
  and g22228 (n15005, pi0174, n15004);
  and g22229 (n15006, pi0224, n_9882);
  and g22230 (n15007, n_219, n14981);
  not g22231 (n_10136, n15006);
  and g22232 (n15008, n6405, n_10136);
  not g22233 (n_10137, n15007);
  and g22234 (n15009, n_10137, n15008);
  not g22235 (n_10138, n15009);
  and g22236 (n15010, n_9902, n_10138);
  not g22237 (n_10139, n15010);
  and g22238 (n15011, n_299, n_10139);
  not g22239 (n_10140, n15005);
  and g22240 (n15012, n_5790, n_10140);
  not g22241 (n_10141, n15011);
  and g22242 (n15013, n_10141, n15012);
  not g22243 (n_10142, n15013);
  and g22244 (n15014, pi0180, n_10142);
  not g22245 (n_10143, n15002);
  and g22246 (n15015, n_10143, n15014);
  not g22247 (n_10144, n14988);
  and g22248 (n15016, n_234, n_10144);
  not g22249 (n_10145, n15015);
  and g22250 (n15017, n_10145, n15016);
  not g22251 (n_10146, n14959);
  not g22252 (n_10147, n14978);
  and g22253 (n15018, n_10146, n_10147);
  not g22254 (n_10148, n15017);
  and g22255 (n15019, n_10148, n15018);
  not g22256 (n_10149, n15019);
  and g22257 (n15020, pi0232, n_10149);
  not g22258 (n_10150, n15020);
  and g22259 (n15021, n14945, n_10150);
  not g22260 (n_10151, n14939);
  and g22261 (n15022, n_161, n_10151);
  not g22262 (n_10152, n15021);
  and g22263 (n15023, n_10152, n15022);
  and g22264 (n15024, pi0038, n_10084);
  not g22265 (n_10153, n15024);
  and g22266 (n15025, n_164, n_10153);
  and g22267 (n15026, n_263, n14521);
  and g22268 (n15027, n_263, n6197);
  not g22269 (n_10154, n15027);
  and g22270 (n15028, n14508, n_10154);
  not g22271 (n_10155, n15026);
  and g22272 (n15029, n_6219, n_10155);
  not g22273 (n_10156, n15028);
  and g22274 (n15030, n_10156, n15029);
  and g22275 (n15031, n_3102, n14508);
  not g22276 (n_10157, n14519);
  not g22277 (n_10158, n15031);
  and g22278 (n15032, n_10157, n_10158);
  not g22279 (n_10159, n15032);
  and g22280 (n15033, n_9782, n_10159);
  and g22281 (n15034, n_263, pi0197);
  not g22282 (n_10160, n15033);
  and g22283 (n15035, n_10160, n15034);
  not g22284 (n_10161, n15030);
  not g22285 (n_10162, n15035);
  and g22286 (n15036, n_10161, n_10162);
  not g22287 (n_10163, n15036);
  and g22288 (n15037, n_10072, n_10163);
  and g22289 (n15038, n_3102, n_9758);
  not g22290 (n_10164, n15038);
  and g22291 (n15039, n_9777, n_10164);
  and g22292 (n15040, n_1362, n15039);
  and g22293 (n15041, n_9757, n_9779);
  and g22294 (n15042, n_9758, n15041);
  not g22295 (n_10165, n15042);
  and g22296 (n15043, pi0172, n_10165);
  not g22302 (n_10168, n15037);
  not g22303 (n_10169, n15046);
  and g22304 (n15047, n_10168, n_10169);
  not g22305 (n_10170, n15047);
  and g22306 (n15048, n9766, n_10170);
  and g22307 (n15049, n14505, n14542);
  not g22308 (n_10171, n15049);
  and g22309 (n15050, n_10164, n_10171);
  and g22310 (n15051, n_263, n15050);
  and g22311 (n15052, n14509, n_9843);
  not g22312 (n_10172, n15052);
  and g22313 (n15053, pi0152, n_10172);
  not g22314 (n_10173, n15051);
  and g22315 (n15054, pi0172, n_10173);
  not g22316 (n_10174, n15053);
  and g22317 (n15055, n_10174, n15054);
  and g22318 (n15056, n_9841, n_10164);
  and g22319 (n15057, pi0152, n15056);
  and g22320 (n15058, n_9822, n_10158);
  not g22321 (n_10175, n15058);
  and g22322 (n15059, n_263, n_10175);
  not g22323 (n_10176, n15059);
  and g22324 (n15060, n_1362, n_10176);
  not g22325 (n_10177, n15057);
  and g22326 (n15061, n_10177, n15060);
  not g22327 (n_10178, n15055);
  and g22328 (n15062, n_6219, n_10178);
  not g22329 (n_10179, n15061);
  and g22330 (n15063, n_10179, n15062);
  and g22331 (n15064, n_9815, n_10164);
  and g22332 (n15065, n_1362, n15064);
  and g22333 (n15066, n_9810, n_10164);
  and g22334 (n15067, pi0172, n15066);
  not g22335 (n_10180, n15067);
  and g22336 (n15068, pi0152, n_10180);
  not g22337 (n_10181, n15065);
  and g22338 (n15069, n_10181, n15068);
  and g22339 (n15070, n6197, n14506);
  not g22340 (n_10182, n15070);
  and g22341 (n15071, n_10159, n_10182);
  and g22342 (n15072, n_263, n_10072);
  not g22343 (n_10183, n15071);
  and g22344 (n15073, n_10183, n15072);
  not g22345 (n_10184, n15073);
  and g22346 (n15074, pi0197, n_10184);
  not g22347 (n_10185, n15069);
  and g22348 (n15075, n_10185, n15074);
  not g22349 (n_10186, n15063);
  and g22350 (n15076, n9760, n_10186);
  not g22351 (n_10187, n15075);
  and g22352 (n15077, n_10187, n15076);
  not g22353 (n_10188, n15048);
  not g22354 (n_10189, n15077);
  and g22355 (n15078, n_10188, n_10189);
  not g22356 (n_10190, n15078);
  and g22357 (n15079, pi0299, n_10190);
  and g22358 (n15080, n_6246, n14508);
  and g22359 (n15081, pi0145, n15039);
  not g22360 (n_10191, n15080);
  and g22361 (n15082, pi0174, n_10191);
  not g22362 (n_10192, n15081);
  and g22363 (n15083, n_10192, n15082);
  and g22364 (n15084, n_9767, n_10158);
  not g22365 (n_10193, n15084);
  and g22366 (n15085, n_6246, n_10193);
  and g22367 (n15086, pi0145, n15033);
  not g22368 (n_10194, n15085);
  and g22369 (n15087, n_299, n_10194);
  not g22370 (n_10195, n15086);
  and g22371 (n15088, n_10195, n15087);
  not g22372 (n_10196, n15083);
  not g22373 (n_10197, n15088);
  and g22374 (n15089, n_10196, n_10197);
  not g22375 (n_10198, n15089);
  and g22376 (n15090, n_5790, n_10198);
  and g22377 (n15091, n_6246, n14537);
  not g22378 (n_10199, n15041);
  not g22379 (n_10200, n15091);
  and g22380 (n15092, n_10199, n_10200);
  not g22381 (n_10201, n15092);
  and g22382 (n15093, n_9758, n_10201);
  not g22383 (n_10202, n15093);
  and g22384 (n15094, pi0174, n_10202);
  and g22385 (n15095, n_9757, n_9755);
  not g22386 (n_10203, n15095);
  and g22387 (n15096, pi0145, n_10203);
  not g22388 (n_10204, n15096);
  and g22389 (n15097, n14542, n_10204);
  not g22390 (n_10205, n15097);
  and g22391 (n15098, n_299, n_10205);
  and g22392 (n15099, n_10164, n15098);
  not g22393 (n_10206, n15099);
  and g22394 (n15100, pi0193, n_10206);
  not g22395 (n_10207, n15094);
  and g22396 (n15101, n_10207, n15100);
  not g22397 (n_10208, n15090);
  not g22398 (n_10209, n15101);
  and g22399 (n15102, n_10208, n_10209);
  not g22400 (n_10210, n15102);
  and g22401 (n15103, n9772, n_10210);
  and g22402 (n15104, pi0193, n15050);
  and g22403 (n15105, n_5790, n_10175);
  not g22404 (n_10211, n15104);
  and g22405 (n15106, n_6246, n_10211);
  not g22406 (n_10212, n15105);
  and g22407 (n15107, n_10212, n15106);
  and g22408 (n15108, pi0145, n_10080);
  and g22409 (n15109, n_10183, n15108);
  not g22410 (n_10213, n15109);
  and g22411 (n15110, n_299, n_10213);
  not g22412 (n_10214, n15107);
  and g22413 (n15111, n_10214, n15110);
  and g22414 (n15112, pi0145, n15066);
  and g22415 (n15113, n_6246, n_10172);
  not g22416 (n_10215, n15113);
  and g22417 (n15114, pi0193, n_10215);
  not g22418 (n_10216, n15112);
  and g22419 (n15115, n_10216, n15114);
  and g22420 (n15116, n_6246, n15056);
  and g22421 (n15117, pi0145, n15064);
  not g22422 (n_10217, n15116);
  and g22423 (n15118, n_5790, n_10217);
  not g22424 (n_10218, n15117);
  and g22425 (n15119, n_10218, n15118);
  not g22426 (n_10219, n15115);
  and g22427 (n15120, pi0174, n_10219);
  not g22428 (n_10220, n15119);
  and g22429 (n15121, n_10220, n15120);
  not g22430 (n_10221, n15111);
  and g22431 (n15122, n9776, n_10221);
  not g22432 (n_10222, n15121);
  and g22433 (n15123, n_10222, n15122);
  not g22434 (n_10223, n15103);
  not g22435 (n_10224, n15123);
  and g22436 (n15124, n_10223, n_10224);
  not g22437 (n_10225, n15124);
  and g22438 (n15125, n_161, n_10225);
  not g22439 (n_10226, n15079);
  not g22440 (n_10227, n15125);
  and g22441 (n15126, n_10226, n_10227);
  not g22442 (n_10228, n15126);
  and g22443 (n15127, n9159, n_10228);
  not g22444 (n_10229, n15023);
  and g22445 (n15128, n_10229, n15025);
  not g22446 (n_10230, n15127);
  and g22447 (n15129, n_10230, n15128);
  not g22448 (n_10231, n14937);
  and g22449 (n15130, n2535, n_10231);
  not g22450 (n_10232, n15129);
  and g22451 (n15131, n_10232, n15130);
  not g22452 (n_10233, n14936);
  and g22458 (n15135, n14456, n_10084);
  not g22459 (n_10236, n15025);
  and g22460 (n15136, n_9744, n_10236);
  and g22461 (n15137, n_9765, n_9843);
  and g22462 (n15138, pi0145, n15137);
  and g22463 (n15139, n14536, n14582);
  not g22464 (n_10237, n15139);
  and g22465 (n15140, n_9765, n_10237);
  and g22466 (n15141, n_6246, n15140);
  not g22467 (n_10238, n15138);
  and g22468 (n15142, n_299, n_10238);
  not g22469 (n_10239, n15141);
  and g22470 (n15143, n_10239, n15142);
  not g22471 (n_10240, n14794);
  and g22472 (n15144, n_9765, n_10240);
  and g22473 (n15145, n_6246, n_9948);
  and g22474 (n15146, n_3102, n_9948);
  not g22475 (n_10241, n15146);
  and g22476 (n15147, n_9764, n_10241);
  and g22477 (n15148, n_9753, n15147);
  not g22478 (n_10242, n15145);
  and g22479 (n15149, n_10242, n15148);
  and g22480 (n15150, n2519, n15149);
  not g22481 (n_10243, n15144);
  and g22482 (n15151, pi0174, n_10243);
  not g22483 (n_10244, n15150);
  and g22484 (n15152, n_10244, n15151);
  not g22485 (n_10245, n15152);
  and g22486 (n15153, pi0193, n_10245);
  not g22487 (n_10246, n15143);
  and g22488 (n15154, n_10246, n15153);
  not g22489 (n_10247, n15149);
  and g22490 (n15155, pi0174, n_10247);
  and g22491 (n15156, n_138, n15138);
  and g22492 (n15157, n_6246, n_9765);
  not g22493 (n_10248, n14785);
  and g22494 (n15158, n_10248, n15157);
  not g22495 (n_10249, n15156);
  and g22496 (n15159, n_299, n_10249);
  not g22497 (n_10250, n15158);
  and g22498 (n15160, n_10250, n15159);
  not g22499 (n_10251, n15155);
  and g22500 (n15161, n_5790, n_10251);
  not g22501 (n_10252, n15160);
  and g22502 (n15162, n_10252, n15161);
  not g22503 (n_10253, n15154);
  and g22504 (n15163, n9772, n_10253);
  not g22505 (n_10254, n15162);
  and g22506 (n15164, n_10254, n15163);
  and g22507 (n15165, pi0145, n_9827);
  and g22508 (n15166, n_299, n_10200);
  and g22509 (n15167, n_6246, pi0174);
  not g22510 (n_10255, n14750);
  and g22511 (n15168, n_10255, n15167);
  not g22512 (n_10256, n15165);
  not g22513 (n_10257, n15168);
  and g22514 (n15169, n_10256, n_10257);
  not g22515 (n_10258, n15166);
  and g22516 (n15170, n_10258, n15169);
  and g22517 (n15171, pi0193, n_9765);
  not g22518 (n_10259, n15170);
  and g22519 (n15172, n_10259, n15171);
  and g22520 (n15173, n_9757, n_9765);
  and g22521 (n15174, pi0145, n14438);
  not g22522 (n_10260, n15174);
  and g22523 (n15175, n_10258, n_10260);
  not g22524 (n_10261, n15175);
  and g22525 (n15176, n15173, n_10261);
  not g22526 (n_10262, n14745);
  and g22527 (n15177, n_9765, n_10262);
  and g22528 (n15178, pi0174, n15177);
  not g22529 (n_10263, n15176);
  not g22530 (n_10264, n15178);
  and g22531 (n15179, n_10263, n_10264);
  not g22532 (n_10265, n15179);
  and g22533 (n15180, n_5790, n_10265);
  not g22534 (n_10266, n15172);
  and g22535 (n15181, n9776, n_10266);
  not g22536 (n_10267, n15180);
  and g22537 (n15182, n_10267, n15181);
  not g22538 (n_10268, n15164);
  not g22539 (n_10269, n15182);
  and g22540 (n15183, n_10268, n_10269);
  not g22541 (n_10270, n15183);
  and g22542 (n15184, n_161, n_10270);
  and g22543 (n15185, n_1362, n14443);
  and g22544 (n15186, n_1362, n15148);
  and g22545 (n15187, n_9765, n_9831);
  and g22546 (n15188, pi0172, n15187);
  not g22547 (n_10271, n15186);
  and g22548 (n15189, pi0152, n_10271);
  not g22549 (n_10272, n15188);
  and g22550 (n15190, n_10272, n15189);
  not g22551 (n_10273, n15137);
  and g22552 (n15191, n_263, n_10273);
  not g22559 (n_10277, n15140);
  and g22560 (n15195, n_263, n_10277);
  and g22561 (n15196, pi0152, n_10243);
  not g22562 (n_10278, n15196);
  and g22563 (n15197, pi0172, n_10278);
  not g22564 (n_10279, n15195);
  and g22565 (n15198, n_10279, n15197);
  and g22566 (n15199, n_263, n14785);
  and g22567 (n15200, n_9763, n_10154);
  not g22568 (n_10280, n15200);
  and g22569 (n15201, n_1362, n_10280);
  not g22570 (n_10281, n15199);
  and g22571 (n15202, n_10281, n15201);
  not g22572 (n_10282, n15198);
  not g22573 (n_10283, n15202);
  and g22574 (n15203, n_10282, n_10283);
  not g22575 (n_10284, n15203);
  and g22576 (n15204, n_6219, n_10284);
  and g22582 (n15208, pi0152, n14597);
  not g22583 (n_10287, n15208);
  and g22584 (n15209, n_9765, n_10287);
  not g22585 (n_10288, n15209);
  and g22586 (n15210, pi0172, n_10288);
  and g22587 (n15211, n_1362, n_10073);
  and g22588 (n15212, n_9834, n15211);
  not g22589 (n_10289, n15210);
  and g22590 (n15213, pi0197, n_10289);
  not g22591 (n_10290, n15212);
  and g22592 (n15214, n_10290, n15213);
  and g22593 (n15215, pi0152, n15177);
  and g22594 (n15216, n_9765, n_9779);
  and g22595 (n15217, n_263, n15216);
  and g22596 (n15218, n_9757, n15217);
  not g22597 (n_10291, n15215);
  and g22598 (n15219, n_1362, n_10291);
  not g22599 (n_10292, n15218);
  and g22600 (n15220, n_10292, n15219);
  and g22601 (n15221, n_9765, n_10255);
  and g22602 (n15222, pi0152, n15221);
  not g22603 (n_10293, n15222);
  and g22604 (n15223, pi0172, n_10293);
  not g22605 (n_10294, n15217);
  and g22606 (n15224, n_10294, n15223);
  not g22607 (n_10295, n15224);
  and g22608 (n15225, n_6219, n_10295);
  not g22609 (n_10296, n15220);
  and g22610 (n15226, n_10296, n15225);
  not g22616 (n_10299, n15207);
  not g22617 (n_10300, n15229);
  and g22618 (n15230, n_10299, n_10300);
  not g22619 (n_10301, n15184);
  and g22620 (n15231, n_10301, n15230);
  not g22621 (n_10302, n15231);
  and g22622 (n15232, n9159, n_10302);
  and g22623 (n15233, n_9724, n14916);
  not g22624 (n_10303, n15233);
  and g22625 (n15234, n_5881, n_10303);
  and g22626 (n15235, n_9876, n_10154);
  and g22627 (n15236, n_263, n14677);
  not g22628 (n_10304, n15235);
  not g22629 (n_10305, n15236);
  and g22630 (n15237, n_10304, n_10305);
  not g22631 (n_10306, n15237);
  and g22632 (n15238, n_1362, n_10306);
  and g22633 (n15239, n_263, n14673);
  and g22634 (n15240, pi0152, n14667);
  not g22635 (n_10307, n15240);
  and g22636 (n15241, pi0172, n_10307);
  not g22637 (n_10308, n15239);
  and g22638 (n15242, n_10308, n15241);
  not g22639 (n_10309, n15238);
  and g22640 (n15243, n9036, n_10309);
  not g22641 (n_10310, n15242);
  and g22642 (n15244, n_10310, n15243);
  not g22643 (n_10311, n15244);
  and g22644 (n15245, n9603, n_10311);
  and g22645 (n15246, pi0152, n_10072);
  and g22646 (n15247, n_9922, n15246);
  and g22647 (n15248, n14684, n15072);
  not g22648 (n_10312, n15247);
  and g22649 (n15249, n9036, n_10312);
  not g22650 (n_10313, n15248);
  and g22651 (n15250, n_10313, n15249);
  not g22652 (n_10314, n15250);
  and g22653 (n15251, n9572, n_10314);
  not g22654 (n_10315, n15245);
  not g22655 (n_10316, n15251);
  and g22656 (n15252, n_10315, n_10316);
  not g22657 (n_10317, n15234);
  not g22658 (n_10318, n15252);
  and g22659 (n15253, n_10317, n_10318);
  and g22660 (n15254, pi0180, n14714);
  and g22661 (n15255, n9051, n14649);
  not g22662 (n_10319, n15255);
  and g22663 (n15256, n14439, n_10319);
  not g22664 (n_10320, n15256);
  and g22665 (n15257, pi0174, n_10320);
  not g22666 (n_10321, n15254);
  and g22667 (n15258, n_10321, n15257);
  and g22668 (n15259, n9051, n14678);
  and g22669 (n15260, n_3102, n_9825);
  not g22670 (n_10322, n15260);
  and g22671 (n15261, n_5891, n_10322);
  and g22672 (n15262, n_138, n15261);
  not g22673 (n_10323, n15259);
  not g22674 (n_10324, n15262);
  and g22675 (n15263, n_10323, n_10324);
  and g22676 (n15264, pi0180, n14683);
  not g22677 (n_10325, n15264);
  and g22678 (n15265, n_299, n_10325);
  and g22679 (n15266, n15263, n15265);
  not g22680 (n_10326, n15258);
  and g22681 (n15267, n_5790, n_10326);
  not g22682 (n_10327, n15266);
  and g22683 (n15268, n_10327, n15267);
  and g22684 (n15269, n_9887, n15261);
  and g22685 (n15270, n9051, n14673);
  not g22686 (n_10328, n15269);
  not g22687 (n_10329, n15270);
  and g22688 (n15271, n_10328, n_10329);
  not g22689 (n_10330, n15271);
  and g22690 (n15272, n_299, n_10330);
  and g22691 (n15273, n_9757, n_10320);
  not g22692 (n_10331, n15273);
  and g22693 (n15274, pi0174, n_10331);
  not g22694 (n_10332, n15274);
  and g22695 (n15275, n_6015, n_10332);
  not g22696 (n_10333, n15272);
  and g22697 (n15276, n_10333, n15275);
  and g22698 (n15277, n9051, n_9890);
  not g22699 (n_10334, n10603);
  and g22700 (n15278, n_10334, n15277);
  not g22701 (n_10335, n15278);
  and g22702 (n15279, n_10328, n_10335);
  not g22703 (n_10336, n15279);
  and g22704 (n15280, n_299, n_10336);
  and g22705 (n15281, n_138, n_9922);
  not g22706 (n_10337, n15281);
  and g22707 (n15282, n6197, n_10337);
  not g22708 (n_10338, n15282);
  and g22709 (n15283, n_10320, n_10338);
  not g22710 (n_10339, n15283);
  and g22711 (n15284, pi0174, n_10339);
  not g22712 (n_10340, n15284);
  and g22713 (n15285, pi0180, n_10340);
  not g22714 (n_10341, n15280);
  and g22715 (n15286, n_10341, n15285);
  not g22716 (n_10342, n15286);
  and g22717 (n15287, pi0193, n_10342);
  not g22718 (n_10343, n15276);
  and g22719 (n15288, n_10343, n15287);
  not g22720 (n_10344, n15268);
  and g22721 (n15289, n_234, n_10344);
  not g22722 (n_10345, n15288);
  and g22723 (n15290, n_10345, n15289);
  not g22724 (n_10346, n15253);
  not g22725 (n_10347, n15290);
  and g22726 (n15291, n_10346, n_10347);
  not g22727 (n_10348, n15291);
  and g22728 (n15292, pi0232, n_10348);
  and g22729 (n15293, n_234, n_10320);
  and g22730 (n15294, n9036, n14649);
  not g22731 (n_10349, n15294);
  and g22732 (n15295, n14439, n_10349);
  not g22733 (n_10350, n15295);
  and g22734 (n15296, pi0299, n_10350);
  not g22735 (n_10351, n15293);
  not g22736 (n_10352, n15296);
  and g22737 (n15297, n_10351, n_10352);
  not g22738 (n_10353, n15297);
  and g22739 (n15298, n_3410, n_10353);
  not g22740 (n_10354, n15298);
  and g22741 (n15299, pi0039, n_10354);
  not g22742 (n_10355, n15292);
  and g22743 (n15300, n_10355, n15299);
  and g22744 (n15301, n_3410, n_9763);
  not g22745 (n_10356, n15301);
  and g22746 (n15302, n_162, n_10356);
  not g22747 (n_10357, n15302);
  and g22748 (n15303, n_161, n_10357);
  not g22749 (n_10358, n15300);
  and g22750 (n15304, n_10358, n15303);
  not g22751 (n_10359, n15136);
  not g22752 (n_10360, n15304);
  and g22753 (n15305, n_10359, n_10360);
  not g22754 (n_10361, n15232);
  and g22755 (n15306, n_10361, n15305);
  and g22756 (n15307, n14468, n_10231);
  not g22757 (n_10362, n15306);
  and g22758 (n15308, n_10362, n15307);
  not g22764 (n_10365, n15311);
  and g22765 (n15312, n_4226, n_10365);
  not g22766 (n_10366, n15134);
  and g22767 (n15313, n_10366, n15312);
  or g22768 (po0282, n14923, n15313);
  and g22769 (n15315, pi0175, n14443);
  and g22770 (n15316, n_301, n14597);
  not g22771 (n_10367, n15315);
  and g22772 (n15317, n_234, n_10367);
  not g22773 (n_10368, n15316);
  and g22774 (n15318, n_10368, n15317);
  and g22775 (n15319, n_138, n_9827);
  not g22776 (n_10369, n10299);
  and g22777 (n15320, n_10369, n_9825);
  not g22778 (n_10370, n15320);
  and g22779 (n15321, n_138, n_10370);
  and g22780 (n15322, pi0153, n14443);
  not g22781 (n_10371, n15321);
  not g22782 (n_10372, n15322);
  and g22783 (n15323, n_10371, n_10372);
  not g22784 (n_10373, n15319);
  not g22785 (n_10374, n15323);
  and g22786 (n15324, n_10373, n_10374);
  not g22787 (n_10375, n15324);
  and g22788 (n15325, pi0299, n_10375);
  not g22789 (n_10376, n15318);
  and g22790 (n15326, pi0232, n_10376);
  not g22791 (n_10377, n15325);
  and g22792 (n15327, n_10377, n15326);
  and g22793 (n15328, n_958, n15327);
  and g22794 (n15329, n_9710, n14435);
  and g22795 (n15330, pi0126, n_9719);
  not g22796 (n_10378, n15329);
  not g22797 (n_10379, n15330);
  and g22798 (n15331, n_10378, n_10379);
  not g22799 (n_10380, n14431);
  not g22800 (n_10381, n15331);
  and g22801 (n15332, n_10380, n_10381);
  and g22802 (n15333, n_958, n14439);
  not g22803 (n_10382, n15332);
  and g22804 (n15334, n_10382, n15333);
  and g22805 (n15335, pi0182, n14714);
  and g22806 (n15336, pi0189, n_10320);
  not g22807 (n_10383, n15335);
  and g22808 (n15337, n_10383, n15336);
  and g22809 (n15338, pi0182, n14683);
  not g22810 (n_10384, n15338);
  and g22811 (n15339, n_301, n_10384);
  and g22812 (n15340, n15263, n15339);
  not g22813 (n_10385, n15337);
  not g22814 (n_10386, n15340);
  and g22815 (n15341, n_10385, n_10386);
  not g22816 (n_10387, n15341);
  and g22817 (n15342, n11765, n_10387);
  and g22818 (n15343, n_301, n_10330);
  and g22819 (n15344, pi0189, n_10331);
  not g22820 (n_10388, n15344);
  and g22821 (n15345, n_7715, n_10388);
  not g22822 (n_10389, n15343);
  and g22823 (n15346, n_10389, n15345);
  and g22824 (n15347, n_301, n_10336);
  and g22825 (n15348, pi0189, n_10339);
  not g22826 (n_10390, n15348);
  and g22827 (n15349, pi0182, n_10390);
  not g22828 (n_10391, n15347);
  and g22829 (n15350, n_10391, n15349);
  not g22830 (n_10392, n15346);
  not g22831 (n_10393, n15350);
  and g22832 (n15351, n_10392, n_10393);
  not g22833 (n_10394, n15351);
  and g22834 (n15352, n11833, n_10394);
  and g22835 (n15353, n_5881, n_10374);
  and g22836 (n15354, n_266, n14684);
  and g22837 (n15355, pi0166, n_9922);
  not g22838 (n_10395, n15354);
  not g22839 (n_10396, n15355);
  and g22840 (n15356, n_10395, n_10396);
  and g22841 (n15357, pi0160, n_10372);
  not g22842 (n_10397, n15356);
  and g22843 (n15358, n_10397, n15357);
  and g22844 (n15359, n_10369, n_9876);
  and g22845 (n15360, n_266, n14677);
  not g22846 (n_10398, n15359);
  not g22847 (n_10399, n15360);
  and g22848 (n15361, n_10398, n_10399);
  not g22849 (n_10400, n15361);
  and g22850 (n15362, n_187, n_10400);
  and g22851 (n15363, n_266, n14673);
  and g22852 (n15364, pi0166, n14667);
  not g22853 (n_10401, n15364);
  and g22854 (n15365, pi0153, n_10401);
  not g22855 (n_10402, n15363);
  and g22856 (n15366, n_10402, n15365);
  not g22857 (n_10403, n15362);
  not g22858 (n_10404, n15366);
  and g22859 (n15367, n_10403, n_10404);
  not g22860 (n_10405, n15367);
  and g22861 (n15368, n_7697, n_10405);
  not g22862 (n_10406, n15358);
  and g22863 (n15369, n9036, n_10406);
  not g22864 (n_10407, n15368);
  and g22865 (n15370, n_10407, n15369);
  not g22866 (n_10408, n15353);
  and g22867 (n15371, pi0299, n_10408);
  not g22868 (n_10409, n15370);
  and g22869 (n15372, n_10409, n15371);
  not g22870 (n_10410, n15342);
  not g22871 (n_10411, n15352);
  and g22872 (n15373, n_10410, n_10411);
  not g22873 (n_10412, n15372);
  and g22874 (n15374, n_10412, n15373);
  not g22875 (n_10413, n15374);
  and g22876 (n15375, pi0232, n_10413);
  not g22877 (n_10414, n15375);
  and g22878 (n15376, n15299, n_10414);
  and g22879 (n15377, n_301, n15173);
  not g22880 (n_10415, n15377);
  and g22881 (n15378, pi0178, n_10415);
  and g22882 (n15379, pi0189, n14516);
  not g22883 (n_10416, n15379);
  and g22884 (n15380, n15378, n_10416);
  and g22885 (n15381, pi0189, n15148);
  and g22886 (n15382, n_9843, n15377);
  not g22887 (n_10417, n15381);
  and g22888 (n15383, n_5708, n_10417);
  not g22889 (n_10418, n15382);
  and g22890 (n15384, n_10418, n15383);
  not g22891 (n_10419, n15380);
  and g22892 (n15385, pi0181, n_10419);
  not g22893 (n_10420, n15384);
  and g22894 (n15386, n_10420, n15385);
  and g22895 (n15387, pi0189, n15177);
  and g22896 (n15388, n_301, n15216);
  not g22897 (n_10421, n15388);
  and g22898 (n15389, pi0178, n_10421);
  not g22899 (n_10422, n15378);
  not g22900 (n_10423, n15389);
  and g22901 (n15390, n_10422, n_10423);
  not g22902 (n_10424, n15387);
  not g22903 (n_10425, n15390);
  and g22904 (n15391, n_10424, n_10425);
  and g22905 (n15392, n_6812, n_9763);
  and g22906 (n15393, n_301, n14785);
  not g22907 (n_10426, n15392);
  not g22908 (n_10427, n15393);
  and g22909 (n15394, n_10426, n_10427);
  not g22910 (n_10428, n15394);
  and g22911 (n15395, n_5708, n_10428);
  not g22912 (n_10429, n15391);
  and g22913 (n15396, n_6429, n_10429);
  not g22914 (n_10430, n15395);
  and g22915 (n15397, n_10430, n15396);
  not g22916 (n_10431, n15386);
  and g22917 (n15398, n11765, n_10431);
  not g22918 (n_10432, n15397);
  and g22919 (n15399, n_10432, n15398);
  and g22920 (n15400, n_301, n_9843);
  and g22921 (n15401, pi0189, n_9831);
  not g22922 (n_10433, n15401);
  and g22923 (n15402, n_5708, n_10433);
  not g22924 (n_10434, n15400);
  and g22925 (n15403, n_10434, n15402);
  and g22926 (n15404, pi0178, n11826);
  and g22927 (n15405, n14596, n15404);
  and g22933 (n15409, pi0189, n15221);
  not g22934 (n_10437, n15409);
  and g22935 (n15410, n15389, n_10437);
  and g22936 (n15411, n_301, n15140);
  and g22937 (n15412, pi0189, n15144);
  not g22938 (n_10438, n15412);
  and g22939 (n15413, n_5708, n_10438);
  not g22940 (n_10439, n15411);
  and g22941 (n15414, n_10439, n15413);
  not g22942 (n_10440, n15410);
  and g22943 (n15415, n_6429, n_10440);
  not g22944 (n_10441, n15414);
  and g22945 (n15416, n_10441, n15415);
  not g22946 (n_10442, n15408);
  and g22947 (n15417, n11833, n_10442);
  not g22948 (n_10443, n15416);
  and g22949 (n15418, n_10443, n15417);
  and g22950 (n15419, pi0166, n14597);
  not g22951 (n_10444, n15419);
  and g22952 (n15420, n_9765, n_10444);
  not g22953 (n_10445, n15420);
  and g22954 (n15421, pi0153, n_10445);
  and g22955 (n15422, n_187, n_10375);
  and g22956 (n15423, n_9834, n15422);
  not g22957 (n_10446, n15421);
  and g22958 (n15424, pi0157, n_10446);
  not g22959 (n_10447, n15423);
  and g22960 (n15425, n_10447, n15424);
  and g22961 (n15426, pi0153, pi0166);
  not g22962 (n_10448, n15187);
  and g22963 (n15427, n_10448, n15426);
  and g22964 (n15428, n_266, n_10273);
  not g22965 (n_10449, n15148);
  and g22966 (n15429, pi0166, n_10449);
  and g22967 (n15430, pi0051, n10299);
  not g22968 (n_10450, n15429);
  not g22969 (n_10451, n15430);
  and g22970 (n15431, n_10450, n_10451);
  not g22971 (n_10452, n15431);
  and g22972 (n15432, n_187, n_10452);
  not g22979 (n_10456, n15425);
  and g22980 (n15436, n9794, n_10456);
  not g22981 (n_10457, n15435);
  and g22982 (n15437, n_10457, n15436);
  not g22983 (n_10458, n15216);
  and g22984 (n15438, n_266, n_10458);
  not g22985 (n_10459, n15177);
  and g22986 (n15439, pi0166, n_10459);
  not g22987 (n_10460, n15439);
  and g22988 (n15440, n_10451, n_10460);
  not g22989 (n_10461, n15440);
  and g22990 (n15441, n_187, n_10461);
  not g22991 (n_10462, n15221);
  and g22992 (n15442, n_10462, n15426);
  and g22999 (n15446, n_266, n_10277);
  and g23000 (n15447, pi0166, n_10243);
  not g23001 (n_10466, n15447);
  and g23002 (n15448, pi0153, n_10466);
  not g23003 (n_10467, n15446);
  and g23004 (n15449, n_10467, n15448);
  and g23005 (n15450, n_266, n14785);
  and g23006 (n15451, n_10369, n_9763);
  not g23007 (n_10468, n15451);
  and g23008 (n15452, n_187, n_10468);
  not g23009 (n_10469, n15450);
  and g23010 (n15453, n_10469, n15452);
  not g23011 (n_10470, n15449);
  not g23012 (n_10471, n15453);
  and g23013 (n15454, n_10470, n_10471);
  not g23014 (n_10472, n15454);
  and g23015 (n15455, n_5686, n_10472);
  not g23016 (n_10473, n15445);
  and g23017 (n15456, n9793, n_10473);
  not g23018 (n_10474, n15455);
  and g23019 (n15457, n_10474, n15456);
  not g23027 (n_10479, n15460);
  and g23028 (n15461, pi0232, n_10479);
  not g23029 (n_10480, n15461);
  and g23030 (n15462, n15302, n_10480);
  not g23031 (n_10481, n15376);
  and g23032 (n15463, n_10382, n_10481);
  not g23033 (n_10482, n15462);
  and g23034 (n15464, n_10482, n15463);
  and g23035 (n15465, n_301, n14982);
  and g23036 (n15466, pi0189, n14984);
  not g23037 (n_10483, n15466);
  and g23038 (n15467, n_7715, n_10483);
  not g23039 (n_10484, n15465);
  and g23040 (n15468, n_10484, n15467);
  and g23041 (n15469, n_9757, n15468);
  and g23042 (n15470, n_301, n14993);
  and g23043 (n15471, pi0189, n_10131);
  not g23044 (n_10485, n15470);
  and g23045 (n15472, pi0182, n_10485);
  not g23046 (n_10486, n15471);
  and g23047 (n15473, n_10486, n15472);
  not g23048 (n_10487, n15469);
  not g23049 (n_10488, n15473);
  and g23050 (n15474, n_10487, n_10488);
  not g23051 (n_10489, n15474);
  and g23052 (n15475, n11833, n_10489);
  and g23053 (n15476, n_301, n_10139);
  and g23054 (n15477, pi0189, n15004);
  not g23055 (n_10490, n15477);
  and g23056 (n15478, pi0182, n_10490);
  not g23057 (n_10491, n15476);
  and g23058 (n15479, n_10491, n15478);
  not g23059 (n_10492, n15468);
  not g23060 (n_10493, n15479);
  and g23061 (n15480, n_10492, n_10493);
  not g23062 (n_10494, n15480);
  and g23063 (n15481, n11765, n_10494);
  and g23064 (n15482, n_7697, pi0216);
  not g23065 (n_10495, n15482);
  and g23066 (n15483, n6379, n_10495);
  not g23067 (n_10496, n15483);
  and g23068 (n15484, n15324, n_10496);
  and g23069 (n15485, n_266, n14659);
  and g23070 (n15486, pi0166, n14776);
  not g23071 (n_10497, n15485);
  and g23072 (n15487, n_187, n_10497);
  not g23073 (n_10498, n15486);
  and g23074 (n15488, n_10498, n15487);
  not g23075 (n_10499, n14965);
  and g23076 (n15489, pi0166, n_10499);
  not g23077 (n_10500, n14962);
  and g23078 (n15490, n_266, n_10500);
  not g23079 (n_10501, n15490);
  and g23080 (n15491, pi0153, n_10501);
  not g23081 (n_10502, n15489);
  and g23082 (n15492, n_10502, n15491);
  not g23083 (n_10503, n15488);
  and g23084 (n15493, pi0160, n_10503);
  not g23085 (n_10504, n15492);
  and g23086 (n15494, n_10504, n15493);
  not g23087 (n_10505, n15494);
  and g23088 (n15495, pi0216, n_10505);
  and g23089 (n15496, n_266, n_10096);
  and g23090 (n15497, pi0166, n_10097);
  not g23091 (n_10506, n15496);
  not g23092 (n_10507, n15497);
  and g23093 (n15498, n_10506, n_10507);
  and g23094 (n15499, pi0051, n_187);
  not g23095 (n_10508, n15498);
  not g23096 (n_10509, n15499);
  and g23097 (n15500, n_10508, n_10509);
  not g23098 (n_10510, n15500);
  and g23099 (n15501, n_20, n_10510);
  not g23100 (n_10511, n15495);
  and g23101 (n15502, n6379, n_10511);
  not g23102 (n_10512, n15501);
  and g23103 (n15503, n_10512, n15502);
  not g23104 (n_10513, n15484);
  and g23105 (n15504, pi0299, n_10513);
  not g23106 (n_10514, n15503);
  and g23107 (n15505, n_10514, n15504);
  not g23108 (n_10515, n15475);
  not g23109 (n_10516, n15481);
  and g23110 (n15506, n_10515, n_10516);
  not g23111 (n_10517, n15505);
  and g23112 (n15507, n_10517, n15506);
  not g23113 (n_10518, n15507);
  and g23114 (n15508, pi0232, n_10518);
  not g23115 (n_10519, n15508);
  and g23116 (n15509, n14945, n_10519);
  and g23117 (n15510, n_187, n15064);
  and g23118 (n15511, pi0153, n15066);
  not g23119 (n_10520, n15511);
  and g23120 (n15512, pi0157, n_10520);
  not g23121 (n_10521, n15510);
  and g23122 (n15513, n_10521, n15512);
  and g23123 (n15514, n_187, n15039);
  and g23124 (n15515, pi0153, n_10165);
  not g23125 (n_10522, n15515);
  and g23126 (n15516, n_5686, n_10522);
  not g23127 (n_10523, n15514);
  and g23128 (n15517, n_10523, n15516);
  not g23129 (n_10524, n15513);
  not g23130 (n_10525, n15517);
  and g23131 (n15518, n_10524, n_10525);
  not g23132 (n_10526, n15518);
  and g23133 (n15519, pi0166, n_10526);
  and g23134 (n15520, pi0157, n15071);
  and g23135 (n15521, n_5686, n15033);
  not g23141 (n_10529, n15519);
  not g23142 (n_10530, n15524);
  and g23143 (n15525, n_10529, n_10530);
  not g23144 (n_10531, n15525);
  and g23145 (n15526, n9794, n_10531);
  and g23146 (n15527, n_266, n15050);
  and g23147 (n15528, pi0166, n_10172);
  not g23148 (n_10532, n15527);
  and g23149 (n15529, pi0153, n_10532);
  not g23150 (n_10533, n15528);
  and g23151 (n15530, n_10533, n15529);
  and g23152 (n15531, pi0166, n15056);
  and g23153 (n15532, n_266, n_10175);
  not g23154 (n_10534, n15532);
  and g23155 (n15533, n_187, n_10534);
  not g23156 (n_10535, n15531);
  and g23157 (n15534, n_10535, n15533);
  not g23158 (n_10536, n15530);
  not g23159 (n_10537, n15534);
  and g23160 (n15535, n_10536, n_10537);
  not g23161 (n_10538, n15535);
  and g23162 (n15536, pi0157, n_10538);
  and g23163 (n15537, pi0166, n14508);
  and g23164 (n15538, n_266, n_10193);
  not g23170 (n_10541, n15536);
  not g23171 (n_10542, n15541);
  and g23172 (n15542, n_10541, n_10542);
  not g23173 (n_10543, n15542);
  and g23174 (n15543, n9793, n_10543);
  and g23175 (n15544, n_301, n_10193);
  and g23176 (n15545, pi0189, n14508);
  not g23177 (n_10544, n15545);
  and g23178 (n15546, n_5708, n_10544);
  and g23179 (n15547, n_9757, n15546);
  not g23180 (n_10545, n15544);
  and g23181 (n15548, n_10545, n15547);
  not g23182 (n_10546, n15548);
  and g23183 (n15549, n_6429, n_10546);
  and g23184 (n15550, pi0189, n_10172);
  and g23185 (n15551, n_301, n15050);
  not g23186 (n_10547, n15551);
  and g23187 (n15552, pi0178, n_10547);
  not g23188 (n_10548, n15550);
  and g23189 (n15553, n_10548, n15552);
  not g23190 (n_10549, n15553);
  and g23191 (n15554, n15549, n_10549);
  and g23192 (n15555, pi0189, n15042);
  and g23193 (n15556, n_301, n_10160);
  and g23194 (n15557, n_9757, n15556);
  not g23195 (n_10550, n15555);
  not g23196 (n_10551, n15557);
  and g23197 (n15558, n_10550, n_10551);
  not g23198 (n_10552, n15558);
  and g23199 (n15559, n_5708, n_10552);
  and g23200 (n15560, n_301, n15071);
  and g23201 (n15561, n15066, n_10415);
  not g23202 (n_10553, n15560);
  and g23203 (n15562, pi0178, n_10553);
  not g23204 (n_10554, n15561);
  and g23205 (n15563, n_10554, n15562);
  not g23206 (n_10555, n15559);
  and g23207 (n15564, pi0181, n_10555);
  not g23208 (n_10556, n15563);
  and g23209 (n15565, n_10556, n15564);
  not g23210 (n_10557, n15554);
  and g23211 (n15566, n11833, n_10557);
  not g23212 (n_10558, n15565);
  and g23213 (n15567, n_10558, n15566);
  and g23214 (n15568, n15084, n15546);
  and g23215 (n15569, n_301, n_10175);
  and g23216 (n15570, pi0189, n15056);
  not g23217 (n_10559, n15569);
  and g23218 (n15571, pi0178, n_10559);
  not g23219 (n_10560, n15570);
  and g23220 (n15572, n_10560, n15571);
  not g23221 (n_10561, n15568);
  and g23222 (n15573, n15549, n_10561);
  not g23223 (n_10562, n15572);
  and g23224 (n15574, n_10562, n15573);
  and g23225 (n15575, pi0189, n15064);
  not g23226 (n_10563, n15575);
  and g23227 (n15576, n_10553, n_10563);
  not g23228 (n_10564, n15576);
  and g23229 (n15577, pi0178, n_10564);
  not g23230 (n_10565, n15039);
  and g23231 (n15578, pi0189, n_10565);
  not g23232 (n_10566, n15556);
  and g23233 (n15579, n_5708, n_10566);
  not g23234 (n_10567, n15578);
  and g23235 (n15580, n_10567, n15579);
  not g23236 (n_10568, n15577);
  not g23237 (n_10569, n15580);
  and g23238 (n15581, n_10568, n_10569);
  not g23239 (n_10570, n15581);
  and g23240 (n15582, pi0181, n_10570);
  not g23241 (n_10571, n15574);
  and g23242 (n15583, n11765, n_10571);
  not g23243 (n_10572, n15582);
  and g23244 (n15584, n_10572, n15583);
  not g23252 (n_10577, n15587);
  and g23253 (n15588, pi0232, n_10577);
  not g23254 (n_10578, n15588);
  and g23255 (n15589, n14939, n_10578);
  not g23256 (n_10579, n15509);
  and g23257 (n15590, n15332, n_10579);
  not g23258 (n_10580, n15589);
  and g23259 (n15591, n_10580, n15590);
  not g23260 (n_10581, n15464);
  and g23261 (n15592, n2608, n_10581);
  not g23262 (n_10582, n15591);
  and g23263 (n15593, n_10582, n15592);
  not g23270 (n_10586, n15327);
  and g23271 (n15597, n14455, n_10586);
  and g23272 (n15598, n_9109, pi0299);
  and g23273 (n15599, n_9132, n_234);
  not g23274 (n_10587, n15598);
  not g23275 (n_10588, n15599);
  and g23276 (n15600, n_10587, n_10588);
  and g23277 (n15601, n7473, n15600);
  not g23278 (n_10589, n15601);
  and g23279 (n15602, pi0087, n_10589);
  not g23280 (n_10590, n15597);
  not g23281 (n_10591, n15602);
  and g23282 (n15603, n_10590, n_10591);
  and g23283 (n15604, n14440, n_10382);
  not g23284 (n_10592, n15603);
  not g23285 (n_10593, n15604);
  and g23286 (n15605, n_10592, n_10593);
  not g23287 (n_10594, n15605);
  and g23288 (n15606, n_4226, n_10594);
  not g23289 (n_10595, n15596);
  and g23290 (n15607, n_10595, n15606);
  and g23291 (n15608, pi0232, n_10373);
  not g23292 (n_10596, n15608);
  and g23293 (n15609, n15332, n_10596);
  and g23294 (n15610, n_3410, n_9724);
  not g23295 (n_10597, n15610);
  and g23296 (n15611, n_10374, n_10597);
  not g23297 (n_10598, n15609);
  and g23298 (n15612, n_10598, n15611);
  not g23299 (n_10599, n15612);
  and g23300 (n15613, n_172, n_10599);
  and g23301 (n15614, pi0087, n_9327);
  not g23302 (n_10600, n15614);
  and g23303 (n15615, po1038, n_10600);
  not g23304 (n_10601, n15613);
  and g23305 (n15616, n_10601, n15615);
  not g23306 (n_10602, n15607);
  not g23307 (n_10603, n15616);
  and g23308 (po0283, n_10602, n_10603);
  and g23309 (n15618, n2537, n8887);
  and g23310 (n15619, n2529, n15618);
  not g23311 (n_10604, n15619);
  and g23312 (n15620, n_824, n_10604);
  not g23313 (n_10605, n15618);
  and g23314 (n15621, n_3243, n_10605);
  and g23315 (n15622, pi0129, n7301);
  and g23316 (n15623, n6323, n15622);
  not g23317 (n_10606, n15623);
  and g23318 (n15624, pi0074, n_10606);
  and g23319 (n15625, pi0054, n2611);
  and g23320 (n15626, n8887, n15625);
  not g23321 (n_10607, pi0129);
  and g23322 (n15627, pi0092, n_10607);
  and g23323 (n15628, pi0075, n15622);
  not g23324 (n_10608, n8965);
  and g23325 (n15629, n_251, n_10608);
  not g23326 (n_10609, n15629);
  and g23327 (n15630, n8887, n_10609);
  not g23328 (n_10610, n2568);
  not g23329 (n_10611, n15630);
  and g23330 (n15631, n_10610, n_10611);
  and g23331 (n15632, pi0129, n6135);
  not g23332 (n_10612, n15632);
  and g23333 (n15633, pi0038, n_10612);
  and g23334 (n15634, pi0039, n8887);
  and g23335 (n15635, n_339, n_628);
  not g23336 (n_10613, n2859);
  and g23337 (n15636, n2788, n_10613);
  not g23338 (n_10614, n15636);
  and g23339 (n15637, n2462, n_10614);
  not g23340 (n_10615, n15637);
  and g23341 (n15638, n2873, n_10615);
  not g23342 (n_10616, n15638);
  and g23343 (n15639, n2785, n_10616);
  not g23344 (n_10617, n15639);
  and g23345 (n15640, n2877, n_10617);
  not g23346 (n_10618, n15640);
  and g23347 (n15641, n2719, n_10618);
  not g23348 (n_10619, n15641);
  and g23349 (n15642, n_333, n_10619);
  not g23350 (n_10620, n15642);
  and g23351 (n15643, n_119, n_10620);
  not g23352 (n_10621, n15643);
  and g23353 (n15644, n2783, n_10621);
  not g23354 (n_10622, n15644);
  and g23355 (n15645, n_122, n_10622);
  not g23356 (n_10623, n15645);
  and g23357 (n15646, n_453, n_10623);
  not g23358 (n_10624, n15646);
  and g23359 (n15647, n_123, n_10624);
  not g23360 (n_10625, n15647);
  and g23361 (n15648, n2775, n_10625);
  not g23362 (n_10626, n15648);
  and g23363 (n15649, n2889, n_10626);
  not g23364 (n_10627, n15649);
  and g23365 (n15650, n_459, n_10627);
  not g23366 (n_10628, n15650);
  and g23367 (n15651, n2765, n_10628);
  not g23368 (n_10629, n15651);
  and g23369 (n15652, n2764, n_10629);
  and g23370 (n15653, po0740, n15652);
  and g23371 (n15654, pi0250, n_4117);
  and g23372 (n15655, n10077, n15654);
  and g23373 (n15656, n2781, n_10622);
  not g23374 (n_10630, n15656);
  and g23375 (n15657, n_453, n_10630);
  not g23376 (n_10631, n15657);
  and g23377 (n15658, n_123, n_10631);
  not g23378 (n_10632, n15658);
  and g23379 (n15659, n2775, n_10632);
  not g23380 (n_10633, n15659);
  and g23381 (n15660, n2889, n_10633);
  not g23382 (n_10634, n15660);
  and g23383 (n15661, n_459, n_10634);
  not g23384 (n_10635, n15661);
  and g23385 (n15662, n2765, n_10635);
  not g23386 (n_10636, n15662);
  and g23387 (n15663, n2764, n_10636);
  and g23388 (n15664, n_3209, n15663);
  not g23389 (n_10637, n15653);
  and g23390 (n15665, n_10637, n15655);
  not g23391 (n_10638, n15664);
  and g23392 (n15666, n_10638, n15665);
  not g23393 (n_10640, pi0127);
  and g23394 (n15667, n_10640, n15652);
  and g23395 (n15668, pi0127, n15663);
  not g23396 (n_10641, n15655);
  not g23397 (n_10642, n15667);
  and g23398 (n15669, n_10641, n_10642);
  not g23399 (n_10643, n15668);
  and g23400 (n15670, n_10643, n15669);
  not g23401 (n_10644, n15666);
  not g23402 (n_10645, n15670);
  and g23403 (n15671, n_10644, n_10645);
  not g23404 (n_10646, n15671);
  and g23405 (n15672, n2757, n_10646);
  not g23406 (n_10647, n15672);
  and g23407 (n15673, n3108, n_10647);
  not g23408 (n_10648, n15673);
  and g23409 (n15674, n2504, n_10648);
  not g23410 (n_10649, n15674);
  and g23411 (n15675, n15635, n_10649);
  not g23412 (n_10650, n15675);
  and g23413 (n15676, n_139, n_10650);
  not g23414 (n_10651, n15676);
  and g23415 (n15677, n_622, n_10651);
  not g23416 (n_10652, n15677);
  and g23417 (n15678, n_138, n_10652);
  not g23418 (n_10653, n15678);
  and g23419 (n15679, n2748, n_10653);
  not g23420 (n_10654, n15679);
  and g23421 (n15680, n3168, n_10654);
  not g23422 (n_10655, n15680);
  and g23423 (n15681, n_348, n_10655);
  not g23424 (n_10656, n15681);
  and g23425 (n15682, n2510, n_10656);
  not g23426 (n_10657, n15682);
  and g23427 (n15683, n3413, n_10657);
  not g23428 (n_10658, n15683);
  and g23429 (n15684, n_144, n_10658);
  not g23434 (n_10660, n15634);
  and g23435 (n15688, n_161, n_10660);
  not g23436 (n_10661, n15687);
  and g23437 (n15689, n_10661, n15688);
  not g23438 (n_10662, n15633);
  not g23439 (n_10663, n15689);
  and g23440 (n15690, n_10662, n_10663);
  not g23441 (n_10664, n15690);
  and g23442 (n15691, n2568, n_10664);
  not g23443 (n_10665, n15631);
  and g23444 (n15692, n_171, n_10665);
  not g23445 (n_10666, n15691);
  and g23446 (n15693, n_10666, n15692);
  not g23447 (n_10667, n15628);
  and g23448 (n15694, n_174, n_10667);
  not g23449 (n_10668, n15693);
  and g23450 (n15695, n_10668, n15694);
  not g23451 (n_10669, n15627);
  and g23452 (n15696, n13654, n_10669);
  not g23453 (n_10670, n15695);
  and g23454 (n15697, n_10670, n15696);
  not g23455 (n_10671, n15626);
  and g23456 (n15698, n_168, n_10671);
  not g23457 (n_10672, n15697);
  and g23458 (n15699, n_10672, n15698);
  not g23459 (n_10673, n15624);
  and g23460 (n15700, n_176, n_10673);
  not g23461 (n_10674, n15699);
  and g23462 (n15701, n_10674, n15700);
  and g23463 (n15702, pi0055, n2570);
  and g23464 (n15703, n15622, n15702);
  not g23465 (n_10675, n15701);
  not g23466 (n_10676, n15703);
  and g23467 (n15704, n_10675, n_10676);
  not g23468 (n_10677, n15704);
  and g23469 (n15705, n_157, n_10677);
  not g23470 (n_10678, n11318);
  and g23471 (n15706, n_7348, n_10678);
  not g23472 (n_10679, n15705);
  and g23473 (n15707, n_10679, n15706);
  not g23474 (n_10680, n15621);
  not g23475 (n_10681, n15707);
  and g23476 (n15708, n_10680, n_10681);
  not g23477 (n_10682, n15708);
  and g23478 (n15709, n3328, n_10682);
  not g23479 (n_10683, n15620);
  and g23480 (n15710, n_3030, n_10683);
  not g23481 (n_10684, n15709);
  and g23482 (po0284, n_10684, n15710);
  and g23483 (n15712, n_3035, n_4025);
  and g23484 (n15713, n8888, n10391);
  and g23485 (n15714, po0740, n15713);
  not g23486 (n_10685, n15713);
  and g23487 (n15715, n_10607, n_10685);
  not g23493 (n_10688, n3418);
  and g23494 (n15719, n_161, n_10688);
  not g23495 (n_10689, n15719);
  and g23496 (n15720, n6137, n_10689);
  and g23497 (n15721, n_3213, n6286);
  not g23498 (n_10690, n15721);
  and g23499 (n15722, n_172, n_10690);
  not g23500 (n_10691, n15720);
  and g23501 (n15723, n_10691, n15722);
  not g23502 (n_10692, n15723);
  and g23503 (n15724, n6133, n_10692);
  not g23504 (n_10693, n15718);
  and g23505 (n15725, n6134, n_10693);
  not g23506 (n_10694, n15724);
  and g23507 (n15726, n_10694, n15725);
  and g23508 (n15727, n_3994, n_4020);
  not g23509 (n_10695, n15726);
  and g23510 (n15728, n_10695, n15727);
  not g23511 (n_10696, n15728);
  and g23512 (n15729, n8879, n_10696);
  not g23513 (n_10697, n15729);
  and g23514 (n15730, n15712, n_10697);
  not g23515 (n_10698, n15730);
  and g23516 (n15731, n_157, n_10698);
  not g23517 (n_10699, n15731);
  and g23518 (n15732, n_3223, n_10699);
  not g23519 (n_10700, n15732);
  and g23520 (n15733, n_158, n_10700);
  not g23521 (n_10701, n15733);
  and g23522 (n15734, n_3227, n_10701);
  not g23523 (n_10702, n15734);
  and g23524 (n15735, n3328, n_10702);
  not g23525 (n_10703, n15735);
  and g23526 (po0286, n6123, n_10703);
  and g23527 (n15737, pi0087, n_6269);
  and g23528 (n15738, n7473, n_5721);
  not g23529 (n_10704, n15738);
  and g23530 (n15739, n14596, n_10704);
  not g23531 (n_10705, n15739);
  and g23532 (n15740, n_10373, n_10705);
  not g23533 (n_10706, n15740);
  and g23534 (n15741, n14455, n_10706);
  not g23535 (n_10707, n15737);
  not g23536 (n_10708, n15741);
  and g23537 (n15742, n_10707, n_10708);
  not g23538 (n_10709, n14440);
  not g23539 (n_10710, n15742);
  and g23540 (n15743, n_10709, n_10710);
  and g23541 (n15744, n_9708, n15329);
  not g23542 (n_10711, n15744);
  and g23543 (n15745, pi0130, n_10711);
  and g23544 (n15746, n_9706, n15744);
  not g23545 (n_10712, n15745);
  not g23546 (n_10713, n15746);
  and g23547 (n15747, n_10712, n_10713);
  not g23548 (n_10714, n14429);
  not g23549 (n_10715, n15747);
  and g23550 (n15748, n_10714, n_10715);
  and g23551 (n15749, pi0100, n15740);
  not g23552 (n_10716, n15749);
  and g23553 (n15750, n2535, n_10716);
  not g23554 (n_10717, n10982);
  and g23555 (n15751, n_10717, n15739);
  and g23556 (n15752, n_138, n_10353);
  not g23557 (n_10718, n15752);
  and g23558 (n15753, n_3410, n_10718);
  not g23559 (n_10719, n15753);
  and g23560 (n15754, n10982, n_10719);
  not g23561 (n_10720, pi0191);
  and g23562 (n15755, n_10720, n_234);
  and g23563 (n15756, n_138, n_10320);
  and g23564 (n15757, pi0140, n15282);
  not g23565 (n_10721, n15757);
  and g23566 (n15758, n15756, n_10721);
  not g23567 (n_10722, n15758);
  and g23568 (n15759, n15755, n_10722);
  and g23569 (n15760, n_138, n15263);
  and g23570 (n15761, pi0140, n14657);
  not g23571 (n_10723, n15761);
  and g23572 (n15762, n15760, n_10723);
  not g23573 (n_10724, n15762);
  and g23574 (n15763, n9020, n_10724);
  and g23575 (n15764, pi0169, n6197);
  and g23576 (n15765, n_5881, n14596);
  not g23577 (n_10725, n15764);
  and g23578 (n15766, n_10725, n15765);
  and g23579 (n15767, pi0162, n9036);
  and g23580 (n15768, n_138, n_9895);
  and g23581 (n15769, n_9878, n15768);
  not g23582 (n_10726, n15769);
  and g23583 (n15770, pi0169, n_10726);
  and g23584 (n15771, n_2027, n_10337);
  not g23585 (n_10727, n15771);
  and g23586 (n15772, n15767, n_10727);
  not g23587 (n_10728, n15770);
  and g23588 (n15773, n_10728, n15772);
  and g23589 (n15774, n_207, n15764);
  and g23590 (n15775, n_9877, n_10725);
  not g23602 (n_10734, n15759);
  not g23603 (n_10735, n15763);
  and g23604 (n15782, n_10734, n_10735);
  not g23605 (n_10736, n15781);
  and g23606 (n15783, n_10736, n15782);
  not g23607 (n_10737, n15783);
  and g23608 (n15784, pi0232, n_10737);
  not g23609 (n_10738, n15784);
  and g23610 (n15785, n15754, n_10738);
  not g23611 (n_10739, n15751);
  and g23612 (n15786, n_164, n_10739);
  not g23613 (n_10740, n15785);
  and g23614 (n15787, n_10740, n15786);
  and g23615 (n15788, n_9740, n15750);
  not g23616 (n_10741, n15787);
  and g23617 (n15789, n_10741, n15788);
  not g23618 (n_10742, n15743);
  not g23619 (n_10743, n15748);
  and g23620 (n15790, n_10742, n_10743);
  not g23621 (n_10744, n15789);
  and g23622 (n15791, n_10744, n15790);
  and g23623 (n15792, n_9893, n_10725);
  and g23624 (n15793, pi0169, n14948);
  not g23625 (n_10745, n15792);
  not g23626 (n_10746, n15793);
  and g23627 (n15794, n_10745, n_10746);
  not g23628 (n_10747, n15794);
  and g23629 (n15795, n_20, n_10747);
  and g23630 (n15796, n_9887, n14962);
  and g23631 (n15797, pi0169, n15796);
  and g23632 (n15798, n_138, n_10107);
  and g23633 (n15799, n_2027, n15798);
  not g23639 (n_10750, n15795);
  not g23640 (n_10751, n15802);
  and g23641 (n15803, n_10750, n_10751);
  not g23642 (n_10752, n15803);
  and g23643 (n15804, n6379, n_10752);
  and g23644 (n15805, pi0169, n14597);
  not g23645 (n_10753, n15805);
  and g23646 (n15806, n_138, n_10753);
  not g23647 (n_10754, n15767);
  and g23648 (n15807, n_4176, n_10754);
  not g23649 (n_10755, n15806);
  and g23650 (n15808, n_10755, n15807);
  not g23651 (n_10756, n15804);
  not g23652 (n_10757, n15808);
  and g23653 (n15809, n_10756, n_10757);
  not g23654 (n_10758, n15809);
  and g23655 (n15810, pi0299, n_10758);
  and g23656 (n15811, n7551, n14675);
  not g23657 (n_10759, n15811);
  and g23658 (n15812, n_138, n_10759);
  and g23659 (n15813, n_6245, n15812);
  and g23660 (n15814, n14675, n14996);
  not g23661 (n_10760, n15814);
  and g23662 (n15815, n_138, n_10760);
  and g23663 (n15816, pi0140, n15815);
  not g23664 (n_10761, n15813);
  and g23665 (n15817, n15755, n_10761);
  not g23666 (n_10762, n15816);
  and g23667 (n15818, n_10762, n15817);
  and g23668 (n15819, n_3102, n_9893);
  not g23669 (n_10763, n15819);
  and g23670 (n15820, n_10095, n_10763);
  not g23671 (n_10764, n15820);
  and g23672 (n15821, n7551, n_10764);
  and g23673 (n15822, n_4165, n_10373);
  not g23674 (n_10765, n15821);
  not g23675 (n_10766, n15822);
  and g23676 (n15823, n_10765, n_10766);
  and g23677 (n15824, n_6245, n15823);
  not g23678 (n_10767, n15796);
  and g23679 (n15825, pi0224, n_10767);
  and g23680 (n15826, n_219, n_10764);
  not g23681 (n_10768, n15825);
  not g23682 (n_10769, n15826);
  and g23683 (n15827, n_10768, n_10769);
  not g23684 (n_10770, n15827);
  and g23685 (n15828, n6405, n_10770);
  and g23686 (n15829, n_9884, n_10373);
  not g23687 (n_10771, n15828);
  not g23688 (n_10772, n15829);
  and g23689 (n15830, n_10771, n_10772);
  and g23690 (n15831, pi0140, n15830);
  not g23691 (n_10773, n15824);
  and g23692 (n15832, n9020, n_10773);
  not g23693 (n_10774, n15831);
  and g23694 (n15833, n_10774, n15832);
  not g23695 (n_10775, n15810);
  not g23696 (n_10776, n15818);
  and g23697 (n15834, n_10775, n_10776);
  not g23698 (n_10777, n15833);
  and g23699 (n15835, n_10777, n15834);
  not g23700 (n_10778, n15835);
  and g23701 (n15836, pi0232, n_10778);
  and g23702 (n15837, n14675, n14942);
  not g23703 (n_10779, n15837);
  and g23704 (n15838, n_138, n_10779);
  not g23705 (n_10780, n15838);
  and g23706 (n15839, n_3410, n_10780);
  not g23707 (n_10781, n15839);
  and g23708 (n15840, pi0039, n_10781);
  not g23709 (n_10782, n15836);
  and g23710 (n15841, n_10782, n15840);
  and g23711 (n15842, n_3410, n_9810);
  not g23712 (n_10783, n15842);
  and g23713 (n15843, n_162, n_10783);
  and g23714 (n15844, n_3102, n14578);
  not g23715 (n_10784, n15844);
  and g23716 (n15845, n_10182, n_10784);
  not g23717 (n_10785, n15845);
  and g23718 (n15846, n_5721, n_10785);
  and g23719 (n15847, n9022, n14578);
  not g23720 (n_10786, n15847);
  and g23721 (n15848, pi0232, n_10786);
  not g23722 (n_10787, n15846);
  and g23723 (n15849, n_10787, n15848);
  not g23724 (n_10788, n15849);
  and g23725 (n15850, n15843, n_10788);
  not g23726 (n_10789, n15841);
  not g23727 (n_10790, n15850);
  and g23728 (n15851, n_10789, n_10790);
  not g23729 (n_10791, n15851);
  and g23730 (n15852, n_161, n_10791);
  and g23731 (n15853, pi0038, n_10706);
  not g23732 (n_10792, n15853);
  and g23733 (n15854, n_164, n_10792);
  not g23734 (n_10793, n15852);
  and g23735 (n15855, n_10793, n15854);
  not g23736 (n_10794, n15855);
  and g23737 (n15856, n15750, n_10794);
  and g23738 (n15857, n15742, n15748);
  not g23739 (n_10795, n15856);
  and g23740 (n15858, n_10795, n15857);
  not g23741 (n_10796, n15791);
  not g23742 (n_10797, n15858);
  and g23743 (n15859, n_10796, n_10797);
  not g23744 (n_10798, n15859);
  and g23745 (n15860, n_4226, n_10798);
  not g23746 (n_10799, n9705);
  and g23747 (n15861, pi0087, n_10799);
  and g23748 (n15862, pi0169, n7473);
  and g23749 (n15863, n_172, n14596);
  not g23750 (n_10800, n15862);
  and g23751 (n15864, n_10800, n15863);
  and g23752 (n15865, n_138, n_172);
  and g23753 (n15866, n_10753, n15865);
  and g23754 (n15867, n15748, n15866);
  not g23761 (n_10804, n15860);
  not g23762 (n_10805, n15870);
  and g23763 (po0287, n_10804, n_10805);
  not g23764 (n_10806, n14009);
  and g23765 (n15872, n_164, n_10806);
  and g23766 (n15873, n_172, n_4013);
  not g23767 (n_10807, n15872);
  and g23768 (n15874, n_10807, n15873);
  not g23769 (n_10808, n15874);
  and g23770 (n15875, n_171, n_10808);
  not g23771 (n_10809, n15875);
  and g23772 (n15876, n_3993, n_10809);
  not g23773 (n_10810, n15876);
  and g23774 (n15877, n_174, n_10810);
  and g23775 (n15878, n8880, n13654);
  not g23776 (n_10811, n15877);
  and g23777 (po0288, n_10811, n15878);
  and g23778 (n15880, pi0164, n14920);
  and g23779 (n15881, pi0051, n_983);
  and g23780 (n15882, n_9173, n_9757);
  not g23781 (n_10812, n15881);
  not g23782 (n_10813, n15882);
  and g23783 (n15883, n_10812, n_10813);
  and g23784 (n15884, n14446, n15883);
  and g23785 (n15885, pi0232, n15884);
  and g23786 (n15886, pi0132, n_10378);
  not g23787 (n_10814, n15886);
  and g23788 (n15887, n_10711, n_10814);
  not g23789 (n_10815, n14430);
  not g23790 (n_10816, n15887);
  and g23791 (n15888, n_10815, n_10816);
  not g23792 (n_10817, n15888);
  and g23793 (n15889, n14439, n_10817);
  not g23794 (n_10818, n15885);
  not g23795 (n_10819, n15889);
  and g23796 (n15890, n_10818, n_10819);
  not g23797 (n_10820, n15890);
  and g23798 (n15891, n_172, n_10820);
  not g23799 (n_10821, n15880);
  and g23800 (n15892, po1038, n_10821);
  not g23801 (n_10822, n15891);
  and g23802 (n15893, n_10822, n15892);
  and g23803 (n15894, pi0173, n14443);
  and g23804 (n15895, pi0190, n14597);
  not g23805 (n_10823, n15894);
  and g23806 (n15896, n_234, n_10823);
  not g23807 (n_10824, n15895);
  and g23808 (n15897, n_10824, n15896);
  not g23809 (n_10825, n15884);
  and g23810 (n15898, pi0299, n_10825);
  not g23811 (n_10826, n15897);
  and g23812 (n15899, pi0232, n_10826);
  not g23813 (n_10827, n15898);
  and g23814 (n15900, n_10827, n15899);
  not g23815 (n_10828, n15900);
  and g23816 (n15901, n14455, n_10828);
  not g23817 (n_10829, n9030);
  and g23818 (n15902, pi0087, n_10829);
  and g23819 (n15903, n_958, n15900);
  and g23820 (n15904, n_9173, n14608);
  and g23821 (n15905, pi0168, n14592);
  not g23822 (n_10830, n15905);
  and g23823 (n15906, n_983, n_10830);
  not g23824 (n_10831, n15904);
  and g23825 (n15907, n_10831, n15906);
  and g23826 (n15908, n_3102, n_9840);
  and g23827 (n15909, pi0168, n_10171);
  not g23828 (n_10832, n15908);
  and g23829 (n15910, n_10832, n15909);
  and g23830 (n15911, n_3102, n14608);
  not g23831 (n_10833, n15911);
  and g23832 (n15912, n14613, n_10833);
  not g23833 (n_10834, n15912);
  and g23834 (n15913, n_2206, n_10834);
  not g23835 (n_10835, n15910);
  and g23836 (n15914, pi0151, n_10835);
  not g23837 (n_10836, n15913);
  and g23838 (n15915, n_10836, n15914);
  not g23839 (n_10837, n15907);
  and g23840 (n15916, n_7697, n_10837);
  not g23841 (n_10838, n15915);
  and g23842 (n15917, n_10838, n15916);
  and g23843 (n15918, pi0151, n14578);
  and g23844 (n15919, n_983, n_9814);
  not g23845 (n_10839, n15918);
  and g23846 (n15920, n_2206, n_10839);
  not g23847 (n_10840, n15919);
  and g23848 (n15921, n_10840, n15920);
  and g23849 (n15922, pi0168, n_10812);
  and g23850 (n15923, n_9756, n15922);
  not g23851 (n_10841, n15923);
  and g23852 (n15924, n6197, n_10841);
  not g23853 (n_10842, n15921);
  and g23854 (n15925, n_10842, n15924);
  and g23855 (n15926, pi0160, n_10832);
  not g23856 (n_10843, n15925);
  and g23857 (n15927, n_10843, n15926);
  not g23858 (n_10844, n15917);
  and g23859 (n15928, pi0299, n_10844);
  not g23860 (n_10845, n15927);
  and g23861 (n15929, n_10845, n15928);
  and g23862 (n15930, pi0190, n_234);
  and g23863 (n15931, pi0051, n_9183);
  and g23864 (n15932, pi0182, n14486);
  not g23865 (n_10846, n15932);
  and g23866 (n15933, n14505, n_10846);
  not g23867 (n_10847, n15931);
  and g23868 (n15934, n6197, n_10847);
  not g23869 (n_10848, n15933);
  and g23870 (n15935, n_10848, n15934);
  not g23871 (n_10849, n15935);
  and g23872 (n15936, n15930, n_10849);
  and g23873 (n15937, n_10833, n15936);
  and g23874 (n15938, n_9199, n_234);
  and g23875 (n15939, n_7715, n14608);
  and g23876 (n15940, pi0182, n_10832);
  and g23877 (n15941, n_9815, n15940);
  not g23878 (n_10850, n15939);
  and g23879 (n15942, n_9183, n_10850);
  not g23880 (n_10851, n15941);
  and g23881 (n15943, n_10851, n15942);
  and g23882 (n15944, n_7715, n_10834);
  and g23883 (n15945, n_9811, n_10833);
  not g23884 (n_10852, n15945);
  and g23885 (n15946, pi0182, n_10852);
  not g23886 (n_10853, n15944);
  and g23887 (n15947, pi0173, n_10853);
  not g23888 (n_10854, n15946);
  and g23889 (n15948, n_10854, n15947);
  not g23890 (n_10855, n15943);
  not g23891 (n_10856, n15948);
  and g23892 (n15949, n_10855, n_10856);
  not g23893 (n_10857, n15949);
  and g23894 (n15950, n15938, n_10857);
  and g23901 (n15954, n_3410, n14608);
  not g23902 (n_10861, n15953);
  not g23903 (n_10862, n15954);
  and g23904 (n15955, n_10861, n_10862);
  not g23905 (n_10863, n15955);
  and g23906 (n15956, n_162, n_10863);
  and g23907 (n15957, n_5709, n14979);
  and g23908 (n15958, pi0183, n_10139);
  and g23909 (n15959, n_5709, n_10120);
  not g23910 (n_10864, n15959);
  and g23911 (n15960, n_9183, n_10864);
  not g23912 (n_10865, n15958);
  and g23913 (n15961, n_10865, n15960);
  and g23914 (n15962, n_5709, n_10126);
  not g23915 (n_10866, n14993);
  and g23916 (n15963, pi0173, n_10866);
  not g23917 (n_10867, n15962);
  and g23918 (n15964, n_10867, n15963);
  not g23919 (n_10868, n15957);
  not g23920 (n_10869, n15964);
  and g23921 (n15965, n_10868, n_10869);
  not g23922 (n_10870, n15961);
  and g23923 (n15966, n_10870, n15965);
  not g23924 (n_10871, n15966);
  and g23925 (n15967, n15930, n_10871);
  and g23926 (n15968, n_5709, n_4165);
  not g23927 (n_10872, n15968);
  and g23928 (n15969, n_9183, n_10872);
  and g23929 (n15970, n15004, n15969);
  and g23930 (n15971, pi0183, n14999);
  and g23931 (n15972, n_5709, n_9757);
  not g23932 (n_10873, n14984);
  and g23933 (n15973, n_10873, n15972);
  not g23934 (n_10874, n15973);
  and g23935 (n15974, pi0173, n_10874);
  not g23936 (n_10875, n15971);
  and g23937 (n15975, n_10875, n15974);
  not g23938 (n_10876, n15970);
  and g23939 (n15976, n15938, n_10876);
  not g23940 (n_10877, n15975);
  and g23941 (n15977, n_10877, n15976);
  and g23942 (n15978, n_5685, pi0216);
  not g23943 (n_10878, n15978);
  and g23944 (n15979, n6379, n_10878);
  not g23945 (n_10879, n15979);
  and g23946 (n15980, n15884, n_10879);
  and g23947 (n15981, n_2206, n14776);
  and g23948 (n15982, pi0168, n14659);
  not g23949 (n_10880, n15982);
  and g23950 (n15983, n_983, n_10880);
  not g23951 (n_10881, n15981);
  and g23952 (n15984, n_10881, n15983);
  and g23953 (n15985, n_2206, n_10499);
  and g23954 (n15986, pi0168, n_10500);
  not g23955 (n_10882, n15986);
  and g23956 (n15987, pi0151, n_10882);
  not g23957 (n_10883, n15985);
  and g23958 (n15988, n_10883, n15987);
  not g23959 (n_10884, n15984);
  and g23960 (n15989, pi0149, n_10884);
  not g23961 (n_10885, n15988);
  and g23962 (n15990, n_10885, n15989);
  not g23963 (n_10886, n15990);
  and g23964 (n15991, pi0216, n_10886);
  and g23965 (n15992, pi0168, n_10096);
  and g23966 (n15993, n_2206, n_10097);
  not g23967 (n_10887, n15992);
  not g23968 (n_10888, n15993);
  and g23969 (n15994, n_10887, n_10888);
  not g23970 (n_10889, n15994);
  and g23971 (n15995, n_10812, n_10889);
  not g23972 (n_10890, n15995);
  and g23973 (n15996, n_20, n_10890);
  not g23974 (n_10891, n15991);
  and g23975 (n15997, n6379, n_10891);
  not g23976 (n_10892, n15996);
  and g23977 (n15998, n_10892, n15997);
  not g23978 (n_10893, n15980);
  and g23979 (n15999, pi0299, n_10893);
  not g23980 (n_10894, n15998);
  and g23981 (n16000, n_10894, n15999);
  not g23982 (n_10895, n15967);
  not g23983 (n_10896, n15977);
  and g23984 (n16001, n_10895, n_10896);
  not g23985 (n_10897, n16000);
  and g23986 (n16002, n_10897, n16001);
  not g23987 (n_10898, n16002);
  and g23988 (n16003, pi0232, n_10898);
  not g23989 (n_10899, n16003);
  and g23990 (n16004, n14945, n_10899);
  not g23991 (n_10900, n15956);
  not g23992 (n_10901, n16004);
  and g23993 (n16005, n_10900, n_10901);
  not g23994 (n_10902, n16005);
  and g23995 (n16006, n2608, n_10902);
  not g23996 (n_10903, n15903);
  and g23997 (n16007, n2535, n_10903);
  not g23998 (n_10904, n16006);
  and g23999 (n16008, n_10904, n16007);
  not g24000 (n_10905, n15902);
  and g24006 (n16012, n14456, n_10828);
  and g24007 (n16013, n_9724, n15898);
  not g24008 (n_10908, n13130);
  not g24009 (n_10909, n16013);
  and g24010 (n16014, n_10908, n_10909);
  not g24011 (n_10910, n14667);
  and g24012 (n16015, n_2206, n_10910);
  and g24013 (n16016, pi0168, n_9891);
  not g24014 (n_10911, n16015);
  and g24015 (n16017, pi0151, n_10911);
  not g24016 (n_10912, n16016);
  and g24017 (n16018, n_10912, n16017);
  and g24018 (n16019, pi0168, n14677);
  and g24019 (n16020, n_9173, n_9876);
  not g24020 (n_10913, n16020);
  and g24021 (n16021, n_983, n_10913);
  not g24022 (n_10914, n16019);
  and g24023 (n16022, n_10914, n16021);
  not g24024 (n_10915, n16022);
  and g24025 (n16023, n_5685, n_10915);
  not g24026 (n_10916, n16018);
  and g24027 (n16024, n_10916, n16023);
  not g24028 (n_10917, n15883);
  and g24029 (n16025, n_9922, n_10917);
  not g24030 (n_10918, n16025);
  and g24031 (n16026, n_2206, n_10918);
  and g24032 (n16027, n_10499, n_10812);
  not g24033 (n_10919, n16027);
  and g24034 (n16028, n_9895, n_10919);
  not g24035 (n_10920, n16028);
  and g24036 (n16029, pi0168, n_10920);
  not g24037 (n_10921, n16026);
  and g24038 (n16030, pi0149, n_10921);
  not g24039 (n_10922, n16029);
  and g24040 (n16031, n_10922, n16030);
  not g24041 (n_10923, n16024);
  and g24042 (n16032, n9036, n_10923);
  not g24043 (n_10924, n16031);
  and g24044 (n16033, n_10924, n16032);
  not g24045 (n_10925, n16014);
  not g24046 (n_10926, n16033);
  and g24047 (n16034, n_10925, n_10926);
  and g24048 (n16035, n_5709, n_10330);
  and g24049 (n16036, pi0183, n_10336);
  not g24050 (n_10927, n16036);
  and g24051 (n16037, pi0173, n_10927);
  not g24052 (n_10928, n16035);
  and g24053 (n16038, n_10928, n16037);
  and g24054 (n16039, pi0183, n14683);
  not g24055 (n_10929, n16039);
  and g24056 (n16040, n_9183, n_10929);
  and g24057 (n16041, n15263, n16040);
  not g24058 (n_10930, n16038);
  not g24059 (n_10931, n16041);
  and g24060 (n16042, n_10930, n_10931);
  not g24061 (n_10932, n16042);
  and g24062 (n16043, n15930, n_10932);
  and g24063 (n16044, pi0183, n14714);
  and g24064 (n16045, n_10823, n15938);
  and g24065 (n16046, n_10320, n16045);
  not g24066 (n_10933, n16044);
  and g24067 (n16047, n_10933, n16046);
  not g24068 (n_10934, n16034);
  not g24069 (n_10935, n16047);
  and g24070 (n16048, n_10934, n_10935);
  not g24071 (n_10936, n16043);
  and g24072 (n16049, n_10936, n16048);
  not g24073 (n_10937, n16049);
  and g24074 (n16050, pi0232, n_10937);
  not g24075 (n_10938, n16050);
  and g24076 (n16051, n_10354, n_10938);
  not g24077 (n_10939, n16051);
  and g24078 (n16052, pi0039, n_10939);
  and g24079 (n16053, n_3410, n14513);
  and g24080 (n16054, pi0182, n15147);
  and g24081 (n16055, n_9948, n16045);
  not g24082 (n_10940, n16054);
  and g24083 (n16056, n_10940, n16055);
  and g24084 (n16057, n_7715, n14537);
  and g24085 (n16058, n_10241, n_10847);
  not g24086 (n_10941, n16057);
  and g24087 (n16059, n_10941, n16058);
  not g24088 (n_10942, n16059);
  and g24089 (n16060, n15930, n_10942);
  and g24090 (n16061, n_2206, n14597);
  not g24091 (n_10943, n16061);
  and g24092 (n16062, n_10241, n_10943);
  not g24093 (n_10944, n16062);
  and g24094 (n16063, pi0151, n_10944);
  and g24095 (n16064, n_983, n_10825);
  not g24096 (n_10945, n15147);
  and g24097 (n16065, n_10945, n16064);
  not g24098 (n_10946, n16063);
  and g24099 (n16066, pi0160, n_10946);
  not g24100 (n_10947, n16065);
  and g24101 (n16067, n_10947, n16066);
  and g24102 (n16068, n_983, n_9948);
  and g24103 (n16069, pi0151, n14750);
  not g24104 (n_10948, n16068);
  and g24105 (n16070, n_2206, n_10948);
  not g24106 (n_10949, n16069);
  and g24107 (n16071, n_10949, n16070);
  and g24108 (n16072, n_983, n14443);
  not g24109 (n_10950, n16072);
  and g24110 (n16073, pi0168, n_10950);
  and g24111 (n16074, n_9779, n16073);
  not g24112 (n_10951, n16071);
  not g24113 (n_10952, n16074);
  and g24114 (n16075, n_10951, n_10952);
  and g24115 (n16076, n_7697, n_10241);
  not g24116 (n_10953, n16075);
  and g24117 (n16077, n_10953, n16076);
  not g24118 (n_10954, n16067);
  and g24119 (n16078, pi0299, n_10954);
  not g24120 (n_10955, n16077);
  and g24121 (n16079, n_10955, n16078);
  not g24128 (n_10959, n16053);
  and g24129 (n16083, n_162, n_10959);
  not g24130 (n_10960, n16082);
  and g24131 (n16084, n_10960, n16083);
  not g24132 (n_10961, n16084);
  and g24133 (n16085, n2608, n_10961);
  not g24134 (n_10962, n16052);
  and g24135 (n16086, n_10962, n16085);
  not g24136 (n_10963, n15333);
  not g24146 (n_10967, n16092);
  and g24147 (n16093, n_4226, n_10967);
  not g24148 (n_10968, n16011);
  and g24149 (n16094, n_10968, n16093);
  or g24150 (po0289, n15893, n16094);
  and g24151 (n16096, n_9716, n_10069);
  and g24152 (n16097, pi0145, n14714);
  not g24153 (n_10969, n16097);
  and g24154 (n16098, n15293, n_10969);
  and g24155 (n16099, pi0197, n14657);
  not g24156 (n_10970, n16099);
  and g24157 (n16100, n15294, n_10970);
  not g24158 (n_10971, n16100);
  and g24159 (n16101, n14439, n_10971);
  not g24160 (n_10972, n16101);
  and g24161 (n16102, pi0299, n_10972);
  not g24162 (n_10973, n16098);
  not g24163 (n_10974, n16102);
  and g24164 (n16103, n_10973, n_10974);
  not g24165 (n_10975, n16103);
  and g24166 (n16104, pi0232, n_10975);
  not g24167 (n_10976, n16104);
  and g24168 (n16105, n15299, n_10976);
  and g24169 (n16106, n_5876, n14503);
  and g24170 (n16107, n_162, n14439);
  not g24171 (n_10977, n16106);
  and g24172 (n16108, n_10977, n16107);
  not g24173 (n_10978, n16108);
  and g24174 (n16109, n_161, n_10978);
  not g24175 (n_10979, n16105);
  and g24176 (n16110, n_10979, n16109);
  not g24177 (n_10980, n16110);
  and g24178 (n16111, n14473, n_10980);
  not g24179 (n_10981, n16111);
  and g24180 (n16112, n14468, n_10981);
  not g24181 (n_10982, n14456);
  not g24182 (n_10983, n16112);
  and g24183 (n16113, n_10982, n_10983);
  not g24184 (n_10984, n16096);
  not g24185 (n_10985, n16113);
  and g24186 (n16114, n_10984, n_10985);
  and g24187 (n16115, n_5709, n_234);
  and g24188 (n16116, n_5685, pi0299);
  not g24189 (n_10986, n16115);
  not g24190 (n_10987, n16116);
  and g24191 (n16117, n_10986, n_10987);
  and g24192 (n16118, n7473, n16117);
  not g24193 (n_10988, n16118);
  and g24194 (n16119, pi0087, n_10988);
  not g24195 (n_10989, n9209);
  and g24196 (n16120, n_10989, n14532);
  and g24197 (n16121, n_3102, n_9775);
  not g24198 (n_10990, n16121);
  and g24199 (n16122, n_9815, n_10990);
  and g24200 (n16123, n9209, n16122);
  not g24206 (n_10993, n5777);
  and g24207 (n16127, n_10993, n_10970);
  not g24208 (n_10994, n16127);
  and g24209 (n16128, n6640, n_10994);
  and g24210 (n16129, n_6246, n_4165);
  not g24211 (n_10995, n16129);
  and g24212 (n16130, n_234, n_10995);
  and g24213 (n16131, n_10135, n16130);
  not g24214 (n_10996, n16128);
  not g24215 (n_10997, n16131);
  and g24216 (n16132, n_10996, n_10997);
  not g24217 (n_10998, n16132);
  and g24218 (n16133, n2521, n_10998);
  not g24219 (n_10999, n16133);
  and g24220 (n16134, pi0232, n_10999);
  not g24221 (n_11000, n16134);
  and g24222 (n16135, n_10093, n_11000);
  not g24223 (n_11001, n16135);
  and g24224 (n16136, pi0039, n_11001);
  and g24225 (n16137, pi0154, pi0232);
  and g24226 (n16138, pi0299, n16137);
  not g24227 (n_11002, n16138);
  and g24228 (n16139, n14532, n_11002);
  and g24229 (n16140, n16122, n16138);
  and g24241 (n16147, n_172, n16096);
  not g24242 (n_11008, n16146);
  and g24243 (n16148, n_11008, n16147);
  not g24244 (n_11009, n16114);
  not g24245 (n_11010, n16119);
  and g24246 (n16149, n_11009, n_11010);
  not g24247 (n_11011, n16148);
  and g24248 (n16150, n_11011, n16149);
  not g24249 (n_11012, n16150);
  and g24250 (n16151, n_4226, n_11012);
  and g24251 (n16152, pi0149, n14920);
  and g24252 (n16153, n14440, n_10984);
  not g24253 (n_11013, n16152);
  and g24254 (n16154, po1038, n_11013);
  not g24255 (n_11014, n16153);
  and g24256 (n16155, n_11014, n16154);
  or g24257 (po0290, n16151, n16155);
  and g24258 (n16157, po1038, n15865);
  and g24259 (n16158, n_9704, n15746);
  and g24260 (n16159, n_9702, n16158);
  not g24261 (n_11015, n16159);
  and g24262 (n16160, pi0134, n_11015);
  not g24263 (n_11016, n16160);
  and g24264 (n16161, n14438, n_11016);
  and g24265 (n16162, pi0171, n6197);
  and g24266 (n16163, n_9825, n16162);
  and g24267 (n16164, pi0232, n16163);
  not g24268 (n_11017, n16164);
  and g24269 (n16165, n16157, n_11017);
  not g24270 (n_11018, n16161);
  and g24271 (n16166, n_11018, n16165);
  and g24272 (n16167, pi0192, n_234);
  and g24273 (n16168, pi0171, pi0299);
  not g24274 (n_11020, n16167);
  not g24275 (n_11021, n16168);
  and g24276 (n16169, n_11020, n_11021);
  not g24277 (n_11022, n16169);
  and g24278 (n16170, n7473, n_11022);
  not g24279 (n_11023, n16170);
  and g24280 (n16171, n14596, n_11023);
  not g24281 (n_11024, n16171);
  and g24282 (n16172, n_10373, n_11024);
  not g24283 (n_11025, n16172);
  and g24284 (n16173, n14455, n_11025);
  and g24285 (n16174, n_958, n16172);
  not g24286 (n_11026, n16174);
  and g24287 (n16175, n2535, n_11026);
  not g24288 (n_11027, n16163);
  and g24289 (n16176, n_138, n_11027);
  and g24290 (n16177, n_5727, pi0216);
  not g24291 (n_11028, n16177);
  and g24292 (n16178, n6379, n_11028);
  not g24293 (n_11029, n16176);
  not g24294 (n_11030, n16178);
  and g24295 (n16179, n_11029, n_11030);
  not g24296 (n_11031, n16162);
  and g24297 (n16180, n_9893, n_11031);
  and g24298 (n16181, pi0171, n14948);
  not g24299 (n_11032, n16180);
  not g24300 (n_11033, n16181);
  and g24301 (n16182, n_11032, n_11033);
  not g24302 (n_11034, n16182);
  and g24303 (n16183, n_20, n_11034);
  and g24304 (n16184, pi0171, n15796);
  and g24305 (n16185, n_1493, n15798);
  not g24311 (n_11037, n16183);
  not g24312 (n_11038, n16188);
  and g24313 (n16189, n_11037, n_11038);
  not g24314 (n_11039, n16189);
  and g24315 (n16190, n6379, n_11039);
  not g24316 (n_11040, n16179);
  not g24317 (n_11041, n16190);
  and g24318 (n16191, n_11040, n_11041);
  not g24319 (n_11042, n16191);
  and g24320 (n16192, pi0299, n_11042);
  not g24321 (n_11043, pi0192);
  and g24322 (n16193, n_11043, n_234);
  not g24323 (n_11044, n15812);
  and g24324 (n16194, n_11044, n16193);
  and g24325 (n16195, pi0039, pi0186);
  not g24326 (n_11045, n15823);
  and g24327 (n16196, n_11045, n16167);
  not g24328 (n_11046, n16194);
  not g24329 (n_11047, n16195);
  and g24330 (n16197, n_11046, n_11047);
  not g24331 (n_11048, n16196);
  and g24332 (n16198, n_11048, n16197);
  not g24333 (n_11049, n15815);
  and g24334 (n16199, n_11049, n16193);
  not g24335 (n_11050, n15830);
  and g24336 (n16200, n_11050, n16167);
  not g24337 (n_11051, n16199);
  and g24338 (n16201, pi0186, n_11051);
  not g24339 (n_11052, n16200);
  and g24340 (n16202, n_11052, n16201);
  not g24341 (n_11053, n16198);
  not g24342 (n_11054, n16202);
  and g24343 (n16203, n_11053, n_11054);
  not g24344 (n_11055, n16192);
  not g24345 (n_11056, n16203);
  and g24346 (n16204, n_11055, n_11056);
  not g24347 (n_11057, n16204);
  and g24348 (n16205, pi0232, n_11057);
  not g24349 (n_11058, n16205);
  and g24350 (n16206, n15840, n_11058);
  and g24351 (n16207, pi0232, n_11022);
  not g24352 (n_11059, n16207);
  and g24353 (n16208, n_9810, n_11059);
  and g24354 (n16209, n15845, n16207);
  not g24355 (n_11060, n16208);
  and g24356 (n16210, n_162, n_11060);
  not g24357 (n_11061, n16209);
  and g24358 (n16211, n_11061, n16210);
  not g24359 (n_11062, n16206);
  and g24360 (n16212, n2608, n_11062);
  not g24361 (n_11063, n16211);
  and g24362 (n16213, n_11063, n16212);
  not g24363 (n_11064, n16213);
  and g24364 (n16214, n16175, n_11064);
  not g24365 (n_11065, n16173);
  and g24366 (n16215, n16160, n_11065);
  not g24367 (n_11066, n16214);
  and g24368 (n16216, n_11066, n16215);
  and g24369 (n16217, n14455, n16171);
  and g24370 (n16218, pi0039, n_5726);
  not g24371 (n_11067, n15760);
  and g24372 (n16219, n_11067, n16167);
  not g24373 (n_11068, n15756);
  and g24374 (n16220, n_11068, n16193);
  not g24375 (n_11069, n16219);
  not g24376 (n_11070, n16220);
  and g24377 (n16221, n_11069, n_11070);
  and g24378 (n16222, n15765, n_11031);
  not g24379 (n_11071, n16222);
  and g24380 (n16223, pi0299, n_11071);
  and g24381 (n16224, n_9877, n_11031);
  and g24382 (n16225, n4192, n6197);
  not g24383 (n_11072, n16224);
  and g24384 (n16226, n9036, n_11072);
  not g24385 (n_11073, n16225);
  and g24386 (n16227, n_11073, n16226);
  not g24387 (n_11074, n16227);
  and g24388 (n16228, n16223, n_11074);
  not g24389 (n_11075, n16228);
  and g24390 (n16229, n16221, n_11075);
  not g24391 (n_11076, n16229);
  and g24392 (n16230, pi0232, n_11076);
  not g24393 (n_11077, n16230);
  and g24394 (n16231, n_10719, n_11077);
  not g24395 (n_11078, n16231);
  and g24396 (n16232, n16218, n_11078);
  and g24397 (n16233, n_162, n_11024);
  and g24398 (n16234, n_9878, n15760);
  not g24399 (n_11079, n16234);
  and g24400 (n16235, n16167, n_11079);
  and g24401 (n16236, n_10338, n15756);
  not g24402 (n_11080, n16236);
  and g24403 (n16237, n16193, n_11080);
  not g24404 (n_11081, n16235);
  not g24405 (n_11082, n16237);
  and g24406 (n16238, n_11081, n_11082);
  and g24407 (n16239, n_11075, n16238);
  not g24408 (n_11083, n16239);
  and g24409 (n16240, pi0232, n_11083);
  not g24410 (n_11084, n16240);
  and g24411 (n16241, n_10719, n_11084);
  not g24412 (n_11085, n16241);
  and g24413 (n16242, n16195, n_11085);
  not g24414 (n_11086, n16233);
  and g24420 (n16246, n_1493, n_10337);
  and g24421 (n16247, pi0171, n_10726);
  not g24422 (n_11089, n16246);
  and g24423 (n16248, n9036, n_11089);
  not g24424 (n_11090, n16247);
  and g24425 (n16249, n_11090, n16248);
  not g24426 (n_11091, n16249);
  and g24427 (n16250, n16223, n_11091);
  not g24428 (n_11092, n16250);
  and g24429 (n16251, n16221, n_11092);
  not g24430 (n_11093, n16251);
  and g24431 (n16252, pi0232, n_11093);
  not g24432 (n_11094, n16252);
  and g24433 (n16253, n_10719, n_11094);
  not g24434 (n_11095, n16253);
  and g24435 (n16254, n16218, n_11095);
  and g24436 (n16255, n16238, n_11092);
  not g24437 (n_11096, n16255);
  and g24438 (n16256, pi0232, n_11096);
  not g24439 (n_11097, n16256);
  and g24440 (n16257, n_10719, n_11097);
  not g24441 (n_11098, n16257);
  and g24442 (n16258, n16195, n_11098);
  not g24448 (n_11101, n16245);
  and g24449 (n16262, n2608, n_11101);
  not g24450 (n_11102, n16261);
  and g24451 (n16263, n_11102, n16262);
  and g24452 (n16264, n_10963, n16175);
  not g24453 (n_11103, n16263);
  and g24454 (n16265, n_11103, n16264);
  not g24455 (n_11104, n16217);
  and g24456 (n16266, n_11016, n_11104);
  not g24457 (n_11105, n16265);
  and g24458 (n16267, n_11105, n16266);
  not g24459 (n_11106, n16216);
  and g24460 (n16268, n_4226, n_11106);
  not g24461 (n_11107, n16267);
  and g24462 (n16269, n_11107, n16268);
  or g24463 (po0291, n16166, n16269);
  not g24464 (n_11108, n16158);
  and g24465 (n16271, pi0135, n_11108);
  and g24466 (n16272, pi0134, n16159);
  not g24467 (n_11109, n16271);
  not g24468 (n_11110, n16272);
  and g24469 (n16273, n_11109, n_11110);
  and g24470 (n16274, pi0170, n6197);
  and g24471 (n16275, n10598, n16274);
  not g24472 (n_11111, n16275);
  and g24473 (n16276, n14596, n_11111);
  and g24474 (n16277, pi0194, n9193);
  not g24475 (n_11113, n16277);
  and g24476 (n16278, n16276, n_11113);
  and g24477 (n16279, n14455, n16278);
  and g24478 (n16280, pi0185, n15282);
  not g24479 (n_11114, n16280);
  and g24480 (n16281, n15756, n_11114);
  and g24481 (n16282, n_10717, n16276);
  not g24482 (n_11115, pi0194);
  not g24483 (n_11116, n16282);
  and g24484 (n16283, n_11115, n_11116);
  not g24485 (n_11117, n16281);
  and g24486 (n16284, n_11117, n16283);
  and g24487 (n16285, n_9132, n15760);
  and g24488 (n16286, pi0170, n7473);
  not g24489 (n_11118, n9193);
  not g24490 (n_11119, n16286);
  and g24491 (n16287, n_11118, n_11119);
  and g24492 (n16288, n14596, n16287);
  and g24493 (n16289, n_10717, n16288);
  not g24494 (n_11120, n16289);
  and g24495 (n16290, pi0194, n_11120);
  and g24496 (n16291, n_11079, n16290);
  not g24497 (n_11121, n16285);
  and g24498 (n16292, n_11121, n16291);
  not g24499 (n_11122, n16284);
  not g24500 (n_11123, n16292);
  and g24501 (n16293, n_11122, n_11123);
  not g24502 (n_11124, n16293);
  and g24503 (n16294, n_234, n_11124);
  not g24504 (n_11125, n16274);
  and g24505 (n16295, n15765, n_11125);
  and g24506 (n16296, pi0150, pi0299);
  and g24507 (n16297, n_1673, n_10337);
  and g24508 (n16298, pi0170, n_10726);
  not g24509 (n_11126, n16297);
  and g24510 (n16299, n9036, n_11126);
  not g24511 (n_11127, n16298);
  and g24512 (n16300, n_11127, n16299);
  not g24513 (n_11128, n16300);
  and g24514 (n16301, n16296, n_11128);
  and g24515 (n16302, n_9877, n_11125);
  and g24516 (n16303, n4415, n6197);
  not g24517 (n_11129, n16302);
  and g24518 (n16304, n9036, n_11129);
  not g24519 (n_11130, n16303);
  and g24520 (n16305, n_11130, n16304);
  not g24521 (n_11131, n16305);
  and g24522 (n16306, n15598, n_11131);
  not g24523 (n_11132, n16301);
  not g24524 (n_11133, n16306);
  and g24525 (n16307, n_11132, n_11133);
  not g24526 (n_11134, n16283);
  not g24527 (n_11135, n16290);
  and g24528 (n16308, n_11134, n_11135);
  not g24529 (n_11136, n16295);
  not g24530 (n_11137, n16308);
  and g24531 (n16309, n_11136, n_11137);
  not g24532 (n_11138, n16307);
  and g24533 (n16310, n_11138, n16309);
  not g24534 (n_11139, n16294);
  not g24535 (n_11140, n16310);
  and g24536 (n16311, n_11139, n_11140);
  not g24537 (n_11141, n16311);
  and g24538 (n16312, pi0232, n_11141);
  not g24539 (n_11142, n15754);
  and g24540 (n16313, n_11142, n_11137);
  not g24541 (n_11143, n16312);
  not g24542 (n_11144, n16313);
  and g24543 (n16314, n_11143, n_11144);
  not g24544 (n_11145, n16314);
  and g24545 (n16315, n_164, n_11145);
  not g24546 (n_11146, n16278);
  and g24547 (n16316, n_10373, n_11146);
  and g24548 (n16317, pi0100, n16316);
  not g24549 (n_11147, n16317);
  and g24550 (n16318, n2535, n_11147);
  and g24551 (n16319, n_9740, n16318);
  not g24552 (n_11148, n16315);
  and g24553 (n16320, n_11148, n16319);
  not g24554 (n_11149, n16279);
  and g24555 (n16321, n16273, n_11149);
  not g24556 (n_11150, n16320);
  and g24557 (n16322, n_11150, n16321);
  not g24558 (n_11151, n16276);
  and g24559 (n16323, n_10373, n_11151);
  not g24560 (n_11152, n16323);
  and g24561 (n16324, pi0038, n_11152);
  and g24562 (n16325, n_9825, n16274);
  not g24563 (n_11153, n16325);
  and g24564 (n16326, n_138, n_11153);
  and g24565 (n16327, n_9917, n16326);
  and g24566 (n16328, pi0170, n14948);
  and g24567 (n16329, n_9893, n_11125);
  not g24568 (n_11154, n16328);
  and g24569 (n16330, n7570, n_11154);
  not g24570 (n_11155, n16329);
  and g24571 (n16331, n_11155, n16330);
  not g24572 (n_11156, n16331);
  and g24573 (n16332, n_5881, n_11156);
  and g24574 (n16333, n_1673, n15798);
  and g24575 (n16334, pi0170, n15796);
  not g24576 (n_11157, n16334);
  and g24577 (n16335, pi0216, n_11157);
  not g24578 (n_11158, n16333);
  and g24579 (n16336, n_11158, n16335);
  not g24580 (n_11159, n16332);
  not g24581 (n_11160, n16336);
  and g24582 (n16337, n_11159, n_11160);
  not g24583 (n_11161, n16327);
  and g24584 (n16338, n16296, n_11161);
  not g24585 (n_11162, n16337);
  and g24586 (n16339, n_11162, n16338);
  and g24587 (n16340, n_4176, n16326);
  not g24588 (n_11163, n16340);
  and g24589 (n16341, n15598, n_11163);
  and g24590 (n16342, n_11156, n16341);
  not g24591 (n_11164, n16339);
  not g24592 (n_11165, n16342);
  and g24593 (n16343, n_11164, n_11165);
  and g24594 (n16344, n_9132, n15812);
  and g24595 (n16345, pi0185, n15815);
  not g24596 (n_11166, n16344);
  and g24597 (n16346, n_234, n_11166);
  not g24598 (n_11167, n16345);
  and g24599 (n16347, n_11167, n16346);
  not g24600 (n_11168, n16347);
  and g24601 (n16348, n16343, n_11168);
  not g24602 (n_11169, n16348);
  and g24603 (n16349, pi0232, n_11169);
  not g24604 (n_11170, n16349);
  and g24605 (n16350, n15840, n_11170);
  and g24606 (n16351, n_234, n_9810);
  and g24607 (n16352, pi0170, n_10785);
  and g24608 (n16353, n_1673, n14578);
  not g24609 (n_11171, n16353);
  and g24610 (n16354, n10598, n_11171);
  not g24611 (n_11172, n16352);
  and g24612 (n16355, n_11172, n16354);
  not g24613 (n_11173, n16355);
  and g24614 (n16356, n15843, n_11173);
  not g24615 (n_11174, n16351);
  and g24616 (n16357, n_11174, n16356);
  not g24617 (n_11175, n16350);
  not g24618 (n_11176, n16357);
  and g24619 (n16358, n_11175, n_11176);
  not g24620 (n_11177, n16358);
  and g24621 (n16359, n_161, n_11177);
  not g24622 (n_11178, n16324);
  and g24623 (n16360, n_11115, n_11178);
  not g24624 (n_11179, n16359);
  and g24625 (n16361, n_11179, n16360);
  not g24626 (n_11180, n16288);
  and g24627 (n16362, n_10373, n_11180);
  not g24628 (n_11181, n16362);
  and g24629 (n16363, pi0038, n_11181);
  and g24630 (n16364, n_9132, n15823);
  and g24631 (n16365, pi0185, n15830);
  not g24632 (n_11182, n16364);
  and g24633 (n16366, n_234, n_11182);
  not g24634 (n_11183, n16365);
  and g24635 (n16367, n_11183, n16366);
  not g24636 (n_11184, n16367);
  and g24637 (n16368, n16343, n_11184);
  not g24638 (n_11185, n16368);
  and g24639 (n16369, pi0232, n_11185);
  not g24640 (n_11186, n16369);
  and g24641 (n16370, n15840, n_11186);
  and g24642 (n16371, n10602, n15845);
  not g24643 (n_11187, n16371);
  and g24644 (n16372, n16356, n_11187);
  not g24645 (n_11188, n16370);
  not g24646 (n_11189, n16372);
  and g24647 (n16373, n_11188, n_11189);
  not g24648 (n_11190, n16373);
  and g24649 (n16374, n_161, n_11190);
  not g24650 (n_11191, n16363);
  and g24651 (n16375, pi0194, n_11191);
  not g24652 (n_11192, n16374);
  and g24653 (n16376, n_11192, n16375);
  not g24654 (n_11193, n16361);
  not g24655 (n_11194, n16376);
  and g24656 (n16377, n_11193, n_11194);
  not g24657 (n_11195, n16377);
  and g24658 (n16378, n_164, n_11195);
  not g24659 (n_11196, n16378);
  and g24660 (n16379, n16318, n_11196);
  not g24661 (n_11197, n16316);
  and g24662 (n16380, n14455, n_11197);
  not g24663 (n_11198, n16273);
  not g24664 (n_11199, n16380);
  and g24665 (n16381, n_11198, n_11199);
  not g24666 (n_11200, n16379);
  and g24667 (n16382, n_11200, n16381);
  not g24668 (n_11201, n16322);
  and g24669 (n16383, n_4226, n_11201);
  not g24670 (n_11202, n16382);
  and g24671 (n16384, n_11202, n16383);
  and g24672 (n16385, n14438, n16273);
  and g24673 (n16386, n_9825, n16286);
  not g24674 (n_11203, n16386);
  and g24675 (n16387, n16157, n_11203);
  not g24676 (n_11204, n16385);
  and g24677 (n16388, n_11204, n16387);
  or g24678 (po0292, n16384, n16388);
  and g24679 (n16390, pi0136, n_10713);
  not g24680 (n_11205, n16390);
  and g24681 (n16391, n_11108, n_11205);
  not g24682 (n_11206, n14428);
  not g24683 (n_11207, n16391);
  and g24684 (n16392, n_11206, n_11207);
  not g24685 (n_11208, n14596);
  and g24686 (n16393, n_11208, n16392);
  and g24687 (n16394, pi0148, n7473);
  not g24688 (n_11209, n16394);
  and g24689 (n16395, n_9825, n_11209);
  not g24690 (n_11210, n16393);
  not g24691 (n_11211, n16395);
  and g24692 (n16396, n_11210, n_11211);
  not g24693 (n_11212, n16396);
  and g24694 (n16397, n16157, n_11212);
  and g24695 (n16398, n9739, n_9825);
  not g24696 (n_11213, n16398);
  and g24697 (n16399, n_138, n_11213);
  and g24698 (n16400, n14455, n16399);
  not g24699 (n_11214, n16399);
  and g24700 (n16401, n_958, n_11214);
  and g24701 (n16402, n_6260, n_10785);
  and g24702 (n16403, n9738, n14578);
  not g24703 (n_11215, n16403);
  and g24704 (n16404, pi0232, n_11215);
  not g24705 (n_11216, n16402);
  and g24706 (n16405, n_11216, n16404);
  not g24707 (n_11217, n16405);
  and g24708 (n16406, n15843, n_11217);
  and g24709 (n16407, n_7617, n15823);
  and g24710 (n16408, pi0184, n15830);
  not g24711 (n_11218, n16407);
  and g24712 (n16409, n9736, n_11218);
  not g24713 (n_11219, n16408);
  and g24714 (n16410, n_11219, n16409);
  not g24715 (n_11220, pi0141);
  and g24716 (n16411, n_11220, n_234);
  and g24717 (n16412, n_7617, n15812);
  and g24718 (n16413, pi0184, n15815);
  not g24719 (n_11221, n16412);
  and g24720 (n16414, n16411, n_11221);
  not g24721 (n_11222, n16413);
  and g24722 (n16415, n_11222, n16414);
  and g24723 (n16416, n_3084, n13665);
  not g24724 (n_11223, n16416);
  and g24725 (n16417, pi0216, n_11223);
  not g24726 (n_11224, n16417);
  and g24727 (n16418, n6379, n_11224);
  and g24728 (n16419, n14675, n16418);
  and g24729 (n16420, n_138, n_1865);
  not g24730 (n_11225, n16419);
  and g24731 (n16421, n_11225, n16420);
  and g24732 (n16422, n_9917, n15319);
  and g24733 (n16423, n_4176, n_10373);
  not g24734 (n_11226, n16423);
  and g24735 (n16424, n_7591, n_11226);
  and g24736 (n16425, pi0163, n6379);
  and g24737 (n16426, n15796, n16425);
  not g24738 (n_11227, n16422);
  not g24739 (n_11228, n16424);
  and g24740 (n16427, n_11227, n_11228);
  not g24741 (n_11229, n16426);
  and g24742 (n16428, n_11229, n16427);
  and g24743 (n16429, n7570, n_10764);
  not g24744 (n_11230, n16428);
  and g24745 (n16430, pi0148, n_11230);
  not g24746 (n_11231, n16429);
  and g24747 (n16431, n_11231, n16430);
  not g24748 (n_11232, n16421);
  and g24749 (n16432, pi0299, n_11232);
  not g24750 (n_11233, n16431);
  and g24751 (n16433, n_11233, n16432);
  not g24752 (n_11234, n16415);
  not g24753 (n_11235, n16433);
  and g24754 (n16434, n_11234, n_11235);
  not g24755 (n_11236, n16410);
  and g24756 (n16435, n_11236, n16434);
  not g24757 (n_11237, n16435);
  and g24758 (n16436, pi0232, n_11237);
  not g24759 (n_11238, n16436);
  and g24760 (n16437, n15840, n_11238);
  not g24761 (n_11239, n16437);
  and g24762 (n16438, n2608, n_11239);
  not g24763 (n_11240, n16406);
  and g24764 (n16439, n_11240, n16438);
  not g24765 (n_11241, n16401);
  and g24766 (n16440, n2535, n_11241);
  not g24767 (n_11242, n16439);
  and g24768 (n16441, n_11242, n16440);
  not g24769 (n_11243, n16400);
  and g24770 (n16442, n16392, n_11243);
  not g24771 (n_11244, n16441);
  and g24772 (n16443, n_11244, n16442);
  and g24773 (n16444, n_9825, n16400);
  and g24774 (n16445, n_7295, n_9825);
  and g24775 (n16446, n16399, n16445);
  and g24776 (n16447, pi0184, n15282);
  not g24777 (n_11245, n16447);
  and g24778 (n16448, n15756, n_11245);
  not g24779 (n_11246, n16448);
  and g24780 (n16449, n16411, n_11246);
  and g24781 (n16450, pi0184, n14657);
  not g24782 (n_11247, n16450);
  and g24783 (n16451, n15760, n_11247);
  not g24784 (n_11248, n16451);
  and g24785 (n16452, n9736, n_11248);
  and g24786 (n16453, n_3102, n15765);
  and g24787 (n16454, n9036, n15768);
  not g24788 (n_11249, n16453);
  and g24789 (n16455, pi0148, n_11249);
  not g24790 (n_11250, n16454);
  and g24791 (n16456, n_11250, n16455);
  and g24792 (n16457, n_138, n15294);
  not g24793 (n_11251, n16457);
  and g24794 (n16458, n_1865, n_11251);
  not g24795 (n_11252, n16458);
  and g24796 (n16459, n_11223, n_11252);
  and g24797 (n16460, n_1865, n14596);
  not g24798 (n_11253, n16459);
  not g24799 (n_11254, n16460);
  and g24800 (n16461, n_11253, n_11254);
  not g24801 (n_11255, n16456);
  not g24802 (n_11256, n16461);
  and g24803 (n16462, n_11255, n_11256);
  not g24804 (n_11257, n16462);
  and g24805 (n16463, pi0299, n_11257);
  not g24806 (n_11258, n16449);
  not g24807 (n_11259, n16452);
  and g24808 (n16464, n_11258, n_11259);
  not g24809 (n_11260, n16463);
  and g24810 (n16465, n_11260, n16464);
  not g24811 (n_11261, n16465);
  and g24812 (n16466, pi0232, n_11261);
  and g24813 (n16467, n_164, n15754);
  not g24814 (n_11262, n16466);
  and g24815 (n16468, n_11262, n16467);
  not g24816 (n_11263, n16446);
  not g24817 (n_11264, n16468);
  and g24818 (n16469, n_11263, n_11264);
  not g24819 (n_11265, n16469);
  and g24820 (n16470, n2535, n_11265);
  not g24821 (n_11266, n16392);
  not g24822 (n_11267, n16444);
  and g24823 (n16471, n_11266, n_11267);
  not g24824 (n_11268, n16470);
  and g24825 (n16472, n_11268, n16471);
  not g24826 (n_11269, n16472);
  and g24827 (n16473, n_4226, n_11269);
  not g24828 (n_11270, n16443);
  and g24829 (n16474, n_11270, n16473);
  or g24830 (po0293, n16397, n16474);
  and g24831 (n16476, n_162, pi0137);
  and g24832 (n16477, n10368, n14873);
  and g24833 (n16478, n6168, n11568);
  and g24834 (n16479, n_234, n_4226);
  and g24835 (n16480, n_305, n11579);
  and g24836 (n16481, n16479, n16480);
  not g24837 (n_11271, n16478);
  not g24838 (n_11272, n16481);
  and g24839 (n16482, n_11271, n_11272);
  not g24840 (n_11273, n16477);
  not g24841 (n_11274, n16482);
  and g24842 (n16483, n_11273, n_11274);
  and g24843 (n16484, n_271, n11568);
  and g24844 (n16485, po1038, n16484);
  not g24845 (n_11275, n16483);
  not g24846 (n_11276, n16485);
  and g24847 (n16486, n_11275, n_11276);
  not g24848 (n_11277, n16486);
  and g24849 (n16487, n10478, n_11277);
  or g24850 (po0294, n16476, n16487);
  and g24851 (n16489, n_6261, n13910);
  not g24852 (n_11278, n16489);
  and g24853 (n16490, n_162, n_11278);
  and g24854 (n16491, n_3410, n_7430);
  and g24855 (n16492, n6198, n6396);
  and g24856 (n16493, n9051, n16492);
  not g24857 (n_11279, n16493);
  and g24858 (n16494, n9736, n_11279);
  and g24859 (n16495, n_3120, n9737);
  and g24860 (n16496, n_6258, n_7430);
  not g24861 (n_11280, n16494);
  not g24862 (n_11281, n16495);
  and g24863 (n16497, n_11280, n_11281);
  not g24864 (n_11282, n16496);
  and g24865 (n16498, n_11282, n16497);
  not g24866 (n_11283, n16498);
  and g24867 (n16499, pi0232, n_11283);
  not g24868 (n_11284, n16491);
  not g24869 (n_11285, n16499);
  and g24870 (n16500, n_11284, n_11285);
  not g24871 (n_11286, n16500);
  and g24872 (n16501, pi0039, n_11286);
  not g24873 (n_11287, n16490);
  and g24874 (n16502, n10200, n_11287);
  not g24875 (n_11288, n16501);
  and g24876 (n16503, n_11288, n16502);
  and g24877 (n16504, n_5671, n16503);
  not g24878 (n_11289, n9282);
  and g24879 (n16505, n9250, n_11289);
  not g24880 (n_11290, n16505);
  and g24881 (n16506, pi0092, n_11290);
  not g24882 (n_11291, n16506);
  and g24883 (n16507, n2532, n_11291);
  not g24884 (n_11292, n9288);
  and g24885 (n16508, n_171, n_11292);
  not g24886 (n_11293, n9326);
  not g24887 (n_11294, n11892);
  and g24888 (n16509, n_11293, n_11294);
  not g24889 (n_11295, n16509);
  and g24890 (n16510, n9337, n_11295);
  not g24891 (n_11296, n16510);
  and g24892 (n16511, n13815, n_11296);
  and g24893 (n16512, n_3162, n_11293);
  and g24894 (n16513, n9036, n_11295);
  not g24895 (n_11297, n16512);
  and g24896 (n16514, n_11297, n16513);
  not g24897 (n_11298, n16514);
  and g24898 (n16515, n9291, n_11298);
  not g24899 (n_11299, n16511);
  not g24900 (n_11300, n16515);
  and g24901 (n16516, n_11299, n_11300);
  not g24902 (n_11301, n16516);
  and g24903 (n16517, n_3410, n_11301);
  and g24904 (n16518, n_11220, n16511);
  and g24905 (n16519, n_9220, n16510);
  not g24906 (n_11302, n16519);
  and g24907 (n16520, n13815, n_11302);
  and g24908 (n16521, pi0141, n16520);
  and g24909 (n16522, n_5889, n_11295);
  not g24910 (n_11303, n16522);
  and g24911 (n16523, n_5882, n_11303);
  not g24912 (n_11304, n16523);
  and g24913 (n16524, pi0148, n_11304);
  and g24914 (n16525, n_6259, n_11300);
  not g24915 (n_11305, n16524);
  not g24916 (n_11306, n16525);
  and g24917 (n16526, n_11305, n_11306);
  not g24918 (n_11307, n16518);
  not g24919 (n_11308, n16521);
  and g24920 (n16527, n_11307, n_11308);
  not g24921 (n_11309, n16526);
  and g24922 (n16528, n_11309, n16527);
  not g24923 (n_11310, n16528);
  and g24924 (n16529, pi0232, n_11310);
  not g24925 (n_11311, n16517);
  not g24926 (n_11312, n16529);
  and g24927 (n16530, n_11311, n_11312);
  not g24928 (n_11313, n16530);
  and g24929 (n16531, pi0039, n_11313);
  not g24930 (n_11314, n9605);
  and g24931 (n16532, pi0299, n_11314);
  and g24932 (n16533, n_234, n_6440);
  not g24933 (n_11315, n16532);
  and g24934 (n16534, n_3410, n_11315);
  not g24935 (n_11316, n16533);
  and g24936 (n16535, n_11316, n16534);
  not g24937 (n_11317, n16535);
  and g24938 (n16536, n_162, n_11317);
  and g24939 (n16537, n_3102, n_6440);
  not g24940 (n_11318, n16537);
  and g24941 (n16538, n_9187, n_11318);
  not g24942 (n_11319, n16538);
  and g24943 (n16539, n_234, n_11319);
  and g24944 (n16540, pi0141, n16539);
  and g24945 (n16541, pi0148, n6197);
  not g24946 (n_11320, n16541);
  and g24947 (n16542, n_11314, n_11320);
  and g24948 (n16543, pi0148, n13737);
  not g24949 (n_11321, n16542);
  not g24950 (n_11322, n16543);
  and g24951 (n16544, n_11321, n_11322);
  not g24952 (n_11323, n16544);
  and g24953 (n16545, pi0299, n_11323);
  and g24954 (n16546, n_11220, n16533);
  not g24961 (n_11327, n16549);
  and g24962 (n16550, n16536, n_11327);
  not g24963 (n_11328, n16531);
  and g24964 (n16551, n2608, n_11328);
  not g24965 (n_11329, n16550);
  and g24966 (n16552, n_11329, n16551);
  not g24967 (n_11330, n16552);
  and g24968 (n16553, n_172, n_11330);
  not g24969 (n_11331, n16553);
  and g24970 (n16554, n16508, n_11331);
  not g24971 (n_11332, n16554);
  and g24972 (n16555, n_174, n_11332);
  not g24973 (n_11333, n16555);
  and g24974 (n16556, n16507, n_11333);
  not g24975 (n_11334, n16556);
  and g24976 (n16557, n_176, n_11334);
  not g24977 (n_11335, n13686);
  and g24978 (n16558, n9251, n_11335);
  not g24979 (n_11336, n16558);
  and g24980 (n16559, pi0055, n_11336);
  not g24981 (n_11337, n16557);
  not g24982 (n_11338, n16559);
  and g24983 (n16560, n_11337, n_11338);
  not g24984 (n_11339, n16560);
  and g24985 (n16561, n2529, n_11339);
  not g24986 (n_11340, n16561);
  and g24987 (n16562, n9883, n_11340);
  and g24988 (n16563, pi0138, n16562);
  and g24989 (n16564, n_5675, n13664);
  and g24990 (n16565, n_5673, n16564);
  not g24991 (n_11341, n16504);
  not g24992 (n_11342, n16565);
  and g24993 (n16566, n_11341, n_11342);
  not g24994 (n_11343, n16563);
  and g24995 (n16567, n_11343, n16566);
  not g24996 (n_11344, n8974);
  and g24997 (n16568, n_5671, n_11344);
  not g24998 (n_11345, n16568);
  and g24999 (n16569, n16503, n_11345);
  and g25000 (n16570, n16562, n16568);
  not g25001 (n_11346, n16569);
  and g25002 (n16571, n16565, n_11346);
  not g25003 (n_11347, n16570);
  and g25004 (n16572, n_11347, n16571);
  not g25005 (n_11348, n16567);
  not g25006 (n_11349, n16572);
  and g25007 (po0295, n_11348, n_11349);
  and g25008 (n16574, n13910, n_10704);
  not g25009 (n_11350, n16574);
  and g25010 (n16575, n_162, n_11350);
  and g25011 (n16576, n_7426, n15755);
  and g25012 (n16577, n_3120, n9021);
  and g25013 (n16578, n9020, n_11279);
  not g25020 (n_11354, n16581);
  and g25021 (n16582, pi0232, n_11354);
  not g25022 (n_11355, n16582);
  and g25023 (n16583, n_11284, n_11355);
  not g25024 (n_11356, n16583);
  and g25025 (n16584, pi0039, n_11356);
  not g25026 (n_11357, n16575);
  and g25027 (n16585, n10200, n_11357);
  not g25028 (n_11358, n16584);
  and g25029 (n16586, n_11358, n16585);
  and g25030 (n16587, n_5673, n16586);
  and g25031 (n16588, n_2027, n9326);
  not g25032 (n_11359, n16588);
  and g25033 (n16589, n_11303, n_11359);
  not g25034 (n_11360, n16589);
  and g25035 (n16590, n9036, n_11360);
  not g25036 (n_11361, n16590);
  and g25037 (n16591, n9291, n_11361);
  and g25038 (n16592, n_10720, n16511);
  and g25039 (n16593, pi0191, n16520);
  not g25040 (n_11362, n16591);
  not g25041 (n_11363, n16592);
  and g25042 (n16594, n_11362, n_11363);
  not g25043 (n_11364, n16593);
  and g25044 (n16595, n_11364, n16594);
  not g25045 (n_11365, n16595);
  and g25046 (n16596, pi0232, n_11365);
  not g25047 (n_11366, n16596);
  and g25048 (n16597, n_11311, n_11366);
  not g25049 (n_11367, n16597);
  and g25050 (n16598, pi0039, n_11367);
  and g25051 (n16599, pi0191, n16539);
  and g25052 (n16600, n_11314, n_10725);
  and g25053 (n16601, pi0169, n13737);
  not g25054 (n_11368, n16600);
  not g25055 (n_11369, n16601);
  and g25056 (n16602, n_11368, n_11369);
  not g25057 (n_11370, n16602);
  and g25058 (n16603, pi0299, n_11370);
  and g25059 (n16604, n_10720, n16533);
  not g25066 (n_11374, n16607);
  and g25067 (n16608, n16536, n_11374);
  not g25068 (n_11375, n16598);
  and g25069 (n16609, n2608, n_11375);
  not g25070 (n_11376, n16608);
  and g25071 (n16610, n_11376, n16609);
  not g25072 (n_11377, n16610);
  and g25073 (n16611, n_172, n_11377);
  not g25074 (n_11378, n16611);
  and g25075 (n16612, n16508, n_11378);
  not g25076 (n_11379, n16612);
  and g25077 (n16613, n_174, n_11379);
  not g25078 (n_11380, n16613);
  and g25079 (n16614, n16507, n_11380);
  not g25080 (n_11381, n16614);
  and g25081 (n16615, n_176, n_11381);
  not g25082 (n_11382, n16615);
  and g25083 (n16616, n_11338, n_11382);
  not g25084 (n_11383, n16616);
  and g25085 (n16617, n2529, n_11383);
  not g25086 (n_11384, n16617);
  and g25087 (n16618, n9883, n_11384);
  and g25088 (n16619, pi0139, n16618);
  not g25089 (n_11385, n16564);
  not g25090 (n_11386, n16587);
  and g25091 (n16620, n_11385, n_11386);
  not g25092 (n_11387, n16619);
  and g25093 (n16621, n_11387, n16620);
  not g25094 (n_11388, n8975);
  and g25095 (n16622, n_5673, n_11388);
  not g25096 (n_11389, n16622);
  and g25097 (n16623, n16586, n_11389);
  and g25098 (n16624, n16618, n16622);
  not g25099 (n_11390, n16623);
  and g25100 (n16625, n16564, n_11390);
  not g25101 (n_11391, n16624);
  and g25102 (n16626, n_11391, n16625);
  not g25103 (n_11392, n16621);
  not g25104 (n_11393, n16626);
  and g25105 (po0296, n_11392, n_11393);
  not g25106 (n_11395, pi0641);
  and g25107 (n16628, n_11395, pi1158);
  not g25108 (n_11397, pi1158);
  and g25109 (n16629, pi0641, n_11397);
  not g25110 (n_11398, n16628);
  not g25111 (n_11399, n16629);
  and g25112 (n16630, n_11398, n_11399);
  not g25113 (n_11401, n16630);
  and g25114 (n16631, pi0788, n_11401);
  not g25115 (n_11403, pi0648);
  and g25116 (n16632, n_11403, pi1159);
  not g25117 (n_11405, pi1159);
  and g25118 (n16633, pi0648, n_11405);
  not g25119 (n_11406, n16632);
  not g25120 (n_11407, n16633);
  and g25121 (n16634, n_11406, n_11407);
  not g25122 (n_11409, n16634);
  and g25123 (n16635, pi0789, n_11409);
  and g25124 (n16636, pi0627, pi1154);
  not g25125 (n_11412, pi0627);
  not g25126 (n_11413, pi1154);
  and g25127 (n16637, n_11412, n_11413);
  not g25128 (n_11415, n16636);
  and g25129 (n16638, pi0781, n_11415);
  not g25130 (n_11416, n16637);
  and g25131 (n16639, n_11416, n16638);
  not g25132 (n_11417, n2571);
  and g25133 (n16640, pi0140, n_11417);
  and g25134 (n16641, n2926, n6284);
  not g25135 (n_11418, n16641);
  and g25136 (n16642, n_6245, n_11418);
  and g25137 (n16643, pi0665, pi1091);
  not g25138 (n_11420, n16643);
  and g25139 (n16644, pi0680, n_11420);
  and g25140 (n16645, n2926, n16644);
  and g25141 (n16646, n6284, n16645);
  not g25142 (n_11421, n16646);
  and g25143 (n16647, pi0038, n_11421);
  not g25144 (n_11422, n16642);
  and g25145 (n16648, n_11422, n16647);
  not g25146 (n_11423, n6184);
  and g25147 (n16649, n_11423, n6380);
  not g25148 (n_11424, n16649);
  and g25149 (n16650, n_9389, n_11424);
  and g25150 (n16651, pi0120, n_207);
  not g25151 (n_11425, n16650);
  not g25152 (n_11426, n16651);
  and g25153 (n16652, n_11425, n_11426);
  and g25154 (n16653, n2926, n16652);
  and g25155 (n16654, n2603, n16653);
  and g25156 (n16655, n16644, n16654);
  and g25157 (n16656, n_3096, n_3098);
  and g25158 (n16657, n_3093, n16656);
  and g25159 (n16658, n_11420, n16653);
  and g25160 (n16659, n_3138, n16658);
  and g25161 (n16660, n_3126, n_11424);
  and g25162 (n16661, n6380, n_6608);
  and g25163 (n16662, pi1092, n16661);
  not g25164 (n_11427, n11031);
  not g25165 (n_11428, n16662);
  and g25166 (n16663, n_11427, n_11428);
  not g25167 (n_11429, n16660);
  not g25168 (n_11430, n16663);
  and g25169 (n16664, n_11429, n_11430);
  and g25170 (n16665, pi1093, n16664);
  not g25171 (n_11431, n16665);
  and g25172 (n16666, n_9389, n_11431);
  and g25173 (n16667, n2521, n2926);
  not g25174 (n_11432, n16667);
  and g25175 (n16668, pi0120, n_11432);
  not g25176 (n_11433, n16668);
  and g25177 (n16669, n_3128, n_11433);
  not g25178 (n_11434, n16666);
  and g25179 (n16670, n_11434, n16669);
  and g25180 (n16671, n2926, n16649);
  and g25181 (n16672, n2923, n16671);
  and g25182 (n16673, pi0829, n_11428);
  not g25183 (n_11435, n16664);
  and g25184 (n16674, n_3127, n_11435);
  not g25185 (n_11436, n16673);
  and g25186 (n16675, n7517, n_11436);
  not g25187 (n_11437, n16674);
  and g25188 (n16676, n_11437, n16675);
  not g25189 (n_11438, n16672);
  not g25190 (n_11439, n16676);
  and g25191 (n16677, n_11438, n_11439);
  not g25192 (n_11440, n16677);
  and g25193 (n16678, pi1091, n_11440);
  not g25194 (n_11441, n16678);
  and g25195 (n16679, n_9389, n_11441);
  not g25196 (n_11442, n16679);
  and g25197 (n16680, n_11433, n_11442);
  not g25198 (n_11443, n16670);
  not g25199 (n_11444, n16680);
  and g25200 (n16681, n_11443, n_11444);
  and g25201 (n16682, n_3102, n16681);
  not g25202 (n_11445, n16653);
  and g25203 (n16683, n6197, n_11445);
  not g25204 (n_11446, n16682);
  not g25205 (n_11447, n16683);
  and g25206 (n16684, n_11446, n_11447);
  and g25207 (n16685, pi0665, n_11443);
  not g25208 (n_11448, n16681);
  not g25209 (n_11449, n16685);
  and g25210 (n16686, n_11448, n_11449);
  not g25211 (n_11450, n16658);
  not g25212 (n_11451, n16686);
  and g25213 (n16687, n_11450, n_11451);
  not g25214 (n_11452, n16687);
  and g25215 (n16688, n16684, n_11452);
  and g25216 (n16689, n6192, n16688);
  not g25217 (n_11453, n16659);
  not g25218 (n_11454, n16689);
  and g25219 (n16690, n_11453, n_11454);
  not g25220 (n_11455, n16657);
  and g25221 (n16691, n_11455, n16690);
  not g25222 (n_11456, n16688);
  and g25223 (n16692, n16657, n_11456);
  not g25224 (n_11457, n16692);
  and g25225 (n16693, pi0680, n_11457);
  not g25226 (n_11458, n16691);
  and g25227 (n16694, n_11458, n16693);
  not g25228 (n_11459, n16694);
  and g25229 (n16695, n6205, n_11459);
  and g25230 (n16696, n6195, n16686);
  and g25231 (n16697, n6197, n_11448);
  and g25232 (n16698, n_3102, n16653);
  not g25233 (n_11460, n16697);
  not g25234 (n_11461, n16698);
  and g25235 (n16699, n_11460, n_11461);
  and g25236 (n16700, n_3138, n16699);
  and g25237 (n16701, n6192, n16681);
  not g25238 (n_11462, n16700);
  not g25239 (n_11463, n16701);
  and g25240 (n16702, n_11462, n_11463);
  and g25241 (n16703, n16644, n16702);
  and g25242 (n16704, n_11455, n16703);
  not g25243 (n_11464, n16696);
  not g25244 (n_11465, n16704);
  and g25245 (n16705, n_11464, n_11465);
  and g25246 (n16706, n_3119, n16705);
  not g25247 (n_11466, n16695);
  and g25248 (n16707, n_9349, n_11466);
  not g25249 (n_11467, n16706);
  and g25250 (n16708, n_11467, n16707);
  not g25251 (n_11468, n16655);
  not g25252 (n_11469, n16708);
  and g25253 (n16709, n_11468, n_11469);
  not g25254 (n_11470, n16709);
  and g25255 (n16710, n_223, n_11470);
  and g25256 (n16711, n6187, n14205);
  not g25257 (n_11471, n16711);
  and g25258 (n16712, n16667, n_11471);
  not g25259 (n_11472, n16712);
  and g25260 (n16713, pi0120, n_11472);
  not g25261 (n_11473, n16671);
  and g25262 (n16714, n_9389, n_11473);
  not g25263 (n_11474, n16713);
  and g25264 (n16715, pi1091, n_11474);
  not g25265 (n_11475, n16714);
  and g25266 (n16716, n_11475, n16715);
  and g25267 (n16717, pi0120, pi0824);
  and g25268 (n16718, n6187, n16717);
  not g25269 (n_11476, n16718);
  and g25270 (n16719, n16669, n_11476);
  and g25271 (n16720, n_11475, n16719);
  not g25272 (n_11477, n16716);
  not g25273 (n_11478, n16720);
  and g25274 (n16721, n_11477, n_11478);
  not g25275 (n_11479, n16721);
  and g25276 (n16722, n6197, n_11479);
  not g25277 (n_11480, n16722);
  and g25278 (n16723, n_11461, n_11480);
  and g25279 (n16724, n_3119, n16723);
  and g25280 (n16725, n_3102, n16721);
  not g25281 (n_11481, n16725);
  and g25282 (n16726, n16658, n_11481);
  not g25283 (n_11482, n16726);
  and g25284 (n16727, n_11453, n_11482);
  not g25285 (n_11483, n16727);
  and g25286 (n16728, pi0680, n_11483);
  not g25287 (n_11484, n16724);
  and g25288 (n16729, n_11484, n16728);
  and g25289 (n16730, n16657, n_11482);
  not g25290 (n_11485, n16730);
  and g25291 (n16731, pi0223, n_11485);
  and g25292 (n16732, n16729, n16731);
  not g25293 (n_11486, n16710);
  not g25294 (n_11487, n16732);
  and g25295 (n16733, n_11486, n_11487);
  not g25296 (n_11488, n16733);
  and g25297 (n16734, n_234, n_11488);
  and g25298 (n16735, n_3162, n16705);
  and g25299 (n16736, n6242, n_11459);
  not g25300 (n_11489, n16735);
  and g25301 (n16737, n_9350, n_11489);
  not g25302 (n_11490, n16736);
  and g25303 (n16738, n_11490, n16737);
  and g25304 (n16739, n16644, n16653);
  and g25305 (n16740, n3448, n16739);
  not g25306 (n_11491, n16738);
  not g25307 (n_11492, n16740);
  and g25308 (n16741, n_11491, n_11492);
  not g25309 (n_11493, n16741);
  and g25310 (n16742, n_36, n_11493);
  and g25311 (n16743, n_3162, n16723);
  not g25312 (n_11494, n16743);
  and g25313 (n16744, n16728, n_11494);
  and g25314 (n16745, pi0215, n_11485);
  and g25315 (n16746, n16744, n16745);
  not g25316 (n_11495, n16742);
  not g25317 (n_11496, n16746);
  and g25318 (n16747, n_11495, n_11496);
  not g25319 (n_11497, n16747);
  and g25320 (n16748, pi0299, n_11497);
  not g25321 (n_11498, n16734);
  not g25322 (n_11499, n16748);
  and g25323 (n16749, n_11498, n_11499);
  not g25324 (n_11500, n16749);
  and g25325 (n16750, pi0140, n_11500);
  and g25326 (n16751, pi0039, pi0140);
  not g25327 (n_11501, n16644);
  and g25328 (n16752, n_11501, n16654);
  not g25329 (n_11502, pi0680);
  not g25330 (n_11503, n16702);
  and g25331 (n16753, n_11502, n_11503);
  and g25332 (n16754, n16643, n16680);
  and g25333 (n16755, n_3441, n16754);
  and g25334 (n16756, n16643, n16698);
  and g25335 (n16757, n_3138, n16756);
  not g25336 (n_11504, n16755);
  not g25337 (n_11505, n16757);
  and g25338 (n16758, n_11504, n_11505);
  not g25339 (n_11506, n16758);
  and g25340 (n16759, n_11455, n_11506);
  and g25341 (n16760, n16657, n16754);
  not g25342 (n_11507, n16760);
  and g25343 (n16761, pi0680, n_11507);
  not g25344 (n_11508, n16759);
  and g25345 (n16762, n_11508, n16761);
  not g25346 (n_11509, n16753);
  not g25347 (n_11510, n16762);
  and g25348 (n16763, n_11509, n_11510);
  not g25349 (n_11511, n16763);
  and g25350 (n16764, n_3119, n_11511);
  and g25351 (n16765, pi0616, n_11445);
  and g25352 (n16766, pi0614, n_11445);
  not g25353 (n_11512, pi0603);
  and g25354 (n16767, n_11512, n_11445);
  not g25355 (n_11513, n16684);
  and g25356 (n16768, pi0603, n_11513);
  not g25357 (n_11514, n16767);
  not g25358 (n_11515, n16768);
  and g25359 (n16769, n_11514, n_11515);
  not g25360 (n_11516, n16769);
  and g25361 (n16770, n_3087, n_11516);
  not g25362 (n_11517, n6190);
  and g25363 (n16771, n_11517, n_11445);
  not g25364 (n_11518, n16770);
  not g25365 (n_11519, n16771);
  and g25366 (n16772, n_11518, n_11519);
  not g25367 (n_11520, n16772);
  and g25368 (n16773, n_3090, n_11520);
  not g25369 (n_11521, n16766);
  not g25370 (n_11522, n16773);
  and g25371 (n16774, n_11521, n_11522);
  not g25372 (n_11523, n16774);
  and g25373 (n16775, n_3091, n_11523);
  not g25374 (n_11524, n16765);
  not g25375 (n_11525, n16775);
  and g25376 (n16776, n_11524, n_11525);
  not g25377 (n_11526, n16776);
  and g25378 (n16777, n_11502, n_11526);
  and g25379 (n16778, n16643, n16653);
  not g25380 (n_11527, n16778);
  and g25381 (n16779, n6197, n_11527);
  not g25382 (n_11528, n16754);
  and g25383 (n16780, n_3102, n_11528);
  not g25384 (n_11529, n16779);
  not g25385 (n_11530, n16780);
  and g25386 (n16781, n_11529, n_11530);
  and g25387 (n16782, n6192, n16781);
  and g25388 (n16783, n_3138, n16778);
  not g25389 (n_11531, n16783);
  and g25390 (n16784, pi0680, n_11531);
  not g25391 (n_11532, n16782);
  and g25392 (n16785, n_11532, n16784);
  not g25393 (n_11533, n16777);
  not g25394 (n_11534, n16785);
  and g25395 (n16786, n_11533, n_11534);
  and g25396 (n16787, n_11455, n16786);
  not g25397 (n_11535, n16781);
  and g25398 (n16788, pi0680, n_11535);
  not g25399 (n_11536, n16788);
  and g25400 (n16789, n16657, n_11536);
  and g25401 (n16790, n_11533, n16789);
  not g25402 (n_11537, n16787);
  not g25403 (n_11538, n16790);
  and g25404 (n16791, n_11537, n_11538);
  and g25405 (n16792, n6205, n16791);
  not g25406 (n_11539, n16764);
  and g25407 (n16793, n_9349, n_11539);
  not g25408 (n_11540, n16792);
  and g25409 (n16794, n_11540, n16793);
  not g25410 (n_11541, n16752);
  and g25411 (n16795, n_223, n_11541);
  not g25412 (n_11542, n16794);
  and g25413 (n16796, n_11542, n16795);
  and g25414 (n16797, n_11447, n_11481);
  not g25415 (n_11543, n16797);
  and g25416 (n16798, n6190, n_11543);
  not g25417 (n_11544, n16798);
  and g25418 (n16799, n_11519, n_11544);
  not g25419 (n_11545, n16799);
  and g25420 (n16800, n_3090, n_11545);
  not g25421 (n_11546, n16800);
  and g25422 (n16801, n_11521, n_11546);
  not g25423 (n_11547, n16801);
  and g25424 (n16802, n_3091, n_11547);
  not g25425 (n_11548, n16802);
  and g25426 (n16803, n_11524, n_11548);
  not g25427 (n_11549, n16803);
  and g25428 (n16804, n_11502, n_11549);
  and g25429 (n16805, pi0665, n16716);
  not g25430 (n_11550, n16805);
  and g25431 (n16806, n_3102, n_11550);
  not g25432 (n_11551, n16806);
  and g25433 (n16807, n_11529, n_11551);
  not g25434 (n_11552, n16807);
  and g25435 (n16808, n6195, n_11552);
  and g25436 (n16809, n16784, n_11552);
  not g25437 (n_11553, n16808);
  not g25438 (n_11554, n16809);
  and g25439 (n16810, n_11553, n_11554);
  not g25440 (n_11555, n16804);
  and g25441 (n16811, n_11555, n16810);
  and g25442 (n16812, n6205, n16811);
  and g25443 (n16813, n_3091, n16800);
  not g25444 (n_11556, n16723);
  not g25445 (n_11557, n16813);
  and g25446 (n16814, n_11556, n_11557);
  not g25447 (n_11558, n16814);
  and g25448 (n16815, n_11502, n_11558);
  and g25449 (n16816, pi0680, n_11550);
  and g25450 (n16817, n_11505, n16816);
  not g25451 (n_11559, n16815);
  not g25452 (n_11560, n16817);
  and g25453 (n16818, n_11559, n_11560);
  and g25454 (n16819, n16810, n16818);
  and g25455 (n16820, n_3119, n16819);
  not g25456 (n_11561, n16812);
  and g25457 (n16821, pi0223, n_11561);
  not g25458 (n_11562, n16820);
  and g25459 (n16822, n_11562, n16821);
  not g25460 (n_11563, n16796);
  not g25461 (n_11564, n16822);
  and g25462 (n16823, n_11563, n_11564);
  not g25463 (n_11565, n16823);
  and g25464 (n16824, n_234, n_11565);
  and g25465 (n16825, n3448, n16652);
  and g25466 (n16826, n2926, n_11501);
  and g25467 (n16827, n16825, n16826);
  and g25468 (n16828, n_3162, n_11511);
  and g25469 (n16829, n6242, n16791);
  not g25470 (n_11566, n16828);
  and g25471 (n16830, n_9350, n_11566);
  not g25472 (n_11567, n16829);
  and g25473 (n16831, n_11567, n16830);
  not g25474 (n_11568, n16827);
  and g25475 (n16832, n_36, n_11568);
  not g25476 (n_11569, n16831);
  and g25477 (n16833, n_11569, n16832);
  and g25478 (n16834, n6242, n16811);
  and g25479 (n16835, n_3162, n16819);
  not g25480 (n_11570, n16834);
  and g25481 (n16836, pi0215, n_11570);
  not g25482 (n_11571, n16835);
  and g25483 (n16837, n_11571, n16836);
  not g25484 (n_11572, n16833);
  not g25485 (n_11573, n16837);
  and g25486 (n16838, n_11572, n_11573);
  not g25487 (n_11574, n16838);
  and g25488 (n16839, pi0299, n_11574);
  not g25489 (n_11575, n16824);
  not g25490 (n_11576, n16839);
  and g25491 (n16840, n_11575, n_11576);
  and g25492 (n16841, pi0039, n16840);
  not g25493 (n_11577, n16751);
  not g25494 (n_11578, n16841);
  and g25495 (n16842, n_11577, n_11578);
  not g25496 (n_11579, n16750);
  not g25497 (n_11580, n16842);
  and g25498 (n16843, n_11579, n_11580);
  not g25499 (n_11581, n11299);
  and g25500 (n16844, n_53, n_11581);
  and g25501 (n16845, n_47, n_369);
  not g25502 (n_11582, n16844);
  and g25503 (n16846, n_11582, n16845);
  and g25504 (n16847, n7438, n12375);
  and g25505 (n16848, n16846, n16847);
  and g25506 (n16849, n8897, n9141);
  and g25507 (n16850, n16848, n16849);
  not g25508 (n_11583, n16850);
  and g25509 (n16851, n_143, n_11583);
  not g25510 (n_11584, n16851);
  and g25511 (n16852, n10289, n_11584);
  not g25512 (n_11585, n16852);
  and g25513 (n16853, n_280, n_11585);
  and g25514 (n16854, n2763, n2938);
  and g25515 (n16855, n8896, n16848);
  not g25516 (n_11586, n16855);
  and g25517 (n16856, n_108, n_11586);
  and g25518 (n16857, pi0314, n10241);
  not g25519 (n_11587, n16857);
  and g25520 (n16858, n16856, n_11587);
  not g25521 (n_11588, n16858);
  and g25522 (n16859, n16854, n_11588);
  not g25523 (n_11589, n16859);
  and g25524 (n16860, n_130, n_11589);
  and g25525 (n16861, n_143, n10274);
  not g25526 (n_11590, n16860);
  and g25527 (n16862, n_11590, n16861);
  and g25528 (n16863, pi0252, n_346);
  not g25529 (n_11591, n16862);
  and g25530 (n16864, n_11591, n16863);
  not g25531 (n_11592, n16853);
  not g25532 (n_11593, n16864);
  and g25533 (n16865, n_11592, n_11593);
  and g25534 (n16866, n2518, n16865);
  not g25535 (n_11594, n12373);
  and g25536 (n16867, pi1092, n_11594);
  and g25537 (n16868, n16866, n16867);
  not g25538 (n_11595, n16846);
  and g25539 (n16869, n_46, n_11595);
  not g25540 (n_11596, n16869);
  and g25541 (n16870, n11020, n_11596);
  and g25542 (n16871, n_280, n9500);
  and g25543 (n16872, n16870, n16871);
  and g25544 (n16873, n2500, n16870);
  and g25545 (n16874, n_108, n_11587);
  not g25546 (n_11597, n16873);
  and g25547 (n16875, n_11597, n16874);
  not g25548 (n_11598, n16875);
  and g25549 (n16876, n16854, n_11598);
  not g25550 (n_11599, n16876);
  and g25551 (n16877, n_130, n_11599);
  and g25552 (n16878, pi0252, n10274);
  not g25553 (n_11600, n16877);
  and g25554 (n16879, n_11600, n16878);
  not g25555 (n_11601, n16872);
  and g25556 (n16880, n_143, n_11601);
  not g25557 (n_11602, n16879);
  and g25558 (n16881, n_11602, n16880);
  and g25559 (n16882, n7417, n10289);
  not g25560 (n_11603, n16881);
  and g25561 (n16883, n_11603, n16882);
  not g25562 (n_11604, n16868);
  not g25563 (n_11605, n16883);
  and g25564 (n16884, n_11604, n_11605);
  not g25565 (n_11606, n16884);
  and g25566 (n16885, pi1093, n_11606);
  not g25567 (n_11607, n16885);
  and g25568 (n16886, n_489, n_11607);
  and g25569 (n16887, pi1092, n2930);
  and g25570 (po1106, n2923, n16887);
  and g25571 (n16889, n16866, po1106);
  not g25572 (n_11609, n16889);
  and g25573 (n16890, n_538, n_11609);
  not g25574 (n_11610, n16886);
  not g25575 (n_11611, n16890);
  and g25576 (n16891, n_11610, n_11611);
  and g25577 (n16892, n_3128, n16885);
  not g25578 (n_11612, n16891);
  not g25579 (n_11613, n16892);
  and g25580 (n16893, n_11612, n_11613);
  and g25581 (n16894, pi0665, n_11613);
  not g25582 (n_11614, n16893);
  not g25583 (n_11615, n16894);
  and g25584 (n16895, n_11614, n_11615);
  not g25585 (n_11616, n16895);
  and g25586 (n16896, n_305, n_11616);
  and g25587 (n16897, n_874, n_11603);
  not g25588 (n_11617, n16897);
  and g25589 (n16898, n_142, n_11617);
  not g25590 (n_11618, n6485);
  and g25591 (n16899, pi0032, n_11618);
  and g25592 (n16900, n_144, n2932);
  not g25593 (n_11619, n16899);
  and g25594 (n16901, n_11619, n16900);
  not g25595 (n_11620, n16898);
  and g25596 (n16902, n_11620, n16901);
  and g25597 (n16903, pi0824, n16902);
  not g25598 (n_11621, n16903);
  and g25599 (n16904, n_11604, n_11621);
  not g25600 (n_11622, n16904);
  and g25601 (n16905, n7626, n_11622);
  not g25602 (n_11623, n16865);
  and g25603 (n16906, n_142, n_11623);
  not g25604 (n_11624, n16906);
  and g25605 (n16907, n16901, n_11624);
  and g25606 (n16908, n_3126, pi0829);
  and g25607 (n16909, n16907, n16908);
  not g25608 (n_11625, n16909);
  and g25609 (n16910, n16904, n_11625);
  not g25610 (n_11626, n16910);
  and g25611 (n16911, pi1093, n_11626);
  not g25612 (n_11627, n16911);
  and g25613 (n16912, n_489, n_11627);
  not g25614 (n_11628, n16912);
  and g25615 (n16913, n_11611, n_11628);
  not g25616 (n_11629, n16905);
  not g25617 (n_11630, n16913);
  and g25618 (n16914, n_11629, n_11630);
  and g25619 (n16915, pi0665, n_11629);
  not g25620 (n_11631, n16914);
  not g25621 (n_11632, n16915);
  and g25622 (n16916, n_11631, n_11632);
  not g25623 (n_11633, n16916);
  and g25624 (n16917, pi0198, n_11633);
  not g25625 (n_11634, n16896);
  not g25626 (n_11635, n16917);
  and g25627 (n16918, n_11634, n_11635);
  and g25628 (n16919, pi0680, n16918);
  not g25629 (n_11636, n16919);
  and g25630 (n16920, n_234, n_11636);
  and g25631 (n16921, pi0210, n_11633);
  and g25632 (n16922, n_271, n_11616);
  not g25633 (n_11637, n16921);
  not g25634 (n_11638, n16922);
  and g25635 (n16923, n_11637, n_11638);
  and g25636 (n16924, pi0680, n16923);
  not g25637 (n_11639, n16924);
  and g25638 (n16925, pi0299, n_11639);
  not g25639 (n_11640, n16920);
  not g25640 (n_11641, n16925);
  and g25641 (n16926, n_11640, n_11641);
  and g25642 (n16927, pi0140, n16926);
  and g25643 (n16928, n_305, n16893);
  and g25644 (n16929, pi0198, n16914);
  not g25645 (n_11642, n16928);
  not g25646 (n_11643, n16929);
  and g25647 (n16930, n_11642, n_11643);
  and g25648 (n16931, pi0665, n16913);
  not g25649 (n_11644, n16931);
  and g25650 (n16932, pi0198, n_11644);
  and g25651 (n16933, pi0665, n16891);
  not g25652 (n_11645, n16933);
  and g25653 (n16934, n_305, n_11645);
  not g25654 (n_11646, n16932);
  not g25655 (n_11647, n16934);
  and g25656 (n16935, n_11646, n_11647);
  not g25657 (n_11648, n16935);
  and g25658 (n16936, pi0680, n_11648);
  not g25659 (n_11649, n16936);
  and g25660 (n16937, n16930, n_11649);
  not g25661 (n_11650, n16937);
  and g25662 (n16938, n_234, n_11650);
  and g25663 (n16939, n_271, n16893);
  and g25664 (n16940, pi0210, n16914);
  not g25665 (n_11651, n16939);
  not g25666 (n_11652, n16940);
  and g25667 (n16941, n_11651, n_11652);
  and g25668 (n16942, n_271, n_11645);
  and g25669 (n16943, pi0210, n_11644);
  not g25670 (n_11653, n16942);
  not g25671 (n_11654, n16943);
  and g25672 (n16944, n_11653, n_11654);
  not g25673 (n_11655, n16944);
  and g25674 (n16945, pi0680, n_11655);
  not g25675 (n_11656, n16945);
  and g25676 (n16946, n16941, n_11656);
  not g25677 (n_11657, n16946);
  and g25678 (n16947, pi0299, n_11657);
  not g25679 (n_11658, n16938);
  not g25680 (n_11659, n16947);
  and g25681 (n16948, n_11658, n_11659);
  not g25682 (n_11660, n16948);
  and g25683 (n16949, n_6245, n_11660);
  not g25684 (n_11661, n16927);
  and g25685 (n16950, n_162, n_11661);
  not g25686 (n_11662, n16949);
  and g25687 (n16951, n_11662, n16950);
  not g25688 (n_11663, n16843);
  not g25689 (n_11664, n16951);
  and g25690 (n16952, n_11663, n_11664);
  not g25691 (n_11665, n16952);
  and g25692 (n16953, n_161, n_11665);
  not g25693 (n_11667, pi0738);
  not g25694 (n_11668, n16648);
  and g25695 (n16954, n_11667, n_11668);
  not g25696 (n_11669, n16953);
  and g25697 (n16955, n_11669, n16954);
  not g25698 (n_11670, n16941);
  and g25699 (n16956, pi0299, n_11670);
  not g25700 (n_11671, n16930);
  and g25701 (n16957, n_234, n_11671);
  not g25702 (n_11672, n16956);
  not g25703 (n_11673, n16957);
  and g25704 (n16958, n_11672, n_11673);
  not g25705 (n_11674, n16958);
  and g25706 (n16959, n_162, n_11674);
  and g25707 (n16960, pi0681, n_11558);
  and g25708 (n16961, pi0661, n16814);
  not g25709 (n_11675, n6193);
  and g25710 (n16962, n_11675, n_11549);
  and g25711 (n16963, n6193, n16721);
  not g25712 (n_11676, n16963);
  and g25713 (n16964, n_3102, n_11676);
  not g25714 (n_11677, n16962);
  and g25715 (n16965, n_11677, n16964);
  not g25716 (n_11678, n16965);
  and g25717 (n16966, n_11480, n_11678);
  not g25718 (n_11679, n16966);
  and g25719 (n16967, n_3096, n_11679);
  not g25720 (n_11680, n16961);
  and g25721 (n16968, n_3098, n_11680);
  not g25722 (n_11681, n16967);
  and g25723 (n16969, n_11681, n16968);
  not g25724 (n_11682, n16960);
  not g25725 (n_11683, n16969);
  and g25726 (n16970, n_11682, n_11683);
  not g25727 (n_11684, n16970);
  and g25728 (n16971, n_3119, n_11684);
  and g25729 (n16972, pi0681, n_11549);
  and g25730 (n16973, pi0680, n_11543);
  and g25731 (n16974, n_11502, n_11445);
  and g25732 (n16975, pi0616, n16657);
  not g25733 (n_11685, n16974);
  and g25734 (n16976, n_11685, n16975);
  not g25735 (n_11686, n16973);
  and g25736 (n16977, n_11686, n16976);
  and g25737 (n16978, pi0616, n16653);
  and g25738 (n16979, n_11455, n16978);
  not g25739 (n_11687, n16977);
  not g25740 (n_11688, n16979);
  and g25741 (n16980, n_11687, n_11688);
  and g25742 (n16981, n_3091, n_11455);
  and g25743 (n16982, n16801, n16981);
  and g25744 (n16983, n_11502, n16802);
  and g25745 (n16984, n_3091, n16657);
  and g25746 (n16985, n_11686, n16984);
  not g25747 (n_11689, n16983);
  and g25748 (n16986, n_11689, n16985);
  not g25749 (n_11690, n16982);
  not g25750 (n_11691, n16986);
  and g25751 (n16987, n_11690, n_11691);
  and g25752 (n16988, n_3098, n16980);
  and g25753 (n16989, n16987, n16988);
  not g25754 (n_11692, n16972);
  not g25755 (n_11693, n16989);
  and g25756 (n16990, n_11692, n_11693);
  not g25757 (n_11694, n16990);
  and g25758 (n16991, n6205, n_11694);
  not g25759 (n_11695, n16971);
  not g25760 (n_11696, n16991);
  and g25761 (n16992, n_11695, n_11696);
  not g25762 (n_11697, n16992);
  and g25763 (n16993, pi0223, n_11697);
  and g25764 (n16994, pi0681, n_11526);
  and g25765 (n16995, pi0680, n_11513);
  and g25766 (n16996, pi0614, n16657);
  and g25767 (n16997, n_11685, n16996);
  not g25768 (n_11698, n16995);
  and g25769 (n16998, n_11698, n16997);
  and g25770 (n16999, pi0614, n16653);
  and g25771 (n17000, n_11455, n16999);
  not g25772 (n_11699, n16998);
  not g25773 (n_11700, n17000);
  and g25774 (n17001, n_11699, n_11700);
  and g25775 (n17002, n_3090, n_3139);
  and g25776 (n17003, n_3091, n_11520);
  and g25777 (n17004, n_11524, n17002);
  not g25778 (n_11701, n17003);
  and g25779 (n17005, n_11701, n17004);
  and g25780 (n17006, n_3090, n6195);
  and g25781 (n17007, n16684, n17006);
  not g25782 (n_11702, n17005);
  not g25783 (n_11703, n17007);
  and g25784 (n17008, n_11702, n_11703);
  and g25785 (n17009, n_3098, n17001);
  and g25786 (n17010, n17008, n17009);
  not g25787 (n_11704, n16994);
  not g25788 (n_11705, n17010);
  and g25789 (n17011, n_11704, n_11705);
  not g25790 (n_11706, n17011);
  and g25791 (n17012, n6205, n_11706);
  and g25792 (n17013, pi0681, n_11503);
  and g25793 (n17014, n6194, n_11448);
  not g25794 (n_11707, n6194);
  and g25795 (n17015, n_11707, n16702);
  not g25796 (n_11708, n17014);
  and g25797 (n17016, n_3098, n_11708);
  not g25798 (n_11709, n17015);
  and g25799 (n17017, n_11709, n17016);
  not g25800 (n_11710, n17013);
  not g25801 (n_11711, n17017);
  and g25802 (n17018, n_11710, n_11711);
  not g25803 (n_11712, n17018);
  and g25804 (n17019, n_3119, n_11712);
  not g25805 (n_11713, n17012);
  not g25806 (n_11714, n17019);
  and g25807 (n17020, n_11713, n_11714);
  and g25808 (n17021, n_9349, n17020);
  not g25809 (n_11715, n16654);
  and g25810 (n17022, n_223, n_11715);
  not g25811 (n_11716, n17021);
  and g25812 (n17023, n_11716, n17022);
  not g25813 (n_11717, n16993);
  not g25814 (n_11718, n17023);
  and g25815 (n17024, n_11717, n_11718);
  not g25816 (n_11719, n17024);
  and g25817 (n17025, n_234, n_11719);
  and g25818 (n17026, n3448, n16653);
  and g25819 (n17027, n6241, n_11706);
  not g25820 (n_11720, n6241);
  and g25821 (n17028, n_11720, n_11712);
  not g25822 (n_11721, n17028);
  and g25823 (n17029, n6236, n_11721);
  not g25824 (n_11722, n17027);
  and g25825 (n17030, n_11722, n17029);
  and g25826 (n17031, n_9350, n17030);
  not g25827 (n_11723, n6236);
  and g25828 (n17032, n_11723, n17018);
  and g25829 (n17033, n_9350, n17032);
  not g25832 (n_11725, n17033);
  not g25834 (n_11726, n17031);
  and g25836 (n17037, n_11723, n16970);
  and g25837 (n17038, n_11720, n_11684);
  and g25838 (n17039, n6241, n_11694);
  not g25839 (n_11727, n17039);
  and g25840 (n17040, n6236, n_11727);
  not g25841 (n_11728, n17038);
  and g25842 (n17041, n_11728, n17040);
  not g25843 (n_11729, n17037);
  not g25844 (n_11730, n17041);
  and g25845 (n17042, n_11729, n_11730);
  and g25846 (n17043, pi0215, n17042);
  not g25847 (n_11731, n17036);
  not g25848 (n_11732, n17043);
  and g25849 (n17044, n_11731, n_11732);
  not g25850 (n_11733, n17044);
  and g25851 (n17045, pi0299, n_11733);
  not g25852 (n_11734, n17025);
  not g25853 (n_11735, n17045);
  and g25854 (n17046, n_11734, n_11735);
  not g25855 (n_11736, n17046);
  and g25856 (n17047, pi0039, n_11736);
  not g25857 (n_11737, n16959);
  not g25858 (n_11738, n17047);
  and g25859 (n17048, n_11737, n_11738);
  not g25860 (n_11739, n17048);
  and g25861 (n17049, n_161, n_11739);
  and g25862 (n17050, n2926, n6135);
  not g25863 (n_11740, n17050);
  and g25864 (n17051, pi0038, n_11740);
  not g25865 (n_11741, n17049);
  not g25866 (n_11742, n17051);
  and g25867 (n17052, n_11741, n_11742);
  and g25868 (n17053, n_6245, pi0738);
  not g25869 (n_11743, n17052);
  and g25870 (n17054, n_11743, n17053);
  not g25871 (n_11744, n17054);
  and g25872 (n17055, n2571, n_11744);
  not g25873 (n_11745, n16955);
  and g25874 (n17056, n_11745, n17055);
  not g25875 (n_11746, n16640);
  not g25876 (n_11747, n17056);
  and g25877 (n17057, n_11746, n_11747);
  not g25878 (n_11749, pi0778);
  not g25879 (n_11750, n17057);
  and g25880 (n17058, n_11749, n_11750);
  and g25881 (n17059, n2571, n17052);
  not g25882 (n_11751, n17059);
  and g25883 (n17060, n_6245, n_11751);
  not g25884 (n_11753, pi0625);
  and g25885 (n17061, n_11753, n17060);
  and g25886 (n17062, pi0625, n17057);
  not g25887 (n_11755, n17061);
  and g25888 (n17063, pi1153, n_11755);
  not g25889 (n_11756, n17062);
  and g25890 (n17064, n_11756, n17063);
  and g25891 (n17065, n_11753, n17057);
  and g25892 (n17066, pi0625, n17060);
  not g25893 (n_11757, pi1153);
  not g25894 (n_11758, n17066);
  and g25895 (n17067, n_11757, n_11758);
  not g25896 (n_11759, n17065);
  and g25897 (n17068, n_11759, n17067);
  not g25898 (n_11760, n17064);
  not g25899 (n_11761, n17068);
  and g25900 (n17069, n_11760, n_11761);
  not g25901 (n_11762, n17069);
  and g25902 (n17070, pi0778, n_11762);
  not g25903 (n_11763, n17058);
  not g25904 (n_11764, n17070);
  and g25905 (n17071, n_11763, n_11764);
  and g25906 (n17072, pi0660, pi1155);
  not g25907 (n_11767, pi0660);
  not g25908 (n_11768, pi1155);
  and g25909 (n17073, n_11767, n_11768);
  not g25910 (n_11770, n17072);
  and g25911 (n17074, pi0785, n_11770);
  not g25912 (n_11771, n17073);
  and g25913 (n17075, n_11771, n17074);
  not g25914 (n_11772, n17071);
  not g25915 (n_11773, n17075);
  and g25916 (n17076, n_11772, n_11773);
  not g25917 (n_11774, n17060);
  and g25918 (n17077, n_11774, n17075);
  not g25919 (n_11775, n17076);
  not g25920 (n_11776, n17077);
  and g25921 (n17078, n_11775, n_11776);
  not g25922 (n_11777, n16639);
  and g25923 (n17079, n_11777, n17078);
  and g25924 (n17080, n16639, n17060);
  not g25925 (n_11778, n17079);
  not g25926 (n_11779, n17080);
  and g25927 (n17081, n_11778, n_11779);
  not g25928 (n_11780, n16635);
  and g25929 (n17082, n_11780, n17081);
  and g25930 (n17083, n16635, n_11774);
  not g25931 (n_11781, n17082);
  not g25932 (n_11782, n17083);
  and g25933 (n17084, n_11781, n_11782);
  not g25934 (n_11783, n16631);
  and g25935 (n17085, n_11783, n17084);
  and g25936 (n17086, n16631, n17060);
  not g25937 (n_11784, n17085);
  not g25938 (n_11785, n17086);
  and g25939 (n17087, n_11784, n_11785);
  not g25940 (n_11787, pi0792);
  and g25941 (n17088, n_11787, n17087);
  not g25942 (n_11789, pi0628);
  and g25943 (n17089, n_11789, n17060);
  not g25944 (n_11790, n17087);
  and g25945 (n17090, pi0628, n_11790);
  not g25946 (n_11792, n17089);
  and g25947 (n17091, pi1156, n_11792);
  not g25948 (n_11793, n17090);
  and g25949 (n17092, n_11793, n17091);
  and g25950 (n17093, pi0628, n17060);
  and g25951 (n17094, n_11789, n_11790);
  not g25952 (n_11794, pi1156);
  not g25953 (n_11795, n17093);
  and g25954 (n17095, n_11794, n_11795);
  not g25955 (n_11796, n17094);
  and g25956 (n17096, n_11796, n17095);
  not g25957 (n_11797, n17092);
  not g25958 (n_11798, n17096);
  and g25959 (n17097, n_11797, n_11798);
  not g25960 (n_11799, n17097);
  and g25961 (n17098, pi0792, n_11799);
  not g25962 (n_11800, n17088);
  not g25963 (n_11801, n17098);
  and g25964 (n17099, n_11800, n_11801);
  not g25965 (n_11803, pi0787);
  not g25966 (n_11804, n17099);
  and g25967 (n17100, n_11803, n_11804);
  not g25968 (n_11806, pi0647);
  and g25969 (n17101, n_11806, n17060);
  and g25970 (n17102, pi0647, n17099);
  not g25971 (n_11808, n17101);
  and g25972 (n17103, pi1157, n_11808);
  not g25973 (n_11809, n17102);
  and g25974 (n17104, n_11809, n17103);
  and g25975 (n17105, n_11806, n17099);
  and g25976 (n17106, pi0647, n17060);
  not g25977 (n_11810, pi1157);
  not g25978 (n_11811, n17106);
  and g25979 (n17107, n_11810, n_11811);
  not g25980 (n_11812, n17105);
  and g25981 (n17108, n_11812, n17107);
  not g25982 (n_11813, n17104);
  not g25983 (n_11814, n17108);
  and g25984 (n17109, n_11813, n_11814);
  not g25985 (n_11815, n17109);
  and g25986 (n17110, pi0787, n_11815);
  not g25987 (n_11816, n17100);
  not g25988 (n_11817, n17110);
  and g25989 (n17111, n_11816, n_11817);
  not g25990 (n_11819, pi0644);
  and g25991 (n17112, n_11819, n17111);
  not g25992 (n_11821, pi0619);
  and g25993 (n17113, n_11821, n17060);
  not g25994 (n_11823, pi0608);
  and g25995 (n17114, n_11823, pi1153);
  and g25996 (n17115, pi0608, n_11757);
  not g25997 (n_11824, n17114);
  not g25998 (n_11825, n17115);
  and g25999 (n17116, n_11824, n_11825);
  not g26000 (n_11826, n17116);
  and g26001 (n17117, pi0778, n_11826);
  and g26002 (n17118, pi0621, n16891);
  not g26003 (n_11828, n17118);
  and g26004 (n17119, n_271, n_11828);
  and g26005 (n17120, pi0621, n16913);
  not g26006 (n_11829, n17120);
  and g26007 (n17121, pi0210, n_11829);
  not g26008 (n_11830, n17119);
  not g26009 (n_11831, n17121);
  and g26010 (n17122, n_11830, n_11831);
  not g26011 (n_11832, n17122);
  and g26012 (n17123, pi0603, n_11832);
  not g26013 (n_11833, n17123);
  and g26014 (n17124, n16941, n_11833);
  not g26015 (n_11834, n17124);
  and g26016 (n17125, pi0299, n_11834);
  and g26017 (n17126, n_305, n_11828);
  and g26018 (n17127, pi0198, n_11829);
  not g26019 (n_11835, n17126);
  not g26020 (n_11836, n17127);
  and g26021 (n17128, n_11835, n_11836);
  and g26022 (n17129, pi0621, n_11613);
  not g26023 (n_11837, n17129);
  and g26024 (n17130, n_11614, n_11837);
  and g26025 (n17131, n_305, n17130);
  and g26026 (n17132, pi0621, n_11629);
  not g26027 (n_11838, n17132);
  and g26028 (n17133, n_11631, n_11838);
  and g26029 (n17134, pi0198, n17133);
  not g26030 (n_11839, n17131);
  not g26031 (n_11840, n17134);
  and g26032 (n17135, n_11839, n_11840);
  not g26033 (n_11841, n17135);
  and g26034 (n17136, n_11512, n_11841);
  not g26035 (n_11842, n17128);
  not g26036 (n_11843, n17136);
  and g26037 (n17137, n_11842, n_11843);
  and g26038 (n17138, n_234, n17137);
  not g26039 (n_11844, n17125);
  not g26040 (n_11845, n17138);
  and g26041 (n17139, n_11844, n_11845);
  not g26042 (n_11846, n17139);
  and g26043 (n17140, n_162, n_11846);
  and g26044 (n17141, n_3139, n_11503);
  and g26045 (n17142, n6195, n16681);
  not g26046 (n_11847, n17141);
  not g26047 (n_11848, n17142);
  and g26048 (n17143, n_11847, n_11848);
  and g26049 (n17144, pi0621, pi1091);
  and g26050 (n17145, n16680, n17144);
  and g26051 (n17146, pi0621, n_11443);
  not g26052 (n_11849, n17146);
  and g26053 (n17147, n_11448, n_11849);
  and g26054 (n17148, n_11512, n17147);
  and g26055 (n17149, n_11512, n16699);
  and g26056 (n17150, n6197, n17145);
  and g26057 (n17151, n16698, n17144);
  not g26058 (n_11850, n17151);
  and g26059 (n17152, pi0603, n_11850);
  not g26060 (n_11851, n17150);
  and g26061 (n17153, n_11851, n17152);
  not g26062 (n_11852, n17149);
  not g26063 (n_11853, n17153);
  and g26064 (n17154, n_11852, n_11853);
  not g26065 (n_11854, n17145);
  not g26066 (n_11855, n17148);
  and g26067 (n17155, n_11854, n_11855);
  not g26068 (n_11856, n17154);
  and g26069 (n17156, n_11856, n17155);
  not g26070 (n_11857, n17156);
  and g26071 (n17157, n17143, n_11857);
  not g26072 (n_11858, n17157);
  and g26073 (n17158, n_3162, n_11858);
  and g26074 (n17159, n16653, n17144);
  not g26075 (n_11859, n17159);
  and g26076 (n17160, n6197, n_11859);
  and g26077 (n17161, n_3102, n_11854);
  not g26078 (n_11860, n17160);
  not g26079 (n_11861, n17161);
  and g26080 (n17162, n_11860, n_11861);
  not g26081 (n_11862, n17162);
  and g26082 (n17163, pi0603, n_11862);
  not g26083 (n_11863, n17163);
  and g26084 (n17164, n16684, n_11863);
  not g26085 (n_11864, n17164);
  and g26086 (n17165, n6195, n_11864);
  and g26087 (n17166, n_3090, n_3087);
  and g26088 (n17167, n_3091, n17166);
  not g26089 (n_11865, n17144);
  and g26090 (n17168, pi0603, n_11865);
  not g26091 (n_11866, n17168);
  and g26092 (n17169, n16653, n_11866);
  not g26093 (n_11867, n17167);
  and g26094 (n17170, n_11867, n17169);
  and g26095 (n17171, n_11514, n17167);
  and g26096 (n17172, n_11863, n17171);
  not g26097 (n_11868, n17170);
  not g26098 (n_11869, n17172);
  and g26099 (n17173, n_11868, n_11869);
  and g26100 (n17174, n_3139, n17173);
  not g26101 (n_11870, n17165);
  not g26102 (n_11871, n17174);
  and g26103 (n17175, n_11870, n_11871);
  not g26104 (n_11872, n17175);
  and g26105 (n17176, n6242, n_11872);
  not g26106 (n_11873, n17158);
  and g26107 (n17177, n_9350, n_11873);
  not g26108 (n_11874, n17176);
  and g26109 (n17178, n_11874, n17177);
  and g26110 (n17179, n3448, n17169);
  not g26111 (n_11875, n17178);
  not g26112 (n_11876, n17179);
  and g26113 (n17180, n_11875, n_11876);
  not g26114 (n_11877, n17180);
  and g26115 (n17181, n_36, n_11877);
  and g26116 (n17182, n2926, n_11866);
  and g26117 (n17183, n_11556, n17182);
  and g26118 (n17184, n6192, n_11477);
  not g26119 (n_11878, n17184);
  and g26120 (n17185, n17183, n_11878);
  not g26121 (n_11879, n17185);
  and g26122 (n17186, n_3139, n_11879);
  and g26123 (n17187, n_11479, n17182);
  not g26124 (n_11880, n17187);
  and g26125 (n17188, n6195, n_11880);
  not g26126 (n_11881, n17186);
  not g26127 (n_11882, n17188);
  and g26128 (n17189, n_11881, n_11882);
  not g26129 (n_11883, n17189);
  and g26130 (n17190, n_3162, n_11883);
  and g26131 (n17191, pi0621, n16716);
  not g26132 (n_11884, n17191);
  and g26133 (n17192, n_3102, n_11884);
  not g26134 (n_11885, n17192);
  and g26135 (n17193, n_11860, n_11885);
  not g26136 (n_11886, n17193);
  and g26137 (n17194, pi0603, n_11886);
  not g26138 (n_11887, n17194);
  and g26139 (n17195, n17171, n_11887);
  not g26140 (n_11888, n17195);
  and g26141 (n17196, n_11868, n_11888);
  not g26142 (n_11889, n17196);
  and g26143 (n17197, n_3139, n_11889);
  and g26144 (n17198, n6195, n16797);
  and g26145 (n17199, n_11887, n17198);
  not g26146 (n_11890, n17197);
  not g26147 (n_11891, n17199);
  and g26148 (n17200, n_11890, n_11891);
  and g26149 (n17201, n6242, n17200);
  not g26150 (n_11892, n17190);
  and g26151 (n17202, pi0215, n_11892);
  not g26152 (n_11893, n17201);
  and g26153 (n17203, n_11893, n17202);
  not g26154 (n_11894, n17181);
  not g26155 (n_11895, n17203);
  and g26156 (n17204, n_11894, n_11895);
  not g26157 (n_11896, n17204);
  and g26158 (n17205, pi0299, n_11896);
  and g26159 (n17206, n_3119, n_11858);
  and g26160 (n17207, n6205, n_11872);
  not g26161 (n_11897, n17206);
  and g26162 (n17208, n_9349, n_11897);
  not g26163 (n_11898, n17207);
  and g26164 (n17209, n_11898, n17208);
  and g26165 (n17210, n2603, n17169);
  not g26166 (n_11899, n17209);
  not g26167 (n_11900, n17210);
  and g26168 (n17211, n_11899, n_11900);
  not g26169 (n_11901, n17211);
  and g26170 (n17212, n_223, n_11901);
  and g26171 (n17213, n_3119, n_11883);
  and g26172 (n17214, n6205, n17200);
  not g26173 (n_11902, n17213);
  and g26174 (n17215, pi0223, n_11902);
  not g26175 (n_11903, n17214);
  and g26176 (n17216, n_11903, n17215);
  not g26177 (n_11904, n17212);
  not g26178 (n_11905, n17216);
  and g26179 (n17217, n_11904, n_11905);
  not g26180 (n_11906, n17217);
  and g26181 (n17218, n_234, n_11906);
  not g26182 (n_11907, n17205);
  not g26183 (n_11908, n17218);
  and g26184 (n17219, n_11907, n_11908);
  and g26185 (n17220, pi0039, n17219);
  not g26186 (n_11909, n17140);
  not g26187 (n_11910, n17220);
  and g26188 (n17221, n_11909, n_11910);
  not g26189 (n_11912, pi0761);
  and g26190 (n17222, n_11912, n17221);
  and g26191 (n17223, pi0761, n17048);
  not g26192 (n_11913, n17222);
  and g26193 (n17224, n_6245, n_11913);
  not g26194 (n_11914, n17223);
  and g26195 (n17225, n_11914, n17224);
  and g26196 (n17226, pi0603, n_11841);
  not g26197 (n_11915, n17226);
  and g26198 (n17227, n_234, n_11915);
  not g26199 (n_11916, n17130);
  and g26200 (n17228, n_271, n_11916);
  not g26201 (n_11917, n17133);
  and g26202 (n17229, pi0210, n_11917);
  not g26203 (n_11918, n17228);
  not g26204 (n_11919, n17229);
  and g26205 (n17230, n_11918, n_11919);
  and g26206 (n17231, pi0603, n17230);
  not g26207 (n_11920, n17231);
  and g26208 (n17232, pi0299, n_11920);
  not g26209 (n_11921, n17227);
  not g26210 (n_11922, n17232);
  and g26211 (n17233, n_11921, n_11922);
  not g26212 (n_11923, n17233);
  and g26213 (n17234, n_162, n_11923);
  and g26214 (n17235, n16653, n17168);
  and g26215 (n17236, n_11481, n17235);
  and g26216 (n17237, n_11556, n17235);
  and g26217 (n17238, n16725, n17167);
  not g26218 (n_11924, n17238);
  and g26219 (n17239, n17237, n_11924);
  and g26220 (n17240, n_3139, n17239);
  not g26221 (n_11925, n17236);
  not g26222 (n_11926, n17240);
  and g26223 (n17241, n_11925, n_11926);
  not g26224 (n_11927, n17241);
  and g26225 (n17242, n_11494, n_11927);
  not g26226 (n_11928, n17242);
  and g26227 (n17243, pi0215, n_11928);
  and g26228 (n17244, n2926, n17168);
  and g26229 (n17245, n16825, n17244);
  and g26230 (n17246, n16684, n17168);
  and g26231 (n17247, n6195, n17246);
  and g26232 (n17248, n_11867, n17235);
  and g26233 (n17249, n17167, n17246);
  not g26234 (n_11929, n17248);
  not g26235 (n_11930, n17249);
  and g26236 (n17250, n_11929, n_11930);
  not g26237 (n_11931, n17250);
  and g26238 (n17251, n_3139, n_11931);
  not g26239 (n_11932, n17247);
  not g26240 (n_11933, n17251);
  and g26241 (n17252, n_11932, n_11933);
  and g26242 (n17253, n6242, n17252);
  and g26243 (n17254, n17143, n17168);
  not g26244 (n_11934, n17254);
  and g26245 (n17255, n_3162, n_11934);
  not g26246 (n_11935, n17253);
  and g26247 (n17256, n_9350, n_11935);
  not g26248 (n_11936, n17255);
  and g26249 (n17257, n_11936, n17256);
  not g26250 (n_11937, n17245);
  and g26251 (n17258, n_36, n_11937);
  not g26252 (n_11938, n17257);
  and g26253 (n17259, n_11938, n17258);
  not g26254 (n_11939, n17243);
  and g26255 (n17260, pi0299, n_11939);
  not g26256 (n_11940, n17259);
  and g26257 (n17261, n_11940, n17260);
  and g26258 (n17262, n_11484, n_11927);
  not g26259 (n_11941, n17262);
  and g26260 (n17263, pi0223, n_11941);
  and g26261 (n17264, n6205, n17252);
  and g26262 (n17265, n_3119, n_11934);
  not g26263 (n_11942, n17264);
  and g26264 (n17266, n_9349, n_11942);
  not g26265 (n_11943, n17265);
  and g26266 (n17267, n_11943, n17266);
  and g26267 (n17268, n16654, n17168);
  not g26268 (n_11944, n17268);
  and g26269 (n17269, n_223, n_11944);
  not g26270 (n_11945, n17267);
  and g26271 (n17270, n_11945, n17269);
  not g26272 (n_11946, n17263);
  and g26273 (n17271, n_234, n_11946);
  not g26274 (n_11947, n17270);
  and g26275 (n17272, n_11947, n17271);
  not g26276 (n_11948, n17261);
  not g26277 (n_11949, n17272);
  and g26278 (n17273, n_11948, n_11949);
  and g26279 (n17274, pi0039, n17273);
  not g26280 (n_11950, n17234);
  not g26281 (n_11951, n17274);
  and g26282 (n17275, n_11950, n_11951);
  and g26283 (n17276, pi0140, n_11912);
  and g26284 (n17277, n17275, n17276);
  not g26285 (n_11952, n17225);
  not g26286 (n_11953, n17277);
  and g26287 (n17278, n_11952, n_11953);
  not g26288 (n_11954, n17278);
  and g26289 (n17279, n_161, n_11954);
  and g26290 (n17280, n6284, n17244);
  and g26291 (n17281, n_11912, n17280);
  not g26292 (n_11955, n17281);
  and g26293 (n17282, n_11422, n_11955);
  not g26294 (n_11956, n17282);
  and g26295 (n17283, pi0038, n_11956);
  not g26296 (n_11957, n17279);
  not g26297 (n_11958, n17283);
  and g26298 (n17284, n_11957, n_11958);
  and g26299 (n17285, n2571, n17284);
  not g26300 (n_11959, n17285);
  and g26301 (n17286, n_11746, n_11959);
  not g26302 (n_11960, n17117);
  not g26303 (n_11961, n17286);
  and g26304 (n17287, n_11960, n_11961);
  and g26305 (n17288, n_11774, n17117);
  not g26306 (n_11962, n17287);
  not g26307 (n_11963, n17288);
  and g26308 (n17289, n_11962, n_11963);
  not g26309 (n_11964, pi0785);
  not g26310 (n_11965, n17289);
  and g26311 (n17290, n_11964, n_11965);
  and g26312 (n17291, pi0609, n_11960);
  not g26313 (n_11967, n17291);
  and g26314 (n17292, n_11774, n_11967);
  and g26315 (n17293, pi0609, n17287);
  not g26316 (n_11968, n17292);
  not g26317 (n_11969, n17293);
  and g26318 (n17294, n_11968, n_11969);
  not g26319 (n_11970, n17294);
  and g26320 (n17295, pi1155, n_11970);
  not g26321 (n_11971, pi0609);
  and g26322 (n17296, n_11971, n_11960);
  not g26323 (n_11972, n17296);
  and g26324 (n17297, n_11774, n_11972);
  and g26325 (n17298, n_11971, n17287);
  not g26326 (n_11973, n17297);
  not g26327 (n_11974, n17298);
  and g26328 (n17299, n_11973, n_11974);
  not g26329 (n_11975, n17299);
  and g26330 (n17300, n_11768, n_11975);
  not g26331 (n_11976, n17295);
  not g26332 (n_11977, n17300);
  and g26333 (n17301, n_11976, n_11977);
  not g26334 (n_11978, n17301);
  and g26335 (n17302, pi0785, n_11978);
  not g26336 (n_11979, n17290);
  not g26337 (n_11980, n17302);
  and g26338 (n17303, n_11979, n_11980);
  not g26339 (n_11981, pi0781);
  not g26340 (n_11982, n17303);
  and g26341 (n17304, n_11981, n_11982);
  not g26342 (n_11984, pi0618);
  and g26343 (n17305, n_11984, n17060);
  and g26344 (n17306, pi0618, n17303);
  not g26345 (n_11985, n17305);
  and g26346 (n17307, pi1154, n_11985);
  not g26347 (n_11986, n17306);
  and g26348 (n17308, n_11986, n17307);
  and g26349 (n17309, n_11984, n17303);
  and g26350 (n17310, pi0618, n17060);
  not g26351 (n_11987, n17310);
  and g26352 (n17311, n_11413, n_11987);
  not g26353 (n_11988, n17309);
  and g26354 (n17312, n_11988, n17311);
  not g26355 (n_11989, n17308);
  not g26356 (n_11990, n17312);
  and g26357 (n17313, n_11989, n_11990);
  not g26358 (n_11991, n17313);
  and g26359 (n17314, pi0781, n_11991);
  not g26360 (n_11992, n17304);
  not g26361 (n_11993, n17314);
  and g26362 (n17315, n_11992, n_11993);
  and g26363 (n17316, pi0619, n17315);
  not g26364 (n_11994, n17113);
  and g26365 (n17317, pi1159, n_11994);
  not g26366 (n_11995, n17316);
  and g26367 (n17318, n_11995, n17317);
  not g26368 (n_11996, n17284);
  and g26369 (n17319, pi0738, n_11996);
  and g26370 (n17320, n_11479, n17235);
  not g26371 (n_11997, n17320);
  and g26372 (n17321, n_11550, n_11997);
  and g26373 (n17322, n6195, n17321);
  and g26374 (n17323, pi0680, n_11455);
  not g26375 (n_11998, n16756);
  and g26376 (n17324, n_11998, n_11550);
  not g26377 (n_11999, n17237);
  and g26378 (n17325, n_11999, n17324);
  and g26379 (n17326, n_11867, n17325);
  and g26380 (n17327, n_11512, n16756);
  not g26381 (n_12000, n17327);
  and g26382 (n17328, n17321, n_12000);
  and g26383 (n17329, n17167, n17328);
  not g26384 (n_12001, n17326);
  not g26385 (n_12002, n17329);
  and g26386 (n17330, n_12001, n_12002);
  not g26387 (n_12003, n17330);
  and g26388 (n17331, n17323, n_12003);
  not g26389 (n_12004, n17322);
  not g26390 (n_12005, n17331);
  and g26391 (n17332, n_12004, n_12005);
  and g26392 (n17333, n_11559, n17332);
  not g26393 (n_12006, n17333);
  and g26394 (n17334, n_3119, n_12006);
  and g26395 (n17335, n16808, n_11925);
  and g26396 (n17336, n_11420, n_11866);
  not g26397 (n_12007, n17336);
  and g26398 (n17337, n16653, n_12007);
  not g26399 (n_12008, n17337);
  and g26400 (n17338, pi0616, n_12008);
  and g26401 (n17339, pi0614, n_12008);
  and g26402 (n17340, pi0642, n_12008);
  not g26406 (n_12009, n17340);
  not g26407 (n_12010, n17343);
  and g26408 (n17344, n_12009, n_12010);
  not g26409 (n_12011, n17344);
  and g26410 (n17345, n_3090, n_12011);
  not g26411 (n_12012, n17339);
  not g26412 (n_12013, n17345);
  and g26413 (n17346, n_12012, n_12013);
  not g26414 (n_12014, n17346);
  and g26415 (n17347, n_3091, n_12014);
  not g26416 (n_12015, n17338);
  not g26417 (n_12016, n17347);
  and g26418 (n17348, n_12015, n_12016);
  not g26419 (n_12017, n17348);
  and g26420 (n17349, n17323, n_12017);
  not g26421 (n_12018, n17335);
  and g26422 (n17350, n_11555, n_12018);
  not g26423 (n_12019, n17349);
  and g26424 (n17351, n_12019, n17350);
  not g26425 (n_12020, n17351);
  and g26426 (n17352, n6205, n_12020);
  not g26427 (n_12021, n17334);
  and g26428 (n17353, pi0223, n_12021);
  not g26429 (n_12022, n17352);
  and g26430 (n17354, n_12022, n17353);
  and g26431 (n17355, pi0680, n17336);
  not g26432 (n_12023, n17355);
  and g26433 (n17356, n16653, n_12023);
  not g26434 (n_12024, n17356);
  and g26435 (n17357, n2603, n_12024);
  and g26436 (n17358, n16769, n_12007);
  not g26437 (n_12025, n17358);
  and g26438 (n17359, n_3087, n_12025);
  not g26439 (n_12026, n17359);
  and g26440 (n17360, n_12009, n_12026);
  not g26441 (n_12027, n17360);
  and g26442 (n17361, n_3090, n_12027);
  not g26443 (n_12028, n17361);
  and g26444 (n17362, n_12012, n_12028);
  not g26445 (n_12029, n17362);
  and g26446 (n17363, n_3091, n_12029);
  not g26447 (n_12030, n17363);
  and g26448 (n17364, n_12015, n_12030);
  not g26449 (n_12031, n17364);
  and g26450 (n17365, n17323, n_12031);
  and g26451 (n17366, n_11512, n_11535);
  not g26452 (n_12032, pi0665);
  and g26453 (n17367, pi0603, n_12032);
  and g26454 (n17368, n17144, n17367);
  not g26455 (n_12033, n17368);
  and g26456 (n17369, n_11515, n_12033);
  not g26457 (n_12034, n17366);
  and g26458 (n17370, n_12034, n17369);
  not g26459 (n_12035, n17370);
  and g26460 (n17371, n6195, n_12035);
  not g26461 (n_12036, n17371);
  and g26462 (n17372, n_11533, n_12036);
  not g26463 (n_12037, n17365);
  and g26464 (n17373, n_12037, n17372);
  and g26465 (n17374, n6205, n17373);
  and g26466 (n17375, pi0603, n17147);
  not g26467 (n_12038, pi0621);
  and g26468 (n17376, pi0603, n_12038);
  not g26469 (n_12039, n17376);
  and g26470 (n17377, n16754, n_12039);
  not g26471 (n_12040, n17377);
  and g26472 (n17378, n6195, n_12040);
  not g26473 (n_12041, n17375);
  and g26474 (n17379, n_12041, n17378);
  and g26475 (n17380, n16702, n_12007);
  not g26476 (n_12042, n17380);
  and g26477 (n17381, n17323, n_12042);
  not g26478 (n_12043, n17379);
  and g26479 (n17382, n_11509, n_12043);
  not g26480 (n_12044, n17381);
  and g26481 (n17383, n_12044, n17382);
  and g26482 (n17384, n_3119, n17383);
  not g26483 (n_12045, n17384);
  and g26484 (n17385, n_9349, n_12045);
  not g26485 (n_12046, n17374);
  and g26486 (n17386, n_12046, n17385);
  not g26487 (n_12047, n17357);
  and g26488 (n17387, n_223, n_12047);
  not g26489 (n_12048, n17386);
  and g26490 (n17388, n_12048, n17387);
  not g26491 (n_12049, n17354);
  not g26492 (n_12050, n17388);
  and g26493 (n17389, n_12049, n_12050);
  not g26494 (n_12051, n17389);
  and g26495 (n17390, n_234, n_12051);
  and g26496 (n17391, n3448, n_12024);
  not g26497 (n_12052, n17383);
  and g26498 (n17392, n_3162, n_12052);
  not g26499 (n_12053, n17373);
  and g26500 (n17393, n6242, n_12053);
  not g26501 (n_12054, n17392);
  not g26502 (n_12055, n17393);
  and g26503 (n17394, n_12054, n_12055);
  not g26504 (n_12056, n17394);
  and g26505 (n17395, n_9350, n_12056);
  not g26506 (n_12057, n17391);
  and g26507 (n17396, n_36, n_12057);
  not g26508 (n_12058, n17395);
  and g26509 (n17397, n_12058, n17396);
  and g26510 (n17398, n6242, n_12020);
  and g26511 (n17399, n_3162, n_12006);
  not g26512 (n_12059, n17399);
  and g26513 (n17400, pi0215, n_12059);
  not g26514 (n_12060, n17398);
  and g26515 (n17401, n_12060, n17400);
  not g26516 (n_12061, n17397);
  not g26517 (n_12062, n17401);
  and g26518 (n17402, n_12061, n_12062);
  not g26519 (n_12063, n17402);
  and g26520 (n17403, pi0299, n_12063);
  not g26521 (n_12064, n17390);
  not g26522 (n_12065, n17403);
  and g26523 (n17404, n_12064, n_12065);
  and g26524 (n17405, n_6245, n17404);
  and g26525 (n17406, n17026, n17355);
  and g26526 (n17407, n_11420, n17169);
  not g26527 (n_12066, n17407);
  and g26528 (n17408, pi0616, n_12066);
  not g26529 (n_12067, n17408);
  and g26530 (n17409, n17323, n_12067);
  not g26531 (n_12068, n17166);
  and g26532 (n17410, n_12068, n17407);
  and g26533 (n17411, pi0603, pi0665);
  and g26534 (n17412, n_11512, n_11450);
  not g26535 (n_12069, n17411);
  not g26536 (n_12070, n17412);
  and g26537 (n17413, n_12069, n_12070);
  and g26538 (n17414, n_11863, n17413);
  and g26539 (n17415, n17166, n17414);
  not g26540 (n_12071, n17410);
  and g26541 (n17416, n_3091, n_12071);
  not g26542 (n_12072, n17415);
  and g26543 (n17417, n_12072, n17416);
  not g26544 (n_12073, n17417);
  and g26545 (n17418, n17409, n_12073);
  and g26546 (n17419, n16684, n17371);
  not g26547 (n_12074, n17418);
  not g26548 (n_12075, n17419);
  and g26549 (n17420, n_12074, n_12075);
  and g26550 (n17421, n6242, n17420);
  and g26551 (n17422, n_11452, n17154);
  not g26552 (n_12076, n17422);
  and g26553 (n17423, pi0616, n_12076);
  and g26554 (n17424, n_12032, n17145);
  not g26555 (n_12077, n17424);
  and g26556 (n17425, pi0603, n_12077);
  not g26557 (n_12078, n16699);
  and g26558 (n17426, n_11452, n_12078);
  not g26559 (n_12079, n17426);
  and g26560 (n17427, n_11512, n_12079);
  not g26561 (n_12080, n17425);
  not g26562 (n_12081, n17427);
  and g26563 (n17428, n_12080, n_12081);
  and g26564 (n17429, n17166, n17428);
  not g26565 (n_12082, n17428);
  and g26566 (n17430, n17167, n_12082);
  not g26567 (n_12083, n17430);
  and g26568 (n17431, n17422, n_12083);
  not g26569 (n_12084, n17429);
  and g26570 (n17432, n_3091, n_12084);
  not g26571 (n_12085, n17431);
  and g26572 (n17433, n_12085, n17432);
  not g26573 (n_12086, n17423);
  not g26574 (n_12087, n17433);
  and g26575 (n17434, n_12086, n_12087);
  not g26576 (n_12088, n17434);
  and g26577 (n17435, n_11455, n_12088);
  and g26578 (n17436, n16696, n_12080);
  not g26579 (n_12089, n17323);
  not g26580 (n_12090, n17436);
  and g26581 (n17437, n_12089, n_12090);
  not g26582 (n_12091, n17435);
  not g26583 (n_12092, n17437);
  and g26584 (n17438, n_12091, n_12092);
  not g26585 (n_12093, n17438);
  and g26586 (n17439, n_3162, n_12093);
  not g26587 (n_12094, n17421);
  and g26588 (n17440, n_9350, n_12094);
  not g26589 (n_12095, n17439);
  and g26590 (n17441, n_12095, n17440);
  not g26591 (n_12096, n17406);
  and g26592 (n17442, n_36, n_12096);
  not g26593 (n_12097, n17441);
  and g26594 (n17443, n_12097, n17442);
  and g26595 (n17444, n_11420, n_11889);
  not g26596 (n_12098, n17444);
  and g26597 (n17445, n_3091, n_12098);
  not g26598 (n_12099, n17445);
  and g26599 (n17446, n17409, n_12099);
  and g26600 (n17447, n17199, n17413);
  not g26601 (n_12100, n17446);
  not g26602 (n_12101, n17447);
  and g26603 (n17448, n_12100, n_12101);
  not g26604 (n_12102, n17448);
  and g26605 (n17449, n6242, n_12102);
  and g26606 (n17450, n17183, n17413);
  not g26607 (n_12103, n17450);
  and g26608 (n17451, pi0616, n_12103);
  and g26609 (n17452, pi0614, n_3091);
  and g26610 (n17453, n_12103, n17452);
  and g26611 (n17454, n_11887, n17413);
  not g26612 (n_12104, n17454);
  and g26613 (n17455, n_3087, n_12104);
  not g26614 (n_12105, n17455);
  and g26615 (n17456, n17450, n_12105);
  not g26616 (n_12106, n17456);
  and g26617 (n17457, n6191, n_12106);
  not g26618 (n_12107, n17453);
  not g26619 (n_12108, n17457);
  and g26620 (n17458, n_12107, n_12108);
  not g26621 (n_12109, n17451);
  and g26622 (n17459, n_12109, n17458);
  not g26623 (n_12110, n17459);
  and g26624 (n17460, n_11455, n_12110);
  and g26625 (n17461, n_11479, n17355);
  not g26626 (n_12111, n17461);
  and g26627 (n17462, n_12089, n_12111);
  not g26628 (n_12112, n17460);
  not g26629 (n_12113, n17462);
  and g26630 (n17463, n_12112, n_12113);
  and g26631 (n17464, n_3162, n17463);
  not g26632 (n_12114, n17449);
  and g26633 (n17465, pi0215, n_12114);
  not g26634 (n_12115, n17464);
  and g26635 (n17466, n_12115, n17465);
  not g26636 (n_12116, n17443);
  not g26637 (n_12117, n17466);
  and g26638 (n17467, n_12116, n_12117);
  not g26639 (n_12118, n17467);
  and g26640 (n17468, pi0299, n_12118);
  and g26641 (n17469, n16645, n_11866);
  not g26642 (n_12119, n17244);
  not g26643 (n_12120, n17469);
  and g26644 (n17470, n_12119, n_12120);
  not g26645 (n_12121, n17470);
  and g26646 (n17471, n16653, n_12121);
  not g26647 (n_12122, n17471);
  and g26648 (n17472, n2603, n_12122);
  and g26649 (n17473, n_3119, n17438);
  not g26650 (n_12123, n17420);
  and g26651 (n17474, n6205, n_12123);
  not g26652 (n_12124, n17474);
  and g26653 (n17475, n_9349, n_12124);
  not g26654 (n_12125, n17473);
  and g26655 (n17476, n_12125, n17475);
  not g26656 (n_12126, n17472);
  and g26657 (n17477, n17269, n_12126);
  not g26658 (n_12127, n17476);
  and g26659 (n17478, n_12127, n17477);
  and g26660 (n17479, n6205, n17448);
  not g26661 (n_12128, n17463);
  and g26662 (n17480, n_3119, n_12128);
  not g26663 (n_12129, n17479);
  and g26664 (n17481, pi0223, n_12129);
  not g26665 (n_12130, n17480);
  and g26666 (n17482, n_12130, n17481);
  not g26667 (n_12131, n17482);
  and g26668 (n17483, n_234, n_12131);
  not g26669 (n_12132, n17478);
  and g26670 (n17484, n_12132, n17483);
  not g26671 (n_12133, n17468);
  not g26672 (n_12134, n17484);
  and g26673 (n17485, n_12133, n_12134);
  and g26674 (n17486, pi0140, n17485);
  not g26675 (n_12135, n17486);
  and g26676 (n17487, pi0761, n_12135);
  not g26677 (n_12136, n17405);
  and g26678 (n17488, n_12136, n17487);
  and g26679 (n17489, n_11501, n_11866);
  and g26680 (n17490, n16667, n17489);
  and g26681 (n17491, n_11425, n17490);
  and g26682 (n17492, n2603, n17491);
  and g26683 (n17493, n16643, n_12039);
  and g26684 (n17494, n_11506, n17493);
  not g26685 (n_12137, n17494);
  and g26686 (n17495, n17323, n_12137);
  and g26687 (n17496, n16702, n_11866);
  not g26688 (n_12138, n17496);
  and g26689 (n17497, n_11502, n_12138);
  not g26690 (n_12139, n17378);
  not g26691 (n_12140, n17495);
  and g26692 (n17498, n_12139, n_12140);
  not g26693 (n_12141, n17497);
  and g26694 (n17499, n_12141, n17498);
  and g26695 (n17500, n_3119, n17499);
  and g26696 (n17501, n_11502, n17173);
  and g26697 (n17502, n16781, n17493);
  not g26698 (n_12142, n17502);
  and g26699 (n17503, n6195, n_12142);
  and g26700 (n17504, n16778, n_12039);
  and g26701 (n17505, n_11867, n17504);
  and g26702 (n17506, n16643, n17172);
  not g26703 (n_12143, n17505);
  and g26704 (n17507, n17323, n_12143);
  not g26705 (n_12144, n17506);
  and g26706 (n17508, n_12144, n17507);
  not g26707 (n_12145, n17501);
  not g26708 (n_12146, n17503);
  and g26709 (n17509, n_12145, n_12146);
  not g26710 (n_12147, n17508);
  and g26711 (n17510, n_12147, n17509);
  and g26712 (n17511, n6205, n17510);
  not g26713 (n_12148, n17500);
  not g26714 (n_12149, n17511);
  and g26715 (n17512, n_12148, n_12149);
  not g26716 (n_12150, n17512);
  and g26717 (n17513, n_9349, n_12150);
  not g26718 (n_12151, n17492);
  and g26719 (n17514, n_223, n_12151);
  not g26720 (n_12152, n17513);
  and g26721 (n17515, n_12152, n17514);
  and g26722 (n17516, n_11501, n17197);
  and g26723 (n17517, n6195, n_12039);
  and g26724 (n17518, n16807, n17517);
  not g26725 (n_12153, n17516);
  not g26726 (n_12154, n17518);
  and g26727 (n17519, n_12153, n_12154);
  not g26728 (n_12155, n17519);
  and g26729 (n17520, n6205, n_12155);
  and g26730 (n17521, n_11502, n_11879);
  not g26731 (n_12156, n16816);
  and g26732 (n17522, n_12156, n_12039);
  not g26733 (n_12157, n17522);
  and g26734 (n17523, n6195, n_12157);
  not g26735 (n_12158, n17324);
  and g26736 (n17524, n_11889, n_12158);
  not g26737 (n_12159, n17524);
  and g26738 (n17525, n17323, n_12159);
  not g26739 (n_12160, n17521);
  not g26740 (n_12161, n17523);
  and g26741 (n17526, n_12160, n_12161);
  not g26742 (n_12162, n17525);
  and g26743 (n17527, n_12162, n17526);
  and g26744 (n17528, n_3119, n17527);
  not g26745 (n_12163, n17520);
  and g26746 (n17529, pi0223, n_12163);
  not g26747 (n_12164, n17528);
  and g26748 (n17530, n_12164, n17529);
  not g26749 (n_12165, n17515);
  not g26750 (n_12166, n17530);
  and g26751 (n17531, n_12165, n_12166);
  not g26752 (n_12167, n17531);
  and g26753 (n17532, n_234, n_12167);
  and g26754 (n17533, n3448, n17491);
  and g26755 (n17534, n_3162, n17499);
  and g26756 (n17535, n6242, n17510);
  not g26757 (n_12168, n17534);
  not g26758 (n_12169, n17535);
  and g26759 (n17536, n_12168, n_12169);
  not g26760 (n_12170, n17536);
  and g26761 (n17537, n_9350, n_12170);
  not g26762 (n_12171, n17533);
  and g26763 (n17538, n_36, n_12171);
  not g26764 (n_12172, n17537);
  and g26765 (n17539, n_12172, n17538);
  and g26766 (n17540, n6242, n_12155);
  and g26767 (n17541, n_3162, n17527);
  not g26768 (n_12173, n17540);
  and g26769 (n17542, pi0215, n_12173);
  not g26770 (n_12174, n17541);
  and g26771 (n17543, n_12174, n17542);
  not g26772 (n_12175, n17539);
  not g26773 (n_12176, n17543);
  and g26774 (n17544, n_12175, n_12176);
  not g26775 (n_12177, n17544);
  and g26776 (n17545, pi0299, n_12177);
  not g26777 (n_12178, n17532);
  not g26778 (n_12179, n17545);
  and g26779 (n17546, n_12178, n_12179);
  not g26780 (n_12180, n17546);
  and g26781 (n17547, n_6245, n_12180);
  not g26782 (n_12181, n17493);
  and g26783 (n17548, n16653, n_12181);
  and g26784 (n17549, n_11867, n17548);
  not g26785 (n_12182, n17549);
  and g26786 (n17550, n17323, n_12182);
  and g26787 (n17551, n16727, n_11925);
  not g26788 (n_12183, n17551);
  and g26789 (n17552, n17167, n_12183);
  not g26790 (n_12184, n17552);
  and g26791 (n17553, n17550, n_12184);
  and g26792 (n17554, pi0680, n_11485);
  not g26793 (n_12185, n17554);
  and g26794 (n17555, n17241, n_12185);
  not g26795 (n_12186, n17553);
  not g26796 (n_12187, n17555);
  and g26797 (n17556, n_12186, n_12187);
  not g26798 (n_12188, n17556);
  and g26799 (n17557, n6205, n_12188);
  and g26800 (n17558, n_11926, n_11997);
  and g26801 (n17559, n16658, n_11556);
  and g26802 (n17560, n_11483, n17554);
  and g26803 (n17561, n17559, n17560);
  not g26804 (n_12189, n17561);
  and g26805 (n17562, n17558, n_12189);
  and g26806 (n17563, n_3119, n17562);
  not g26807 (n_12190, n17563);
  and g26808 (n17564, pi0223, n_12190);
  not g26809 (n_12191, n17557);
  and g26810 (n17565, n_12191, n17564);
  and g26811 (n17566, n_11502, n17250);
  not g26812 (n_12192, n17246);
  not g26813 (n_12193, n17414);
  and g26814 (n17567, n_12192, n_12193);
  not g26815 (n_12194, n17567);
  and g26816 (n17568, n17167, n_12194);
  not g26817 (n_12195, n17568);
  and g26818 (n17569, n17550, n_12195);
  and g26819 (n17570, n6195, n_11456);
  and g26820 (n17571, n_12192, n17570);
  not g26821 (n_12196, n17566);
  not g26822 (n_12197, n17571);
  and g26823 (n17572, n_12196, n_12197);
  not g26824 (n_12198, n17569);
  and g26825 (n17573, n_12198, n17572);
  and g26826 (n17574, n6205, n17573);
  and g26827 (n17575, n_12041, n_12082);
  not g26828 (n_12199, n17575);
  and g26829 (n17576, n17167, n_12199);
  and g26830 (n17577, n_12078, n17168);
  not g26831 (n_12200, n17577);
  and g26832 (n17578, n_12079, n_12200);
  not g26833 (n_12201, n17578);
  and g26834 (n17579, n_11867, n_12201);
  not g26835 (n_12202, n17579);
  and g26836 (n17580, n17323, n_12202);
  not g26837 (n_12203, n17576);
  and g26838 (n17581, n_12203, n17580);
  and g26839 (n17582, n_11464, n_12089);
  and g26840 (n17583, n_11934, n17582);
  not g26841 (n_12204, n17581);
  not g26842 (n_12205, n17583);
  and g26843 (n17584, n_12204, n_12205);
  and g26844 (n17585, n_3119, n17584);
  not g26845 (n_12206, n17574);
  and g26846 (n17586, n_9349, n_12206);
  not g26847 (n_12207, n17585);
  and g26848 (n17587, n_12207, n17586);
  and g26849 (n17588, n_223, n_12126);
  not g26850 (n_12208, n17587);
  and g26851 (n17589, n_12208, n17588);
  not g26852 (n_12209, n17565);
  and g26853 (n17590, n_234, n_12209);
  not g26854 (n_12210, n17589);
  and g26855 (n17591, n_12210, n17590);
  and g26856 (n17592, n3448, n17471);
  and g26857 (n17593, n_3162, n17584);
  and g26858 (n17594, n6242, n17573);
  not g26859 (n_12211, n17593);
  not g26860 (n_12212, n17594);
  and g26861 (n17595, n_12211, n_12212);
  not g26862 (n_12213, n17595);
  and g26863 (n17596, n_9350, n_12213);
  not g26864 (n_12214, n17592);
  and g26865 (n17597, n_36, n_12214);
  not g26866 (n_12215, n17596);
  and g26867 (n17598, n_12215, n17597);
  not g26868 (n_12216, n17562);
  and g26869 (n17599, n_3162, n_12216);
  and g26870 (n17600, n6242, n17556);
  not g26871 (n_12217, n17599);
  and g26872 (n17601, pi0215, n_12217);
  not g26873 (n_12218, n17600);
  and g26874 (n17602, n_12218, n17601);
  not g26875 (n_12219, n17598);
  not g26876 (n_12220, n17602);
  and g26877 (n17603, n_12219, n_12220);
  not g26878 (n_12221, n17603);
  and g26879 (n17604, pi0299, n_12221);
  not g26880 (n_12222, n17591);
  not g26881 (n_12223, n17604);
  and g26882 (n17605, n_12222, n_12223);
  and g26883 (n17606, pi0140, n17605);
  not g26884 (n_12224, n17547);
  and g26885 (n17607, n_11912, n_12224);
  not g26886 (n_12225, n17606);
  and g26887 (n17608, n_12225, n17607);
  not g26888 (n_12226, n17488);
  not g26889 (n_12227, n17608);
  and g26890 (n17609, n_12226, n_12227);
  not g26891 (n_12228, n17609);
  and g26892 (n17610, pi0039, n_12228);
  and g26893 (n17611, pi0680, n17233);
  not g26894 (n_12229, n17611);
  and g26895 (n17612, n_11660, n_12229);
  not g26896 (n_12230, n17612);
  and g26897 (n17613, n_6245, n_12230);
  and g26898 (n17614, pi0603, n_11842);
  not g26899 (n_12231, n16918);
  and g26900 (n17615, n_11512, n_12231);
  not g26901 (n_12232, n17614);
  and g26902 (n17616, n_12069, n_12232);
  not g26903 (n_12233, n17615);
  and g26904 (n17617, n_12233, n17616);
  and g26905 (n17618, pi0680, n17617);
  not g26906 (n_12234, n17618);
  and g26907 (n17619, n_234, n_12234);
  not g26908 (n_12235, n16923);
  and g26909 (n17620, n_11512, n_12235);
  and g26910 (n17621, n_11833, n_12069);
  not g26911 (n_12236, n17620);
  and g26912 (n17622, n_12236, n17621);
  and g26913 (n17623, pi0680, n17622);
  not g26914 (n_12237, n17623);
  and g26915 (n17624, pi0299, n_12237);
  not g26916 (n_12238, n17619);
  not g26917 (n_12239, n17624);
  and g26918 (n17625, n_12238, n_12239);
  not g26919 (n_12240, n17625);
  and g26920 (n17626, pi0140, n_12240);
  not g26921 (n_12241, n17613);
  and g26922 (n17627, pi0761, n_12241);
  not g26923 (n_12242, n17626);
  and g26924 (n17628, n_12242, n17627);
  and g26925 (n17629, n16948, n17139);
  and g26926 (n17630, n_6245, n17629);
  not g26927 (n_12243, n16926);
  and g26928 (n17631, n_12243, n_11923);
  and g26929 (n17632, pi0140, n17631);
  not g26930 (n_12244, n17632);
  and g26931 (n17633, n_11912, n_12244);
  not g26932 (n_12245, n17630);
  and g26933 (n17634, n_12245, n17633);
  not g26934 (n_12246, n17634);
  and g26935 (n17635, n_162, n_12246);
  not g26936 (n_12247, n17628);
  and g26937 (n17636, n_12247, n17635);
  not g26938 (n_12248, n17636);
  and g26939 (n17637, n_161, n_12248);
  not g26940 (n_12249, n17610);
  and g26941 (n17638, n_12249, n17637);
  and g26942 (n17639, pi0140, n_12121);
  and g26943 (n17640, n2521, n17639);
  not g26944 (n_12250, n17490);
  and g26945 (n17641, n_6245, n_12250);
  not g26946 (n_12251, n17640);
  and g26947 (n17642, n_11912, n_12251);
  not g26948 (n_12252, n17641);
  and g26949 (n17643, n_12252, n17642);
  and g26950 (n17644, n_6245, n_11432);
  and g26951 (n17645, n16667, n17355);
  not g26952 (n_12253, n17644);
  and g26953 (n17646, pi0761, n_12253);
  not g26954 (n_12254, n17645);
  and g26955 (n17647, n_12254, n17646);
  not g26956 (n_12255, n17643);
  not g26957 (n_12256, n17647);
  and g26958 (n17648, n_12255, n_12256);
  not g26959 (n_12257, n17648);
  and g26960 (n17649, n_162, n_12257);
  and g26961 (n17650, pi0038, n_11577);
  not g26962 (n_12258, n17649);
  and g26963 (n17651, n_12258, n17650);
  not g26964 (n_12259, n17638);
  not g26965 (n_12260, n17651);
  and g26966 (n17652, n_12259, n_12260);
  not g26967 (n_12261, n17652);
  and g26968 (n17653, n_11667, n_12261);
  not g26969 (n_12262, n17319);
  and g26970 (n17654, n2571, n_12262);
  not g26971 (n_12263, n17653);
  and g26972 (n17655, n_12263, n17654);
  not g26973 (n_12264, n17655);
  and g26974 (n17656, n_11746, n_12264);
  and g26975 (n17657, n_11753, n17656);
  and g26976 (n17658, pi0625, n17286);
  not g26977 (n_12265, n17658);
  and g26978 (n17659, n_11757, n_12265);
  not g26979 (n_12266, n17657);
  and g26980 (n17660, n_12266, n17659);
  and g26981 (n17661, n_11823, n_11760);
  not g26982 (n_12267, n17660);
  and g26983 (n17662, n_12267, n17661);
  and g26984 (n17663, n_11753, n17286);
  and g26985 (n17664, pi0625, n17656);
  not g26986 (n_12268, n17663);
  and g26987 (n17665, pi1153, n_12268);
  not g26988 (n_12269, n17664);
  and g26989 (n17666, n_12269, n17665);
  and g26990 (n17667, pi0608, n_11761);
  not g26991 (n_12270, n17666);
  and g26992 (n17668, n_12270, n17667);
  not g26993 (n_12271, n17662);
  not g26994 (n_12272, n17668);
  and g26995 (n17669, n_12271, n_12272);
  not g26996 (n_12273, n17669);
  and g26997 (n17670, pi0778, n_12273);
  and g26998 (n17671, n_11749, n17656);
  not g26999 (n_12274, n17670);
  not g27000 (n_12275, n17671);
  and g27001 (n17672, n_12274, n_12275);
  not g27002 (n_12276, n17672);
  and g27003 (n17673, n_11971, n_12276);
  and g27004 (n17674, pi0609, n17071);
  not g27005 (n_12277, n17674);
  and g27006 (n17675, n_11768, n_12277);
  not g27007 (n_12278, n17673);
  and g27008 (n17676, n_12278, n17675);
  and g27009 (n17677, n_11767, n_11976);
  not g27010 (n_12279, n17676);
  and g27011 (n17678, n_12279, n17677);
  and g27012 (n17679, n_11971, n17071);
  and g27013 (n17680, pi0609, n_12276);
  not g27014 (n_12280, n17679);
  and g27015 (n17681, pi1155, n_12280);
  not g27016 (n_12281, n17680);
  and g27017 (n17682, n_12281, n17681);
  and g27018 (n17683, pi0660, n_11977);
  not g27019 (n_12282, n17682);
  and g27020 (n17684, n_12282, n17683);
  not g27021 (n_12283, n17678);
  not g27022 (n_12284, n17684);
  and g27023 (n17685, n_12283, n_12284);
  not g27024 (n_12285, n17685);
  and g27025 (n17686, pi0785, n_12285);
  and g27026 (n17687, n_11964, n_12276);
  not g27027 (n_12286, n17686);
  not g27028 (n_12287, n17687);
  and g27029 (n17688, n_12286, n_12287);
  not g27030 (n_12288, n17688);
  and g27031 (n17689, n_11984, n_12288);
  and g27032 (n17690, pi0618, n17078);
  not g27033 (n_12289, n17690);
  and g27034 (n17691, n_11413, n_12289);
  not g27035 (n_12290, n17689);
  and g27036 (n17692, n_12290, n17691);
  and g27037 (n17693, n_11412, n_11989);
  not g27038 (n_12291, n17692);
  and g27039 (n17694, n_12291, n17693);
  and g27040 (n17695, n_11984, n17078);
  and g27041 (n17696, pi0618, n_12288);
  not g27042 (n_12292, n17695);
  and g27043 (n17697, pi1154, n_12292);
  not g27044 (n_12293, n17696);
  and g27045 (n17698, n_12293, n17697);
  and g27046 (n17699, pi0627, n_11990);
  not g27047 (n_12294, n17698);
  and g27048 (n17700, n_12294, n17699);
  not g27049 (n_12295, n17694);
  not g27050 (n_12296, n17700);
  and g27051 (n17701, n_12295, n_12296);
  not g27052 (n_12297, n17701);
  and g27053 (n17702, pi0781, n_12297);
  and g27054 (n17703, n_11981, n_12288);
  not g27055 (n_12298, n17702);
  not g27056 (n_12299, n17703);
  and g27057 (n17704, n_12298, n_12299);
  not g27058 (n_12300, n17704);
  and g27059 (n17705, n_11821, n_12300);
  not g27060 (n_12301, n17081);
  and g27061 (n17706, pi0619, n_12301);
  not g27062 (n_12302, n17706);
  and g27063 (n17707, n_11405, n_12302);
  not g27064 (n_12303, n17705);
  and g27065 (n17708, n_12303, n17707);
  not g27066 (n_12304, n17318);
  and g27067 (n17709, n_11403, n_12304);
  not g27068 (n_12305, n17708);
  and g27069 (n17710, n_12305, n17709);
  and g27070 (n17711, n_11821, n17315);
  and g27071 (n17712, pi0619, n17060);
  not g27072 (n_12306, n17712);
  and g27073 (n17713, n_11405, n_12306);
  not g27074 (n_12307, n17711);
  and g27075 (n17714, n_12307, n17713);
  and g27076 (n17715, pi0619, n_12300);
  and g27077 (n17716, n_11821, n_12301);
  not g27078 (n_12308, n17716);
  and g27079 (n17717, pi1159, n_12308);
  not g27080 (n_12309, n17715);
  and g27081 (n17718, n_12309, n17717);
  not g27082 (n_12310, n17714);
  and g27083 (n17719, pi0648, n_12310);
  not g27084 (n_12311, n17718);
  and g27085 (n17720, n_12311, n17719);
  not g27086 (n_12312, n17710);
  not g27087 (n_12313, n17720);
  and g27088 (n17721, n_12312, n_12313);
  not g27089 (n_12314, n17721);
  and g27090 (n17722, pi0789, n_12314);
  not g27091 (n_12315, pi0789);
  and g27092 (n17723, n_12315, n_12300);
  not g27093 (n_12316, n17722);
  not g27094 (n_12317, n17723);
  and g27095 (n17724, n_12316, n_12317);
  not g27096 (n_12318, pi0788);
  and g27097 (n17725, n_12318, n17724);
  not g27098 (n_12320, pi0626);
  and g27099 (n17726, n_12320, n17724);
  not g27100 (n_12321, n17084);
  and g27101 (n17727, pi0626, n_12321);
  not g27102 (n_12322, n17727);
  and g27103 (n17728, n_11395, n_12322);
  not g27104 (n_12323, n17726);
  and g27105 (n17729, n_12323, n17728);
  and g27106 (n17730, n_11395, n_11397);
  not g27107 (n_12324, n17315);
  and g27108 (n17731, n_12315, n_12324);
  and g27109 (n17732, n_12304, n_12310);
  not g27110 (n_12325, n17732);
  and g27111 (n17733, pi0789, n_12325);
  not g27112 (n_12326, n17731);
  not g27113 (n_12327, n17733);
  and g27114 (n17734, n_12326, n_12327);
  and g27115 (n17735, n_12320, n17734);
  and g27116 (n17736, pi0626, n17060);
  not g27117 (n_12328, n17736);
  and g27118 (n17737, n_11397, n_12328);
  not g27119 (n_12329, n17735);
  and g27120 (n17738, n_12329, n17737);
  not g27121 (n_12330, n17730);
  not g27122 (n_12331, n17738);
  and g27123 (n17739, n_12330, n_12331);
  not g27124 (n_12332, n17729);
  not g27125 (n_12333, n17739);
  and g27126 (n17740, n_12332, n_12333);
  and g27127 (n17741, pi0626, n17724);
  and g27128 (n17742, n_12320, n_12321);
  not g27129 (n_12334, n17742);
  and g27130 (n17743, pi0641, n_12334);
  not g27131 (n_12335, n17741);
  and g27132 (n17744, n_12335, n17743);
  and g27133 (n17745, pi0641, pi1158);
  and g27134 (n17746, n_12320, n17060);
  and g27135 (n17747, pi0626, n17734);
  not g27136 (n_12336, n17746);
  and g27137 (n17748, pi1158, n_12336);
  not g27138 (n_12337, n17747);
  and g27139 (n17749, n_12337, n17748);
  not g27140 (n_12338, n17745);
  not g27141 (n_12339, n17749);
  and g27142 (n17750, n_12338, n_12339);
  not g27143 (n_12340, n17744);
  not g27144 (n_12341, n17750);
  and g27145 (n17751, n_12340, n_12341);
  not g27146 (n_12342, n17740);
  not g27147 (n_12343, n17751);
  and g27148 (n17752, n_12342, n_12343);
  not g27149 (n_12344, n17752);
  and g27150 (n17753, pi0788, n_12344);
  not g27151 (n_12345, n17725);
  not g27152 (n_12346, n17753);
  and g27153 (n17754, n_12345, n_12346);
  and g27154 (n17755, n_11789, n17754);
  and g27155 (n17756, n_12331, n_12339);
  not g27156 (n_12347, n17756);
  and g27157 (n17757, pi0788, n_12347);
  not g27158 (n_12348, n17734);
  and g27159 (n17758, n_12318, n_12348);
  not g27160 (n_12349, n17757);
  not g27161 (n_12350, n17758);
  and g27162 (n17759, n_12349, n_12350);
  and g27163 (n17760, pi0628, n17759);
  not g27164 (n_12351, n17760);
  and g27165 (n17761, n_11794, n_12351);
  not g27166 (n_12352, n17755);
  and g27167 (n17762, n_12352, n17761);
  not g27168 (n_12354, pi0629);
  and g27169 (n17763, n_12354, n_11797);
  not g27170 (n_12355, n17762);
  and g27171 (n17764, n_12355, n17763);
  and g27172 (n17765, pi0628, n17754);
  and g27173 (n17766, n_11789, n17759);
  not g27174 (n_12356, n17766);
  and g27175 (n17767, pi1156, n_12356);
  not g27176 (n_12357, n17765);
  and g27177 (n17768, n_12357, n17767);
  and g27178 (n17769, pi0629, n_11798);
  not g27179 (n_12358, n17768);
  and g27180 (n17770, n_12358, n17769);
  not g27181 (n_12359, n17764);
  not g27182 (n_12360, n17770);
  and g27183 (n17771, n_12359, n_12360);
  not g27184 (n_12361, n17771);
  and g27185 (n17772, pi0792, n_12361);
  and g27186 (n17773, n_11787, n17754);
  not g27187 (n_12362, n17772);
  not g27188 (n_12363, n17773);
  and g27189 (n17774, n_12362, n_12363);
  not g27190 (n_12364, n17774);
  and g27191 (n17775, n_11806, n_12364);
  and g27192 (n17776, n_12354, pi1156);
  and g27193 (n17777, pi0629, n_11794);
  not g27194 (n_12365, n17776);
  not g27195 (n_12366, n17777);
  and g27196 (n17778, n_12365, n_12366);
  not g27197 (n_12367, n17778);
  and g27198 (n17779, pi0792, n_12367);
  not g27199 (n_12368, n17779);
  and g27200 (n17780, n17759, n_12368);
  and g27201 (n17781, n17060, n17779);
  not g27202 (n_12369, n17780);
  not g27203 (n_12370, n17781);
  and g27204 (n17782, n_12369, n_12370);
  not g27205 (n_12371, n17782);
  and g27206 (n17783, pi0647, n_12371);
  not g27207 (n_12372, n17783);
  and g27208 (n17784, n_11810, n_12372);
  not g27209 (n_12373, n17775);
  and g27210 (n17785, n_12373, n17784);
  not g27211 (n_12375, pi0630);
  and g27212 (n17786, n_12375, n_11813);
  not g27213 (n_12376, n17785);
  and g27214 (n17787, n_12376, n17786);
  and g27215 (n17788, pi0647, n_12364);
  and g27216 (n17789, n_11806, n_12371);
  not g27217 (n_12377, n17789);
  and g27218 (n17790, pi1157, n_12377);
  not g27219 (n_12378, n17788);
  and g27220 (n17791, n_12378, n17790);
  and g27221 (n17792, pi0630, n_11814);
  not g27222 (n_12379, n17791);
  and g27223 (n17793, n_12379, n17792);
  not g27224 (n_12380, n17787);
  not g27225 (n_12381, n17793);
  and g27226 (n17794, n_12380, n_12381);
  not g27227 (n_12382, n17794);
  and g27228 (n17795, pi0787, n_12382);
  and g27229 (n17796, n_11803, n_12364);
  not g27230 (n_12383, n17795);
  not g27231 (n_12384, n17796);
  and g27232 (n17797, n_12383, n_12384);
  not g27233 (n_12385, n17797);
  and g27234 (n17798, pi0644, n_12385);
  not g27235 (n_12387, n17112);
  and g27236 (n17799, pi0715, n_12387);
  not g27237 (n_12388, n17798);
  and g27238 (n17800, n_12388, n17799);
  and g27239 (n17801, n_12375, pi1157);
  and g27240 (n17802, pi0630, n_11810);
  not g27241 (n_12389, n17801);
  not g27242 (n_12390, n17802);
  and g27243 (n17803, n_12389, n_12390);
  not g27244 (n_12391, n17803);
  and g27245 (n17804, pi0787, n_12391);
  not g27246 (n_12392, n17804);
  and g27247 (n17805, n17782, n_12392);
  and g27248 (n17806, n_11774, n17804);
  not g27249 (n_12393, n17805);
  not g27250 (n_12394, n17806);
  and g27251 (n17807, n_12393, n_12394);
  and g27252 (n17808, pi0644, n17807);
  and g27253 (n17809, n_11819, n17060);
  not g27254 (n_12395, pi0715);
  not g27255 (n_12396, n17809);
  and g27256 (n17810, n_12395, n_12396);
  not g27257 (n_12397, n17808);
  and g27258 (n17811, n_12397, n17810);
  not g27259 (n_12399, n17811);
  and g27260 (n17812, pi1160, n_12399);
  not g27261 (n_12400, n17800);
  and g27262 (n17813, n_12400, n17812);
  and g27263 (n17814, n_11819, n_12385);
  and g27264 (n17815, pi0644, n17111);
  not g27265 (n_12401, n17815);
  and g27266 (n17816, n_12395, n_12401);
  not g27267 (n_12402, n17814);
  and g27268 (n17817, n_12402, n17816);
  and g27269 (n17818, n_11819, n17807);
  and g27270 (n17819, pi0644, n17060);
  not g27271 (n_12403, n17819);
  and g27272 (n17820, pi0715, n_12403);
  not g27273 (n_12404, n17818);
  and g27274 (n17821, n_12404, n17820);
  not g27275 (n_12405, pi1160);
  not g27276 (n_12406, n17821);
  and g27277 (n17822, n_12405, n_12406);
  not g27278 (n_12407, n17817);
  and g27279 (n17823, n_12407, n17822);
  not g27280 (n_12409, n17813);
  and g27281 (n17824, pi0790, n_12409);
  not g27282 (n_12410, n17823);
  and g27283 (n17825, n_12410, n17824);
  not g27284 (n_12411, pi0790);
  and g27285 (n17826, n_12411, n17797);
  not g27286 (n_12412, n17826);
  and g27287 (n17827, n_4226, n_12412);
  not g27288 (n_12413, n17825);
  and g27289 (n17828, n_12413, n17827);
  and g27290 (n17829, n_6245, po1038);
  not g27291 (n_12415, pi0832);
  not g27292 (n_12416, n17829);
  and g27293 (n17830, n_12415, n_12416);
  not g27294 (n_12417, n17828);
  and g27295 (n17831, n_12417, n17830);
  not g27296 (n_12418, n2926);
  and g27297 (n17832, n_6245, n_12418);
  and g27298 (n17833, n_11806, n17832);
  and g27299 (n17834, n_11667, n16645);
  not g27300 (n_12419, n17832);
  not g27301 (n_12420, n17834);
  and g27302 (n17835, n_12419, n_12420);
  and g27303 (n17836, n_11749, n17835);
  and g27304 (n17837, n_11753, n17834);
  not g27305 (n_12421, n17835);
  not g27306 (n_12422, n17837);
  and g27307 (n17838, n_12421, n_12422);
  not g27308 (n_12423, n17838);
  and g27309 (n17839, pi1153, n_12423);
  and g27310 (n17840, n_11757, n_12419);
  and g27311 (n17841, n_12422, n17840);
  not g27312 (n_12424, n17839);
  not g27313 (n_12425, n17841);
  and g27314 (n17842, n_12424, n_12425);
  not g27315 (n_12426, n17842);
  and g27316 (n17843, pi0778, n_12426);
  not g27317 (n_12427, n17836);
  not g27318 (n_12428, n17843);
  and g27319 (n17844, n_12427, n_12428);
  and g27320 (n17845, n2926, n17075);
  not g27321 (n_12429, n17845);
  and g27322 (n17846, n17844, n_12429);
  and g27323 (n17847, n2926, n16639);
  not g27324 (n_12430, n17847);
  and g27325 (n17848, n17846, n_12430);
  and g27326 (n17849, n2926, n16635);
  not g27327 (n_12431, n17849);
  and g27328 (n17850, n17848, n_12431);
  and g27329 (n17851, n2926, n16631);
  not g27330 (n_12432, n17851);
  and g27331 (n17852, n17850, n_12432);
  and g27332 (n17853, n_11789, pi1156);
  and g27333 (n17854, pi0628, n_11794);
  not g27334 (n_12433, n17853);
  not g27335 (n_12434, n17854);
  and g27336 (n17855, n_12433, n_12434);
  not g27337 (n_12435, n17855);
  and g27338 (n17856, pi0792, n_12435);
  and g27339 (n17857, n2926, n17856);
  not g27340 (n_12436, n17857);
  and g27341 (n17858, n17852, n_12436);
  and g27342 (n17859, pi0647, n17858);
  not g27343 (n_12437, n17833);
  and g27344 (n17860, pi1157, n_12437);
  not g27345 (n_12438, n17859);
  and g27346 (n17861, n_12438, n17860);
  and g27347 (n17862, n_11789, n2926);
  not g27348 (n_12439, n17862);
  and g27349 (n17863, n17852, n_12439);
  not g27350 (n_12440, n17863);
  and g27351 (n17864, pi1156, n_12440);
  and g27352 (n17865, n_12320, pi1158);
  and g27353 (n17866, pi0626, n_11397);
  not g27354 (n_12441, n17865);
  not g27355 (n_12442, n17866);
  and g27356 (n17867, n_12441, n_12442);
  and g27357 (n17868, n_12320, pi0641);
  and g27358 (n17869, pi0626, n_11395);
  not g27359 (n_12443, n17868);
  not g27360 (n_12444, n17869);
  and g27361 (n17870, n_12443, n_12444);
  not g27362 (n_12445, n17867);
  not g27363 (n_12446, n17870);
  and g27364 (n17871, n_12445, n_12446);
  and g27365 (n17872, n17850, n17871);
  and g27366 (n17873, n_12320, n17832);
  and g27367 (n17874, n2926, n17117);
  and g27368 (n17875, n_11912, n17244);
  not g27369 (n_12447, n17875);
  and g27370 (n17876, n_12419, n_12447);
  not g27371 (n_12448, n17874);
  not g27372 (n_12449, n17876);
  and g27373 (n17877, n_12448, n_12449);
  not g27374 (n_12450, n17877);
  and g27375 (n17878, n_11964, n_12450);
  and g27376 (n17879, n2926, n_11967);
  not g27377 (n_12451, n17879);
  and g27378 (n17880, n_12449, n_12451);
  not g27379 (n_12452, n17880);
  and g27380 (n17881, pi1155, n_12452);
  and g27381 (n17882, pi0609, n2926);
  not g27382 (n_12453, n17882);
  and g27383 (n17883, n17877, n_12453);
  not g27384 (n_12454, n17883);
  and g27385 (n17884, n_11768, n_12454);
  not g27386 (n_12455, n17881);
  not g27387 (n_12456, n17884);
  and g27388 (n17885, n_12455, n_12456);
  not g27389 (n_12457, n17885);
  and g27390 (n17886, pi0785, n_12457);
  not g27391 (n_12458, n17878);
  not g27392 (n_12459, n17886);
  and g27393 (n17887, n_12458, n_12459);
  not g27394 (n_12460, n17887);
  and g27395 (n17888, n_11981, n_12460);
  and g27396 (n17889, n_11984, n2926);
  not g27397 (n_12461, n17889);
  and g27398 (n17890, n17887, n_12461);
  not g27399 (n_12462, n17890);
  and g27400 (n17891, pi1154, n_12462);
  and g27401 (n17892, pi0618, n2926);
  not g27402 (n_12463, n17892);
  and g27403 (n17893, n17887, n_12463);
  not g27404 (n_12464, n17893);
  and g27405 (n17894, n_11413, n_12464);
  not g27406 (n_12465, n17891);
  not g27407 (n_12466, n17894);
  and g27408 (n17895, n_12465, n_12466);
  not g27409 (n_12467, n17895);
  and g27410 (n17896, pi0781, n_12467);
  not g27411 (n_12468, n17888);
  not g27412 (n_12469, n17896);
  and g27413 (n17897, n_12468, n_12469);
  not g27414 (n_12470, n17897);
  and g27415 (n17898, n_12315, n_12470);
  and g27416 (n17899, n_11821, n17832);
  and g27417 (n17900, pi0619, n17897);
  not g27418 (n_12471, n17899);
  and g27419 (n17901, pi1159, n_12471);
  not g27420 (n_12472, n17900);
  and g27421 (n17902, n_12472, n17901);
  and g27422 (n17903, n_11821, n17897);
  and g27423 (n17904, pi0619, n17832);
  not g27424 (n_12473, n17904);
  and g27425 (n17905, n_11405, n_12473);
  not g27426 (n_12474, n17903);
  and g27427 (n17906, n_12474, n17905);
  not g27428 (n_12475, n17902);
  not g27429 (n_12476, n17906);
  and g27430 (n17907, n_12475, n_12476);
  not g27431 (n_12477, n17907);
  and g27432 (n17908, pi0789, n_12477);
  not g27433 (n_12478, n17898);
  not g27434 (n_12479, n17908);
  and g27435 (n17909, n_12478, n_12479);
  and g27436 (n17910, pi0626, n17909);
  not g27437 (n_12480, n17873);
  and g27438 (n17911, pi1158, n_12480);
  not g27439 (n_12481, n17910);
  and g27440 (n17912, n_12481, n17911);
  and g27441 (n17913, n_12320, n17909);
  and g27442 (n17914, pi0626, n17832);
  not g27443 (n_12482, n17914);
  and g27444 (n17915, n_11397, n_12482);
  not g27445 (n_12483, n17913);
  and g27446 (n17916, n_12483, n17915);
  not g27447 (n_12484, n17912);
  not g27448 (n_12485, n17916);
  and g27449 (n17917, n_12484, n_12485);
  and g27450 (n17918, n_11401, n17917);
  not g27451 (n_12486, n17872);
  not g27452 (n_12487, n17918);
  and g27453 (n17919, n_12486, n_12487);
  not g27454 (n_12488, n17919);
  and g27455 (n17920, pi0788, n_12488);
  and g27456 (n17921, pi0618, n17846);
  and g27457 (n17922, pi0609, n17844);
  and g27458 (n17923, n_11866, n_12421);
  and g27459 (n17924, pi0625, n17923);
  not g27460 (n_12489, n17923);
  and g27461 (n17925, n17876, n_12489);
  not g27462 (n_12490, n17924);
  not g27463 (n_12491, n17925);
  and g27464 (n17926, n_12490, n_12491);
  not g27465 (n_12492, n17926);
  and g27466 (n17927, n17840, n_12492);
  and g27467 (n17928, n_11823, n_12424);
  not g27468 (n_12493, n17927);
  and g27469 (n17929, n_12493, n17928);
  and g27470 (n17930, pi1153, n17876);
  and g27471 (n17931, n_12490, n17930);
  and g27472 (n17932, pi0608, n_12425);
  not g27473 (n_12494, n17931);
  and g27474 (n17933, n_12494, n17932);
  not g27475 (n_12495, n17929);
  not g27476 (n_12496, n17933);
  and g27477 (n17934, n_12495, n_12496);
  not g27478 (n_12497, n17934);
  and g27479 (n17935, pi0778, n_12497);
  and g27480 (n17936, n_11749, n_12491);
  not g27481 (n_12498, n17935);
  not g27482 (n_12499, n17936);
  and g27483 (n17937, n_12498, n_12499);
  not g27484 (n_12500, n17937);
  and g27485 (n17938, n_11971, n_12500);
  not g27486 (n_12501, n17922);
  and g27487 (n17939, n_11768, n_12501);
  not g27488 (n_12502, n17938);
  and g27489 (n17940, n_12502, n17939);
  and g27490 (n17941, n_11767, n_12455);
  not g27491 (n_12503, n17940);
  and g27492 (n17942, n_12503, n17941);
  and g27493 (n17943, n_11971, n17844);
  and g27494 (n17944, pi0609, n_12500);
  not g27495 (n_12504, n17943);
  and g27496 (n17945, pi1155, n_12504);
  not g27497 (n_12505, n17944);
  and g27498 (n17946, n_12505, n17945);
  and g27499 (n17947, pi0660, n_12456);
  not g27500 (n_12506, n17946);
  and g27501 (n17948, n_12506, n17947);
  not g27502 (n_12507, n17942);
  not g27503 (n_12508, n17948);
  and g27504 (n17949, n_12507, n_12508);
  not g27505 (n_12509, n17949);
  and g27506 (n17950, pi0785, n_12509);
  and g27507 (n17951, n_11964, n_12500);
  not g27508 (n_12510, n17950);
  not g27509 (n_12511, n17951);
  and g27510 (n17952, n_12510, n_12511);
  not g27511 (n_12512, n17952);
  and g27512 (n17953, n_11984, n_12512);
  not g27513 (n_12513, n17921);
  and g27514 (n17954, n_11413, n_12513);
  not g27515 (n_12514, n17953);
  and g27516 (n17955, n_12514, n17954);
  and g27517 (n17956, n_11412, n_12465);
  not g27518 (n_12515, n17955);
  and g27519 (n17957, n_12515, n17956);
  and g27520 (n17958, n_11984, n17846);
  and g27521 (n17959, pi0618, n_12512);
  not g27522 (n_12516, n17958);
  and g27523 (n17960, pi1154, n_12516);
  not g27524 (n_12517, n17959);
  and g27525 (n17961, n_12517, n17960);
  and g27526 (n17962, pi0627, n_12466);
  not g27527 (n_12518, n17961);
  and g27528 (n17963, n_12518, n17962);
  not g27529 (n_12519, n17957);
  not g27530 (n_12520, n17963);
  and g27531 (n17964, n_12519, n_12520);
  not g27532 (n_12521, n17964);
  and g27533 (n17965, pi0781, n_12521);
  and g27534 (n17966, n_11981, n_12512);
  not g27535 (n_12522, n17965);
  not g27536 (n_12523, n17966);
  and g27537 (n17967, n_12522, n_12523);
  and g27538 (n17968, n_12315, n17967);
  and g27539 (n17969, pi0788, n_12445);
  not g27540 (n_12524, n17969);
  and g27541 (n17970, n_11783, n_12524);
  not g27542 (n_12525, n17967);
  and g27543 (n17971, n_11821, n_12525);
  and g27544 (n17972, pi0619, n17848);
  not g27545 (n_12526, n17972);
  and g27546 (n17973, n_11405, n_12526);
  not g27547 (n_12527, n17971);
  and g27548 (n17974, n_12527, n17973);
  and g27549 (n17975, n_11403, n_12475);
  not g27550 (n_12528, n17974);
  and g27551 (n17976, n_12528, n17975);
  and g27552 (n17977, n_11821, n17848);
  and g27553 (n17978, pi0619, n_12525);
  not g27554 (n_12529, n17977);
  and g27555 (n17979, pi1159, n_12529);
  not g27556 (n_12530, n17978);
  and g27557 (n17980, n_12530, n17979);
  and g27558 (n17981, pi0648, n_12476);
  not g27559 (n_12531, n17980);
  and g27560 (n17982, n_12531, n17981);
  not g27561 (n_12532, n17976);
  and g27562 (n17983, pi0789, n_12532);
  not g27563 (n_12533, n17982);
  and g27564 (n17984, n_12533, n17983);
  not g27565 (n_12534, n17968);
  and g27566 (n17985, n_12534, n17970);
  not g27567 (n_12535, n17984);
  and g27568 (n17986, n_12535, n17985);
  not g27569 (n_12536, n17920);
  not g27570 (n_12537, n17986);
  and g27571 (n17987, n_12536, n_12537);
  not g27572 (n_12538, n17987);
  and g27573 (n17988, n_11789, n_12538);
  not g27574 (n_12539, n17909);
  and g27575 (n17989, n_12318, n_12539);
  not g27576 (n_12540, n17917);
  and g27577 (n17990, pi0788, n_12540);
  not g27578 (n_12541, n17989);
  not g27579 (n_12542, n17990);
  and g27580 (n17991, n_12541, n_12542);
  and g27581 (n17992, pi0628, n17991);
  not g27582 (n_12543, n17992);
  and g27583 (n17993, n_11794, n_12543);
  not g27584 (n_12544, n17988);
  and g27585 (n17994, n_12544, n17993);
  not g27586 (n_12545, n17864);
  and g27587 (n17995, n_12354, n_12545);
  not g27588 (n_12546, n17994);
  and g27589 (n17996, n_12546, n17995);
  and g27590 (n17997, pi0628, n2926);
  not g27591 (n_12547, n17997);
  and g27592 (n17998, n17852, n_12547);
  not g27593 (n_12548, n17998);
  and g27594 (n17999, n_11794, n_12548);
  and g27595 (n18000, n_11789, n17991);
  and g27596 (n18001, pi0628, n_12538);
  not g27597 (n_12549, n18000);
  and g27598 (n18002, pi1156, n_12549);
  not g27599 (n_12550, n18001);
  and g27600 (n18003, n_12550, n18002);
  not g27601 (n_12551, n17999);
  and g27602 (n18004, pi0629, n_12551);
  not g27603 (n_12552, n18003);
  and g27604 (n18005, n_12552, n18004);
  not g27605 (n_12553, n17996);
  not g27606 (n_12554, n18005);
  and g27607 (n18006, n_12553, n_12554);
  not g27608 (n_12555, n18006);
  and g27609 (n18007, pi0792, n_12555);
  and g27610 (n18008, n_11787, n_12538);
  not g27611 (n_12556, n18007);
  not g27612 (n_12557, n18008);
  and g27613 (n18009, n_12556, n_12557);
  not g27614 (n_12558, n18009);
  and g27615 (n18010, n_11806, n_12558);
  and g27616 (n18011, n_12368, n17991);
  and g27617 (n18012, n17779, n17832);
  not g27618 (n_12559, n18011);
  not g27619 (n_12560, n18012);
  and g27620 (n18013, n_12559, n_12560);
  not g27621 (n_12561, n18013);
  and g27622 (n18014, pi0647, n_12561);
  not g27623 (n_12562, n18014);
  and g27624 (n18015, n_11810, n_12562);
  not g27625 (n_12563, n18010);
  and g27626 (n18016, n_12563, n18015);
  not g27627 (n_12564, n17861);
  and g27628 (n18017, n_12375, n_12564);
  not g27629 (n_12565, n18016);
  and g27630 (n18018, n_12565, n18017);
  and g27631 (n18019, n_11806, n17858);
  and g27632 (n18020, pi0647, n17832);
  not g27633 (n_12566, n18020);
  and g27634 (n18021, n_11810, n_12566);
  not g27635 (n_12567, n18019);
  and g27636 (n18022, n_12567, n18021);
  and g27637 (n18023, pi0647, n_12558);
  and g27638 (n18024, n_11806, n_12561);
  not g27639 (n_12568, n18024);
  and g27640 (n18025, pi1157, n_12568);
  not g27641 (n_12569, n18023);
  and g27642 (n18026, n_12569, n18025);
  not g27643 (n_12570, n18022);
  and g27644 (n18027, pi0630, n_12570);
  not g27645 (n_12571, n18026);
  and g27646 (n18028, n_12571, n18027);
  not g27647 (n_12572, n18018);
  not g27648 (n_12573, n18028);
  and g27649 (n18029, n_12572, n_12573);
  not g27650 (n_12574, n18029);
  and g27651 (n18030, pi0787, n_12574);
  and g27652 (n18031, n_11803, n_12558);
  not g27653 (n_12575, n18030);
  not g27654 (n_12576, n18031);
  and g27655 (n18032, n_12575, n_12576);
  not g27656 (n_12577, n18032);
  and g27657 (n18033, n_12411, n_12577);
  not g27658 (n_12578, n17858);
  and g27659 (n18034, n_11803, n_12578);
  and g27660 (n18035, n_12564, n_12570);
  not g27661 (n_12579, n18035);
  and g27662 (n18036, pi0787, n_12579);
  not g27663 (n_12580, n18034);
  not g27664 (n_12581, n18036);
  and g27665 (n18037, n_12580, n_12581);
  and g27666 (n18038, n_11819, n18037);
  and g27667 (n18039, pi0644, n_12577);
  not g27668 (n_12582, n18038);
  and g27669 (n18040, pi0715, n_12582);
  not g27670 (n_12583, n18039);
  and g27671 (n18041, n_12583, n18040);
  and g27672 (n18042, n17804, n_12419);
  and g27673 (n18043, n_12392, n18013);
  not g27674 (n_12584, n18042);
  not g27675 (n_12585, n18043);
  and g27676 (n18044, n_12584, n_12585);
  and g27677 (n18045, pi0644, n18044);
  and g27678 (n18046, n_11819, n17832);
  not g27679 (n_12586, n18046);
  and g27680 (n18047, n_12395, n_12586);
  not g27681 (n_12587, n18045);
  and g27682 (n18048, n_12587, n18047);
  not g27683 (n_12588, n18048);
  and g27684 (n18049, pi1160, n_12588);
  not g27685 (n_12589, n18041);
  and g27686 (n18050, n_12589, n18049);
  and g27687 (n18051, n_11819, n18044);
  and g27688 (n18052, pi0644, n17832);
  not g27689 (n_12590, n18052);
  and g27690 (n18053, pi0715, n_12590);
  not g27691 (n_12591, n18051);
  and g27692 (n18054, n_12591, n18053);
  and g27693 (n18055, pi0644, n18037);
  and g27694 (n18056, n_11819, n_12577);
  not g27695 (n_12592, n18055);
  and g27696 (n18057, n_12395, n_12592);
  not g27697 (n_12593, n18056);
  and g27698 (n18058, n_12593, n18057);
  not g27699 (n_12594, n18054);
  and g27700 (n18059, n_12405, n_12594);
  not g27701 (n_12595, n18058);
  and g27702 (n18060, n_12595, n18059);
  not g27703 (n_12596, n18050);
  not g27704 (n_12597, n18060);
  and g27705 (n18061, n_12596, n_12597);
  not g27706 (n_12598, n18061);
  and g27707 (n18062, pi0790, n_12598);
  not g27708 (n_12599, n18033);
  and g27709 (n18063, pi0832, n_12599);
  not g27710 (n_12600, n18062);
  and g27711 (n18064, n_12600, n18063);
  not g27712 (n_12601, n17831);
  not g27713 (n_12602, n18064);
  and g27714 (po0297, n_12601, n_12602);
  and g27715 (n18066, n_11220, n_11751);
  not g27716 (n_12603, n18066);
  and g27717 (n18067, n16635, n_12603);
  and g27718 (n18068, pi0141, n_11417);
  and g27719 (n18069, n_11220, n_11418);
  not g27720 (n_12604, n18069);
  and g27721 (n18070, n16647, n_12604);
  and g27722 (n18071, n_162, n16948);
  not g27723 (n_12605, n18071);
  and g27724 (n18072, n_11578, n_12605);
  and g27725 (n18073, n_11220, n18072);
  and g27726 (n18074, pi0039, n_11500);
  and g27727 (n18075, n_162, n16926);
  not g27728 (n_12606, n18074);
  not g27729 (n_12607, n18075);
  and g27730 (n18076, n_12606, n_12607);
  not g27731 (n_12608, n18076);
  and g27732 (n18077, pi0141, n_12608);
  not g27733 (n_12609, n18077);
  and g27734 (n18078, n_161, n_12609);
  not g27735 (n_12610, n18073);
  and g27736 (n18079, n_12610, n18078);
  not g27737 (n_12612, n18070);
  and g27738 (n18080, pi0706, n_12612);
  not g27739 (n_12613, n18079);
  and g27740 (n18081, n_12613, n18080);
  not g27741 (n_12614, pi0706);
  and g27742 (n18082, n_11220, n_12614);
  and g27743 (n18083, n_11743, n18082);
  not g27744 (n_12615, n18083);
  and g27745 (n18084, n2571, n_12615);
  not g27746 (n_12616, n18081);
  and g27747 (n18085, n_12616, n18084);
  not g27748 (n_12617, n18068);
  not g27749 (n_12618, n18085);
  and g27750 (n18086, n_12617, n_12618);
  not g27751 (n_12619, n18086);
  and g27752 (n18087, n_11749, n_12619);
  and g27753 (n18088, n_11753, n18066);
  and g27754 (n18089, pi0625, n18086);
  not g27755 (n_12620, n18088);
  and g27756 (n18090, pi1153, n_12620);
  not g27757 (n_12621, n18089);
  and g27758 (n18091, n_12621, n18090);
  and g27759 (n18092, n_11753, n18086);
  and g27760 (n18093, pi0625, n18066);
  not g27761 (n_12622, n18093);
  and g27762 (n18094, n_11757, n_12622);
  not g27763 (n_12623, n18092);
  and g27764 (n18095, n_12623, n18094);
  not g27765 (n_12624, n18091);
  not g27766 (n_12625, n18095);
  and g27767 (n18096, n_12624, n_12625);
  not g27768 (n_12626, n18096);
  and g27769 (n18097, pi0778, n_12626);
  not g27770 (n_12627, n18087);
  not g27771 (n_12628, n18097);
  and g27772 (n18098, n_12627, n_12628);
  not g27773 (n_12629, n18098);
  and g27774 (n18099, n_11773, n_12629);
  and g27775 (n18100, n17075, n_12603);
  not g27776 (n_12630, n18099);
  not g27777 (n_12631, n18100);
  and g27778 (n18101, n_12630, n_12631);
  and g27779 (n18102, n_11777, n18101);
  and g27780 (n18103, n16639, n18066);
  not g27781 (n_12632, n18102);
  not g27782 (n_12633, n18103);
  and g27783 (n18104, n_12632, n_12633);
  and g27784 (n18105, n_11780, n18104);
  not g27785 (n_12634, n18067);
  not g27786 (n_12635, n18105);
  and g27787 (n18106, n_12634, n_12635);
  and g27788 (n18107, n_11783, n18106);
  and g27789 (n18108, n16631, n18066);
  not g27790 (n_12636, n18107);
  not g27791 (n_12637, n18108);
  and g27792 (n18109, n_12636, n_12637);
  and g27793 (n18110, n_11787, n18109);
  and g27794 (n18111, n_11789, n18066);
  not g27795 (n_12638, n18109);
  and g27796 (n18112, pi0628, n_12638);
  not g27797 (n_12639, n18111);
  and g27798 (n18113, pi1156, n_12639);
  not g27799 (n_12640, n18112);
  and g27800 (n18114, n_12640, n18113);
  and g27801 (n18115, pi0628, n18066);
  and g27802 (n18116, n_11789, n_12638);
  not g27803 (n_12641, n18115);
  and g27804 (n18117, n_11794, n_12641);
  not g27805 (n_12642, n18116);
  and g27806 (n18118, n_12642, n18117);
  not g27807 (n_12643, n18114);
  not g27808 (n_12644, n18118);
  and g27809 (n18119, n_12643, n_12644);
  not g27810 (n_12645, n18119);
  and g27811 (n18120, pi0792, n_12645);
  not g27812 (n_12646, n18110);
  not g27813 (n_12647, n18120);
  and g27814 (n18121, n_12646, n_12647);
  not g27815 (n_12648, n18121);
  and g27816 (n18122, n_11803, n_12648);
  and g27817 (n18123, n_11806, n18066);
  and g27818 (n18124, pi0647, n18121);
  not g27819 (n_12649, n18123);
  and g27820 (n18125, pi1157, n_12649);
  not g27821 (n_12650, n18124);
  and g27822 (n18126, n_12650, n18125);
  and g27823 (n18127, n_11806, n18121);
  and g27824 (n18128, pi0647, n18066);
  not g27825 (n_12651, n18128);
  and g27826 (n18129, n_11810, n_12651);
  not g27827 (n_12652, n18127);
  and g27828 (n18130, n_12652, n18129);
  not g27829 (n_12653, n18126);
  not g27830 (n_12654, n18130);
  and g27831 (n18131, n_12653, n_12654);
  not g27832 (n_12655, n18131);
  and g27833 (n18132, pi0787, n_12655);
  not g27834 (n_12656, n18122);
  not g27835 (n_12657, n18132);
  and g27836 (n18133, n_12656, n_12657);
  and g27837 (n18134, n_11819, n18133);
  and g27838 (n18135, n_11984, n18066);
  and g27839 (n18136, pi0749, n17280);
  not g27840 (n_12659, n18136);
  and g27841 (n18137, n_12604, n_12659);
  not g27842 (n_12660, n18137);
  and g27843 (n18138, pi0038, n_12660);
  not g27844 (n_12661, pi0749);
  and g27845 (n18139, n_12661, n17046);
  and g27846 (n18140, pi0141, n17273);
  not g27847 (n_12662, n18139);
  not g27848 (n_12663, n18140);
  and g27849 (n18141, n_12662, n_12663);
  not g27850 (n_12664, n18141);
  and g27851 (n18142, pi0039, n_12664);
  and g27852 (n18143, n_11220, n17221);
  and g27853 (n18144, pi0141, n17234);
  not g27854 (n_12665, n18144);
  and g27855 (n18145, pi0749, n_12665);
  not g27856 (n_12666, n18143);
  and g27857 (n18146, n_12666, n18145);
  and g27858 (n18147, n_162, n16958);
  and g27859 (n18148, n_11220, n_12661);
  not g27860 (n_12667, n18147);
  and g27861 (n18149, n_12667, n18148);
  not g27862 (n_12668, n18146);
  not g27863 (n_12669, n18149);
  and g27864 (n18150, n_12668, n_12669);
  not g27865 (n_12670, n18150);
  and g27866 (n18151, n_161, n_12670);
  not g27867 (n_12671, n18142);
  and g27868 (n18152, n_12671, n18151);
  not g27869 (n_12672, n18138);
  not g27870 (n_12673, n18152);
  and g27871 (n18153, n_12672, n_12673);
  and g27872 (n18154, n2571, n18153);
  not g27873 (n_12674, n18154);
  and g27874 (n18155, n_12617, n_12674);
  not g27875 (n_12675, n18155);
  and g27876 (n18156, n_11960, n_12675);
  and g27877 (n18157, n17117, n_12603);
  not g27878 (n_12676, n18156);
  not g27879 (n_12677, n18157);
  and g27880 (n18158, n_12676, n_12677);
  not g27881 (n_12678, n18158);
  and g27882 (n18159, n_11964, n_12678);
  and g27883 (n18160, n_11967, n_12603);
  and g27884 (n18161, pi0609, n18156);
  not g27885 (n_12679, n18160);
  not g27886 (n_12680, n18161);
  and g27887 (n18162, n_12679, n_12680);
  not g27888 (n_12681, n18162);
  and g27889 (n18163, pi1155, n_12681);
  and g27890 (n18164, n_11972, n_12603);
  and g27891 (n18165, n_11971, n18156);
  not g27892 (n_12682, n18164);
  not g27893 (n_12683, n18165);
  and g27894 (n18166, n_12682, n_12683);
  not g27895 (n_12684, n18166);
  and g27896 (n18167, n_11768, n_12684);
  not g27897 (n_12685, n18163);
  not g27898 (n_12686, n18167);
  and g27899 (n18168, n_12685, n_12686);
  not g27900 (n_12687, n18168);
  and g27901 (n18169, pi0785, n_12687);
  not g27902 (n_12688, n18159);
  not g27903 (n_12689, n18169);
  and g27904 (n18170, n_12688, n_12689);
  and g27905 (n18171, pi0618, n18170);
  not g27906 (n_12690, n18135);
  and g27907 (n18172, pi1154, n_12690);
  not g27908 (n_12691, n18171);
  and g27909 (n18173, n_12691, n18172);
  not g27910 (n_12692, n18153);
  and g27911 (n18174, n_12614, n_12692);
  and g27912 (n18175, n_162, n17645);
  not g27913 (n_12693, n18175);
  and g27914 (n18176, pi0038, n_12693);
  and g27915 (n18177, n18137, n18176);
  not g27916 (n_12694, n17629);
  and g27917 (n18178, n_11220, n_12694);
  not g27918 (n_12695, n17631);
  and g27919 (n18179, pi0141, n_12695);
  not g27920 (n_12696, n18179);
  and g27921 (n18180, pi0749, n_12696);
  not g27922 (n_12697, n18178);
  and g27923 (n18181, n_12697, n18180);
  and g27924 (n18182, n_11220, n17612);
  and g27925 (n18183, pi0141, n17625);
  not g27926 (n_12698, n18182);
  and g27927 (n18184, n_12661, n_12698);
  not g27928 (n_12699, n18183);
  and g27929 (n18185, n_12699, n18184);
  not g27930 (n_12700, n18181);
  and g27931 (n18186, n_162, n_12700);
  not g27932 (n_12701, n18185);
  and g27933 (n18187, n_12701, n18186);
  and g27934 (n18188, pi0141, n17605);
  and g27935 (n18189, n_11220, n_12180);
  not g27936 (n_12702, n18189);
  and g27937 (n18190, pi0749, n_12702);
  not g27938 (n_12703, n18188);
  and g27939 (n18191, n_12703, n18190);
  and g27940 (n18192, n_11220, n17404);
  and g27941 (n18193, pi0141, n17485);
  not g27942 (n_12704, n18193);
  and g27943 (n18194, n_12661, n_12704);
  not g27944 (n_12705, n18192);
  and g27945 (n18195, n_12705, n18194);
  not g27946 (n_12706, n18191);
  and g27947 (n18196, pi0039, n_12706);
  not g27948 (n_12707, n18195);
  and g27949 (n18197, n_12707, n18196);
  not g27950 (n_12708, n18187);
  and g27951 (n18198, n_161, n_12708);
  not g27952 (n_12709, n18197);
  and g27953 (n18199, n_12709, n18198);
  not g27954 (n_12710, n18177);
  and g27955 (n18200, pi0706, n_12710);
  not g27956 (n_12711, n18199);
  and g27957 (n18201, n_12711, n18200);
  not g27958 (n_12712, n18174);
  and g27959 (n18202, n2571, n_12712);
  not g27960 (n_12713, n18201);
  and g27961 (n18203, n_12713, n18202);
  not g27962 (n_12714, n18203);
  and g27963 (n18204, n_12617, n_12714);
  and g27964 (n18205, n_11753, n18204);
  and g27965 (n18206, pi0625, n18155);
  not g27966 (n_12715, n18206);
  and g27967 (n18207, n_11757, n_12715);
  not g27968 (n_12716, n18205);
  and g27969 (n18208, n_12716, n18207);
  and g27970 (n18209, n_11823, n_12624);
  not g27971 (n_12717, n18208);
  and g27972 (n18210, n_12717, n18209);
  and g27973 (n18211, n_11753, n18155);
  and g27974 (n18212, pi0625, n18204);
  not g27975 (n_12718, n18211);
  and g27976 (n18213, pi1153, n_12718);
  not g27977 (n_12719, n18212);
  and g27978 (n18214, n_12719, n18213);
  and g27979 (n18215, pi0608, n_12625);
  not g27980 (n_12720, n18214);
  and g27981 (n18216, n_12720, n18215);
  not g27982 (n_12721, n18210);
  not g27983 (n_12722, n18216);
  and g27984 (n18217, n_12721, n_12722);
  not g27985 (n_12723, n18217);
  and g27986 (n18218, pi0778, n_12723);
  and g27987 (n18219, n_11749, n18204);
  not g27988 (n_12724, n18218);
  not g27989 (n_12725, n18219);
  and g27990 (n18220, n_12724, n_12725);
  not g27991 (n_12726, n18220);
  and g27992 (n18221, n_11971, n_12726);
  and g27993 (n18222, pi0609, n18098);
  not g27994 (n_12727, n18222);
  and g27995 (n18223, n_11768, n_12727);
  not g27996 (n_12728, n18221);
  and g27997 (n18224, n_12728, n18223);
  and g27998 (n18225, n_11767, n_12685);
  not g27999 (n_12729, n18224);
  and g28000 (n18226, n_12729, n18225);
  and g28001 (n18227, n_11971, n18098);
  and g28002 (n18228, pi0609, n_12726);
  not g28003 (n_12730, n18227);
  and g28004 (n18229, pi1155, n_12730);
  not g28005 (n_12731, n18228);
  and g28006 (n18230, n_12731, n18229);
  and g28007 (n18231, pi0660, n_12686);
  not g28008 (n_12732, n18230);
  and g28009 (n18232, n_12732, n18231);
  not g28010 (n_12733, n18226);
  not g28011 (n_12734, n18232);
  and g28012 (n18233, n_12733, n_12734);
  not g28013 (n_12735, n18233);
  and g28014 (n18234, pi0785, n_12735);
  and g28015 (n18235, n_11964, n_12726);
  not g28016 (n_12736, n18234);
  not g28017 (n_12737, n18235);
  and g28018 (n18236, n_12736, n_12737);
  not g28019 (n_12738, n18236);
  and g28020 (n18237, n_11984, n_12738);
  and g28021 (n18238, pi0618, n18101);
  not g28022 (n_12739, n18238);
  and g28023 (n18239, n_11413, n_12739);
  not g28024 (n_12740, n18237);
  and g28025 (n18240, n_12740, n18239);
  not g28026 (n_12741, n18173);
  and g28027 (n18241, n_11412, n_12741);
  not g28028 (n_12742, n18240);
  and g28029 (n18242, n_12742, n18241);
  and g28030 (n18243, n_11984, n18170);
  and g28031 (n18244, pi0618, n18066);
  not g28032 (n_12743, n18244);
  and g28033 (n18245, n_11413, n_12743);
  not g28034 (n_12744, n18243);
  and g28035 (n18246, n_12744, n18245);
  and g28036 (n18247, n_11984, n18101);
  and g28037 (n18248, pi0618, n_12738);
  not g28038 (n_12745, n18247);
  and g28039 (n18249, pi1154, n_12745);
  not g28040 (n_12746, n18248);
  and g28041 (n18250, n_12746, n18249);
  not g28042 (n_12747, n18246);
  and g28043 (n18251, pi0627, n_12747);
  not g28044 (n_12748, n18250);
  and g28045 (n18252, n_12748, n18251);
  not g28046 (n_12749, n18242);
  not g28047 (n_12750, n18252);
  and g28048 (n18253, n_12749, n_12750);
  not g28049 (n_12751, n18253);
  and g28050 (n18254, pi0781, n_12751);
  and g28051 (n18255, n_11981, n_12738);
  not g28052 (n_12752, n18254);
  not g28053 (n_12753, n18255);
  and g28054 (n18256, n_12752, n_12753);
  not g28055 (n_12754, n18256);
  and g28056 (n18257, n_11821, n_12754);
  not g28057 (n_12755, n18104);
  and g28058 (n18258, pi0619, n_12755);
  not g28059 (n_12756, n18258);
  and g28060 (n18259, n_11405, n_12756);
  not g28061 (n_12757, n18257);
  and g28062 (n18260, n_12757, n18259);
  and g28063 (n18261, n_11821, n18066);
  not g28064 (n_12758, n18170);
  and g28065 (n18262, n_11981, n_12758);
  and g28066 (n18263, n_12741, n_12747);
  not g28067 (n_12759, n18263);
  and g28068 (n18264, pi0781, n_12759);
  not g28069 (n_12760, n18262);
  not g28070 (n_12761, n18264);
  and g28071 (n18265, n_12760, n_12761);
  and g28072 (n18266, pi0619, n18265);
  not g28073 (n_12762, n18261);
  and g28074 (n18267, pi1159, n_12762);
  not g28075 (n_12763, n18266);
  and g28076 (n18268, n_12763, n18267);
  not g28077 (n_12764, n18268);
  and g28078 (n18269, n_11403, n_12764);
  not g28079 (n_12765, n18260);
  and g28080 (n18270, n_12765, n18269);
  and g28081 (n18271, pi0619, n_12754);
  and g28082 (n18272, n_11821, n_12755);
  not g28083 (n_12766, n18272);
  and g28084 (n18273, pi1159, n_12766);
  not g28085 (n_12767, n18271);
  and g28086 (n18274, n_12767, n18273);
  and g28087 (n18275, n_11821, n18265);
  and g28088 (n18276, pi0619, n18066);
  not g28089 (n_12768, n18276);
  and g28090 (n18277, n_11405, n_12768);
  not g28091 (n_12769, n18275);
  and g28092 (n18278, n_12769, n18277);
  not g28093 (n_12770, n18278);
  and g28094 (n18279, pi0648, n_12770);
  not g28095 (n_12771, n18274);
  and g28096 (n18280, n_12771, n18279);
  not g28097 (n_12772, n18270);
  not g28098 (n_12773, n18280);
  and g28099 (n18281, n_12772, n_12773);
  not g28100 (n_12774, n18281);
  and g28101 (n18282, pi0789, n_12774);
  and g28102 (n18283, n_12315, n_12754);
  not g28103 (n_12775, n18282);
  not g28104 (n_12776, n18283);
  and g28105 (n18284, n_12775, n_12776);
  and g28106 (n18285, n_12318, n18284);
  and g28107 (n18286, n_12320, n18284);
  not g28108 (n_12777, n18106);
  and g28109 (n18287, pi0626, n_12777);
  not g28110 (n_12778, n18287);
  and g28111 (n18288, n_11395, n_12778);
  not g28112 (n_12779, n18286);
  and g28113 (n18289, n_12779, n18288);
  not g28114 (n_12780, n18265);
  and g28115 (n18290, n_12315, n_12780);
  and g28116 (n18291, n_12764, n_12770);
  not g28117 (n_12781, n18291);
  and g28118 (n18292, pi0789, n_12781);
  not g28119 (n_12782, n18290);
  not g28120 (n_12783, n18292);
  and g28121 (n18293, n_12782, n_12783);
  and g28122 (n18294, n_12320, n18293);
  and g28123 (n18295, pi0626, n18066);
  not g28124 (n_12784, n18295);
  and g28125 (n18296, n_11397, n_12784);
  not g28126 (n_12785, n18294);
  and g28127 (n18297, n_12785, n18296);
  not g28128 (n_12786, n18297);
  and g28129 (n18298, n_12330, n_12786);
  not g28130 (n_12787, n18289);
  not g28131 (n_12788, n18298);
  and g28132 (n18299, n_12787, n_12788);
  and g28133 (n18300, pi0626, n18284);
  and g28134 (n18301, n_12320, n_12777);
  not g28135 (n_12789, n18301);
  and g28136 (n18302, pi0641, n_12789);
  not g28137 (n_12790, n18300);
  and g28138 (n18303, n_12790, n18302);
  and g28139 (n18304, n_12320, n18066);
  and g28140 (n18305, pi0626, n18293);
  not g28141 (n_12791, n18304);
  and g28142 (n18306, pi1158, n_12791);
  not g28143 (n_12792, n18305);
  and g28144 (n18307, n_12792, n18306);
  not g28145 (n_12793, n18307);
  and g28146 (n18308, n_12338, n_12793);
  not g28147 (n_12794, n18303);
  not g28148 (n_12795, n18308);
  and g28149 (n18309, n_12794, n_12795);
  not g28150 (n_12796, n18299);
  not g28151 (n_12797, n18309);
  and g28152 (n18310, n_12796, n_12797);
  not g28153 (n_12798, n18310);
  and g28154 (n18311, pi0788, n_12798);
  not g28155 (n_12799, n18285);
  not g28156 (n_12800, n18311);
  and g28157 (n18312, n_12799, n_12800);
  and g28158 (n18313, n_11789, n18312);
  and g28159 (n18314, n_12786, n_12793);
  not g28160 (n_12801, n18314);
  and g28161 (n18315, pi0788, n_12801);
  not g28162 (n_12802, n18293);
  and g28163 (n18316, n_12318, n_12802);
  not g28164 (n_12803, n18315);
  not g28165 (n_12804, n18316);
  and g28166 (n18317, n_12803, n_12804);
  and g28167 (n18318, pi0628, n18317);
  not g28168 (n_12805, n18318);
  and g28169 (n18319, n_11794, n_12805);
  not g28170 (n_12806, n18313);
  and g28171 (n18320, n_12806, n18319);
  and g28172 (n18321, n_12354, n_12643);
  not g28173 (n_12807, n18320);
  and g28174 (n18322, n_12807, n18321);
  and g28175 (n18323, pi0628, n18312);
  and g28176 (n18324, n_11789, n18317);
  not g28177 (n_12808, n18324);
  and g28178 (n18325, pi1156, n_12808);
  not g28179 (n_12809, n18323);
  and g28180 (n18326, n_12809, n18325);
  and g28181 (n18327, pi0629, n_12644);
  not g28182 (n_12810, n18326);
  and g28183 (n18328, n_12810, n18327);
  not g28184 (n_12811, n18322);
  not g28185 (n_12812, n18328);
  and g28186 (n18329, n_12811, n_12812);
  not g28187 (n_12813, n18329);
  and g28188 (n18330, pi0792, n_12813);
  and g28189 (n18331, n_11787, n18312);
  not g28190 (n_12814, n18330);
  not g28191 (n_12815, n18331);
  and g28192 (n18332, n_12814, n_12815);
  not g28193 (n_12816, n18332);
  and g28194 (n18333, n_11806, n_12816);
  and g28195 (n18334, n_12368, n18317);
  and g28196 (n18335, n17779, n18066);
  not g28197 (n_12817, n18334);
  not g28198 (n_12818, n18335);
  and g28199 (n18336, n_12817, n_12818);
  not g28200 (n_12819, n18336);
  and g28201 (n18337, pi0647, n_12819);
  not g28202 (n_12820, n18337);
  and g28203 (n18338, n_11810, n_12820);
  not g28204 (n_12821, n18333);
  and g28205 (n18339, n_12821, n18338);
  and g28206 (n18340, n_12375, n_12653);
  not g28207 (n_12822, n18339);
  and g28208 (n18341, n_12822, n18340);
  and g28209 (n18342, pi0647, n_12816);
  and g28210 (n18343, n_11806, n_12819);
  not g28211 (n_12823, n18343);
  and g28212 (n18344, pi1157, n_12823);
  not g28213 (n_12824, n18342);
  and g28214 (n18345, n_12824, n18344);
  and g28215 (n18346, pi0630, n_12654);
  not g28216 (n_12825, n18345);
  and g28217 (n18347, n_12825, n18346);
  not g28218 (n_12826, n18341);
  not g28219 (n_12827, n18347);
  and g28220 (n18348, n_12826, n_12827);
  not g28221 (n_12828, n18348);
  and g28222 (n18349, pi0787, n_12828);
  and g28223 (n18350, n_11803, n_12816);
  not g28224 (n_12829, n18349);
  not g28225 (n_12830, n18350);
  and g28226 (n18351, n_12829, n_12830);
  not g28227 (n_12831, n18351);
  and g28228 (n18352, pi0644, n_12831);
  not g28229 (n_12832, n18134);
  and g28230 (n18353, pi0715, n_12832);
  not g28231 (n_12833, n18352);
  and g28232 (n18354, n_12833, n18353);
  and g28233 (n18355, n17804, n_12603);
  and g28234 (n18356, n_12392, n18336);
  not g28235 (n_12834, n18355);
  not g28236 (n_12835, n18356);
  and g28237 (n18357, n_12834, n_12835);
  and g28238 (n18358, pi0644, n18357);
  and g28239 (n18359, n_11819, n18066);
  not g28240 (n_12836, n18359);
  and g28241 (n18360, n_12395, n_12836);
  not g28242 (n_12837, n18358);
  and g28243 (n18361, n_12837, n18360);
  not g28244 (n_12838, n18361);
  and g28245 (n18362, pi1160, n_12838);
  not g28246 (n_12839, n18354);
  and g28247 (n18363, n_12839, n18362);
  and g28248 (n18364, n_11819, n_12831);
  and g28249 (n18365, pi0644, n18133);
  not g28250 (n_12840, n18365);
  and g28251 (n18366, n_12395, n_12840);
  not g28252 (n_12841, n18364);
  and g28253 (n18367, n_12841, n18366);
  and g28254 (n18368, n_11819, n18357);
  and g28255 (n18369, pi0644, n18066);
  not g28256 (n_12842, n18369);
  and g28257 (n18370, pi0715, n_12842);
  not g28258 (n_12843, n18368);
  and g28259 (n18371, n_12843, n18370);
  not g28260 (n_12844, n18371);
  and g28261 (n18372, n_12405, n_12844);
  not g28262 (n_12845, n18367);
  and g28263 (n18373, n_12845, n18372);
  not g28264 (n_12846, n18363);
  and g28265 (n18374, pi0790, n_12846);
  not g28266 (n_12847, n18373);
  and g28267 (n18375, n_12847, n18374);
  and g28268 (n18376, n_12411, n18351);
  not g28269 (n_12848, n18376);
  and g28270 (n18377, n_4226, n_12848);
  not g28271 (n_12849, n18375);
  and g28272 (n18378, n_12849, n18377);
  and g28273 (n18379, n_11220, po1038);
  not g28274 (n_12850, n18379);
  and g28275 (n18380, n_12415, n_12850);
  not g28276 (n_12851, n18378);
  and g28277 (n18381, n_12851, n18380);
  and g28278 (n18382, n_11220, n_12418);
  and g28279 (n18383, n_11806, n18382);
  and g28280 (n18384, pi0706, n16645);
  not g28281 (n_12852, n18382);
  not g28282 (n_12853, n18384);
  and g28283 (n18385, n_12852, n_12853);
  and g28284 (n18386, n_11749, n18385);
  and g28285 (n18387, n_11753, n18384);
  not g28286 (n_12854, n18385);
  not g28287 (n_12855, n18387);
  and g28288 (n18388, n_12854, n_12855);
  not g28289 (n_12856, n18388);
  and g28290 (n18389, pi1153, n_12856);
  and g28291 (n18390, n_11757, n_12852);
  and g28292 (n18391, n_12855, n18390);
  not g28293 (n_12857, n18389);
  not g28294 (n_12858, n18391);
  and g28295 (n18392, n_12857, n_12858);
  not g28296 (n_12859, n18392);
  and g28297 (n18393, pi0778, n_12859);
  not g28298 (n_12860, n18386);
  not g28299 (n_12861, n18393);
  and g28300 (n18394, n_12860, n_12861);
  and g28301 (n18395, n_12429, n18394);
  and g28302 (n18396, n_12430, n18395);
  and g28303 (n18397, n_12431, n18396);
  and g28304 (n18398, n_12432, n18397);
  and g28305 (n18399, n_12436, n18398);
  and g28306 (n18400, pi0647, n18399);
  not g28307 (n_12862, n18383);
  and g28308 (n18401, pi1157, n_12862);
  not g28309 (n_12863, n18400);
  and g28310 (n18402, n_12863, n18401);
  and g28311 (n18403, n_12439, n18398);
  not g28312 (n_12864, n18403);
  and g28313 (n18404, pi1156, n_12864);
  and g28314 (n18405, n17871, n18397);
  and g28315 (n18406, n_12320, n18382);
  and g28316 (n18407, pi0749, n17244);
  not g28317 (n_12865, n18407);
  and g28318 (n18408, n_12852, n_12865);
  not g28319 (n_12866, n18408);
  and g28320 (n18409, n_12448, n_12866);
  not g28321 (n_12867, n18409);
  and g28322 (n18410, n_11964, n_12867);
  and g28323 (n18411, n_12451, n_12866);
  not g28324 (n_12868, n18411);
  and g28325 (n18412, pi1155, n_12868);
  and g28326 (n18413, n_12453, n18409);
  not g28327 (n_12869, n18413);
  and g28328 (n18414, n_11768, n_12869);
  not g28329 (n_12870, n18412);
  not g28330 (n_12871, n18414);
  and g28331 (n18415, n_12870, n_12871);
  not g28332 (n_12872, n18415);
  and g28333 (n18416, pi0785, n_12872);
  not g28334 (n_12873, n18410);
  not g28335 (n_12874, n18416);
  and g28336 (n18417, n_12873, n_12874);
  not g28337 (n_12875, n18417);
  and g28338 (n18418, n_11981, n_12875);
  and g28339 (n18419, n_12461, n18417);
  not g28340 (n_12876, n18419);
  and g28341 (n18420, pi1154, n_12876);
  and g28342 (n18421, n_12463, n18417);
  not g28343 (n_12877, n18421);
  and g28344 (n18422, n_11413, n_12877);
  not g28345 (n_12878, n18420);
  not g28346 (n_12879, n18422);
  and g28347 (n18423, n_12878, n_12879);
  not g28348 (n_12880, n18423);
  and g28349 (n18424, pi0781, n_12880);
  not g28350 (n_12881, n18418);
  not g28351 (n_12882, n18424);
  and g28352 (n18425, n_12881, n_12882);
  not g28353 (n_12883, n18425);
  and g28354 (n18426, n_12315, n_12883);
  and g28355 (n18427, n_11821, n18382);
  and g28356 (n18428, pi0619, n18425);
  not g28357 (n_12884, n18427);
  and g28358 (n18429, pi1159, n_12884);
  not g28359 (n_12885, n18428);
  and g28360 (n18430, n_12885, n18429);
  and g28361 (n18431, n_11821, n18425);
  and g28362 (n18432, pi0619, n18382);
  not g28363 (n_12886, n18432);
  and g28364 (n18433, n_11405, n_12886);
  not g28365 (n_12887, n18431);
  and g28366 (n18434, n_12887, n18433);
  not g28367 (n_12888, n18430);
  not g28368 (n_12889, n18434);
  and g28369 (n18435, n_12888, n_12889);
  not g28370 (n_12890, n18435);
  and g28371 (n18436, pi0789, n_12890);
  not g28372 (n_12891, n18426);
  not g28373 (n_12892, n18436);
  and g28374 (n18437, n_12891, n_12892);
  and g28375 (n18438, pi0626, n18437);
  not g28376 (n_12893, n18406);
  and g28377 (n18439, pi1158, n_12893);
  not g28378 (n_12894, n18438);
  and g28379 (n18440, n_12894, n18439);
  and g28380 (n18441, n_12320, n18437);
  and g28381 (n18442, pi0626, n18382);
  not g28382 (n_12895, n18442);
  and g28383 (n18443, n_11397, n_12895);
  not g28384 (n_12896, n18441);
  and g28385 (n18444, n_12896, n18443);
  not g28386 (n_12897, n18440);
  not g28387 (n_12898, n18444);
  and g28388 (n18445, n_12897, n_12898);
  and g28389 (n18446, n_11401, n18445);
  not g28390 (n_12899, n18405);
  not g28391 (n_12900, n18446);
  and g28392 (n18447, n_12899, n_12900);
  not g28393 (n_12901, n18447);
  and g28394 (n18448, pi0788, n_12901);
  and g28395 (n18449, pi0618, n18395);
  and g28396 (n18450, pi0609, n18394);
  and g28397 (n18451, n_11866, n_12854);
  and g28398 (n18452, pi0625, n18451);
  not g28399 (n_12902, n18451);
  and g28400 (n18453, n18408, n_12902);
  not g28401 (n_12903, n18452);
  not g28402 (n_12904, n18453);
  and g28403 (n18454, n_12903, n_12904);
  not g28404 (n_12905, n18454);
  and g28405 (n18455, n18390, n_12905);
  and g28406 (n18456, n_11823, n_12857);
  not g28407 (n_12906, n18455);
  and g28408 (n18457, n_12906, n18456);
  and g28409 (n18458, pi1153, n18408);
  and g28410 (n18459, n_12903, n18458);
  and g28411 (n18460, pi0608, n_12858);
  not g28412 (n_12907, n18459);
  and g28413 (n18461, n_12907, n18460);
  not g28414 (n_12908, n18457);
  not g28415 (n_12909, n18461);
  and g28416 (n18462, n_12908, n_12909);
  not g28417 (n_12910, n18462);
  and g28418 (n18463, pi0778, n_12910);
  and g28419 (n18464, n_11749, n_12904);
  not g28420 (n_12911, n18463);
  not g28421 (n_12912, n18464);
  and g28422 (n18465, n_12911, n_12912);
  not g28423 (n_12913, n18465);
  and g28424 (n18466, n_11971, n_12913);
  not g28425 (n_12914, n18450);
  and g28426 (n18467, n_11768, n_12914);
  not g28427 (n_12915, n18466);
  and g28428 (n18468, n_12915, n18467);
  and g28429 (n18469, n_11767, n_12870);
  not g28430 (n_12916, n18468);
  and g28431 (n18470, n_12916, n18469);
  and g28432 (n18471, n_11971, n18394);
  and g28433 (n18472, pi0609, n_12913);
  not g28434 (n_12917, n18471);
  and g28435 (n18473, pi1155, n_12917);
  not g28436 (n_12918, n18472);
  and g28437 (n18474, n_12918, n18473);
  and g28438 (n18475, pi0660, n_12871);
  not g28439 (n_12919, n18474);
  and g28440 (n18476, n_12919, n18475);
  not g28441 (n_12920, n18470);
  not g28442 (n_12921, n18476);
  and g28443 (n18477, n_12920, n_12921);
  not g28444 (n_12922, n18477);
  and g28445 (n18478, pi0785, n_12922);
  and g28446 (n18479, n_11964, n_12913);
  not g28447 (n_12923, n18478);
  not g28448 (n_12924, n18479);
  and g28449 (n18480, n_12923, n_12924);
  not g28450 (n_12925, n18480);
  and g28451 (n18481, n_11984, n_12925);
  not g28452 (n_12926, n18449);
  and g28453 (n18482, n_11413, n_12926);
  not g28454 (n_12927, n18481);
  and g28455 (n18483, n_12927, n18482);
  and g28456 (n18484, n_11412, n_12878);
  not g28457 (n_12928, n18483);
  and g28458 (n18485, n_12928, n18484);
  and g28459 (n18486, n_11984, n18395);
  and g28460 (n18487, pi0618, n_12925);
  not g28461 (n_12929, n18486);
  and g28462 (n18488, pi1154, n_12929);
  not g28463 (n_12930, n18487);
  and g28464 (n18489, n_12930, n18488);
  and g28465 (n18490, pi0627, n_12879);
  not g28466 (n_12931, n18489);
  and g28467 (n18491, n_12931, n18490);
  not g28468 (n_12932, n18485);
  not g28469 (n_12933, n18491);
  and g28470 (n18492, n_12932, n_12933);
  not g28471 (n_12934, n18492);
  and g28472 (n18493, pi0781, n_12934);
  and g28473 (n18494, n_11981, n_12925);
  not g28474 (n_12935, n18493);
  not g28475 (n_12936, n18494);
  and g28476 (n18495, n_12935, n_12936);
  and g28477 (n18496, n_12315, n18495);
  not g28478 (n_12937, n18495);
  and g28479 (n18497, n_11821, n_12937);
  and g28480 (n18498, pi0619, n18396);
  not g28481 (n_12938, n18498);
  and g28482 (n18499, n_11405, n_12938);
  not g28483 (n_12939, n18497);
  and g28484 (n18500, n_12939, n18499);
  and g28485 (n18501, n_11403, n_12888);
  not g28486 (n_12940, n18500);
  and g28487 (n18502, n_12940, n18501);
  and g28488 (n18503, n_11821, n18396);
  and g28489 (n18504, pi0619, n_12937);
  not g28490 (n_12941, n18503);
  and g28491 (n18505, pi1159, n_12941);
  not g28492 (n_12942, n18504);
  and g28493 (n18506, n_12942, n18505);
  and g28494 (n18507, pi0648, n_12889);
  not g28495 (n_12943, n18506);
  and g28496 (n18508, n_12943, n18507);
  not g28497 (n_12944, n18502);
  and g28498 (n18509, pi0789, n_12944);
  not g28499 (n_12945, n18508);
  and g28500 (n18510, n_12945, n18509);
  not g28501 (n_12946, n18496);
  and g28502 (n18511, n17970, n_12946);
  not g28503 (n_12947, n18510);
  and g28504 (n18512, n_12947, n18511);
  not g28505 (n_12948, n18448);
  not g28506 (n_12949, n18512);
  and g28507 (n18513, n_12948, n_12949);
  not g28508 (n_12950, n18513);
  and g28509 (n18514, n_11789, n_12950);
  not g28510 (n_12951, n18437);
  and g28511 (n18515, n_12318, n_12951);
  not g28512 (n_12952, n18445);
  and g28513 (n18516, pi0788, n_12952);
  not g28514 (n_12953, n18515);
  not g28515 (n_12954, n18516);
  and g28516 (n18517, n_12953, n_12954);
  and g28517 (n18518, pi0628, n18517);
  not g28518 (n_12955, n18518);
  and g28519 (n18519, n_11794, n_12955);
  not g28520 (n_12956, n18514);
  and g28521 (n18520, n_12956, n18519);
  not g28522 (n_12957, n18404);
  and g28523 (n18521, n_12354, n_12957);
  not g28524 (n_12958, n18520);
  and g28525 (n18522, n_12958, n18521);
  and g28526 (n18523, n_12547, n18398);
  not g28527 (n_12959, n18523);
  and g28528 (n18524, n_11794, n_12959);
  and g28529 (n18525, n_11789, n18517);
  and g28530 (n18526, pi0628, n_12950);
  not g28531 (n_12960, n18525);
  and g28532 (n18527, pi1156, n_12960);
  not g28533 (n_12961, n18526);
  and g28534 (n18528, n_12961, n18527);
  not g28535 (n_12962, n18524);
  and g28536 (n18529, pi0629, n_12962);
  not g28537 (n_12963, n18528);
  and g28538 (n18530, n_12963, n18529);
  not g28539 (n_12964, n18522);
  not g28540 (n_12965, n18530);
  and g28541 (n18531, n_12964, n_12965);
  not g28542 (n_12966, n18531);
  and g28543 (n18532, pi0792, n_12966);
  and g28544 (n18533, n_11787, n_12950);
  not g28545 (n_12967, n18532);
  not g28546 (n_12968, n18533);
  and g28547 (n18534, n_12967, n_12968);
  not g28548 (n_12969, n18534);
  and g28549 (n18535, n_11806, n_12969);
  and g28550 (n18536, n_12368, n18517);
  and g28551 (n18537, n17779, n18382);
  not g28552 (n_12970, n18536);
  not g28553 (n_12971, n18537);
  and g28554 (n18538, n_12970, n_12971);
  not g28555 (n_12972, n18538);
  and g28556 (n18539, pi0647, n_12972);
  not g28557 (n_12973, n18539);
  and g28558 (n18540, n_11810, n_12973);
  not g28559 (n_12974, n18535);
  and g28560 (n18541, n_12974, n18540);
  not g28561 (n_12975, n18402);
  and g28562 (n18542, n_12375, n_12975);
  not g28563 (n_12976, n18541);
  and g28564 (n18543, n_12976, n18542);
  and g28565 (n18544, n_11806, n18399);
  and g28566 (n18545, pi0647, n18382);
  not g28567 (n_12977, n18545);
  and g28568 (n18546, n_11810, n_12977);
  not g28569 (n_12978, n18544);
  and g28570 (n18547, n_12978, n18546);
  and g28571 (n18548, pi0647, n_12969);
  and g28572 (n18549, n_11806, n_12972);
  not g28573 (n_12979, n18549);
  and g28574 (n18550, pi1157, n_12979);
  not g28575 (n_12980, n18548);
  and g28576 (n18551, n_12980, n18550);
  not g28577 (n_12981, n18547);
  and g28578 (n18552, pi0630, n_12981);
  not g28579 (n_12982, n18551);
  and g28580 (n18553, n_12982, n18552);
  not g28581 (n_12983, n18543);
  not g28582 (n_12984, n18553);
  and g28583 (n18554, n_12983, n_12984);
  not g28584 (n_12985, n18554);
  and g28585 (n18555, pi0787, n_12985);
  and g28586 (n18556, n_11803, n_12969);
  not g28587 (n_12986, n18555);
  not g28588 (n_12987, n18556);
  and g28589 (n18557, n_12986, n_12987);
  not g28590 (n_12988, n18557);
  and g28591 (n18558, n_12411, n_12988);
  not g28592 (n_12989, n18399);
  and g28593 (n18559, n_11803, n_12989);
  and g28594 (n18560, n_12975, n_12981);
  not g28595 (n_12990, n18560);
  and g28596 (n18561, pi0787, n_12990);
  not g28597 (n_12991, n18559);
  not g28598 (n_12992, n18561);
  and g28599 (n18562, n_12991, n_12992);
  and g28600 (n18563, n_11819, n18562);
  and g28601 (n18564, pi0644, n_12988);
  not g28602 (n_12993, n18563);
  and g28603 (n18565, pi0715, n_12993);
  not g28604 (n_12994, n18564);
  and g28605 (n18566, n_12994, n18565);
  and g28606 (n18567, n17804, n_12852);
  and g28607 (n18568, n_12392, n18538);
  not g28608 (n_12995, n18567);
  not g28609 (n_12996, n18568);
  and g28610 (n18569, n_12995, n_12996);
  and g28611 (n18570, pi0644, n18569);
  and g28612 (n18571, n_11819, n18382);
  not g28613 (n_12997, n18571);
  and g28614 (n18572, n_12395, n_12997);
  not g28615 (n_12998, n18570);
  and g28616 (n18573, n_12998, n18572);
  not g28617 (n_12999, n18573);
  and g28618 (n18574, pi1160, n_12999);
  not g28619 (n_13000, n18566);
  and g28620 (n18575, n_13000, n18574);
  and g28621 (n18576, n_11819, n18569);
  and g28622 (n18577, pi0644, n18382);
  not g28623 (n_13001, n18577);
  and g28624 (n18578, pi0715, n_13001);
  not g28625 (n_13002, n18576);
  and g28626 (n18579, n_13002, n18578);
  and g28627 (n18580, pi0644, n18562);
  and g28628 (n18581, n_11819, n_12988);
  not g28629 (n_13003, n18580);
  and g28630 (n18582, n_12395, n_13003);
  not g28631 (n_13004, n18581);
  and g28632 (n18583, n_13004, n18582);
  not g28633 (n_13005, n18579);
  and g28634 (n18584, n_12405, n_13005);
  not g28635 (n_13006, n18583);
  and g28636 (n18585, n_13006, n18584);
  not g28637 (n_13007, n18575);
  not g28638 (n_13008, n18585);
  and g28639 (n18586, n_13007, n_13008);
  not g28640 (n_13009, n18586);
  and g28641 (n18587, pi0790, n_13009);
  not g28642 (n_13010, n18558);
  and g28643 (n18588, pi0832, n_13010);
  not g28644 (n_13011, n18587);
  and g28645 (n18589, n_13011, n18588);
  not g28646 (n_13012, n18381);
  not g28647 (n_13013, n18589);
  and g28648 (po0298, n_13012, n_13013);
  and g28649 (n18591, n2571, n_11742);
  not g28650 (n_13014, n18591);
  and g28651 (n18592, pi0142, n_13014);
  and g28652 (n18593, pi0039, n_11734);
  and g28653 (n18594, pi0142, n_12667);
  not g28654 (n_13015, n18593);
  and g28655 (n18595, n_13015, n18594);
  and g28656 (n18596, pi0142, n_11684);
  not g28657 (n_13016, n18596);
  and g28658 (n18597, n_3162, n_13016);
  and g28659 (n18598, pi0142, n_11694);
  not g28660 (n_13017, n18598);
  and g28661 (n18599, n6242, n_13017);
  not g28662 (n_13018, n18599);
  and g28663 (n18600, pi0215, n_13018);
  not g28664 (n_13019, n18597);
  and g28665 (n18601, n_13019, n18600);
  and g28666 (n18602, pi0142, n_11445);
  not g28667 (n_13020, n18602);
  and g28668 (n18603, n3448, n_13020);
  and g28669 (n18604, pi0142, n_11712);
  not g28670 (n_13021, n18604);
  and g28671 (n18605, n_3162, n_13021);
  and g28672 (n18606, pi0142, n_11706);
  not g28673 (n_13022, n18606);
  and g28674 (n18607, n6242, n_13022);
  not g28675 (n_13023, n18605);
  not g28676 (n_13024, n18607);
  and g28677 (n18608, n_13023, n_13024);
  not g28678 (n_13025, n18608);
  and g28679 (n18609, n_9350, n_13025);
  not g28680 (n_13026, n18603);
  and g28681 (n18610, n_36, n_13026);
  not g28682 (n_13027, n18609);
  and g28683 (n18611, n_13027, n18610);
  not g28684 (n_13028, n18601);
  not g28685 (n_13029, n18611);
  and g28686 (n18612, n_13028, n_13029);
  and g28687 (n18613, pi0039, pi0299);
  not g28688 (n_13030, n18612);
  and g28689 (n18614, n_13030, n18613);
  not g28690 (n_13031, n18595);
  not g28691 (n_13032, n18614);
  and g28692 (n18615, n_13031, n_13032);
  not g28693 (n_13033, n18615);
  and g28694 (n18616, n14873, n_13033);
  not g28695 (n_13034, n18592);
  not g28696 (n_13035, n18616);
  and g28697 (n18617, n_13034, n_13035);
  not g28698 (n_13036, n18617);
  and g28699 (n18618, n16639, n_13036);
  and g28700 (n18619, pi0142, n_11417);
  and g28701 (n18620, pi0039, pi0142);
  not g28702 (n_13037, n18620);
  and g28703 (n18621, pi0038, n_13037);
  and g28704 (n18622, pi0142, n_11432);
  and g28705 (n18623, pi0735, n16645);
  and g28706 (n18624, n2521, n18623);
  not g28707 (n_13039, n18622);
  not g28708 (n_13040, n18624);
  and g28709 (n18625, n_13039, n_13040);
  not g28710 (n_13041, n18625);
  and g28711 (n18626, n_162, n_13041);
  not g28712 (n_13042, n18626);
  and g28713 (n18627, n18621, n_13042);
  and g28714 (n18628, n_738, n_12243);
  and g28715 (n18629, pi0142, n16948);
  not g28716 (n_13043, n18628);
  and g28717 (n18630, pi0735, n_13043);
  not g28718 (n_13044, n18629);
  and g28719 (n18631, n_13044, n18630);
  not g28720 (n_13045, pi0735);
  and g28721 (n18632, pi0142, n_13045);
  and g28722 (n18633, n_11674, n18632);
  not g28723 (n_13046, n18631);
  not g28724 (n_13047, n18633);
  and g28725 (n18634, n_13046, n_13047);
  not g28726 (n_13048, n18634);
  and g28727 (n18635, n_162, n_13048);
  and g28728 (n18636, n16652, n18623);
  not g28729 (n_13049, n18636);
  and g28730 (n18637, n_13020, n_13049);
  and g28731 (n18638, n3448, n18637);
  and g28732 (n18639, n_738, n_11459);
  not g28733 (n_13050, n16791);
  and g28734 (n18640, pi0142, n_13050);
  not g28735 (n_13051, n18639);
  not g28736 (n_13052, n18640);
  and g28737 (n18641, n_13051, n_13052);
  not g28738 (n_13053, n18641);
  and g28739 (n18642, pi0735, n_13053);
  and g28740 (n18643, n_13045, n_13022);
  not g28741 (n_13054, n18642);
  not g28742 (n_13055, n18643);
  and g28743 (n18644, n_13054, n_13055);
  and g28744 (n18645, n6242, n18644);
  and g28745 (n18646, n_738, n16705);
  and g28746 (n18647, pi0142, n16763);
  not g28747 (n_13056, n18646);
  not g28748 (n_13057, n18647);
  and g28749 (n18648, n_13056, n_13057);
  not g28750 (n_13058, n18648);
  and g28751 (n18649, pi0735, n_13058);
  and g28752 (n18650, n_13045, n_13021);
  not g28753 (n_13059, n18649);
  not g28754 (n_13060, n18650);
  and g28755 (n18651, n_13059, n_13060);
  and g28756 (n18652, n_3162, n18651);
  not g28757 (n_13061, n18652);
  and g28758 (n18653, n_9350, n_13061);
  not g28759 (n_13062, n18645);
  and g28760 (n18654, n_13062, n18653);
  not g28761 (n_13063, n18638);
  and g28762 (n18655, n_36, n_13063);
  not g28763 (n_13064, n18654);
  and g28764 (n18656, n_13064, n18655);
  and g28765 (n18657, n_13045, n_13017);
  and g28766 (n18658, n_738, n17560);
  not g28767 (n_13065, n16811);
  and g28768 (n18659, pi0142, n_13065);
  not g28769 (n_13066, n18658);
  and g28770 (n18660, pi0735, n_13066);
  not g28771 (n_13067, n18659);
  and g28772 (n18661, n_13067, n18660);
  not g28773 (n_13068, n18657);
  not g28774 (n_13069, n18661);
  and g28775 (n18662, n_13068, n_13069);
  not g28776 (n_13070, n18662);
  and g28777 (n18663, n6242, n_13070);
  and g28778 (n18664, n_13045, n_13016);
  not g28779 (n_13071, n16819);
  and g28780 (n18665, pi0142, n_13071);
  and g28781 (n18666, n17559, n18658);
  not g28782 (n_13072, n18666);
  and g28783 (n18667, pi0735, n_13072);
  not g28784 (n_13073, n18665);
  and g28785 (n18668, n_13073, n18667);
  not g28786 (n_13074, n18664);
  not g28787 (n_13075, n18668);
  and g28788 (n18669, n_13074, n_13075);
  not g28789 (n_13076, n18669);
  and g28790 (n18670, n_3162, n_13076);
  not g28791 (n_13077, n18663);
  and g28792 (n18671, pi0215, n_13077);
  not g28793 (n_13078, n18670);
  and g28794 (n18672, n_13078, n18671);
  not g28795 (n_13079, n18672);
  and g28796 (n18673, pi0299, n_13079);
  not g28797 (n_13080, n18656);
  and g28798 (n18674, n_13080, n18673);
  and g28799 (n18675, n6205, n_13070);
  and g28800 (n18676, n_3119, n_13076);
  not g28801 (n_13081, n18675);
  and g28802 (n18677, pi0223, n_13081);
  not g28803 (n_13082, n18676);
  and g28804 (n18678, n_13082, n18677);
  and g28805 (n18679, n2603, n18637);
  and g28806 (n18680, n6205, n18644);
  and g28807 (n18681, n_3119, n18651);
  not g28808 (n_13083, n18681);
  and g28809 (n18682, n_9349, n_13083);
  not g28810 (n_13084, n18680);
  and g28811 (n18683, n_13084, n18682);
  not g28812 (n_13085, n18679);
  and g28813 (n18684, n_223, n_13085);
  not g28814 (n_13086, n18683);
  and g28815 (n18685, n_13086, n18684);
  not g28816 (n_13087, n18678);
  and g28817 (n18686, n_234, n_13087);
  not g28818 (n_13088, n18685);
  and g28819 (n18687, n_13088, n18686);
  not g28820 (n_13089, n18674);
  and g28821 (n18688, pi0039, n_13089);
  not g28822 (n_13090, n18687);
  and g28823 (n18689, n_13090, n18688);
  not g28824 (n_13091, n18635);
  and g28825 (n18690, n_161, n_13091);
  not g28826 (n_13092, n18689);
  and g28827 (n18691, n_13092, n18690);
  not g28828 (n_13093, n18627);
  and g28829 (n18692, n2571, n_13093);
  not g28830 (n_13094, n18691);
  and g28831 (n18693, n_13094, n18692);
  not g28832 (n_13095, n18619);
  not g28833 (n_13096, n18693);
  and g28834 (n18694, n_13095, n_13096);
  not g28835 (n_13097, n18694);
  and g28836 (n18695, n_11749, n_13097);
  and g28837 (n18696, n_11753, n18694);
  and g28838 (n18697, pi0625, n18617);
  not g28839 (n_13098, n18697);
  and g28840 (n18698, n_11757, n_13098);
  not g28841 (n_13099, n18696);
  and g28842 (n18699, n_13099, n18698);
  and g28843 (n18700, n_11753, n18617);
  and g28844 (n18701, pi0625, n18694);
  not g28845 (n_13100, n18700);
  and g28846 (n18702, pi1153, n_13100);
  not g28847 (n_13101, n18701);
  and g28848 (n18703, n_13101, n18702);
  not g28849 (n_13102, n18699);
  not g28850 (n_13103, n18703);
  and g28851 (n18704, n_13102, n_13103);
  not g28852 (n_13104, n18704);
  and g28853 (n18705, pi0778, n_13104);
  not g28854 (n_13105, n18695);
  not g28855 (n_13106, n18705);
  and g28856 (n18706, n_13105, n_13106);
  and g28857 (n18707, n_11773, n18706);
  and g28858 (n18708, n17075, n18617);
  not g28859 (n_13107, n18707);
  not g28860 (n_13108, n18708);
  and g28861 (n18709, n_13107, n_13108);
  and g28862 (n18710, n_11777, n18709);
  not g28863 (n_13109, n18618);
  not g28864 (n_13110, n18710);
  and g28865 (n18711, n_13109, n_13110);
  and g28866 (n18712, n_11780, n18711);
  and g28867 (n18713, n16635, n18617);
  not g28868 (n_13111, n18712);
  not g28869 (n_13112, n18713);
  and g28870 (n18714, n_13111, n_13112);
  not g28871 (n_13113, n18714);
  and g28872 (n18715, n_11783, n_13113);
  and g28873 (n18716, n16631, n18617);
  not g28874 (n_13114, n18715);
  not g28875 (n_13115, n18716);
  and g28876 (n18717, n_13114, n_13115);
  and g28877 (n18718, n_11787, n18717);
  and g28878 (n18719, n_11789, n18617);
  not g28879 (n_13116, n18717);
  and g28880 (n18720, pi0628, n_13116);
  not g28881 (n_13117, n18719);
  and g28882 (n18721, pi1156, n_13117);
  not g28883 (n_13118, n18720);
  and g28884 (n18722, n_13118, n18721);
  and g28885 (n18723, pi0628, n18617);
  and g28886 (n18724, n_11789, n_13116);
  not g28887 (n_13119, n18723);
  and g28888 (n18725, n_11794, n_13119);
  not g28889 (n_13120, n18724);
  and g28890 (n18726, n_13120, n18725);
  not g28891 (n_13121, n18722);
  not g28892 (n_13122, n18726);
  and g28893 (n18727, n_13121, n_13122);
  not g28894 (n_13123, n18727);
  and g28895 (n18728, pi0792, n_13123);
  not g28896 (n_13124, n18718);
  not g28897 (n_13125, n18728);
  and g28898 (n18729, n_13124, n_13125);
  not g28899 (n_13126, n18729);
  and g28900 (n18730, n_11803, n_13126);
  and g28901 (n18731, n_11806, n18617);
  and g28902 (n18732, pi0647, n18729);
  not g28903 (n_13127, n18731);
  and g28904 (n18733, pi1157, n_13127);
  not g28905 (n_13128, n18732);
  and g28906 (n18734, n_13128, n18733);
  and g28907 (n18735, n_11806, n18729);
  and g28908 (n18736, pi0647, n18617);
  not g28909 (n_13129, n18736);
  and g28910 (n18737, n_11810, n_13129);
  not g28911 (n_13130, n18735);
  and g28912 (n18738, n_13130, n18737);
  not g28913 (n_13131, n18734);
  not g28914 (n_13132, n18738);
  and g28915 (n18739, n_13131, n_13132);
  not g28916 (n_13133, n18739);
  and g28917 (n18740, pi0787, n_13133);
  not g28918 (n_13134, n18730);
  not g28919 (n_13135, n18740);
  and g28920 (n18741, n_13134, n_13135);
  and g28921 (n18742, n_11819, n18741);
  and g28922 (n18743, n_11984, n18617);
  and g28923 (n18744, pi0743, n17244);
  and g28924 (n18745, n2521, n18744);
  not g28925 (n_13137, n18745);
  and g28926 (n18746, n_13039, n_13137);
  not g28927 (n_13138, n18746);
  and g28928 (n18747, n_162, n_13138);
  not g28929 (n_13139, n18747);
  and g28930 (n18748, n18621, n_13139);
  not g28931 (n_13140, pi0743);
  and g28932 (n18749, pi0142, n_13140);
  and g28933 (n18750, n_11671, n18749);
  and g28934 (n18751, n_738, n_11915);
  not g28935 (n_13141, n17137);
  and g28936 (n18752, pi0142, n_13141);
  not g28937 (n_13142, n18751);
  and g28938 (n18753, pi0743, n_13142);
  not g28939 (n_13143, n18752);
  and g28940 (n18754, n_13143, n18753);
  not g28941 (n_13144, n18750);
  and g28942 (n18755, n_234, n_13144);
  not g28943 (n_13145, n18754);
  and g28944 (n18756, n_13145, n18755);
  and g28945 (n18757, n_738, n_11920);
  and g28946 (n18758, pi0142, n_11670);
  not g28947 (n_13146, n18758);
  and g28948 (n18759, n_13140, n_13146);
  and g28949 (n18760, pi0142, n17124);
  not g28950 (n_13147, n18757);
  not g28951 (n_13148, n18759);
  and g28952 (n18761, n_13147, n_13148);
  not g28953 (n_13149, n18760);
  and g28954 (n18762, n_13149, n18761);
  not g28955 (n_13150, n18762);
  and g28956 (n18763, pi0299, n_13150);
  not g28957 (n_13151, n18756);
  not g28958 (n_13152, n18763);
  and g28959 (n18764, n_13151, n_13152);
  and g28960 (n18765, n_162, n18764);
  and g28961 (n18766, n_13140, n_13016);
  and g28962 (n18767, pi0142, n_11883);
  and g28963 (n18768, pi0743, n17558);
  not g28964 (n_13153, n18767);
  and g28965 (n18769, n_13153, n18768);
  not g28966 (n_13154, n18766);
  not g28967 (n_13155, n18769);
  and g28968 (n18770, n_13154, n_13155);
  not g28969 (n_13156, n18770);
  and g28970 (n18771, n_3119, n_13156);
  and g28971 (n18772, n_13140, n_13017);
  and g28972 (n18773, pi0142, n17200);
  and g28973 (n18774, pi0743, n17241);
  not g28974 (n_13157, n18773);
  and g28975 (n18775, n_13157, n18774);
  not g28976 (n_13158, n18772);
  not g28977 (n_13159, n18775);
  and g28978 (n18776, n_13158, n_13159);
  not g28979 (n_13160, n18776);
  and g28980 (n18777, n6205, n_13160);
  not g28981 (n_13161, n18777);
  and g28982 (n18778, pi0223, n_13161);
  not g28983 (n_13162, n18771);
  and g28984 (n18779, n_13162, n18778);
  and g28985 (n18780, n_13140, n_13021);
  and g28986 (n18781, pi0142, n_11858);
  and g28987 (n18782, pi0743, n_11934);
  not g28988 (n_13163, n18781);
  and g28989 (n18783, n_13163, n18782);
  not g28990 (n_13164, n18780);
  not g28991 (n_13165, n18783);
  and g28992 (n18784, n_13164, n_13165);
  and g28993 (n18785, n_3119, n18784);
  and g28994 (n18786, n_738, n17252);
  and g28995 (n18787, pi0142, n17175);
  not g28996 (n_13166, n18786);
  not g28997 (n_13167, n18787);
  and g28998 (n18788, n_13166, n_13167);
  not g28999 (n_13168, n18788);
  and g29000 (n18789, pi0743, n_13168);
  and g29001 (n18790, n_13140, n_13022);
  not g29002 (n_13169, n18789);
  not g29003 (n_13170, n18790);
  and g29004 (n18791, n_13169, n_13170);
  and g29005 (n18792, n6205, n18791);
  not g29006 (n_13171, n18785);
  and g29007 (n18793, n_9349, n_13171);
  not g29008 (n_13172, n18792);
  and g29009 (n18794, n_13172, n18793);
  and g29010 (n18795, pi0743, n17235);
  not g29011 (n_13173, n18795);
  and g29012 (n18796, n_13020, n_13173);
  and g29013 (n18797, n2603, n18796);
  not g29014 (n_13174, n18797);
  and g29015 (n18798, n_223, n_13174);
  not g29016 (n_13175, n18794);
  and g29017 (n18799, n_13175, n18798);
  not g29018 (n_13176, n18779);
  and g29019 (n18800, n_234, n_13176);
  not g29020 (n_13177, n18799);
  and g29021 (n18801, n_13177, n18800);
  not g29022 (n_13178, n18796);
  and g29023 (n18802, n3448, n_13178);
  and g29024 (n18803, n_3162, n18784);
  and g29025 (n18804, n6242, n18791);
  not g29026 (n_13179, n18803);
  not g29027 (n_13180, n18804);
  and g29028 (n18805, n_13179, n_13180);
  not g29029 (n_13181, n18805);
  and g29030 (n18806, n_9350, n_13181);
  not g29031 (n_13182, n18802);
  and g29032 (n18807, n_36, n_13182);
  not g29033 (n_13183, n18806);
  and g29034 (n18808, n_13183, n18807);
  and g29035 (n18809, n_3162, n18770);
  and g29036 (n18810, n6242, n18776);
  not g29037 (n_13184, n18810);
  and g29038 (n18811, pi0215, n_13184);
  not g29039 (n_13185, n18809);
  and g29040 (n18812, n_13185, n18811);
  not g29041 (n_13186, n18808);
  not g29042 (n_13187, n18812);
  and g29043 (n18813, n_13186, n_13187);
  not g29044 (n_13188, n18813);
  and g29045 (n18814, pi0299, n_13188);
  not g29046 (n_13189, n18801);
  and g29047 (n18815, pi0039, n_13189);
  not g29048 (n_13190, n18814);
  and g29049 (n18816, n_13190, n18815);
  not g29050 (n_13191, n18765);
  and g29051 (n18817, n_161, n_13191);
  not g29052 (n_13192, n18816);
  and g29053 (n18818, n_13192, n18817);
  not g29054 (n_13193, n18748);
  and g29055 (n18819, n2571, n_13193);
  not g29056 (n_13194, n18818);
  and g29057 (n18820, n_13194, n18819);
  not g29058 (n_13195, n18820);
  and g29059 (n18821, n_13095, n_13195);
  not g29060 (n_13196, n18821);
  and g29061 (n18822, n_11960, n_13196);
  and g29062 (n18823, n17117, n_13036);
  not g29063 (n_13197, n18822);
  not g29064 (n_13198, n18823);
  and g29065 (n18824, n_13197, n_13198);
  not g29066 (n_13199, n18824);
  and g29067 (n18825, n_11964, n_13199);
  and g29068 (n18826, n_11967, n_13036);
  and g29069 (n18827, pi0609, n18822);
  not g29070 (n_13200, n18826);
  not g29071 (n_13201, n18827);
  and g29072 (n18828, n_13200, n_13201);
  not g29073 (n_13202, n18828);
  and g29074 (n18829, pi1155, n_13202);
  and g29075 (n18830, n_11972, n_13036);
  and g29076 (n18831, n_11971, n18822);
  not g29077 (n_13203, n18830);
  not g29078 (n_13204, n18831);
  and g29079 (n18832, n_13203, n_13204);
  not g29080 (n_13205, n18832);
  and g29081 (n18833, n_11768, n_13205);
  not g29082 (n_13206, n18829);
  not g29083 (n_13207, n18833);
  and g29084 (n18834, n_13206, n_13207);
  not g29085 (n_13208, n18834);
  and g29086 (n18835, pi0785, n_13208);
  not g29087 (n_13209, n18825);
  not g29088 (n_13210, n18835);
  and g29089 (n18836, n_13209, n_13210);
  and g29090 (n18837, pi0618, n18836);
  not g29091 (n_13211, n18743);
  and g29092 (n18838, pi1154, n_13211);
  not g29093 (n_13212, n18837);
  and g29094 (n18839, n_13212, n18838);
  and g29095 (n18840, pi0609, n18706);
  and g29096 (n18841, n_11753, n18821);
  and g29097 (n18842, n_13045, n18764);
  and g29098 (n18843, n16937, n18752);
  and g29099 (n18844, n_11636, n18751);
  not g29100 (n_13213, n18843);
  not g29101 (n_13214, n18844);
  and g29102 (n18845, n_13213, n_13214);
  not g29103 (n_13215, n18845);
  and g29104 (n18846, pi0743, n_13215);
  and g29105 (n18847, pi0142, n_11650);
  and g29106 (n18848, n_11915, n18847);
  and g29107 (n18849, n_738, n17618);
  not g29108 (n_13216, n18848);
  and g29109 (n18850, n_13140, n_13216);
  not g29110 (n_13217, n18849);
  and g29111 (n18851, n_13217, n18850);
  not g29112 (n_13218, n18851);
  and g29113 (n18852, n_234, n_13218);
  not g29114 (n_13219, n18846);
  and g29115 (n18853, n_13219, n18852);
  and g29116 (n18854, n_11639, n18757);
  and g29117 (n18855, n_11656, n18760);
  not g29118 (n_13220, n18854);
  not g29119 (n_13221, n18855);
  and g29120 (n18856, n_13220, n_13221);
  not g29121 (n_13222, n18856);
  and g29122 (n18857, pi0743, n_13222);
  and g29123 (n18858, n_738, n17623);
  and g29124 (n18859, pi0142, n_11657);
  and g29125 (n18860, n_11920, n18859);
  not g29126 (n_13223, n18860);
  and g29127 (n18861, n_13140, n_13223);
  not g29128 (n_13224, n18858);
  and g29129 (n18862, n_13224, n18861);
  not g29130 (n_13225, n18857);
  and g29131 (n18863, pi0299, n_13225);
  not g29132 (n_13226, n18862);
  and g29133 (n18864, n_13226, n18863);
  not g29134 (n_13227, n18853);
  not g29135 (n_13228, n18864);
  and g29136 (n18865, n_13227, n_13228);
  not g29137 (n_13229, n18865);
  and g29138 (n18866, pi0735, n_13229);
  not g29139 (n_13230, n18842);
  and g29140 (n18867, n_162, n_13230);
  not g29141 (n_13231, n18866);
  and g29142 (n18868, n_13231, n18867);
  and g29143 (n18869, n_738, n_12188);
  and g29144 (n18870, pi0142, n_12155);
  not g29145 (n_13232, n18869);
  and g29146 (n18871, pi0743, n_13232);
  not g29147 (n_13233, n18870);
  and g29148 (n18872, n_13233, n18871);
  and g29149 (n18873, n_738, n17448);
  and g29150 (n18874, pi0142, n17351);
  not g29151 (n_13234, n18873);
  and g29152 (n18875, n_13140, n_13234);
  not g29153 (n_13235, n18874);
  and g29154 (n18876, n_13235, n18875);
  not g29155 (n_13236, n18872);
  not g29156 (n_13237, n18876);
  and g29157 (n18877, n_13236, n_13237);
  not g29158 (n_13238, n18877);
  and g29159 (n18878, pi0735, n_13238);
  and g29160 (n18879, n_13045, n18776);
  not g29161 (n_13239, n18878);
  not g29162 (n_13240, n18879);
  and g29163 (n18880, n_13239, n_13240);
  and g29164 (n18881, n6205, n18880);
  and g29165 (n18882, n_738, n17562);
  and g29166 (n18883, pi0142, n17527);
  not g29167 (n_13241, n18882);
  and g29168 (n18884, pi0743, n_13241);
  not g29169 (n_13242, n18883);
  and g29170 (n18885, n_13242, n18884);
  and g29171 (n18886, n_738, n_12128);
  and g29172 (n18887, pi0142, n17333);
  not g29173 (n_13243, n18887);
  and g29174 (n18888, n_13140, n_13243);
  not g29175 (n_13244, n18886);
  and g29176 (n18889, n_13244, n18888);
  not g29177 (n_13245, n18885);
  not g29178 (n_13246, n18889);
  and g29179 (n18890, n_13245, n_13246);
  not g29180 (n_13247, n18890);
  and g29181 (n18891, pi0735, n_13247);
  and g29182 (n18892, n_13045, n18770);
  not g29183 (n_13248, n18891);
  not g29184 (n_13249, n18892);
  and g29185 (n18893, n_13248, n_13249);
  and g29186 (n18894, n_3119, n18893);
  not g29187 (n_13250, n18881);
  and g29188 (n18895, pi0223, n_13250);
  not g29189 (n_13251, n18894);
  and g29190 (n18896, n_13251, n18895);
  and g29191 (n18897, n_13045, n18796);
  and g29192 (n18898, n_12254, n18746);
  not g29193 (n_13252, n18898);
  and g29194 (n18899, n_11425, n_13252);
  not g29195 (n_13253, n18899);
  and g29196 (n18900, pi0735, n_13253);
  and g29197 (n18901, n_13020, n18900);
  not g29198 (n_13254, n18897);
  not g29199 (n_13255, n18901);
  and g29200 (n18902, n_13254, n_13255);
  not g29201 (n_13256, n18902);
  and g29202 (n18903, n2603, n_13256);
  and g29203 (n18904, pi0142, n17510);
  not g29204 (n_13257, n17573);
  and g29205 (n18905, n_738, n_13257);
  not g29206 (n_13258, n18904);
  and g29207 (n18906, pi0743, n_13258);
  not g29208 (n_13259, n18905);
  and g29209 (n18907, n_13259, n18906);
  and g29210 (n18908, n_738, n17420);
  and g29211 (n18909, pi0142, n17373);
  not g29212 (n_13260, n18908);
  and g29213 (n18910, n_13140, n_13260);
  not g29214 (n_13261, n18909);
  and g29215 (n18911, n_13261, n18910);
  not g29216 (n_13262, n18907);
  not g29217 (n_13263, n18911);
  and g29218 (n18912, n_13262, n_13263);
  not g29219 (n_13264, n18912);
  and g29220 (n18913, pi0735, n_13264);
  and g29221 (n18914, n_13045, n18791);
  not g29222 (n_13265, n18913);
  not g29223 (n_13266, n18914);
  and g29224 (n18915, n_13265, n_13266);
  not g29225 (n_13267, n18915);
  and g29226 (n18916, n6205, n_13267);
  not g29227 (n_13268, n17584);
  and g29228 (n18917, n_738, n_13268);
  and g29229 (n18918, pi0142, n17499);
  not g29230 (n_13269, n18918);
  and g29231 (n18919, pi0743, n_13269);
  not g29232 (n_13270, n18917);
  and g29233 (n18920, n_13270, n18919);
  and g29234 (n18921, n_738, n_12093);
  and g29235 (n18922, pi0142, n17383);
  not g29236 (n_13271, n18922);
  and g29237 (n18923, n_13140, n_13271);
  not g29238 (n_13272, n18921);
  and g29239 (n18924, n_13272, n18923);
  not g29240 (n_13273, n18920);
  not g29241 (n_13274, n18924);
  and g29242 (n18925, n_13273, n_13274);
  not g29243 (n_13275, n18925);
  and g29244 (n18926, pi0735, n_13275);
  and g29245 (n18927, n_13045, n18784);
  not g29246 (n_13276, n18926);
  not g29247 (n_13277, n18927);
  and g29248 (n18928, n_13276, n_13277);
  not g29249 (n_13278, n18928);
  and g29250 (n18929, n_3119, n_13278);
  not g29251 (n_13279, n18929);
  and g29252 (n18930, n_9349, n_13279);
  not g29253 (n_13280, n18916);
  and g29254 (n18931, n_13280, n18930);
  not g29255 (n_13281, n18903);
  and g29256 (n18932, n_223, n_13281);
  not g29257 (n_13282, n18931);
  and g29258 (n18933, n_13282, n18932);
  not g29259 (n_13283, n18896);
  not g29260 (n_13284, n18933);
  and g29261 (n18934, n_13283, n_13284);
  not g29262 (n_13285, n18934);
  and g29263 (n18935, n_234, n_13285);
  and g29264 (n18936, n6242, n18880);
  and g29265 (n18937, n_3162, n18893);
  not g29266 (n_13286, n18936);
  and g29267 (n18938, pi0215, n_13286);
  not g29268 (n_13287, n18937);
  and g29269 (n18939, n_13287, n18938);
  and g29270 (n18940, n3448, n_13256);
  and g29271 (n18941, n_3162, n_13278);
  and g29272 (n18942, n6242, n_13267);
  not g29273 (n_13288, n18941);
  and g29274 (n18943, n_9350, n_13288);
  not g29275 (n_13289, n18942);
  and g29276 (n18944, n_13289, n18943);
  not g29277 (n_13290, n18940);
  and g29278 (n18945, n_36, n_13290);
  not g29279 (n_13291, n18944);
  and g29280 (n18946, n_13291, n18945);
  not g29281 (n_13292, n18939);
  not g29282 (n_13293, n18946);
  and g29283 (n18947, n_13292, n_13293);
  not g29284 (n_13294, n18947);
  and g29285 (n18948, pi0299, n_13294);
  not g29286 (n_13295, n18935);
  and g29287 (n18949, pi0039, n_13295);
  not g29288 (n_13296, n18948);
  and g29289 (n18950, n_13296, n18949);
  not g29290 (n_13297, n18868);
  not g29291 (n_13298, n18950);
  and g29292 (n18951, n_13297, n_13298);
  not g29293 (n_13299, n18951);
  and g29294 (n18952, n_161, n_13299);
  and g29295 (n18953, pi0735, n17645);
  not g29296 (n_13300, n18953);
  and g29297 (n18954, n18746, n_13300);
  not g29298 (n_13301, n18954);
  and g29299 (n18955, n_162, n_13301);
  not g29300 (n_13302, n18955);
  and g29301 (n18956, n18621, n_13302);
  not g29302 (n_13303, n18956);
  and g29303 (n18957, n2571, n_13303);
  not g29304 (n_13304, n18952);
  and g29305 (n18958, n_13304, n18957);
  not g29306 (n_13305, n18958);
  and g29307 (n18959, n_13095, n_13305);
  and g29308 (n18960, pi0625, n18959);
  not g29309 (n_13306, n18841);
  and g29310 (n18961, pi1153, n_13306);
  not g29311 (n_13307, n18960);
  and g29312 (n18962, n_13307, n18961);
  and g29313 (n18963, pi0608, n_13102);
  not g29314 (n_13308, n18962);
  and g29315 (n18964, n_13308, n18963);
  and g29316 (n18965, n_11753, n18959);
  and g29317 (n18966, pi0625, n18821);
  not g29318 (n_13309, n18966);
  and g29319 (n18967, n_11757, n_13309);
  not g29320 (n_13310, n18965);
  and g29321 (n18968, n_13310, n18967);
  and g29322 (n18969, n_11823, n_13103);
  not g29323 (n_13311, n18968);
  and g29324 (n18970, n_13311, n18969);
  not g29325 (n_13312, n18964);
  not g29326 (n_13313, n18970);
  and g29327 (n18971, n_13312, n_13313);
  not g29328 (n_13314, n18971);
  and g29329 (n18972, pi0778, n_13314);
  and g29330 (n18973, n_11749, n18959);
  not g29331 (n_13315, n18972);
  not g29332 (n_13316, n18973);
  and g29333 (n18974, n_13315, n_13316);
  not g29334 (n_13317, n18974);
  and g29335 (n18975, n_11971, n_13317);
  not g29336 (n_13318, n18840);
  and g29337 (n18976, n_11768, n_13318);
  not g29338 (n_13319, n18975);
  and g29339 (n18977, n_13319, n18976);
  and g29340 (n18978, n_11767, n_13206);
  not g29341 (n_13320, n18977);
  and g29342 (n18979, n_13320, n18978);
  and g29343 (n18980, n_11971, n18706);
  and g29344 (n18981, pi0609, n_13317);
  not g29345 (n_13321, n18980);
  and g29346 (n18982, pi1155, n_13321);
  not g29347 (n_13322, n18981);
  and g29348 (n18983, n_13322, n18982);
  and g29349 (n18984, pi0660, n_13207);
  not g29350 (n_13323, n18983);
  and g29351 (n18985, n_13323, n18984);
  not g29352 (n_13324, n18979);
  not g29353 (n_13325, n18985);
  and g29354 (n18986, n_13324, n_13325);
  not g29355 (n_13326, n18986);
  and g29356 (n18987, pi0785, n_13326);
  and g29357 (n18988, n_11964, n_13317);
  not g29358 (n_13327, n18987);
  not g29359 (n_13328, n18988);
  and g29360 (n18989, n_13327, n_13328);
  not g29361 (n_13329, n18989);
  and g29362 (n18990, n_11984, n_13329);
  not g29363 (n_13330, n18709);
  and g29364 (n18991, pi0618, n_13330);
  not g29365 (n_13331, n18991);
  and g29366 (n18992, n_11413, n_13331);
  not g29367 (n_13332, n18990);
  and g29368 (n18993, n_13332, n18992);
  not g29369 (n_13333, n18839);
  and g29370 (n18994, n_11412, n_13333);
  not g29371 (n_13334, n18993);
  and g29372 (n18995, n_13334, n18994);
  and g29373 (n18996, n_11984, n18836);
  and g29374 (n18997, pi0618, n18617);
  not g29375 (n_13335, n18997);
  and g29376 (n18998, n_11413, n_13335);
  not g29377 (n_13336, n18996);
  and g29378 (n18999, n_13336, n18998);
  and g29379 (n19000, pi0618, n_13329);
  and g29380 (n19001, n_11984, n_13330);
  not g29381 (n_13337, n19001);
  and g29382 (n19002, pi1154, n_13337);
  not g29383 (n_13338, n19000);
  and g29384 (n19003, n_13338, n19002);
  not g29385 (n_13339, n18999);
  and g29386 (n19004, pi0627, n_13339);
  not g29387 (n_13340, n19003);
  and g29388 (n19005, n_13340, n19004);
  not g29389 (n_13341, n18995);
  not g29390 (n_13342, n19005);
  and g29391 (n19006, n_13341, n_13342);
  not g29392 (n_13343, n19006);
  and g29393 (n19007, pi0781, n_13343);
  and g29394 (n19008, n_11981, n_13329);
  not g29395 (n_13344, n19007);
  not g29396 (n_13345, n19008);
  and g29397 (n19009, n_13344, n_13345);
  not g29398 (n_13346, n19009);
  and g29399 (n19010, n_11821, n_13346);
  and g29400 (n19011, pi0619, n18711);
  not g29401 (n_13347, n19011);
  and g29402 (n19012, n_11405, n_13347);
  not g29403 (n_13348, n19010);
  and g29404 (n19013, n_13348, n19012);
  and g29405 (n19014, n_11821, n18617);
  not g29406 (n_13349, n18836);
  and g29407 (n19015, n_11981, n_13349);
  and g29408 (n19016, n_13333, n_13339);
  not g29409 (n_13350, n19016);
  and g29410 (n19017, pi0781, n_13350);
  not g29411 (n_13351, n19015);
  not g29412 (n_13352, n19017);
  and g29413 (n19018, n_13351, n_13352);
  and g29414 (n19019, pi0619, n19018);
  not g29415 (n_13353, n19014);
  and g29416 (n19020, pi1159, n_13353);
  not g29417 (n_13354, n19019);
  and g29418 (n19021, n_13354, n19020);
  not g29419 (n_13355, n19021);
  and g29420 (n19022, n_11403, n_13355);
  not g29421 (n_13356, n19013);
  and g29422 (n19023, n_13356, n19022);
  and g29423 (n19024, pi0619, n_13346);
  and g29424 (n19025, n_11821, n18711);
  not g29425 (n_13357, n19025);
  and g29426 (n19026, pi1159, n_13357);
  not g29427 (n_13358, n19024);
  and g29428 (n19027, n_13358, n19026);
  and g29429 (n19028, n_11821, n19018);
  and g29430 (n19029, pi0619, n18617);
  not g29431 (n_13359, n19029);
  and g29432 (n19030, n_11405, n_13359);
  not g29433 (n_13360, n19028);
  and g29434 (n19031, n_13360, n19030);
  not g29435 (n_13361, n19031);
  and g29436 (n19032, pi0648, n_13361);
  not g29437 (n_13362, n19027);
  and g29438 (n19033, n_13362, n19032);
  not g29439 (n_13363, n19023);
  not g29440 (n_13364, n19033);
  and g29441 (n19034, n_13363, n_13364);
  not g29442 (n_13365, n19034);
  and g29443 (n19035, pi0789, n_13365);
  and g29444 (n19036, n_12315, n_13346);
  not g29445 (n_13366, n19035);
  not g29446 (n_13367, n19036);
  and g29447 (n19037, n_13366, n_13367);
  and g29448 (n19038, n_12318, n19037);
  and g29449 (n19039, n_12320, n19037);
  and g29450 (n19040, pi0626, n18714);
  not g29451 (n_13368, n19040);
  and g29452 (n19041, n_11395, n_13368);
  not g29453 (n_13369, n19039);
  and g29454 (n19042, n_13369, n19041);
  not g29455 (n_13370, n19018);
  and g29456 (n19043, n_12315, n_13370);
  and g29457 (n19044, n_13355, n_13361);
  not g29458 (n_13371, n19044);
  and g29459 (n19045, pi0789, n_13371);
  not g29460 (n_13372, n19043);
  not g29461 (n_13373, n19045);
  and g29462 (n19046, n_13372, n_13373);
  and g29463 (n19047, n_12320, n19046);
  and g29464 (n19048, pi0626, n18617);
  not g29465 (n_13374, n19048);
  and g29466 (n19049, n_11397, n_13374);
  not g29467 (n_13375, n19047);
  and g29468 (n19050, n_13375, n19049);
  not g29469 (n_13376, n19050);
  and g29470 (n19051, n_12330, n_13376);
  not g29471 (n_13377, n19042);
  not g29472 (n_13378, n19051);
  and g29473 (n19052, n_13377, n_13378);
  and g29474 (n19053, pi0626, n19037);
  and g29475 (n19054, n_12320, n18714);
  not g29476 (n_13379, n19054);
  and g29477 (n19055, pi0641, n_13379);
  not g29478 (n_13380, n19053);
  and g29479 (n19056, n_13380, n19055);
  and g29480 (n19057, n_12320, n18617);
  and g29481 (n19058, pi0626, n19046);
  not g29482 (n_13381, n19057);
  and g29483 (n19059, pi1158, n_13381);
  not g29484 (n_13382, n19058);
  and g29485 (n19060, n_13382, n19059);
  not g29486 (n_13383, n19060);
  and g29487 (n19061, n_12338, n_13383);
  not g29488 (n_13384, n19056);
  not g29489 (n_13385, n19061);
  and g29490 (n19062, n_13384, n_13385);
  not g29491 (n_13386, n19052);
  not g29492 (n_13387, n19062);
  and g29493 (n19063, n_13386, n_13387);
  not g29494 (n_13388, n19063);
  and g29495 (n19064, pi0788, n_13388);
  not g29496 (n_13389, n19038);
  not g29497 (n_13390, n19064);
  and g29498 (n19065, n_13389, n_13390);
  and g29499 (n19066, n_11789, n19065);
  and g29500 (n19067, n_13376, n_13383);
  not g29501 (n_13391, n19067);
  and g29502 (n19068, pi0788, n_13391);
  not g29503 (n_13392, n19046);
  and g29504 (n19069, n_12318, n_13392);
  not g29505 (n_13393, n19068);
  not g29506 (n_13394, n19069);
  and g29507 (n19070, n_13393, n_13394);
  and g29508 (n19071, pi0628, n19070);
  not g29509 (n_13395, n19071);
  and g29510 (n19072, n_11794, n_13395);
  not g29511 (n_13396, n19066);
  and g29512 (n19073, n_13396, n19072);
  and g29513 (n19074, n_12354, n_13121);
  not g29514 (n_13397, n19073);
  and g29515 (n19075, n_13397, n19074);
  and g29516 (n19076, pi0628, n19065);
  and g29517 (n19077, n_11789, n19070);
  not g29518 (n_13398, n19077);
  and g29519 (n19078, pi1156, n_13398);
  not g29520 (n_13399, n19076);
  and g29521 (n19079, n_13399, n19078);
  and g29522 (n19080, pi0629, n_13122);
  not g29523 (n_13400, n19079);
  and g29524 (n19081, n_13400, n19080);
  not g29525 (n_13401, n19075);
  not g29526 (n_13402, n19081);
  and g29527 (n19082, n_13401, n_13402);
  not g29528 (n_13403, n19082);
  and g29529 (n19083, pi0792, n_13403);
  and g29530 (n19084, n_11787, n19065);
  not g29531 (n_13404, n19083);
  not g29532 (n_13405, n19084);
  and g29533 (n19085, n_13404, n_13405);
  not g29534 (n_13406, n19085);
  and g29535 (n19086, n_11806, n_13406);
  and g29536 (n19087, n_12368, n19070);
  and g29537 (n19088, n17779, n18617);
  not g29538 (n_13407, n19087);
  not g29539 (n_13408, n19088);
  and g29540 (n19089, n_13407, n_13408);
  not g29541 (n_13409, n19089);
  and g29542 (n19090, pi0647, n_13409);
  not g29543 (n_13410, n19090);
  and g29544 (n19091, n_11810, n_13410);
  not g29545 (n_13411, n19086);
  and g29546 (n19092, n_13411, n19091);
  and g29547 (n19093, n_12375, n_13131);
  not g29548 (n_13412, n19092);
  and g29549 (n19094, n_13412, n19093);
  and g29550 (n19095, pi0647, n_13406);
  and g29551 (n19096, n_11806, n_13409);
  not g29552 (n_13413, n19096);
  and g29553 (n19097, pi1157, n_13413);
  not g29554 (n_13414, n19095);
  and g29555 (n19098, n_13414, n19097);
  and g29556 (n19099, pi0630, n_13132);
  not g29557 (n_13415, n19098);
  and g29558 (n19100, n_13415, n19099);
  not g29559 (n_13416, n19094);
  not g29560 (n_13417, n19100);
  and g29561 (n19101, n_13416, n_13417);
  not g29562 (n_13418, n19101);
  and g29563 (n19102, pi0787, n_13418);
  and g29564 (n19103, n_11803, n_13406);
  not g29565 (n_13419, n19102);
  not g29566 (n_13420, n19103);
  and g29567 (n19104, n_13419, n_13420);
  not g29568 (n_13421, n19104);
  and g29569 (n19105, pi0644, n_13421);
  not g29570 (n_13422, n18742);
  and g29571 (n19106, pi0715, n_13422);
  not g29572 (n_13423, n19105);
  and g29573 (n19107, n_13423, n19106);
  and g29574 (n19108, n17804, n_13036);
  and g29575 (n19109, n_12392, n19089);
  not g29576 (n_13424, n19108);
  not g29577 (n_13425, n19109);
  and g29578 (n19110, n_13424, n_13425);
  and g29579 (n19111, pi0644, n19110);
  and g29580 (n19112, n_11819, n18617);
  not g29581 (n_13426, n19112);
  and g29582 (n19113, n_12395, n_13426);
  not g29583 (n_13427, n19111);
  and g29584 (n19114, n_13427, n19113);
  not g29585 (n_13428, n19114);
  and g29586 (n19115, pi1160, n_13428);
  not g29587 (n_13429, n19107);
  and g29588 (n19116, n_13429, n19115);
  and g29589 (n19117, n_11819, n_13421);
  and g29590 (n19118, pi0644, n18741);
  not g29591 (n_13430, n19118);
  and g29592 (n19119, n_12395, n_13430);
  not g29593 (n_13431, n19117);
  and g29594 (n19120, n_13431, n19119);
  and g29595 (n19121, n_11819, n19110);
  and g29596 (n19122, pi0644, n18617);
  not g29597 (n_13432, n19122);
  and g29598 (n19123, pi0715, n_13432);
  not g29599 (n_13433, n19121);
  and g29600 (n19124, n_13433, n19123);
  not g29601 (n_13434, n19124);
  and g29602 (n19125, n_12405, n_13434);
  not g29603 (n_13435, n19120);
  and g29604 (n19126, n_13435, n19125);
  not g29605 (n_13436, n19116);
  and g29606 (n19127, pi0790, n_13436);
  not g29607 (n_13437, n19126);
  and g29608 (n19128, n_13437, n19127);
  and g29609 (n19129, n_12411, n19104);
  not g29610 (n_13438, n19129);
  and g29611 (n19130, n6305, n_13438);
  not g29612 (n_13439, n19128);
  and g29613 (n19131, n_13439, n19130);
  and g29614 (n19132, n_738, n_3232);
  not g29615 (n_13440, n19132);
  and g29616 (n19133, n_796, n_13440);
  not g29617 (n_13441, n19131);
  and g29618 (n19134, n_13441, n19133);
  and g29619 (n19135, pi0057, pi0142);
  not g29620 (n_13442, n19135);
  and g29621 (n19136, n_12415, n_13442);
  not g29622 (n_13443, n19134);
  and g29623 (n19137, n_13443, n19136);
  and g29624 (n19138, pi0142, n_12418);
  and g29625 (n19139, pi0628, pi1156);
  and g29626 (n19140, n_11789, n_11794);
  not g29627 (n_13444, n19139);
  and g29628 (n19141, pi0792, n_13444);
  not g29629 (n_13445, n19140);
  and g29630 (n19142, n_13445, n19141);
  and g29631 (n19143, n_11753, pi1153);
  and g29632 (n19144, pi0625, n_11757);
  not g29633 (n_13446, n19143);
  not g29634 (n_13447, n19144);
  and g29635 (n19145, n_13446, n_13447);
  not g29636 (n_13448, n19145);
  and g29637 (n19146, pi0778, n_13448);
  not g29638 (n_13449, n19146);
  and g29639 (n19147, n18623, n_13449);
  not g29640 (n_13450, n19138);
  not g29641 (n_13451, n19147);
  and g29642 (n19148, n_13450, n_13451);
  and g29643 (n19149, n_11783, n_11780);
  and g29644 (n19150, n_11777, n_11773);
  and g29645 (n19151, n19149, n19150);
  not g29646 (n_13452, n19148);
  and g29647 (n19152, n_13452, n19151);
  not g29648 (n_13453, n19142);
  and g29649 (n19153, n_13453, n19152);
  and g29650 (n19154, pi0647, n19153);
  and g29651 (n19155, pi1157, n_13450);
  not g29652 (n_13454, n19154);
  and g29653 (n19156, n_13454, n19155);
  and g29654 (n19157, pi0628, n19152);
  not g29655 (n_13455, n19157);
  and g29656 (n19158, n_13450, n_13455);
  not g29657 (n_13456, n19158);
  and g29658 (n19159, pi1156, n_13456);
  and g29659 (n19160, n_12320, n19138);
  and g29660 (n19161, n_11960, n18744);
  and g29661 (n19162, pi0609, n19161);
  and g29662 (n19163, pi1155, n_13450);
  not g29663 (n_13457, n19162);
  and g29664 (n19164, n_13457, n19163);
  and g29665 (n19165, n_11971, n19161);
  and g29666 (n19166, n_11768, n_13450);
  not g29667 (n_13458, n19165);
  and g29668 (n19167, n_13458, n19166);
  not g29669 (n_13459, n19164);
  not g29670 (n_13460, n19167);
  and g29671 (n19168, n_13459, n_13460);
  not g29672 (n_13461, n19168);
  and g29673 (n19169, pi0785, n_13461);
  and g29674 (n19170, n_11964, n_13450);
  not g29675 (n_13462, n19161);
  and g29676 (n19171, n_13462, n19170);
  not g29677 (n_13463, n19169);
  not g29678 (n_13464, n19171);
  and g29679 (n19172, n_13463, n_13464);
  not g29680 (n_13465, n19172);
  and g29681 (n19173, n_11981, n_13465);
  and g29682 (n19174, n_11984, n19138);
  and g29683 (n19175, pi0618, n19172);
  not g29684 (n_13466, n19174);
  and g29685 (n19176, pi1154, n_13466);
  not g29686 (n_13467, n19175);
  and g29687 (n19177, n_13467, n19176);
  and g29688 (n19178, n_11984, n19172);
  and g29689 (n19179, pi0618, n19138);
  not g29690 (n_13468, n19179);
  and g29691 (n19180, n_11413, n_13468);
  not g29692 (n_13469, n19178);
  and g29693 (n19181, n_13469, n19180);
  not g29694 (n_13470, n19177);
  not g29695 (n_13471, n19181);
  and g29696 (n19182, n_13470, n_13471);
  not g29697 (n_13472, n19182);
  and g29698 (n19183, pi0781, n_13472);
  not g29699 (n_13473, n19173);
  not g29700 (n_13474, n19183);
  and g29701 (n19184, n_13473, n_13474);
  not g29702 (n_13475, n19184);
  and g29703 (n19185, n_12315, n_13475);
  and g29704 (n19186, n_11821, n19138);
  and g29705 (n19187, pi0619, n19184);
  not g29706 (n_13476, n19186);
  and g29707 (n19188, pi1159, n_13476);
  not g29708 (n_13477, n19187);
  and g29709 (n19189, n_13477, n19188);
  and g29710 (n19190, n_11821, n19184);
  and g29711 (n19191, pi0619, n19138);
  not g29712 (n_13478, n19191);
  and g29713 (n19192, n_11405, n_13478);
  not g29714 (n_13479, n19190);
  and g29715 (n19193, n_13479, n19192);
  not g29716 (n_13480, n19189);
  not g29717 (n_13481, n19193);
  and g29718 (n19194, n_13480, n_13481);
  not g29719 (n_13482, n19194);
  and g29720 (n19195, pi0789, n_13482);
  not g29721 (n_13483, n19185);
  not g29722 (n_13484, n19195);
  and g29723 (n19196, n_13483, n_13484);
  and g29724 (n19197, pi0626, n19196);
  not g29725 (n_13485, n19160);
  and g29726 (n19198, pi1158, n_13485);
  not g29727 (n_13486, n19197);
  and g29728 (n19199, n_13486, n19198);
  and g29729 (n19200, n_12320, n19196);
  and g29730 (n19201, pi0626, n19138);
  not g29731 (n_13487, n19201);
  and g29732 (n19202, n_11397, n_13487);
  not g29733 (n_13488, n19200);
  and g29734 (n19203, n_13488, n19202);
  not g29735 (n_13489, n19199);
  not g29736 (n_13490, n19203);
  and g29737 (n19204, n_13489, n_13490);
  and g29738 (n19205, n_11401, n19204);
  and g29739 (n19206, n16635, n_13450);
  and g29740 (n19207, n_11773, n_13452);
  and g29741 (n19208, n_11777, n19207);
  not g29742 (n_13491, n19208);
  and g29743 (n19209, n_13450, n_13491);
  not g29744 (n_13492, n19206);
  and g29745 (n19210, n17871, n_13492);
  not g29746 (n_13493, n19209);
  and g29747 (n19211, n_13493, n19210);
  not g29748 (n_13494, n19205);
  not g29749 (n_13495, n19211);
  and g29750 (n19212, n_13494, n_13495);
  not g29751 (n_13496, n19212);
  and g29752 (n19213, pi0788, n_13496);
  not g29753 (n_13497, n19207);
  and g29754 (n19214, n_13450, n_13497);
  not g29755 (n_13498, n19214);
  and g29756 (n19215, pi0618, n_13498);
  and g29757 (n19216, pi0625, n18623);
  and g29758 (n19217, pi1153, n_13450);
  not g29759 (n_13499, n19216);
  and g29760 (n19218, n_13499, n19217);
  and g29761 (n19219, pi0735, n17469);
  and g29762 (n19220, pi0625, n19219);
  not g29763 (n_13500, n18744);
  and g29764 (n19221, n_13500, n_13450);
  not g29765 (n_13501, n19219);
  and g29766 (n19222, n_13501, n19221);
  not g29767 (n_13502, n19220);
  not g29768 (n_13503, n19222);
  and g29769 (n19223, n_13502, n_13503);
  not g29770 (n_13504, n19223);
  and g29771 (n19224, n_11757, n_13504);
  not g29772 (n_13505, n19218);
  and g29773 (n19225, n_11823, n_13505);
  not g29774 (n_13506, n19224);
  and g29775 (n19226, n_13506, n19225);
  and g29776 (n19227, n_13500, n_13502);
  not g29777 (n_13507, n19227);
  and g29778 (n19228, pi1153, n_13507);
  and g29779 (n19229, n_11753, n_11757);
  and g29780 (n19230, n18623, n19229);
  not g29781 (n_13508, n19230);
  and g29782 (n19231, n_13450, n_13508);
  not g29783 (n_13509, n19228);
  and g29784 (n19232, n_13509, n19231);
  not g29785 (n_13510, n19232);
  and g29786 (n19233, pi0608, n_13510);
  not g29787 (n_13511, n19226);
  not g29788 (n_13512, n19233);
  and g29789 (n19234, n_13511, n_13512);
  not g29790 (n_13513, n19234);
  and g29791 (n19235, pi0778, n_13513);
  and g29792 (n19236, n_11749, n_13503);
  not g29793 (n_13514, n19235);
  not g29794 (n_13515, n19236);
  and g29795 (n19237, n_13514, n_13515);
  not g29796 (n_13516, n19237);
  and g29797 (n19238, n_11971, n_13516);
  and g29798 (n19239, pi0609, n_13452);
  not g29799 (n_13517, n19239);
  and g29800 (n19240, n_11768, n_13517);
  not g29801 (n_13518, n19238);
  and g29802 (n19241, n_13518, n19240);
  and g29803 (n19242, n_11767, n_13459);
  not g29804 (n_13519, n19241);
  and g29805 (n19243, n_13519, n19242);
  and g29806 (n19244, pi0609, n_13516);
  and g29807 (n19245, n_11971, n_13452);
  not g29808 (n_13520, n19245);
  and g29809 (n19246, pi1155, n_13520);
  not g29810 (n_13521, n19244);
  and g29811 (n19247, n_13521, n19246);
  and g29812 (n19248, pi0660, n_13460);
  not g29813 (n_13522, n19247);
  and g29814 (n19249, n_13522, n19248);
  not g29815 (n_13523, n19243);
  not g29816 (n_13524, n19249);
  and g29817 (n19250, n_13523, n_13524);
  not g29818 (n_13525, n19250);
  and g29819 (n19251, pi0785, n_13525);
  and g29820 (n19252, n_11964, n_13516);
  not g29821 (n_13526, n19251);
  not g29822 (n_13527, n19252);
  and g29823 (n19253, n_13526, n_13527);
  not g29824 (n_13528, n19253);
  and g29825 (n19254, n_11984, n_13528);
  not g29826 (n_13529, n19215);
  and g29827 (n19255, n_11413, n_13529);
  not g29828 (n_13530, n19254);
  and g29829 (n19256, n_13530, n19255);
  and g29830 (n19257, n_11412, n_13470);
  not g29831 (n_13531, n19256);
  and g29832 (n19258, n_13531, n19257);
  and g29833 (n19259, n_11984, n_13498);
  and g29834 (n19260, pi0618, n_13528);
  not g29835 (n_13532, n19259);
  and g29836 (n19261, pi1154, n_13532);
  not g29837 (n_13533, n19260);
  and g29838 (n19262, n_13533, n19261);
  and g29839 (n19263, pi0627, n_13471);
  not g29840 (n_13534, n19262);
  and g29841 (n19264, n_13534, n19263);
  not g29842 (n_13535, n19258);
  not g29843 (n_13536, n19264);
  and g29844 (n19265, n_13535, n_13536);
  not g29845 (n_13537, n19265);
  and g29846 (n19266, pi0781, n_13537);
  and g29847 (n19267, n_11981, n_13528);
  not g29848 (n_13538, n19266);
  not g29849 (n_13539, n19267);
  and g29850 (n19268, n_13538, n_13539);
  and g29851 (n19269, n_12315, n19268);
  not g29852 (n_13540, n19268);
  and g29853 (n19270, n_11821, n_13540);
  and g29854 (n19271, pi0619, n_13493);
  not g29855 (n_13541, n19271);
  and g29856 (n19272, n_11405, n_13541);
  not g29857 (n_13542, n19270);
  and g29858 (n19273, n_13542, n19272);
  and g29859 (n19274, n_11403, n_13480);
  not g29860 (n_13543, n19273);
  and g29861 (n19275, n_13543, n19274);
  and g29862 (n19276, pi0619, n_13540);
  and g29863 (n19277, n_11821, n_13493);
  not g29864 (n_13544, n19277);
  and g29865 (n19278, pi1159, n_13544);
  not g29866 (n_13545, n19276);
  and g29867 (n19279, n_13545, n19278);
  and g29868 (n19280, pi0648, n_13481);
  not g29869 (n_13546, n19279);
  and g29870 (n19281, n_13546, n19280);
  not g29871 (n_13547, n19275);
  and g29872 (n19282, pi0789, n_13547);
  not g29873 (n_13548, n19281);
  and g29874 (n19283, n_13548, n19282);
  not g29875 (n_13549, n19269);
  and g29876 (n19284, n17970, n_13549);
  not g29877 (n_13550, n19283);
  and g29878 (n19285, n_13550, n19284);
  not g29879 (n_13551, n19213);
  not g29880 (n_13552, n19285);
  and g29881 (n19286, n_13551, n_13552);
  and g29882 (n19287, n_11789, n19286);
  not g29883 (n_13553, n19196);
  and g29884 (n19288, n_12318, n_13553);
  not g29885 (n_13554, n19204);
  and g29886 (n19289, pi0788, n_13554);
  not g29887 (n_13555, n19288);
  not g29888 (n_13556, n19289);
  and g29889 (n19290, n_13555, n_13556);
  not g29890 (n_13557, n19290);
  and g29891 (n19291, pi0628, n_13557);
  not g29892 (n_13558, n19291);
  and g29893 (n19292, n_11794, n_13558);
  not g29894 (n_13559, n19287);
  and g29895 (n19293, n_13559, n19292);
  not g29896 (n_13560, n19159);
  and g29897 (n19294, n_12354, n_13560);
  not g29898 (n_13561, n19293);
  and g29899 (n19295, n_13561, n19294);
  and g29900 (n19296, n_11789, n19152);
  not g29901 (n_13562, n19296);
  and g29902 (n19297, n_13450, n_13562);
  not g29903 (n_13563, n19297);
  and g29904 (n19298, n_11794, n_13563);
  and g29905 (n19299, pi0628, n19286);
  and g29906 (n19300, n_11789, n_13557);
  not g29907 (n_13564, n19300);
  and g29908 (n19301, pi1156, n_13564);
  not g29909 (n_13565, n19299);
  and g29910 (n19302, n_13565, n19301);
  not g29911 (n_13566, n19298);
  and g29912 (n19303, pi0629, n_13566);
  not g29913 (n_13567, n19302);
  and g29914 (n19304, n_13567, n19303);
  not g29915 (n_13568, n19295);
  not g29916 (n_13569, n19304);
  and g29917 (n19305, n_13568, n_13569);
  not g29918 (n_13570, n19305);
  and g29919 (n19306, pi0792, n_13570);
  and g29920 (n19307, n_11787, n19286);
  not g29921 (n_13571, n19306);
  not g29922 (n_13572, n19307);
  and g29923 (n19308, n_13571, n_13572);
  and g29924 (n19309, n_11806, n19308);
  and g29925 (n19310, n_12368, n19290);
  and g29926 (n19311, n17779, n19138);
  not g29927 (n_13573, n19310);
  not g29928 (n_13574, n19311);
  and g29929 (n19312, n_13573, n_13574);
  not g29930 (n_13575, n19312);
  and g29931 (n19313, pi0647, n_13575);
  not g29932 (n_13576, n19313);
  and g29933 (n19314, n_11810, n_13576);
  not g29934 (n_13577, n19309);
  and g29935 (n19315, n_13577, n19314);
  not g29936 (n_13578, n19156);
  and g29937 (n19316, n_12375, n_13578);
  not g29938 (n_13579, n19315);
  and g29939 (n19317, n_13579, n19316);
  and g29940 (n19318, n_11806, n19153);
  and g29941 (n19319, n_11810, n_13450);
  not g29942 (n_13580, n19318);
  and g29943 (n19320, n_13580, n19319);
  and g29944 (n19321, n_11806, n_13575);
  and g29945 (n19322, pi0647, n19308);
  not g29946 (n_13581, n19321);
  and g29947 (n19323, pi1157, n_13581);
  not g29948 (n_13582, n19322);
  and g29949 (n19324, n_13582, n19323);
  not g29950 (n_13583, n19320);
  and g29951 (n19325, pi0630, n_13583);
  not g29952 (n_13584, n19324);
  and g29953 (n19326, n_13584, n19325);
  not g29954 (n_13585, n19317);
  not g29955 (n_13586, n19326);
  and g29956 (n19327, n_13585, n_13586);
  not g29957 (n_13587, n19327);
  and g29958 (n19328, pi0787, n_13587);
  and g29959 (n19329, n_11803, n19308);
  not g29960 (n_13588, n19328);
  not g29961 (n_13589, n19329);
  and g29962 (n19330, n_13588, n_13589);
  not g29963 (n_13590, n19330);
  and g29964 (n19331, n_12411, n_13590);
  and g29965 (n19332, n17804, n_13450);
  and g29966 (n19333, n_12392, n19312);
  not g29967 (n_13591, n19332);
  not g29968 (n_13592, n19333);
  and g29969 (n19334, n_13591, n_13592);
  and g29970 (n19335, pi0644, n19334);
  and g29971 (n19336, n_11819, n19138);
  not g29972 (n_13593, n19336);
  and g29973 (n19337, n_12395, n_13593);
  not g29974 (n_13594, n19335);
  and g29975 (n19338, n_13594, n19337);
  and g29976 (n19339, n_11806, pi1157);
  and g29977 (n19340, pi0647, n_11810);
  not g29978 (n_13595, n19339);
  not g29979 (n_13596, n19340);
  and g29980 (n19341, n_13595, n_13596);
  not g29981 (n_13597, n19341);
  and g29982 (n19342, pi0787, n_13597);
  not g29983 (n_13598, n19342);
  and g29984 (n19343, n19153, n_13598);
  not g29985 (n_13599, n19343);
  and g29986 (n19344, n_13450, n_13599);
  not g29987 (n_13600, n19344);
  and g29988 (n19345, n_11819, n_13600);
  and g29989 (n19346, pi0644, n_13590);
  not g29990 (n_13601, n19345);
  and g29991 (n19347, pi0715, n_13601);
  not g29992 (n_13602, n19346);
  and g29993 (n19348, n_13602, n19347);
  not g29994 (n_13603, n19338);
  and g29995 (n19349, pi1160, n_13603);
  not g29996 (n_13604, n19348);
  and g29997 (n19350, n_13604, n19349);
  and g29998 (n19351, n_11819, n19334);
  and g29999 (n19352, pi0644, n19138);
  not g30000 (n_13605, n19352);
  and g30001 (n19353, pi0715, n_13605);
  not g30002 (n_13606, n19351);
  and g30003 (n19354, n_13606, n19353);
  and g30004 (n19355, pi0644, n_13600);
  and g30005 (n19356, n_11819, n_13590);
  not g30006 (n_13607, n19355);
  and g30007 (n19357, n_12395, n_13607);
  not g30008 (n_13608, n19356);
  and g30009 (n19358, n_13608, n19357);
  not g30010 (n_13609, n19354);
  and g30011 (n19359, n_12405, n_13609);
  not g30012 (n_13610, n19358);
  and g30013 (n19360, n_13610, n19359);
  not g30014 (n_13611, n19350);
  not g30015 (n_13612, n19360);
  and g30016 (n19361, n_13611, n_13612);
  not g30017 (n_13613, n19361);
  and g30018 (n19362, pi0790, n_13613);
  not g30019 (n_13614, n19331);
  and g30020 (n19363, pi0832, n_13614);
  not g30021 (n_13615, n19362);
  and g30022 (n19364, n_13615, n19363);
  not g30023 (n_13616, n19137);
  not g30024 (n_13617, n19364);
  and g30025 (po0299, n_13616, n_13617);
  and g30026 (n19366, n_9141, n_11751);
  not g30027 (n_13618, n19366);
  and g30028 (n19367, n16635, n_13618);
  and g30029 (n19368, pi0143, n_11417);
  and g30030 (n19369, n_9141, n_11743);
  not g30031 (n_13620, pi0687);
  and g30032 (n19370, n_13620, n19369);
  and g30033 (n19371, n_9141, n_11418);
  not g30034 (n_13621, n19371);
  and g30035 (n19372, n16647, n_13621);
  and g30036 (n19373, n_9141, n18072);
  and g30037 (n19374, pi0143, n_12608);
  not g30038 (n_13622, n19374);
  and g30039 (n19375, n_161, n_13622);
  not g30040 (n_13623, n19373);
  and g30041 (n19376, n_13623, n19375);
  not g30042 (n_13624, n19372);
  and g30043 (n19377, pi0687, n_13624);
  not g30044 (n_13625, n19376);
  and g30045 (n19378, n_13625, n19377);
  not g30046 (n_13626, n19370);
  and g30047 (n19379, n2571, n_13626);
  not g30048 (n_13627, n19378);
  and g30049 (n19380, n_13627, n19379);
  not g30050 (n_13628, n19368);
  not g30051 (n_13629, n19380);
  and g30052 (n19381, n_13628, n_13629);
  not g30053 (n_13630, n19381);
  and g30054 (n19382, n_11749, n_13630);
  and g30055 (n19383, n_11753, n19366);
  and g30056 (n19384, pi0625, n19381);
  not g30057 (n_13631, n19383);
  and g30058 (n19385, pi1153, n_13631);
  not g30059 (n_13632, n19384);
  and g30060 (n19386, n_13632, n19385);
  and g30061 (n19387, n_11753, n19381);
  and g30062 (n19388, pi0625, n19366);
  not g30063 (n_13633, n19388);
  and g30064 (n19389, n_11757, n_13633);
  not g30065 (n_13634, n19387);
  and g30066 (n19390, n_13634, n19389);
  not g30067 (n_13635, n19386);
  not g30068 (n_13636, n19390);
  and g30069 (n19391, n_13635, n_13636);
  not g30070 (n_13637, n19391);
  and g30071 (n19392, pi0778, n_13637);
  not g30072 (n_13638, n19382);
  not g30073 (n_13639, n19392);
  and g30074 (n19393, n_13638, n_13639);
  not g30075 (n_13640, n19393);
  and g30076 (n19394, n_11773, n_13640);
  and g30077 (n19395, n17075, n_13618);
  not g30078 (n_13641, n19394);
  not g30079 (n_13642, n19395);
  and g30080 (n19396, n_13641, n_13642);
  and g30081 (n19397, n_11777, n19396);
  and g30082 (n19398, n16639, n19366);
  not g30083 (n_13643, n19397);
  not g30084 (n_13644, n19398);
  and g30085 (n19399, n_13643, n_13644);
  and g30086 (n19400, n_11780, n19399);
  not g30087 (n_13645, n19367);
  not g30088 (n_13646, n19400);
  and g30089 (n19401, n_13645, n_13646);
  and g30090 (n19402, n_11783, n19401);
  and g30091 (n19403, n16631, n19366);
  not g30092 (n_13647, n19402);
  not g30093 (n_13648, n19403);
  and g30094 (n19404, n_13647, n_13648);
  and g30095 (n19405, n_11787, n19404);
  and g30096 (n19406, n_11789, n19366);
  not g30097 (n_13649, n19404);
  and g30098 (n19407, pi0628, n_13649);
  not g30099 (n_13650, n19406);
  and g30100 (n19408, pi1156, n_13650);
  not g30101 (n_13651, n19407);
  and g30102 (n19409, n_13651, n19408);
  and g30103 (n19410, pi0628, n19366);
  and g30104 (n19411, n_11789, n_13649);
  not g30105 (n_13652, n19410);
  and g30106 (n19412, n_11794, n_13652);
  not g30107 (n_13653, n19411);
  and g30108 (n19413, n_13653, n19412);
  not g30109 (n_13654, n19409);
  not g30110 (n_13655, n19413);
  and g30111 (n19414, n_13654, n_13655);
  not g30112 (n_13656, n19414);
  and g30113 (n19415, pi0792, n_13656);
  not g30114 (n_13657, n19405);
  not g30115 (n_13658, n19415);
  and g30116 (n19416, n_13657, n_13658);
  not g30117 (n_13659, n19416);
  and g30118 (n19417, n_11803, n_13659);
  and g30119 (n19418, n_11806, n19366);
  and g30120 (n19419, pi0647, n19416);
  not g30121 (n_13660, n19418);
  and g30122 (n19420, pi1157, n_13660);
  not g30123 (n_13661, n19419);
  and g30124 (n19421, n_13661, n19420);
  and g30125 (n19422, n_11806, n19416);
  and g30126 (n19423, pi0647, n19366);
  not g30127 (n_13662, n19423);
  and g30128 (n19424, n_11810, n_13662);
  not g30129 (n_13663, n19422);
  and g30130 (n19425, n_13663, n19424);
  not g30131 (n_13664, n19421);
  not g30132 (n_13665, n19425);
  and g30133 (n19426, n_13664, n_13665);
  not g30134 (n_13666, n19426);
  and g30135 (n19427, pi0787, n_13666);
  not g30136 (n_13667, n19417);
  not g30137 (n_13668, n19427);
  and g30138 (n19428, n_13667, n_13668);
  and g30139 (n19429, n_11819, n19428);
  and g30140 (n19430, n_11984, n19366);
  not g30141 (n_13670, n19369);
  and g30142 (n19431, pi0774, n_13670);
  and g30143 (n19432, n6135, n17244);
  and g30144 (n19433, pi0038, n19432);
  and g30145 (n19434, n_161, n17275);
  not g30146 (n_13671, n19434);
  and g30147 (n19435, pi0143, n_13671);
  not g30148 (n_13672, n17221);
  and g30149 (n19436, n_161, n_13672);
  and g30150 (n19437, n6284, n17182);
  not g30151 (n_13673, n19437);
  and g30152 (n19438, pi0038, n_13673);
  not g30153 (n_13674, n19436);
  not g30154 (n_13675, n19438);
  and g30155 (n19439, n_13674, n_13675);
  not g30156 (n_13676, pi0774);
  and g30157 (n19440, n_9141, n_13676);
  and g30158 (n19441, n19439, n19440);
  not g30159 (n_13677, n19435);
  not g30160 (n_13678, n19441);
  and g30161 (n19442, n_13677, n_13678);
  not g30162 (n_13679, n19433);
  not g30163 (n_13680, n19442);
  and g30164 (n19443, n_13679, n_13680);
  not g30165 (n_13681, n19431);
  not g30166 (n_13682, n19443);
  and g30167 (n19444, n_13681, n_13682);
  not g30168 (n_13683, n19444);
  and g30169 (n19445, n2571, n_13683);
  not g30170 (n_13684, n19445);
  and g30171 (n19446, n_13628, n_13684);
  not g30172 (n_13685, n19446);
  and g30173 (n19447, n_11960, n_13685);
  and g30174 (n19448, n17117, n_13618);
  not g30175 (n_13686, n19447);
  not g30176 (n_13687, n19448);
  and g30177 (n19449, n_13686, n_13687);
  not g30178 (n_13688, n19449);
  and g30179 (n19450, n_11964, n_13688);
  and g30180 (n19451, n_11967, n_13618);
  and g30181 (n19452, pi0609, n19447);
  not g30182 (n_13689, n19451);
  not g30183 (n_13690, n19452);
  and g30184 (n19453, n_13689, n_13690);
  not g30185 (n_13691, n19453);
  and g30186 (n19454, pi1155, n_13691);
  and g30187 (n19455, n_11972, n_13618);
  and g30188 (n19456, n_11971, n19447);
  not g30189 (n_13692, n19455);
  not g30190 (n_13693, n19456);
  and g30191 (n19457, n_13692, n_13693);
  not g30192 (n_13694, n19457);
  and g30193 (n19458, n_11768, n_13694);
  not g30194 (n_13695, n19454);
  not g30195 (n_13696, n19458);
  and g30196 (n19459, n_13695, n_13696);
  not g30197 (n_13697, n19459);
  and g30198 (n19460, pi0785, n_13697);
  not g30199 (n_13698, n19450);
  not g30200 (n_13699, n19460);
  and g30201 (n19461, n_13698, n_13699);
  and g30202 (n19462, pi0618, n19461);
  not g30203 (n_13700, n19430);
  and g30204 (n19463, pi1154, n_13700);
  not g30205 (n_13701, n19462);
  and g30206 (n19464, n_13701, n19463);
  and g30207 (n19465, n_162, n_12240);
  not g30208 (n_13702, n17485);
  and g30209 (n19466, pi0039, n_13702);
  not g30210 (n_13703, n19465);
  not g30211 (n_13704, n19466);
  and g30212 (n19467, n_13703, n_13704);
  and g30213 (n19468, n_161, n19467);
  and g30214 (n19469, pi0143, n19468);
  and g30215 (n19470, pi0038, n18175);
  and g30216 (n19471, n16641, n_12023);
  and g30217 (n19472, pi0038, n19471);
  not g30218 (n_13705, n17404);
  and g30219 (n19473, pi0039, n_13705);
  and g30220 (n19474, n_162, n_12230);
  not g30221 (n_13706, n19473);
  not g30222 (n_13707, n19474);
  and g30223 (n19475, n_13706, n_13707);
  not g30224 (n_13708, n19475);
  and g30225 (n19476, n_161, n_13708);
  not g30226 (n_13709, n19472);
  not g30227 (n_13710, n19476);
  and g30228 (n19477, n_13709, n_13710);
  and g30229 (n19478, n_9141, n19477);
  not g30230 (n_13711, n19470);
  and g30236 (n19482, n_162, n_12694);
  and g30237 (n19483, n_161, n19482);
  and g30238 (n19484, pi0039, n_12180);
  and g30239 (n19485, n_162, n17490);
  not g30240 (n_13714, n19485);
  and g30241 (n19486, pi0038, n_13714);
  not g30242 (n_13715, n19483);
  not g30243 (n_13716, n19486);
  and g30244 (n19487, n_13715, n_13716);
  not g30245 (n_13717, n19484);
  and g30246 (n19488, n_13717, n19487);
  not g30247 (n_13718, n19488);
  and g30248 (n19489, n_9141, n_13718);
  and g30249 (n19490, n6284, n_12121);
  not g30250 (n_13719, n19490);
  and g30251 (n19491, pi0038, n_13719);
  not g30252 (n_13720, n17605);
  and g30253 (n19492, pi0039, n_13720);
  and g30254 (n19493, n_12243, n17234);
  not g30255 (n_13721, n19492);
  not g30256 (n_13722, n19493);
  and g30257 (n19494, n_13721, n_13722);
  not g30258 (n_13723, n19494);
  and g30259 (n19495, n_161, n_13723);
  not g30260 (n_13724, n19491);
  not g30261 (n_13725, n19495);
  and g30262 (n19496, n_13724, n_13725);
  and g30263 (n19497, pi0143, n19496);
  not g30264 (n_13726, n19489);
  and g30265 (n19498, n_13676, n_13726);
  not g30266 (n_13727, n19497);
  and g30267 (n19499, n_13727, n19498);
  not g30268 (n_13728, n19499);
  and g30269 (n19500, pi0687, n_13728);
  not g30270 (n_13729, n19481);
  and g30271 (n19501, n_13729, n19500);
  and g30272 (n19502, n_13620, n19444);
  not g30273 (n_13730, n19501);
  and g30274 (n19503, n2571, n_13730);
  not g30275 (n_13731, n19502);
  and g30276 (n19504, n_13731, n19503);
  not g30277 (n_13732, n19504);
  and g30278 (n19505, n_13628, n_13732);
  and g30279 (n19506, n_11753, n19505);
  and g30280 (n19507, pi0625, n19446);
  not g30281 (n_13733, n19507);
  and g30282 (n19508, n_11757, n_13733);
  not g30283 (n_13734, n19506);
  and g30284 (n19509, n_13734, n19508);
  and g30285 (n19510, n_11823, n_13635);
  not g30286 (n_13735, n19509);
  and g30287 (n19511, n_13735, n19510);
  and g30288 (n19512, n_11753, n19446);
  and g30289 (n19513, pi0625, n19505);
  not g30290 (n_13736, n19512);
  and g30291 (n19514, pi1153, n_13736);
  not g30292 (n_13737, n19513);
  and g30293 (n19515, n_13737, n19514);
  and g30294 (n19516, pi0608, n_13636);
  not g30295 (n_13738, n19515);
  and g30296 (n19517, n_13738, n19516);
  not g30297 (n_13739, n19511);
  not g30298 (n_13740, n19517);
  and g30299 (n19518, n_13739, n_13740);
  not g30300 (n_13741, n19518);
  and g30301 (n19519, pi0778, n_13741);
  and g30302 (n19520, n_11749, n19505);
  not g30303 (n_13742, n19519);
  not g30304 (n_13743, n19520);
  and g30305 (n19521, n_13742, n_13743);
  not g30306 (n_13744, n19521);
  and g30307 (n19522, n_11971, n_13744);
  and g30308 (n19523, pi0609, n19393);
  not g30309 (n_13745, n19523);
  and g30310 (n19524, n_11768, n_13745);
  not g30311 (n_13746, n19522);
  and g30312 (n19525, n_13746, n19524);
  and g30313 (n19526, n_11767, n_13695);
  not g30314 (n_13747, n19525);
  and g30315 (n19527, n_13747, n19526);
  and g30316 (n19528, n_11971, n19393);
  and g30317 (n19529, pi0609, n_13744);
  not g30318 (n_13748, n19528);
  and g30319 (n19530, pi1155, n_13748);
  not g30320 (n_13749, n19529);
  and g30321 (n19531, n_13749, n19530);
  and g30322 (n19532, pi0660, n_13696);
  not g30323 (n_13750, n19531);
  and g30324 (n19533, n_13750, n19532);
  not g30325 (n_13751, n19527);
  not g30326 (n_13752, n19533);
  and g30327 (n19534, n_13751, n_13752);
  not g30328 (n_13753, n19534);
  and g30329 (n19535, pi0785, n_13753);
  and g30330 (n19536, n_11964, n_13744);
  not g30331 (n_13754, n19535);
  not g30332 (n_13755, n19536);
  and g30333 (n19537, n_13754, n_13755);
  not g30334 (n_13756, n19537);
  and g30335 (n19538, n_11984, n_13756);
  and g30336 (n19539, pi0618, n19396);
  not g30337 (n_13757, n19539);
  and g30338 (n19540, n_11413, n_13757);
  not g30339 (n_13758, n19538);
  and g30340 (n19541, n_13758, n19540);
  not g30341 (n_13759, n19464);
  and g30342 (n19542, n_11412, n_13759);
  not g30343 (n_13760, n19541);
  and g30344 (n19543, n_13760, n19542);
  and g30345 (n19544, n_11984, n19461);
  and g30346 (n19545, pi0618, n19366);
  not g30347 (n_13761, n19545);
  and g30348 (n19546, n_11413, n_13761);
  not g30349 (n_13762, n19544);
  and g30350 (n19547, n_13762, n19546);
  and g30351 (n19548, n_11984, n19396);
  and g30352 (n19549, pi0618, n_13756);
  not g30353 (n_13763, n19548);
  and g30354 (n19550, pi1154, n_13763);
  not g30355 (n_13764, n19549);
  and g30356 (n19551, n_13764, n19550);
  not g30357 (n_13765, n19547);
  and g30358 (n19552, pi0627, n_13765);
  not g30359 (n_13766, n19551);
  and g30360 (n19553, n_13766, n19552);
  not g30361 (n_13767, n19543);
  not g30362 (n_13768, n19553);
  and g30363 (n19554, n_13767, n_13768);
  not g30364 (n_13769, n19554);
  and g30365 (n19555, pi0781, n_13769);
  and g30366 (n19556, n_11981, n_13756);
  not g30367 (n_13770, n19555);
  not g30368 (n_13771, n19556);
  and g30369 (n19557, n_13770, n_13771);
  not g30370 (n_13772, n19557);
  and g30371 (n19558, n_11821, n_13772);
  not g30372 (n_13773, n19399);
  and g30373 (n19559, pi0619, n_13773);
  not g30374 (n_13774, n19559);
  and g30375 (n19560, n_11405, n_13774);
  not g30376 (n_13775, n19558);
  and g30377 (n19561, n_13775, n19560);
  and g30378 (n19562, n_11821, n19366);
  not g30379 (n_13776, n19461);
  and g30380 (n19563, n_11981, n_13776);
  and g30381 (n19564, n_13759, n_13765);
  not g30382 (n_13777, n19564);
  and g30383 (n19565, pi0781, n_13777);
  not g30384 (n_13778, n19563);
  not g30385 (n_13779, n19565);
  and g30386 (n19566, n_13778, n_13779);
  and g30387 (n19567, pi0619, n19566);
  not g30388 (n_13780, n19562);
  and g30389 (n19568, pi1159, n_13780);
  not g30390 (n_13781, n19567);
  and g30391 (n19569, n_13781, n19568);
  not g30392 (n_13782, n19569);
  and g30393 (n19570, n_11403, n_13782);
  not g30394 (n_13783, n19561);
  and g30395 (n19571, n_13783, n19570);
  and g30396 (n19572, pi0619, n_13772);
  and g30397 (n19573, n_11821, n_13773);
  not g30398 (n_13784, n19573);
  and g30399 (n19574, pi1159, n_13784);
  not g30400 (n_13785, n19572);
  and g30401 (n19575, n_13785, n19574);
  and g30402 (n19576, n_11821, n19566);
  and g30403 (n19577, pi0619, n19366);
  not g30404 (n_13786, n19577);
  and g30405 (n19578, n_11405, n_13786);
  not g30406 (n_13787, n19576);
  and g30407 (n19579, n_13787, n19578);
  not g30408 (n_13788, n19579);
  and g30409 (n19580, pi0648, n_13788);
  not g30410 (n_13789, n19575);
  and g30411 (n19581, n_13789, n19580);
  not g30412 (n_13790, n19571);
  not g30413 (n_13791, n19581);
  and g30414 (n19582, n_13790, n_13791);
  not g30415 (n_13792, n19582);
  and g30416 (n19583, pi0789, n_13792);
  and g30417 (n19584, n_12315, n_13772);
  not g30418 (n_13793, n19583);
  not g30419 (n_13794, n19584);
  and g30420 (n19585, n_13793, n_13794);
  and g30421 (n19586, n_12318, n19585);
  and g30422 (n19587, n_12320, n19585);
  not g30423 (n_13795, n19401);
  and g30424 (n19588, pi0626, n_13795);
  not g30425 (n_13796, n19588);
  and g30426 (n19589, n_11395, n_13796);
  not g30427 (n_13797, n19587);
  and g30428 (n19590, n_13797, n19589);
  not g30429 (n_13798, n19566);
  and g30430 (n19591, n_12315, n_13798);
  and g30431 (n19592, n_13782, n_13788);
  not g30432 (n_13799, n19592);
  and g30433 (n19593, pi0789, n_13799);
  not g30434 (n_13800, n19591);
  not g30435 (n_13801, n19593);
  and g30436 (n19594, n_13800, n_13801);
  and g30437 (n19595, n_12320, n19594);
  and g30438 (n19596, pi0626, n19366);
  not g30439 (n_13802, n19596);
  and g30440 (n19597, n_11397, n_13802);
  not g30441 (n_13803, n19595);
  and g30442 (n19598, n_13803, n19597);
  not g30443 (n_13804, n19598);
  and g30444 (n19599, n_12330, n_13804);
  not g30445 (n_13805, n19590);
  not g30446 (n_13806, n19599);
  and g30447 (n19600, n_13805, n_13806);
  and g30448 (n19601, pi0626, n19585);
  and g30449 (n19602, n_12320, n_13795);
  not g30450 (n_13807, n19602);
  and g30451 (n19603, pi0641, n_13807);
  not g30452 (n_13808, n19601);
  and g30453 (n19604, n_13808, n19603);
  and g30454 (n19605, n_12320, n19366);
  and g30455 (n19606, pi0626, n19594);
  not g30456 (n_13809, n19605);
  and g30457 (n19607, pi1158, n_13809);
  not g30458 (n_13810, n19606);
  and g30459 (n19608, n_13810, n19607);
  not g30460 (n_13811, n19608);
  and g30461 (n19609, n_12338, n_13811);
  not g30462 (n_13812, n19604);
  not g30463 (n_13813, n19609);
  and g30464 (n19610, n_13812, n_13813);
  not g30465 (n_13814, n19600);
  not g30466 (n_13815, n19610);
  and g30467 (n19611, n_13814, n_13815);
  not g30468 (n_13816, n19611);
  and g30469 (n19612, pi0788, n_13816);
  not g30470 (n_13817, n19586);
  not g30471 (n_13818, n19612);
  and g30472 (n19613, n_13817, n_13818);
  and g30473 (n19614, n_11789, n19613);
  and g30474 (n19615, n_13804, n_13811);
  not g30475 (n_13819, n19615);
  and g30476 (n19616, pi0788, n_13819);
  not g30477 (n_13820, n19594);
  and g30478 (n19617, n_12318, n_13820);
  not g30479 (n_13821, n19616);
  not g30480 (n_13822, n19617);
  and g30481 (n19618, n_13821, n_13822);
  and g30482 (n19619, pi0628, n19618);
  not g30483 (n_13823, n19619);
  and g30484 (n19620, n_11794, n_13823);
  not g30485 (n_13824, n19614);
  and g30486 (n19621, n_13824, n19620);
  and g30487 (n19622, n_12354, n_13654);
  not g30488 (n_13825, n19621);
  and g30489 (n19623, n_13825, n19622);
  and g30490 (n19624, pi0628, n19613);
  and g30491 (n19625, n_11789, n19618);
  not g30492 (n_13826, n19625);
  and g30493 (n19626, pi1156, n_13826);
  not g30494 (n_13827, n19624);
  and g30495 (n19627, n_13827, n19626);
  and g30496 (n19628, pi0629, n_13655);
  not g30497 (n_13828, n19627);
  and g30498 (n19629, n_13828, n19628);
  not g30499 (n_13829, n19623);
  not g30500 (n_13830, n19629);
  and g30501 (n19630, n_13829, n_13830);
  not g30502 (n_13831, n19630);
  and g30503 (n19631, pi0792, n_13831);
  and g30504 (n19632, n_11787, n19613);
  not g30505 (n_13832, n19631);
  not g30506 (n_13833, n19632);
  and g30507 (n19633, n_13832, n_13833);
  not g30508 (n_13834, n19633);
  and g30509 (n19634, n_11806, n_13834);
  and g30510 (n19635, n_12368, n19618);
  and g30511 (n19636, n17779, n19366);
  not g30512 (n_13835, n19635);
  not g30513 (n_13836, n19636);
  and g30514 (n19637, n_13835, n_13836);
  not g30515 (n_13837, n19637);
  and g30516 (n19638, pi0647, n_13837);
  not g30517 (n_13838, n19638);
  and g30518 (n19639, n_11810, n_13838);
  not g30519 (n_13839, n19634);
  and g30520 (n19640, n_13839, n19639);
  and g30521 (n19641, n_12375, n_13664);
  not g30522 (n_13840, n19640);
  and g30523 (n19642, n_13840, n19641);
  and g30524 (n19643, pi0647, n_13834);
  and g30525 (n19644, n_11806, n_13837);
  not g30526 (n_13841, n19644);
  and g30527 (n19645, pi1157, n_13841);
  not g30528 (n_13842, n19643);
  and g30529 (n19646, n_13842, n19645);
  and g30530 (n19647, pi0630, n_13665);
  not g30531 (n_13843, n19646);
  and g30532 (n19648, n_13843, n19647);
  not g30533 (n_13844, n19642);
  not g30534 (n_13845, n19648);
  and g30535 (n19649, n_13844, n_13845);
  not g30536 (n_13846, n19649);
  and g30537 (n19650, pi0787, n_13846);
  and g30538 (n19651, n_11803, n_13834);
  not g30539 (n_13847, n19650);
  not g30540 (n_13848, n19651);
  and g30541 (n19652, n_13847, n_13848);
  not g30542 (n_13849, n19652);
  and g30543 (n19653, pi0644, n_13849);
  not g30544 (n_13850, n19429);
  and g30545 (n19654, pi0715, n_13850);
  not g30546 (n_13851, n19653);
  and g30547 (n19655, n_13851, n19654);
  and g30548 (n19656, n17804, n_13618);
  and g30549 (n19657, n_12392, n19637);
  not g30550 (n_13852, n19656);
  not g30551 (n_13853, n19657);
  and g30552 (n19658, n_13852, n_13853);
  and g30553 (n19659, pi0644, n19658);
  and g30554 (n19660, n_11819, n19366);
  not g30555 (n_13854, n19660);
  and g30556 (n19661, n_12395, n_13854);
  not g30557 (n_13855, n19659);
  and g30558 (n19662, n_13855, n19661);
  not g30559 (n_13856, n19662);
  and g30560 (n19663, pi1160, n_13856);
  not g30561 (n_13857, n19655);
  and g30562 (n19664, n_13857, n19663);
  and g30563 (n19665, n_11819, n_13849);
  and g30564 (n19666, pi0644, n19428);
  not g30565 (n_13858, n19666);
  and g30566 (n19667, n_12395, n_13858);
  not g30567 (n_13859, n19665);
  and g30568 (n19668, n_13859, n19667);
  and g30569 (n19669, n_11819, n19658);
  and g30570 (n19670, pi0644, n19366);
  not g30571 (n_13860, n19670);
  and g30572 (n19671, pi0715, n_13860);
  not g30573 (n_13861, n19669);
  and g30574 (n19672, n_13861, n19671);
  not g30575 (n_13862, n19672);
  and g30576 (n19673, n_12405, n_13862);
  not g30577 (n_13863, n19668);
  and g30578 (n19674, n_13863, n19673);
  not g30579 (n_13864, n19664);
  and g30580 (n19675, pi0790, n_13864);
  not g30581 (n_13865, n19674);
  and g30582 (n19676, n_13865, n19675);
  and g30583 (n19677, n_12411, n19652);
  not g30584 (n_13866, n19677);
  and g30585 (n19678, n_4226, n_13866);
  not g30586 (n_13867, n19676);
  and g30587 (n19679, n_13867, n19678);
  and g30588 (n19680, n_9141, po1038);
  not g30589 (n_13868, n19680);
  and g30590 (n19681, n_12415, n_13868);
  not g30591 (n_13869, n19679);
  and g30592 (n19682, n_13869, n19681);
  and g30593 (n19683, n_9141, n_12418);
  and g30594 (n19684, n_11806, n19683);
  and g30595 (n19685, pi0687, n16645);
  not g30596 (n_13870, n19683);
  not g30597 (n_13871, n19685);
  and g30598 (n19686, n_13870, n_13871);
  and g30599 (n19687, n_11749, n19686);
  and g30600 (n19688, n_11753, n19685);
  not g30601 (n_13872, n19686);
  not g30602 (n_13873, n19688);
  and g30603 (n19689, n_13872, n_13873);
  not g30604 (n_13874, n19689);
  and g30605 (n19690, pi1153, n_13874);
  and g30606 (n19691, n_11757, n_13870);
  and g30607 (n19692, n_13873, n19691);
  not g30608 (n_13875, n19690);
  not g30609 (n_13876, n19692);
  and g30610 (n19693, n_13875, n_13876);
  not g30611 (n_13877, n19693);
  and g30612 (n19694, pi0778, n_13877);
  not g30613 (n_13878, n19687);
  not g30614 (n_13879, n19694);
  and g30615 (n19695, n_13878, n_13879);
  and g30616 (n19696, n_12429, n19695);
  and g30617 (n19697, n_12430, n19696);
  and g30618 (n19698, n_12431, n19697);
  and g30619 (n19699, n_12432, n19698);
  and g30620 (n19700, n_12436, n19699);
  and g30621 (n19701, pi0647, n19700);
  not g30622 (n_13880, n19684);
  and g30623 (n19702, pi1157, n_13880);
  not g30624 (n_13881, n19701);
  and g30625 (n19703, n_13881, n19702);
  and g30626 (n19704, n_12439, n19699);
  not g30627 (n_13882, n19704);
  and g30628 (n19705, pi1156, n_13882);
  and g30629 (n19706, n17871, n19698);
  and g30630 (n19707, n_12320, n19683);
  and g30631 (n19708, n_13676, n17244);
  not g30632 (n_13883, n19708);
  and g30633 (n19709, n_13870, n_13883);
  not g30634 (n_13884, n19709);
  and g30635 (n19710, n_12448, n_13884);
  not g30636 (n_13885, n19710);
  and g30637 (n19711, n_11964, n_13885);
  and g30638 (n19712, n_12451, n_13884);
  not g30639 (n_13886, n19712);
  and g30640 (n19713, pi1155, n_13886);
  and g30641 (n19714, n_12453, n19710);
  not g30642 (n_13887, n19714);
  and g30643 (n19715, n_11768, n_13887);
  not g30644 (n_13888, n19713);
  not g30645 (n_13889, n19715);
  and g30646 (n19716, n_13888, n_13889);
  not g30647 (n_13890, n19716);
  and g30648 (n19717, pi0785, n_13890);
  not g30649 (n_13891, n19711);
  not g30650 (n_13892, n19717);
  and g30651 (n19718, n_13891, n_13892);
  not g30652 (n_13893, n19718);
  and g30653 (n19719, n_11981, n_13893);
  and g30654 (n19720, n_12461, n19718);
  not g30655 (n_13894, n19720);
  and g30656 (n19721, pi1154, n_13894);
  and g30657 (n19722, n_12463, n19718);
  not g30658 (n_13895, n19722);
  and g30659 (n19723, n_11413, n_13895);
  not g30660 (n_13896, n19721);
  not g30661 (n_13897, n19723);
  and g30662 (n19724, n_13896, n_13897);
  not g30663 (n_13898, n19724);
  and g30664 (n19725, pi0781, n_13898);
  not g30665 (n_13899, n19719);
  not g30666 (n_13900, n19725);
  and g30667 (n19726, n_13899, n_13900);
  not g30668 (n_13901, n19726);
  and g30669 (n19727, n_12315, n_13901);
  and g30670 (n19728, n_11821, n19683);
  and g30671 (n19729, pi0619, n19726);
  not g30672 (n_13902, n19728);
  and g30673 (n19730, pi1159, n_13902);
  not g30674 (n_13903, n19729);
  and g30675 (n19731, n_13903, n19730);
  and g30676 (n19732, n_11821, n19726);
  and g30677 (n19733, pi0619, n19683);
  not g30678 (n_13904, n19733);
  and g30679 (n19734, n_11405, n_13904);
  not g30680 (n_13905, n19732);
  and g30681 (n19735, n_13905, n19734);
  not g30682 (n_13906, n19731);
  not g30683 (n_13907, n19735);
  and g30684 (n19736, n_13906, n_13907);
  not g30685 (n_13908, n19736);
  and g30686 (n19737, pi0789, n_13908);
  not g30687 (n_13909, n19727);
  not g30688 (n_13910, n19737);
  and g30689 (n19738, n_13909, n_13910);
  and g30690 (n19739, pi0626, n19738);
  not g30691 (n_13911, n19707);
  and g30692 (n19740, pi1158, n_13911);
  not g30693 (n_13912, n19739);
  and g30694 (n19741, n_13912, n19740);
  and g30695 (n19742, n_12320, n19738);
  and g30696 (n19743, pi0626, n19683);
  not g30697 (n_13913, n19743);
  and g30698 (n19744, n_11397, n_13913);
  not g30699 (n_13914, n19742);
  and g30700 (n19745, n_13914, n19744);
  not g30701 (n_13915, n19741);
  not g30702 (n_13916, n19745);
  and g30703 (n19746, n_13915, n_13916);
  and g30704 (n19747, n_11401, n19746);
  not g30705 (n_13917, n19706);
  not g30706 (n_13918, n19747);
  and g30707 (n19748, n_13917, n_13918);
  not g30708 (n_13919, n19748);
  and g30709 (n19749, pi0788, n_13919);
  and g30710 (n19750, pi0618, n19696);
  and g30711 (n19751, pi0609, n19695);
  and g30712 (n19752, n_11866, n_13872);
  and g30713 (n19753, pi0625, n19752);
  not g30714 (n_13920, n19752);
  and g30715 (n19754, n19709, n_13920);
  not g30716 (n_13921, n19753);
  not g30717 (n_13922, n19754);
  and g30718 (n19755, n_13921, n_13922);
  not g30719 (n_13923, n19755);
  and g30720 (n19756, n19691, n_13923);
  and g30721 (n19757, n_11823, n_13875);
  not g30722 (n_13924, n19756);
  and g30723 (n19758, n_13924, n19757);
  and g30724 (n19759, pi1153, n19709);
  and g30725 (n19760, n_13921, n19759);
  and g30726 (n19761, pi0608, n_13876);
  not g30727 (n_13925, n19760);
  and g30728 (n19762, n_13925, n19761);
  not g30729 (n_13926, n19758);
  not g30730 (n_13927, n19762);
  and g30731 (n19763, n_13926, n_13927);
  not g30732 (n_13928, n19763);
  and g30733 (n19764, pi0778, n_13928);
  and g30734 (n19765, n_11749, n_13922);
  not g30735 (n_13929, n19764);
  not g30736 (n_13930, n19765);
  and g30737 (n19766, n_13929, n_13930);
  not g30738 (n_13931, n19766);
  and g30739 (n19767, n_11971, n_13931);
  not g30740 (n_13932, n19751);
  and g30741 (n19768, n_11768, n_13932);
  not g30742 (n_13933, n19767);
  and g30743 (n19769, n_13933, n19768);
  and g30744 (n19770, n_11767, n_13888);
  not g30745 (n_13934, n19769);
  and g30746 (n19771, n_13934, n19770);
  and g30747 (n19772, n_11971, n19695);
  and g30748 (n19773, pi0609, n_13931);
  not g30749 (n_13935, n19772);
  and g30750 (n19774, pi1155, n_13935);
  not g30751 (n_13936, n19773);
  and g30752 (n19775, n_13936, n19774);
  and g30753 (n19776, pi0660, n_13889);
  not g30754 (n_13937, n19775);
  and g30755 (n19777, n_13937, n19776);
  not g30756 (n_13938, n19771);
  not g30757 (n_13939, n19777);
  and g30758 (n19778, n_13938, n_13939);
  not g30759 (n_13940, n19778);
  and g30760 (n19779, pi0785, n_13940);
  and g30761 (n19780, n_11964, n_13931);
  not g30762 (n_13941, n19779);
  not g30763 (n_13942, n19780);
  and g30764 (n19781, n_13941, n_13942);
  not g30765 (n_13943, n19781);
  and g30766 (n19782, n_11984, n_13943);
  not g30767 (n_13944, n19750);
  and g30768 (n19783, n_11413, n_13944);
  not g30769 (n_13945, n19782);
  and g30770 (n19784, n_13945, n19783);
  and g30771 (n19785, n_11412, n_13896);
  not g30772 (n_13946, n19784);
  and g30773 (n19786, n_13946, n19785);
  and g30774 (n19787, n_11984, n19696);
  and g30775 (n19788, pi0618, n_13943);
  not g30776 (n_13947, n19787);
  and g30777 (n19789, pi1154, n_13947);
  not g30778 (n_13948, n19788);
  and g30779 (n19790, n_13948, n19789);
  and g30780 (n19791, pi0627, n_13897);
  not g30781 (n_13949, n19790);
  and g30782 (n19792, n_13949, n19791);
  not g30783 (n_13950, n19786);
  not g30784 (n_13951, n19792);
  and g30785 (n19793, n_13950, n_13951);
  not g30786 (n_13952, n19793);
  and g30787 (n19794, pi0781, n_13952);
  and g30788 (n19795, n_11981, n_13943);
  not g30789 (n_13953, n19794);
  not g30790 (n_13954, n19795);
  and g30791 (n19796, n_13953, n_13954);
  and g30792 (n19797, n_12315, n19796);
  not g30793 (n_13955, n19796);
  and g30794 (n19798, n_11821, n_13955);
  and g30795 (n19799, pi0619, n19697);
  not g30796 (n_13956, n19799);
  and g30797 (n19800, n_11405, n_13956);
  not g30798 (n_13957, n19798);
  and g30799 (n19801, n_13957, n19800);
  and g30800 (n19802, n_11403, n_13906);
  not g30801 (n_13958, n19801);
  and g30802 (n19803, n_13958, n19802);
  and g30803 (n19804, n_11821, n19697);
  and g30804 (n19805, pi0619, n_13955);
  not g30805 (n_13959, n19804);
  and g30806 (n19806, pi1159, n_13959);
  not g30807 (n_13960, n19805);
  and g30808 (n19807, n_13960, n19806);
  and g30809 (n19808, pi0648, n_13907);
  not g30810 (n_13961, n19807);
  and g30811 (n19809, n_13961, n19808);
  not g30812 (n_13962, n19803);
  and g30813 (n19810, pi0789, n_13962);
  not g30814 (n_13963, n19809);
  and g30815 (n19811, n_13963, n19810);
  not g30816 (n_13964, n19797);
  and g30817 (n19812, n17970, n_13964);
  not g30818 (n_13965, n19811);
  and g30819 (n19813, n_13965, n19812);
  not g30820 (n_13966, n19749);
  not g30821 (n_13967, n19813);
  and g30822 (n19814, n_13966, n_13967);
  not g30823 (n_13968, n19814);
  and g30824 (n19815, n_11789, n_13968);
  not g30825 (n_13969, n19738);
  and g30826 (n19816, n_12318, n_13969);
  not g30827 (n_13970, n19746);
  and g30828 (n19817, pi0788, n_13970);
  not g30829 (n_13971, n19816);
  not g30830 (n_13972, n19817);
  and g30831 (n19818, n_13971, n_13972);
  and g30832 (n19819, pi0628, n19818);
  not g30833 (n_13973, n19819);
  and g30834 (n19820, n_11794, n_13973);
  not g30835 (n_13974, n19815);
  and g30836 (n19821, n_13974, n19820);
  not g30837 (n_13975, n19705);
  and g30838 (n19822, n_12354, n_13975);
  not g30839 (n_13976, n19821);
  and g30840 (n19823, n_13976, n19822);
  and g30841 (n19824, n_12547, n19699);
  not g30842 (n_13977, n19824);
  and g30843 (n19825, n_11794, n_13977);
  and g30844 (n19826, n_11789, n19818);
  and g30845 (n19827, pi0628, n_13968);
  not g30846 (n_13978, n19826);
  and g30847 (n19828, pi1156, n_13978);
  not g30848 (n_13979, n19827);
  and g30849 (n19829, n_13979, n19828);
  not g30850 (n_13980, n19825);
  and g30851 (n19830, pi0629, n_13980);
  not g30852 (n_13981, n19829);
  and g30853 (n19831, n_13981, n19830);
  not g30854 (n_13982, n19823);
  not g30855 (n_13983, n19831);
  and g30856 (n19832, n_13982, n_13983);
  not g30857 (n_13984, n19832);
  and g30858 (n19833, pi0792, n_13984);
  and g30859 (n19834, n_11787, n_13968);
  not g30860 (n_13985, n19833);
  not g30861 (n_13986, n19834);
  and g30862 (n19835, n_13985, n_13986);
  not g30863 (n_13987, n19835);
  and g30864 (n19836, n_11806, n_13987);
  and g30865 (n19837, n_12368, n19818);
  and g30866 (n19838, n17779, n19683);
  not g30867 (n_13988, n19837);
  not g30868 (n_13989, n19838);
  and g30869 (n19839, n_13988, n_13989);
  not g30870 (n_13990, n19839);
  and g30871 (n19840, pi0647, n_13990);
  not g30872 (n_13991, n19840);
  and g30873 (n19841, n_11810, n_13991);
  not g30874 (n_13992, n19836);
  and g30875 (n19842, n_13992, n19841);
  not g30876 (n_13993, n19703);
  and g30877 (n19843, n_12375, n_13993);
  not g30878 (n_13994, n19842);
  and g30879 (n19844, n_13994, n19843);
  and g30880 (n19845, n_11806, n19700);
  and g30881 (n19846, pi0647, n19683);
  not g30882 (n_13995, n19846);
  and g30883 (n19847, n_11810, n_13995);
  not g30884 (n_13996, n19845);
  and g30885 (n19848, n_13996, n19847);
  and g30886 (n19849, pi0647, n_13987);
  and g30887 (n19850, n_11806, n_13990);
  not g30888 (n_13997, n19850);
  and g30889 (n19851, pi1157, n_13997);
  not g30890 (n_13998, n19849);
  and g30891 (n19852, n_13998, n19851);
  not g30892 (n_13999, n19848);
  and g30893 (n19853, pi0630, n_13999);
  not g30894 (n_14000, n19852);
  and g30895 (n19854, n_14000, n19853);
  not g30896 (n_14001, n19844);
  not g30897 (n_14002, n19854);
  and g30898 (n19855, n_14001, n_14002);
  not g30899 (n_14003, n19855);
  and g30900 (n19856, pi0787, n_14003);
  and g30901 (n19857, n_11803, n_13987);
  not g30902 (n_14004, n19856);
  not g30903 (n_14005, n19857);
  and g30904 (n19858, n_14004, n_14005);
  not g30905 (n_14006, n19858);
  and g30906 (n19859, n_12411, n_14006);
  not g30907 (n_14007, n19700);
  and g30908 (n19860, n_11803, n_14007);
  and g30909 (n19861, n_13993, n_13999);
  not g30910 (n_14008, n19861);
  and g30911 (n19862, pi0787, n_14008);
  not g30912 (n_14009, n19860);
  not g30913 (n_14010, n19862);
  and g30914 (n19863, n_14009, n_14010);
  and g30915 (n19864, n_11819, n19863);
  and g30916 (n19865, pi0644, n_14006);
  not g30917 (n_14011, n19864);
  and g30918 (n19866, pi0715, n_14011);
  not g30919 (n_14012, n19865);
  and g30920 (n19867, n_14012, n19866);
  and g30921 (n19868, n17804, n_13870);
  and g30922 (n19869, n_12392, n19839);
  not g30923 (n_14013, n19868);
  not g30924 (n_14014, n19869);
  and g30925 (n19870, n_14013, n_14014);
  and g30926 (n19871, pi0644, n19870);
  and g30927 (n19872, n_11819, n19683);
  not g30928 (n_14015, n19872);
  and g30929 (n19873, n_12395, n_14015);
  not g30930 (n_14016, n19871);
  and g30931 (n19874, n_14016, n19873);
  not g30932 (n_14017, n19874);
  and g30933 (n19875, pi1160, n_14017);
  not g30934 (n_14018, n19867);
  and g30935 (n19876, n_14018, n19875);
  and g30936 (n19877, n_11819, n19870);
  and g30937 (n19878, pi0644, n19683);
  not g30938 (n_14019, n19878);
  and g30939 (n19879, pi0715, n_14019);
  not g30940 (n_14020, n19877);
  and g30941 (n19880, n_14020, n19879);
  and g30942 (n19881, pi0644, n19863);
  and g30943 (n19882, n_11819, n_14006);
  not g30944 (n_14021, n19881);
  and g30945 (n19883, n_12395, n_14021);
  not g30946 (n_14022, n19882);
  and g30947 (n19884, n_14022, n19883);
  not g30948 (n_14023, n19880);
  and g30949 (n19885, n_12405, n_14023);
  not g30950 (n_14024, n19884);
  and g30951 (n19886, n_14024, n19885);
  not g30952 (n_14025, n19876);
  not g30953 (n_14026, n19886);
  and g30954 (n19887, n_14025, n_14026);
  not g30955 (n_14027, n19887);
  and g30956 (n19888, pi0790, n_14027);
  not g30957 (n_14028, n19859);
  and g30958 (n19889, pi0832, n_14028);
  not g30959 (n_14029, n19888);
  and g30960 (n19890, n_14029, n19889);
  not g30961 (n_14030, n19682);
  not g30962 (n_14031, n19890);
  and g30963 (po0300, n_14030, n_14031);
  and g30964 (n19892, pi0144, n_11751);
  not g30965 (n_14032, n19892);
  and g30966 (n19893, n16635, n_14032);
  and g30967 (n19894, n17075, n_14032);
  and g30968 (n19895, pi0736, n2571);
  not g30969 (n_14034, n19895);
  and g30970 (n19896, n_14032, n_14034);
  and g30971 (n19897, n_298, n_11418);
  and g30972 (n19898, n16641, n_11501);
  not g30973 (n_14035, n19898);
  and g30974 (n19899, pi0038, n_14035);
  not g30975 (n_14036, n19897);
  and g30976 (n19900, n_14036, n19899);
  and g30977 (n19901, n_298, n18076);
  not g30978 (n_14037, n18072);
  and g30979 (n19902, pi0144, n_14037);
  not g30980 (n_14038, n19901);
  and g30981 (n19903, n_161, n_14038);
  not g30982 (n_14039, n19902);
  and g30983 (n19904, n_14039, n19903);
  not g30984 (n_14040, n19900);
  and g30985 (n19905, n19895, n_14040);
  not g30986 (n_14041, n19904);
  and g30987 (n19906, n_14041, n19905);
  not g30988 (n_14042, n19896);
  not g30989 (n_14043, n19906);
  and g30990 (n19907, n_14042, n_14043);
  and g30991 (n19908, n_11749, n19907);
  and g30992 (n19909, n_11753, n_14032);
  not g30993 (n_14044, n19907);
  and g30994 (n19910, pi0625, n_14044);
  not g30995 (n_14045, n19909);
  and g30996 (n19911, pi1153, n_14045);
  not g30997 (n_14046, n19910);
  and g30998 (n19912, n_14046, n19911);
  and g30999 (n19913, n_11753, n_14044);
  and g31000 (n19914, pi0625, n_14032);
  not g31001 (n_14047, n19914);
  and g31002 (n19915, n_11757, n_14047);
  not g31003 (n_14048, n19913);
  and g31004 (n19916, n_14048, n19915);
  not g31005 (n_14049, n19912);
  not g31006 (n_14050, n19916);
  and g31007 (n19917, n_14049, n_14050);
  not g31008 (n_14051, n19917);
  and g31009 (n19918, pi0778, n_14051);
  not g31010 (n_14052, n19908);
  not g31011 (n_14053, n19918);
  and g31012 (n19919, n_14052, n_14053);
  and g31013 (n19920, n_11773, n19919);
  not g31014 (n_14054, n19894);
  not g31015 (n_14055, n19920);
  and g31016 (n19921, n_14054, n_14055);
  and g31017 (n19922, n_11777, n19921);
  and g31018 (n19923, n16639, n19892);
  not g31019 (n_14056, n19922);
  not g31020 (n_14057, n19923);
  and g31021 (n19924, n_14056, n_14057);
  and g31022 (n19925, n_11780, n19924);
  not g31023 (n_14058, n19893);
  not g31024 (n_14059, n19925);
  and g31025 (n19926, n_14058, n_14059);
  and g31026 (n19927, n_11783, n19926);
  and g31027 (n19928, n16631, n19892);
  not g31028 (n_14060, n19927);
  not g31029 (n_14061, n19928);
  and g31030 (n19929, n_14060, n_14061);
  not g31031 (n_14062, n19929);
  and g31032 (n19930, n_11787, n_14062);
  and g31033 (n19931, n_11789, n_14032);
  and g31034 (n19932, pi0628, n19929);
  not g31035 (n_14063, n19931);
  and g31036 (n19933, pi1156, n_14063);
  not g31037 (n_14064, n19932);
  and g31038 (n19934, n_14064, n19933);
  and g31039 (n19935, pi0628, n_14032);
  and g31040 (n19936, n_11789, n19929);
  not g31041 (n_14065, n19935);
  and g31042 (n19937, n_11794, n_14065);
  not g31043 (n_14066, n19936);
  and g31044 (n19938, n_14066, n19937);
  not g31045 (n_14067, n19934);
  not g31046 (n_14068, n19938);
  and g31047 (n19939, n_14067, n_14068);
  not g31048 (n_14069, n19939);
  and g31049 (n19940, pi0792, n_14069);
  not g31050 (n_14070, n19930);
  not g31051 (n_14071, n19940);
  and g31052 (n19941, n_14070, n_14071);
  not g31053 (n_14072, n19941);
  and g31054 (n19942, n_11803, n_14072);
  and g31055 (n19943, n_11806, n_14032);
  and g31056 (n19944, pi0647, n19941);
  not g31057 (n_14073, n19943);
  and g31058 (n19945, pi1157, n_14073);
  not g31059 (n_14074, n19944);
  and g31060 (n19946, n_14074, n19945);
  and g31061 (n19947, pi0647, n_14032);
  and g31062 (n19948, n_11806, n19941);
  not g31063 (n_14075, n19947);
  and g31064 (n19949, n_11810, n_14075);
  not g31065 (n_14076, n19948);
  and g31066 (n19950, n_14076, n19949);
  not g31067 (n_14077, n19946);
  not g31068 (n_14078, n19950);
  and g31069 (n19951, n_14077, n_14078);
  not g31070 (n_14079, n19951);
  and g31071 (n19952, pi0787, n_14079);
  not g31072 (n_14080, n19942);
  not g31073 (n_14081, n19952);
  and g31074 (n19953, n_14080, n_14081);
  and g31075 (n19954, n_11819, n19953);
  and g31076 (n19955, n_11821, n_14032);
  and g31077 (n19956, n17117, n_14032);
  and g31078 (n19957, pi0144, n_11417);
  not g31079 (n_14083, pi0758);
  and g31080 (n19958, n_14083, n_11736);
  and g31081 (n19959, pi0758, n17219);
  not g31082 (n_14084, n19958);
  not g31083 (n_14085, n19959);
  and g31084 (n19960, n_14084, n_14085);
  not g31085 (n_14086, n19960);
  and g31086 (n19961, pi0039, n_14086);
  and g31087 (n19962, n_14083, n16958);
  and g31088 (n19963, pi0758, n17139);
  not g31089 (n_14087, n19962);
  and g31090 (n19964, n_162, n_14087);
  not g31091 (n_14088, n19963);
  and g31092 (n19965, n_14088, n19964);
  not g31093 (n_14089, n19961);
  not g31094 (n_14090, n19965);
  and g31095 (n19966, n_14089, n_14090);
  not g31096 (n_14091, n19966);
  and g31097 (n19967, pi0144, n_14091);
  and g31098 (n19968, n_298, pi0758);
  and g31099 (n19969, n17275, n19968);
  not g31100 (n_14092, n19967);
  not g31101 (n_14093, n19969);
  and g31102 (n19970, n_14092, n_14093);
  not g31103 (n_14094, n19970);
  and g31104 (n19971, n_161, n_14094);
  and g31105 (n19972, pi0758, n17168);
  not g31106 (n_14095, n19972);
  and g31107 (n19973, n16641, n_14095);
  and g31108 (n19974, pi0038, n_14036);
  not g31109 (n_14096, n19973);
  and g31110 (n19975, n_14096, n19974);
  not g31111 (n_14097, n19971);
  not g31112 (n_14098, n19975);
  and g31113 (n19976, n_14097, n_14098);
  not g31114 (n_14099, n19976);
  and g31115 (n19977, n2571, n_14099);
  not g31116 (n_14100, n19957);
  not g31117 (n_14101, n19977);
  and g31118 (n19978, n_14100, n_14101);
  and g31119 (n19979, n_11960, n19978);
  not g31120 (n_14102, n19956);
  not g31121 (n_14103, n19979);
  and g31122 (n19980, n_14102, n_14103);
  and g31123 (n19981, n_11964, n19980);
  and g31124 (n19982, n_11971, n_14032);
  not g31125 (n_14104, n19980);
  and g31126 (n19983, pi0609, n_14104);
  not g31127 (n_14105, n19982);
  and g31128 (n19984, pi1155, n_14105);
  not g31129 (n_14106, n19983);
  and g31130 (n19985, n_14106, n19984);
  and g31131 (n19986, n_11971, n_14104);
  and g31132 (n19987, pi0609, n_14032);
  not g31133 (n_14107, n19987);
  and g31134 (n19988, n_11768, n_14107);
  not g31135 (n_14108, n19986);
  and g31136 (n19989, n_14108, n19988);
  not g31137 (n_14109, n19985);
  not g31138 (n_14110, n19989);
  and g31139 (n19990, n_14109, n_14110);
  not g31140 (n_14111, n19990);
  and g31141 (n19991, pi0785, n_14111);
  not g31142 (n_14112, n19981);
  not g31143 (n_14113, n19991);
  and g31144 (n19992, n_14112, n_14113);
  not g31145 (n_14114, n19992);
  and g31146 (n19993, n_11981, n_14114);
  and g31147 (n19994, n_11984, n_14032);
  and g31148 (n19995, pi0618, n19992);
  not g31149 (n_14115, n19994);
  and g31150 (n19996, pi1154, n_14115);
  not g31151 (n_14116, n19995);
  and g31152 (n19997, n_14116, n19996);
  and g31153 (n19998, pi0618, n_14032);
  and g31154 (n19999, n_11984, n19992);
  not g31155 (n_14117, n19998);
  and g31156 (n20000, n_11413, n_14117);
  not g31157 (n_14118, n19999);
  and g31158 (n20001, n_14118, n20000);
  not g31159 (n_14119, n19997);
  not g31160 (n_14120, n20001);
  and g31161 (n20002, n_14119, n_14120);
  not g31162 (n_14121, n20002);
  and g31163 (n20003, pi0781, n_14121);
  not g31164 (n_14122, n19993);
  not g31165 (n_14123, n20003);
  and g31166 (n20004, n_14122, n_14123);
  and g31167 (n20005, pi0619, n20004);
  not g31168 (n_14124, n19955);
  and g31169 (n20006, pi1159, n_14124);
  not g31170 (n_14125, n20005);
  and g31171 (n20007, n_14125, n20006);
  not g31172 (n_14126, pi0736);
  and g31173 (n20008, n_14126, n19976);
  and g31174 (n20009, n_298, n_13720);
  and g31175 (n20010, pi0144, n17546);
  not g31176 (n_14127, n20010);
  and g31177 (n20011, pi0758, n_14127);
  not g31178 (n_14128, n20009);
  and g31179 (n20012, n_14128, n20011);
  and g31180 (n20013, pi0144, n_13705);
  and g31181 (n20014, n_298, n_13702);
  not g31182 (n_14129, n20014);
  and g31183 (n20015, n_14083, n_14129);
  not g31184 (n_14130, n20013);
  and g31185 (n20016, n_14130, n20015);
  not g31186 (n_14131, n20012);
  and g31187 (n20017, pi0039, n_14131);
  not g31188 (n_14132, n20016);
  and g31189 (n20018, n_14132, n20017);
  and g31190 (n20019, n_298, n17631);
  and g31191 (n20020, pi0144, n17629);
  not g31192 (n_14133, n20019);
  and g31193 (n20021, pi0758, n_14133);
  not g31194 (n_14134, n20020);
  and g31195 (n20022, n_14134, n20021);
  and g31196 (n20023, n_298, n_12240);
  and g31197 (n20024, pi0144, n_12230);
  not g31198 (n_14135, n20023);
  and g31199 (n20025, n_14083, n_14135);
  not g31200 (n_14136, n20024);
  and g31201 (n20026, n_14136, n20025);
  not g31202 (n_14137, n20022);
  and g31203 (n20027, n_162, n_14137);
  not g31204 (n_14138, n20026);
  and g31205 (n20028, n_14138, n20027);
  not g31206 (n_14139, n20028);
  and g31207 (n20029, n_161, n_14139);
  not g31208 (n_14140, n20018);
  and g31209 (n20030, n_14140, n20029);
  not g31214 (n_14142, n20033);
  and g31215 (n20034, n2571, n_14142);
  not g31216 (n_14143, n20008);
  and g31217 (n20035, n_14143, n20034);
  not g31218 (n_14144, n20035);
  and g31219 (n20036, n_14100, n_14144);
  and g31220 (n20037, n_11753, n20036);
  and g31221 (n20038, pi0625, n19978);
  not g31222 (n_14145, n20038);
  and g31223 (n20039, n_11757, n_14145);
  not g31224 (n_14146, n20037);
  and g31225 (n20040, n_14146, n20039);
  and g31226 (n20041, n_11823, n_14049);
  not g31227 (n_14147, n20040);
  and g31228 (n20042, n_14147, n20041);
  and g31229 (n20043, n_11753, n19978);
  and g31230 (n20044, pi0625, n20036);
  not g31231 (n_14148, n20043);
  and g31232 (n20045, pi1153, n_14148);
  not g31233 (n_14149, n20044);
  and g31234 (n20046, n_14149, n20045);
  and g31235 (n20047, pi0608, n_14050);
  not g31236 (n_14150, n20046);
  and g31237 (n20048, n_14150, n20047);
  not g31238 (n_14151, n20042);
  not g31239 (n_14152, n20048);
  and g31240 (n20049, n_14151, n_14152);
  not g31241 (n_14153, n20049);
  and g31242 (n20050, pi0778, n_14153);
  and g31243 (n20051, n_11749, n20036);
  not g31244 (n_14154, n20050);
  not g31245 (n_14155, n20051);
  and g31246 (n20052, n_14154, n_14155);
  not g31247 (n_14156, n20052);
  and g31248 (n20053, n_11971, n_14156);
  and g31249 (n20054, pi0609, n19919);
  not g31250 (n_14157, n20054);
  and g31251 (n20055, n_11768, n_14157);
  not g31252 (n_14158, n20053);
  and g31253 (n20056, n_14158, n20055);
  and g31254 (n20057, n_11767, n_14109);
  not g31255 (n_14159, n20056);
  and g31256 (n20058, n_14159, n20057);
  and g31257 (n20059, n_11971, n19919);
  and g31258 (n20060, pi0609, n_14156);
  not g31259 (n_14160, n20059);
  and g31260 (n20061, pi1155, n_14160);
  not g31261 (n_14161, n20060);
  and g31262 (n20062, n_14161, n20061);
  and g31263 (n20063, pi0660, n_14110);
  not g31264 (n_14162, n20062);
  and g31265 (n20064, n_14162, n20063);
  not g31266 (n_14163, n20058);
  not g31267 (n_14164, n20064);
  and g31268 (n20065, n_14163, n_14164);
  not g31269 (n_14165, n20065);
  and g31270 (n20066, pi0785, n_14165);
  and g31271 (n20067, n_11964, n_14156);
  not g31272 (n_14166, n20066);
  not g31273 (n_14167, n20067);
  and g31274 (n20068, n_14166, n_14167);
  not g31275 (n_14168, n20068);
  and g31276 (n20069, n_11984, n_14168);
  not g31277 (n_14169, n19921);
  and g31278 (n20070, pi0618, n_14169);
  not g31279 (n_14170, n20070);
  and g31280 (n20071, n_11413, n_14170);
  not g31281 (n_14171, n20069);
  and g31282 (n20072, n_14171, n20071);
  and g31283 (n20073, n_11412, n_14119);
  not g31284 (n_14172, n20072);
  and g31285 (n20074, n_14172, n20073);
  and g31286 (n20075, pi0618, n_14168);
  and g31287 (n20076, n_11984, n_14169);
  not g31288 (n_14173, n20076);
  and g31289 (n20077, pi1154, n_14173);
  not g31290 (n_14174, n20075);
  and g31291 (n20078, n_14174, n20077);
  and g31292 (n20079, pi0627, n_14120);
  not g31293 (n_14175, n20078);
  and g31294 (n20080, n_14175, n20079);
  not g31295 (n_14176, n20074);
  not g31296 (n_14177, n20080);
  and g31297 (n20081, n_14176, n_14177);
  not g31298 (n_14178, n20081);
  and g31299 (n20082, pi0781, n_14178);
  and g31300 (n20083, n_11981, n_14168);
  not g31301 (n_14179, n20082);
  not g31302 (n_14180, n20083);
  and g31303 (n20084, n_14179, n_14180);
  not g31304 (n_14181, n20084);
  and g31305 (n20085, n_11821, n_14181);
  and g31306 (n20086, pi0619, n19924);
  not g31307 (n_14182, n20086);
  and g31308 (n20087, n_11405, n_14182);
  not g31309 (n_14183, n20085);
  and g31310 (n20088, n_14183, n20087);
  not g31311 (n_14184, n20007);
  and g31312 (n20089, n_11403, n_14184);
  not g31313 (n_14185, n20088);
  and g31314 (n20090, n_14185, n20089);
  and g31315 (n20091, pi0619, n_14032);
  and g31316 (n20092, n_11821, n20004);
  not g31317 (n_14186, n20091);
  and g31318 (n20093, n_11405, n_14186);
  not g31319 (n_14187, n20092);
  and g31320 (n20094, n_14187, n20093);
  and g31321 (n20095, n_11821, n19924);
  and g31322 (n20096, pi0619, n_14181);
  not g31323 (n_14188, n20095);
  and g31324 (n20097, pi1159, n_14188);
  not g31325 (n_14189, n20096);
  and g31326 (n20098, n_14189, n20097);
  not g31327 (n_14190, n20094);
  and g31328 (n20099, pi0648, n_14190);
  not g31329 (n_14191, n20098);
  and g31330 (n20100, n_14191, n20099);
  not g31331 (n_14192, n20090);
  not g31332 (n_14193, n20100);
  and g31333 (n20101, n_14192, n_14193);
  not g31334 (n_14194, n20101);
  and g31335 (n20102, pi0789, n_14194);
  and g31336 (n20103, n_12315, n_14181);
  not g31337 (n_14195, n20102);
  not g31338 (n_14196, n20103);
  and g31339 (n20104, n_14195, n_14196);
  and g31340 (n20105, n_12318, n20104);
  and g31341 (n20106, n_12320, n20104);
  and g31342 (n20107, pi0626, n19926);
  not g31343 (n_14197, n20107);
  and g31344 (n20108, n_11395, n_14197);
  not g31345 (n_14198, n20106);
  and g31346 (n20109, n_14198, n20108);
  not g31347 (n_14199, n20004);
  and g31348 (n20110, n_12315, n_14199);
  and g31349 (n20111, n_14184, n_14190);
  not g31350 (n_14200, n20111);
  and g31351 (n20112, pi0789, n_14200);
  not g31352 (n_14201, n20110);
  not g31353 (n_14202, n20112);
  and g31354 (n20113, n_14201, n_14202);
  and g31355 (n20114, n_12320, n20113);
  and g31356 (n20115, pi0626, n_14032);
  not g31357 (n_14203, n20115);
  and g31358 (n20116, n_11397, n_14203);
  not g31359 (n_14204, n20114);
  and g31360 (n20117, n_14204, n20116);
  not g31361 (n_14205, n20117);
  and g31362 (n20118, n_12330, n_14205);
  not g31363 (n_14206, n20109);
  not g31364 (n_14207, n20118);
  and g31365 (n20119, n_14206, n_14207);
  and g31366 (n20120, pi0626, n20104);
  and g31367 (n20121, n_12320, n19926);
  not g31368 (n_14208, n20121);
  and g31369 (n20122, pi0641, n_14208);
  not g31370 (n_14209, n20120);
  and g31371 (n20123, n_14209, n20122);
  and g31372 (n20124, pi0626, n20113);
  and g31373 (n20125, n_12320, n_14032);
  not g31374 (n_14210, n20125);
  and g31375 (n20126, pi1158, n_14210);
  not g31376 (n_14211, n20124);
  and g31377 (n20127, n_14211, n20126);
  not g31378 (n_14212, n20127);
  and g31379 (n20128, n_12338, n_14212);
  not g31380 (n_14213, n20123);
  not g31381 (n_14214, n20128);
  and g31382 (n20129, n_14213, n_14214);
  not g31383 (n_14215, n20119);
  not g31384 (n_14216, n20129);
  and g31385 (n20130, n_14215, n_14216);
  not g31386 (n_14217, n20130);
  and g31387 (n20131, pi0788, n_14217);
  not g31388 (n_14218, n20105);
  not g31389 (n_14219, n20131);
  and g31390 (n20132, n_14218, n_14219);
  and g31391 (n20133, n_11789, n20132);
  and g31392 (n20134, n_14205, n_14212);
  not g31393 (n_14220, n20134);
  and g31394 (n20135, pi0788, n_14220);
  not g31395 (n_14221, n20113);
  and g31396 (n20136, n_12318, n_14221);
  not g31397 (n_14222, n20135);
  not g31398 (n_14223, n20136);
  and g31399 (n20137, n_14222, n_14223);
  and g31400 (n20138, pi0628, n20137);
  not g31401 (n_14224, n20138);
  and g31402 (n20139, n_11794, n_14224);
  not g31403 (n_14225, n20133);
  and g31404 (n20140, n_14225, n20139);
  and g31405 (n20141, n_12354, n_14067);
  not g31406 (n_14226, n20140);
  and g31407 (n20142, n_14226, n20141);
  and g31408 (n20143, pi0628, n20132);
  and g31409 (n20144, n_11789, n20137);
  not g31410 (n_14227, n20144);
  and g31411 (n20145, pi1156, n_14227);
  not g31412 (n_14228, n20143);
  and g31413 (n20146, n_14228, n20145);
  and g31414 (n20147, pi0629, n_14068);
  not g31415 (n_14229, n20146);
  and g31416 (n20148, n_14229, n20147);
  not g31417 (n_14230, n20142);
  not g31418 (n_14231, n20148);
  and g31419 (n20149, n_14230, n_14231);
  not g31420 (n_14232, n20149);
  and g31421 (n20150, pi0792, n_14232);
  and g31422 (n20151, n_11787, n20132);
  not g31423 (n_14233, n20150);
  not g31424 (n_14234, n20151);
  and g31425 (n20152, n_14233, n_14234);
  not g31426 (n_14235, n20152);
  and g31427 (n20153, n_11806, n_14235);
  not g31428 (n_14236, n20137);
  and g31429 (n20154, n_12368, n_14236);
  and g31430 (n20155, n17779, n19892);
  not g31431 (n_14237, n20154);
  not g31432 (n_14238, n20155);
  and g31433 (n20156, n_14237, n_14238);
  and g31434 (n20157, pi0647, n20156);
  not g31435 (n_14239, n20157);
  and g31436 (n20158, n_11810, n_14239);
  not g31437 (n_14240, n20153);
  and g31438 (n20159, n_14240, n20158);
  and g31439 (n20160, n_12375, n_14077);
  not g31440 (n_14241, n20159);
  and g31441 (n20161, n_14241, n20160);
  and g31442 (n20162, pi0647, n_14235);
  and g31443 (n20163, n_11806, n20156);
  not g31444 (n_14242, n20163);
  and g31445 (n20164, pi1157, n_14242);
  not g31446 (n_14243, n20162);
  and g31447 (n20165, n_14243, n20164);
  and g31448 (n20166, pi0630, n_14078);
  not g31449 (n_14244, n20165);
  and g31450 (n20167, n_14244, n20166);
  not g31451 (n_14245, n20161);
  not g31452 (n_14246, n20167);
  and g31453 (n20168, n_14245, n_14246);
  not g31454 (n_14247, n20168);
  and g31455 (n20169, pi0787, n_14247);
  and g31456 (n20170, n_11803, n_14235);
  not g31457 (n_14248, n20169);
  not g31458 (n_14249, n20170);
  and g31459 (n20171, n_14248, n_14249);
  not g31460 (n_14250, n20171);
  and g31461 (n20172, pi0644, n_14250);
  not g31462 (n_14251, n19954);
  and g31463 (n20173, pi0715, n_14251);
  not g31464 (n_14252, n20172);
  and g31465 (n20174, n_14252, n20173);
  and g31466 (n20175, n17804, n_14032);
  and g31467 (n20176, n_12392, n20156);
  not g31468 (n_14253, n20175);
  not g31469 (n_14254, n20176);
  and g31470 (n20177, n_14253, n_14254);
  not g31471 (n_14255, n20177);
  and g31472 (n20178, pi0644, n_14255);
  and g31473 (n20179, n_11819, n_14032);
  not g31474 (n_14256, n20179);
  and g31475 (n20180, n_12395, n_14256);
  not g31476 (n_14257, n20178);
  and g31477 (n20181, n_14257, n20180);
  not g31478 (n_14258, n20181);
  and g31479 (n20182, pi1160, n_14258);
  not g31480 (n_14259, n20174);
  and g31481 (n20183, n_14259, n20182);
  and g31482 (n20184, n_11819, n_14250);
  and g31483 (n20185, pi0644, n19953);
  not g31484 (n_14260, n20185);
  and g31485 (n20186, n_12395, n_14260);
  not g31486 (n_14261, n20184);
  and g31487 (n20187, n_14261, n20186);
  and g31488 (n20188, n_11819, n_14255);
  and g31489 (n20189, pi0644, n_14032);
  not g31490 (n_14262, n20189);
  and g31491 (n20190, pi0715, n_14262);
  not g31492 (n_14263, n20188);
  and g31493 (n20191, n_14263, n20190);
  not g31494 (n_14264, n20191);
  and g31495 (n20192, n_12405, n_14264);
  not g31496 (n_14265, n20187);
  and g31497 (n20193, n_14265, n20192);
  not g31498 (n_14266, n20183);
  and g31499 (n20194, pi0790, n_14266);
  not g31500 (n_14267, n20193);
  and g31501 (n20195, n_14267, n20194);
  and g31502 (n20196, n_12411, n20171);
  not g31503 (n_14268, n20196);
  and g31504 (n20197, n6305, n_14268);
  not g31505 (n_14269, n20195);
  and g31506 (n20198, n_14269, n20197);
  and g31507 (n20199, n_298, n_3232);
  not g31508 (n_14270, n20199);
  and g31509 (n20200, n_796, n_14270);
  not g31510 (n_14271, n20198);
  and g31511 (n20201, n_14271, n20200);
  and g31512 (n20202, pi0057, pi0144);
  not g31513 (n_14272, n20202);
  and g31514 (n20203, n_12415, n_14272);
  not g31515 (n_14273, n20201);
  and g31516 (n20204, n_14273, n20203);
  and g31517 (n20205, n17803, n19341);
  not g31518 (n_14274, n20205);
  and g31519 (n20206, pi0787, n_14274);
  and g31520 (n20207, pi0144, n_12418);
  and g31521 (n20208, pi0736, n16645);
  not g31522 (n_14275, n20207);
  not g31523 (n_14276, n20208);
  and g31524 (n20209, n_14275, n_14276);
  and g31525 (n20210, n_11749, n20209);
  and g31526 (n20211, pi0625, n20208);
  not g31527 (n_14277, n20209);
  not g31528 (n_14278, n20211);
  and g31529 (n20212, n_14277, n_14278);
  not g31530 (n_14279, n20212);
  and g31531 (n20213, n_11757, n_14279);
  and g31532 (n20214, pi1153, n_14275);
  and g31533 (n20215, n_14278, n20214);
  not g31534 (n_14280, n20213);
  not g31535 (n_14281, n20215);
  and g31536 (n20216, n_14280, n_14281);
  not g31537 (n_14282, n20216);
  and g31538 (n20217, pi0778, n_14282);
  not g31539 (n_14283, n20210);
  not g31540 (n_14284, n20217);
  and g31541 (n20218, n_14283, n_14284);
  and g31542 (n20219, n19151, n20218);
  and g31543 (n20220, n_11789, n20219);
  not g31544 (n_14285, n20220);
  and g31545 (n20221, pi0629, n_14285);
  and g31546 (n20222, n_11971, n_11768);
  and g31547 (n20223, pi0609, pi1155);
  not g31548 (n_14286, n20222);
  and g31549 (n20224, pi0785, n_14286);
  not g31550 (n_14287, n20223);
  and g31551 (n20225, n_14287, n20224);
  and g31552 (n20226, pi0758, n17244);
  not g31553 (n_14288, n20225);
  and g31554 (n20227, n_14288, n20226);
  and g31555 (n20228, n_11821, pi1159);
  and g31556 (n20229, pi0619, n_11405);
  not g31557 (n_14289, n20228);
  not g31558 (n_14290, n20229);
  and g31559 (n20230, n_14289, n_14290);
  not g31560 (n_14291, n20230);
  and g31561 (n20231, pi0789, n_14291);
  and g31562 (n20232, n_11984, n_11413);
  and g31563 (n20233, pi0618, pi1154);
  not g31564 (n_14292, n20232);
  and g31565 (n20234, pi0781, n_14292);
  not g31566 (n_14293, n20233);
  and g31567 (n20235, n_14293, n20234);
  not g31568 (n_14294, n20231);
  and g31569 (n20236, n_11960, n_14294);
  not g31570 (n_14295, n20235);
  and g31571 (n20237, n_14295, n20236);
  and g31572 (n20238, n20227, n20237);
  and g31573 (n20239, n_12524, n20238);
  not g31574 (n_14296, n20239);
  and g31575 (n20240, pi0628, n_14296);
  not g31576 (n_14297, n20221);
  not g31577 (n_14298, n20240);
  and g31578 (n20241, n_14297, n_14298);
  not g31579 (n_14299, n20241);
  and g31580 (n20242, n_11794, n_14299);
  and g31581 (n20243, pi0628, n20219);
  and g31582 (n20244, n_11789, n_14296);
  not g31583 (n_14300, n20244);
  and g31584 (n20245, pi0629, n_14300);
  not g31585 (n_14301, n20245);
  and g31586 (n20246, pi1156, n_14301);
  not g31587 (n_14302, n20243);
  and g31588 (n20247, n_14302, n20246);
  not g31589 (n_14303, n20242);
  not g31590 (n_14304, n20247);
  and g31591 (n20248, n_14303, n_14304);
  not g31592 (n_14305, n20248);
  and g31593 (n20249, n_14275, n_14305);
  and g31594 (n20250, pi0792, n20249);
  and g31595 (n20251, n16635, n_14275);
  and g31596 (n20252, n_11773, n20218);
  and g31597 (n20253, n_11777, n20252);
  not g31598 (n_14306, n20253);
  and g31599 (n20254, n_14275, n_14306);
  not g31600 (n_14307, n20251);
  not g31601 (n_14308, n20254);
  and g31602 (n20255, n_14307, n_14308);
  and g31603 (n20256, n17865, n20255);
  and g31604 (n20257, n_12320, n20238);
  not g31605 (n_14309, n20257);
  and g31606 (n20258, n_14275, n_14309);
  not g31607 (n_14310, n20258);
  and g31608 (n20259, n_11397, n_14310);
  not g31609 (n_14311, n20259);
  and g31610 (n20260, pi0641, n_14311);
  not g31611 (n_14312, n20256);
  and g31612 (n20261, n_14312, n20260);
  and g31613 (n20262, pi0626, n20238);
  not g31614 (n_14313, n20262);
  and g31615 (n20263, n_14275, n_14313);
  not g31616 (n_14314, n20263);
  and g31617 (n20264, pi1158, n_14314);
  and g31618 (n20265, n17866, n20255);
  not g31619 (n_14315, n20264);
  and g31620 (n20266, n_11395, n_14315);
  not g31621 (n_14316, n20265);
  and g31622 (n20267, n_14316, n20266);
  not g31623 (n_14317, n20261);
  and g31624 (n20268, pi0788, n_14317);
  not g31625 (n_14318, n20267);
  and g31626 (n20269, n_14318, n20268);
  and g31627 (n20270, pi0618, n_11960);
  and g31628 (n20271, n20227, n20270);
  and g31629 (n20272, pi1154, n_14275);
  not g31630 (n_14319, n20271);
  and g31631 (n20273, n_14319, n20272);
  not g31632 (n_14320, n20252);
  and g31633 (n20274, n_14275, n_14320);
  not g31634 (n_14321, n20274);
  and g31635 (n20275, pi0618, n_14321);
  and g31636 (n20276, n17291, n20226);
  and g31637 (n20277, pi1155, n_14275);
  not g31638 (n_14322, n20276);
  and g31639 (n20278, n_14322, n20277);
  and g31640 (n20279, pi0609, n20218);
  not g31641 (n_14323, n20226);
  and g31642 (n20280, n_14275, n_14323);
  and g31643 (n20281, pi0736, n17469);
  not g31644 (n_14324, n20281);
  and g31645 (n20282, n20280, n_14324);
  and g31646 (n20283, pi0625, n20281);
  not g31647 (n_14325, n20282);
  not g31648 (n_14326, n20283);
  and g31649 (n20284, n_14325, n_14326);
  not g31650 (n_14327, n20284);
  and g31651 (n20285, n_11757, n_14327);
  and g31652 (n20286, n_11823, n_14281);
  not g31653 (n_14328, n20285);
  and g31654 (n20287, n_14328, n20286);
  and g31655 (n20288, pi1153, n20280);
  and g31656 (n20289, n_14326, n20288);
  and g31657 (n20290, pi0608, n_14280);
  not g31658 (n_14329, n20289);
  and g31659 (n20291, n_14329, n20290);
  not g31660 (n_14330, n20287);
  not g31661 (n_14331, n20291);
  and g31662 (n20292, n_14330, n_14331);
  not g31663 (n_14332, n20292);
  and g31664 (n20293, pi0778, n_14332);
  and g31665 (n20294, n_11749, n_14325);
  not g31666 (n_14333, n20293);
  not g31667 (n_14334, n20294);
  and g31668 (n20295, n_14333, n_14334);
  not g31669 (n_14335, n20295);
  and g31670 (n20296, n_11971, n_14335);
  not g31671 (n_14336, n20279);
  and g31672 (n20297, n_11768, n_14336);
  not g31673 (n_14337, n20296);
  and g31674 (n20298, n_14337, n20297);
  not g31675 (n_14338, n20278);
  and g31676 (n20299, n_11767, n_14338);
  not g31677 (n_14339, n20298);
  and g31678 (n20300, n_14339, n20299);
  and g31679 (n20301, n17296, n20226);
  and g31680 (n20302, n_11768, n_14275);
  not g31681 (n_14340, n20301);
  and g31682 (n20303, n_14340, n20302);
  and g31683 (n20304, n_11971, n20218);
  and g31684 (n20305, pi0609, n_14335);
  not g31685 (n_14341, n20304);
  and g31686 (n20306, pi1155, n_14341);
  not g31687 (n_14342, n20305);
  and g31688 (n20307, n_14342, n20306);
  not g31689 (n_14343, n20303);
  and g31690 (n20308, pi0660, n_14343);
  not g31691 (n_14344, n20307);
  and g31692 (n20309, n_14344, n20308);
  not g31693 (n_14345, n20300);
  not g31694 (n_14346, n20309);
  and g31695 (n20310, n_14345, n_14346);
  not g31696 (n_14347, n20310);
  and g31697 (n20311, pi0785, n_14347);
  and g31698 (n20312, n_11964, n_14335);
  not g31699 (n_14348, n20311);
  not g31700 (n_14349, n20312);
  and g31701 (n20313, n_14348, n_14349);
  not g31702 (n_14350, n20313);
  and g31703 (n20314, n_11984, n_14350);
  not g31704 (n_14351, n20275);
  and g31705 (n20315, n_11413, n_14351);
  not g31706 (n_14352, n20314);
  and g31707 (n20316, n_14352, n20315);
  not g31708 (n_14353, n20273);
  and g31709 (n20317, n_11412, n_14353);
  not g31710 (n_14354, n20316);
  and g31711 (n20318, n_14354, n20317);
  and g31712 (n20319, n_11984, n_11960);
  and g31713 (n20320, n20227, n20319);
  and g31714 (n20321, n_11413, n_14275);
  not g31715 (n_14355, n20320);
  and g31716 (n20322, n_14355, n20321);
  and g31717 (n20323, n_11984, n_14321);
  and g31718 (n20324, pi0618, n_14350);
  not g31719 (n_14356, n20323);
  and g31720 (n20325, pi1154, n_14356);
  not g31721 (n_14357, n20324);
  and g31722 (n20326, n_14357, n20325);
  not g31723 (n_14358, n20322);
  and g31724 (n20327, pi0627, n_14358);
  not g31725 (n_14359, n20326);
  and g31726 (n20328, n_14359, n20327);
  not g31727 (n_14360, n20318);
  not g31728 (n_14361, n20328);
  and g31729 (n20329, n_14360, n_14361);
  not g31730 (n_14362, n20329);
  and g31731 (n20330, pi0781, n_14362);
  and g31732 (n20331, n_11981, n_14350);
  not g31733 (n_14363, n20330);
  not g31734 (n_14364, n20331);
  and g31735 (n20332, n_14363, n_14364);
  and g31736 (n20333, n_12315, n20332);
  and g31737 (n20334, n20227, n_14295);
  and g31738 (n20335, pi0619, n_11960);
  and g31739 (n20336, n20334, n20335);
  and g31740 (n20337, pi1159, n_14275);
  not g31741 (n_14365, n20336);
  and g31742 (n20338, n_14365, n20337);
  and g31743 (n20339, pi0619, n_14308);
  not g31744 (n_14366, n20332);
  and g31745 (n20340, n_11821, n_14366);
  not g31746 (n_14367, n20339);
  and g31747 (n20341, n_11405, n_14367);
  not g31748 (n_14368, n20340);
  and g31749 (n20342, n_14368, n20341);
  not g31750 (n_14369, n20338);
  and g31751 (n20343, n_11403, n_14369);
  not g31752 (n_14370, n20342);
  and g31753 (n20344, n_14370, n20343);
  and g31754 (n20345, n_11821, n_11960);
  and g31755 (n20346, n20334, n20345);
  and g31756 (n20347, n_11405, n_14275);
  not g31757 (n_14371, n20346);
  and g31758 (n20348, n_14371, n20347);
  and g31759 (n20349, n_11821, n_14308);
  and g31760 (n20350, pi0619, n_14366);
  not g31761 (n_14372, n20349);
  and g31762 (n20351, pi1159, n_14372);
  not g31763 (n_14373, n20350);
  and g31764 (n20352, n_14373, n20351);
  not g31765 (n_14374, n20348);
  and g31766 (n20353, pi0648, n_14374);
  not g31767 (n_14375, n20352);
  and g31768 (n20354, n_14375, n20353);
  not g31769 (n_14376, n20344);
  and g31770 (n20355, pi0789, n_14376);
  not g31771 (n_14377, n20354);
  and g31772 (n20356, n_14377, n20355);
  not g31773 (n_14378, n20333);
  and g31774 (n20357, n17970, n_14378);
  not g31775 (n_14379, n20356);
  and g31776 (n20358, n_14379, n20357);
  not g31777 (n_14380, n20269);
  not g31778 (n_14381, n20358);
  and g31779 (n20359, n_14380, n_14381);
  not g31780 (n_14382, n20250);
  not g31781 (n_14383, n20359);
  and g31782 (n20360, n_14382, n_14383);
  and g31783 (n20361, pi0629, n19139);
  and g31784 (n20362, n_12354, n19140);
  not g31785 (n_14384, n20361);
  and g31786 (n20363, pi0792, n_14384);
  not g31787 (n_14385, n20362);
  and g31788 (n20364, n_14385, n20363);
  not g31789 (n_14386, n20249);
  and g31790 (n20365, n_14386, n20364);
  not g31791 (n_14387, n20206);
  not g31792 (n_14388, n20365);
  and g31793 (n20366, n_14387, n_14388);
  not g31794 (n_14389, n20360);
  and g31795 (n20367, n_14389, n20366);
  and g31796 (n20368, n_12368, n20239);
  and g31797 (n20369, n_12375, n20368);
  not g31798 (n_14390, n20369);
  and g31799 (n20370, pi0647, n_14390);
  and g31800 (n20371, n_13453, n20219);
  not g31801 (n_14391, n20371);
  and g31802 (n20372, pi0630, n_14391);
  not g31803 (n_14392, n20370);
  not g31804 (n_14393, n20372);
  and g31805 (n20373, n_14392, n_14393);
  not g31806 (n_14394, n20373);
  and g31807 (n20374, n_11810, n_14394);
  and g31808 (n20375, pi0630, n20368);
  and g31809 (n20376, n_12375, n_14391);
  not g31810 (n_14395, n20376);
  and g31811 (n20377, pi0647, n_14395);
  not g31812 (n_14396, n20375);
  and g31813 (n20378, pi1157, n_14396);
  not g31814 (n_14397, n20377);
  and g31815 (n20379, n_14397, n20378);
  not g31816 (n_14398, n20374);
  not g31817 (n_14399, n20379);
  and g31818 (n20380, n_14398, n_14399);
  and g31819 (n20381, pi0787, n_14275);
  not g31820 (n_14400, n20380);
  and g31821 (n20382, n_14400, n20381);
  not g31822 (n_14401, n20367);
  not g31823 (n_14402, n20382);
  and g31824 (n20383, n_14401, n_14402);
  and g31825 (n20384, n_12411, n20383);
  and g31826 (n20385, n_12392, n20368);
  and g31827 (n20386, pi0644, n20385);
  and g31828 (n20387, n_12395, n_14275);
  not g31829 (n_14403, n20386);
  and g31830 (n20388, n_14403, n20387);
  and g31831 (n20389, n_13598, n20371);
  not g31832 (n_14404, n20389);
  and g31833 (n20390, n_14275, n_14404);
  not g31834 (n_14405, n20390);
  and g31835 (n20391, n_11819, n_14405);
  and g31836 (n20392, pi0644, n20383);
  not g31837 (n_14406, n20391);
  and g31838 (n20393, pi0715, n_14406);
  not g31839 (n_14407, n20392);
  and g31840 (n20394, n_14407, n20393);
  not g31841 (n_14408, n20388);
  and g31842 (n20395, pi1160, n_14408);
  not g31843 (n_14409, n20394);
  and g31844 (n20396, n_14409, n20395);
  and g31845 (n20397, n_11819, n20385);
  and g31846 (n20398, pi0715, n_14275);
  not g31847 (n_14410, n20397);
  and g31848 (n20399, n_14410, n20398);
  and g31849 (n20400, n_11819, n20383);
  and g31850 (n20401, pi0644, n_14405);
  not g31851 (n_14411, n20401);
  and g31852 (n20402, n_12395, n_14411);
  not g31853 (n_14412, n20400);
  and g31854 (n20403, n_14412, n20402);
  not g31855 (n_14413, n20399);
  and g31856 (n20404, n_12405, n_14413);
  not g31857 (n_14414, n20403);
  and g31858 (n20405, n_14414, n20404);
  not g31859 (n_14415, n20396);
  not g31860 (n_14416, n20405);
  and g31861 (n20406, n_14415, n_14416);
  not g31862 (n_14417, n20406);
  and g31863 (n20407, pi0790, n_14417);
  not g31864 (n_14418, n20384);
  and g31865 (n20408, pi0832, n_14418);
  not g31866 (n_14419, n20407);
  and g31867 (n20409, n_14419, n20408);
  not g31868 (n_14420, n20204);
  not g31869 (n_14421, n20409);
  and g31870 (po0301, n_14420, n_14421);
  and g31871 (n20411, n_6246, po1038);
  and g31872 (n20412, n_6246, n_11751);
  not g31873 (n_14422, n20412);
  and g31874 (n20413, n16635, n_14422);
  not g31875 (n_14424, pi0698);
  and g31876 (n20414, n_14424, n2571);
  not g31877 (n_14425, n20414);
  and g31878 (n20415, n20412, n_14425);
  and g31879 (n20416, n_6246, n_11418);
  not g31880 (n_14426, n20416);
  and g31881 (n20417, n16647, n_14426);
  and g31882 (n20418, pi0145, n_12608);
  not g31883 (n_14427, n20418);
  and g31884 (n20419, n_161, n_14427);
  not g31885 (n_14428, n20419);
  and g31886 (n20420, n2571, n_14428);
  and g31887 (n20421, n_6246, n18072);
  not g31888 (n_14429, n20420);
  not g31889 (n_14430, n20421);
  and g31890 (n20422, n_14429, n_14430);
  not g31891 (n_14431, n20417);
  and g31892 (n20423, n_14424, n_14431);
  not g31893 (n_14432, n20422);
  and g31894 (n20424, n_14432, n20423);
  not g31895 (n_14433, n20415);
  not g31896 (n_14434, n20424);
  and g31897 (n20425, n_14433, n_14434);
  and g31898 (n20426, n_11749, n20425);
  and g31899 (n20427, n_11753, n20412);
  not g31900 (n_14435, n20425);
  and g31901 (n20428, pi0625, n_14435);
  not g31902 (n_14436, n20427);
  and g31903 (n20429, pi1153, n_14436);
  not g31904 (n_14437, n20428);
  and g31905 (n20430, n_14437, n20429);
  and g31906 (n20431, pi0625, n20412);
  and g31907 (n20432, n_11753, n_14435);
  not g31908 (n_14438, n20431);
  and g31909 (n20433, n_11757, n_14438);
  not g31910 (n_14439, n20432);
  and g31911 (n20434, n_14439, n20433);
  not g31912 (n_14440, n20430);
  not g31913 (n_14441, n20434);
  and g31914 (n20435, n_14440, n_14441);
  not g31915 (n_14442, n20435);
  and g31916 (n20436, pi0778, n_14442);
  not g31917 (n_14443, n20426);
  not g31918 (n_14444, n20436);
  and g31919 (n20437, n_14443, n_14444);
  not g31920 (n_14445, n20437);
  and g31921 (n20438, n_11773, n_14445);
  and g31922 (n20439, n17075, n_14422);
  not g31923 (n_14446, n20438);
  not g31924 (n_14447, n20439);
  and g31925 (n20440, n_14446, n_14447);
  and g31926 (n20441, n_11777, n20440);
  and g31927 (n20442, n16639, n20412);
  not g31928 (n_14448, n20441);
  not g31929 (n_14449, n20442);
  and g31930 (n20443, n_14448, n_14449);
  and g31931 (n20444, n_11780, n20443);
  not g31932 (n_14450, n20413);
  not g31933 (n_14451, n20444);
  and g31934 (n20445, n_14450, n_14451);
  and g31935 (n20446, n_11783, n20445);
  and g31936 (n20447, n16631, n20412);
  not g31937 (n_14452, n20446);
  not g31938 (n_14453, n20447);
  and g31939 (n20448, n_14452, n_14453);
  and g31940 (n20449, n_11787, n20448);
  not g31941 (n_14454, n20448);
  and g31942 (n20450, pi0628, n_14454);
  and g31943 (n20451, n_11789, n20412);
  not g31944 (n_14455, n20451);
  and g31945 (n20452, pi1156, n_14455);
  not g31946 (n_14456, n20450);
  and g31947 (n20453, n_14456, n20452);
  and g31948 (n20454, pi0628, n20412);
  and g31949 (n20455, n_11789, n_14454);
  not g31950 (n_14457, n20454);
  and g31951 (n20456, n_11794, n_14457);
  not g31952 (n_14458, n20455);
  and g31953 (n20457, n_14458, n20456);
  not g31954 (n_14459, n20453);
  not g31955 (n_14460, n20457);
  and g31956 (n20458, n_14459, n_14460);
  not g31957 (n_14461, n20458);
  and g31958 (n20459, pi0792, n_14461);
  not g31959 (n_14462, n20449);
  not g31960 (n_14463, n20459);
  and g31961 (n20460, n_14462, n_14463);
  not g31962 (n_14464, n20460);
  and g31963 (n20461, n_11806, n_14464);
  and g31964 (n20462, pi0647, n_14422);
  not g31965 (n_14465, n20461);
  not g31966 (n_14466, n20462);
  and g31967 (n20463, n_14465, n_14466);
  and g31968 (n20464, n_11810, n20463);
  and g31969 (n20465, pi0647, n_14464);
  and g31970 (n20466, n_11806, n_14422);
  not g31971 (n_14467, n20465);
  not g31972 (n_14468, n20466);
  and g31973 (n20467, n_14467, n_14468);
  and g31974 (n20468, pi1157, n20467);
  not g31975 (n_14469, n20464);
  not g31976 (n_14470, n20468);
  and g31977 (n20469, n_14469, n_14470);
  not g31978 (n_14471, n20469);
  and g31979 (n20470, pi0787, n_14471);
  and g31980 (n20471, n_11803, n20460);
  not g31981 (n_14472, n20470);
  not g31982 (n_14473, n20471);
  and g31983 (n20472, n_14472, n_14473);
  not g31984 (n_14474, n20472);
  and g31985 (n20473, n_11819, n_14474);
  not g31986 (n_14475, n20473);
  and g31987 (n20474, pi0715, n_14475);
  and g31988 (n20475, pi0145, n_11417);
  not g31989 (n_14476, n17275);
  and g31990 (n20476, pi0145, n_14476);
  and g31991 (n20477, n_6246, n_11739);
  not g31992 (n_14478, n20477);
  and g31993 (n20478, pi0767, n_14478);
  not g31994 (n_14479, pi0767);
  and g31995 (n20479, n_6246, n_14479);
  and g31996 (n20480, n17221, n20479);
  not g31997 (n_14480, n20476);
  not g31998 (n_14481, n20480);
  and g31999 (n20481, n_14480, n_14481);
  not g32000 (n_14482, n20478);
  and g32001 (n20482, n_14482, n20481);
  not g32002 (n_14483, n20482);
  and g32003 (n20483, n_161, n_14483);
  and g32004 (n20484, n_14479, n17280);
  and g32005 (n20485, pi0038, n_14426);
  not g32006 (n_14484, n20484);
  and g32007 (n20486, n_14484, n20485);
  not g32008 (n_14485, n20483);
  not g32009 (n_14486, n20486);
  and g32010 (n20487, n_14485, n_14486);
  not g32011 (n_14487, n20487);
  and g32012 (n20488, n2571, n_14487);
  not g32013 (n_14488, n20475);
  not g32014 (n_14489, n20488);
  and g32015 (n20489, n_14488, n_14489);
  not g32016 (n_14490, n20489);
  and g32017 (n20490, n_11960, n_14490);
  and g32018 (n20491, n17117, n_14422);
  not g32019 (n_14491, n20490);
  not g32020 (n_14492, n20491);
  and g32021 (n20492, n_14491, n_14492);
  not g32022 (n_14493, n20492);
  and g32023 (n20493, n_11964, n_14493);
  and g32024 (n20494, n_11967, n_14422);
  and g32025 (n20495, pi0609, n20490);
  not g32026 (n_14494, n20494);
  not g32027 (n_14495, n20495);
  and g32028 (n20496, n_14494, n_14495);
  not g32029 (n_14496, n20496);
  and g32030 (n20497, pi1155, n_14496);
  and g32031 (n20498, n_11972, n_14422);
  and g32032 (n20499, n_11971, n20490);
  not g32033 (n_14497, n20498);
  not g32034 (n_14498, n20499);
  and g32035 (n20500, n_14497, n_14498);
  not g32036 (n_14499, n20500);
  and g32037 (n20501, n_11768, n_14499);
  not g32038 (n_14500, n20497);
  not g32039 (n_14501, n20501);
  and g32040 (n20502, n_14500, n_14501);
  not g32041 (n_14502, n20502);
  and g32042 (n20503, pi0785, n_14502);
  not g32043 (n_14503, n20493);
  not g32044 (n_14504, n20503);
  and g32045 (n20504, n_14503, n_14504);
  not g32046 (n_14505, n20504);
  and g32047 (n20505, n_11981, n_14505);
  and g32048 (n20506, n_11984, n20412);
  and g32049 (n20507, pi0618, n20504);
  not g32050 (n_14506, n20506);
  and g32051 (n20508, pi1154, n_14506);
  not g32052 (n_14507, n20507);
  and g32053 (n20509, n_14507, n20508);
  and g32054 (n20510, n_11984, n20504);
  and g32055 (n20511, pi0618, n20412);
  not g32056 (n_14508, n20511);
  and g32057 (n20512, n_11413, n_14508);
  not g32058 (n_14509, n20510);
  and g32059 (n20513, n_14509, n20512);
  not g32060 (n_14510, n20509);
  not g32061 (n_14511, n20513);
  and g32062 (n20514, n_14510, n_14511);
  not g32063 (n_14512, n20514);
  and g32064 (n20515, pi0781, n_14512);
  not g32065 (n_14513, n20505);
  not g32066 (n_14514, n20515);
  and g32067 (n20516, n_14513, n_14514);
  not g32068 (n_14515, n20516);
  and g32069 (n20517, n_12315, n_14515);
  and g32070 (n20518, n_11821, n20412);
  and g32071 (n20519, pi0619, n20516);
  not g32072 (n_14516, n20518);
  and g32073 (n20520, pi1159, n_14516);
  not g32074 (n_14517, n20519);
  and g32075 (n20521, n_14517, n20520);
  and g32076 (n20522, n_11821, n20516);
  and g32077 (n20523, pi0619, n20412);
  not g32078 (n_14518, n20523);
  and g32079 (n20524, n_11405, n_14518);
  not g32080 (n_14519, n20522);
  and g32081 (n20525, n_14519, n20524);
  not g32082 (n_14520, n20521);
  not g32083 (n_14521, n20525);
  and g32084 (n20526, n_14520, n_14521);
  not g32085 (n_14522, n20526);
  and g32086 (n20527, pi0789, n_14522);
  not g32087 (n_14523, n20517);
  not g32088 (n_14524, n20527);
  and g32089 (n20528, n_14523, n_14524);
  not g32090 (n_14525, n20528);
  and g32091 (n20529, n_12318, n_14525);
  and g32092 (n20530, n_12320, n20412);
  and g32093 (n20531, pi0626, n20528);
  not g32094 (n_14526, n20530);
  and g32095 (n20532, pi1158, n_14526);
  not g32096 (n_14527, n20531);
  and g32097 (n20533, n_14527, n20532);
  and g32098 (n20534, n_12320, n20528);
  and g32099 (n20535, pi0626, n20412);
  not g32100 (n_14528, n20535);
  and g32101 (n20536, n_11397, n_14528);
  not g32102 (n_14529, n20534);
  and g32103 (n20537, n_14529, n20536);
  not g32104 (n_14530, n20533);
  not g32105 (n_14531, n20537);
  and g32106 (n20538, n_14530, n_14531);
  not g32107 (n_14532, n20538);
  and g32108 (n20539, pi0788, n_14532);
  not g32109 (n_14533, n20529);
  not g32110 (n_14534, n20539);
  and g32111 (n20540, n_14533, n_14534);
  and g32112 (n20541, n_12368, n20540);
  and g32113 (n20542, n17779, n20412);
  not g32114 (n_14535, n20541);
  not g32115 (n_14536, n20542);
  and g32116 (n20543, n_14535, n_14536);
  not g32117 (n_14537, n20543);
  and g32118 (n20544, n_12392, n_14537);
  and g32119 (n20545, n17804, n20412);
  not g32120 (n_14538, n20544);
  not g32121 (n_14539, n20545);
  and g32122 (n20546, n_14538, n_14539);
  not g32123 (n_14540, n20546);
  and g32124 (n20547, pi0644, n_14540);
  and g32125 (n20548, n_11819, n20412);
  not g32126 (n_14541, n20548);
  and g32127 (n20549, n_12395, n_14541);
  not g32128 (n_14542, n20547);
  and g32129 (n20550, n_14542, n20549);
  not g32130 (n_14543, n20550);
  and g32131 (n20551, pi1160, n_14543);
  not g32132 (n_14544, n20474);
  and g32133 (n20552, n_14544, n20551);
  and g32134 (n20553, pi0644, n_14474);
  not g32135 (n_14545, n20463);
  and g32136 (n20554, n17802, n_14545);
  and g32137 (n20555, pi0630, n_11806);
  and g32138 (n20556, pi1157, n20555);
  and g32139 (n20557, n_12375, pi0647);
  and g32140 (n20558, n_11810, n20557);
  not g32141 (n_14546, n20556);
  not g32142 (n_14547, n20558);
  and g32143 (n20559, n_14546, n_14547);
  not g32144 (n_14548, n20559);
  and g32145 (n20560, n20543, n_14548);
  not g32146 (n_14549, n20467);
  and g32147 (n20561, n17801, n_14549);
  not g32148 (n_14550, n20554);
  not g32149 (n_14551, n20561);
  and g32150 (n20562, n_14550, n_14551);
  not g32151 (n_14552, n20560);
  and g32152 (n20563, n_14552, n20562);
  not g32153 (n_14553, n20563);
  and g32154 (n20564, pi0787, n_14553);
  and g32155 (n20565, n_12354, n20453);
  and g32156 (n20566, n_11789, pi0629);
  and g32157 (n20567, pi1156, n20566);
  and g32158 (n20568, pi0628, n_12354);
  and g32159 (n20569, n_11794, n20568);
  not g32160 (n_14554, n20567);
  not g32161 (n_14555, n20569);
  and g32162 (n20570, n_14554, n_14555);
  not g32163 (n_14556, n20540);
  not g32164 (n_14557, n20570);
  and g32165 (n20571, n_14556, n_14557);
  and g32166 (n20572, pi0629, n20457);
  not g32167 (n_14558, n20565);
  not g32168 (n_14559, n20572);
  and g32169 (n20573, n_14558, n_14559);
  not g32170 (n_14560, n20571);
  and g32171 (n20574, n_14560, n20573);
  not g32172 (n_14561, n20574);
  and g32173 (n20575, pi0792, n_14561);
  and g32174 (n20576, pi0609, n20437);
  and g32175 (n20577, pi0145, n_12240);
  and g32176 (n20578, n_6246, n_12230);
  not g32177 (n_14562, n20577);
  and g32178 (n20579, pi0767, n_14562);
  not g32179 (n_14563, n20578);
  and g32180 (n20580, n_14563, n20579);
  and g32181 (n20581, n_6246, n17629);
  and g32182 (n20582, pi0145, n17631);
  not g32183 (n_14564, n20582);
  and g32184 (n20583, n_14479, n_14564);
  not g32185 (n_14565, n20581);
  and g32186 (n20584, n_14565, n20583);
  not g32187 (n_14566, n20580);
  not g32188 (n_14567, n20584);
  and g32189 (n20585, n_14566, n_14567);
  not g32190 (n_14568, n20585);
  and g32191 (n20586, n_162, n_14568);
  and g32192 (n20587, pi0145, n17605);
  and g32193 (n20588, n_6246, n_12180);
  not g32194 (n_14569, n20588);
  and g32195 (n20589, n_14479, n_14569);
  not g32196 (n_14570, n20587);
  and g32197 (n20590, n_14570, n20589);
  and g32198 (n20591, n_6246, n17404);
  and g32199 (n20592, pi0145, n17485);
  not g32200 (n_14571, n20592);
  and g32201 (n20593, pi0767, n_14571);
  not g32202 (n_14572, n20591);
  and g32203 (n20594, n_14572, n20593);
  not g32204 (n_14573, n20590);
  and g32205 (n20595, pi0039, n_14573);
  not g32206 (n_14574, n20594);
  and g32207 (n20596, n_14574, n20595);
  not g32208 (n_14575, n20586);
  and g32209 (n20597, n_161, n_14575);
  not g32210 (n_14576, n20596);
  and g32211 (n20598, n_14576, n20597);
  and g32212 (n20599, n_14479, n_12250);
  not g32213 (n_14577, n20599);
  and g32214 (n20600, n19471, n_14577);
  not g32215 (n_14578, n20600);
  and g32216 (n20601, n_6246, n_14578);
  and g32217 (n20602, n_14479, n17244);
  not g32218 (n_14579, n20602);
  and g32219 (n20603, n_12120, n_14579);
  not g32220 (n_14580, n20603);
  and g32221 (n20604, pi0145, n_14580);
  and g32222 (n20605, n6284, n20604);
  not g32223 (n_14581, n20605);
  and g32224 (n20606, pi0038, n_14581);
  not g32225 (n_14582, n20601);
  and g32226 (n20607, n_14582, n20606);
  not g32227 (n_14583, n20607);
  and g32228 (n20608, n_14424, n_14583);
  not g32229 (n_14584, n20598);
  and g32230 (n20609, n_14584, n20608);
  and g32231 (n20610, pi0698, n20487);
  not g32232 (n_14585, n20609);
  and g32233 (n20611, n2571, n_14585);
  not g32234 (n_14586, n20610);
  and g32235 (n20612, n_14586, n20611);
  not g32236 (n_14587, n20612);
  and g32237 (n20613, n_14488, n_14587);
  and g32238 (n20614, n_11753, n20613);
  and g32239 (n20615, pi0625, n20489);
  not g32240 (n_14588, n20615);
  and g32241 (n20616, n_11757, n_14588);
  not g32242 (n_14589, n20614);
  and g32243 (n20617, n_14589, n20616);
  and g32244 (n20618, n_11823, n_14440);
  not g32245 (n_14590, n20617);
  and g32246 (n20619, n_14590, n20618);
  and g32247 (n20620, n_11753, n20489);
  and g32248 (n20621, pi0625, n20613);
  not g32249 (n_14591, n20620);
  and g32250 (n20622, pi1153, n_14591);
  not g32251 (n_14592, n20621);
  and g32252 (n20623, n_14592, n20622);
  and g32253 (n20624, pi0608, n_14441);
  not g32254 (n_14593, n20623);
  and g32255 (n20625, n_14593, n20624);
  not g32256 (n_14594, n20619);
  not g32257 (n_14595, n20625);
  and g32258 (n20626, n_14594, n_14595);
  not g32259 (n_14596, n20626);
  and g32260 (n20627, pi0778, n_14596);
  and g32261 (n20628, n_11749, n20613);
  not g32262 (n_14597, n20627);
  not g32263 (n_14598, n20628);
  and g32264 (n20629, n_14597, n_14598);
  not g32265 (n_14599, n20629);
  and g32266 (n20630, n_11971, n_14599);
  not g32267 (n_14600, n20576);
  and g32268 (n20631, n_11768, n_14600);
  not g32269 (n_14601, n20630);
  and g32270 (n20632, n_14601, n20631);
  and g32271 (n20633, n_11767, n_14500);
  not g32272 (n_14602, n20632);
  and g32273 (n20634, n_14602, n20633);
  and g32274 (n20635, n_11971, n20437);
  and g32275 (n20636, pi0609, n_14599);
  not g32276 (n_14603, n20635);
  and g32277 (n20637, pi1155, n_14603);
  not g32278 (n_14604, n20636);
  and g32279 (n20638, n_14604, n20637);
  and g32280 (n20639, pi0660, n_14501);
  not g32281 (n_14605, n20638);
  and g32282 (n20640, n_14605, n20639);
  not g32283 (n_14606, n20634);
  not g32284 (n_14607, n20640);
  and g32285 (n20641, n_14606, n_14607);
  not g32286 (n_14608, n20641);
  and g32287 (n20642, pi0785, n_14608);
  and g32288 (n20643, n_11964, n_14599);
  not g32289 (n_14609, n20642);
  not g32290 (n_14610, n20643);
  and g32291 (n20644, n_14609, n_14610);
  not g32292 (n_14611, n20644);
  and g32293 (n20645, n_11984, n_14611);
  and g32294 (n20646, pi0618, n20440);
  not g32295 (n_14612, n20646);
  and g32296 (n20647, n_11413, n_14612);
  not g32297 (n_14613, n20645);
  and g32298 (n20648, n_14613, n20647);
  and g32299 (n20649, n_11412, n_14510);
  not g32300 (n_14614, n20648);
  and g32301 (n20650, n_14614, n20649);
  and g32302 (n20651, n_11984, n20440);
  and g32303 (n20652, pi0618, n_14611);
  not g32304 (n_14615, n20651);
  and g32305 (n20653, pi1154, n_14615);
  not g32306 (n_14616, n20652);
  and g32307 (n20654, n_14616, n20653);
  and g32308 (n20655, pi0627, n_14511);
  not g32309 (n_14617, n20654);
  and g32310 (n20656, n_14617, n20655);
  not g32311 (n_14618, n20650);
  not g32312 (n_14619, n20656);
  and g32313 (n20657, n_14618, n_14619);
  not g32314 (n_14620, n20657);
  and g32315 (n20658, pi0781, n_14620);
  and g32316 (n20659, n_11981, n_14611);
  not g32317 (n_14621, n20658);
  not g32318 (n_14622, n20659);
  and g32319 (n20660, n_14621, n_14622);
  and g32320 (n20661, n_12315, n20660);
  not g32321 (n_14623, n20443);
  and g32322 (n20662, pi0619, n_14623);
  not g32323 (n_14624, n20660);
  and g32324 (n20663, n_11821, n_14624);
  not g32325 (n_14625, n20662);
  and g32326 (n20664, n_11405, n_14625);
  not g32327 (n_14626, n20663);
  and g32328 (n20665, n_14626, n20664);
  and g32329 (n20666, n_11403, n_14520);
  not g32330 (n_14627, n20665);
  and g32331 (n20667, n_14627, n20666);
  and g32332 (n20668, pi0619, n_14624);
  and g32333 (n20669, n_11821, n_14623);
  not g32334 (n_14628, n20669);
  and g32335 (n20670, pi1159, n_14628);
  not g32336 (n_14629, n20668);
  and g32337 (n20671, n_14629, n20670);
  and g32338 (n20672, pi0648, n_14521);
  not g32339 (n_14630, n20671);
  and g32340 (n20673, n_14630, n20672);
  not g32341 (n_14631, n20667);
  and g32342 (n20674, pi0789, n_14631);
  not g32343 (n_14632, n20673);
  and g32344 (n20675, n_14632, n20674);
  not g32345 (n_14633, n20661);
  and g32346 (n20676, n17970, n_14633);
  not g32347 (n_14634, n20675);
  and g32348 (n20677, n_14634, n20676);
  and g32349 (n20678, n17871, n20445);
  and g32350 (n20679, n_11401, n20538);
  not g32351 (n_14635, n20678);
  not g32352 (n_14636, n20679);
  and g32353 (n20680, n_14635, n_14636);
  not g32354 (n_14637, n20680);
  and g32355 (n20681, pi0788, n_14637);
  not g32356 (n_14638, n20364);
  not g32357 (n_14639, n20681);
  and g32358 (n20682, n_14638, n_14639);
  not g32359 (n_14640, n20677);
  and g32360 (n20683, n_14640, n20682);
  not g32361 (n_14641, n20575);
  not g32362 (n_14642, n20683);
  and g32363 (n20684, n_14641, n_14642);
  not g32364 (n_14643, n20684);
  and g32365 (n20685, n_14387, n_14643);
  not g32366 (n_14644, n20564);
  not g32367 (n_14645, n20685);
  and g32368 (n20686, n_14644, n_14645);
  and g32369 (n20687, n_11819, n20686);
  not g32370 (n_14646, n20553);
  and g32371 (n20688, n_12395, n_14646);
  not g32372 (n_14647, n20687);
  and g32373 (n20689, n_14647, n20688);
  and g32374 (n20690, pi0644, n20412);
  and g32375 (n20691, n_11819, n_14540);
  not g32376 (n_14648, n20690);
  and g32377 (n20692, pi0715, n_14648);
  not g32378 (n_14649, n20691);
  and g32379 (n20693, n_14649, n20692);
  not g32380 (n_14650, n20693);
  and g32381 (n20694, n_12405, n_14650);
  not g32382 (n_14651, n20689);
  and g32383 (n20695, n_14651, n20694);
  not g32384 (n_14652, n20552);
  not g32385 (n_14653, n20695);
  and g32386 (n20696, n_14652, n_14653);
  not g32387 (n_14654, n20696);
  and g32388 (n20697, pi0790, n_14654);
  and g32389 (n20698, pi0644, n20551);
  not g32390 (n_14655, n20698);
  and g32391 (n20699, pi0790, n_14655);
  not g32392 (n_14656, n20699);
  and g32393 (n20700, n20686, n_14656);
  not g32394 (n_14657, n20697);
  not g32395 (n_14658, n20700);
  and g32396 (n20701, n_14657, n_14658);
  not g32397 (n_14659, n20701);
  and g32398 (n20702, n_4226, n_14659);
  not g32399 (n_14660, n20411);
  and g32400 (n20703, n_12415, n_14660);
  not g32401 (n_14661, n20702);
  and g32402 (n20704, n_14661, n20703);
  and g32403 (n20705, n_6246, n_12418);
  and g32404 (n20706, n_14424, n16645);
  not g32405 (n_14662, n20705);
  not g32406 (n_14663, n20706);
  and g32407 (n20707, n_14662, n_14663);
  and g32408 (n20708, n_11749, n20707);
  and g32409 (n20709, n_11753, n20706);
  not g32410 (n_14664, n20707);
  not g32411 (n_14665, n20709);
  and g32412 (n20710, n_14664, n_14665);
  not g32413 (n_14666, n20710);
  and g32414 (n20711, pi1153, n_14666);
  and g32415 (n20712, n_11757, n_14662);
  and g32416 (n20713, n_14665, n20712);
  not g32417 (n_14667, n20711);
  not g32418 (n_14668, n20713);
  and g32419 (n20714, n_14667, n_14668);
  not g32420 (n_14669, n20714);
  and g32421 (n20715, pi0778, n_14669);
  not g32422 (n_14670, n20708);
  not g32423 (n_14671, n20715);
  and g32424 (n20716, n_14670, n_14671);
  and g32425 (n20717, n_12429, n20716);
  and g32426 (n20718, n_12430, n20717);
  and g32427 (n20719, n_12431, n20718);
  and g32428 (n20720, n_12432, n20719);
  and g32429 (n20721, n_12436, n20720);
  and g32430 (n20722, n_11806, n20721);
  and g32431 (n20723, pi0647, n20705);
  not g32432 (n_14672, n20723);
  and g32433 (n20724, n_11810, n_14672);
  not g32434 (n_14673, n20722);
  and g32435 (n20725, n_14673, n20724);
  and g32436 (n20726, pi0630, n20725);
  and g32437 (n20727, n_14579, n_14662);
  not g32438 (n_14674, n20727);
  and g32439 (n20728, n_12448, n_14674);
  not g32440 (n_14675, n20728);
  and g32441 (n20729, n_11964, n_14675);
  and g32442 (n20730, n_12451, n_14674);
  not g32443 (n_14676, n20730);
  and g32444 (n20731, pi1155, n_14676);
  and g32445 (n20732, n_12453, n20728);
  not g32446 (n_14677, n20732);
  and g32447 (n20733, n_11768, n_14677);
  not g32448 (n_14678, n20731);
  not g32449 (n_14679, n20733);
  and g32450 (n20734, n_14678, n_14679);
  not g32451 (n_14680, n20734);
  and g32452 (n20735, pi0785, n_14680);
  not g32453 (n_14681, n20729);
  not g32454 (n_14682, n20735);
  and g32455 (n20736, n_14681, n_14682);
  not g32456 (n_14683, n20736);
  and g32457 (n20737, n_11981, n_14683);
  and g32458 (n20738, n_12461, n20736);
  not g32459 (n_14684, n20738);
  and g32460 (n20739, pi1154, n_14684);
  and g32461 (n20740, n_12463, n20736);
  not g32462 (n_14685, n20740);
  and g32463 (n20741, n_11413, n_14685);
  not g32464 (n_14686, n20739);
  not g32465 (n_14687, n20741);
  and g32466 (n20742, n_14686, n_14687);
  not g32467 (n_14688, n20742);
  and g32468 (n20743, pi0781, n_14688);
  not g32469 (n_14689, n20737);
  not g32470 (n_14690, n20743);
  and g32471 (n20744, n_14689, n_14690);
  not g32472 (n_14691, n20744);
  and g32473 (n20745, n_12315, n_14691);
  and g32474 (n20746, n_11821, n20705);
  and g32475 (n20747, pi0619, n20744);
  not g32476 (n_14692, n20746);
  and g32477 (n20748, pi1159, n_14692);
  not g32478 (n_14693, n20747);
  and g32479 (n20749, n_14693, n20748);
  and g32480 (n20750, n_11821, n20744);
  and g32481 (n20751, pi0619, n20705);
  not g32482 (n_14694, n20751);
  and g32483 (n20752, n_11405, n_14694);
  not g32484 (n_14695, n20750);
  and g32485 (n20753, n_14695, n20752);
  not g32486 (n_14696, n20749);
  not g32487 (n_14697, n20753);
  and g32488 (n20754, n_14696, n_14697);
  not g32489 (n_14698, n20754);
  and g32490 (n20755, pi0789, n_14698);
  not g32491 (n_14699, n20745);
  not g32492 (n_14700, n20755);
  and g32493 (n20756, n_14699, n_14700);
  not g32494 (n_14701, n20756);
  and g32495 (n20757, n_12318, n_14701);
  and g32496 (n20758, n_12320, n20705);
  and g32497 (n20759, pi0626, n20756);
  not g32498 (n_14702, n20758);
  and g32499 (n20760, pi1158, n_14702);
  not g32500 (n_14703, n20759);
  and g32501 (n20761, n_14703, n20760);
  and g32502 (n20762, n_12320, n20756);
  and g32503 (n20763, pi0626, n20705);
  not g32504 (n_14704, n20763);
  and g32505 (n20764, n_11397, n_14704);
  not g32506 (n_14705, n20762);
  and g32507 (n20765, n_14705, n20764);
  not g32508 (n_14706, n20761);
  not g32509 (n_14707, n20765);
  and g32510 (n20766, n_14706, n_14707);
  not g32511 (n_14708, n20766);
  and g32512 (n20767, pi0788, n_14708);
  not g32513 (n_14709, n20757);
  not g32514 (n_14710, n20767);
  and g32515 (n20768, n_14709, n_14710);
  and g32516 (n20769, n_12368, n20768);
  and g32517 (n20770, n17779, n20705);
  not g32518 (n_14711, n20769);
  not g32519 (n_14712, n20770);
  and g32520 (n20771, n_14711, n_14712);
  and g32521 (n20772, n_14548, n20771);
  not g32522 (n_14713, n20721);
  and g32523 (n20773, pi0647, n_14713);
  and g32524 (n20774, n_11806, n_14662);
  not g32525 (n_14714, n20773);
  not g32526 (n_14715, n20774);
  and g32527 (n20775, n_14714, n_14715);
  not g32528 (n_14716, n20775);
  and g32529 (n20776, n17801, n_14716);
  not g32530 (n_14717, n20726);
  not g32531 (n_14718, n20776);
  and g32532 (n20777, n_14717, n_14718);
  not g32533 (n_14719, n20772);
  and g32534 (n20778, n_14719, n20777);
  not g32535 (n_14720, n20778);
  and g32536 (n20779, pi0787, n_14720);
  and g32537 (n20780, n17871, n20719);
  and g32538 (n20781, n_11401, n20766);
  not g32539 (n_14721, n20780);
  not g32540 (n_14722, n20781);
  and g32541 (n20782, n_14721, n_14722);
  not g32542 (n_14723, n20782);
  and g32543 (n20783, pi0788, n_14723);
  and g32544 (n20784, pi0618, n20717);
  and g32545 (n20785, pi0609, n20716);
  and g32546 (n20786, n_11866, n_14664);
  and g32547 (n20787, pi0625, n20786);
  not g32548 (n_14724, n20786);
  and g32549 (n20788, n20727, n_14724);
  not g32550 (n_14725, n20787);
  not g32551 (n_14726, n20788);
  and g32552 (n20789, n_14725, n_14726);
  not g32553 (n_14727, n20789);
  and g32554 (n20790, n20712, n_14727);
  and g32555 (n20791, n_11823, n_14667);
  not g32556 (n_14728, n20790);
  and g32557 (n20792, n_14728, n20791);
  and g32558 (n20793, pi1153, n20727);
  and g32559 (n20794, n_14725, n20793);
  and g32560 (n20795, pi0608, n_14668);
  not g32561 (n_14729, n20794);
  and g32562 (n20796, n_14729, n20795);
  not g32563 (n_14730, n20792);
  not g32564 (n_14731, n20796);
  and g32565 (n20797, n_14730, n_14731);
  not g32566 (n_14732, n20797);
  and g32567 (n20798, pi0778, n_14732);
  and g32568 (n20799, n_11749, n_14726);
  not g32569 (n_14733, n20798);
  not g32570 (n_14734, n20799);
  and g32571 (n20800, n_14733, n_14734);
  not g32572 (n_14735, n20800);
  and g32573 (n20801, n_11971, n_14735);
  not g32574 (n_14736, n20785);
  and g32575 (n20802, n_11768, n_14736);
  not g32576 (n_14737, n20801);
  and g32577 (n20803, n_14737, n20802);
  and g32578 (n20804, n_11767, n_14678);
  not g32579 (n_14738, n20803);
  and g32580 (n20805, n_14738, n20804);
  and g32581 (n20806, n_11971, n20716);
  and g32582 (n20807, pi0609, n_14735);
  not g32583 (n_14739, n20806);
  and g32584 (n20808, pi1155, n_14739);
  not g32585 (n_14740, n20807);
  and g32586 (n20809, n_14740, n20808);
  and g32587 (n20810, pi0660, n_14679);
  not g32588 (n_14741, n20809);
  and g32589 (n20811, n_14741, n20810);
  not g32590 (n_14742, n20805);
  not g32591 (n_14743, n20811);
  and g32592 (n20812, n_14742, n_14743);
  not g32593 (n_14744, n20812);
  and g32594 (n20813, pi0785, n_14744);
  and g32595 (n20814, n_11964, n_14735);
  not g32596 (n_14745, n20813);
  not g32597 (n_14746, n20814);
  and g32598 (n20815, n_14745, n_14746);
  not g32599 (n_14747, n20815);
  and g32600 (n20816, n_11984, n_14747);
  not g32601 (n_14748, n20784);
  and g32602 (n20817, n_11413, n_14748);
  not g32603 (n_14749, n20816);
  and g32604 (n20818, n_14749, n20817);
  and g32605 (n20819, n_11412, n_14686);
  not g32606 (n_14750, n20818);
  and g32607 (n20820, n_14750, n20819);
  and g32608 (n20821, n_11984, n20717);
  and g32609 (n20822, pi0618, n_14747);
  not g32610 (n_14751, n20821);
  and g32611 (n20823, pi1154, n_14751);
  not g32612 (n_14752, n20822);
  and g32613 (n20824, n_14752, n20823);
  and g32614 (n20825, pi0627, n_14687);
  not g32615 (n_14753, n20824);
  and g32616 (n20826, n_14753, n20825);
  not g32617 (n_14754, n20820);
  not g32618 (n_14755, n20826);
  and g32619 (n20827, n_14754, n_14755);
  not g32620 (n_14756, n20827);
  and g32621 (n20828, pi0781, n_14756);
  and g32622 (n20829, n_11981, n_14747);
  not g32623 (n_14757, n20828);
  not g32624 (n_14758, n20829);
  and g32625 (n20830, n_14757, n_14758);
  and g32626 (n20831, n_12315, n20830);
  not g32627 (n_14759, n20830);
  and g32628 (n20832, n_11821, n_14759);
  and g32629 (n20833, pi0619, n20718);
  not g32630 (n_14760, n20833);
  and g32631 (n20834, n_11405, n_14760);
  not g32632 (n_14761, n20832);
  and g32633 (n20835, n_14761, n20834);
  and g32634 (n20836, n_11403, n_14696);
  not g32635 (n_14762, n20835);
  and g32636 (n20837, n_14762, n20836);
  and g32637 (n20838, n_11821, n20718);
  and g32638 (n20839, pi0619, n_14759);
  not g32639 (n_14763, n20838);
  and g32640 (n20840, pi1159, n_14763);
  not g32641 (n_14764, n20839);
  and g32642 (n20841, n_14764, n20840);
  and g32643 (n20842, pi0648, n_14697);
  not g32644 (n_14765, n20841);
  and g32645 (n20843, n_14765, n20842);
  not g32646 (n_14766, n20837);
  and g32647 (n20844, pi0789, n_14766);
  not g32648 (n_14767, n20843);
  and g32649 (n20845, n_14767, n20844);
  not g32650 (n_14768, n20831);
  and g32651 (n20846, n17970, n_14768);
  not g32652 (n_14769, n20845);
  and g32653 (n20847, n_14769, n20846);
  not g32654 (n_14770, n20783);
  not g32655 (n_14771, n20847);
  and g32656 (n20848, n_14770, n_14771);
  not g32657 (n_14772, n20848);
  and g32658 (n20849, n_14638, n_14772);
  and g32659 (n20850, n17854, n20768);
  and g32660 (n20851, pi1156, n_12439);
  and g32661 (n20852, n20720, n20851);
  not g32662 (n_14773, n20850);
  not g32663 (n_14774, n20852);
  and g32664 (n20853, n_14773, n_14774);
  not g32665 (n_14775, n20853);
  and g32666 (n20854, n_12354, n_14775);
  and g32667 (n20855, n_11794, n_12547);
  and g32668 (n20856, n20720, n20855);
  and g32669 (n20857, n17853, n20768);
  not g32670 (n_14776, n20856);
  not g32671 (n_14777, n20857);
  and g32672 (n20858, n_14776, n_14777);
  not g32673 (n_14778, n20858);
  and g32674 (n20859, pi0629, n_14778);
  not g32675 (n_14779, n20854);
  not g32676 (n_14780, n20859);
  and g32677 (n20860, n_14779, n_14780);
  not g32678 (n_14781, n20860);
  and g32679 (n20861, pi0792, n_14781);
  not g32680 (n_14782, n20861);
  and g32681 (n20862, n_14387, n_14782);
  not g32682 (n_14783, n20849);
  and g32683 (n20863, n_14783, n20862);
  not g32684 (n_14784, n20779);
  not g32685 (n_14785, n20863);
  and g32686 (n20864, n_14784, n_14785);
  and g32687 (n20865, n_12411, n20864);
  and g32688 (n20866, n_11803, n_14713);
  and g32689 (n20867, pi1157, n_14716);
  not g32690 (n_14786, n20725);
  not g32691 (n_14787, n20867);
  and g32692 (n20868, n_14786, n_14787);
  not g32693 (n_14788, n20868);
  and g32694 (n20869, pi0787, n_14788);
  not g32695 (n_14789, n20866);
  not g32696 (n_14790, n20869);
  and g32697 (n20870, n_14789, n_14790);
  and g32698 (n20871, n_11819, n20870);
  and g32699 (n20872, pi0644, n20864);
  not g32700 (n_14791, n20871);
  and g32701 (n20873, pi0715, n_14791);
  not g32702 (n_14792, n20872);
  and g32703 (n20874, n_14792, n20873);
  not g32704 (n_14793, n20771);
  and g32705 (n20875, n_12392, n_14793);
  and g32706 (n20876, n17804, n20705);
  not g32707 (n_14794, n20875);
  not g32708 (n_14795, n20876);
  and g32709 (n20877, n_14794, n_14795);
  not g32710 (n_14796, n20877);
  and g32711 (n20878, pi0644, n_14796);
  and g32712 (n20879, n_11819, n20705);
  not g32713 (n_14797, n20879);
  and g32714 (n20880, n_12395, n_14797);
  not g32715 (n_14798, n20878);
  and g32716 (n20881, n_14798, n20880);
  not g32717 (n_14799, n20881);
  and g32718 (n20882, pi1160, n_14799);
  not g32719 (n_14800, n20874);
  and g32720 (n20883, n_14800, n20882);
  and g32721 (n20884, n_11819, n_14796);
  and g32722 (n20885, pi0644, n20705);
  not g32723 (n_14801, n20885);
  and g32724 (n20886, pi0715, n_14801);
  not g32725 (n_14802, n20884);
  and g32726 (n20887, n_14802, n20886);
  and g32727 (n20888, pi0644, n20870);
  and g32728 (n20889, n_11819, n20864);
  not g32729 (n_14803, n20888);
  and g32730 (n20890, n_12395, n_14803);
  not g32731 (n_14804, n20889);
  and g32732 (n20891, n_14804, n20890);
  not g32733 (n_14805, n20887);
  and g32734 (n20892, n_12405, n_14805);
  not g32735 (n_14806, n20891);
  and g32736 (n20893, n_14806, n20892);
  not g32737 (n_14807, n20883);
  not g32738 (n_14808, n20893);
  and g32739 (n20894, n_14807, n_14808);
  not g32740 (n_14809, n20894);
  and g32741 (n20895, pi0790, n_14809);
  not g32742 (n_14810, n20865);
  and g32743 (n20896, pi0832, n_14810);
  not g32744 (n_14811, n20895);
  and g32745 (n20897, n_14811, n20896);
  not g32746 (n_14812, n20704);
  not g32747 (n_14813, n20897);
  and g32748 (po0302, n_14812, n_14813);
  not g32749 (n_14814, n10197);
  and g32750 (n20899, n_268, n_14814);
  and g32751 (n20900, n_268, n_11418);
  and g32752 (n20901, pi0743, pi0947);
  and g32753 (n20902, pi0907, n_3149);
  and g32754 (n20903, pi0735, n20902);
  not g32755 (n_14815, n20901);
  not g32756 (n_14816, n20903);
  and g32757 (n20904, n_14815, n_14816);
  and g32758 (n20905, n2926, n20904);
  and g32759 (n20906, n6284, n20905);
  not g32760 (n_14817, n20906);
  and g32761 (n20907, pi0038, n_14817);
  not g32762 (n_14818, n20900);
  and g32763 (n20908, n_14818, n20907);
  and g32764 (n20909, n_268, n_11670);
  and g32765 (n20910, n16941, n20904);
  not g32766 (n_14819, n20909);
  and g32767 (n20911, pi0299, n_14819);
  not g32768 (n_14820, n20910);
  and g32769 (n20912, n_14820, n20911);
  and g32770 (n20913, n_268, n_11671);
  and g32771 (n20914, n16930, n20904);
  not g32772 (n_14821, n20913);
  and g32773 (n20915, n_234, n_14821);
  not g32774 (n_14822, n20914);
  and g32775 (n20916, n_14822, n20915);
  not g32776 (n_14823, n20912);
  and g32777 (n20917, n_162, n_14823);
  not g32778 (n_14824, n20916);
  and g32779 (n20918, n_14824, n20917);
  not g32780 (n_14825, n20904);
  and g32781 (n20919, n16653, n_14825);
  and g32782 (n20920, pi0146, n_11445);
  not g32783 (n_14826, n20919);
  not g32784 (n_14827, n20920);
  and g32785 (n20921, n_14826, n_14827);
  not g32786 (n_14828, n20921);
  and g32787 (n20922, n3448, n_14828);
  and g32788 (n20923, n_3148, n6241);
  and g32789 (n20924, pi0146, n_11712);
  not g32790 (n_14829, n20923);
  and g32791 (n20925, n_14829, n20924);
  and g32792 (n20926, pi0735, pi0907);
  and g32793 (n20927, n17018, n20926);
  and g32794 (n20928, pi0146, n_11706);
  and g32795 (n20929, n20923, n20928);
  not g32796 (n_14830, n20927);
  and g32797 (n20930, n_3149, n_14830);
  not g32798 (n_14831, n20929);
  and g32799 (n20931, n_14831, n20930);
  and g32800 (n20932, pi0743, n17018);
  not g32801 (n_14832, n20924);
  and g32802 (n20933, pi0947, n_14832);
  not g32803 (n_14833, n20932);
  and g32804 (n20934, n_14833, n20933);
  not g32805 (n_14834, n20931);
  not g32806 (n_14835, n20934);
  and g32807 (n20935, n_14834, n_14835);
  not g32808 (n_14836, n20925);
  not g32809 (n_14837, n20935);
  and g32810 (n20936, n_14836, n_14837);
  not g32811 (n_14838, n20936);
  and g32812 (n20937, n_9350, n_14838);
  not g32813 (n_14839, n20922);
  and g32814 (n20938, n_36, n_14839);
  not g32815 (n_14840, n20937);
  and g32816 (n20939, n_14840, n20938);
  and g32817 (n20940, n16970, n_14825);
  and g32818 (n20941, pi0146, n17042);
  not g32819 (n_14841, n20940);
  and g32820 (n20942, pi0215, n_14841);
  not g32821 (n_14842, n20941);
  and g32822 (n20943, n_14842, n20942);
  not g32823 (n_14843, n20939);
  not g32824 (n_14844, n20943);
  and g32825 (n20944, n_14843, n_14844);
  not g32826 (n_14845, n20944);
  and g32827 (n20945, pi0299, n_14845);
  and g32828 (n20946, pi0146, n_11684);
  not g32829 (n_14846, n20946);
  and g32830 (n20947, n_14841, n_14846);
  not g32831 (n_14847, n20947);
  and g32832 (n20948, n_3119, n_14847);
  and g32833 (n20949, n_268, n_11694);
  and g32834 (n20950, n16990, n20904);
  not g32835 (n_14848, n20949);
  and g32836 (n20951, n6205, n_14848);
  not g32837 (n_14849, n20950);
  and g32838 (n20952, n_14849, n20951);
  not g32839 (n_14850, n20948);
  not g32840 (n_14851, n20952);
  and g32841 (n20953, n_14850, n_14851);
  not g32842 (n_14852, n20953);
  and g32843 (n20954, pi0223, n_14852);
  and g32844 (n20955, n2603, n20921);
  and g32845 (n20956, n17018, n_14825);
  and g32846 (n20957, n_3119, n_14832);
  not g32847 (n_14853, n20956);
  and g32848 (n20958, n_14853, n20957);
  and g32849 (n20959, n17011, n_14825);
  not g32850 (n_14854, n20928);
  and g32851 (n20960, n6205, n_14854);
  not g32852 (n_14855, n20959);
  and g32853 (n20961, n_14855, n20960);
  not g32854 (n_14856, n20958);
  not g32855 (n_14857, n20961);
  and g32856 (n20962, n_14856, n_14857);
  not g32857 (n_14858, n20962);
  and g32858 (n20963, n_9349, n_14858);
  not g32859 (n_14859, n20955);
  and g32860 (n20964, n_223, n_14859);
  not g32861 (n_14860, n20963);
  and g32862 (n20965, n_14860, n20964);
  not g32863 (n_14861, n20954);
  and g32864 (n20966, n_234, n_14861);
  not g32865 (n_14862, n20965);
  and g32866 (n20967, n_14862, n20966);
  not g32867 (n_14863, n20945);
  not g32868 (n_14864, n20967);
  and g32869 (n20968, n_14863, n_14864);
  not g32870 (n_14865, n20968);
  and g32871 (n20969, pi0039, n_14865);
  not g32872 (n_14866, n20918);
  and g32873 (n20970, n_161, n_14866);
  not g32874 (n_14867, n20969);
  and g32875 (n20971, n_14867, n20970);
  not g32876 (n_14868, n20908);
  and g32877 (n20972, n10197, n_14868);
  not g32878 (n_14869, n20971);
  and g32879 (n20973, n_14869, n20972);
  not g32880 (n_14870, n20899);
  and g32881 (n20974, n_12415, n_14870);
  not g32882 (n_14871, n20973);
  and g32883 (n20975, n_14871, n20974);
  and g32884 (n20976, n_268, n_12418);
  not g32885 (n_14872, n20976);
  and g32886 (n20977, pi0832, n_14872);
  not g32887 (n_14873, n20905);
  and g32888 (n20978, n_14873, n20977);
  or g32889 (po0303, n20975, n20978);
  and g32890 (n20980, n_7628, n_12418);
  not g32891 (n_14875, pi0770);
  and g32892 (n20981, n_14875, pi0947);
  and g32893 (n20982, pi0726, n20902);
  not g32894 (n_14877, n20981);
  not g32895 (n_14878, n20982);
  and g32896 (n20983, n_14877, n_14878);
  not g32897 (n_14879, n20983);
  and g32898 (n20984, n2926, n_14879);
  not g32899 (n_14880, n20980);
  and g32900 (n20985, pi0832, n_14880);
  not g32901 (n_14881, n20984);
  and g32902 (n20986, n_14881, n20985);
  and g32903 (n20987, n_7628, n_14814);
  and g32904 (n20988, n_3149, n16958);
  not g32905 (n_14882, n20988);
  and g32906 (n20989, n_162, n_14882);
  and g32907 (n20990, n_234, n17024);
  and g32908 (n20991, pi0947, n20990);
  and g32909 (n20992, n_3149, n17026);
  and g32910 (n20993, n17018, n20902);
  not g32911 (n_14883, n17030);
  not g32912 (n_14884, n20993);
  and g32913 (n20994, n_14883, n_14884);
  not g32914 (n_14885, n20994);
  and g32915 (n20995, n_9350, n_14885);
  not g32916 (n_14886, n20995);
  and g32917 (n20996, n_36, n_14886);
  not g32918 (n_14887, n20992);
  and g32919 (n20997, n_14887, n20996);
  and g32920 (n20998, pi0215, n_11730);
  and g32921 (n20999, n16970, n20902);
  not g32922 (n_14888, n20999);
  and g32923 (n21000, n20998, n_14888);
  not g32924 (n_14889, n20997);
  not g32925 (n_14890, n21000);
  and g32926 (n21001, n_14889, n_14890);
  not g32927 (n_14891, n21001);
  and g32928 (n21002, pi0299, n_14891);
  not g32929 (n_14892, n21002);
  and g32930 (n21003, n_11734, n_14892);
  not g32931 (n_14893, n20991);
  and g32932 (n21004, n_14893, n21003);
  not g32933 (n_14894, n21004);
  and g32934 (n21005, pi0039, n_14894);
  not g32935 (n_14895, n20989);
  not g32936 (n_14896, n21005);
  and g32937 (n21006, n_14895, n_14896);
  and g32938 (n21007, n_161, n21006);
  and g32939 (n21008, pi0038, n_3149);
  and g32940 (n21009, n17050, n21008);
  not g32941 (n_14897, n21007);
  not g32942 (n_14898, n21009);
  and g32943 (n21010, n_14897, n_14898);
  and g32944 (n21011, n_14875, n21010);
  and g32945 (n21012, pi0770, n_11743);
  not g32946 (n_14899, n21011);
  not g32947 (n_14900, n21012);
  and g32948 (n21013, n_14899, n_14900);
  not g32949 (n_14901, n21013);
  and g32950 (n21014, n_7628, n_14901);
  and g32951 (n21015, n_11742, n_14898);
  and g32952 (n21016, pi0947, n16958);
  not g32953 (n_14902, n21016);
  and g32954 (n21017, n_162, n_14902);
  and g32955 (n21018, pi0947, n17024);
  not g32956 (n_14903, n21018);
  and g32957 (n21019, n_234, n_14903);
  and g32958 (n21020, pi0215, pi0947);
  and g32959 (n21021, n16970, n21020);
  not g32960 (n_14904, n21021);
  and g32961 (n21022, pi0299, n_14904);
  and g32962 (n21023, pi0947, n17018);
  not g32963 (n_14905, n21023);
  and g32964 (n21024, n_9350, n_14905);
  and g32965 (n21025, pi0947, n16653);
  not g32966 (n_14906, n21025);
  and g32967 (n21026, n3448, n_14906);
  not g32968 (n_14907, n21026);
  and g32969 (n21027, n_36, n_14907);
  not g32970 (n_14908, n21024);
  and g32971 (n21028, n_14908, n21027);
  not g32972 (n_14909, n21028);
  and g32973 (n21029, n21022, n_14909);
  not g32974 (n_14910, n21019);
  not g32975 (n_14911, n21029);
  and g32976 (n21030, n_14910, n_14911);
  not g32977 (n_14912, n21030);
  and g32978 (n21031, pi0039, n_14912);
  not g32979 (n_14913, n21017);
  not g32980 (n_14914, n21031);
  and g32981 (n21032, n_14913, n_14914);
  not g32982 (n_14915, n21032);
  and g32983 (n21033, n_161, n_14915);
  not g32984 (n_14916, n21033);
  and g32985 (n21034, n21015, n_14916);
  and g32986 (n21035, pi0147, n_14875);
  and g32987 (n21036, n21034, n21035);
  not g32988 (n_14917, pi0726);
  not g32989 (n_14918, n21036);
  and g32990 (n21037, n_14917, n_14918);
  not g32991 (n_14919, n21014);
  and g32992 (n21038, n_14919, n21037);
  and g32993 (n21039, n6236, n17050);
  not g32994 (n_14920, n21039);
  and g32995 (n21040, n_7628, n_14920);
  and g32996 (n21041, n_11723, n16641);
  not g32997 (n_14921, n21041);
  and g32998 (n21042, pi0038, n_14921);
  not g32999 (n_14922, n21040);
  and g33000 (n21043, n_14922, n21042);
  and g33001 (n21044, pi0299, pi0947);
  not g33002 (n_14923, n20902);
  and g33003 (n21045, n17026, n_14923);
  and g33004 (n21046, n_14883, n_14905);
  not g33005 (n_14924, n21046);
  and g33006 (n21047, n_9350, n_14924);
  not g33007 (n_14925, n21047);
  and g33008 (n21048, n_36, n_14925);
  not g33009 (n_14926, n21045);
  and g33010 (n21049, n_14926, n21048);
  not g33011 (n_14927, n20998);
  not g33012 (n_14928, n21049);
  and g33013 (n21050, n_14927, n_14928);
  not g33014 (n_14929, n21050);
  and g33015 (n21051, pi0299, n_14929);
  and g33016 (n21052, n_3149, n16992);
  not g33017 (n_14930, n21052);
  and g33018 (n21053, pi0223, n_14930);
  and g33019 (n21054, n16992, n_14923);
  not g33020 (n_14931, n21054);
  and g33021 (n21055, pi0223, n_14931);
  and g33022 (n21056, n2521, n16654);
  not g33023 (n_14932, n21056);
  and g33024 (n21057, n_11716, n_14932);
  not g33025 (n_14933, n21057);
  and g33026 (n21058, n6236, n_14933);
  not g33027 (n_14934, n21058);
  and g33028 (n21059, n_223, n_14934);
  not g33029 (n_14935, n21053);
  not g33030 (n_14936, n21055);
  and g33031 (n21060, n_14935, n_14936);
  not g33032 (n_14937, n21059);
  and g33033 (n21061, n_14937, n21060);
  not g33034 (n_14938, n21061);
  and g33035 (n21062, n_234, n_14938);
  not g33036 (n_14939, n21044);
  not g33037 (n_14940, n21051);
  and g33038 (n21063, n_14939, n_14940);
  not g33039 (n_14941, n21062);
  and g33040 (n21064, n_14941, n21063);
  and g33041 (n21065, pi0039, n21064);
  and g33042 (n21066, n_11723, n16958);
  not g33043 (n_14942, n21066);
  and g33044 (n21067, n_162, n_14942);
  and g33045 (n21068, n16958, n21067);
  not g33046 (n_14943, n21065);
  not g33047 (n_14944, n21068);
  and g33048 (n21069, n_14943, n_14944);
  and g33049 (n21070, n_7628, n21069);
  and g33050 (n21071, n_11723, n17024);
  and g33051 (n21072, n_234, n21071);
  and g33052 (n21073, pi0215, n_11729);
  and g33053 (n21074, n_11723, n16653);
  and g33054 (n21075, n3448, n21074);
  not g33055 (n_14945, n21075);
  and g33056 (n21076, n_36, n_14945);
  and g33057 (n21077, n_11725, n21076);
  not g33058 (n_14946, n21073);
  and g33059 (n21078, pi0299, n_14946);
  not g33060 (n_14947, n21077);
  and g33061 (n21079, n_14947, n21078);
  not g33062 (n_14948, n21072);
  not g33063 (n_14949, n21079);
  and g33064 (n21080, n_14948, n_14949);
  and g33065 (n21081, pi0039, n21080);
  not g33066 (n_14950, n21067);
  not g33067 (n_14951, n21081);
  and g33068 (n21082, n_14950, n_14951);
  and g33069 (n21083, pi0147, n21082);
  not g33070 (n_14952, n21083);
  and g33071 (n21084, n_161, n_14952);
  not g33072 (n_14953, n21070);
  and g33073 (n21085, n_14953, n21084);
  not g33074 (n_14954, n21043);
  and g33075 (n21086, n_14875, n_14954);
  not g33076 (n_14955, n21085);
  and g33077 (n21087, n_14955, n21086);
  and g33078 (n21088, n_7628, n_11418);
  and g33079 (n21089, n16641, n20902);
  not g33080 (n_14956, n21089);
  and g33081 (n21090, pi0038, n_14956);
  not g33082 (n_14957, n21088);
  and g33083 (n21091, n_14957, n21090);
  and g33084 (n21092, n_14904, n_14929);
  not g33085 (n_14958, n21092);
  and g33086 (n21093, pi0299, n_14958);
  and g33087 (n21094, n_14923, n20990);
  not g33088 (n_14959, n21093);
  not g33089 (n_14960, n21094);
  and g33090 (n21095, n_14959, n_14960);
  not g33091 (n_14961, n21095);
  and g33092 (n21096, pi0039, n_14961);
  and g33093 (n21097, n16958, n_14923);
  and g33094 (n21098, n_162, n21097);
  not g33095 (n_14962, n21096);
  not g33096 (n_14963, n21098);
  and g33097 (n21099, n_14962, n_14963);
  and g33098 (n21100, n_7628, n21099);
  and g33099 (n21101, pi0215, n_14888);
  and g33100 (n21102, n_9350, n_14884);
  and g33101 (n21103, pi0907, n16653);
  and g33102 (n21104, n_3149, n21103);
  not g33103 (n_14964, n21104);
  and g33104 (n21105, n3448, n_14964);
  not g33105 (n_14965, n21102);
  not g33106 (n_14966, n21105);
  and g33107 (n21106, n_14965, n_14966);
  not g33108 (n_14967, n21106);
  and g33109 (n21107, n_36, n_14967);
  not g33110 (n_14968, n21101);
  not g33111 (n_14969, n21107);
  and g33112 (n21108, n_14968, n_14969);
  not g33113 (n_14970, n21108);
  and g33114 (n21109, pi0299, n_14970);
  and g33115 (n21110, n17024, n20902);
  not g33116 (n_14971, n21110);
  and g33117 (n21111, n_234, n_14971);
  not g33118 (n_14972, n21109);
  not g33119 (n_14973, n21111);
  and g33120 (n21112, n_14972, n_14973);
  not g33121 (n_14974, n21112);
  and g33122 (n21113, pi0039, n_14974);
  and g33123 (n21114, n16958, n20902);
  not g33124 (n_14975, n21114);
  and g33125 (n21115, n_162, n_14975);
  not g33126 (n_14976, n21113);
  not g33127 (n_14977, n21115);
  and g33128 (n21116, n_14976, n_14977);
  and g33129 (n21117, pi0147, n21116);
  not g33130 (n_14978, n21117);
  and g33131 (n21118, n_161, n_14978);
  not g33132 (n_14979, n21100);
  and g33133 (n21119, n_14979, n21118);
  not g33134 (n_14980, n21091);
  and g33135 (n21120, pi0770, n_14980);
  not g33136 (n_14981, n21119);
  and g33137 (n21121, n_14981, n21120);
  not g33138 (n_14982, n21087);
  and g33139 (n21122, pi0726, n_14982);
  not g33140 (n_14983, n21121);
  and g33141 (n21123, n_14983, n21122);
  not g33142 (n_14984, n21123);
  and g33143 (n21124, n10197, n_14984);
  not g33144 (n_14985, n21038);
  and g33145 (n21125, n_14985, n21124);
  not g33146 (n_14986, n20987);
  and g33147 (n21126, n_12415, n_14986);
  not g33148 (n_14987, n21125);
  and g33149 (n21127, n_14987, n21126);
  not g33150 (n_14988, n20986);
  not g33151 (n_14989, n21127);
  and g33152 (po0304, n_14988, n_14989);
  and g33153 (n21129, pi0057, pi0148);
  and g33154 (n21130, n2571, n6305);
  not g33155 (n_14990, n21130);
  and g33156 (n21131, n_1865, n_14990);
  and g33157 (n21132, n_12661, pi0947);
  not g33158 (n_14991, n21132);
  and g33159 (n21133, n21041, n_14991);
  and g33160 (n21134, n_1865, n_11418);
  not g33161 (n_14992, n21133);
  not g33162 (n_14993, n21134);
  and g33163 (n21135, n_14992, n_14993);
  not g33164 (n_14994, n21135);
  and g33165 (n21136, pi0038, n_14994);
  and g33166 (n21137, n_11734, n_14972);
  not g33167 (n_14995, n21137);
  and g33168 (n21138, pi0148, n_14995);
  and g33169 (n21139, n_6259, n_14961);
  not g33170 (n_14996, n21138);
  and g33171 (n21140, n_12661, n_14996);
  not g33172 (n_14997, n21139);
  and g33173 (n21141, n_14997, n21140);
  and g33174 (n21142, n_1865, n21064);
  and g33175 (n21143, pi0148, n21080);
  not g33176 (n_14998, n21143);
  and g33177 (n21144, pi0749, n_14998);
  not g33178 (n_14999, n21142);
  and g33179 (n21145, n_14999, n21144);
  not g33180 (n_15000, n21141);
  and g33181 (n21146, pi0039, n_15000);
  not g33182 (n_15001, n21145);
  and g33183 (n21147, n_15001, n21146);
  and g33184 (n21148, n_1865, n_11674);
  not g33185 (n_15002, n21148);
  and g33186 (n21149, n_162, n_15002);
  and g33187 (n21150, n21066, n_14991);
  not g33188 (n_15003, n21150);
  and g33189 (n21151, n21149, n_15003);
  not g33190 (n_15004, n21151);
  and g33191 (n21152, n_161, n_15004);
  not g33192 (n_15005, n21147);
  and g33193 (n21153, n_15005, n21152);
  not g33194 (n_15006, n21136);
  and g33195 (n21154, pi0706, n_15006);
  not g33196 (n_15007, n21153);
  and g33197 (n21155, n_15007, n21154);
  and g33198 (n21156, pi0749, pi0947);
  and g33199 (n21157, n16958, n21156);
  not g33200 (n_15008, n21157);
  and g33201 (n21158, n21149, n_15008);
  and g33202 (n21159, n_1865, n_12661);
  and g33203 (n21160, n_11736, n21159);
  and g33204 (n21161, n_1865, n_14891);
  and g33205 (n21162, n_14904, n_14909);
  not g33206 (n_15009, n21162);
  and g33207 (n21163, pi0148, n_15009);
  not g33208 (n_15010, n21163);
  and g33209 (n21164, pi0299, n_15010);
  not g33210 (n_15011, n21161);
  and g33211 (n21165, n_15011, n21164);
  and g33212 (n21166, n_1865, n_11719);
  not g33213 (n_15012, n21166);
  and g33214 (n21167, n21019, n_15012);
  not g33215 (n_15013, n21167);
  and g33216 (n21168, pi0749, n_15013);
  not g33217 (n_15014, n21165);
  and g33218 (n21169, n_15014, n21168);
  not g33219 (n_15015, n21160);
  and g33220 (n21170, pi0039, n_15015);
  not g33221 (n_15016, n21169);
  and g33222 (n21171, n_15016, n21170);
  not g33223 (n_15017, n21158);
  and g33224 (n21172, n_161, n_15017);
  not g33225 (n_15018, n21171);
  and g33226 (n21173, n_15018, n21172);
  not g33227 (n_15019, n21156);
  and g33228 (n21174, n16641, n_15019);
  and g33229 (n21175, pi0148, n_11740);
  not g33230 (n_15020, n21174);
  and g33231 (n21176, pi0038, n_15020);
  not g33232 (n_15021, n21175);
  and g33233 (n21177, n_15021, n21176);
  not g33234 (n_15022, n21177);
  and g33235 (n21178, n_12614, n_15022);
  not g33236 (n_15023, n21173);
  and g33237 (n21179, n_15023, n21178);
  not g33238 (n_15024, n21179);
  and g33239 (n21180, n21130, n_15024);
  not g33240 (n_15025, n21155);
  and g33241 (n21181, n_15025, n21180);
  not g33242 (n_15026, n21131);
  and g33243 (n21182, n_796, n_15026);
  not g33244 (n_15027, n21181);
  and g33245 (n21183, n_15027, n21182);
  not g33246 (n_15028, n21129);
  and g33247 (n21184, n_12415, n_15028);
  not g33248 (n_15029, n21183);
  and g33249 (n21185, n_15029, n21184);
  and g33250 (n21186, pi0706, n20902);
  and g33251 (n21187, n2926, n_15019);
  not g33252 (n_15030, n21186);
  and g33253 (n21188, n_15030, n21187);
  and g33254 (n21189, pi0148, n_12418);
  not g33255 (n_15031, n21189);
  and g33256 (n21190, pi0832, n_15031);
  not g33257 (n_15032, n21188);
  and g33258 (n21191, n_15032, n21190);
  or g33259 (po0305, n21185, n21191);
  and g33260 (n21193, n_5685, n_12418);
  not g33261 (n_15034, pi0755);
  and g33262 (n21194, n_15034, pi0947);
  not g33263 (n_15036, pi0725);
  and g33264 (n21195, n_15036, n20902);
  not g33265 (n_15037, n21194);
  not g33266 (n_15038, n21195);
  and g33267 (n21196, n_15037, n_15038);
  not g33268 (n_15039, n21196);
  and g33269 (n21197, n2926, n_15039);
  not g33270 (n_15040, n21193);
  and g33271 (n21198, pi0832, n_15040);
  not g33272 (n_15041, n21197);
  and g33273 (n21199, n_15041, n21198);
  and g33274 (n21200, n_5685, n_14814);
  and g33275 (n21201, n16641, n_15037);
  and g33276 (n21202, pi0149, n_11740);
  not g33277 (n_15042, n21201);
  and g33278 (n21203, pi0038, n_15042);
  not g33279 (n_15043, n21202);
  and g33280 (n21204, n_15043, n21203);
  and g33281 (n21205, n_5685, n_11674);
  and g33282 (n21206, n16958, n21194);
  not g33283 (n_15044, n21205);
  and g33284 (n21207, n_162, n_15044);
  not g33285 (n_15045, n21206);
  and g33286 (n21208, n_15045, n21207);
  and g33287 (n21209, n_5685, n_11719);
  not g33288 (n_15046, n21209);
  and g33289 (n21210, n21019, n_15046);
  and g33290 (n21211, n_5685, n_14891);
  and g33291 (n21212, n_10987, n_14911);
  not g33292 (n_15047, n21211);
  not g33293 (n_15048, n21212);
  and g33294 (n21213, n_15047, n_15048);
  not g33295 (n_15049, n21210);
  and g33296 (n21214, n_15034, n_15049);
  not g33297 (n_15050, n21213);
  and g33298 (n21215, n_15050, n21214);
  and g33299 (n21216, n_5685, pi0755);
  and g33300 (n21217, n_11736, n21216);
  not g33301 (n_15051, n21217);
  and g33302 (n21218, pi0039, n_15051);
  not g33303 (n_15052, n21215);
  and g33304 (n21219, n_15052, n21218);
  not g33305 (n_15053, n21208);
  and g33306 (n21220, n_161, n_15053);
  not g33307 (n_15054, n21219);
  and g33308 (n21221, n_15054, n21220);
  not g33309 (n_15055, n21204);
  not g33310 (n_15056, n21221);
  and g33311 (n21222, n_15055, n_15056);
  not g33312 (n_15057, n21222);
  and g33313 (n21223, pi0725, n_15057);
  and g33314 (n21224, n_14975, n21208);
  and g33315 (n21225, n_5685, n21064);
  and g33316 (n21226, pi0149, n21080);
  not g33317 (n_15058, n21226);
  and g33318 (n21227, n_15034, n_15058);
  not g33319 (n_15059, n21225);
  and g33320 (n21228, n_15059, n21227);
  and g33321 (n21229, n_5685, n21093);
  and g33322 (n21230, pi0149, n_14995);
  not g33328 (n_15062, n21233);
  and g33329 (n21234, pi0039, n_15062);
  not g33330 (n_15063, n21228);
  and g33331 (n21235, n_15063, n21234);
  not g33332 (n_15064, n21224);
  not g33333 (n_15065, n21235);
  and g33334 (n21236, n_15064, n_15065);
  not g33335 (n_15066, n21236);
  and g33336 (n21237, n_161, n_15066);
  and g33337 (n21238, n_5685, n_11418);
  and g33338 (n21239, n_11723, n16667);
  and g33339 (n21240, pi0755, pi0947);
  not g33340 (n_15067, n21240);
  and g33341 (n21241, n_162, n_15067);
  and g33342 (n21242, n21239, n21241);
  not g33343 (n_15068, n21238);
  and g33344 (n21243, pi0038, n_15068);
  not g33345 (n_15069, n21242);
  and g33346 (n21244, n_15069, n21243);
  not g33347 (n_15070, n21244);
  and g33348 (n21245, n_15036, n_15070);
  not g33349 (n_15071, n21237);
  and g33350 (n21246, n_15071, n21245);
  not g33351 (n_15072, n21223);
  not g33352 (n_15073, n21246);
  and g33353 (n21247, n_15072, n_15073);
  not g33354 (n_15074, n21247);
  and g33355 (n21248, n10197, n_15074);
  not g33356 (n_15075, n21200);
  and g33357 (n21249, n_12415, n_15075);
  not g33358 (n_15076, n21248);
  and g33359 (n21250, n_15076, n21249);
  not g33360 (n_15077, n21199);
  not g33361 (n_15078, n21250);
  and g33362 (po0306, n_15077, n_15078);
  and g33363 (n21252, n_9109, n_14814);
  and g33364 (n21253, pi0150, n_11740);
  not g33365 (n_15080, pi0751);
  and g33366 (n21254, n_15080, pi0947);
  not g33367 (n_15081, n21254);
  and g33368 (n21255, n16641, n_15081);
  not g33369 (n_15082, n21253);
  not g33370 (n_15083, n21255);
  and g33371 (n21256, n_15082, n_15083);
  not g33372 (n_15084, n21256);
  and g33373 (n21257, pi0038, n_15084);
  and g33374 (n21258, pi0150, n_11674);
  and g33375 (n21259, pi0751, n16958);
  not g33376 (n_15085, n21258);
  not g33377 (n_15086, n21259);
  and g33378 (n21260, n_15085, n_15086);
  and g33379 (n21261, n20989, n21260);
  and g33380 (n21262, n_9109, n21004);
  and g33381 (n21263, pi0150, n_14912);
  not g33382 (n_15087, n21263);
  and g33383 (n21264, n_15080, n_15087);
  not g33384 (n_15088, n21262);
  and g33385 (n21265, n_15088, n21264);
  and g33386 (n21266, n_9109, pi0751);
  and g33387 (n21267, n_11736, n21266);
  not g33388 (n_15089, n21265);
  not g33389 (n_15090, n21267);
  and g33390 (n21268, n_15089, n_15090);
  not g33391 (n_15091, n21268);
  and g33392 (n21269, pi0039, n_15091);
  not g33393 (n_15092, n21261);
  and g33394 (n21270, n_161, n_15092);
  not g33395 (n_15093, n21269);
  and g33396 (n21271, n_15093, n21270);
  not g33397 (n_15095, n21257);
  and g33398 (n21272, pi0701, n_15095);
  not g33399 (n_15096, n21271);
  and g33400 (n21273, n_15096, n21272);
  and g33401 (n21274, n_9109, n_11418);
  and g33402 (n21275, pi0751, pi0947);
  not g33403 (n_15097, n21275);
  and g33404 (n21276, n_162, n_15097);
  and g33405 (n21277, n21239, n21276);
  not g33406 (n_15098, n21274);
  and g33407 (n21278, pi0038, n_15098);
  not g33408 (n_15099, n21277);
  and g33409 (n21279, n_15099, n21278);
  and g33410 (n21280, n21097, n_15081);
  and g33411 (n21281, n_162, n_15085);
  not g33412 (n_15100, n21280);
  and g33413 (n21282, n_15100, n21281);
  and g33414 (n21283, n_9109, n_14961);
  and g33415 (n21284, pi0150, n_14974);
  not g33416 (n_15101, n21284);
  and g33417 (n21285, pi0751, n_15101);
  not g33418 (n_15102, n21283);
  and g33419 (n21286, n_15102, n21285);
  and g33420 (n21287, n_9109, n21064);
  and g33421 (n21288, pi0150, n21080);
  not g33422 (n_15103, n21288);
  and g33423 (n21289, n_15080, n_15103);
  not g33424 (n_15104, n21287);
  and g33425 (n21290, n_15104, n21289);
  not g33426 (n_15105, n21286);
  not g33427 (n_15106, n21290);
  and g33428 (n21291, n_15105, n_15106);
  not g33429 (n_15107, n21291);
  and g33430 (n21292, pi0039, n_15107);
  not g33431 (n_15108, n21282);
  and g33432 (n21293, n_161, n_15108);
  not g33433 (n_15109, n21292);
  and g33434 (n21294, n_15109, n21293);
  not g33435 (n_15110, pi0701);
  not g33436 (n_15111, n21279);
  and g33437 (n21295, n_15110, n_15111);
  not g33438 (n_15112, n21294);
  and g33439 (n21296, n_15112, n21295);
  not g33440 (n_15113, n21273);
  not g33441 (n_15114, n21296);
  and g33442 (n21297, n_15113, n_15114);
  not g33443 (n_15115, n21297);
  and g33444 (n21298, n10197, n_15115);
  not g33445 (n_15116, n21252);
  and g33446 (n21299, n_12415, n_15116);
  not g33447 (n_15117, n21298);
  and g33448 (n21300, n_15117, n21299);
  and g33449 (n21301, n_9109, n_12418);
  and g33450 (n21302, n_15110, n20902);
  not g33451 (n_15118, n21302);
  and g33452 (n21303, n_15081, n_15118);
  not g33453 (n_15119, n21303);
  and g33454 (n21304, n2926, n_15119);
  not g33455 (n_15120, n21301);
  and g33456 (n21305, pi0832, n_15120);
  not g33457 (n_15121, n21304);
  and g33458 (n21306, n_15121, n21305);
  not g33459 (n_15122, n21300);
  not g33460 (n_15123, n21306);
  and g33461 (po0307, n_15122, n_15123);
  and g33462 (n21308, n_983, n_12418);
  not g33463 (n_15125, pi0745);
  and g33464 (n21309, n_15125, pi0947);
  not g33465 (n_15127, pi0723);
  and g33466 (n21310, n_15127, n20902);
  not g33467 (n_15128, n21309);
  not g33468 (n_15129, n21310);
  and g33469 (n21311, n_15128, n_15129);
  not g33470 (n_15130, n21311);
  and g33471 (n21312, n2926, n_15130);
  not g33472 (n_15131, n21308);
  and g33473 (n21313, pi0832, n_15131);
  not g33474 (n_15132, n21312);
  and g33475 (n21314, n_15132, n21313);
  and g33476 (n21315, n_983, n_14814);
  and g33477 (n21316, n_983, n_11418);
  and g33478 (n21317, pi0745, pi0947);
  not g33479 (n_15133, n21317);
  and g33480 (n21318, n_162, n_15133);
  and g33481 (n21319, n21239, n21318);
  not g33482 (n_15134, n21316);
  and g33483 (n21320, pi0038, n_15134);
  not g33484 (n_15135, n21319);
  and g33485 (n21321, n_15135, n21320);
  and g33486 (n21322, n_983, n_11674);
  and g33487 (n21323, n_15125, n21016);
  not g33488 (n_15136, n21322);
  not g33489 (n_15137, n21323);
  and g33490 (n21324, n_15136, n_15137);
  and g33491 (n21325, n21115, n21324);
  and g33492 (n21326, n_11730, n_14888);
  and g33493 (n21327, n_983, n21326);
  not g33494 (n_15138, n21327);
  and g33495 (n21328, n_11729, n_15138);
  not g33496 (n_15139, n21328);
  and g33497 (n21329, pi0215, n_15139);
  and g33498 (n21330, pi0151, n_9350);
  not g33499 (n_15140, n17032);
  and g33500 (n21331, n_15140, n21330);
  not g33501 (n_15141, n21331);
  and g33502 (n21332, n_11726, n_15141);
  and g33503 (n21333, n_983, n_11445);
  not g33504 (n_15142, n21333);
  and g33505 (n21334, n21105, n_15142);
  not g33506 (n_15143, n21074);
  and g33507 (n21335, n_15143, n21334);
  not g33508 (n_15144, n21335);
  and g33509 (n21336, n_36, n_15144);
  and g33510 (n21337, n21332, n21336);
  not g33511 (n_15145, n21329);
  not g33512 (n_15146, n21337);
  and g33513 (n21338, n_15145, n_15146);
  not g33514 (n_15147, n21338);
  and g33515 (n21339, pi0299, n_15147);
  not g33516 (n_15148, n21071);
  and g33517 (n21340, pi0151, n_15148);
  not g33518 (n_15149, n21340);
  and g33519 (n21341, n21062, n_15149);
  not g33520 (n_15150, n21339);
  not g33521 (n_15151, n21341);
  and g33522 (n21342, n_15150, n_15151);
  not g33523 (n_15152, n21342);
  and g33524 (n21343, n_15125, n_15152);
  not g33525 (n_15153, n21334);
  and g33526 (n21344, n21332, n_15153);
  and g33527 (n21345, n21048, n21344);
  not g33528 (n_15154, n21345);
  and g33529 (n21346, n_15145, n_15154);
  not g33530 (n_15155, n21346);
  and g33531 (n21347, n_14904, n_15155);
  not g33532 (n_15156, n21347);
  and g33533 (n21348, pi0299, n_15156);
  and g33534 (n21349, n_983, n_11719);
  not g33535 (n_15157, n21349);
  and g33536 (n21350, n21111, n_15157);
  not g33537 (n_15158, n21350);
  and g33538 (n21351, pi0745, n_15158);
  not g33539 (n_15159, n21348);
  and g33540 (n21352, n_15159, n21351);
  not g33541 (n_15160, n21352);
  and g33542 (n21353, pi0039, n_15160);
  not g33543 (n_15161, n21343);
  and g33544 (n21354, n_15161, n21353);
  not g33545 (n_15162, n21325);
  not g33546 (n_15163, n21354);
  and g33547 (n21355, n_15162, n_15163);
  not g33548 (n_15164, n21355);
  and g33549 (n21356, n_161, n_15164);
  not g33550 (n_15165, n21321);
  and g33551 (n21357, n_15127, n_15165);
  not g33552 (n_15166, n21356);
  and g33553 (n21358, n_15166, n21357);
  and g33554 (n21359, pi0151, n_11740);
  and g33555 (n21360, n16641, n_15128);
  not g33556 (n_15167, n21359);
  not g33557 (n_15168, n21360);
  and g33558 (n21361, n_15167, n_15168);
  not g33559 (n_15169, n21361);
  and g33560 (n21362, pi0038, n_15169);
  not g33561 (n_15170, n21324);
  and g33562 (n21363, n_162, n_15170);
  and g33563 (n21364, n_15125, n_11734);
  and g33564 (n21365, n_983, n_11736);
  not g33565 (n_15171, n21364);
  and g33566 (n21366, n_15171, n21365);
  and g33567 (n21367, n21026, n_15142);
  not g33568 (n_15172, n21367);
  and g33569 (n21368, n21332, n_15172);
  and g33570 (n21369, n20996, n21368);
  and g33571 (n21370, n21101, n_15139);
  not g33572 (n_15173, n21370);
  and g33573 (n21371, pi0299, n_15173);
  not g33574 (n_15174, n21369);
  and g33575 (n21372, n_15174, n21371);
  and g33576 (n21373, n_15125, n_14910);
  not g33577 (n_15175, n21372);
  and g33578 (n21374, n_15175, n21373);
  not g33579 (n_15176, n21366);
  not g33580 (n_15177, n21374);
  and g33581 (n21375, n_15176, n_15177);
  not g33582 (n_15178, n21375);
  and g33583 (n21376, pi0039, n_15178);
  not g33584 (n_15179, n21363);
  and g33585 (n21377, n_161, n_15179);
  not g33586 (n_15180, n21376);
  and g33587 (n21378, n_15180, n21377);
  not g33588 (n_15181, n21362);
  and g33589 (n21379, pi0723, n_15181);
  not g33590 (n_15182, n21378);
  and g33591 (n21380, n_15182, n21379);
  not g33592 (n_15183, n21358);
  not g33593 (n_15184, n21380);
  and g33594 (n21381, n_15183, n_15184);
  not g33595 (n_15185, n21381);
  and g33596 (n21382, n10197, n_15185);
  not g33597 (n_15186, n21315);
  and g33598 (n21383, n_12415, n_15186);
  not g33599 (n_15187, n21382);
  and g33600 (n21384, n_15187, n21383);
  not g33601 (n_15188, n21314);
  not g33602 (n_15189, n21384);
  and g33603 (po0308, n_15188, n_15189);
  and g33604 (n21386, n_263, n_14814);
  and g33605 (n21387, n_263, n_11418);
  and g33606 (n21388, pi0759, pi0947);
  not g33607 (n_15191, n21388);
  and g33608 (n21389, n_162, n_15191);
  and g33609 (n21390, n16667, n_14923);
  and g33610 (n21391, n21389, n21390);
  not g33611 (n_15192, n21387);
  and g33612 (n21392, pi0038, n_15192);
  not g33613 (n_15193, n21391);
  and g33614 (n21393, n_15193, n21392);
  and g33615 (n21394, pi0152, n_11674);
  not g33616 (n_15194, n21389);
  and g33617 (n21395, n_11737, n_15194);
  not g33618 (n_15195, n21394);
  not g33619 (n_15196, n21395);
  and g33620 (n21396, n_15195, n_15196);
  and g33621 (n21397, n_14975, n21396);
  and g33622 (n21398, n_263, n_11729);
  not g33623 (n_15197, n21398);
  and g33624 (n21399, n20998, n_15197);
  and g33625 (n21400, n_14923, n_14946);
  not g33626 (n_15198, n21400);
  and g33627 (n21401, n21399, n_15198);
  and g33628 (n21402, pi0152, n21046);
  not g33629 (n_15199, n21402);
  and g33630 (n21403, n21102, n_15199);
  and g33631 (n21404, pi0152, n_11445);
  not g33632 (n_15200, n21404);
  and g33633 (n21405, n_15143, n_15200);
  and g33634 (n21406, n3448, n21405);
  not g33635 (n_15201, n21406);
  and g33636 (n21407, n_36, n_15201);
  and g33637 (n21408, n_14926, n21407);
  not g33638 (n_15202, n21403);
  and g33639 (n21409, n_15202, n21408);
  not g33640 (n_15203, n21401);
  and g33641 (n21410, pi0299, n_15203);
  not g33642 (n_15204, n21409);
  and g33643 (n21411, n_15204, n21410);
  and g33644 (n21412, n_14964, n_15200);
  not g33645 (n_15205, n21412);
  and g33646 (n21413, n2603, n_15205);
  not g33647 (n_15206, n17020);
  and g33648 (n21414, n_263, n_15206);
  and g33649 (n21415, n17020, n_14923);
  not g33650 (n_15207, n21415);
  and g33651 (n21416, n_9349, n_15207);
  not g33652 (n_15208, n21414);
  and g33653 (n21417, n_15208, n21416);
  not g33654 (n_15209, n21413);
  not g33655 (n_15210, n21417);
  and g33656 (n21418, n_15209, n_15210);
  not g33657 (n_15211, n21418);
  and g33658 (n21419, n_223, n_15211);
  and g33659 (n21420, n_263, n_11697);
  not g33660 (n_15212, n21420);
  and g33661 (n21421, n21055, n_15212);
  not g33662 (n_15213, n21421);
  and g33663 (n21422, n_234, n_15213);
  not g33664 (n_15214, n21419);
  and g33665 (n21423, n_15214, n21422);
  not g33666 (n_15215, pi0759);
  not g33667 (n_15216, n21411);
  and g33668 (n21424, n_15215, n_15216);
  not g33669 (n_15217, n21423);
  and g33670 (n21425, n_15217, n21424);
  and g33671 (n21426, n_15140, n21403);
  not g33672 (n_15218, n21426);
  and g33673 (n21427, n21407, n_15218);
  not g33674 (n_15219, n21399);
  and g33675 (n21428, pi0299, n_15219);
  not g33676 (n_15220, n21427);
  and g33677 (n21429, n_15220, n21428);
  and g33678 (n21430, n2603, n21405);
  and g33679 (n21431, n_3149, n17020);
  not g33680 (n_15221, n21431);
  and g33681 (n21432, n_9349, n_15221);
  and g33682 (n21433, n_15208, n21432);
  and g33683 (n21434, n_11723, n17020);
  not g33684 (n_15222, n21434);
  and g33685 (n21435, n_9349, n_15222);
  not g33686 (n_15223, n21433);
  and g33687 (n21436, n_15223, n21435);
  not g33688 (n_15224, n21430);
  and g33689 (n21437, n_223, n_15224);
  not g33690 (n_15225, n21436);
  and g33691 (n21438, n_15225, n21437);
  and g33692 (n21439, n21053, n_15212);
  not g33693 (n_15226, n21439);
  and g33694 (n21440, n_234, n_15226);
  and g33695 (n21441, n_15213, n21440);
  not g33696 (n_15227, n21438);
  and g33697 (n21442, n_15227, n21441);
  not g33698 (n_15228, n21429);
  and g33699 (n21443, pi0759, n_15228);
  not g33700 (n_15229, n21442);
  and g33701 (n21444, n_15229, n21443);
  not g33702 (n_15230, n21425);
  and g33703 (n21445, pi0039, n_15230);
  not g33704 (n_15231, n21444);
  and g33705 (n21446, n_15231, n21445);
  not g33706 (n_15232, n21397);
  and g33707 (n21447, n_161, n_15232);
  not g33708 (n_15233, n21446);
  and g33709 (n21448, n_15233, n21447);
  not g33710 (n_15235, n21393);
  and g33711 (n21449, pi0696, n_15235);
  not g33712 (n_15236, n21448);
  and g33713 (n21450, n_15236, n21449);
  and g33714 (n21451, n_263, n_11740);
  and g33715 (n21452, n16641, n_15191);
  not g33716 (n_15237, n21452);
  and g33717 (n21453, pi0038, n_15237);
  not g33718 (n_15238, n21451);
  and g33719 (n21454, n_15238, n21453);
  and g33720 (n21455, n_14906, n_15200);
  not g33721 (n_15239, n21455);
  and g33722 (n21456, n2603, n_15239);
  not g33723 (n_15240, n21456);
  and g33724 (n21457, n_15223, n_15240);
  not g33725 (n_15241, n21457);
  and g33726 (n21458, n_223, n_15241);
  not g33727 (n_15242, n21458);
  and g33728 (n21459, n21440, n_15242);
  and g33729 (n21460, pi0152, n21000);
  and g33730 (n21461, n3448, n21455);
  and g33731 (n21462, n_14886, n_15202);
  not g33732 (n_15243, n21462);
  and g33733 (n21463, n_14905, n_15243);
  not g33734 (n_15244, n21461);
  and g33735 (n21464, n_36, n_15244);
  not g33736 (n_15245, n21463);
  and g33737 (n21465, n_15245, n21464);
  not g33738 (n_15246, n21460);
  and g33739 (n21466, n21022, n_15246);
  not g33740 (n_15247, n21465);
  and g33741 (n21467, n_15247, n21466);
  not g33742 (n_15248, n21459);
  and g33743 (n21468, pi0759, n_15248);
  not g33744 (n_15249, n21467);
  and g33745 (n21469, n_15249, n21468);
  and g33746 (n21470, n_15215, n_11736);
  and g33747 (n21471, pi0152, n21470);
  not g33748 (n_15250, n21471);
  and g33749 (n21472, pi0039, n_15250);
  not g33750 (n_15251, n21469);
  and g33751 (n21473, n_15251, n21472);
  not g33752 (n_15252, n21396);
  and g33753 (n21474, n_161, n_15252);
  not g33754 (n_15253, n21473);
  and g33755 (n21475, n_15253, n21474);
  not g33756 (n_15254, pi0696);
  not g33757 (n_15255, n21454);
  and g33758 (n21476, n_15254, n_15255);
  not g33759 (n_15256, n21475);
  and g33760 (n21477, n_15256, n21476);
  not g33761 (n_15257, n21450);
  not g33762 (n_15258, n21477);
  and g33763 (n21478, n_15257, n_15258);
  not g33764 (n_15259, n21478);
  and g33765 (n21479, n10197, n_15259);
  not g33766 (n_15260, n21386);
  and g33767 (n21480, n_12415, n_15260);
  not g33768 (n_15261, n21479);
  and g33769 (n21481, n_15261, n21480);
  and g33770 (n21482, n_263, n_12418);
  and g33771 (n21483, pi0696, n20902);
  and g33772 (n21484, n2926, n_15191);
  not g33773 (n_15262, n21483);
  and g33774 (n21485, n_15262, n21484);
  not g33775 (n_15263, n21482);
  and g33776 (n21486, pi0832, n_15263);
  not g33777 (n_15264, n21485);
  and g33778 (n21487, n_15264, n21486);
  or g33779 (po0309, n21481, n21487);
  and g33780 (n21489, pi0153, n_12418);
  and g33781 (n21490, pi0766, pi0947);
  not g33782 (n_15266, n21490);
  and g33783 (n21491, n2926, n_15266);
  and g33784 (n21492, pi0700, n20902);
  not g33785 (n_15268, n21492);
  and g33786 (n21493, n21491, n_15268);
  not g33787 (n_15269, n21489);
  and g33788 (n21494, pi0832, n_15269);
  not g33789 (n_15270, n21493);
  and g33790 (n21495, n_15270, n21494);
  and g33791 (n21496, pi0057, pi0153);
  and g33792 (n21497, n_187, n_14990);
  and g33793 (n21498, n_187, n_11674);
  not g33794 (n_15271, pi0766);
  and g33795 (n21499, n_15271, n18147);
  not g33796 (n_15272, n21499);
  and g33797 (n21500, n_14913, n_15272);
  not g33798 (n_15273, n21498);
  not g33799 (n_15274, n21500);
  and g33800 (n21501, n_15273, n_15274);
  and g33801 (n21502, n_14975, n21501);
  and g33802 (n21503, n_187, n_11719);
  not g33803 (n_15275, n21503);
  and g33804 (n21504, n21111, n_15275);
  and g33805 (n21505, pi0153, n_11729);
  not g33806 (n_15276, n21505);
  and g33807 (n21506, n20998, n_15276);
  not g33808 (n_15277, n21506);
  and g33809 (n21507, n21073, n_15277);
  and g33810 (n21508, pi0153, n_9350);
  and g33811 (n21509, n_15140, n21508);
  not g33812 (n_15278, n21509);
  and g33813 (n21510, n_11726, n_15278);
  and g33814 (n21511, n_187, n_11445);
  not g33815 (n_15279, n21511);
  and g33816 (n21512, n21105, n_15279);
  not g33817 (n_15280, n21512);
  and g33818 (n21513, n_14925, n_15280);
  and g33819 (n21514, n21510, n21513);
  not g33820 (n_15281, n21514);
  and g33821 (n21515, n_36, n_15281);
  not g33822 (n_15282, n21507);
  and g33823 (n21516, n_14904, n_15282);
  not g33824 (n_15283, n21515);
  and g33825 (n21517, n_15283, n21516);
  not g33826 (n_15284, n21517);
  and g33827 (n21518, pi0299, n_15284);
  not g33828 (n_15285, n21504);
  and g33829 (n21519, n_15271, n_15285);
  not g33830 (n_15286, n21518);
  and g33831 (n21520, n_15286, n21519);
  and g33832 (n21521, n21026, n_15279);
  not g33833 (n_15287, n21103);
  and g33834 (n21522, n_15287, n21521);
  not g33835 (n_15288, n21522);
  and g33836 (n21523, n_36, n_15288);
  and g33837 (n21524, n21510, n21523);
  not g33838 (n_15289, n21524);
  and g33839 (n21525, n_15277, n_15289);
  not g33840 (n_15290, n21525);
  and g33841 (n21526, pi0299, n_15290);
  and g33842 (n21527, pi0153, n_15148);
  not g33843 (n_15291, n21527);
  and g33844 (n21528, n21062, n_15291);
  not g33845 (n_15292, n21526);
  not g33846 (n_15293, n21528);
  and g33847 (n21529, n_15292, n_15293);
  not g33848 (n_15294, n21529);
  and g33849 (n21530, pi0766, n_15294);
  not g33850 (n_15295, n21520);
  and g33851 (n21531, pi0039, n_15295);
  not g33852 (n_15296, n21530);
  and g33853 (n21532, n_15296, n21531);
  not g33854 (n_15297, n21502);
  not g33855 (n_15298, n21532);
  and g33856 (n21533, n_15297, n_15298);
  not g33857 (n_15299, n21533);
  and g33858 (n21534, n_161, n_15299);
  and g33859 (n21535, n_187, n_11418);
  and g33860 (n21536, n_15271, pi0947);
  not g33861 (n_15300, n21536);
  and g33862 (n21537, n_162, n_15300);
  and g33863 (n21538, n21239, n21537);
  not g33864 (n_15301, n21535);
  and g33865 (n21539, pi0038, n_15301);
  not g33866 (n_15302, n21538);
  and g33867 (n21540, n_15302, n21539);
  not g33868 (n_15303, n21534);
  not g33869 (n_15304, n21540);
  and g33870 (n21541, n_15303, n_15304);
  not g33871 (n_15305, n21541);
  and g33872 (n21542, pi0700, n_15305);
  and g33873 (n21543, n6284, n21491);
  and g33874 (n21544, pi0153, n_11740);
  not g33875 (n_15306, n21543);
  and g33876 (n21545, pi0038, n_15306);
  not g33877 (n_15307, n21544);
  and g33878 (n21546, n_15307, n21545);
  and g33879 (n21547, n21019, n_15275);
  and g33880 (n21548, n21000, n_15276);
  not g33881 (n_15308, n21521);
  and g33882 (n21549, n21510, n_15308);
  and g33883 (n21550, n20996, n21549);
  not g33884 (n_15309, n21548);
  and g33885 (n21551, pi0299, n_15309);
  not g33886 (n_15310, n21550);
  and g33887 (n21552, n_15310, n21551);
  not g33888 (n_15311, n21552);
  and g33889 (n21553, pi0766, n_15311);
  not g33890 (n_15312, n21547);
  and g33891 (n21554, n_15312, n21553);
  and g33892 (n21555, n_187, n_15271);
  and g33893 (n21556, n_11736, n21555);
  not g33894 (n_15313, n21556);
  and g33895 (n21557, pi0039, n_15313);
  not g33896 (n_15314, n21554);
  and g33897 (n21558, n_15314, n21557);
  not g33898 (n_15315, n21501);
  and g33899 (n21559, n_161, n_15315);
  not g33900 (n_15316, n21558);
  and g33901 (n21560, n_15316, n21559);
  not g33902 (n_15317, pi0700);
  not g33903 (n_15318, n21546);
  and g33904 (n21561, n_15317, n_15318);
  not g33905 (n_15319, n21560);
  and g33906 (n21562, n_15319, n21561);
  not g33907 (n_15320, n21562);
  and g33908 (n21563, n21130, n_15320);
  not g33909 (n_15321, n21542);
  and g33910 (n21564, n_15321, n21563);
  not g33911 (n_15322, n21497);
  and g33912 (n21565, n_796, n_15322);
  not g33913 (n_15323, n21564);
  and g33914 (n21566, n_15323, n21565);
  not g33915 (n_15324, n21496);
  and g33916 (n21567, n_12415, n_15324);
  not g33917 (n_15325, n21566);
  and g33918 (n21568, n_15325, n21567);
  or g33919 (po0310, n21495, n21568);
  and g33920 (n21570, n_820, n_12418);
  not g33921 (n_15327, pi0742);
  and g33922 (n21571, n_15327, pi0947);
  not g33923 (n_15329, pi0704);
  and g33924 (n21572, n_15329, n20902);
  not g33925 (n_15330, n21571);
  not g33926 (n_15331, n21572);
  and g33927 (n21573, n_15330, n_15331);
  not g33928 (n_15332, n21573);
  and g33929 (n21574, n2926, n_15332);
  not g33930 (n_15333, n21570);
  and g33931 (n21575, pi0832, n_15333);
  not g33932 (n_15334, n21574);
  and g33933 (n21576, n_15334, n21575);
  and g33934 (n21577, n_820, n_14814);
  and g33935 (n21578, n_820, n_11418);
  not g33936 (n_15335, n21578);
  and g33937 (n21579, n21090, n_15335);
  and g33938 (n21580, n_820, n_11674);
  not g33939 (n_15336, n21580);
  and g33940 (n21581, n21115, n_15336);
  and g33941 (n21582, n_820, n21095);
  and g33942 (n21583, pi0154, n21112);
  not g33943 (n_15337, n21583);
  and g33944 (n21584, pi0039, n_15337);
  not g33945 (n_15338, n21582);
  and g33946 (n21585, n_15338, n21584);
  not g33947 (n_15339, n21581);
  not g33948 (n_15340, n21585);
  and g33949 (n21586, n_15339, n_15340);
  not g33950 (n_15341, n21586);
  and g33951 (n21587, n_161, n_15341);
  not g33952 (n_15342, n21579);
  and g33953 (n21588, pi0742, n_15342);
  not g33954 (n_15343, n21587);
  and g33955 (n21589, n_15343, n21588);
  and g33956 (n21590, n21042, n_15335);
  and g33957 (n21591, n_14942, n21581);
  not g33958 (n_15344, n21064);
  and g33959 (n21592, n_820, n_15344);
  not g33960 (n_15345, n21080);
  and g33961 (n21593, pi0154, n_15345);
  not g33962 (n_15346, n21593);
  and g33963 (n21594, pi0039, n_15346);
  not g33964 (n_15347, n21592);
  and g33965 (n21595, n_15347, n21594);
  not g33966 (n_15348, n21591);
  not g33967 (n_15349, n21595);
  and g33968 (n21596, n_15348, n_15349);
  not g33969 (n_15350, n21596);
  and g33970 (n21597, n_161, n_15350);
  not g33971 (n_15351, n21590);
  and g33972 (n21598, n_15327, n_15351);
  not g33973 (n_15352, n21597);
  and g33974 (n21599, n_15352, n21598);
  not g33975 (n_15353, n21589);
  and g33976 (n21600, n_15329, n_15353);
  not g33977 (n_15354, n21599);
  and g33978 (n21601, n_15354, n21600);
  and g33979 (n21602, n_820, n_11740);
  not g33980 (n_15355, n21015);
  not g33981 (n_15356, n21602);
  and g33982 (n21603, n_15355, n_15356);
  and g33983 (n21604, n21017, n_15336);
  and g33984 (n21605, pi0154, n21030);
  and g33985 (n21606, n_820, n_14894);
  not g33986 (n_15357, n21605);
  and g33987 (n21607, pi0039, n_15357);
  not g33988 (n_15358, n21606);
  and g33989 (n21608, n_15358, n21607);
  not g33990 (n_15359, n21604);
  not g33991 (n_15360, n21608);
  and g33992 (n21609, n_15359, n_15360);
  not g33993 (n_15361, n21609);
  and g33994 (n21610, n_161, n_15361);
  not g33995 (n_15362, n21603);
  and g33996 (n21611, n_15327, n_15362);
  not g33997 (n_15363, n21610);
  and g33998 (n21612, n_15363, n21611);
  and g33999 (n21613, n_820, pi0742);
  and g34000 (n21614, n_11743, n21613);
  not g34001 (n_15364, n21614);
  and g34002 (n21615, pi0704, n_15364);
  not g34003 (n_15365, n21612);
  and g34004 (n21616, n_15365, n21615);
  not g34005 (n_15366, n21616);
  and g34006 (n21617, n10197, n_15366);
  not g34007 (n_15367, n21601);
  and g34008 (n21618, n_15367, n21617);
  not g34009 (n_15368, n21577);
  and g34010 (n21619, n_12415, n_15368);
  not g34011 (n_15369, n21618);
  and g34012 (n21620, n_15369, n21619);
  not g34013 (n_15370, n21576);
  not g34014 (n_15371, n21620);
  and g34015 (po0311, n_15370, n_15371);
  not g34016 (n_15373, pi0757);
  and g34017 (n21622, n_15373, n21034);
  not g34018 (n_15375, n21622);
  and g34019 (n21623, pi0686, n_15375);
  not g34020 (n_15376, n21082);
  and g34021 (n21624, n_161, n_15376);
  not g34022 (n_15377, n21042);
  not g34023 (n_15378, n21624);
  and g34024 (n21625, n_15377, n_15378);
  and g34025 (n21626, n_15373, n21625);
  not g34026 (n_15379, n21116);
  and g34027 (n21627, n_161, n_15379);
  not g34028 (n_15380, n21090);
  not g34029 (n_15381, n21627);
  and g34030 (n21628, n_15380, n_15381);
  and g34031 (n21629, pi0757, n21628);
  not g34032 (n_15382, pi0686);
  not g34033 (n_15383, n21626);
  and g34034 (n21630, n_15382, n_15383);
  not g34035 (n_15384, n21629);
  and g34036 (n21631, n_15384, n21630);
  not g34037 (n_15385, n21623);
  and g34038 (n21632, n10197, n_15385);
  not g34039 (n_15386, n21631);
  and g34040 (n21633, n_15386, n21632);
  not g34041 (n_15387, n21633);
  and g34042 (n21634, pi0155, n_15387);
  not g34043 (n_15388, n21069);
  and g34044 (n21635, n_161, n_15388);
  and g34045 (n21636, pi0038, n21039);
  not g34046 (n_15389, n21635);
  not g34047 (n_15390, n21636);
  and g34048 (n21637, n_15389, n_15390);
  and g34049 (n21638, n_15373, n21637);
  not g34050 (n_15391, n21099);
  and g34051 (n21639, n_161, n_15391);
  and g34052 (n21640, n16641, n21090);
  not g34053 (n_15392, n21639);
  not g34054 (n_15393, n21640);
  and g34055 (n21641, n_15392, n_15393);
  and g34056 (n21642, pi0757, n21641);
  not g34057 (n_15394, n21638);
  and g34058 (n21643, n_15382, n_15394);
  not g34059 (n_15395, n21642);
  and g34060 (n21644, n_15395, n21643);
  and g34061 (n21645, n_15373, n21010);
  and g34062 (n21646, pi0757, n_11743);
  not g34063 (n_15396, n21646);
  and g34064 (n21647, pi0686, n_15396);
  not g34065 (n_15397, n21645);
  and g34066 (n21648, n_15397, n21647);
  not g34067 (n_15398, n21644);
  not g34068 (n_15399, n21648);
  and g34069 (n21649, n_15398, n_15399);
  and g34070 (n21650, n_6284, n10197);
  not g34071 (n_15400, n21649);
  and g34072 (n21651, n_15400, n21650);
  not g34073 (n_15401, n21634);
  not g34074 (n_15402, n21651);
  and g34075 (n21652, n_15401, n_15402);
  not g34076 (n_15403, n21652);
  and g34077 (n21653, n_12415, n_15403);
  and g34078 (n21654, n_6284, n_12418);
  and g34079 (n21655, n_15373, pi0947);
  and g34080 (n21656, n_15382, n20902);
  not g34081 (n_15404, n21655);
  not g34082 (n_15405, n21656);
  and g34083 (n21657, n_15404, n_15405);
  not g34084 (n_15406, n21657);
  and g34085 (n21658, n2926, n_15406);
  not g34086 (n_15407, n21654);
  and g34087 (n21659, pi0832, n_15407);
  not g34088 (n_15408, n21658);
  and g34089 (n21660, n_15408, n21659);
  not g34090 (n_15409, n21653);
  not g34091 (n_15410, n21660);
  and g34092 (po0312, n_15409, n_15410);
  and g34093 (n21662, n_7638, n_12418);
  not g34094 (n_15412, pi0741);
  and g34095 (n21663, n_15412, pi0947);
  not g34096 (n_15414, pi0724);
  and g34097 (n21664, n_15414, n20902);
  not g34098 (n_15415, n21663);
  not g34099 (n_15416, n21664);
  and g34100 (n21665, n_15415, n_15416);
  not g34101 (n_15417, n21665);
  and g34102 (n21666, n2926, n_15417);
  not g34103 (n_15418, n21662);
  and g34104 (n21667, pi0832, n_15418);
  not g34105 (n_15419, n21666);
  and g34106 (n21668, n_15419, n21667);
  not g34107 (n_15420, n21637);
  and g34108 (n21669, n_15412, n_15420);
  not g34109 (n_15421, n21641);
  and g34110 (n21670, pi0741, n_15421);
  not g34111 (n_15422, n21669);
  and g34112 (n21671, n_15414, n_15422);
  not g34113 (n_15423, n21670);
  and g34114 (n21672, n_15423, n21671);
  not g34115 (n_15424, n21010);
  and g34116 (n21673, n_15412, n_15424);
  and g34117 (n21674, pi0741, n17052);
  not g34118 (n_15425, n21674);
  and g34119 (n21675, pi0724, n_15425);
  not g34120 (n_15426, n21673);
  and g34121 (n21676, n_15426, n21675);
  not g34122 (n_15427, n21676);
  and g34123 (n21677, n10197, n_15427);
  not g34124 (n_15428, n21672);
  and g34125 (n21678, n_15428, n21677);
  not g34126 (n_15429, n21678);
  and g34127 (n21679, n_7638, n_15429);
  not g34128 (n_15430, n21625);
  and g34129 (n21680, n_15412, n_15430);
  not g34130 (n_15431, n21628);
  and g34131 (n21681, pi0741, n_15431);
  not g34132 (n_15432, n21680);
  and g34133 (n21682, n_15414, n_15432);
  not g34134 (n_15433, n21681);
  and g34135 (n21683, n_15433, n21682);
  and g34136 (n21684, pi0724, n_15412);
  and g34137 (n21685, n21034, n21684);
  not g34138 (n_15434, n21683);
  not g34139 (n_15435, n21685);
  and g34140 (n21686, n_15434, n_15435);
  and g34141 (n21687, pi0156, n10197);
  not g34142 (n_15436, n21686);
  and g34143 (n21688, n_15436, n21687);
  not g34144 (n_15437, n21688);
  and g34145 (n21689, n_12415, n_15437);
  not g34146 (n_15438, n21679);
  and g34147 (n21690, n_15438, n21689);
  not g34148 (n_15439, n21668);
  not g34149 (n_15440, n21690);
  and g34150 (po0313, n_15439, n_15440);
  and g34151 (n21692, n_5686, n_12418);
  not g34152 (n_15442, pi0760);
  and g34153 (n21693, n_15442, pi0947);
  not g34154 (n_15444, pi0688);
  and g34155 (n21694, n_15444, n20902);
  not g34156 (n_15445, n21693);
  not g34157 (n_15446, n21694);
  and g34158 (n21695, n_15445, n_15446);
  not g34159 (n_15447, n21695);
  and g34160 (n21696, n2926, n_15447);
  not g34161 (n_15448, n21692);
  and g34162 (n21697, pi0832, n_15448);
  not g34163 (n_15449, n21696);
  and g34164 (n21698, n_15449, n21697);
  and g34165 (n21699, n_5686, n_14814);
  and g34166 (n21700, n16641, n_15445);
  and g34167 (n21701, pi0157, n_11740);
  not g34168 (n_15450, n21700);
  and g34169 (n21702, pi0038, n_15450);
  not g34170 (n_15451, n21701);
  and g34171 (n21703, n_15451, n21702);
  and g34172 (n21704, n_5686, pi0760);
  and g34173 (n21705, n_11736, n21704);
  and g34174 (n21706, n_5686, n_11719);
  not g34175 (n_15452, n21706);
  and g34176 (n21707, n21019, n_15452);
  and g34177 (n21708, n_5686, n_14891);
  and g34178 (n21709, n_9149, n_14911);
  not g34179 (n_15453, n21708);
  not g34180 (n_15454, n21709);
  and g34181 (n21710, n_15453, n_15454);
  not g34182 (n_15455, n21707);
  and g34183 (n21711, n_15442, n_15455);
  not g34184 (n_15456, n21710);
  and g34185 (n21712, n_15456, n21711);
  not g34186 (n_15457, n21705);
  and g34187 (n21713, pi0039, n_15457);
  not g34188 (n_15458, n21712);
  and g34189 (n21714, n_15458, n21713);
  and g34190 (n21715, n_5686, n_11674);
  and g34191 (n21716, n16958, n21693);
  not g34192 (n_15459, n21715);
  and g34193 (n21717, n_162, n_15459);
  not g34194 (n_15460, n21716);
  and g34195 (n21718, n_15460, n21717);
  not g34196 (n_15461, n21718);
  and g34197 (n21719, n_161, n_15461);
  not g34198 (n_15462, n21714);
  and g34199 (n21720, n_15462, n21719);
  not g34200 (n_15463, n21703);
  not g34201 (n_15464, n21720);
  and g34202 (n21721, n_15463, n_15464);
  not g34203 (n_15465, n21721);
  and g34204 (n21722, pi0688, n_15465);
  and g34205 (n21723, n_14975, n21718);
  and g34206 (n21724, n_15442, n21080);
  and g34207 (n21725, pi0760, n_14974);
  not g34208 (n_15466, n21724);
  and g34209 (n21726, pi0157, n_15466);
  not g34210 (n_15467, n21725);
  and g34211 (n21727, n_15467, n21726);
  and g34212 (n21728, pi0760, n_14961);
  and g34213 (n21729, n_15442, n21064);
  not g34214 (n_15468, n21728);
  and g34215 (n21730, n_5686, n_15468);
  not g34216 (n_15469, n21729);
  and g34217 (n21731, n_15469, n21730);
  not g34218 (n_15470, n21727);
  and g34219 (n21732, pi0039, n_15470);
  not g34220 (n_15471, n21731);
  and g34221 (n21733, n_15471, n21732);
  not g34222 (n_15472, n21723);
  not g34223 (n_15473, n21733);
  and g34224 (n21734, n_15472, n_15473);
  not g34225 (n_15474, n21734);
  and g34226 (n21735, n_161, n_15474);
  and g34227 (n21736, n_5686, n_11418);
  and g34228 (n21737, pi0760, pi0947);
  not g34229 (n_15475, n21737);
  and g34230 (n21738, n_162, n_15475);
  and g34231 (n21739, n21239, n21738);
  not g34232 (n_15476, n21736);
  and g34233 (n21740, pi0038, n_15476);
  not g34234 (n_15477, n21739);
  and g34235 (n21741, n_15477, n21740);
  not g34236 (n_15478, n21741);
  and g34237 (n21742, n_15444, n_15478);
  not g34238 (n_15479, n21735);
  and g34239 (n21743, n_15479, n21742);
  not g34240 (n_15480, n21722);
  not g34241 (n_15481, n21743);
  and g34242 (n21744, n_15480, n_15481);
  not g34243 (n_15482, n21744);
  and g34244 (n21745, n10197, n_15482);
  not g34245 (n_15483, n21699);
  and g34246 (n21746, n_12415, n_15483);
  not g34247 (n_15484, n21745);
  and g34248 (n21747, n_15484, n21746);
  not g34249 (n_15485, n21698);
  not g34250 (n_15486, n21747);
  and g34251 (po0314, n_15485, n_15486);
  and g34252 (n21749, n_6143, n_14814);
  and g34253 (n21750, pi0158, n_11740);
  not g34254 (n_15488, pi0753);
  and g34255 (n21751, n_15488, pi0947);
  not g34256 (n_15489, n21751);
  and g34257 (n21752, n16641, n_15489);
  not g34258 (n_15490, n21750);
  not g34259 (n_15491, n21752);
  and g34260 (n21753, n_15490, n_15491);
  not g34261 (n_15492, n21753);
  and g34262 (n21754, pi0038, n_15492);
  and g34263 (n21755, pi0158, n_11674);
  and g34264 (n21756, pi0753, n16958);
  not g34265 (n_15493, n21755);
  not g34266 (n_15494, n21756);
  and g34267 (n21757, n_15493, n_15494);
  and g34268 (n21758, n20989, n21757);
  and g34269 (n21759, n_6143, n21004);
  and g34270 (n21760, pi0158, n_14912);
  not g34271 (n_15495, n21760);
  and g34272 (n21761, n_15488, n_15495);
  not g34273 (n_15496, n21759);
  and g34274 (n21762, n_15496, n21761);
  and g34275 (n21763, n_6143, pi0753);
  and g34276 (n21764, n_11736, n21763);
  not g34277 (n_15497, n21762);
  not g34278 (n_15498, n21764);
  and g34279 (n21765, n_15497, n_15498);
  not g34280 (n_15499, n21765);
  and g34281 (n21766, pi0039, n_15499);
  not g34282 (n_15500, n21758);
  and g34283 (n21767, n_161, n_15500);
  not g34284 (n_15501, n21766);
  and g34285 (n21768, n_15501, n21767);
  not g34286 (n_15503, n21754);
  and g34287 (n21769, pi0702, n_15503);
  not g34288 (n_15504, n21768);
  and g34289 (n21770, n_15504, n21769);
  and g34290 (n21771, n_6143, n_11418);
  and g34291 (n21772, pi0753, pi0947);
  not g34292 (n_15505, n21772);
  and g34293 (n21773, n_162, n_15505);
  and g34294 (n21774, n21239, n21773);
  not g34295 (n_15506, n21771);
  and g34296 (n21775, pi0038, n_15506);
  not g34297 (n_15507, n21774);
  and g34298 (n21776, n_15507, n21775);
  and g34299 (n21777, n21097, n_15489);
  and g34300 (n21778, n_162, n_15493);
  not g34301 (n_15508, n21777);
  and g34302 (n21779, n_15508, n21778);
  and g34303 (n21780, n_6143, n_14961);
  and g34304 (n21781, pi0158, n_14974);
  not g34305 (n_15509, n21781);
  and g34306 (n21782, pi0753, n_15509);
  not g34307 (n_15510, n21780);
  and g34308 (n21783, n_15510, n21782);
  and g34309 (n21784, n_6143, n21064);
  and g34310 (n21785, pi0158, n21080);
  not g34311 (n_15511, n21785);
  and g34312 (n21786, n_15488, n_15511);
  not g34313 (n_15512, n21784);
  and g34314 (n21787, n_15512, n21786);
  not g34315 (n_15513, n21783);
  not g34316 (n_15514, n21787);
  and g34317 (n21788, n_15513, n_15514);
  not g34318 (n_15515, n21788);
  and g34319 (n21789, pi0039, n_15515);
  not g34320 (n_15516, n21779);
  and g34321 (n21790, n_161, n_15516);
  not g34322 (n_15517, n21789);
  and g34323 (n21791, n_15517, n21790);
  not g34324 (n_15518, pi0702);
  not g34325 (n_15519, n21776);
  and g34326 (n21792, n_15518, n_15519);
  not g34327 (n_15520, n21791);
  and g34328 (n21793, n_15520, n21792);
  not g34329 (n_15521, n21770);
  not g34330 (n_15522, n21793);
  and g34331 (n21794, n_15521, n_15522);
  not g34332 (n_15523, n21794);
  and g34333 (n21795, n10197, n_15523);
  not g34334 (n_15524, n21749);
  and g34335 (n21796, n_12415, n_15524);
  not g34336 (n_15525, n21795);
  and g34337 (n21797, n_15525, n21796);
  and g34338 (n21798, n_6143, n_12418);
  and g34339 (n21799, n_15518, n20902);
  not g34340 (n_15526, n21799);
  and g34341 (n21800, n_15489, n_15526);
  not g34342 (n_15527, n21800);
  and g34343 (n21801, n2926, n_15527);
  not g34344 (n_15528, n21798);
  and g34345 (n21802, pi0832, n_15528);
  not g34346 (n_15529, n21801);
  and g34347 (n21803, n_15529, n21802);
  not g34348 (n_15530, n21797);
  not g34349 (n_15531, n21803);
  and g34350 (po0315, n_15530, n_15531);
  and g34351 (n21805, n_6307, n_14814);
  and g34352 (n21806, pi0159, n_11740);
  not g34353 (n_15533, pi0754);
  and g34354 (n21807, n_15533, pi0947);
  not g34355 (n_15534, n21807);
  and g34356 (n21808, n16641, n_15534);
  not g34357 (n_15535, n21806);
  not g34358 (n_15536, n21808);
  and g34359 (n21809, n_15535, n_15536);
  not g34360 (n_15537, n21809);
  and g34361 (n21810, pi0038, n_15537);
  and g34362 (n21811, pi0159, n_11674);
  and g34363 (n21812, pi0754, n16958);
  not g34364 (n_15538, n21811);
  not g34365 (n_15539, n21812);
  and g34366 (n21813, n_15538, n_15539);
  and g34367 (n21814, n20989, n21813);
  and g34368 (n21815, n_6307, n21004);
  and g34369 (n21816, pi0159, n_14912);
  not g34370 (n_15540, n21816);
  and g34371 (n21817, n_15533, n_15540);
  not g34372 (n_15541, n21815);
  and g34373 (n21818, n_15541, n21817);
  and g34374 (n21819, n_6307, pi0754);
  and g34375 (n21820, n_11736, n21819);
  not g34376 (n_15542, n21818);
  not g34377 (n_15543, n21820);
  and g34378 (n21821, n_15542, n_15543);
  not g34379 (n_15544, n21821);
  and g34380 (n21822, pi0039, n_15544);
  not g34381 (n_15545, n21814);
  and g34382 (n21823, n_161, n_15545);
  not g34383 (n_15546, n21822);
  and g34384 (n21824, n_15546, n21823);
  not g34385 (n_15548, n21810);
  and g34386 (n21825, pi0709, n_15548);
  not g34387 (n_15549, n21824);
  and g34388 (n21826, n_15549, n21825);
  and g34389 (n21827, n_6307, n_11418);
  and g34390 (n21828, pi0754, pi0947);
  not g34391 (n_15550, n21828);
  and g34392 (n21829, n_162, n_15550);
  and g34393 (n21830, n21239, n21829);
  not g34394 (n_15551, n21827);
  and g34395 (n21831, pi0038, n_15551);
  not g34396 (n_15552, n21830);
  and g34397 (n21832, n_15552, n21831);
  and g34398 (n21833, n21097, n_15534);
  and g34399 (n21834, n_162, n_15538);
  not g34400 (n_15553, n21833);
  and g34401 (n21835, n_15553, n21834);
  and g34402 (n21836, n_6307, n_14961);
  and g34403 (n21837, pi0159, n_14974);
  not g34404 (n_15554, n21837);
  and g34405 (n21838, pi0754, n_15554);
  not g34406 (n_15555, n21836);
  and g34407 (n21839, n_15555, n21838);
  and g34408 (n21840, n_6307, n21064);
  and g34409 (n21841, pi0159, n21080);
  not g34410 (n_15556, n21841);
  and g34411 (n21842, n_15533, n_15556);
  not g34412 (n_15557, n21840);
  and g34413 (n21843, n_15557, n21842);
  not g34414 (n_15558, n21839);
  not g34415 (n_15559, n21843);
  and g34416 (n21844, n_15558, n_15559);
  not g34417 (n_15560, n21844);
  and g34418 (n21845, pi0039, n_15560);
  not g34419 (n_15561, n21835);
  and g34420 (n21846, n_161, n_15561);
  not g34421 (n_15562, n21845);
  and g34422 (n21847, n_15562, n21846);
  not g34423 (n_15563, pi0709);
  not g34424 (n_15564, n21832);
  and g34425 (n21848, n_15563, n_15564);
  not g34426 (n_15565, n21847);
  and g34427 (n21849, n_15565, n21848);
  not g34428 (n_15566, n21826);
  not g34429 (n_15567, n21849);
  and g34430 (n21850, n_15566, n_15567);
  not g34431 (n_15568, n21850);
  and g34432 (n21851, n10197, n_15568);
  not g34433 (n_15569, n21805);
  and g34434 (n21852, n_12415, n_15569);
  not g34435 (n_15570, n21851);
  and g34436 (n21853, n_15570, n21852);
  and g34437 (n21854, n_6307, n_12418);
  and g34438 (n21855, n_15563, n20902);
  not g34439 (n_15571, n21855);
  and g34440 (n21856, n_15534, n_15571);
  not g34441 (n_15572, n21856);
  and g34442 (n21857, n2926, n_15572);
  not g34443 (n_15573, n21854);
  and g34444 (n21858, pi0832, n_15573);
  not g34445 (n_15574, n21857);
  and g34446 (n21859, n_15574, n21858);
  not g34447 (n_15575, n21853);
  not g34448 (n_15576, n21859);
  and g34449 (po0316, n_15575, n_15576);
  and g34450 (n21861, n_7697, n_12418);
  not g34451 (n_15578, pi0756);
  and g34452 (n21862, n_15578, pi0947);
  not g34453 (n_15580, pi0734);
  and g34454 (n21863, n_15580, n20902);
  not g34455 (n_15581, n21862);
  not g34456 (n_15582, n21863);
  and g34457 (n21864, n_15581, n_15582);
  not g34458 (n_15583, n21864);
  and g34459 (n21865, n2926, n_15583);
  not g34460 (n_15584, n21861);
  and g34461 (n21866, pi0832, n_15584);
  not g34462 (n_15585, n21865);
  and g34463 (n21867, n_15585, n21866);
  and g34464 (n21868, n_7697, n_14814);
  and g34465 (n21869, n16641, n_15581);
  and g34466 (n21870, pi0160, n_11740);
  not g34467 (n_15586, n21869);
  and g34468 (n21871, pi0038, n_15586);
  not g34469 (n_15587, n21870);
  and g34470 (n21872, n_15587, n21871);
  and g34471 (n21873, n_7697, n_11674);
  and g34472 (n21874, n16958, n21862);
  not g34473 (n_15588, n21873);
  and g34474 (n21875, n_162, n_15588);
  not g34475 (n_15589, n21874);
  and g34476 (n21876, n_15589, n21875);
  and g34477 (n21877, n_7697, n_14891);
  and g34478 (n21878, pi0160, n_15009);
  not g34479 (n_15590, n21878);
  and g34480 (n21879, pi0299, n_15590);
  not g34481 (n_15591, n21877);
  and g34482 (n21880, n_15591, n21879);
  and g34483 (n21881, n_7697, n_11719);
  not g34484 (n_15592, n21881);
  and g34485 (n21882, n21019, n_15592);
  not g34486 (n_15593, n21882);
  and g34487 (n21883, n_15578, n_15593);
  not g34488 (n_15594, n21880);
  and g34489 (n21884, n_15594, n21883);
  and g34490 (n21885, n_7697, pi0756);
  and g34491 (n21886, n_11736, n21885);
  not g34492 (n_15595, n21886);
  and g34493 (n21887, pi0039, n_15595);
  not g34494 (n_15596, n21884);
  and g34495 (n21888, n_15596, n21887);
  not g34496 (n_15597, n21876);
  and g34497 (n21889, n_161, n_15597);
  not g34498 (n_15598, n21888);
  and g34499 (n21890, n_15598, n21889);
  not g34500 (n_15599, n21872);
  not g34501 (n_15600, n21890);
  and g34502 (n21891, n_15599, n_15600);
  not g34503 (n_15601, n21891);
  and g34504 (n21892, pi0734, n_15601);
  and g34505 (n21893, n_14975, n21876);
  and g34506 (n21894, n_7697, n21064);
  and g34507 (n21895, pi0160, n21080);
  not g34508 (n_15602, n21895);
  and g34509 (n21896, n_15578, n_15602);
  not g34510 (n_15603, n21894);
  and g34511 (n21897, n_15603, n21896);
  and g34512 (n21898, pi0160, n_14995);
  and g34513 (n21899, n_7697, n21093);
  not g34519 (n_15606, n21902);
  and g34520 (n21903, pi0039, n_15606);
  not g34521 (n_15607, n21897);
  and g34522 (n21904, n_15607, n21903);
  not g34523 (n_15608, n21893);
  not g34524 (n_15609, n21904);
  and g34525 (n21905, n_15608, n_15609);
  not g34526 (n_15610, n21905);
  and g34527 (n21906, n_161, n_15610);
  and g34528 (n21907, n_7697, n_11418);
  and g34529 (n21908, pi0756, pi0947);
  not g34530 (n_15611, n21908);
  and g34531 (n21909, n_162, n_15611);
  and g34532 (n21910, n21239, n21909);
  not g34533 (n_15612, n21907);
  and g34534 (n21911, pi0038, n_15612);
  not g34535 (n_15613, n21910);
  and g34536 (n21912, n_15613, n21911);
  not g34537 (n_15614, n21912);
  and g34538 (n21913, n_15580, n_15614);
  not g34539 (n_15615, n21906);
  and g34540 (n21914, n_15615, n21913);
  not g34541 (n_15616, n21892);
  not g34542 (n_15617, n21914);
  and g34543 (n21915, n_15616, n_15617);
  not g34544 (n_15618, n21915);
  and g34545 (n21916, n10197, n_15618);
  not g34546 (n_15619, n21868);
  and g34547 (n21917, n_12415, n_15619);
  not g34548 (n_15620, n21916);
  and g34549 (n21918, n_15620, n21917);
  not g34550 (n_15621, n21867);
  not g34551 (n_15622, n21918);
  and g34552 (po0317, n_15621, n_15622);
  and g34553 (n21920, n_264, n_14814);
  and g34554 (n21921, n_264, n_11418);
  and g34555 (n21922, pi0758, pi0947);
  not g34556 (n_15623, n21922);
  and g34557 (n21923, n_162, n_15623);
  and g34558 (n21924, n21390, n21923);
  not g34559 (n_15624, n21921);
  and g34560 (n21925, pi0038, n_15624);
  not g34561 (n_15625, n21924);
  and g34562 (n21926, n_15625, n21925);
  and g34563 (n21927, n16958, n21922);
  and g34564 (n21928, pi0161, n_11674);
  not g34565 (n_15626, n21927);
  and g34566 (n21929, n_162, n_15626);
  not g34567 (n_15627, n21928);
  and g34568 (n21930, n_15627, n21929);
  and g34569 (n21931, n_14975, n21930);
  and g34570 (n21932, n_264, n_11729);
  not g34571 (n_15628, n21932);
  and g34572 (n21933, n20998, n_15628);
  and g34573 (n21934, n_15198, n21933);
  and g34574 (n21935, pi0161, n21046);
  not g34575 (n_15629, n21935);
  and g34576 (n21936, n21102, n_15629);
  and g34577 (n21937, pi0161, n_11445);
  not g34578 (n_15630, n21937);
  and g34579 (n21938, n_15143, n_15630);
  and g34580 (n21939, n3448, n21938);
  not g34581 (n_15631, n21939);
  and g34582 (n21940, n_36, n_15631);
  and g34583 (n21941, n_14926, n21940);
  not g34584 (n_15632, n21936);
  and g34585 (n21942, n_15632, n21941);
  not g34586 (n_15633, n21934);
  and g34587 (n21943, pi0299, n_15633);
  not g34588 (n_15634, n21942);
  and g34589 (n21944, n_15634, n21943);
  and g34590 (n21945, n_14964, n_15630);
  not g34591 (n_15635, n21945);
  and g34592 (n21946, n2603, n_15635);
  and g34593 (n21947, n_264, n_15206);
  not g34594 (n_15636, n21947);
  and g34595 (n21948, n21416, n_15636);
  not g34596 (n_15637, n21946);
  not g34597 (n_15638, n21948);
  and g34598 (n21949, n_15637, n_15638);
  not g34599 (n_15639, n21949);
  and g34600 (n21950, n_223, n_15639);
  and g34601 (n21951, n_264, n_11697);
  not g34602 (n_15640, n21951);
  and g34603 (n21952, n21055, n_15640);
  not g34604 (n_15641, n21952);
  and g34605 (n21953, n_234, n_15641);
  not g34606 (n_15642, n21950);
  and g34607 (n21954, n_15642, n21953);
  not g34608 (n_15643, n21944);
  and g34609 (n21955, n_14083, n_15643);
  not g34610 (n_15644, n21954);
  and g34611 (n21956, n_15644, n21955);
  and g34612 (n21957, n_15140, n21936);
  not g34613 (n_15645, n21957);
  and g34614 (n21958, n21940, n_15645);
  not g34615 (n_15646, n21933);
  and g34616 (n21959, pi0299, n_15646);
  not g34617 (n_15647, n21958);
  and g34618 (n21960, n_15647, n21959);
  and g34619 (n21961, n2603, n21938);
  and g34620 (n21962, n21432, n_15636);
  not g34621 (n_15648, n21962);
  and g34622 (n21963, n21435, n_15648);
  not g34623 (n_15649, n21961);
  and g34624 (n21964, n_223, n_15649);
  not g34625 (n_15650, n21963);
  and g34626 (n21965, n_15650, n21964);
  and g34627 (n21966, n21053, n_15640);
  not g34628 (n_15651, n21966);
  and g34629 (n21967, n_234, n_15651);
  and g34630 (n21968, n_15641, n21967);
  not g34631 (n_15652, n21965);
  and g34632 (n21969, n_15652, n21968);
  not g34633 (n_15653, n21960);
  and g34634 (n21970, pi0758, n_15653);
  not g34635 (n_15654, n21969);
  and g34636 (n21971, n_15654, n21970);
  not g34637 (n_15655, n21956);
  and g34638 (n21972, pi0039, n_15655);
  not g34639 (n_15656, n21971);
  and g34640 (n21973, n_15656, n21972);
  not g34641 (n_15657, n21931);
  and g34642 (n21974, n_161, n_15657);
  not g34643 (n_15658, n21973);
  and g34644 (n21975, n_15658, n21974);
  not g34645 (n_15659, n21926);
  and g34646 (n21976, pi0736, n_15659);
  not g34647 (n_15660, n21975);
  and g34648 (n21977, n_15660, n21976);
  and g34649 (n21978, n_264, n_11740);
  and g34650 (n21979, n16641, n_15623);
  not g34651 (n_15661, n21979);
  and g34652 (n21980, pi0038, n_15661);
  not g34653 (n_15662, n21978);
  and g34654 (n21981, n_15662, n21980);
  and g34655 (n21982, n_14906, n_15630);
  not g34656 (n_15663, n21982);
  and g34657 (n21983, n2603, n_15663);
  not g34658 (n_15664, n21983);
  and g34659 (n21984, n_15648, n_15664);
  not g34660 (n_15665, n21984);
  and g34661 (n21985, n_223, n_15665);
  not g34662 (n_15666, n21985);
  and g34663 (n21986, n21967, n_15666);
  and g34664 (n21987, pi0161, n21000);
  and g34665 (n21988, n3448, n21982);
  and g34666 (n21989, n_14886, n_15632);
  not g34667 (n_15667, n21989);
  and g34668 (n21990, n_14905, n_15667);
  not g34669 (n_15668, n21988);
  and g34670 (n21991, n_36, n_15668);
  not g34671 (n_15669, n21990);
  and g34672 (n21992, n_15669, n21991);
  not g34673 (n_15670, n21987);
  and g34674 (n21993, n21022, n_15670);
  not g34675 (n_15671, n21992);
  and g34676 (n21994, n_15671, n21993);
  not g34677 (n_15672, n21986);
  and g34678 (n21995, pi0758, n_15672);
  not g34679 (n_15673, n21994);
  and g34680 (n21996, n_15673, n21995);
  and g34681 (n21997, pi0161, n19958);
  not g34682 (n_15674, n21997);
  and g34683 (n21998, pi0039, n_15674);
  not g34684 (n_15675, n21996);
  and g34685 (n21999, n_15675, n21998);
  not g34686 (n_15676, n21930);
  and g34687 (n22000, n_161, n_15676);
  not g34688 (n_15677, n21999);
  and g34689 (n22001, n_15677, n22000);
  not g34690 (n_15678, n21981);
  and g34691 (n22002, n_14126, n_15678);
  not g34692 (n_15679, n22001);
  and g34693 (n22003, n_15679, n22002);
  not g34694 (n_15680, n21977);
  not g34695 (n_15681, n22003);
  and g34696 (n22004, n_15680, n_15681);
  not g34697 (n_15682, n22004);
  and g34698 (n22005, n10197, n_15682);
  not g34699 (n_15683, n21920);
  and g34700 (n22006, n_12415, n_15683);
  not g34701 (n_15684, n22005);
  and g34702 (n22007, n_15684, n22006);
  and g34703 (n22008, n_264, n_12418);
  and g34704 (n22009, pi0736, n20902);
  and g34705 (n22010, n2926, n_15623);
  not g34706 (n_15685, n22009);
  and g34707 (n22011, n_15685, n22010);
  not g34708 (n_15686, n22008);
  and g34709 (n22012, pi0832, n_15686);
  not g34710 (n_15687, n22011);
  and g34711 (n22013, n_15687, n22012);
  or g34712 (po0318, n22007, n22013);
  and g34713 (n22015, n_6224, n_14814);
  and g34714 (n22016, n_11912, pi0947);
  not g34715 (n_15688, n22016);
  and g34716 (n22017, n16641, n_15688);
  and g34717 (n22018, pi0162, n_11740);
  not g34718 (n_15689, n22017);
  and g34719 (n22019, pi0038, n_15689);
  not g34720 (n_15690, n22018);
  and g34721 (n22020, n_15690, n22019);
  and g34722 (n22021, n_6224, n_11674);
  and g34723 (n22022, n16958, n22016);
  not g34724 (n_15691, n22021);
  and g34725 (n22023, n_162, n_15691);
  not g34726 (n_15692, n22022);
  and g34727 (n22024, n_15692, n22023);
  and g34728 (n22025, n14933, n_15009);
  not g34729 (n_15693, n22025);
  and g34730 (n22026, n_14893, n_15693);
  not g34731 (n_15694, n22026);
  and g34732 (n22027, n_11912, n_15694);
  and g34733 (n22028, n_11912, n21003);
  and g34734 (n22029, pi0761, n17046);
  not g34735 (n_15695, n22029);
  and g34736 (n22030, n_6224, n_15695);
  not g34737 (n_15696, n22028);
  and g34738 (n22031, n_15696, n22030);
  not g34739 (n_15697, n22027);
  and g34740 (n22032, pi0039, n_15697);
  not g34741 (n_15698, n22031);
  and g34742 (n22033, n_15698, n22032);
  not g34743 (n_15699, n22024);
  and g34744 (n22034, n_161, n_15699);
  not g34745 (n_15700, n22033);
  and g34746 (n22035, n_15700, n22034);
  not g34747 (n_15701, n22020);
  not g34748 (n_15702, n22035);
  and g34749 (n22036, n_15701, n_15702);
  not g34750 (n_15703, n22036);
  and g34751 (n22037, pi0738, n_15703);
  and g34752 (n22038, n_14975, n22024);
  and g34753 (n22039, pi0162, n_14995);
  and g34754 (n22040, n_10086, n_14961);
  not g34755 (n_15704, n22039);
  and g34756 (n22041, pi0761, n_15704);
  not g34757 (n_15705, n22040);
  and g34758 (n22042, n_15705, n22041);
  and g34759 (n22043, n_6224, n21064);
  and g34760 (n22044, pi0162, n21080);
  not g34761 (n_15706, n22044);
  and g34762 (n22045, n_11912, n_15706);
  not g34763 (n_15707, n22043);
  and g34764 (n22046, n_15707, n22045);
  not g34765 (n_15708, n22042);
  and g34766 (n22047, pi0039, n_15708);
  not g34767 (n_15709, n22046);
  and g34768 (n22048, n_15709, n22047);
  not g34769 (n_15710, n22038);
  not g34770 (n_15711, n22048);
  and g34771 (n22049, n_15710, n_15711);
  not g34772 (n_15712, n22049);
  and g34773 (n22050, n_161, n_15712);
  and g34774 (n22051, n_6224, n_11418);
  and g34775 (n22052, pi0761, pi0947);
  not g34776 (n_15713, n22052);
  and g34777 (n22053, n_162, n_15713);
  and g34778 (n22054, n21239, n22053);
  not g34779 (n_15714, n22051);
  and g34780 (n22055, pi0038, n_15714);
  not g34781 (n_15715, n22054);
  and g34782 (n22056, n_15715, n22055);
  not g34783 (n_15716, n22056);
  and g34784 (n22057, n_11667, n_15716);
  not g34785 (n_15717, n22050);
  and g34786 (n22058, n_15717, n22057);
  not g34787 (n_15718, n22037);
  not g34788 (n_15719, n22058);
  and g34789 (n22059, n_15718, n_15719);
  not g34790 (n_15720, n22059);
  and g34791 (n22060, n10197, n_15720);
  not g34792 (n_15721, n22015);
  and g34793 (n22061, n_12415, n_15721);
  not g34794 (n_15722, n22060);
  and g34795 (n22062, n_15722, n22061);
  and g34796 (n22063, n_6224, n_12418);
  and g34797 (n22064, n_11667, n20902);
  not g34798 (n_15723, n22064);
  and g34799 (n22065, n_15688, n_15723);
  not g34800 (n_15724, n22065);
  and g34801 (n22066, n2926, n_15724);
  not g34802 (n_15725, n22063);
  and g34803 (n22067, pi0832, n_15725);
  not g34804 (n_15726, n22066);
  and g34805 (n22068, n_15726, n22067);
  not g34806 (n_15727, n22062);
  not g34807 (n_15728, n22068);
  and g34808 (po0319, n_15727, n_15728);
  and g34809 (n22070, n_7591, n_12418);
  not g34810 (n_15730, pi0777);
  and g34811 (n22071, n_15730, pi0947);
  not g34812 (n_15732, pi0737);
  and g34813 (n22072, n_15732, n20902);
  not g34814 (n_15733, n22071);
  not g34815 (n_15734, n22072);
  and g34816 (n22073, n_15733, n_15734);
  not g34817 (n_15735, n22073);
  and g34818 (n22074, n2926, n_15735);
  not g34819 (n_15736, n22070);
  and g34820 (n22075, pi0832, n_15736);
  not g34821 (n_15737, n22074);
  and g34822 (n22076, n_15737, n22075);
  and g34823 (n22077, n_7591, n_14814);
  and g34824 (n22078, n16641, n_15733);
  and g34825 (n22079, pi0163, n_11740);
  not g34826 (n_15738, n22078);
  and g34827 (n22080, pi0038, n_15738);
  not g34828 (n_15739, n22079);
  and g34829 (n22081, n_15739, n22080);
  and g34830 (n22082, n_7591, n_11674);
  and g34831 (n22083, n16958, n22071);
  not g34832 (n_15740, n22082);
  and g34833 (n22084, n_162, n_15740);
  not g34834 (n_15741, n22083);
  and g34835 (n22085, n_15741, n22084);
  and g34836 (n22086, n_7591, n_11719);
  not g34837 (n_15742, n22086);
  and g34838 (n22087, n21019, n_15742);
  and g34839 (n22088, n_7591, n_14891);
  and g34840 (n22089, n_9943, n_14911);
  not g34841 (n_15743, n22088);
  not g34842 (n_15744, n22089);
  and g34843 (n22090, n_15743, n_15744);
  not g34844 (n_15745, n22087);
  and g34845 (n22091, n_15730, n_15745);
  not g34846 (n_15746, n22090);
  and g34847 (n22092, n_15746, n22091);
  and g34848 (n22093, n_7591, pi0777);
  and g34849 (n22094, n_11736, n22093);
  not g34850 (n_15747, n22094);
  and g34851 (n22095, pi0039, n_15747);
  not g34852 (n_15748, n22092);
  and g34853 (n22096, n_15748, n22095);
  not g34854 (n_15749, n22085);
  and g34855 (n22097, n_161, n_15749);
  not g34856 (n_15750, n22096);
  and g34857 (n22098, n_15750, n22097);
  not g34858 (n_15751, n22081);
  not g34859 (n_15752, n22098);
  and g34860 (n22099, n_15751, n_15752);
  not g34861 (n_15753, n22099);
  and g34862 (n22100, pi0737, n_15753);
  and g34863 (n22101, n_14975, n22085);
  and g34864 (n22102, n_7591, n21064);
  and g34865 (n22103, pi0163, n21080);
  not g34866 (n_15754, n22103);
  and g34867 (n22104, n_15730, n_15754);
  not g34868 (n_15755, n22102);
  and g34869 (n22105, n_15755, n22104);
  and g34870 (n22106, n_7591, n21093);
  and g34871 (n22107, pi0163, n_14995);
  not g34877 (n_15758, n22110);
  and g34878 (n22111, pi0039, n_15758);
  not g34879 (n_15759, n22105);
  and g34880 (n22112, n_15759, n22111);
  not g34881 (n_15760, n22101);
  not g34882 (n_15761, n22112);
  and g34883 (n22113, n_15760, n_15761);
  not g34884 (n_15762, n22113);
  and g34885 (n22114, n_161, n_15762);
  and g34886 (n22115, n_7591, n_11418);
  and g34887 (n22116, pi0777, pi0947);
  not g34888 (n_15763, n22116);
  and g34889 (n22117, n_162, n_15763);
  and g34890 (n22118, n21239, n22117);
  not g34891 (n_15764, n22115);
  and g34892 (n22119, pi0038, n_15764);
  not g34893 (n_15765, n22118);
  and g34894 (n22120, n_15765, n22119);
  not g34895 (n_15766, n22120);
  and g34896 (n22121, n_15732, n_15766);
  not g34897 (n_15767, n22114);
  and g34898 (n22122, n_15767, n22121);
  not g34899 (n_15768, n22100);
  not g34900 (n_15769, n22122);
  and g34901 (n22123, n_15768, n_15769);
  not g34902 (n_15770, n22123);
  and g34903 (n22124, n10197, n_15770);
  not g34904 (n_15771, n22077);
  and g34905 (n22125, n_12415, n_15771);
  not g34906 (n_15772, n22124);
  and g34907 (n22126, n_15772, n22125);
  not g34908 (n_15773, n22076);
  not g34909 (n_15774, n22126);
  and g34910 (po0320, n_15773, n_15774);
  and g34911 (n22128, n_5727, n_12418);
  not g34912 (n_15776, pi0752);
  and g34913 (n22129, n_15776, pi0947);
  and g34914 (n22130, pi0703, n20902);
  not g34915 (n_15778, n22129);
  not g34916 (n_15779, n22130);
  and g34917 (n22131, n_15778, n_15779);
  not g34918 (n_15780, n22131);
  and g34919 (n22132, n2926, n_15780);
  not g34920 (n_15781, n22128);
  and g34921 (n22133, pi0832, n_15781);
  not g34922 (n_15782, n22132);
  and g34923 (n22134, n_15782, n22133);
  and g34924 (n22135, n_5727, n_14814);
  and g34925 (n22136, n_5727, n_14920);
  not g34926 (n_15783, n22136);
  and g34927 (n22137, n21042, n_15783);
  and g34928 (n22138, n_5727, n21069);
  and g34929 (n22139, pi0164, n21082);
  not g34930 (n_15784, n22139);
  and g34931 (n22140, n_161, n_15784);
  not g34932 (n_15785, n22138);
  and g34933 (n22141, n_15785, n22140);
  not g34934 (n_15786, n22137);
  and g34935 (n22142, n_15776, n_15786);
  not g34936 (n_15787, n22141);
  and g34937 (n22143, n_15787, n22142);
  and g34938 (n22144, n_5727, n_11418);
  not g34939 (n_15788, n22144);
  and g34940 (n22145, n21090, n_15788);
  and g34941 (n22146, n_5727, n21099);
  and g34942 (n22147, pi0164, n21116);
  not g34943 (n_15789, n22147);
  and g34944 (n22148, n_161, n_15789);
  not g34945 (n_15790, n22146);
  and g34946 (n22149, n_15790, n22148);
  not g34947 (n_15791, n22145);
  and g34948 (n22150, pi0752, n_15791);
  not g34949 (n_15792, n22149);
  and g34950 (n22151, n_15792, n22150);
  not g34951 (n_15793, n22143);
  not g34952 (n_15794, n22151);
  and g34953 (n22152, n_15793, n_15794);
  not g34954 (n_15795, n22152);
  and g34955 (n22153, pi0703, n_15795);
  and g34956 (n22154, pi0752, n17052);
  and g34957 (n22155, n_15776, n21034);
  not g34958 (n_15796, n22155);
  and g34959 (n22156, pi0164, n_15796);
  and g34960 (n22157, pi0164, n_14898);
  not g34961 (n_15797, n22157);
  and g34962 (n22158, n_15776, n_15797);
  and g34963 (n22159, n_15424, n22158);
  not g34964 (n_15798, pi0703);
  not g34971 (n_15802, n22153);
  not g34972 (n_15803, n22162);
  and g34973 (n22163, n_15802, n_15803);
  not g34974 (n_15804, n22163);
  and g34975 (n22164, n10197, n_15804);
  not g34976 (n_15805, n22135);
  and g34977 (n22165, n_12415, n_15805);
  not g34978 (n_15806, n22164);
  and g34979 (n22166, n_15806, n22165);
  not g34980 (n_15807, n22134);
  not g34981 (n_15808, n22166);
  and g34982 (po0321, n_15807, n_15808);
  and g34983 (n22168, n_9142, n_12418);
  and g34984 (n22169, n_13676, pi0947);
  and g34985 (n22170, pi0687, n20902);
  not g34986 (n_15809, n22169);
  not g34987 (n_15810, n22170);
  and g34988 (n22171, n_15809, n_15810);
  not g34989 (n_15811, n22171);
  and g34990 (n22172, n2926, n_15811);
  not g34991 (n_15812, n22168);
  and g34992 (n22173, pi0832, n_15812);
  not g34993 (n_15813, n22172);
  and g34994 (n22174, n_15813, n22173);
  and g34995 (n22175, n_9142, n_14814);
  and g34996 (n22176, n_9142, n_14920);
  not g34997 (n_15814, n22176);
  and g34998 (n22177, n21042, n_15814);
  and g34999 (n22178, n_9142, n21069);
  and g35000 (n22179, pi0165, n21082);
  not g35001 (n_15815, n22179);
  and g35002 (n22180, n_161, n_15815);
  not g35003 (n_15816, n22178);
  and g35004 (n22181, n_15816, n22180);
  not g35005 (n_15817, n22177);
  and g35006 (n22182, n_13676, n_15817);
  not g35007 (n_15818, n22181);
  and g35008 (n22183, n_15818, n22182);
  and g35009 (n22184, n_9142, n_11418);
  not g35010 (n_15819, n22184);
  and g35011 (n22185, n21090, n_15819);
  and g35012 (n22186, n_9142, n21099);
  and g35013 (n22187, pi0165, n21116);
  not g35014 (n_15820, n22187);
  and g35015 (n22188, n_161, n_15820);
  not g35016 (n_15821, n22186);
  and g35017 (n22189, n_15821, n22188);
  not g35018 (n_15822, n22185);
  and g35019 (n22190, pi0774, n_15822);
  not g35020 (n_15823, n22189);
  and g35021 (n22191, n_15823, n22190);
  not g35022 (n_15824, n22183);
  not g35023 (n_15825, n22191);
  and g35024 (n22192, n_15824, n_15825);
  not g35025 (n_15826, n22192);
  and g35026 (n22193, pi0687, n_15826);
  and g35027 (n22194, pi0774, n17052);
  and g35028 (n22195, n_13676, n21034);
  not g35029 (n_15827, n22195);
  and g35030 (n22196, pi0165, n_15827);
  and g35031 (n22197, pi0165, n_14898);
  not g35032 (n_15828, n22197);
  and g35033 (n22198, n_13676, n_15828);
  and g35034 (n22199, n_15424, n22198);
  not g35041 (n_15832, n22193);
  not g35042 (n_15833, n22202);
  and g35043 (n22203, n_15832, n_15833);
  not g35044 (n_15834, n22203);
  and g35045 (n22204, n10197, n_15834);
  not g35046 (n_15835, n22175);
  and g35047 (n22205, n_12415, n_15835);
  not g35048 (n_15836, n22204);
  and g35049 (n22206, n_15836, n22205);
  not g35050 (n_15837, n22174);
  not g35051 (n_15838, n22206);
  and g35052 (po0322, n_15837, n_15838);
  and g35053 (n22208, n_266, n_14814);
  and g35054 (n22209, n_266, n_11740);
  and g35055 (n22210, pi0772, pi0947);
  not g35056 (n_15840, n22210);
  and g35057 (n22211, n16641, n_15840);
  not g35058 (n_15841, n22211);
  and g35059 (n22212, pi0038, n_15841);
  not g35060 (n_15842, n22209);
  and g35061 (n22213, n_15842, n22212);
  and g35062 (n22214, pi0166, n_11674);
  and g35063 (n22215, n_162, n_15840);
  not g35064 (n_15843, n22215);
  and g35065 (n22216, n_11737, n_15843);
  not g35066 (n_15844, n22214);
  not g35067 (n_15845, n22216);
  and g35068 (n22217, n_15844, n_15845);
  and g35069 (n22218, n_266, n_11697);
  not g35070 (n_15846, n22218);
  and g35071 (n22219, n21053, n_15846);
  not g35072 (n_15847, n22219);
  and g35073 (n22220, n_234, n_15847);
  and g35074 (n22221, pi0166, n_11445);
  not g35075 (n_15848, n22221);
  and g35076 (n22222, n_14906, n_15848);
  not g35077 (n_15849, n22222);
  and g35078 (n22223, n2603, n_15849);
  and g35079 (n22224, n_266, n_15206);
  not g35080 (n_15850, n22224);
  and g35081 (n22225, n21432, n_15850);
  not g35082 (n_15851, n22223);
  not g35083 (n_15852, n22225);
  and g35084 (n22226, n_15851, n_15852);
  not g35085 (n_15853, n22226);
  and g35086 (n22227, n_223, n_15853);
  not g35087 (n_15854, n22227);
  and g35088 (n22228, n22220, n_15854);
  and g35089 (n22229, pi0166, n21000);
  and g35090 (n22230, n3448, n22222);
  and g35091 (n22231, pi0166, n21046);
  not g35092 (n_15855, n22231);
  and g35093 (n22232, n21102, n_15855);
  not g35094 (n_15856, n22232);
  and g35095 (n22233, n_14886, n_15856);
  not g35096 (n_15857, n22233);
  and g35097 (n22234, n_14905, n_15857);
  not g35098 (n_15858, n22230);
  and g35099 (n22235, n_36, n_15858);
  not g35100 (n_15859, n22234);
  and g35101 (n22236, n_15859, n22235);
  not g35102 (n_15860, n22229);
  and g35103 (n22237, n21022, n_15860);
  not g35104 (n_15861, n22236);
  and g35105 (n22238, n_15861, n22237);
  not g35106 (n_15862, n22228);
  and g35107 (n22239, pi0772, n_15862);
  not g35108 (n_15863, n22238);
  and g35109 (n22240, n_15863, n22239);
  not g35110 (n_15864, pi0772);
  and g35111 (n22241, n_15864, n_11736);
  and g35112 (n22242, pi0166, n22241);
  not g35113 (n_15865, n22242);
  and g35114 (n22243, pi0039, n_15865);
  not g35115 (n_15866, n22240);
  and g35116 (n22244, n_15866, n22243);
  not g35117 (n_15867, n22217);
  and g35118 (n22245, n_161, n_15867);
  not g35119 (n_15868, n22244);
  and g35120 (n22246, n_15868, n22245);
  not g35121 (n_15870, pi0727);
  not g35122 (n_15871, n22213);
  and g35123 (n22247, n_15870, n_15871);
  not g35124 (n_15872, n22246);
  and g35125 (n22248, n_15872, n22247);
  and g35126 (n22249, n21390, n22215);
  and g35127 (n22250, n_266, n_11418);
  not g35128 (n_15873, n22249);
  and g35129 (n22251, pi0038, n_15873);
  not g35130 (n_15874, n22250);
  and g35131 (n22252, n_15874, n22251);
  and g35132 (n22253, n_14975, n22217);
  and g35133 (n22254, n_11723, n16992);
  not g35134 (n_15875, n22254);
  and g35135 (n22255, n_266, n_15875);
  not g35136 (n_15876, n22255);
  and g35137 (n22256, n21055, n_15876);
  and g35138 (n22257, n_15143, n_15848);
  and g35139 (n22258, n2603, n22257);
  not g35140 (n_15877, n22258);
  and g35141 (n22259, n_223, n_15877);
  and g35142 (n22260, n_15207, n_15850);
  not g35143 (n_15878, n22260);
  and g35144 (n22261, n21435, n_15878);
  not g35145 (n_15879, n22261);
  and g35146 (n22262, n22259, n_15879);
  not g35147 (n_15880, n22256);
  and g35148 (n22263, n22220, n_15880);
  not g35149 (n_15881, n22262);
  and g35150 (n22264, n_15881, n22263);
  and g35151 (n22265, n_266, n_11729);
  not g35152 (n_15882, n22265);
  and g35153 (n22266, n20998, n_15882);
  and g35154 (n22267, n3448, n22257);
  not g35155 (n_15883, n22267);
  and g35156 (n22268, n_36, n_15883);
  and g35157 (n22269, n_15140, n22232);
  not g35158 (n_15884, n22269);
  and g35159 (n22270, n22268, n_15884);
  not g35160 (n_15885, n22266);
  and g35161 (n22271, pi0299, n_15885);
  not g35162 (n_15886, n22270);
  and g35163 (n22272, n_15886, n22271);
  not g35164 (n_15887, n22264);
  and g35165 (n22273, pi0772, n_15887);
  not g35166 (n_15888, n22272);
  and g35167 (n22274, n_15888, n22273);
  and g35168 (n22275, n_9349, n_15878);
  and g35169 (n22276, n2603, n21025);
  not g35170 (n_15889, n22276);
  and g35171 (n22277, n22259, n_15889);
  not g35172 (n_15890, n22275);
  and g35173 (n22278, n_15890, n22277);
  and g35174 (n22279, n_234, n_15880);
  not g35175 (n_15891, n22278);
  and g35176 (n22280, n_15891, n22279);
  and g35177 (n22281, n_14926, n22268);
  and g35178 (n22282, n_15856, n22281);
  and g35179 (n22283, n_15198, n22266);
  not g35180 (n_15892, n22283);
  and g35181 (n22284, pi0299, n_15892);
  not g35182 (n_15893, n22282);
  and g35183 (n22285, n_15893, n22284);
  not g35184 (n_15894, n22280);
  and g35185 (n22286, n_15864, n_15894);
  not g35186 (n_15895, n22285);
  and g35187 (n22287, n_15895, n22286);
  not g35188 (n_15896, n22274);
  and g35189 (n22288, pi0039, n_15896);
  not g35190 (n_15897, n22287);
  and g35191 (n22289, n_15897, n22288);
  not g35192 (n_15898, n22253);
  and g35193 (n22290, n_161, n_15898);
  not g35194 (n_15899, n22289);
  and g35195 (n22291, n_15899, n22290);
  not g35196 (n_15900, n22252);
  and g35197 (n22292, pi0727, n_15900);
  not g35198 (n_15901, n22291);
  and g35199 (n22293, n_15901, n22292);
  not g35200 (n_15902, n22248);
  not g35201 (n_15903, n22293);
  and g35202 (n22294, n_15902, n_15903);
  not g35203 (n_15904, n22294);
  and g35204 (n22295, n10197, n_15904);
  not g35205 (n_15905, n22208);
  and g35206 (n22296, n_12415, n_15905);
  not g35207 (n_15906, n22295);
  and g35208 (n22297, n_15906, n22296);
  and g35209 (n22298, n_266, n_12418);
  and g35210 (n22299, pi0727, n20902);
  and g35211 (n22300, n2926, n_15840);
  not g35212 (n_15907, n22299);
  and g35213 (n22301, n_15907, n22300);
  not g35214 (n_15908, n22298);
  and g35215 (n22302, pi0832, n_15908);
  not g35216 (n_15909, n22301);
  and g35217 (n22303, n_15909, n22302);
  or g35218 (po0323, n22297, n22303);
  and g35219 (n22305, n_6273, n_12418);
  not g35220 (n_15911, pi0768);
  and g35221 (n22306, n_15911, pi0947);
  and g35222 (n22307, pi0705, n20902);
  not g35223 (n_15913, n22306);
  not g35224 (n_15914, n22307);
  and g35225 (n22308, n_15913, n_15914);
  not g35226 (n_15915, n22308);
  and g35227 (n22309, n2926, n_15915);
  not g35228 (n_15916, n22305);
  and g35229 (n22310, pi0832, n_15916);
  not g35230 (n_15917, n22309);
  and g35231 (n22311, n_15917, n22310);
  and g35232 (n22312, n_6273, n_14814);
  and g35233 (n22313, pi0768, n_11743);
  and g35234 (n22314, n_6273, n22313);
  and g35235 (n22315, n_6273, n_11740);
  not g35236 (n_15918, n22315);
  and g35237 (n22316, n_15355, n_15918);
  and g35238 (n22317, pi0167, n21032);
  not g35239 (n_15919, n21006);
  and g35240 (n22318, n_6273, n_15919);
  not g35241 (n_15920, n22317);
  and g35242 (n22319, n_161, n_15920);
  not g35243 (n_15921, n22318);
  and g35244 (n22320, n_15921, n22319);
  not g35245 (n_15922, n22316);
  and g35246 (n22321, n_15911, n_15922);
  not g35247 (n_15923, n22320);
  and g35248 (n22322, n_15923, n22321);
  not g35249 (n_15924, pi0705);
  not g35250 (n_15925, n22314);
  and g35251 (n22323, n_15924, n_15925);
  not g35252 (n_15926, n22322);
  and g35253 (n22324, n_15926, n22323);
  and g35254 (n22325, n_6273, n_11418);
  not g35255 (n_15927, n22325);
  and g35256 (n22326, n21090, n_15927);
  and g35257 (n22327, n_6273, n21099);
  and g35258 (n22328, pi0167, n21116);
  not g35259 (n_15928, n22328);
  and g35260 (n22329, n_161, n_15928);
  not g35261 (n_15929, n22327);
  and g35262 (n22330, n_15929, n22329);
  not g35263 (n_15930, n22326);
  and g35264 (n22331, pi0768, n_15930);
  not g35265 (n_15931, n22330);
  and g35266 (n22332, n_15931, n22331);
  and g35267 (n22333, n_6273, n_14920);
  not g35268 (n_15932, n22333);
  and g35269 (n22334, n21042, n_15932);
  and g35270 (n22335, n_6273, n21069);
  and g35271 (n22336, pi0167, n21082);
  not g35272 (n_15933, n22336);
  and g35273 (n22337, n_161, n_15933);
  not g35274 (n_15934, n22335);
  and g35275 (n22338, n_15934, n22337);
  not g35276 (n_15935, n22334);
  and g35277 (n22339, n_15911, n_15935);
  not g35278 (n_15936, n22338);
  and g35279 (n22340, n_15936, n22339);
  not g35280 (n_15937, n22332);
  and g35281 (n22341, pi0705, n_15937);
  not g35282 (n_15938, n22340);
  and g35283 (n22342, n_15938, n22341);
  not g35284 (n_15939, n22324);
  and g35285 (n22343, n10197, n_15939);
  not g35286 (n_15940, n22342);
  and g35287 (n22344, n_15940, n22343);
  not g35288 (n_15941, n22312);
  and g35289 (n22345, n_12415, n_15941);
  not g35290 (n_15942, n22344);
  and g35291 (n22346, n_15942, n22345);
  not g35292 (n_15943, n22311);
  not g35293 (n_15944, n22346);
  and g35294 (po0324, n_15943, n_15944);
  and g35295 (n22348, pi0168, n_12418);
  and g35296 (n22349, pi0763, pi0947);
  not g35297 (n_15946, n22349);
  and g35298 (n22350, n2926, n_15946);
  and g35299 (n22351, pi0699, n20902);
  not g35300 (n_15948, n22351);
  and g35301 (n22352, n22350, n_15948);
  not g35302 (n_15949, n22348);
  and g35303 (n22353, pi0832, n_15949);
  not g35304 (n_15950, n22352);
  and g35305 (n22354, n_15950, n22353);
  and g35306 (n22355, pi0057, pi0168);
  and g35307 (n22356, n_2206, n_14990);
  and g35308 (n22357, n_2206, n_11674);
  not g35309 (n_15951, pi0763);
  and g35310 (n22358, n_15951, n18147);
  not g35311 (n_15952, n22358);
  and g35312 (n22359, n_14913, n_15952);
  not g35313 (n_15953, n22357);
  not g35314 (n_15954, n22359);
  and g35315 (n22360, n_15953, n_15954);
  and g35316 (n22361, n_14975, n22360);
  and g35317 (n22362, n_2206, n_11719);
  not g35318 (n_15955, n22362);
  and g35319 (n22363, n21111, n_15955);
  and g35320 (n22364, pi0168, n_11729);
  not g35321 (n_15956, n22364);
  and g35322 (n22365, n20998, n_15956);
  not g35323 (n_15957, n22365);
  and g35324 (n22366, n21073, n_15957);
  and g35325 (n22367, pi0168, n_9350);
  and g35326 (n22368, n_15140, n22367);
  not g35327 (n_15958, n22368);
  and g35328 (n22369, n_11726, n_15958);
  and g35329 (n22370, n_2206, n_11445);
  not g35330 (n_15959, n22370);
  and g35331 (n22371, n21105, n_15959);
  not g35332 (n_15960, n22371);
  and g35333 (n22372, n_14925, n_15960);
  and g35334 (n22373, n22369, n22372);
  not g35335 (n_15961, n22373);
  and g35336 (n22374, n_36, n_15961);
  not g35337 (n_15962, n22366);
  and g35338 (n22375, n_14904, n_15962);
  not g35339 (n_15963, n22374);
  and g35340 (n22376, n_15963, n22375);
  not g35341 (n_15964, n22376);
  and g35342 (n22377, pi0299, n_15964);
  not g35343 (n_15965, n22363);
  and g35344 (n22378, n_15951, n_15965);
  not g35345 (n_15966, n22377);
  and g35346 (n22379, n_15966, n22378);
  and g35347 (n22380, n21026, n_15959);
  and g35348 (n22381, n_15287, n22380);
  not g35349 (n_15967, n22381);
  and g35350 (n22382, n_36, n_15967);
  and g35351 (n22383, n22369, n22382);
  not g35352 (n_15968, n22383);
  and g35353 (n22384, n_15957, n_15968);
  not g35354 (n_15969, n22384);
  and g35355 (n22385, pi0299, n_15969);
  and g35356 (n22386, pi0168, n_15148);
  not g35357 (n_15970, n22386);
  and g35358 (n22387, n21062, n_15970);
  not g35359 (n_15971, n22385);
  not g35360 (n_15972, n22387);
  and g35361 (n22388, n_15971, n_15972);
  not g35362 (n_15973, n22388);
  and g35363 (n22389, pi0763, n_15973);
  not g35364 (n_15974, n22379);
  and g35365 (n22390, pi0039, n_15974);
  not g35366 (n_15975, n22389);
  and g35367 (n22391, n_15975, n22390);
  not g35368 (n_15976, n22361);
  not g35369 (n_15977, n22391);
  and g35370 (n22392, n_15976, n_15977);
  not g35371 (n_15978, n22392);
  and g35372 (n22393, n_161, n_15978);
  and g35373 (n22394, n_2206, n_11418);
  and g35374 (n22395, n_15951, pi0947);
  not g35375 (n_15979, n22395);
  and g35376 (n22396, n_162, n_15979);
  and g35377 (n22397, n21239, n22396);
  not g35378 (n_15980, n22394);
  and g35379 (n22398, pi0038, n_15980);
  not g35380 (n_15981, n22397);
  and g35381 (n22399, n_15981, n22398);
  not g35382 (n_15982, n22393);
  not g35383 (n_15983, n22399);
  and g35384 (n22400, n_15982, n_15983);
  not g35385 (n_15984, n22400);
  and g35386 (n22401, pi0699, n_15984);
  and g35387 (n22402, n6284, n22350);
  and g35388 (n22403, pi0168, n_11740);
  not g35389 (n_15985, n22402);
  and g35390 (n22404, pi0038, n_15985);
  not g35391 (n_15986, n22403);
  and g35392 (n22405, n_15986, n22404);
  and g35393 (n22406, n21019, n_15955);
  and g35394 (n22407, n21000, n_15956);
  not g35395 (n_15987, n22380);
  and g35396 (n22408, n22369, n_15987);
  and g35397 (n22409, n20996, n22408);
  not g35398 (n_15988, n22407);
  and g35399 (n22410, pi0299, n_15988);
  not g35400 (n_15989, n22409);
  and g35401 (n22411, n_15989, n22410);
  not g35402 (n_15990, n22411);
  and g35403 (n22412, pi0763, n_15990);
  not g35404 (n_15991, n22406);
  and g35405 (n22413, n_15991, n22412);
  and g35406 (n22414, n_2206, n_15951);
  and g35407 (n22415, n_11736, n22414);
  not g35408 (n_15992, n22415);
  and g35409 (n22416, pi0039, n_15992);
  not g35410 (n_15993, n22413);
  and g35411 (n22417, n_15993, n22416);
  not g35412 (n_15994, n22360);
  and g35413 (n22418, n_161, n_15994);
  not g35414 (n_15995, n22417);
  and g35415 (n22419, n_15995, n22418);
  not g35416 (n_15996, pi0699);
  not g35417 (n_15997, n22405);
  and g35418 (n22420, n_15996, n_15997);
  not g35419 (n_15998, n22419);
  and g35420 (n22421, n_15998, n22420);
  not g35421 (n_15999, n22421);
  and g35422 (n22422, n21130, n_15999);
  not g35423 (n_16000, n22401);
  and g35424 (n22423, n_16000, n22422);
  not g35425 (n_16001, n22356);
  and g35426 (n22424, n_796, n_16001);
  not g35427 (n_16002, n22423);
  and g35428 (n22425, n_16002, n22424);
  not g35429 (n_16003, n22355);
  and g35430 (n22426, n_12415, n_16003);
  not g35431 (n_16004, n22425);
  and g35432 (n22427, n_16004, n22426);
  or g35433 (po0325, n22354, n22427);
  and g35434 (n22429, pi0169, n_12418);
  and g35435 (n22430, pi0746, pi0947);
  not g35436 (n_16006, n22430);
  and g35437 (n22431, n2926, n_16006);
  and g35438 (n22432, pi0729, n20902);
  not g35439 (n_16008, n22432);
  and g35440 (n22433, n22431, n_16008);
  not g35441 (n_16009, n22429);
  and g35442 (n22434, pi0832, n_16009);
  not g35443 (n_16010, n22433);
  and g35444 (n22435, n_16010, n22434);
  and g35445 (n22436, pi0057, pi0169);
  and g35446 (n22437, n_2027, n_14990);
  and g35447 (n22438, n_2027, n_11674);
  not g35448 (n_16011, pi0746);
  and g35449 (n22439, n_16011, n18147);
  not g35450 (n_16012, n22439);
  and g35451 (n22440, n_14913, n_16012);
  not g35452 (n_16013, n22438);
  not g35453 (n_16014, n22440);
  and g35454 (n22441, n_16013, n_16014);
  and g35455 (n22442, n_14975, n22441);
  and g35456 (n22443, n_2027, n_11719);
  not g35457 (n_16015, n22443);
  and g35458 (n22444, n21111, n_16015);
  and g35459 (n22445, pi0169, n_11729);
  not g35460 (n_16016, n22445);
  and g35461 (n22446, n20998, n_16016);
  not g35462 (n_16017, n22446);
  and g35463 (n22447, n21073, n_16017);
  and g35464 (n22448, pi0169, n_9350);
  and g35465 (n22449, n_15140, n22448);
  not g35466 (n_16018, n22449);
  and g35467 (n22450, n_11726, n_16018);
  and g35468 (n22451, n_2027, n_11445);
  not g35469 (n_16019, n22451);
  and g35470 (n22452, n21105, n_16019);
  not g35471 (n_16020, n22452);
  and g35472 (n22453, n_14925, n_16020);
  and g35473 (n22454, n22450, n22453);
  not g35474 (n_16021, n22454);
  and g35475 (n22455, n_36, n_16021);
  not g35476 (n_16022, n22447);
  and g35477 (n22456, n_14904, n_16022);
  not g35478 (n_16023, n22455);
  and g35479 (n22457, n_16023, n22456);
  not g35480 (n_16024, n22457);
  and g35481 (n22458, pi0299, n_16024);
  not g35482 (n_16025, n22444);
  and g35483 (n22459, n_16011, n_16025);
  not g35484 (n_16026, n22458);
  and g35485 (n22460, n_16026, n22459);
  and g35486 (n22461, n21026, n_16019);
  and g35487 (n22462, n_15287, n22461);
  not g35488 (n_16027, n22462);
  and g35489 (n22463, n_36, n_16027);
  and g35490 (n22464, n22450, n22463);
  not g35491 (n_16028, n22464);
  and g35492 (n22465, n_16017, n_16028);
  not g35493 (n_16029, n22465);
  and g35494 (n22466, pi0299, n_16029);
  and g35495 (n22467, pi0169, n_15148);
  not g35496 (n_16030, n22467);
  and g35497 (n22468, n21062, n_16030);
  not g35498 (n_16031, n22466);
  not g35499 (n_16032, n22468);
  and g35500 (n22469, n_16031, n_16032);
  not g35501 (n_16033, n22469);
  and g35502 (n22470, pi0746, n_16033);
  not g35503 (n_16034, n22460);
  and g35504 (n22471, pi0039, n_16034);
  not g35505 (n_16035, n22470);
  and g35506 (n22472, n_16035, n22471);
  not g35507 (n_16036, n22442);
  not g35508 (n_16037, n22472);
  and g35509 (n22473, n_16036, n_16037);
  not g35510 (n_16038, n22473);
  and g35511 (n22474, n_161, n_16038);
  and g35512 (n22475, n_2027, n_11418);
  and g35513 (n22476, n_16011, pi0947);
  not g35514 (n_16039, n22476);
  and g35515 (n22477, n_162, n_16039);
  and g35516 (n22478, n21239, n22477);
  not g35517 (n_16040, n22475);
  and g35518 (n22479, pi0038, n_16040);
  not g35519 (n_16041, n22478);
  and g35520 (n22480, n_16041, n22479);
  not g35521 (n_16042, n22474);
  not g35522 (n_16043, n22480);
  and g35523 (n22481, n_16042, n_16043);
  not g35524 (n_16044, n22481);
  and g35525 (n22482, pi0729, n_16044);
  and g35526 (n22483, n6284, n22431);
  and g35527 (n22484, pi0169, n_11740);
  not g35528 (n_16045, n22483);
  and g35529 (n22485, pi0038, n_16045);
  not g35530 (n_16046, n22484);
  and g35531 (n22486, n_16046, n22485);
  and g35532 (n22487, n21019, n_16015);
  and g35533 (n22488, n21000, n_16016);
  not g35534 (n_16047, n22461);
  and g35535 (n22489, n22450, n_16047);
  and g35536 (n22490, n20996, n22489);
  not g35537 (n_16048, n22488);
  and g35538 (n22491, pi0299, n_16048);
  not g35539 (n_16049, n22490);
  and g35540 (n22492, n_16049, n22491);
  not g35541 (n_16050, n22492);
  and g35542 (n22493, pi0746, n_16050);
  not g35543 (n_16051, n22487);
  and g35544 (n22494, n_16051, n22493);
  and g35545 (n22495, n_2027, n_16011);
  and g35546 (n22496, n_11736, n22495);
  not g35547 (n_16052, n22496);
  and g35548 (n22497, pi0039, n_16052);
  not g35549 (n_16053, n22494);
  and g35550 (n22498, n_16053, n22497);
  not g35551 (n_16054, n22441);
  and g35552 (n22499, n_161, n_16054);
  not g35553 (n_16055, n22498);
  and g35554 (n22500, n_16055, n22499);
  not g35555 (n_16056, pi0729);
  not g35556 (n_16057, n22486);
  and g35557 (n22501, n_16056, n_16057);
  not g35558 (n_16058, n22500);
  and g35559 (n22502, n_16058, n22501);
  not g35560 (n_16059, n22502);
  and g35561 (n22503, n21130, n_16059);
  not g35562 (n_16060, n22482);
  and g35563 (n22504, n_16060, n22503);
  not g35564 (n_16061, n22437);
  and g35565 (n22505, n_796, n_16061);
  not g35566 (n_16062, n22504);
  and g35567 (n22506, n_16062, n22505);
  not g35568 (n_16063, n22436);
  and g35569 (n22507, n_12415, n_16063);
  not g35570 (n_16064, n22506);
  and g35571 (n22508, n_16064, n22507);
  or g35572 (po0326, n22435, n22508);
  and g35573 (n22510, pi0730, n20902);
  and g35574 (n22511, pi0748, pi0947);
  not g35575 (n_16067, n22511);
  and g35576 (n22512, n2926, n_16067);
  not g35577 (n_16068, n22510);
  and g35578 (n22513, n_16068, n22512);
  and g35579 (n22514, pi0170, n_12418);
  not g35580 (n_16069, n22514);
  and g35581 (n22515, pi0832, n_16069);
  not g35582 (n_16070, n22513);
  and g35583 (n22516, n_16070, n22515);
  and g35584 (n22517, pi0057, pi0170);
  and g35585 (n22518, n_1673, n_14990);
  and g35586 (n22519, n_1673, n_11418);
  not g35587 (n_16071, n22519);
  and g35588 (n22520, n21090, n_16071);
  and g35589 (n22521, pi0170, n_11729);
  not g35590 (n_16072, n22521);
  and g35591 (n22522, n20998, n_16072);
  not g35592 (n_16073, n22522);
  and g35593 (n22523, n21073, n_16073);
  and g35594 (n22524, pi0170, n_9350);
  and g35595 (n22525, n_15140, n22524);
  not g35596 (n_16074, n22525);
  and g35597 (n22526, n_11726, n_16074);
  and g35598 (n22527, n_1673, n_11445);
  not g35599 (n_16075, n22527);
  and g35600 (n22528, n21105, n_16075);
  not g35601 (n_16076, n22528);
  and g35602 (n22529, n_14925, n_16076);
  and g35603 (n22530, n22526, n22529);
  not g35604 (n_16077, n22530);
  and g35605 (n22531, n_36, n_16077);
  not g35606 (n_16078, n22523);
  and g35607 (n22532, n_14904, n_16078);
  not g35608 (n_16079, n22531);
  and g35609 (n22533, n_16079, n22532);
  not g35610 (n_16080, n22533);
  and g35611 (n22534, pi0299, n_16080);
  and g35612 (n22535, n_1673, n_11719);
  not g35613 (n_16081, n22535);
  and g35614 (n22536, n_234, n_16081);
  and g35615 (n22537, n_14971, n22536);
  not g35616 (n_16082, n22534);
  not g35617 (n_16083, n22537);
  and g35618 (n22538, n_16082, n_16083);
  not g35619 (n_16084, n22538);
  and g35620 (n22539, pi0039, n_16084);
  and g35621 (n22540, n_1673, n_11674);
  not g35622 (n_16085, n22540);
  and g35623 (n22541, n21115, n_16085);
  not g35624 (n_16086, n22539);
  not g35625 (n_16087, n22541);
  and g35626 (n22542, n_16086, n_16087);
  not g35627 (n_16088, n22542);
  and g35628 (n22543, n_161, n_16088);
  not g35629 (n_16089, pi0748);
  not g35630 (n_16090, n22520);
  and g35631 (n22544, n_16089, n_16090);
  not g35632 (n_16091, n22543);
  and g35633 (n22545, n_16091, n22544);
  and g35634 (n22546, n21042, n_16071);
  and g35635 (n22547, n21067, n_16085);
  and g35636 (n22548, n21026, n_16075);
  and g35637 (n22549, n_15287, n22548);
  not g35638 (n_16092, n22549);
  and g35639 (n22550, n_36, n_16092);
  and g35640 (n22551, n22526, n22550);
  not g35641 (n_16093, n22551);
  and g35642 (n22552, n_16073, n_16093);
  not g35643 (n_16094, n22552);
  and g35644 (n22553, pi0299, n_16094);
  and g35645 (n22554, pi0170, n_15148);
  not g35646 (n_16095, n22554);
  and g35647 (n22555, n21062, n_16095);
  not g35648 (n_16096, n22553);
  and g35649 (n22556, pi0039, n_16096);
  not g35650 (n_16097, n22555);
  and g35651 (n22557, n_16097, n22556);
  not g35652 (n_16098, n22547);
  not g35653 (n_16099, n22557);
  and g35654 (n22558, n_16098, n_16099);
  not g35655 (n_16100, n22558);
  and g35656 (n22559, n_161, n_16100);
  not g35657 (n_16101, n22546);
  and g35658 (n22560, pi0748, n_16101);
  not g35659 (n_16102, n22559);
  and g35660 (n22561, n_16102, n22560);
  not g35661 (n_16103, n22561);
  and g35662 (n22562, pi0730, n_16103);
  not g35663 (n_16104, n22545);
  and g35664 (n22563, n_16104, n22562);
  and g35665 (n22564, n_1673, n_11740);
  not g35666 (n_16105, n22564);
  and g35667 (n22565, n_15355, n_16105);
  and g35668 (n22566, n21017, n_16085);
  and g35669 (n22567, n21000, n_16072);
  not g35670 (n_16106, n22548);
  and g35671 (n22568, n22526, n_16106);
  and g35672 (n22569, n20996, n22568);
  not g35673 (n_16107, n22567);
  and g35674 (n22570, pi0299, n_16107);
  not g35675 (n_16108, n22569);
  and g35676 (n22571, n_16108, n22570);
  and g35677 (n22572, n_14903, n22536);
  not g35678 (n_16109, n22571);
  not g35679 (n_16110, n22572);
  and g35680 (n22573, n_16109, n_16110);
  not g35681 (n_16111, n22573);
  and g35682 (n22574, pi0039, n_16111);
  not g35683 (n_16112, n22566);
  not g35684 (n_16113, n22574);
  and g35685 (n22575, n_16112, n_16113);
  not g35686 (n_16114, n22575);
  and g35687 (n22576, n_161, n_16114);
  not g35688 (n_16115, n22565);
  and g35689 (n22577, pi0748, n_16115);
  not g35690 (n_16116, n22576);
  and g35691 (n22578, n_16116, n22577);
  and g35692 (n22579, n_1673, n_16089);
  and g35693 (n22580, n_11743, n22579);
  not g35694 (n_16117, pi0730);
  not g35695 (n_16118, n22580);
  and g35696 (n22581, n_16117, n_16118);
  not g35697 (n_16119, n22578);
  and g35698 (n22582, n_16119, n22581);
  not g35699 (n_16120, n22582);
  and g35700 (n22583, n21130, n_16120);
  not g35701 (n_16121, n22563);
  and g35702 (n22584, n_16121, n22583);
  not g35703 (n_16122, n22518);
  and g35704 (n22585, n_796, n_16122);
  not g35705 (n_16123, n22584);
  and g35706 (n22586, n_16123, n22585);
  not g35707 (n_16124, n22517);
  and g35708 (n22587, n_12415, n_16124);
  not g35709 (n_16125, n22586);
  and g35710 (n22588, n_16125, n22587);
  or g35711 (po0327, n22516, n22588);
  and g35712 (n22590, pi0171, n_12418);
  and g35713 (n22591, pi0764, pi0947);
  not g35714 (n_16127, n22591);
  and g35715 (n22592, n2926, n_16127);
  and g35716 (n22593, pi0691, n20902);
  not g35717 (n_16129, n22593);
  and g35718 (n22594, n22592, n_16129);
  not g35719 (n_16130, n22590);
  and g35720 (n22595, pi0832, n_16130);
  not g35721 (n_16131, n22594);
  and g35722 (n22596, n_16131, n22595);
  and g35723 (n22597, pi0057, pi0171);
  and g35724 (n22598, n_1493, n_14990);
  and g35725 (n22599, n_1493, n_11674);
  not g35726 (n_16132, pi0764);
  and g35727 (n22600, n_16132, n18147);
  not g35728 (n_16133, n22600);
  and g35729 (n22601, n_14913, n_16133);
  not g35730 (n_16134, n22599);
  not g35731 (n_16135, n22601);
  and g35732 (n22602, n_16134, n_16135);
  and g35733 (n22603, n_14975, n22602);
  and g35734 (n22604, n_1493, n_11719);
  not g35735 (n_16136, n22604);
  and g35736 (n22605, n21111, n_16136);
  and g35737 (n22606, pi0171, n_11729);
  not g35738 (n_16137, n22606);
  and g35739 (n22607, n20998, n_16137);
  not g35740 (n_16138, n22607);
  and g35741 (n22608, n21073, n_16138);
  and g35742 (n22609, pi0171, n_9350);
  and g35743 (n22610, n_15140, n22609);
  not g35744 (n_16139, n22610);
  and g35745 (n22611, n_11726, n_16139);
  and g35746 (n22612, n_1493, n_11445);
  not g35747 (n_16140, n22612);
  and g35748 (n22613, n21105, n_16140);
  not g35749 (n_16141, n22613);
  and g35750 (n22614, n_14925, n_16141);
  and g35751 (n22615, n22611, n22614);
  not g35752 (n_16142, n22615);
  and g35753 (n22616, n_36, n_16142);
  not g35754 (n_16143, n22608);
  and g35755 (n22617, n_14904, n_16143);
  not g35756 (n_16144, n22616);
  and g35757 (n22618, n_16144, n22617);
  not g35758 (n_16145, n22618);
  and g35759 (n22619, pi0299, n_16145);
  not g35760 (n_16146, n22605);
  and g35761 (n22620, n_16132, n_16146);
  not g35762 (n_16147, n22619);
  and g35763 (n22621, n_16147, n22620);
  and g35764 (n22622, n21026, n_16140);
  and g35765 (n22623, n_15287, n22622);
  not g35766 (n_16148, n22623);
  and g35767 (n22624, n_36, n_16148);
  and g35768 (n22625, n22611, n22624);
  not g35769 (n_16149, n22625);
  and g35770 (n22626, n_16138, n_16149);
  not g35771 (n_16150, n22626);
  and g35772 (n22627, pi0299, n_16150);
  and g35773 (n22628, pi0171, n_15148);
  not g35774 (n_16151, n22628);
  and g35775 (n22629, n21062, n_16151);
  not g35776 (n_16152, n22627);
  not g35777 (n_16153, n22629);
  and g35778 (n22630, n_16152, n_16153);
  not g35779 (n_16154, n22630);
  and g35780 (n22631, pi0764, n_16154);
  not g35781 (n_16155, n22621);
  and g35782 (n22632, pi0039, n_16155);
  not g35783 (n_16156, n22631);
  and g35784 (n22633, n_16156, n22632);
  not g35785 (n_16157, n22603);
  not g35786 (n_16158, n22633);
  and g35787 (n22634, n_16157, n_16158);
  not g35788 (n_16159, n22634);
  and g35789 (n22635, n_161, n_16159);
  and g35790 (n22636, n_1493, n_11418);
  and g35791 (n22637, n_16132, pi0947);
  not g35792 (n_16160, n22637);
  and g35793 (n22638, n_162, n_16160);
  and g35794 (n22639, n21239, n22638);
  not g35795 (n_16161, n22636);
  and g35796 (n22640, pi0038, n_16161);
  not g35797 (n_16162, n22639);
  and g35798 (n22641, n_16162, n22640);
  not g35799 (n_16163, n22635);
  not g35800 (n_16164, n22641);
  and g35801 (n22642, n_16163, n_16164);
  not g35802 (n_16165, n22642);
  and g35803 (n22643, pi0691, n_16165);
  and g35804 (n22644, n6284, n22592);
  and g35805 (n22645, pi0171, n_11740);
  not g35806 (n_16166, n22644);
  and g35807 (n22646, pi0038, n_16166);
  not g35808 (n_16167, n22645);
  and g35809 (n22647, n_16167, n22646);
  and g35810 (n22648, n21019, n_16136);
  and g35811 (n22649, n21000, n_16137);
  not g35812 (n_16168, n22622);
  and g35813 (n22650, n22611, n_16168);
  and g35814 (n22651, n20996, n22650);
  not g35815 (n_16169, n22649);
  and g35816 (n22652, pi0299, n_16169);
  not g35817 (n_16170, n22651);
  and g35818 (n22653, n_16170, n22652);
  not g35819 (n_16171, n22653);
  and g35820 (n22654, pi0764, n_16171);
  not g35821 (n_16172, n22648);
  and g35822 (n22655, n_16172, n22654);
  and g35823 (n22656, n_1493, n_16132);
  and g35824 (n22657, n_11736, n22656);
  not g35825 (n_16173, n22657);
  and g35826 (n22658, pi0039, n_16173);
  not g35827 (n_16174, n22655);
  and g35828 (n22659, n_16174, n22658);
  not g35829 (n_16175, n22602);
  and g35830 (n22660, n_161, n_16175);
  not g35831 (n_16176, n22659);
  and g35832 (n22661, n_16176, n22660);
  not g35833 (n_16177, pi0691);
  not g35834 (n_16178, n22647);
  and g35835 (n22662, n_16177, n_16178);
  not g35836 (n_16179, n22661);
  and g35837 (n22663, n_16179, n22662);
  not g35838 (n_16180, n22663);
  and g35839 (n22664, n21130, n_16180);
  not g35840 (n_16181, n22643);
  and g35841 (n22665, n_16181, n22664);
  not g35842 (n_16182, n22598);
  and g35843 (n22666, n_796, n_16182);
  not g35844 (n_16183, n22665);
  and g35845 (n22667, n_16183, n22666);
  not g35846 (n_16184, n22597);
  and g35847 (n22668, n_12415, n_16184);
  not g35848 (n_16185, n22667);
  and g35849 (n22669, n_16185, n22668);
  or g35850 (po0328, n22596, n22669);
  and g35851 (n22671, pi0172, n_12418);
  and g35852 (n22672, pi0739, pi0947);
  not g35853 (n_16187, n22672);
  and g35854 (n22673, n2926, n_16187);
  and g35855 (n22674, pi0690, n20902);
  not g35856 (n_16189, n22674);
  and g35857 (n22675, n22673, n_16189);
  not g35858 (n_16190, n22671);
  and g35859 (n22676, pi0832, n_16190);
  not g35860 (n_16191, n22675);
  and g35861 (n22677, n_16191, n22676);
  and g35862 (n22678, pi0057, pi0172);
  and g35863 (n22679, n_1362, n_14990);
  and g35864 (n22680, n_1362, n_11674);
  and g35865 (n22681, n16958, n22672);
  not g35866 (n_16192, n22680);
  and g35867 (n22682, n_162, n_16192);
  not g35868 (n_16193, n22681);
  and g35869 (n22683, n_16193, n22682);
  and g35870 (n22684, n_14975, n22683);
  and g35871 (n22685, n_1362, n_11719);
  not g35872 (n_16194, n22685);
  and g35873 (n22686, n21111, n_16194);
  and g35874 (n22687, pi0172, n_11729);
  not g35875 (n_16195, n22687);
  and g35876 (n22688, n20998, n_16195);
  not g35877 (n_16196, n22688);
  and g35878 (n22689, n21073, n_16196);
  and g35879 (n22690, pi0172, n_9350);
  and g35880 (n22691, n_15140, n22690);
  not g35881 (n_16197, n22691);
  and g35882 (n22692, n_11726, n_16197);
  and g35883 (n22693, n_1362, n_11445);
  not g35884 (n_16198, n22693);
  and g35885 (n22694, n21105, n_16198);
  not g35886 (n_16199, n22694);
  and g35887 (n22695, n_14925, n_16199);
  and g35888 (n22696, n22692, n22695);
  not g35889 (n_16200, n22696);
  and g35890 (n22697, n_36, n_16200);
  not g35891 (n_16201, n22689);
  and g35892 (n22698, n_14904, n_16201);
  not g35893 (n_16202, n22697);
  and g35894 (n22699, n_16202, n22698);
  not g35895 (n_16203, n22699);
  and g35896 (n22700, pi0299, n_16203);
  not g35897 (n_16204, pi0739);
  not g35898 (n_16205, n22686);
  and g35899 (n22701, n_16204, n_16205);
  not g35900 (n_16206, n22700);
  and g35901 (n22702, n_16206, n22701);
  and g35902 (n22703, n21026, n_16198);
  and g35903 (n22704, n_15287, n22703);
  not g35904 (n_16207, n22704);
  and g35905 (n22705, n_36, n_16207);
  and g35906 (n22706, n22692, n22705);
  not g35907 (n_16208, n22706);
  and g35908 (n22707, n_16196, n_16208);
  not g35909 (n_16209, n22707);
  and g35910 (n22708, pi0299, n_16209);
  and g35911 (n22709, pi0172, n_15148);
  not g35912 (n_16210, n22709);
  and g35913 (n22710, n21062, n_16210);
  not g35914 (n_16211, n22708);
  not g35915 (n_16212, n22710);
  and g35916 (n22711, n_16211, n_16212);
  not g35917 (n_16213, n22711);
  and g35918 (n22712, pi0739, n_16213);
  not g35919 (n_16214, n22702);
  and g35920 (n22713, pi0039, n_16214);
  not g35921 (n_16215, n22712);
  and g35922 (n22714, n_16215, n22713);
  not g35923 (n_16216, n22684);
  not g35924 (n_16217, n22714);
  and g35925 (n22715, n_16216, n_16217);
  not g35926 (n_16218, n22715);
  and g35927 (n22716, n_161, n_16218);
  and g35928 (n22717, n_1362, n_11418);
  and g35929 (n22718, n_16204, pi0947);
  not g35930 (n_16219, n22718);
  and g35931 (n22719, n_162, n_16219);
  and g35932 (n22720, n21239, n22719);
  not g35933 (n_16220, n22717);
  and g35934 (n22721, pi0038, n_16220);
  not g35935 (n_16221, n22720);
  and g35936 (n22722, n_16221, n22721);
  not g35937 (n_16222, n22716);
  not g35938 (n_16223, n22722);
  and g35939 (n22723, n_16222, n_16223);
  not g35940 (n_16224, n22723);
  and g35941 (n22724, pi0690, n_16224);
  and g35942 (n22725, n6284, n22673);
  and g35943 (n22726, pi0172, n_11740);
  not g35944 (n_16225, n22725);
  and g35945 (n22727, pi0038, n_16225);
  not g35946 (n_16226, n22726);
  and g35947 (n22728, n_16226, n22727);
  and g35948 (n22729, n21019, n_16194);
  and g35949 (n22730, n21000, n_16195);
  not g35950 (n_16227, n22703);
  and g35951 (n22731, n22692, n_16227);
  and g35952 (n22732, n20996, n22731);
  not g35953 (n_16228, n22730);
  and g35954 (n22733, pi0299, n_16228);
  not g35955 (n_16229, n22732);
  and g35956 (n22734, n_16229, n22733);
  not g35957 (n_16230, n22734);
  and g35958 (n22735, pi0739, n_16230);
  not g35959 (n_16231, n22729);
  and g35960 (n22736, n_16231, n22735);
  and g35961 (n22737, n_1362, n_16204);
  and g35962 (n22738, n_11736, n22737);
  not g35963 (n_16232, n22738);
  and g35964 (n22739, pi0039, n_16232);
  not g35965 (n_16233, n22736);
  and g35966 (n22740, n_16233, n22739);
  not g35967 (n_16234, n22683);
  and g35968 (n22741, n_161, n_16234);
  not g35969 (n_16235, n22740);
  and g35970 (n22742, n_16235, n22741);
  not g35971 (n_16236, pi0690);
  not g35972 (n_16237, n22728);
  and g35973 (n22743, n_16236, n_16237);
  not g35974 (n_16238, n22742);
  and g35975 (n22744, n_16238, n22743);
  not g35976 (n_16239, n22744);
  and g35977 (n22745, n21130, n_16239);
  not g35978 (n_16240, n22724);
  and g35979 (n22746, n_16240, n22745);
  not g35980 (n_16241, n22679);
  and g35981 (n22747, n_796, n_16241);
  not g35982 (n_16242, n22746);
  and g35983 (n22748, n_16242, n22747);
  not g35984 (n_16243, n22678);
  and g35985 (n22749, n_12415, n_16243);
  not g35986 (n_16244, n22748);
  and g35987 (n22750, n_16244, n22749);
  or g35988 (po0329, n22677, n22750);
  and g35989 (n22752, n_9183, po1038);
  and g35990 (n22753, n_9183, n_11751);
  not g35991 (n_16245, n22753);
  and g35992 (n22754, n16635, n_16245);
  and g35993 (n22755, n_15127, n2571);
  not g35994 (n_16246, n22755);
  and g35995 (n22756, n22753, n_16246);
  and g35996 (n22757, n_9183, n_11418);
  not g35997 (n_16247, n22757);
  and g35998 (n22758, n16647, n_16247);
  and g35999 (n22759, pi0173, n_12608);
  not g36000 (n_16248, n22759);
  and g36001 (n22760, n_161, n_16248);
  not g36002 (n_16249, n22760);
  and g36003 (n22761, n2571, n_16249);
  and g36004 (n22762, n_9183, n18072);
  not g36005 (n_16250, n22761);
  not g36006 (n_16251, n22762);
  and g36007 (n22763, n_16250, n_16251);
  not g36008 (n_16252, n22758);
  and g36009 (n22764, n_15127, n_16252);
  not g36010 (n_16253, n22763);
  and g36011 (n22765, n_16253, n22764);
  not g36012 (n_16254, n22756);
  not g36013 (n_16255, n22765);
  and g36014 (n22766, n_16254, n_16255);
  and g36015 (n22767, n_11749, n22766);
  and g36016 (n22768, n_11753, n22753);
  not g36017 (n_16256, n22766);
  and g36018 (n22769, pi0625, n_16256);
  not g36019 (n_16257, n22768);
  and g36020 (n22770, pi1153, n_16257);
  not g36021 (n_16258, n22769);
  and g36022 (n22771, n_16258, n22770);
  and g36023 (n22772, pi0625, n22753);
  and g36024 (n22773, n_11753, n_16256);
  not g36025 (n_16259, n22772);
  and g36026 (n22774, n_11757, n_16259);
  not g36027 (n_16260, n22773);
  and g36028 (n22775, n_16260, n22774);
  not g36029 (n_16261, n22771);
  not g36030 (n_16262, n22775);
  and g36031 (n22776, n_16261, n_16262);
  not g36032 (n_16263, n22776);
  and g36033 (n22777, pi0778, n_16263);
  not g36034 (n_16264, n22767);
  not g36035 (n_16265, n22777);
  and g36036 (n22778, n_16264, n_16265);
  not g36037 (n_16266, n22778);
  and g36038 (n22779, n_11773, n_16266);
  and g36039 (n22780, n17075, n_16245);
  not g36040 (n_16267, n22779);
  not g36041 (n_16268, n22780);
  and g36042 (n22781, n_16267, n_16268);
  and g36043 (n22782, n_11777, n22781);
  and g36044 (n22783, n16639, n22753);
  not g36045 (n_16269, n22782);
  not g36046 (n_16270, n22783);
  and g36047 (n22784, n_16269, n_16270);
  and g36048 (n22785, n_11780, n22784);
  not g36049 (n_16271, n22754);
  not g36050 (n_16272, n22785);
  and g36051 (n22786, n_16271, n_16272);
  and g36052 (n22787, n_11783, n22786);
  and g36053 (n22788, n16631, n22753);
  not g36054 (n_16273, n22787);
  not g36055 (n_16274, n22788);
  and g36056 (n22789, n_16273, n_16274);
  and g36057 (n22790, n_11787, n22789);
  not g36058 (n_16275, n22789);
  and g36059 (n22791, pi0628, n_16275);
  and g36060 (n22792, n_11789, n22753);
  not g36061 (n_16276, n22792);
  and g36062 (n22793, pi1156, n_16276);
  not g36063 (n_16277, n22791);
  and g36064 (n22794, n_16277, n22793);
  and g36065 (n22795, pi0628, n22753);
  and g36066 (n22796, n_11789, n_16275);
  not g36067 (n_16278, n22795);
  and g36068 (n22797, n_11794, n_16278);
  not g36069 (n_16279, n22796);
  and g36070 (n22798, n_16279, n22797);
  not g36071 (n_16280, n22794);
  not g36072 (n_16281, n22798);
  and g36073 (n22799, n_16280, n_16281);
  not g36074 (n_16282, n22799);
  and g36075 (n22800, pi0792, n_16282);
  not g36076 (n_16283, n22790);
  not g36077 (n_16284, n22800);
  and g36078 (n22801, n_16283, n_16284);
  not g36079 (n_16285, n22801);
  and g36080 (n22802, n_11806, n_16285);
  and g36081 (n22803, pi0647, n_16245);
  not g36082 (n_16286, n22802);
  not g36083 (n_16287, n22803);
  and g36084 (n22804, n_16286, n_16287);
  and g36085 (n22805, n_11810, n22804);
  and g36086 (n22806, pi0647, n_16285);
  and g36087 (n22807, n_11806, n_16245);
  not g36088 (n_16288, n22806);
  not g36089 (n_16289, n22807);
  and g36090 (n22808, n_16288, n_16289);
  and g36091 (n22809, pi1157, n22808);
  not g36092 (n_16290, n22805);
  not g36093 (n_16291, n22809);
  and g36094 (n22810, n_16290, n_16291);
  not g36095 (n_16292, n22810);
  and g36096 (n22811, pi0787, n_16292);
  and g36097 (n22812, n_11803, n22801);
  not g36098 (n_16293, n22811);
  not g36099 (n_16294, n22812);
  and g36100 (n22813, n_16293, n_16294);
  not g36101 (n_16295, n22813);
  and g36102 (n22814, n_11819, n_16295);
  not g36103 (n_16296, n22814);
  and g36104 (n22815, pi0715, n_16296);
  and g36105 (n22816, pi0173, n_11417);
  and g36106 (n22817, pi0173, n_14476);
  and g36107 (n22818, n_9183, n_11739);
  not g36108 (n_16297, n22818);
  and g36109 (n22819, pi0745, n_16297);
  and g36110 (n22820, n_9183, n_15125);
  and g36111 (n22821, n17221, n22820);
  not g36112 (n_16298, n22817);
  not g36113 (n_16299, n22821);
  and g36114 (n22822, n_16298, n_16299);
  not g36115 (n_16300, n22819);
  and g36116 (n22823, n_16300, n22822);
  not g36117 (n_16301, n22823);
  and g36118 (n22824, n_161, n_16301);
  and g36119 (n22825, n_15125, n17280);
  and g36120 (n22826, pi0038, n_16247);
  not g36121 (n_16302, n22825);
  and g36122 (n22827, n_16302, n22826);
  not g36123 (n_16303, n22824);
  not g36124 (n_16304, n22827);
  and g36125 (n22828, n_16303, n_16304);
  not g36126 (n_16305, n22828);
  and g36127 (n22829, n2571, n_16305);
  not g36128 (n_16306, n22816);
  not g36129 (n_16307, n22829);
  and g36130 (n22830, n_16306, n_16307);
  not g36131 (n_16308, n22830);
  and g36132 (n22831, n_11960, n_16308);
  and g36133 (n22832, n17117, n_16245);
  not g36134 (n_16309, n22831);
  not g36135 (n_16310, n22832);
  and g36136 (n22833, n_16309, n_16310);
  not g36137 (n_16311, n22833);
  and g36138 (n22834, n_11964, n_16311);
  and g36139 (n22835, n_11967, n_16245);
  and g36140 (n22836, pi0609, n22831);
  not g36141 (n_16312, n22835);
  not g36142 (n_16313, n22836);
  and g36143 (n22837, n_16312, n_16313);
  not g36144 (n_16314, n22837);
  and g36145 (n22838, pi1155, n_16314);
  and g36146 (n22839, n_11972, n_16245);
  and g36147 (n22840, n_11971, n22831);
  not g36148 (n_16315, n22839);
  not g36149 (n_16316, n22840);
  and g36150 (n22841, n_16315, n_16316);
  not g36151 (n_16317, n22841);
  and g36152 (n22842, n_11768, n_16317);
  not g36153 (n_16318, n22838);
  not g36154 (n_16319, n22842);
  and g36155 (n22843, n_16318, n_16319);
  not g36156 (n_16320, n22843);
  and g36157 (n22844, pi0785, n_16320);
  not g36158 (n_16321, n22834);
  not g36159 (n_16322, n22844);
  and g36160 (n22845, n_16321, n_16322);
  not g36161 (n_16323, n22845);
  and g36162 (n22846, n_11981, n_16323);
  and g36163 (n22847, n_11984, n22753);
  and g36164 (n22848, pi0618, n22845);
  not g36165 (n_16324, n22847);
  and g36166 (n22849, pi1154, n_16324);
  not g36167 (n_16325, n22848);
  and g36168 (n22850, n_16325, n22849);
  and g36169 (n22851, n_11984, n22845);
  and g36170 (n22852, pi0618, n22753);
  not g36171 (n_16326, n22852);
  and g36172 (n22853, n_11413, n_16326);
  not g36173 (n_16327, n22851);
  and g36174 (n22854, n_16327, n22853);
  not g36175 (n_16328, n22850);
  not g36176 (n_16329, n22854);
  and g36177 (n22855, n_16328, n_16329);
  not g36178 (n_16330, n22855);
  and g36179 (n22856, pi0781, n_16330);
  not g36180 (n_16331, n22846);
  not g36181 (n_16332, n22856);
  and g36182 (n22857, n_16331, n_16332);
  not g36183 (n_16333, n22857);
  and g36184 (n22858, n_12315, n_16333);
  and g36185 (n22859, n_11821, n22753);
  and g36186 (n22860, pi0619, n22857);
  not g36187 (n_16334, n22859);
  and g36188 (n22861, pi1159, n_16334);
  not g36189 (n_16335, n22860);
  and g36190 (n22862, n_16335, n22861);
  and g36191 (n22863, n_11821, n22857);
  and g36192 (n22864, pi0619, n22753);
  not g36193 (n_16336, n22864);
  and g36194 (n22865, n_11405, n_16336);
  not g36195 (n_16337, n22863);
  and g36196 (n22866, n_16337, n22865);
  not g36197 (n_16338, n22862);
  not g36198 (n_16339, n22866);
  and g36199 (n22867, n_16338, n_16339);
  not g36200 (n_16340, n22867);
  and g36201 (n22868, pi0789, n_16340);
  not g36202 (n_16341, n22858);
  not g36203 (n_16342, n22868);
  and g36204 (n22869, n_16341, n_16342);
  not g36205 (n_16343, n22869);
  and g36206 (n22870, n_12318, n_16343);
  and g36207 (n22871, n_12320, n22753);
  and g36208 (n22872, pi0626, n22869);
  not g36209 (n_16344, n22871);
  and g36210 (n22873, pi1158, n_16344);
  not g36211 (n_16345, n22872);
  and g36212 (n22874, n_16345, n22873);
  and g36213 (n22875, n_12320, n22869);
  and g36214 (n22876, pi0626, n22753);
  not g36215 (n_16346, n22876);
  and g36216 (n22877, n_11397, n_16346);
  not g36217 (n_16347, n22875);
  and g36218 (n22878, n_16347, n22877);
  not g36219 (n_16348, n22874);
  not g36220 (n_16349, n22878);
  and g36221 (n22879, n_16348, n_16349);
  not g36222 (n_16350, n22879);
  and g36223 (n22880, pi0788, n_16350);
  not g36224 (n_16351, n22870);
  not g36225 (n_16352, n22880);
  and g36226 (n22881, n_16351, n_16352);
  and g36227 (n22882, n_12368, n22881);
  and g36228 (n22883, n17779, n22753);
  not g36229 (n_16353, n22882);
  not g36230 (n_16354, n22883);
  and g36231 (n22884, n_16353, n_16354);
  not g36232 (n_16355, n22884);
  and g36233 (n22885, n_12392, n_16355);
  and g36234 (n22886, n17804, n22753);
  not g36235 (n_16356, n22885);
  not g36236 (n_16357, n22886);
  and g36237 (n22887, n_16356, n_16357);
  not g36238 (n_16358, n22887);
  and g36239 (n22888, pi0644, n_16358);
  and g36240 (n22889, n_11819, n22753);
  not g36241 (n_16359, n22889);
  and g36242 (n22890, n_12395, n_16359);
  not g36243 (n_16360, n22888);
  and g36244 (n22891, n_16360, n22890);
  not g36245 (n_16361, n22891);
  and g36246 (n22892, pi1160, n_16361);
  not g36247 (n_16362, n22815);
  and g36248 (n22893, n_16362, n22892);
  and g36249 (n22894, pi0644, n_16295);
  not g36250 (n_16363, n22804);
  and g36251 (n22895, n17802, n_16363);
  and g36252 (n22896, n_14548, n22884);
  not g36253 (n_16364, n22808);
  and g36254 (n22897, n17801, n_16364);
  not g36255 (n_16365, n22895);
  not g36256 (n_16366, n22897);
  and g36257 (n22898, n_16365, n_16366);
  not g36258 (n_16367, n22896);
  and g36259 (n22899, n_16367, n22898);
  not g36260 (n_16368, n22899);
  and g36261 (n22900, pi0787, n_16368);
  and g36262 (n22901, n_12354, n22794);
  not g36263 (n_16369, n22881);
  and g36264 (n22902, n_14557, n_16369);
  and g36265 (n22903, pi0629, n22798);
  not g36266 (n_16370, n22901);
  not g36267 (n_16371, n22903);
  and g36268 (n22904, n_16370, n_16371);
  not g36269 (n_16372, n22902);
  and g36270 (n22905, n_16372, n22904);
  not g36271 (n_16373, n22905);
  and g36272 (n22906, pi0792, n_16373);
  and g36273 (n22907, pi0609, n22778);
  and g36274 (n22908, pi0173, n_12240);
  and g36275 (n22909, n_9183, n_12230);
  not g36276 (n_16374, n22908);
  and g36277 (n22910, pi0745, n_16374);
  not g36278 (n_16375, n22909);
  and g36279 (n22911, n_16375, n22910);
  and g36280 (n22912, n_9183, n17629);
  and g36281 (n22913, pi0173, n17631);
  not g36282 (n_16376, n22913);
  and g36283 (n22914, n_15125, n_16376);
  not g36284 (n_16377, n22912);
  and g36285 (n22915, n_16377, n22914);
  not g36286 (n_16378, n22911);
  not g36287 (n_16379, n22915);
  and g36288 (n22916, n_16378, n_16379);
  not g36289 (n_16380, n22916);
  and g36290 (n22917, n_162, n_16380);
  and g36291 (n22918, pi0173, n17605);
  and g36292 (n22919, n_9183, n_12180);
  not g36293 (n_16381, n22919);
  and g36294 (n22920, n_15125, n_16381);
  not g36295 (n_16382, n22918);
  and g36296 (n22921, n_16382, n22920);
  and g36297 (n22922, n_9183, n17404);
  and g36298 (n22923, pi0173, n17485);
  not g36299 (n_16383, n22923);
  and g36300 (n22924, pi0745, n_16383);
  not g36301 (n_16384, n22922);
  and g36302 (n22925, n_16384, n22924);
  not g36303 (n_16385, n22921);
  and g36304 (n22926, pi0039, n_16385);
  not g36305 (n_16386, n22925);
  and g36306 (n22927, n_16386, n22926);
  not g36307 (n_16387, n22917);
  and g36308 (n22928, n_161, n_16387);
  not g36309 (n_16388, n22927);
  and g36310 (n22929, n_16388, n22928);
  and g36311 (n22930, n_15125, n_12250);
  not g36312 (n_16389, n22930);
  and g36313 (n22931, n19471, n_16389);
  not g36314 (n_16390, n22931);
  and g36315 (n22932, n_9183, n_16390);
  and g36316 (n22933, n_15125, n17244);
  not g36317 (n_16391, n22933);
  and g36318 (n22934, n_12120, n_16391);
  not g36319 (n_16392, n22934);
  and g36320 (n22935, pi0173, n_16392);
  and g36321 (n22936, n6284, n22935);
  not g36322 (n_16393, n22936);
  and g36323 (n22937, pi0038, n_16393);
  not g36324 (n_16394, n22932);
  and g36325 (n22938, n_16394, n22937);
  not g36326 (n_16395, n22938);
  and g36327 (n22939, n_15127, n_16395);
  not g36328 (n_16396, n22929);
  and g36329 (n22940, n_16396, n22939);
  and g36330 (n22941, pi0723, n22828);
  not g36331 (n_16397, n22940);
  and g36332 (n22942, n2571, n_16397);
  not g36333 (n_16398, n22941);
  and g36334 (n22943, n_16398, n22942);
  not g36335 (n_16399, n22943);
  and g36336 (n22944, n_16306, n_16399);
  and g36337 (n22945, n_11753, n22944);
  and g36338 (n22946, pi0625, n22830);
  not g36339 (n_16400, n22946);
  and g36340 (n22947, n_11757, n_16400);
  not g36341 (n_16401, n22945);
  and g36342 (n22948, n_16401, n22947);
  and g36343 (n22949, n_11823, n_16261);
  not g36344 (n_16402, n22948);
  and g36345 (n22950, n_16402, n22949);
  and g36346 (n22951, n_11753, n22830);
  and g36347 (n22952, pi0625, n22944);
  not g36348 (n_16403, n22951);
  and g36349 (n22953, pi1153, n_16403);
  not g36350 (n_16404, n22952);
  and g36351 (n22954, n_16404, n22953);
  and g36352 (n22955, pi0608, n_16262);
  not g36353 (n_16405, n22954);
  and g36354 (n22956, n_16405, n22955);
  not g36355 (n_16406, n22950);
  not g36356 (n_16407, n22956);
  and g36357 (n22957, n_16406, n_16407);
  not g36358 (n_16408, n22957);
  and g36359 (n22958, pi0778, n_16408);
  and g36360 (n22959, n_11749, n22944);
  not g36361 (n_16409, n22958);
  not g36362 (n_16410, n22959);
  and g36363 (n22960, n_16409, n_16410);
  not g36364 (n_16411, n22960);
  and g36365 (n22961, n_11971, n_16411);
  not g36366 (n_16412, n22907);
  and g36367 (n22962, n_11768, n_16412);
  not g36368 (n_16413, n22961);
  and g36369 (n22963, n_16413, n22962);
  and g36370 (n22964, n_11767, n_16318);
  not g36371 (n_16414, n22963);
  and g36372 (n22965, n_16414, n22964);
  and g36373 (n22966, n_11971, n22778);
  and g36374 (n22967, pi0609, n_16411);
  not g36375 (n_16415, n22966);
  and g36376 (n22968, pi1155, n_16415);
  not g36377 (n_16416, n22967);
  and g36378 (n22969, n_16416, n22968);
  and g36379 (n22970, pi0660, n_16319);
  not g36380 (n_16417, n22969);
  and g36381 (n22971, n_16417, n22970);
  not g36382 (n_16418, n22965);
  not g36383 (n_16419, n22971);
  and g36384 (n22972, n_16418, n_16419);
  not g36385 (n_16420, n22972);
  and g36386 (n22973, pi0785, n_16420);
  and g36387 (n22974, n_11964, n_16411);
  not g36388 (n_16421, n22973);
  not g36389 (n_16422, n22974);
  and g36390 (n22975, n_16421, n_16422);
  not g36391 (n_16423, n22975);
  and g36392 (n22976, n_11984, n_16423);
  and g36393 (n22977, pi0618, n22781);
  not g36394 (n_16424, n22977);
  and g36395 (n22978, n_11413, n_16424);
  not g36396 (n_16425, n22976);
  and g36397 (n22979, n_16425, n22978);
  and g36398 (n22980, n_11412, n_16328);
  not g36399 (n_16426, n22979);
  and g36400 (n22981, n_16426, n22980);
  and g36401 (n22982, n_11984, n22781);
  and g36402 (n22983, pi0618, n_16423);
  not g36403 (n_16427, n22982);
  and g36404 (n22984, pi1154, n_16427);
  not g36405 (n_16428, n22983);
  and g36406 (n22985, n_16428, n22984);
  and g36407 (n22986, pi0627, n_16329);
  not g36408 (n_16429, n22985);
  and g36409 (n22987, n_16429, n22986);
  not g36410 (n_16430, n22981);
  not g36411 (n_16431, n22987);
  and g36412 (n22988, n_16430, n_16431);
  not g36413 (n_16432, n22988);
  and g36414 (n22989, pi0781, n_16432);
  and g36415 (n22990, n_11981, n_16423);
  not g36416 (n_16433, n22989);
  not g36417 (n_16434, n22990);
  and g36418 (n22991, n_16433, n_16434);
  and g36419 (n22992, n_12315, n22991);
  not g36420 (n_16435, n22784);
  and g36421 (n22993, pi0619, n_16435);
  not g36422 (n_16436, n22991);
  and g36423 (n22994, n_11821, n_16436);
  not g36424 (n_16437, n22993);
  and g36425 (n22995, n_11405, n_16437);
  not g36426 (n_16438, n22994);
  and g36427 (n22996, n_16438, n22995);
  and g36428 (n22997, n_11403, n_16338);
  not g36429 (n_16439, n22996);
  and g36430 (n22998, n_16439, n22997);
  and g36431 (n22999, pi0619, n_16436);
  and g36432 (n23000, n_11821, n_16435);
  not g36433 (n_16440, n23000);
  and g36434 (n23001, pi1159, n_16440);
  not g36435 (n_16441, n22999);
  and g36436 (n23002, n_16441, n23001);
  and g36437 (n23003, pi0648, n_16339);
  not g36438 (n_16442, n23002);
  and g36439 (n23004, n_16442, n23003);
  not g36440 (n_16443, n22998);
  and g36441 (n23005, pi0789, n_16443);
  not g36442 (n_16444, n23004);
  and g36443 (n23006, n_16444, n23005);
  not g36444 (n_16445, n22992);
  and g36445 (n23007, n17970, n_16445);
  not g36446 (n_16446, n23006);
  and g36447 (n23008, n_16446, n23007);
  and g36448 (n23009, n17871, n22786);
  and g36449 (n23010, n_11401, n22879);
  not g36450 (n_16447, n23009);
  not g36451 (n_16448, n23010);
  and g36452 (n23011, n_16447, n_16448);
  not g36453 (n_16449, n23011);
  and g36454 (n23012, pi0788, n_16449);
  not g36455 (n_16450, n23012);
  and g36456 (n23013, n_14638, n_16450);
  not g36457 (n_16451, n23008);
  and g36458 (n23014, n_16451, n23013);
  not g36459 (n_16452, n22906);
  not g36460 (n_16453, n23014);
  and g36461 (n23015, n_16452, n_16453);
  not g36462 (n_16454, n23015);
  and g36463 (n23016, n_14387, n_16454);
  not g36464 (n_16455, n22900);
  not g36465 (n_16456, n23016);
  and g36466 (n23017, n_16455, n_16456);
  and g36467 (n23018, n_11819, n23017);
  not g36468 (n_16457, n22894);
  and g36469 (n23019, n_12395, n_16457);
  not g36470 (n_16458, n23018);
  and g36471 (n23020, n_16458, n23019);
  and g36472 (n23021, pi0644, n22753);
  and g36473 (n23022, n_11819, n_16358);
  not g36474 (n_16459, n23021);
  and g36475 (n23023, pi0715, n_16459);
  not g36476 (n_16460, n23022);
  and g36477 (n23024, n_16460, n23023);
  not g36478 (n_16461, n23024);
  and g36479 (n23025, n_12405, n_16461);
  not g36480 (n_16462, n23020);
  and g36481 (n23026, n_16462, n23025);
  not g36482 (n_16463, n22893);
  not g36483 (n_16464, n23026);
  and g36484 (n23027, n_16463, n_16464);
  not g36485 (n_16465, n23027);
  and g36486 (n23028, pi0790, n_16465);
  and g36487 (n23029, pi0644, n22892);
  not g36488 (n_16466, n23029);
  and g36489 (n23030, pi0790, n_16466);
  not g36490 (n_16467, n23030);
  and g36491 (n23031, n23017, n_16467);
  not g36492 (n_16468, n23028);
  not g36493 (n_16469, n23031);
  and g36494 (n23032, n_16468, n_16469);
  not g36495 (n_16470, n23032);
  and g36496 (n23033, n_4226, n_16470);
  not g36497 (n_16471, n22752);
  and g36498 (n23034, n_12415, n_16471);
  not g36499 (n_16472, n23033);
  and g36500 (n23035, n_16472, n23034);
  and g36501 (n23036, n_9183, n_12418);
  and g36502 (n23037, n_15127, n16645);
  not g36503 (n_16473, n23036);
  not g36504 (n_16474, n23037);
  and g36505 (n23038, n_16473, n_16474);
  not g36506 (n_16475, n23038);
  and g36507 (n23039, n_11749, n_16475);
  and g36508 (n23040, n_11753, n23037);
  not g36509 (n_16476, n23040);
  and g36510 (n23041, n_16475, n_16476);
  not g36511 (n_16477, n23041);
  and g36512 (n23042, pi1153, n_16477);
  and g36513 (n23043, n_11757, n_16473);
  and g36514 (n23044, n_16476, n23043);
  not g36515 (n_16478, n23044);
  and g36516 (n23045, pi0778, n_16478);
  not g36517 (n_16479, n23042);
  and g36518 (n23046, n_16479, n23045);
  not g36519 (n_16480, n23039);
  not g36520 (n_16481, n23046);
  and g36521 (n23047, n_16480, n_16481);
  not g36522 (n_16482, n23047);
  and g36523 (n23048, n_12429, n_16482);
  and g36524 (n23049, n_12430, n23048);
  and g36525 (n23050, n_12431, n23049);
  and g36526 (n23051, n_12432, n23050);
  and g36527 (n23052, n_12436, n23051);
  and g36528 (n23053, n_11806, n23052);
  and g36529 (n23054, pi0647, n23036);
  not g36530 (n_16483, n23054);
  and g36531 (n23055, n_11810, n_16483);
  not g36532 (n_16484, n23053);
  and g36533 (n23056, n_16484, n23055);
  and g36534 (n23057, pi0630, n23056);
  and g36535 (n23058, n_16391, n_16473);
  not g36536 (n_16485, n23058);
  and g36537 (n23059, n_12448, n_16485);
  not g36538 (n_16486, n23059);
  and g36539 (n23060, n_11964, n_16486);
  and g36540 (n23061, n17296, n22933);
  not g36541 (n_16487, n23061);
  and g36542 (n23062, n23059, n_16487);
  not g36543 (n_16488, n23062);
  and g36544 (n23063, pi1155, n_16488);
  and g36545 (n23064, n_11768, n_16473);
  and g36546 (n23065, n_16487, n23064);
  not g36547 (n_16489, n23063);
  not g36548 (n_16490, n23065);
  and g36549 (n23066, n_16489, n_16490);
  not g36550 (n_16491, n23066);
  and g36551 (n23067, pi0785, n_16491);
  not g36552 (n_16492, n23060);
  not g36553 (n_16493, n23067);
  and g36554 (n23068, n_16492, n_16493);
  not g36555 (n_16494, n23068);
  and g36556 (n23069, n_11981, n_16494);
  and g36557 (n23070, n_12461, n23068);
  not g36558 (n_16495, n23070);
  and g36559 (n23071, pi1154, n_16495);
  and g36560 (n23072, n_12463, n23068);
  not g36561 (n_16496, n23072);
  and g36562 (n23073, n_11413, n_16496);
  not g36563 (n_16497, n23071);
  not g36564 (n_16498, n23073);
  and g36565 (n23074, n_16497, n_16498);
  not g36566 (n_16499, n23074);
  and g36567 (n23075, pi0781, n_16499);
  not g36568 (n_16500, n23069);
  not g36569 (n_16501, n23075);
  and g36570 (n23076, n_16500, n_16501);
  not g36571 (n_16502, n23076);
  and g36572 (n23077, n_12315, n_16502);
  and g36573 (n23078, n_11821, n2926);
  not g36574 (n_16503, n23078);
  and g36575 (n23079, n23076, n_16503);
  not g36576 (n_16504, n23079);
  and g36577 (n23080, pi1159, n_16504);
  and g36578 (n23081, pi0619, n2926);
  not g36579 (n_16505, n23081);
  and g36580 (n23082, n23076, n_16505);
  not g36581 (n_16506, n23082);
  and g36582 (n23083, n_11405, n_16506);
  not g36583 (n_16507, n23080);
  not g36584 (n_16508, n23083);
  and g36585 (n23084, n_16507, n_16508);
  not g36586 (n_16509, n23084);
  and g36587 (n23085, pi0789, n_16509);
  not g36588 (n_16510, n23077);
  not g36589 (n_16511, n23085);
  and g36590 (n23086, n_16510, n_16511);
  not g36591 (n_16512, n23086);
  and g36592 (n23087, n_12318, n_16512);
  and g36593 (n23088, n_12320, n23036);
  and g36594 (n23089, pi0626, n23086);
  not g36595 (n_16513, n23088);
  and g36596 (n23090, pi1158, n_16513);
  not g36597 (n_16514, n23089);
  and g36598 (n23091, n_16514, n23090);
  and g36599 (n23092, n_12320, n23086);
  and g36600 (n23093, pi0626, n23036);
  not g36601 (n_16515, n23093);
  and g36602 (n23094, n_11397, n_16515);
  not g36603 (n_16516, n23092);
  and g36604 (n23095, n_16516, n23094);
  not g36605 (n_16517, n23091);
  not g36606 (n_16518, n23095);
  and g36607 (n23096, n_16517, n_16518);
  not g36608 (n_16519, n23096);
  and g36609 (n23097, pi0788, n_16519);
  not g36610 (n_16520, n23087);
  not g36611 (n_16521, n23097);
  and g36612 (n23098, n_16520, n_16521);
  and g36613 (n23099, n_12368, n23098);
  and g36614 (n23100, n17779, n23036);
  not g36615 (n_16522, n23099);
  not g36616 (n_16523, n23100);
  and g36617 (n23101, n_16522, n_16523);
  and g36618 (n23102, n_14548, n23101);
  not g36619 (n_16524, n23052);
  and g36620 (n23103, pi0647, n_16524);
  and g36621 (n23104, n_11806, n_16473);
  not g36622 (n_16525, n23103);
  not g36623 (n_16526, n23104);
  and g36624 (n23105, n_16525, n_16526);
  not g36625 (n_16527, n23105);
  and g36626 (n23106, n17801, n_16527);
  not g36627 (n_16528, n23057);
  not g36628 (n_16529, n23106);
  and g36629 (n23107, n_16528, n_16529);
  not g36630 (n_16530, n23102);
  and g36631 (n23108, n_16530, n23107);
  not g36632 (n_16531, n23108);
  and g36633 (n23109, pi0787, n_16531);
  and g36634 (n23110, n17871, n23050);
  and g36635 (n23111, n_11401, n23096);
  not g36636 (n_16532, n23110);
  not g36637 (n_16533, n23111);
  and g36638 (n23112, n_16532, n_16533);
  not g36639 (n_16534, n23112);
  and g36640 (n23113, pi0788, n_16534);
  and g36641 (n23114, pi0618, n23048);
  and g36642 (n23115, n_11866, n_16475);
  and g36643 (n23116, pi0625, n23115);
  not g36644 (n_16535, n23115);
  and g36645 (n23117, n23058, n_16535);
  not g36646 (n_16536, n23116);
  not g36647 (n_16537, n23117);
  and g36648 (n23118, n_16536, n_16537);
  not g36649 (n_16538, n23118);
  and g36650 (n23119, n23043, n_16538);
  and g36651 (n23120, n_11823, n_16479);
  not g36652 (n_16539, n23119);
  and g36653 (n23121, n_16539, n23120);
  and g36654 (n23122, pi1153, n23058);
  and g36655 (n23123, n_16536, n23122);
  and g36656 (n23124, pi0608, n_16478);
  not g36657 (n_16540, n23123);
  and g36658 (n23125, n_16540, n23124);
  not g36659 (n_16541, n23121);
  not g36660 (n_16542, n23125);
  and g36661 (n23126, n_16541, n_16542);
  not g36662 (n_16543, n23126);
  and g36663 (n23127, pi0778, n_16543);
  and g36664 (n23128, n_11749, n_16537);
  not g36665 (n_16544, n23127);
  not g36666 (n_16545, n23128);
  and g36667 (n23129, n_16544, n_16545);
  not g36668 (n_16546, n23129);
  and g36669 (n23130, n_11971, n_16546);
  and g36670 (n23131, pi0609, n_16482);
  not g36671 (n_16547, n23131);
  and g36672 (n23132, n_11768, n_16547);
  not g36673 (n_16548, n23130);
  and g36674 (n23133, n_16548, n23132);
  and g36675 (n23134, n_11767, n_16489);
  not g36676 (n_16549, n23133);
  and g36677 (n23135, n_16549, n23134);
  and g36678 (n23136, pi0609, n_16546);
  and g36679 (n23137, n_11971, n_16482);
  not g36680 (n_16550, n23137);
  and g36681 (n23138, pi1155, n_16550);
  not g36682 (n_16551, n23136);
  and g36683 (n23139, n_16551, n23138);
  and g36684 (n23140, pi0660, n_16490);
  not g36685 (n_16552, n23139);
  and g36686 (n23141, n_16552, n23140);
  not g36687 (n_16553, n23135);
  not g36688 (n_16554, n23141);
  and g36689 (n23142, n_16553, n_16554);
  not g36690 (n_16555, n23142);
  and g36691 (n23143, pi0785, n_16555);
  and g36692 (n23144, n_11964, n_16546);
  not g36693 (n_16556, n23143);
  not g36694 (n_16557, n23144);
  and g36695 (n23145, n_16556, n_16557);
  not g36696 (n_16558, n23145);
  and g36697 (n23146, n_11984, n_16558);
  not g36698 (n_16559, n23114);
  and g36699 (n23147, n_11413, n_16559);
  not g36700 (n_16560, n23146);
  and g36701 (n23148, n_16560, n23147);
  and g36702 (n23149, n_11412, n_16497);
  not g36703 (n_16561, n23148);
  and g36704 (n23150, n_16561, n23149);
  and g36705 (n23151, n_11984, n23048);
  and g36706 (n23152, pi0618, n_16558);
  not g36707 (n_16562, n23151);
  and g36708 (n23153, pi1154, n_16562);
  not g36709 (n_16563, n23152);
  and g36710 (n23154, n_16563, n23153);
  and g36711 (n23155, pi0627, n_16498);
  not g36712 (n_16564, n23154);
  and g36713 (n23156, n_16564, n23155);
  not g36714 (n_16565, n23150);
  not g36715 (n_16566, n23156);
  and g36716 (n23157, n_16565, n_16566);
  not g36717 (n_16567, n23157);
  and g36718 (n23158, pi0781, n_16567);
  and g36719 (n23159, n_11981, n_16558);
  not g36720 (n_16568, n23158);
  not g36721 (n_16569, n23159);
  and g36722 (n23160, n_16568, n_16569);
  and g36723 (n23161, n_12315, n23160);
  not g36724 (n_16570, n23160);
  and g36725 (n23162, n_11821, n_16570);
  and g36726 (n23163, pi0619, n23049);
  not g36727 (n_16571, n23163);
  and g36728 (n23164, n_11405, n_16571);
  not g36729 (n_16572, n23162);
  and g36730 (n23165, n_16572, n23164);
  and g36731 (n23166, n_11403, n_16507);
  not g36732 (n_16573, n23165);
  and g36733 (n23167, n_16573, n23166);
  and g36734 (n23168, n_11821, n23049);
  and g36735 (n23169, pi0619, n_16570);
  not g36736 (n_16574, n23168);
  and g36737 (n23170, pi1159, n_16574);
  not g36738 (n_16575, n23169);
  and g36739 (n23171, n_16575, n23170);
  and g36740 (n23172, pi0648, n_16508);
  not g36741 (n_16576, n23171);
  and g36742 (n23173, n_16576, n23172);
  not g36743 (n_16577, n23167);
  and g36744 (n23174, pi0789, n_16577);
  not g36745 (n_16578, n23173);
  and g36746 (n23175, n_16578, n23174);
  not g36747 (n_16579, n23161);
  and g36748 (n23176, n17970, n_16579);
  not g36749 (n_16580, n23175);
  and g36750 (n23177, n_16580, n23176);
  not g36751 (n_16581, n23113);
  not g36752 (n_16582, n23177);
  and g36753 (n23178, n_16581, n_16582);
  not g36754 (n_16583, n23178);
  and g36755 (n23179, n_14638, n_16583);
  and g36756 (n23180, n17854, n23098);
  and g36757 (n23181, n20851, n23051);
  not g36758 (n_16584, n23180);
  not g36759 (n_16585, n23181);
  and g36760 (n23182, n_16584, n_16585);
  not g36761 (n_16586, n23182);
  and g36762 (n23183, n_12354, n_16586);
  and g36763 (n23184, n20855, n23051);
  and g36764 (n23185, n17853, n23098);
  not g36765 (n_16587, n23184);
  not g36766 (n_16588, n23185);
  and g36767 (n23186, n_16587, n_16588);
  not g36768 (n_16589, n23186);
  and g36769 (n23187, pi0629, n_16589);
  not g36770 (n_16590, n23183);
  not g36771 (n_16591, n23187);
  and g36772 (n23188, n_16590, n_16591);
  not g36773 (n_16592, n23188);
  and g36774 (n23189, pi0792, n_16592);
  not g36775 (n_16593, n23189);
  and g36776 (n23190, n_14387, n_16593);
  not g36777 (n_16594, n23179);
  and g36778 (n23191, n_16594, n23190);
  not g36779 (n_16595, n23109);
  not g36780 (n_16596, n23191);
  and g36781 (n23192, n_16595, n_16596);
  and g36782 (n23193, n_12411, n23192);
  and g36783 (n23194, n_11803, n_16524);
  and g36784 (n23195, pi1157, n_16527);
  not g36785 (n_16597, n23056);
  not g36786 (n_16598, n23195);
  and g36787 (n23196, n_16597, n_16598);
  not g36788 (n_16599, n23196);
  and g36789 (n23197, pi0787, n_16599);
  not g36790 (n_16600, n23194);
  not g36791 (n_16601, n23197);
  and g36792 (n23198, n_16600, n_16601);
  and g36793 (n23199, n_11819, n23198);
  and g36794 (n23200, pi0644, n23192);
  not g36795 (n_16602, n23199);
  and g36796 (n23201, pi0715, n_16602);
  not g36797 (n_16603, n23200);
  and g36798 (n23202, n_16603, n23201);
  not g36799 (n_16604, n23101);
  and g36800 (n23203, n_12392, n_16604);
  and g36801 (n23204, n17804, n23036);
  not g36802 (n_16605, n23203);
  not g36803 (n_16606, n23204);
  and g36804 (n23205, n_16605, n_16606);
  not g36805 (n_16607, n23205);
  and g36806 (n23206, pi0644, n_16607);
  and g36807 (n23207, n_11819, n23036);
  not g36808 (n_16608, n23207);
  and g36809 (n23208, n_12395, n_16608);
  not g36810 (n_16609, n23206);
  and g36811 (n23209, n_16609, n23208);
  not g36812 (n_16610, n23209);
  and g36813 (n23210, pi1160, n_16610);
  not g36814 (n_16611, n23202);
  and g36815 (n23211, n_16611, n23210);
  and g36816 (n23212, n_11819, n_16607);
  and g36817 (n23213, pi0644, n23036);
  not g36818 (n_16612, n23213);
  and g36819 (n23214, pi0715, n_16612);
  not g36820 (n_16613, n23212);
  and g36821 (n23215, n_16613, n23214);
  and g36822 (n23216, pi0644, n23198);
  and g36823 (n23217, n_11819, n23192);
  not g36824 (n_16614, n23216);
  and g36825 (n23218, n_12395, n_16614);
  not g36826 (n_16615, n23217);
  and g36827 (n23219, n_16615, n23218);
  not g36828 (n_16616, n23215);
  and g36829 (n23220, n_12405, n_16616);
  not g36830 (n_16617, n23219);
  and g36831 (n23221, n_16617, n23220);
  not g36832 (n_16618, n23211);
  not g36833 (n_16619, n23221);
  and g36834 (n23222, n_16618, n_16619);
  not g36835 (n_16620, n23222);
  and g36836 (n23223, pi0790, n_16620);
  not g36837 (n_16621, n23193);
  and g36838 (n23224, pi0832, n_16621);
  not g36839 (n_16622, n23223);
  and g36840 (n23225, n_16622, n23224);
  not g36841 (n_16623, n23035);
  not g36842 (n_16624, n23225);
  and g36843 (po0330, n_16623, n_16624);
  and g36844 (n23227, pi0174, n_11751);
  not g36845 (n_16625, n23227);
  and g36846 (n23228, n16635, n_16625);
  and g36847 (n23229, n17075, n_16625);
  and g36848 (n23230, pi0696, n2571);
  not g36849 (n_16626, n23230);
  and g36850 (n23231, n_16625, n_16626);
  and g36851 (n23232, n_299, n_11418);
  not g36852 (n_16627, n23232);
  and g36853 (n23233, n19899, n_16627);
  and g36854 (n23234, n_299, n18076);
  and g36855 (n23235, pi0174, n_14037);
  not g36856 (n_16628, n23234);
  and g36857 (n23236, n_161, n_16628);
  not g36858 (n_16629, n23235);
  and g36859 (n23237, n_16629, n23236);
  not g36860 (n_16630, n23233);
  and g36861 (n23238, n23230, n_16630);
  not g36862 (n_16631, n23237);
  and g36863 (n23239, n_16631, n23238);
  not g36864 (n_16632, n23231);
  not g36865 (n_16633, n23239);
  and g36866 (n23240, n_16632, n_16633);
  and g36867 (n23241, n_11749, n23240);
  and g36868 (n23242, n_11753, n_16625);
  not g36869 (n_16634, n23240);
  and g36870 (n23243, pi0625, n_16634);
  not g36871 (n_16635, n23242);
  and g36872 (n23244, pi1153, n_16635);
  not g36873 (n_16636, n23243);
  and g36874 (n23245, n_16636, n23244);
  and g36875 (n23246, n_11753, n_16634);
  and g36876 (n23247, pi0625, n_16625);
  not g36877 (n_16637, n23247);
  and g36878 (n23248, n_11757, n_16637);
  not g36879 (n_16638, n23246);
  and g36880 (n23249, n_16638, n23248);
  not g36881 (n_16639, n23245);
  not g36882 (n_16640, n23249);
  and g36883 (n23250, n_16639, n_16640);
  not g36884 (n_16641, n23250);
  and g36885 (n23251, pi0778, n_16641);
  not g36886 (n_16642, n23241);
  not g36887 (n_16643, n23251);
  and g36888 (n23252, n_16642, n_16643);
  and g36889 (n23253, n_11773, n23252);
  not g36890 (n_16644, n23229);
  not g36891 (n_16645, n23253);
  and g36892 (n23254, n_16644, n_16645);
  and g36893 (n23255, n_11777, n23254);
  and g36894 (n23256, n16639, n23227);
  not g36895 (n_16646, n23255);
  not g36896 (n_16647, n23256);
  and g36897 (n23257, n_16646, n_16647);
  and g36898 (n23258, n_11780, n23257);
  not g36899 (n_16648, n23228);
  not g36900 (n_16649, n23258);
  and g36901 (n23259, n_16648, n_16649);
  and g36902 (n23260, n_11783, n23259);
  and g36903 (n23261, n16631, n23227);
  not g36904 (n_16650, n23260);
  not g36905 (n_16651, n23261);
  and g36906 (n23262, n_16650, n_16651);
  not g36907 (n_16652, n23262);
  and g36908 (n23263, n_11787, n_16652);
  and g36909 (n23264, n_11789, n_16625);
  and g36910 (n23265, pi0628, n23262);
  not g36911 (n_16653, n23264);
  and g36912 (n23266, pi1156, n_16653);
  not g36913 (n_16654, n23265);
  and g36914 (n23267, n_16654, n23266);
  and g36915 (n23268, pi0628, n_16625);
  and g36916 (n23269, n_11789, n23262);
  not g36917 (n_16655, n23268);
  and g36918 (n23270, n_11794, n_16655);
  not g36919 (n_16656, n23269);
  and g36920 (n23271, n_16656, n23270);
  not g36921 (n_16657, n23267);
  not g36922 (n_16658, n23271);
  and g36923 (n23272, n_16657, n_16658);
  not g36924 (n_16659, n23272);
  and g36925 (n23273, pi0792, n_16659);
  not g36926 (n_16660, n23263);
  not g36927 (n_16661, n23273);
  and g36928 (n23274, n_16660, n_16661);
  not g36929 (n_16662, n23274);
  and g36930 (n23275, n_11803, n_16662);
  and g36931 (n23276, n_11806, n_16625);
  and g36932 (n23277, pi0647, n23274);
  not g36933 (n_16663, n23276);
  and g36934 (n23278, pi1157, n_16663);
  not g36935 (n_16664, n23277);
  and g36936 (n23279, n_16664, n23278);
  and g36937 (n23280, pi0647, n_16625);
  and g36938 (n23281, n_11806, n23274);
  not g36939 (n_16665, n23280);
  and g36940 (n23282, n_11810, n_16665);
  not g36941 (n_16666, n23281);
  and g36942 (n23283, n_16666, n23282);
  not g36943 (n_16667, n23279);
  not g36944 (n_16668, n23283);
  and g36945 (n23284, n_16667, n_16668);
  not g36946 (n_16669, n23284);
  and g36947 (n23285, pi0787, n_16669);
  not g36948 (n_16670, n23275);
  not g36949 (n_16671, n23285);
  and g36950 (n23286, n_16670, n_16671);
  and g36951 (n23287, n_11819, n23286);
  and g36952 (n23288, n_11821, n_16625);
  and g36953 (n23289, n17117, n_16625);
  and g36954 (n23290, pi0174, n_11417);
  and g36955 (n23291, pi0759, n17219);
  not g36956 (n_16672, n21470);
  not g36957 (n_16673, n23291);
  and g36958 (n23292, n_16672, n_16673);
  not g36959 (n_16674, n23292);
  and g36960 (n23293, pi0039, n_16674);
  and g36961 (n23294, n_15215, n16958);
  and g36962 (n23295, pi0759, n17139);
  not g36963 (n_16675, n23294);
  and g36964 (n23296, n_162, n_16675);
  not g36965 (n_16676, n23295);
  and g36966 (n23297, n_16676, n23296);
  not g36967 (n_16677, n23293);
  not g36968 (n_16678, n23297);
  and g36969 (n23298, n_16677, n_16678);
  not g36970 (n_16679, n23298);
  and g36971 (n23299, pi0174, n_16679);
  and g36972 (n23300, n_299, pi0759);
  and g36973 (n23301, n17275, n23300);
  not g36974 (n_16680, n23299);
  not g36975 (n_16681, n23301);
  and g36976 (n23302, n_16680, n_16681);
  not g36977 (n_16682, n23302);
  and g36978 (n23303, n_161, n_16682);
  and g36979 (n23304, pi0759, n17168);
  not g36980 (n_16683, n23304);
  and g36981 (n23305, n16641, n_16683);
  and g36982 (n23306, pi0038, n_16627);
  not g36983 (n_16684, n23305);
  and g36984 (n23307, n_16684, n23306);
  not g36985 (n_16685, n23303);
  not g36986 (n_16686, n23307);
  and g36987 (n23308, n_16685, n_16686);
  not g36988 (n_16687, n23308);
  and g36989 (n23309, n2571, n_16687);
  not g36990 (n_16688, n23290);
  not g36991 (n_16689, n23309);
  and g36992 (n23310, n_16688, n_16689);
  and g36993 (n23311, n_11960, n23310);
  not g36994 (n_16690, n23289);
  not g36995 (n_16691, n23311);
  and g36996 (n23312, n_16690, n_16691);
  and g36997 (n23313, n_11964, n23312);
  and g36998 (n23314, n_11971, n_16625);
  not g36999 (n_16692, n23312);
  and g37000 (n23315, pi0609, n_16692);
  not g37001 (n_16693, n23314);
  and g37002 (n23316, pi1155, n_16693);
  not g37003 (n_16694, n23315);
  and g37004 (n23317, n_16694, n23316);
  and g37005 (n23318, n_11971, n_16692);
  and g37006 (n23319, pi0609, n_16625);
  not g37007 (n_16695, n23319);
  and g37008 (n23320, n_11768, n_16695);
  not g37009 (n_16696, n23318);
  and g37010 (n23321, n_16696, n23320);
  not g37011 (n_16697, n23317);
  not g37012 (n_16698, n23321);
  and g37013 (n23322, n_16697, n_16698);
  not g37014 (n_16699, n23322);
  and g37015 (n23323, pi0785, n_16699);
  not g37016 (n_16700, n23313);
  not g37017 (n_16701, n23323);
  and g37018 (n23324, n_16700, n_16701);
  not g37019 (n_16702, n23324);
  and g37020 (n23325, n_11981, n_16702);
  and g37021 (n23326, n_11984, n_16625);
  and g37022 (n23327, pi0618, n23324);
  not g37023 (n_16703, n23326);
  and g37024 (n23328, pi1154, n_16703);
  not g37025 (n_16704, n23327);
  and g37026 (n23329, n_16704, n23328);
  and g37027 (n23330, pi0618, n_16625);
  and g37028 (n23331, n_11984, n23324);
  not g37029 (n_16705, n23330);
  and g37030 (n23332, n_11413, n_16705);
  not g37031 (n_16706, n23331);
  and g37032 (n23333, n_16706, n23332);
  not g37033 (n_16707, n23329);
  not g37034 (n_16708, n23333);
  and g37035 (n23334, n_16707, n_16708);
  not g37036 (n_16709, n23334);
  and g37037 (n23335, pi0781, n_16709);
  not g37038 (n_16710, n23325);
  not g37039 (n_16711, n23335);
  and g37040 (n23336, n_16710, n_16711);
  and g37041 (n23337, pi0619, n23336);
  not g37042 (n_16712, n23288);
  and g37043 (n23338, pi1159, n_16712);
  not g37044 (n_16713, n23337);
  and g37045 (n23339, n_16713, n23338);
  and g37046 (n23340, n_15254, n23308);
  and g37047 (n23341, n_299, n_13720);
  and g37048 (n23342, pi0174, n17546);
  not g37049 (n_16714, n23342);
  and g37050 (n23343, pi0759, n_16714);
  not g37051 (n_16715, n23341);
  and g37052 (n23344, n_16715, n23343);
  and g37053 (n23345, pi0174, n_13705);
  and g37054 (n23346, n_299, n_13702);
  not g37055 (n_16716, n23346);
  and g37056 (n23347, n_15215, n_16716);
  not g37057 (n_16717, n23345);
  and g37058 (n23348, n_16717, n23347);
  not g37059 (n_16718, n23344);
  and g37060 (n23349, pi0039, n_16718);
  not g37061 (n_16719, n23348);
  and g37062 (n23350, n_16719, n23349);
  and g37063 (n23351, n_299, n17631);
  and g37064 (n23352, pi0174, n17629);
  not g37065 (n_16720, n23351);
  and g37066 (n23353, pi0759, n_16720);
  not g37067 (n_16721, n23352);
  and g37068 (n23354, n_16721, n23353);
  and g37069 (n23355, n_299, n_12240);
  and g37070 (n23356, pi0174, n_12230);
  not g37071 (n_16722, n23355);
  and g37072 (n23357, n_15215, n_16722);
  not g37073 (n_16723, n23356);
  and g37074 (n23358, n_16723, n23357);
  not g37075 (n_16724, n23354);
  and g37076 (n23359, n_162, n_16724);
  not g37077 (n_16725, n23358);
  and g37078 (n23360, n_16725, n23359);
  not g37079 (n_16726, n23360);
  and g37080 (n23361, n_161, n_16726);
  not g37081 (n_16727, n23350);
  and g37082 (n23362, n_16727, n23361);
  not g37087 (n_16729, n23365);
  and g37088 (n23366, n2571, n_16729);
  not g37089 (n_16730, n23340);
  and g37090 (n23367, n_16730, n23366);
  not g37091 (n_16731, n23367);
  and g37092 (n23368, n_16688, n_16731);
  and g37093 (n23369, n_11753, n23368);
  and g37094 (n23370, pi0625, n23310);
  not g37095 (n_16732, n23370);
  and g37096 (n23371, n_11757, n_16732);
  not g37097 (n_16733, n23369);
  and g37098 (n23372, n_16733, n23371);
  and g37099 (n23373, n_11823, n_16639);
  not g37100 (n_16734, n23372);
  and g37101 (n23374, n_16734, n23373);
  and g37102 (n23375, n_11753, n23310);
  and g37103 (n23376, pi0625, n23368);
  not g37104 (n_16735, n23375);
  and g37105 (n23377, pi1153, n_16735);
  not g37106 (n_16736, n23376);
  and g37107 (n23378, n_16736, n23377);
  and g37108 (n23379, pi0608, n_16640);
  not g37109 (n_16737, n23378);
  and g37110 (n23380, n_16737, n23379);
  not g37111 (n_16738, n23374);
  not g37112 (n_16739, n23380);
  and g37113 (n23381, n_16738, n_16739);
  not g37114 (n_16740, n23381);
  and g37115 (n23382, pi0778, n_16740);
  and g37116 (n23383, n_11749, n23368);
  not g37117 (n_16741, n23382);
  not g37118 (n_16742, n23383);
  and g37119 (n23384, n_16741, n_16742);
  not g37120 (n_16743, n23384);
  and g37121 (n23385, n_11971, n_16743);
  and g37122 (n23386, pi0609, n23252);
  not g37123 (n_16744, n23386);
  and g37124 (n23387, n_11768, n_16744);
  not g37125 (n_16745, n23385);
  and g37126 (n23388, n_16745, n23387);
  and g37127 (n23389, n_11767, n_16697);
  not g37128 (n_16746, n23388);
  and g37129 (n23390, n_16746, n23389);
  and g37130 (n23391, n_11971, n23252);
  and g37131 (n23392, pi0609, n_16743);
  not g37132 (n_16747, n23391);
  and g37133 (n23393, pi1155, n_16747);
  not g37134 (n_16748, n23392);
  and g37135 (n23394, n_16748, n23393);
  and g37136 (n23395, pi0660, n_16698);
  not g37137 (n_16749, n23394);
  and g37138 (n23396, n_16749, n23395);
  not g37139 (n_16750, n23390);
  not g37140 (n_16751, n23396);
  and g37141 (n23397, n_16750, n_16751);
  not g37142 (n_16752, n23397);
  and g37143 (n23398, pi0785, n_16752);
  and g37144 (n23399, n_11964, n_16743);
  not g37145 (n_16753, n23398);
  not g37146 (n_16754, n23399);
  and g37147 (n23400, n_16753, n_16754);
  not g37148 (n_16755, n23400);
  and g37149 (n23401, n_11984, n_16755);
  not g37150 (n_16756, n23254);
  and g37151 (n23402, pi0618, n_16756);
  not g37152 (n_16757, n23402);
  and g37153 (n23403, n_11413, n_16757);
  not g37154 (n_16758, n23401);
  and g37155 (n23404, n_16758, n23403);
  and g37156 (n23405, n_11412, n_16707);
  not g37157 (n_16759, n23404);
  and g37158 (n23406, n_16759, n23405);
  and g37159 (n23407, pi0618, n_16755);
  and g37160 (n23408, n_11984, n_16756);
  not g37161 (n_16760, n23408);
  and g37162 (n23409, pi1154, n_16760);
  not g37163 (n_16761, n23407);
  and g37164 (n23410, n_16761, n23409);
  and g37165 (n23411, pi0627, n_16708);
  not g37166 (n_16762, n23410);
  and g37167 (n23412, n_16762, n23411);
  not g37168 (n_16763, n23406);
  not g37169 (n_16764, n23412);
  and g37170 (n23413, n_16763, n_16764);
  not g37171 (n_16765, n23413);
  and g37172 (n23414, pi0781, n_16765);
  and g37173 (n23415, n_11981, n_16755);
  not g37174 (n_16766, n23414);
  not g37175 (n_16767, n23415);
  and g37176 (n23416, n_16766, n_16767);
  not g37177 (n_16768, n23416);
  and g37178 (n23417, n_11821, n_16768);
  and g37179 (n23418, pi0619, n23257);
  not g37180 (n_16769, n23418);
  and g37181 (n23419, n_11405, n_16769);
  not g37182 (n_16770, n23417);
  and g37183 (n23420, n_16770, n23419);
  not g37184 (n_16771, n23339);
  and g37185 (n23421, n_11403, n_16771);
  not g37186 (n_16772, n23420);
  and g37187 (n23422, n_16772, n23421);
  and g37188 (n23423, pi0619, n_16625);
  and g37189 (n23424, n_11821, n23336);
  not g37190 (n_16773, n23423);
  and g37191 (n23425, n_11405, n_16773);
  not g37192 (n_16774, n23424);
  and g37193 (n23426, n_16774, n23425);
  and g37194 (n23427, n_11821, n23257);
  and g37195 (n23428, pi0619, n_16768);
  not g37196 (n_16775, n23427);
  and g37197 (n23429, pi1159, n_16775);
  not g37198 (n_16776, n23428);
  and g37199 (n23430, n_16776, n23429);
  not g37200 (n_16777, n23426);
  and g37201 (n23431, pi0648, n_16777);
  not g37202 (n_16778, n23430);
  and g37203 (n23432, n_16778, n23431);
  not g37204 (n_16779, n23422);
  not g37205 (n_16780, n23432);
  and g37206 (n23433, n_16779, n_16780);
  not g37207 (n_16781, n23433);
  and g37208 (n23434, pi0789, n_16781);
  and g37209 (n23435, n_12315, n_16768);
  not g37210 (n_16782, n23434);
  not g37211 (n_16783, n23435);
  and g37212 (n23436, n_16782, n_16783);
  and g37213 (n23437, n_12318, n23436);
  and g37214 (n23438, n_12320, n23436);
  and g37215 (n23439, pi0626, n23259);
  not g37216 (n_16784, n23439);
  and g37217 (n23440, n_11395, n_16784);
  not g37218 (n_16785, n23438);
  and g37219 (n23441, n_16785, n23440);
  not g37220 (n_16786, n23336);
  and g37221 (n23442, n_12315, n_16786);
  and g37222 (n23443, n_16771, n_16777);
  not g37223 (n_16787, n23443);
  and g37224 (n23444, pi0789, n_16787);
  not g37225 (n_16788, n23442);
  not g37226 (n_16789, n23444);
  and g37227 (n23445, n_16788, n_16789);
  not g37228 (n_16790, n23445);
  and g37229 (n23446, n_12320, n_16790);
  and g37230 (n23447, pi0626, n23227);
  not g37231 (n_16791, n23447);
  and g37232 (n23448, pi0641, n_16791);
  not g37233 (n_16792, n23446);
  and g37234 (n23449, n_16792, n23448);
  not g37235 (n_16793, n23449);
  and g37236 (n23450, n_11397, n_16793);
  not g37237 (n_16794, n23441);
  and g37238 (n23451, n_16794, n23450);
  and g37239 (n23452, pi0626, n23436);
  and g37240 (n23453, n_12320, n23259);
  not g37241 (n_16795, n23453);
  and g37242 (n23454, pi0641, n_16795);
  not g37243 (n_16796, n23452);
  and g37244 (n23455, n_16796, n23454);
  and g37245 (n23456, pi0626, n_16790);
  and g37246 (n23457, n_12320, n23227);
  not g37247 (n_16797, n23457);
  and g37248 (n23458, n_11395, n_16797);
  not g37249 (n_16798, n23456);
  and g37250 (n23459, n_16798, n23458);
  not g37251 (n_16799, n23459);
  and g37252 (n23460, pi1158, n_16799);
  not g37253 (n_16800, n23455);
  and g37254 (n23461, n_16800, n23460);
  not g37255 (n_16801, n23451);
  not g37256 (n_16802, n23461);
  and g37257 (n23462, n_16801, n_16802);
  not g37258 (n_16803, n23462);
  and g37259 (n23463, pi0788, n_16803);
  not g37260 (n_16804, n23437);
  not g37261 (n_16805, n23463);
  and g37262 (n23464, n_16804, n_16805);
  and g37263 (n23465, n_11789, n23464);
  and g37264 (n23466, n_12524, n_16790);
  and g37265 (n23467, n17969, n23227);
  not g37266 (n_16806, n23466);
  not g37267 (n_16807, n23467);
  and g37268 (n23468, n_16806, n_16807);
  and g37269 (n23469, pi0628, n23468);
  not g37270 (n_16808, n23469);
  and g37271 (n23470, n_11794, n_16808);
  not g37272 (n_16809, n23465);
  and g37273 (n23471, n_16809, n23470);
  and g37274 (n23472, n_12354, n_16657);
  not g37275 (n_16810, n23471);
  and g37276 (n23473, n_16810, n23472);
  and g37277 (n23474, pi0628, n23464);
  and g37278 (n23475, n_11789, n23468);
  not g37279 (n_16811, n23475);
  and g37280 (n23476, pi1156, n_16811);
  not g37281 (n_16812, n23474);
  and g37282 (n23477, n_16812, n23476);
  and g37283 (n23478, pi0629, n_16658);
  not g37284 (n_16813, n23477);
  and g37285 (n23479, n_16813, n23478);
  not g37286 (n_16814, n23473);
  not g37287 (n_16815, n23479);
  and g37288 (n23480, n_16814, n_16815);
  not g37289 (n_16816, n23480);
  and g37290 (n23481, pi0792, n_16816);
  and g37291 (n23482, n_11787, n23464);
  not g37292 (n_16817, n23481);
  not g37293 (n_16818, n23482);
  and g37294 (n23483, n_16817, n_16818);
  not g37295 (n_16819, n23483);
  and g37296 (n23484, n_11806, n_16819);
  not g37297 (n_16820, n23468);
  and g37298 (n23485, n_12368, n_16820);
  and g37299 (n23486, n17779, n23227);
  not g37300 (n_16821, n23485);
  not g37301 (n_16822, n23486);
  and g37302 (n23487, n_16821, n_16822);
  and g37303 (n23488, pi0647, n23487);
  not g37304 (n_16823, n23488);
  and g37305 (n23489, n_11810, n_16823);
  not g37306 (n_16824, n23484);
  and g37307 (n23490, n_16824, n23489);
  and g37308 (n23491, n_12375, n_16667);
  not g37309 (n_16825, n23490);
  and g37310 (n23492, n_16825, n23491);
  and g37311 (n23493, pi0647, n_16819);
  and g37312 (n23494, n_11806, n23487);
  not g37313 (n_16826, n23494);
  and g37314 (n23495, pi1157, n_16826);
  not g37315 (n_16827, n23493);
  and g37316 (n23496, n_16827, n23495);
  and g37317 (n23497, pi0630, n_16668);
  not g37318 (n_16828, n23496);
  and g37319 (n23498, n_16828, n23497);
  not g37320 (n_16829, n23492);
  not g37321 (n_16830, n23498);
  and g37322 (n23499, n_16829, n_16830);
  not g37323 (n_16831, n23499);
  and g37324 (n23500, pi0787, n_16831);
  and g37325 (n23501, n_11803, n_16819);
  not g37326 (n_16832, n23500);
  not g37327 (n_16833, n23501);
  and g37328 (n23502, n_16832, n_16833);
  not g37329 (n_16834, n23502);
  and g37330 (n23503, pi0644, n_16834);
  not g37331 (n_16835, n23287);
  and g37332 (n23504, pi0715, n_16835);
  not g37333 (n_16836, n23503);
  and g37334 (n23505, n_16836, n23504);
  and g37335 (n23506, n17804, n_16625);
  and g37336 (n23507, n_12392, n23487);
  not g37337 (n_16837, n23506);
  not g37338 (n_16838, n23507);
  and g37339 (n23508, n_16837, n_16838);
  not g37340 (n_16839, n23508);
  and g37341 (n23509, pi0644, n_16839);
  and g37342 (n23510, n_11819, n_16625);
  not g37343 (n_16840, n23510);
  and g37344 (n23511, n_12395, n_16840);
  not g37345 (n_16841, n23509);
  and g37346 (n23512, n_16841, n23511);
  not g37347 (n_16842, n23512);
  and g37348 (n23513, pi1160, n_16842);
  not g37349 (n_16843, n23505);
  and g37350 (n23514, n_16843, n23513);
  and g37351 (n23515, n_11819, n_16834);
  and g37352 (n23516, pi0644, n23286);
  not g37353 (n_16844, n23516);
  and g37354 (n23517, n_12395, n_16844);
  not g37355 (n_16845, n23515);
  and g37356 (n23518, n_16845, n23517);
  and g37357 (n23519, n_11819, n_16839);
  and g37358 (n23520, pi0644, n_16625);
  not g37359 (n_16846, n23520);
  and g37360 (n23521, pi0715, n_16846);
  not g37361 (n_16847, n23519);
  and g37362 (n23522, n_16847, n23521);
  not g37363 (n_16848, n23522);
  and g37364 (n23523, n_12405, n_16848);
  not g37365 (n_16849, n23518);
  and g37366 (n23524, n_16849, n23523);
  not g37367 (n_16850, n23514);
  and g37368 (n23525, pi0790, n_16850);
  not g37369 (n_16851, n23524);
  and g37370 (n23526, n_16851, n23525);
  and g37371 (n23527, n_12411, n23502);
  not g37372 (n_16852, n23527);
  and g37373 (n23528, n6305, n_16852);
  not g37374 (n_16853, n23526);
  and g37375 (n23529, n_16853, n23528);
  and g37376 (n23530, n_299, n_3232);
  not g37377 (n_16854, n23530);
  and g37378 (n23531, n_796, n_16854);
  not g37379 (n_16855, n23529);
  and g37380 (n23532, n_16855, n23531);
  and g37381 (n23533, pi0057, pi0174);
  not g37382 (n_16856, n23533);
  and g37383 (n23534, n_12415, n_16856);
  not g37384 (n_16857, n23532);
  and g37385 (n23535, n_16857, n23534);
  and g37386 (n23536, pi0174, n_12418);
  and g37387 (n23537, pi0759, n17244);
  and g37388 (n23538, n17291, n23537);
  not g37389 (n_16858, n23536);
  and g37390 (n23539, pi1155, n_16858);
  not g37391 (n_16859, n23538);
  and g37392 (n23540, n_16859, n23539);
  and g37393 (n23541, pi0696, n16645);
  not g37394 (n_16860, n23541);
  and g37395 (n23542, n_16858, n_16860);
  and g37396 (n23543, n_11749, n23542);
  and g37397 (n23544, pi0625, n23541);
  not g37398 (n_16861, n23542);
  not g37399 (n_16862, n23544);
  and g37400 (n23545, n_16861, n_16862);
  not g37401 (n_16863, n23545);
  and g37402 (n23546, n_11757, n_16863);
  and g37403 (n23547, pi1153, n_16858);
  and g37404 (n23548, n_16862, n23547);
  not g37405 (n_16864, n23546);
  not g37406 (n_16865, n23548);
  and g37407 (n23549, n_16864, n_16865);
  not g37408 (n_16866, n23549);
  and g37409 (n23550, pi0778, n_16866);
  not g37410 (n_16867, n23543);
  not g37411 (n_16868, n23550);
  and g37412 (n23551, n_16867, n_16868);
  and g37413 (n23552, pi0609, n23551);
  not g37414 (n_16869, n23537);
  and g37415 (n23553, n_16858, n_16869);
  and g37416 (n23554, pi0696, n17469);
  not g37417 (n_16870, n23554);
  and g37418 (n23555, n23553, n_16870);
  and g37419 (n23556, pi0625, n23554);
  not g37420 (n_16871, n23555);
  not g37421 (n_16872, n23556);
  and g37422 (n23557, n_16871, n_16872);
  not g37423 (n_16873, n23557);
  and g37424 (n23558, n_11757, n_16873);
  and g37425 (n23559, n_11823, n_16865);
  not g37426 (n_16874, n23558);
  and g37427 (n23560, n_16874, n23559);
  and g37428 (n23561, pi1153, n23553);
  and g37429 (n23562, n_16872, n23561);
  and g37430 (n23563, pi0608, n_16864);
  not g37431 (n_16875, n23562);
  and g37432 (n23564, n_16875, n23563);
  not g37433 (n_16876, n23560);
  not g37434 (n_16877, n23564);
  and g37435 (n23565, n_16876, n_16877);
  not g37436 (n_16878, n23565);
  and g37437 (n23566, pi0778, n_16878);
  and g37438 (n23567, n_11749, n_16871);
  not g37439 (n_16879, n23566);
  not g37440 (n_16880, n23567);
  and g37441 (n23568, n_16879, n_16880);
  not g37442 (n_16881, n23568);
  and g37443 (n23569, n_11971, n_16881);
  not g37444 (n_16882, n23552);
  and g37445 (n23570, n_11768, n_16882);
  not g37446 (n_16883, n23569);
  and g37447 (n23571, n_16883, n23570);
  not g37448 (n_16884, n23540);
  and g37449 (n23572, n_11767, n_16884);
  not g37450 (n_16885, n23571);
  and g37451 (n23573, n_16885, n23572);
  and g37452 (n23574, n17296, n23537);
  and g37453 (n23575, n_11768, n_16858);
  not g37454 (n_16886, n23574);
  and g37455 (n23576, n_16886, n23575);
  and g37456 (n23577, n_11971, n23551);
  and g37457 (n23578, pi0609, n_16881);
  not g37458 (n_16887, n23577);
  and g37459 (n23579, pi1155, n_16887);
  not g37460 (n_16888, n23578);
  and g37461 (n23580, n_16888, n23579);
  not g37462 (n_16889, n23576);
  and g37463 (n23581, pi0660, n_16889);
  not g37464 (n_16890, n23580);
  and g37465 (n23582, n_16890, n23581);
  not g37466 (n_16891, n23573);
  not g37467 (n_16892, n23582);
  and g37468 (n23583, n_16891, n_16892);
  not g37469 (n_16893, n23583);
  and g37470 (n23584, pi0785, n_16893);
  and g37471 (n23585, n_11964, n_16881);
  not g37472 (n_16894, n23584);
  not g37473 (n_16895, n23585);
  and g37474 (n23586, n_16894, n_16895);
  not g37475 (n_16896, n23586);
  and g37476 (n23587, n_11981, n_16896);
  and g37477 (n23588, n_14288, n23537);
  and g37478 (n23589, n20270, n23588);
  and g37479 (n23590, pi1154, n_16858);
  not g37480 (n_16897, n23589);
  and g37481 (n23591, n_16897, n23590);
  and g37482 (n23592, n_11773, n23551);
  not g37483 (n_16898, n23592);
  and g37484 (n23593, n_16858, n_16898);
  not g37485 (n_16899, n23593);
  and g37486 (n23594, pi0618, n_16899);
  and g37487 (n23595, n_11984, n_16896);
  not g37488 (n_16900, n23594);
  and g37489 (n23596, n_11413, n_16900);
  not g37490 (n_16901, n23595);
  and g37491 (n23597, n_16901, n23596);
  not g37492 (n_16902, n23591);
  and g37493 (n23598, n_11412, n_16902);
  not g37494 (n_16903, n23597);
  and g37495 (n23599, n_16903, n23598);
  and g37496 (n23600, n20319, n23588);
  and g37497 (n23601, n_11413, n_16858);
  not g37498 (n_16904, n23600);
  and g37499 (n23602, n_16904, n23601);
  and g37500 (n23603, n_11984, n_16899);
  and g37501 (n23604, pi0618, n_16896);
  not g37502 (n_16905, n23603);
  and g37503 (n23605, pi1154, n_16905);
  not g37504 (n_16906, n23604);
  and g37505 (n23606, n_16906, n23605);
  not g37506 (n_16907, n23602);
  and g37507 (n23607, pi0627, n_16907);
  not g37508 (n_16908, n23606);
  and g37509 (n23608, n_16908, n23607);
  not g37510 (n_16909, n23599);
  not g37511 (n_16910, n23608);
  and g37512 (n23609, n_16909, n_16910);
  not g37513 (n_16911, n23609);
  and g37514 (n23610, pi0781, n_16911);
  and g37515 (n23611, pi0648, n20228);
  and g37516 (n23612, n_11403, n20229);
  not g37517 (n_16912, n23611);
  not g37518 (n_16913, n23612);
  and g37519 (n23613, n_16912, n_16913);
  and g37520 (n23614, n16634, n23613);
  not g37521 (n_16914, n23614);
  and g37522 (n23615, pi0789, n_16914);
  not g37523 (n_16915, n23587);
  not g37524 (n_16916, n23615);
  and g37525 (n23616, n_16915, n_16916);
  not g37526 (n_16917, n23610);
  and g37527 (n23617, n_16917, n23616);
  and g37528 (n23618, n_14295, n23588);
  and g37529 (n23619, n20345, n23618);
  not g37530 (n_16918, n23619);
  and g37531 (n23620, n16633, n_16918);
  and g37532 (n23621, n19150, n23551);
  not g37533 (n_16919, n23613);
  not g37534 (n_16920, n23621);
  and g37535 (n23622, n_16919, n_16920);
  and g37536 (n23623, n20335, n23618);
  not g37537 (n_16921, n23623);
  and g37538 (n23624, n16632, n_16921);
  not g37539 (n_16922, n23620);
  not g37540 (n_16923, n23624);
  and g37541 (n23625, n_16922, n_16923);
  not g37542 (n_16924, n23622);
  and g37543 (n23626, n_16924, n23625);
  and g37544 (n23627, pi0789, n_16858);
  not g37545 (n_16925, n23626);
  and g37546 (n23628, n_16925, n23627);
  not g37547 (n_16926, n23628);
  and g37548 (n23629, n17970, n_16926);
  not g37549 (n_16927, n23617);
  and g37550 (n23630, n_16927, n23629);
  and g37551 (n23631, n20237, n23588);
  and g37552 (n23632, n_12320, n23631);
  not g37553 (n_16928, n23632);
  and g37554 (n23633, n_16858, n_16928);
  not g37555 (n_16929, n23633);
  and g37556 (n23634, n_11397, n_16929);
  and g37557 (n23635, n_11780, n23621);
  not g37558 (n_16930, n23635);
  and g37559 (n23636, n_16858, n_16930);
  not g37560 (n_16931, n23636);
  and g37561 (n23637, n17865, n_16931);
  not g37562 (n_16932, n23634);
  and g37563 (n23638, pi0641, n_16932);
  not g37564 (n_16933, n23637);
  and g37565 (n23639, n_16933, n23638);
  and g37566 (n23640, n17866, n_16931);
  and g37567 (n23641, pi0626, n23631);
  not g37568 (n_16934, n23641);
  and g37569 (n23642, n_16858, n_16934);
  not g37570 (n_16935, n23642);
  and g37571 (n23643, pi1158, n_16935);
  not g37572 (n_16936, n23643);
  and g37573 (n23644, n_11395, n_16936);
  not g37574 (n_16937, n23640);
  and g37575 (n23645, n_16937, n23644);
  not g37576 (n_16938, n23639);
  and g37577 (n23646, pi0788, n_16938);
  not g37578 (n_16939, n23645);
  and g37579 (n23647, n_16939, n23646);
  not g37580 (n_16940, n23647);
  and g37581 (n23648, n_14638, n_16940);
  not g37582 (n_16941, n23630);
  and g37583 (n23649, n_16941, n23648);
  and g37584 (n23650, n_12524, n23631);
  and g37585 (n23651, n_12354, n23650);
  not g37586 (n_16942, n23651);
  and g37587 (n23652, pi0628, n_16942);
  and g37588 (n23653, n19151, n23551);
  not g37589 (n_16943, n23653);
  and g37590 (n23654, pi0629, n_16943);
  not g37591 (n_16944, n23652);
  not g37592 (n_16945, n23654);
  and g37593 (n23655, n_16944, n_16945);
  not g37594 (n_16946, n23655);
  and g37595 (n23656, n_11794, n_16946);
  not g37596 (n_16947, n23650);
  and g37597 (n23657, n_11789, n_16947);
  not g37598 (n_16948, n23657);
  and g37599 (n23658, pi0629, n_16948);
  and g37600 (n23659, pi0628, n23653);
  not g37601 (n_16949, n23658);
  and g37602 (n23660, pi1156, n_16949);
  not g37603 (n_16950, n23659);
  and g37604 (n23661, n_16950, n23660);
  not g37605 (n_16951, n23656);
  not g37606 (n_16952, n23661);
  and g37607 (n23662, n_16951, n_16952);
  and g37608 (n23663, pi0792, n_16858);
  not g37609 (n_16953, n23662);
  and g37610 (n23664, n_16953, n23663);
  not g37611 (n_16954, n23649);
  not g37612 (n_16955, n23664);
  and g37613 (n23665, n_16954, n_16955);
  not g37614 (n_16956, n23665);
  and g37615 (n23666, n_14387, n_16956);
  and g37616 (n23667, n_12368, n23650);
  and g37617 (n23668, n_12375, n23667);
  not g37618 (n_16957, n23668);
  and g37619 (n23669, pi0647, n_16957);
  and g37620 (n23670, n_13453, n23653);
  not g37621 (n_16958, n23670);
  and g37622 (n23671, pi0630, n_16958);
  not g37623 (n_16959, n23669);
  not g37624 (n_16960, n23671);
  and g37625 (n23672, n_16959, n_16960);
  not g37626 (n_16961, n23672);
  and g37627 (n23673, n_11810, n_16961);
  and g37628 (n23674, pi0630, n23667);
  and g37629 (n23675, n_12375, n_16958);
  not g37630 (n_16962, n23675);
  and g37631 (n23676, pi0647, n_16962);
  not g37632 (n_16963, n23674);
  and g37633 (n23677, pi1157, n_16963);
  not g37634 (n_16964, n23676);
  and g37635 (n23678, n_16964, n23677);
  not g37636 (n_16965, n23673);
  not g37637 (n_16966, n23678);
  and g37638 (n23679, n_16965, n_16966);
  and g37639 (n23680, pi0787, n_16858);
  not g37640 (n_16967, n23679);
  and g37641 (n23681, n_16967, n23680);
  not g37642 (n_16968, n23666);
  not g37643 (n_16969, n23681);
  and g37644 (n23682, n_16968, n_16969);
  and g37645 (n23683, n_12411, n23682);
  and g37646 (n23684, n_12368, n_12392);
  and g37647 (n23685, n23650, n23684);
  and g37648 (n23686, pi0644, n23685);
  and g37649 (n23687, n_12395, n_16858);
  not g37650 (n_16970, n23686);
  and g37651 (n23688, n_16970, n23687);
  and g37652 (n23689, n_13598, n23670);
  not g37653 (n_16971, n23689);
  and g37654 (n23690, n_16858, n_16971);
  not g37655 (n_16972, n23690);
  and g37656 (n23691, n_11819, n_16972);
  and g37657 (n23692, pi0644, n23682);
  not g37658 (n_16973, n23691);
  and g37659 (n23693, pi0715, n_16973);
  not g37660 (n_16974, n23692);
  and g37661 (n23694, n_16974, n23693);
  not g37662 (n_16975, n23688);
  and g37663 (n23695, pi1160, n_16975);
  not g37664 (n_16976, n23694);
  and g37665 (n23696, n_16976, n23695);
  and g37666 (n23697, n_11819, n23685);
  and g37667 (n23698, pi0715, n_16858);
  not g37668 (n_16977, n23697);
  and g37669 (n23699, n_16977, n23698);
  and g37670 (n23700, n_11819, n23682);
  and g37671 (n23701, pi0644, n_16972);
  not g37672 (n_16978, n23701);
  and g37673 (n23702, n_12395, n_16978);
  not g37674 (n_16979, n23700);
  and g37675 (n23703, n_16979, n23702);
  not g37676 (n_16980, n23699);
  and g37677 (n23704, n_12405, n_16980);
  not g37678 (n_16981, n23703);
  and g37679 (n23705, n_16981, n23704);
  not g37680 (n_16982, n23696);
  not g37681 (n_16983, n23705);
  and g37682 (n23706, n_16982, n_16983);
  not g37683 (n_16984, n23706);
  and g37684 (n23707, pi0790, n_16984);
  not g37685 (n_16985, n23683);
  and g37686 (n23708, pi0832, n_16985);
  not g37687 (n_16986, n23707);
  and g37688 (n23709, n_16986, n23708);
  not g37689 (n_16987, n23535);
  not g37690 (n_16988, n23709);
  and g37691 (po0331, n_16987, n_16988);
  and g37692 (n23711, n_7662, n_12418);
  and g37693 (n23712, pi0700, n16645);
  not g37694 (n_16989, n23711);
  not g37695 (n_16990, n23712);
  and g37696 (n23713, n_16989, n_16990);
  not g37697 (n_16991, n23713);
  and g37698 (n23714, n_11749, n_16991);
  and g37699 (n23715, n_11753, n23712);
  not g37700 (n_16992, n23715);
  and g37701 (n23716, n_16991, n_16992);
  not g37702 (n_16993, n23716);
  and g37703 (n23717, pi1153, n_16993);
  and g37704 (n23718, n_11757, n_16989);
  and g37705 (n23719, n_16992, n23718);
  not g37706 (n_16994, n23719);
  and g37707 (n23720, pi0778, n_16994);
  not g37708 (n_16995, n23717);
  and g37709 (n23721, n_16995, n23720);
  not g37710 (n_16996, n23714);
  not g37711 (n_16997, n23721);
  and g37712 (n23722, n_16996, n_16997);
  not g37713 (n_16998, n23722);
  and g37714 (n23723, n_12429, n_16998);
  and g37715 (n23724, n_12430, n23723);
  and g37716 (n23725, n_12431, n23724);
  and g37717 (n23726, n_12432, n23725);
  and g37718 (n23727, n_12436, n23726);
  and g37719 (n23728, n_11806, n23727);
  and g37720 (n23729, pi0647, n23711);
  not g37721 (n_16999, n23729);
  and g37722 (n23730, n_11810, n_16999);
  not g37723 (n_17000, n23728);
  and g37724 (n23731, n_17000, n23730);
  and g37725 (n23732, pi0630, n23731);
  and g37726 (n23733, pi0766, n17244);
  not g37727 (n_17001, n23733);
  and g37728 (n23734, n_16989, n_17001);
  not g37729 (n_17002, n23734);
  and g37730 (n23735, n_12448, n_17002);
  not g37731 (n_17003, n23735);
  and g37732 (n23736, n_11964, n_17003);
  and g37733 (n23737, n17296, n23733);
  not g37734 (n_17004, n23737);
  and g37735 (n23738, n23735, n_17004);
  not g37736 (n_17005, n23738);
  and g37737 (n23739, pi1155, n_17005);
  and g37738 (n23740, n_11768, n_16989);
  and g37739 (n23741, n_17004, n23740);
  not g37740 (n_17006, n23739);
  not g37741 (n_17007, n23741);
  and g37742 (n23742, n_17006, n_17007);
  not g37743 (n_17008, n23742);
  and g37744 (n23743, pi0785, n_17008);
  not g37745 (n_17009, n23736);
  not g37746 (n_17010, n23743);
  and g37747 (n23744, n_17009, n_17010);
  not g37748 (n_17011, n23744);
  and g37749 (n23745, n_11981, n_17011);
  and g37750 (n23746, n_12461, n23744);
  not g37751 (n_17012, n23746);
  and g37752 (n23747, pi1154, n_17012);
  and g37753 (n23748, n_12463, n23744);
  not g37754 (n_17013, n23748);
  and g37755 (n23749, n_11413, n_17013);
  not g37756 (n_17014, n23747);
  not g37757 (n_17015, n23749);
  and g37758 (n23750, n_17014, n_17015);
  not g37759 (n_17016, n23750);
  and g37760 (n23751, pi0781, n_17016);
  not g37761 (n_17017, n23745);
  not g37762 (n_17018, n23751);
  and g37763 (n23752, n_17017, n_17018);
  not g37764 (n_17019, n23752);
  and g37765 (n23753, n_12315, n_17019);
  and g37766 (n23754, n_16503, n23752);
  not g37767 (n_17020, n23754);
  and g37768 (n23755, pi1159, n_17020);
  and g37769 (n23756, n_16505, n23752);
  not g37770 (n_17021, n23756);
  and g37771 (n23757, n_11405, n_17021);
  not g37772 (n_17022, n23755);
  not g37773 (n_17023, n23757);
  and g37774 (n23758, n_17022, n_17023);
  not g37775 (n_17024, n23758);
  and g37776 (n23759, pi0789, n_17024);
  not g37777 (n_17025, n23753);
  not g37778 (n_17026, n23759);
  and g37779 (n23760, n_17025, n_17026);
  and g37780 (n23761, n_12524, n23760);
  and g37781 (n23762, n17969, n23711);
  not g37782 (n_17027, n23761);
  not g37783 (n_17028, n23762);
  and g37784 (n23763, n_17027, n_17028);
  not g37785 (n_17029, n23763);
  and g37786 (n23764, n_12368, n_17029);
  and g37787 (n23765, n17779, n23711);
  not g37788 (n_17030, n23764);
  not g37789 (n_17031, n23765);
  and g37790 (n23766, n_17030, n_17031);
  and g37791 (n23767, n_14548, n23766);
  not g37792 (n_17032, n23727);
  and g37793 (n23768, pi0647, n_17032);
  and g37794 (n23769, n_11806, n_16989);
  not g37795 (n_17033, n23768);
  not g37796 (n_17034, n23769);
  and g37797 (n23770, n_17033, n_17034);
  not g37798 (n_17035, n23770);
  and g37799 (n23771, n17801, n_17035);
  not g37800 (n_17036, n23732);
  not g37801 (n_17037, n23771);
  and g37802 (n23772, n_17036, n_17037);
  not g37803 (n_17038, n23767);
  and g37804 (n23773, n_17038, n23772);
  not g37805 (n_17039, n23773);
  and g37806 (n23774, pi0787, n_17039);
  and g37807 (n23775, n17871, n23725);
  not g37808 (n_17040, n23760);
  and g37809 (n23776, n_12320, n_17040);
  and g37810 (n23777, pi0626, n_16989);
  not g37811 (n_17041, n23777);
  and g37812 (n23778, n16629, n_17041);
  not g37813 (n_17042, n23776);
  and g37814 (n23779, n_17042, n23778);
  and g37815 (n23780, pi0626, n_17040);
  and g37816 (n23781, n_12320, n_16989);
  not g37817 (n_17043, n23781);
  and g37818 (n23782, n16628, n_17043);
  not g37819 (n_17044, n23780);
  and g37820 (n23783, n_17044, n23782);
  not g37821 (n_17045, n23775);
  not g37822 (n_17046, n23779);
  and g37823 (n23784, n_17045, n_17046);
  not g37824 (n_17047, n23783);
  and g37825 (n23785, n_17047, n23784);
  not g37826 (n_17048, n23785);
  and g37827 (n23786, pi0788, n_17048);
  and g37828 (n23787, pi0618, n23723);
  and g37829 (n23788, n_11866, n_16991);
  and g37830 (n23789, pi0625, n23788);
  not g37831 (n_17049, n23788);
  and g37832 (n23790, n23734, n_17049);
  not g37833 (n_17050, n23789);
  not g37834 (n_17051, n23790);
  and g37835 (n23791, n_17050, n_17051);
  not g37836 (n_17052, n23791);
  and g37837 (n23792, n23718, n_17052);
  and g37838 (n23793, n_11823, n_16995);
  not g37839 (n_17053, n23792);
  and g37840 (n23794, n_17053, n23793);
  and g37841 (n23795, pi1153, n23734);
  and g37842 (n23796, n_17050, n23795);
  and g37843 (n23797, pi0608, n_16994);
  not g37844 (n_17054, n23796);
  and g37845 (n23798, n_17054, n23797);
  not g37846 (n_17055, n23794);
  not g37847 (n_17056, n23798);
  and g37848 (n23799, n_17055, n_17056);
  not g37849 (n_17057, n23799);
  and g37850 (n23800, pi0778, n_17057);
  and g37851 (n23801, n_11749, n_17051);
  not g37852 (n_17058, n23800);
  not g37853 (n_17059, n23801);
  and g37854 (n23802, n_17058, n_17059);
  not g37855 (n_17060, n23802);
  and g37856 (n23803, n_11971, n_17060);
  and g37857 (n23804, pi0609, n_16998);
  not g37858 (n_17061, n23804);
  and g37859 (n23805, n_11768, n_17061);
  not g37860 (n_17062, n23803);
  and g37861 (n23806, n_17062, n23805);
  and g37862 (n23807, n_11767, n_17006);
  not g37863 (n_17063, n23806);
  and g37864 (n23808, n_17063, n23807);
  and g37865 (n23809, pi0609, n_17060);
  and g37866 (n23810, n_11971, n_16998);
  not g37867 (n_17064, n23810);
  and g37868 (n23811, pi1155, n_17064);
  not g37869 (n_17065, n23809);
  and g37870 (n23812, n_17065, n23811);
  and g37871 (n23813, pi0660, n_17007);
  not g37872 (n_17066, n23812);
  and g37873 (n23814, n_17066, n23813);
  not g37874 (n_17067, n23808);
  not g37875 (n_17068, n23814);
  and g37876 (n23815, n_17067, n_17068);
  not g37877 (n_17069, n23815);
  and g37878 (n23816, pi0785, n_17069);
  and g37879 (n23817, n_11964, n_17060);
  not g37880 (n_17070, n23816);
  not g37881 (n_17071, n23817);
  and g37882 (n23818, n_17070, n_17071);
  not g37883 (n_17072, n23818);
  and g37884 (n23819, n_11984, n_17072);
  not g37885 (n_17073, n23787);
  and g37886 (n23820, n_11413, n_17073);
  not g37887 (n_17074, n23819);
  and g37888 (n23821, n_17074, n23820);
  and g37889 (n23822, n_11412, n_17014);
  not g37890 (n_17075, n23821);
  and g37891 (n23823, n_17075, n23822);
  and g37892 (n23824, n_11984, n23723);
  and g37893 (n23825, pi0618, n_17072);
  not g37894 (n_17076, n23824);
  and g37895 (n23826, pi1154, n_17076);
  not g37896 (n_17077, n23825);
  and g37897 (n23827, n_17077, n23826);
  and g37898 (n23828, pi0627, n_17015);
  not g37899 (n_17078, n23827);
  and g37900 (n23829, n_17078, n23828);
  not g37901 (n_17079, n23823);
  not g37902 (n_17080, n23829);
  and g37903 (n23830, n_17079, n_17080);
  not g37904 (n_17081, n23830);
  and g37905 (n23831, pi0781, n_17081);
  and g37906 (n23832, n_11981, n_17072);
  not g37907 (n_17082, n23831);
  not g37908 (n_17083, n23832);
  and g37909 (n23833, n_17082, n_17083);
  and g37910 (n23834, n_12315, n23833);
  not g37911 (n_17084, n23833);
  and g37912 (n23835, n_11821, n_17084);
  and g37913 (n23836, pi0619, n23724);
  not g37914 (n_17085, n23836);
  and g37915 (n23837, n_11405, n_17085);
  not g37916 (n_17086, n23835);
  and g37917 (n23838, n_17086, n23837);
  and g37918 (n23839, n_11403, n_17022);
  not g37919 (n_17087, n23838);
  and g37920 (n23840, n_17087, n23839);
  and g37921 (n23841, pi0619, n_17084);
  and g37922 (n23842, n_11821, n23724);
  not g37923 (n_17088, n23842);
  and g37924 (n23843, pi1159, n_17088);
  not g37925 (n_17089, n23841);
  and g37926 (n23844, n_17089, n23843);
  and g37927 (n23845, pi0648, n_17023);
  not g37928 (n_17090, n23844);
  and g37929 (n23846, n_17090, n23845);
  not g37930 (n_17091, n23840);
  and g37931 (n23847, pi0789, n_17091);
  not g37932 (n_17092, n23846);
  and g37933 (n23848, n_17092, n23847);
  not g37934 (n_17093, n23834);
  and g37935 (n23849, n17970, n_17093);
  not g37936 (n_17094, n23848);
  and g37937 (n23850, n_17094, n23849);
  not g37938 (n_17095, n23786);
  not g37939 (n_17096, n23850);
  and g37940 (n23851, n_17095, n_17096);
  not g37941 (n_17097, n23851);
  and g37942 (n23852, n_14638, n_17097);
  and g37943 (n23853, n17854, n_17029);
  and g37944 (n23854, n20851, n23726);
  not g37945 (n_17098, n23853);
  not g37946 (n_17099, n23854);
  and g37947 (n23855, n_17098, n_17099);
  not g37948 (n_17100, n23855);
  and g37949 (n23856, n_12354, n_17100);
  and g37950 (n23857, n20855, n23726);
  and g37951 (n23858, n17853, n_17029);
  not g37952 (n_17101, n23857);
  not g37953 (n_17102, n23858);
  and g37954 (n23859, n_17101, n_17102);
  not g37955 (n_17103, n23859);
  and g37956 (n23860, pi0629, n_17103);
  not g37957 (n_17104, n23856);
  not g37958 (n_17105, n23860);
  and g37959 (n23861, n_17104, n_17105);
  not g37960 (n_17106, n23861);
  and g37961 (n23862, pi0792, n_17106);
  not g37962 (n_17107, n23862);
  and g37963 (n23863, n_14387, n_17107);
  not g37964 (n_17108, n23852);
  and g37965 (n23864, n_17108, n23863);
  not g37966 (n_17109, n23774);
  not g37967 (n_17110, n23864);
  and g37968 (n23865, n_17109, n_17110);
  and g37969 (n23866, n_12411, n23865);
  and g37970 (n23867, n_11803, n_17032);
  and g37971 (n23868, pi1157, n_17035);
  not g37972 (n_17111, n23731);
  not g37973 (n_17112, n23868);
  and g37974 (n23869, n_17111, n_17112);
  not g37975 (n_17113, n23869);
  and g37976 (n23870, pi0787, n_17113);
  not g37977 (n_17114, n23867);
  not g37978 (n_17115, n23870);
  and g37979 (n23871, n_17114, n_17115);
  and g37980 (n23872, n_11819, n23871);
  and g37981 (n23873, pi0644, n23865);
  not g37982 (n_17116, n23872);
  and g37983 (n23874, pi0715, n_17116);
  not g37984 (n_17117, n23873);
  and g37985 (n23875, n_17117, n23874);
  not g37986 (n_17118, n23766);
  and g37987 (n23876, n_12392, n_17118);
  and g37988 (n23877, n17804, n23711);
  not g37989 (n_17119, n23876);
  not g37990 (n_17120, n23877);
  and g37991 (n23878, n_17119, n_17120);
  not g37992 (n_17121, n23878);
  and g37993 (n23879, pi0644, n_17121);
  and g37994 (n23880, n_11819, n23711);
  not g37995 (n_17122, n23880);
  and g37996 (n23881, n_12395, n_17122);
  not g37997 (n_17123, n23879);
  and g37998 (n23882, n_17123, n23881);
  not g37999 (n_17124, n23882);
  and g38000 (n23883, pi1160, n_17124);
  not g38001 (n_17125, n23875);
  and g38002 (n23884, n_17125, n23883);
  and g38003 (n23885, n_11819, n_17121);
  and g38004 (n23886, pi0644, n23711);
  not g38005 (n_17126, n23886);
  and g38006 (n23887, pi0715, n_17126);
  not g38007 (n_17127, n23885);
  and g38008 (n23888, n_17127, n23887);
  and g38009 (n23889, pi0644, n23871);
  and g38010 (n23890, n_11819, n23865);
  not g38011 (n_17128, n23889);
  and g38012 (n23891, n_12395, n_17128);
  not g38013 (n_17129, n23890);
  and g38014 (n23892, n_17129, n23891);
  not g38015 (n_17130, n23888);
  and g38016 (n23893, n_12405, n_17130);
  not g38017 (n_17131, n23892);
  and g38018 (n23894, n_17131, n23893);
  not g38019 (n_17132, n23884);
  not g38020 (n_17133, n23894);
  and g38021 (n23895, n_17132, n_17133);
  not g38022 (n_17134, n23895);
  and g38023 (n23896, pi0790, n_17134);
  not g38024 (n_17135, n23866);
  and g38025 (n23897, pi0832, n_17135);
  not g38026 (n_17136, n23896);
  and g38027 (n23898, n_17136, n23897);
  and g38028 (n23899, n_7662, po1038);
  and g38029 (n23900, n_7662, n_11751);
  not g38030 (n_17137, n23900);
  and g38031 (n23901, n16635, n_17137);
  and g38032 (n23902, pi0175, n_11417);
  and g38033 (n23903, n_7662, n_11418);
  not g38034 (n_17138, n23903);
  and g38035 (n23904, n16647, n_17138);
  and g38036 (n23905, n_7662, n18072);
  and g38037 (n23906, pi0175, n_12608);
  not g38038 (n_17139, n23906);
  and g38039 (n23907, n_161, n_17139);
  not g38040 (n_17140, n23905);
  and g38041 (n23908, n_17140, n23907);
  not g38042 (n_17141, n23904);
  and g38043 (n23909, pi0700, n_17141);
  not g38044 (n_17142, n23908);
  and g38045 (n23910, n_17142, n23909);
  and g38046 (n23911, n_7662, n_15317);
  and g38047 (n23912, n_11743, n23911);
  not g38048 (n_17143, n23912);
  and g38049 (n23913, n2571, n_17143);
  not g38050 (n_17144, n23910);
  and g38051 (n23914, n_17144, n23913);
  not g38052 (n_17145, n23902);
  not g38053 (n_17146, n23914);
  and g38054 (n23915, n_17145, n_17146);
  not g38055 (n_17147, n23915);
  and g38056 (n23916, n_11749, n_17147);
  and g38057 (n23917, n_11753, n23900);
  and g38058 (n23918, pi0625, n23915);
  not g38059 (n_17148, n23917);
  and g38060 (n23919, pi1153, n_17148);
  not g38061 (n_17149, n23918);
  and g38062 (n23920, n_17149, n23919);
  and g38063 (n23921, n_11753, n23915);
  and g38064 (n23922, pi0625, n23900);
  not g38065 (n_17150, n23922);
  and g38066 (n23923, n_11757, n_17150);
  not g38067 (n_17151, n23921);
  and g38068 (n23924, n_17151, n23923);
  not g38069 (n_17152, n23920);
  not g38070 (n_17153, n23924);
  and g38071 (n23925, n_17152, n_17153);
  not g38072 (n_17154, n23925);
  and g38073 (n23926, pi0778, n_17154);
  not g38074 (n_17155, n23916);
  not g38075 (n_17156, n23926);
  and g38076 (n23927, n_17155, n_17156);
  not g38077 (n_17157, n23927);
  and g38078 (n23928, n_11773, n_17157);
  and g38079 (n23929, n17075, n_17137);
  not g38080 (n_17158, n23928);
  not g38081 (n_17159, n23929);
  and g38082 (n23930, n_17158, n_17159);
  and g38083 (n23931, n_11777, n23930);
  and g38084 (n23932, n16639, n23900);
  not g38085 (n_17160, n23931);
  not g38086 (n_17161, n23932);
  and g38087 (n23933, n_17160, n_17161);
  and g38088 (n23934, n_11780, n23933);
  not g38089 (n_17162, n23901);
  not g38090 (n_17163, n23934);
  and g38091 (n23935, n_17162, n_17163);
  and g38092 (n23936, n_11783, n23935);
  and g38093 (n23937, n16631, n23900);
  not g38094 (n_17164, n23936);
  not g38095 (n_17165, n23937);
  and g38096 (n23938, n_17164, n_17165);
  not g38097 (n_17166, n23938);
  and g38098 (n23939, n_11789, n_17166);
  and g38099 (n23940, pi0628, n23900);
  not g38100 (n_17167, n23939);
  not g38101 (n_17168, n23940);
  and g38102 (n23941, n_17167, n_17168);
  not g38103 (n_17169, n23941);
  and g38104 (n23942, n_11794, n_17169);
  and g38105 (n23943, pi0628, n_17166);
  and g38106 (n23944, n_11789, n23900);
  not g38107 (n_17170, n23943);
  not g38108 (n_17171, n23944);
  and g38109 (n23945, n_17170, n_17171);
  not g38110 (n_17172, n23945);
  and g38111 (n23946, pi1156, n_17172);
  not g38112 (n_17173, n23942);
  not g38113 (n_17174, n23946);
  and g38114 (n23947, n_17173, n_17174);
  not g38115 (n_17175, n23947);
  and g38116 (n23948, pi0792, n_17175);
  and g38117 (n23949, n_11787, n_17166);
  not g38118 (n_17176, n23948);
  not g38119 (n_17177, n23949);
  and g38120 (n23950, n_17176, n_17177);
  not g38121 (n_17178, n23950);
  and g38122 (n23951, n_11806, n_17178);
  and g38123 (n23952, pi0647, n23900);
  not g38124 (n_17179, n23951);
  not g38125 (n_17180, n23952);
  and g38126 (n23953, n_17179, n_17180);
  not g38127 (n_17181, n23953);
  and g38128 (n23954, n_11810, n_17181);
  and g38129 (n23955, pi0647, n_17178);
  and g38130 (n23956, n_11806, n23900);
  not g38131 (n_17182, n23955);
  not g38132 (n_17183, n23956);
  and g38133 (n23957, n_17182, n_17183);
  not g38134 (n_17184, n23957);
  and g38135 (n23958, pi1157, n_17184);
  not g38136 (n_17185, n23954);
  not g38137 (n_17186, n23958);
  and g38138 (n23959, n_17185, n_17186);
  not g38139 (n_17187, n23959);
  and g38140 (n23960, pi0787, n_17187);
  and g38141 (n23961, n_11803, n_17178);
  not g38142 (n_17188, n23960);
  not g38143 (n_17189, n23961);
  and g38144 (n23962, n_17188, n_17189);
  not g38145 (n_17190, n23962);
  and g38146 (n23963, n_11819, n_17190);
  not g38147 (n_17191, n23963);
  and g38148 (n23964, pi0715, n_17191);
  and g38149 (n23965, n_15271, n17046);
  and g38150 (n23966, pi0175, n17273);
  not g38151 (n_17192, n23965);
  not g38152 (n_17193, n23966);
  and g38153 (n23967, n_17192, n_17193);
  not g38154 (n_17194, n23967);
  and g38155 (n23968, pi0039, n_17194);
  and g38156 (n23969, pi0766, n_11950);
  not g38157 (n_17195, n23969);
  and g38158 (n23970, pi0175, n_17195);
  and g38159 (n23971, n_7662, pi0766);
  and g38160 (n23972, n17221, n23971);
  not g38167 (n_17199, n23975);
  and g38168 (n23976, n_161, n_17199);
  and g38169 (n23977, pi0766, n17280);
  and g38170 (n23978, pi0038, n_17138);
  not g38171 (n_17200, n23977);
  and g38172 (n23979, n_17200, n23978);
  not g38173 (n_17201, n23976);
  not g38174 (n_17202, n23979);
  and g38175 (n23980, n_17201, n_17202);
  not g38176 (n_17203, n23980);
  and g38177 (n23981, n2571, n_17203);
  not g38178 (n_17204, n23981);
  and g38179 (n23982, n_17145, n_17204);
  not g38180 (n_17205, n23982);
  and g38181 (n23983, n_11960, n_17205);
  and g38182 (n23984, n17117, n_17137);
  not g38183 (n_17206, n23983);
  not g38184 (n_17207, n23984);
  and g38185 (n23985, n_17206, n_17207);
  not g38186 (n_17208, n23985);
  and g38187 (n23986, n_11964, n_17208);
  and g38188 (n23987, n_11967, n_17137);
  and g38189 (n23988, pi0609, n23983);
  not g38190 (n_17209, n23987);
  not g38191 (n_17210, n23988);
  and g38192 (n23989, n_17209, n_17210);
  not g38193 (n_17211, n23989);
  and g38194 (n23990, pi1155, n_17211);
  and g38195 (n23991, n_11972, n_17137);
  and g38196 (n23992, n_11971, n23983);
  not g38197 (n_17212, n23991);
  not g38198 (n_17213, n23992);
  and g38199 (n23993, n_17212, n_17213);
  not g38200 (n_17214, n23993);
  and g38201 (n23994, n_11768, n_17214);
  not g38202 (n_17215, n23990);
  not g38203 (n_17216, n23994);
  and g38204 (n23995, n_17215, n_17216);
  not g38205 (n_17217, n23995);
  and g38206 (n23996, pi0785, n_17217);
  not g38207 (n_17218, n23986);
  not g38208 (n_17219, n23996);
  and g38209 (n23997, n_17218, n_17219);
  not g38210 (n_17220, n23997);
  and g38211 (n23998, n_11981, n_17220);
  and g38212 (n23999, n_11984, n23900);
  and g38213 (n24000, pi0618, n23997);
  not g38214 (n_17221, n23999);
  and g38215 (n24001, pi1154, n_17221);
  not g38216 (n_17222, n24000);
  and g38217 (n24002, n_17222, n24001);
  and g38218 (n24003, n_11984, n23997);
  and g38219 (n24004, pi0618, n23900);
  not g38220 (n_17223, n24004);
  and g38221 (n24005, n_11413, n_17223);
  not g38222 (n_17224, n24003);
  and g38223 (n24006, n_17224, n24005);
  not g38224 (n_17225, n24002);
  not g38225 (n_17226, n24006);
  and g38226 (n24007, n_17225, n_17226);
  not g38227 (n_17227, n24007);
  and g38228 (n24008, pi0781, n_17227);
  not g38229 (n_17228, n23998);
  not g38230 (n_17229, n24008);
  and g38231 (n24009, n_17228, n_17229);
  not g38232 (n_17230, n24009);
  and g38233 (n24010, n_12315, n_17230);
  and g38234 (n24011, n_11821, n23900);
  and g38235 (n24012, pi0619, n24009);
  not g38236 (n_17231, n24011);
  and g38237 (n24013, pi1159, n_17231);
  not g38238 (n_17232, n24012);
  and g38239 (n24014, n_17232, n24013);
  and g38240 (n24015, n_11821, n24009);
  and g38241 (n24016, pi0619, n23900);
  not g38242 (n_17233, n24016);
  and g38243 (n24017, n_11405, n_17233);
  not g38244 (n_17234, n24015);
  and g38245 (n24018, n_17234, n24017);
  not g38246 (n_17235, n24014);
  not g38247 (n_17236, n24018);
  and g38248 (n24019, n_17235, n_17236);
  not g38249 (n_17237, n24019);
  and g38250 (n24020, pi0789, n_17237);
  not g38251 (n_17238, n24010);
  not g38252 (n_17239, n24020);
  and g38253 (n24021, n_17238, n_17239);
  and g38254 (n24022, n_12524, n24021);
  and g38255 (n24023, n17969, n23900);
  not g38256 (n_17240, n24022);
  not g38257 (n_17241, n24023);
  and g38258 (n24024, n_17240, n_17241);
  not g38259 (n_17242, n24024);
  and g38260 (n24025, n_12368, n_17242);
  and g38261 (n24026, n17779, n23900);
  not g38262 (n_17243, n24025);
  not g38263 (n_17244, n24026);
  and g38264 (n24027, n_17243, n_17244);
  not g38265 (n_17245, n24027);
  and g38266 (n24028, n_12392, n_17245);
  and g38267 (n24029, n17804, n23900);
  not g38268 (n_17246, n24028);
  not g38269 (n_17247, n24029);
  and g38270 (n24030, n_17246, n_17247);
  not g38271 (n_17248, n24030);
  and g38272 (n24031, pi0644, n_17248);
  and g38273 (n24032, n_11819, n23900);
  not g38274 (n_17249, n24032);
  and g38275 (n24033, n_12395, n_17249);
  not g38276 (n_17250, n24031);
  and g38277 (n24034, n_17250, n24033);
  not g38278 (n_17251, n24034);
  and g38279 (n24035, pi1160, n_17251);
  not g38280 (n_17252, n23964);
  and g38281 (n24036, n_17252, n24035);
  and g38282 (n24037, pi0644, n_17190);
  not g38283 (n_17253, n24037);
  and g38284 (n24038, n_12395, n_17253);
  and g38285 (n24039, n_11819, n_17248);
  and g38286 (n24040, pi0644, n23900);
  not g38287 (n_17254, n24040);
  and g38288 (n24041, pi0715, n_17254);
  not g38289 (n_17255, n24039);
  and g38290 (n24042, n_17255, n24041);
  not g38291 (n_17256, n24042);
  and g38292 (n24043, n_12405, n_17256);
  not g38293 (n_17257, n24038);
  and g38294 (n24044, n_17257, n24043);
  not g38295 (n_17258, n24036);
  not g38296 (n_17259, n24044);
  and g38297 (n24045, n_17258, n_17259);
  not g38298 (n_17260, n24045);
  and g38299 (n24046, pi0790, n_17260);
  and g38300 (n24047, n17777, n23941);
  and g38301 (n24048, n_14557, n24024);
  and g38302 (n24049, n17776, n23945);
  not g38303 (n_17261, n24047);
  not g38304 (n_17262, n24049);
  and g38305 (n24050, n_17261, n_17262);
  not g38306 (n_17263, n24048);
  and g38307 (n24051, n_17263, n24050);
  not g38308 (n_17264, n24051);
  and g38309 (n24052, pi0792, n_17264);
  and g38310 (n24053, pi0609, n23927);
  and g38311 (n24054, n_15317, n23980);
  and g38312 (n24055, n16667, n_12007);
  and g38313 (n24056, n_15271, n24055);
  not g38314 (n_17265, n24056);
  and g38315 (n24057, n_12250, n_17265);
  not g38316 (n_17266, n24057);
  and g38317 (n24058, n_162, n_17266);
  not g38318 (n_17267, n24058);
  and g38319 (n24059, n_7662, n_17267);
  and g38320 (n24060, n_12120, n_17001);
  not g38321 (n_17268, n24060);
  and g38322 (n24061, pi0175, n_17268);
  and g38323 (n24062, n6284, n24061);
  not g38324 (n_17269, n24062);
  and g38325 (n24063, pi0038, n_17269);
  not g38326 (n_17270, n24059);
  and g38327 (n24064, n_17270, n24063);
  and g38328 (n24065, n_7662, n_12694);
  and g38329 (n24066, pi0175, n_12695);
  not g38330 (n_17271, n24066);
  and g38331 (n24067, pi0766, n_17271);
  not g38332 (n_17272, n24065);
  and g38333 (n24068, n_17272, n24067);
  and g38334 (n24069, n_7662, n17612);
  and g38335 (n24070, pi0175, n17625);
  not g38336 (n_17273, n24069);
  and g38337 (n24071, n_15271, n_17273);
  not g38338 (n_17274, n24070);
  and g38339 (n24072, n_17274, n24071);
  not g38340 (n_17275, n24068);
  and g38341 (n24073, n_162, n_17275);
  not g38342 (n_17276, n24072);
  and g38343 (n24074, n_17276, n24073);
  and g38344 (n24075, pi0175, n17605);
  and g38345 (n24076, n_7662, n_12180);
  not g38346 (n_17277, n24076);
  and g38347 (n24077, pi0766, n_17277);
  not g38348 (n_17278, n24075);
  and g38349 (n24078, n_17278, n24077);
  and g38350 (n24079, n_7662, n17404);
  and g38351 (n24080, pi0175, n17485);
  not g38352 (n_17279, n24080);
  and g38353 (n24081, n_15271, n_17279);
  not g38354 (n_17280, n24079);
  and g38355 (n24082, n_17280, n24081);
  not g38356 (n_17281, n24078);
  and g38357 (n24083, pi0039, n_17281);
  not g38358 (n_17282, n24082);
  and g38359 (n24084, n_17282, n24083);
  not g38360 (n_17283, n24074);
  and g38361 (n24085, n_161, n_17283);
  not g38362 (n_17284, n24084);
  and g38363 (n24086, n_17284, n24085);
  not g38364 (n_17285, n24064);
  and g38365 (n24087, pi0700, n_17285);
  not g38366 (n_17286, n24086);
  and g38367 (n24088, n_17286, n24087);
  not g38368 (n_17287, n24088);
  and g38369 (n24089, n2571, n_17287);
  not g38370 (n_17288, n24054);
  and g38371 (n24090, n_17288, n24089);
  not g38372 (n_17289, n24090);
  and g38373 (n24091, n_17145, n_17289);
  and g38374 (n24092, n_11753, n24091);
  and g38375 (n24093, pi0625, n23982);
  not g38376 (n_17290, n24093);
  and g38377 (n24094, n_11757, n_17290);
  not g38378 (n_17291, n24092);
  and g38379 (n24095, n_17291, n24094);
  and g38380 (n24096, n_11823, n_17152);
  not g38381 (n_17292, n24095);
  and g38382 (n24097, n_17292, n24096);
  and g38383 (n24098, n_11753, n23982);
  and g38384 (n24099, pi0625, n24091);
  not g38385 (n_17293, n24098);
  and g38386 (n24100, pi1153, n_17293);
  not g38387 (n_17294, n24099);
  and g38388 (n24101, n_17294, n24100);
  and g38389 (n24102, pi0608, n_17153);
  not g38390 (n_17295, n24101);
  and g38391 (n24103, n_17295, n24102);
  not g38392 (n_17296, n24097);
  not g38393 (n_17297, n24103);
  and g38394 (n24104, n_17296, n_17297);
  not g38395 (n_17298, n24104);
  and g38396 (n24105, pi0778, n_17298);
  and g38397 (n24106, n_11749, n24091);
  not g38398 (n_17299, n24105);
  not g38399 (n_17300, n24106);
  and g38400 (n24107, n_17299, n_17300);
  not g38401 (n_17301, n24107);
  and g38402 (n24108, n_11971, n_17301);
  not g38403 (n_17302, n24053);
  and g38404 (n24109, n_11768, n_17302);
  not g38405 (n_17303, n24108);
  and g38406 (n24110, n_17303, n24109);
  and g38407 (n24111, n_11767, n_17215);
  not g38408 (n_17304, n24110);
  and g38409 (n24112, n_17304, n24111);
  and g38410 (n24113, n_11971, n23927);
  and g38411 (n24114, pi0609, n_17301);
  not g38412 (n_17305, n24113);
  and g38413 (n24115, pi1155, n_17305);
  not g38414 (n_17306, n24114);
  and g38415 (n24116, n_17306, n24115);
  and g38416 (n24117, pi0660, n_17216);
  not g38417 (n_17307, n24116);
  and g38418 (n24118, n_17307, n24117);
  not g38419 (n_17308, n24112);
  not g38420 (n_17309, n24118);
  and g38421 (n24119, n_17308, n_17309);
  not g38422 (n_17310, n24119);
  and g38423 (n24120, pi0785, n_17310);
  and g38424 (n24121, n_11964, n_17301);
  not g38425 (n_17311, n24120);
  not g38426 (n_17312, n24121);
  and g38427 (n24122, n_17311, n_17312);
  not g38428 (n_17313, n24122);
  and g38429 (n24123, n_11984, n_17313);
  and g38430 (n24124, pi0618, n23930);
  not g38431 (n_17314, n24124);
  and g38432 (n24125, n_11413, n_17314);
  not g38433 (n_17315, n24123);
  and g38434 (n24126, n_17315, n24125);
  and g38435 (n24127, n_11412, n_17225);
  not g38436 (n_17316, n24126);
  and g38437 (n24128, n_17316, n24127);
  and g38438 (n24129, n_11984, n23930);
  and g38439 (n24130, pi0618, n_17313);
  not g38440 (n_17317, n24129);
  and g38441 (n24131, pi1154, n_17317);
  not g38442 (n_17318, n24130);
  and g38443 (n24132, n_17318, n24131);
  and g38444 (n24133, pi0627, n_17226);
  not g38445 (n_17319, n24132);
  and g38446 (n24134, n_17319, n24133);
  not g38447 (n_17320, n24128);
  not g38448 (n_17321, n24134);
  and g38449 (n24135, n_17320, n_17321);
  not g38450 (n_17322, n24135);
  and g38451 (n24136, pi0781, n_17322);
  and g38452 (n24137, n_11981, n_17313);
  not g38453 (n_17323, n24136);
  not g38454 (n_17324, n24137);
  and g38455 (n24138, n_17323, n_17324);
  and g38456 (n24139, n_12315, n24138);
  not g38457 (n_17325, n23933);
  and g38458 (n24140, pi0619, n_17325);
  not g38459 (n_17326, n24138);
  and g38460 (n24141, n_11821, n_17326);
  not g38461 (n_17327, n24140);
  and g38462 (n24142, n_11405, n_17327);
  not g38463 (n_17328, n24141);
  and g38464 (n24143, n_17328, n24142);
  and g38465 (n24144, n_11403, n_17235);
  not g38466 (n_17329, n24143);
  and g38467 (n24145, n_17329, n24144);
  and g38468 (n24146, n_11821, n_17325);
  and g38469 (n24147, pi0619, n_17326);
  not g38470 (n_17330, n24146);
  and g38471 (n24148, pi1159, n_17330);
  not g38472 (n_17331, n24147);
  and g38473 (n24149, n_17331, n24148);
  and g38474 (n24150, pi0648, n_17236);
  not g38475 (n_17332, n24149);
  and g38476 (n24151, n_17332, n24150);
  not g38477 (n_17333, n24145);
  and g38478 (n24152, pi0789, n_17333);
  not g38479 (n_17334, n24151);
  and g38480 (n24153, n_17334, n24152);
  not g38481 (n_17335, n24139);
  and g38482 (n24154, n17970, n_17335);
  not g38483 (n_17336, n24153);
  and g38484 (n24155, n_17336, n24154);
  and g38485 (n24156, n17871, n23935);
  not g38486 (n_17337, n24021);
  and g38487 (n24157, n_12320, n_17337);
  and g38488 (n24158, pi0626, n_17137);
  not g38489 (n_17338, n24158);
  and g38490 (n24159, n16629, n_17338);
  not g38491 (n_17339, n24157);
  and g38492 (n24160, n_17339, n24159);
  and g38493 (n24161, pi0626, n_17337);
  and g38494 (n24162, n_12320, n_17137);
  not g38495 (n_17340, n24162);
  and g38496 (n24163, n16628, n_17340);
  not g38497 (n_17341, n24161);
  and g38498 (n24164, n_17341, n24163);
  not g38499 (n_17342, n24156);
  not g38500 (n_17343, n24160);
  and g38501 (n24165, n_17342, n_17343);
  not g38502 (n_17344, n24164);
  and g38503 (n24166, n_17344, n24165);
  not g38504 (n_17345, n24166);
  and g38505 (n24167, pi0788, n_17345);
  not g38506 (n_17346, n24167);
  and g38507 (n24168, n_14638, n_17346);
  not g38508 (n_17347, n24155);
  and g38509 (n24169, n_17347, n24168);
  not g38510 (n_17348, n24052);
  not g38511 (n_17349, n24169);
  and g38512 (n24170, n_17348, n_17349);
  not g38513 (n_17350, n24170);
  and g38514 (n24171, n_14387, n_17350);
  and g38515 (n24172, n17802, n23953);
  and g38516 (n24173, n_14548, n24027);
  and g38517 (n24174, n17801, n23957);
  not g38518 (n_17351, n24172);
  not g38519 (n_17352, n24173);
  and g38520 (n24175, n_17351, n_17352);
  not g38521 (n_17353, n24174);
  and g38522 (n24176, n_17353, n24175);
  not g38523 (n_17354, n24176);
  and g38524 (n24177, pi0787, n_17354);
  and g38525 (n24178, n_11819, n24043);
  and g38526 (n24179, pi0644, n24035);
  not g38527 (n_17355, n24178);
  and g38528 (n24180, pi0790, n_17355);
  not g38529 (n_17356, n24179);
  and g38530 (n24181, n_17356, n24180);
  not g38531 (n_17357, n24171);
  not g38532 (n_17358, n24177);
  and g38533 (n24182, n_17357, n_17358);
  not g38534 (n_17359, n24181);
  and g38535 (n24183, n_17359, n24182);
  not g38536 (n_17360, n24046);
  not g38537 (n_17361, n24183);
  and g38538 (n24184, n_17360, n_17361);
  not g38539 (n_17362, n24184);
  and g38540 (n24185, n_4226, n_17362);
  not g38541 (n_17363, n23899);
  and g38542 (n24186, n_12415, n_17363);
  not g38543 (n_17364, n24185);
  and g38544 (n24187, n_17364, n24186);
  not g38545 (n_17365, n23898);
  not g38546 (n_17366, n24187);
  and g38547 (po0332, n_17365, n_17366);
  and g38548 (n24189, n_5742, n_12418);
  and g38549 (n24190, n_15329, n16645);
  not g38550 (n_17367, n24189);
  not g38551 (n_17368, n24190);
  and g38552 (n24191, n_17367, n_17368);
  and g38553 (n24192, n_11749, n24191);
  and g38554 (n24193, n_11753, n24190);
  not g38555 (n_17369, n24191);
  not g38556 (n_17370, n24193);
  and g38557 (n24194, n_17369, n_17370);
  not g38558 (n_17371, n24194);
  and g38559 (n24195, pi1153, n_17371);
  and g38560 (n24196, n_11757, n_17367);
  and g38561 (n24197, n_17370, n24196);
  not g38562 (n_17372, n24195);
  not g38563 (n_17373, n24197);
  and g38564 (n24198, n_17372, n_17373);
  not g38565 (n_17374, n24198);
  and g38566 (n24199, pi0778, n_17374);
  not g38567 (n_17375, n24192);
  not g38568 (n_17376, n24199);
  and g38569 (n24200, n_17375, n_17376);
  and g38570 (n24201, n_12429, n24200);
  and g38571 (n24202, n_12430, n24201);
  and g38572 (n24203, n_12431, n24202);
  and g38573 (n24204, n_12432, n24203);
  and g38574 (n24205, n_12436, n24204);
  and g38575 (n24206, n_11806, n24205);
  and g38576 (n24207, pi0647, n24189);
  not g38577 (n_17377, n24207);
  and g38578 (n24208, n_11810, n_17377);
  not g38579 (n_17378, n24206);
  and g38580 (n24209, n_17378, n24208);
  and g38581 (n24210, pi0630, n24209);
  and g38582 (n24211, n_15327, n17244);
  not g38583 (n_17379, n24211);
  and g38584 (n24212, n_17367, n_17379);
  not g38585 (n_17380, n24212);
  and g38586 (n24213, n_12448, n_17380);
  not g38587 (n_17381, n24213);
  and g38588 (n24214, n_11964, n_17381);
  and g38589 (n24215, n_12451, n_17380);
  not g38590 (n_17382, n24215);
  and g38591 (n24216, pi1155, n_17382);
  and g38592 (n24217, n_12453, n24213);
  not g38593 (n_17383, n24217);
  and g38594 (n24218, n_11768, n_17383);
  not g38595 (n_17384, n24216);
  not g38596 (n_17385, n24218);
  and g38597 (n24219, n_17384, n_17385);
  not g38598 (n_17386, n24219);
  and g38599 (n24220, pi0785, n_17386);
  not g38600 (n_17387, n24214);
  not g38601 (n_17388, n24220);
  and g38602 (n24221, n_17387, n_17388);
  not g38603 (n_17389, n24221);
  and g38604 (n24222, n_11981, n_17389);
  and g38605 (n24223, n_12461, n24221);
  not g38606 (n_17390, n24223);
  and g38607 (n24224, pi1154, n_17390);
  and g38608 (n24225, n_12463, n24221);
  not g38609 (n_17391, n24225);
  and g38610 (n24226, n_11413, n_17391);
  not g38611 (n_17392, n24224);
  not g38612 (n_17393, n24226);
  and g38613 (n24227, n_17392, n_17393);
  not g38614 (n_17394, n24227);
  and g38615 (n24228, pi0781, n_17394);
  not g38616 (n_17395, n24222);
  not g38617 (n_17396, n24228);
  and g38618 (n24229, n_17395, n_17396);
  not g38619 (n_17397, n24229);
  and g38620 (n24230, n_12315, n_17397);
  and g38621 (n24231, n_11821, n24189);
  and g38622 (n24232, pi0619, n24229);
  not g38623 (n_17398, n24231);
  and g38624 (n24233, pi1159, n_17398);
  not g38625 (n_17399, n24232);
  and g38626 (n24234, n_17399, n24233);
  and g38627 (n24235, n_11821, n24229);
  and g38628 (n24236, pi0619, n24189);
  not g38629 (n_17400, n24236);
  and g38630 (n24237, n_11405, n_17400);
  not g38631 (n_17401, n24235);
  and g38632 (n24238, n_17401, n24237);
  not g38633 (n_17402, n24234);
  not g38634 (n_17403, n24238);
  and g38635 (n24239, n_17402, n_17403);
  not g38636 (n_17404, n24239);
  and g38637 (n24240, pi0789, n_17404);
  not g38638 (n_17405, n24230);
  not g38639 (n_17406, n24240);
  and g38640 (n24241, n_17405, n_17406);
  and g38641 (n24242, n_12524, n24241);
  and g38642 (n24243, n17969, n24189);
  not g38643 (n_17407, n24242);
  not g38644 (n_17408, n24243);
  and g38645 (n24244, n_17407, n_17408);
  not g38646 (n_17409, n24244);
  and g38647 (n24245, n_12368, n_17409);
  and g38648 (n24246, n17779, n24189);
  not g38649 (n_17410, n24245);
  not g38650 (n_17411, n24246);
  and g38651 (n24247, n_17410, n_17411);
  and g38652 (n24248, n_14548, n24247);
  not g38653 (n_17412, n24205);
  and g38654 (n24249, pi0647, n_17412);
  and g38655 (n24250, n_11806, n_17367);
  not g38656 (n_17413, n24249);
  not g38657 (n_17414, n24250);
  and g38658 (n24251, n_17413, n_17414);
  not g38659 (n_17415, n24251);
  and g38660 (n24252, n17801, n_17415);
  not g38661 (n_17416, n24210);
  not g38662 (n_17417, n24252);
  and g38663 (n24253, n_17416, n_17417);
  not g38664 (n_17418, n24248);
  and g38665 (n24254, n_17418, n24253);
  not g38666 (n_17419, n24254);
  and g38667 (n24255, pi0787, n_17419);
  and g38668 (n24256, n17871, n24203);
  not g38669 (n_17420, n24241);
  and g38670 (n24257, n_12320, n_17420);
  and g38671 (n24258, pi0626, n_17367);
  not g38672 (n_17421, n24258);
  and g38673 (n24259, n16629, n_17421);
  not g38674 (n_17422, n24257);
  and g38675 (n24260, n_17422, n24259);
  and g38676 (n24261, pi0626, n_17420);
  and g38677 (n24262, n_12320, n_17367);
  not g38678 (n_17423, n24262);
  and g38679 (n24263, n16628, n_17423);
  not g38680 (n_17424, n24261);
  and g38681 (n24264, n_17424, n24263);
  not g38682 (n_17425, n24256);
  not g38683 (n_17426, n24260);
  and g38684 (n24265, n_17425, n_17426);
  not g38685 (n_17427, n24264);
  and g38686 (n24266, n_17427, n24265);
  not g38687 (n_17428, n24266);
  and g38688 (n24267, pi0788, n_17428);
  and g38689 (n24268, pi0618, n24201);
  and g38690 (n24269, pi0609, n24200);
  and g38691 (n24270, n_11866, n_17369);
  and g38692 (n24271, pi0625, n24270);
  not g38693 (n_17429, n24270);
  and g38694 (n24272, n24212, n_17429);
  not g38695 (n_17430, n24271);
  not g38696 (n_17431, n24272);
  and g38697 (n24273, n_17430, n_17431);
  not g38698 (n_17432, n24273);
  and g38699 (n24274, n24196, n_17432);
  and g38700 (n24275, n_11823, n_17372);
  not g38701 (n_17433, n24274);
  and g38702 (n24276, n_17433, n24275);
  and g38703 (n24277, pi1153, n24212);
  and g38704 (n24278, n_17430, n24277);
  and g38705 (n24279, pi0608, n_17373);
  not g38706 (n_17434, n24278);
  and g38707 (n24280, n_17434, n24279);
  not g38708 (n_17435, n24276);
  not g38709 (n_17436, n24280);
  and g38710 (n24281, n_17435, n_17436);
  not g38711 (n_17437, n24281);
  and g38712 (n24282, pi0778, n_17437);
  and g38713 (n24283, n_11749, n_17431);
  not g38714 (n_17438, n24282);
  not g38715 (n_17439, n24283);
  and g38716 (n24284, n_17438, n_17439);
  not g38717 (n_17440, n24284);
  and g38718 (n24285, n_11971, n_17440);
  not g38719 (n_17441, n24269);
  and g38720 (n24286, n_11768, n_17441);
  not g38721 (n_17442, n24285);
  and g38722 (n24287, n_17442, n24286);
  and g38723 (n24288, n_11767, n_17384);
  not g38724 (n_17443, n24287);
  and g38725 (n24289, n_17443, n24288);
  and g38726 (n24290, n_11971, n24200);
  and g38727 (n24291, pi0609, n_17440);
  not g38728 (n_17444, n24290);
  and g38729 (n24292, pi1155, n_17444);
  not g38730 (n_17445, n24291);
  and g38731 (n24293, n_17445, n24292);
  and g38732 (n24294, pi0660, n_17385);
  not g38733 (n_17446, n24293);
  and g38734 (n24295, n_17446, n24294);
  not g38735 (n_17447, n24289);
  not g38736 (n_17448, n24295);
  and g38737 (n24296, n_17447, n_17448);
  not g38738 (n_17449, n24296);
  and g38739 (n24297, pi0785, n_17449);
  and g38740 (n24298, n_11964, n_17440);
  not g38741 (n_17450, n24297);
  not g38742 (n_17451, n24298);
  and g38743 (n24299, n_17450, n_17451);
  not g38744 (n_17452, n24299);
  and g38745 (n24300, n_11984, n_17452);
  not g38746 (n_17453, n24268);
  and g38747 (n24301, n_11413, n_17453);
  not g38748 (n_17454, n24300);
  and g38749 (n24302, n_17454, n24301);
  and g38750 (n24303, n_11412, n_17392);
  not g38751 (n_17455, n24302);
  and g38752 (n24304, n_17455, n24303);
  and g38753 (n24305, n_11984, n24201);
  and g38754 (n24306, pi0618, n_17452);
  not g38755 (n_17456, n24305);
  and g38756 (n24307, pi1154, n_17456);
  not g38757 (n_17457, n24306);
  and g38758 (n24308, n_17457, n24307);
  and g38759 (n24309, pi0627, n_17393);
  not g38760 (n_17458, n24308);
  and g38761 (n24310, n_17458, n24309);
  not g38762 (n_17459, n24304);
  not g38763 (n_17460, n24310);
  and g38764 (n24311, n_17459, n_17460);
  not g38765 (n_17461, n24311);
  and g38766 (n24312, pi0781, n_17461);
  and g38767 (n24313, n_11981, n_17452);
  not g38768 (n_17462, n24312);
  not g38769 (n_17463, n24313);
  and g38770 (n24314, n_17462, n_17463);
  and g38771 (n24315, n_12315, n24314);
  not g38772 (n_17464, n24314);
  and g38773 (n24316, n_11821, n_17464);
  and g38774 (n24317, pi0619, n24202);
  not g38775 (n_17465, n24317);
  and g38776 (n24318, n_11405, n_17465);
  not g38777 (n_17466, n24316);
  and g38778 (n24319, n_17466, n24318);
  and g38779 (n24320, n_11403, n_17402);
  not g38780 (n_17467, n24319);
  and g38781 (n24321, n_17467, n24320);
  and g38782 (n24322, pi0619, n_17464);
  and g38783 (n24323, n_11821, n24202);
  not g38784 (n_17468, n24323);
  and g38785 (n24324, pi1159, n_17468);
  not g38786 (n_17469, n24322);
  and g38787 (n24325, n_17469, n24324);
  and g38788 (n24326, pi0648, n_17403);
  not g38789 (n_17470, n24325);
  and g38790 (n24327, n_17470, n24326);
  not g38791 (n_17471, n24321);
  and g38792 (n24328, pi0789, n_17471);
  not g38793 (n_17472, n24327);
  and g38794 (n24329, n_17472, n24328);
  not g38795 (n_17473, n24315);
  and g38796 (n24330, n17970, n_17473);
  not g38797 (n_17474, n24329);
  and g38798 (n24331, n_17474, n24330);
  not g38799 (n_17475, n24267);
  not g38800 (n_17476, n24331);
  and g38801 (n24332, n_17475, n_17476);
  not g38802 (n_17477, n24332);
  and g38803 (n24333, n_14638, n_17477);
  and g38804 (n24334, n17854, n_17409);
  and g38805 (n24335, n20851, n24204);
  not g38806 (n_17478, n24334);
  not g38807 (n_17479, n24335);
  and g38808 (n24336, n_17478, n_17479);
  not g38809 (n_17480, n24336);
  and g38810 (n24337, n_12354, n_17480);
  and g38811 (n24338, n20855, n24204);
  and g38812 (n24339, n17853, n_17409);
  not g38813 (n_17481, n24338);
  not g38814 (n_17482, n24339);
  and g38815 (n24340, n_17481, n_17482);
  not g38816 (n_17483, n24340);
  and g38817 (n24341, pi0629, n_17483);
  not g38818 (n_17484, n24337);
  not g38819 (n_17485, n24341);
  and g38820 (n24342, n_17484, n_17485);
  not g38821 (n_17486, n24342);
  and g38822 (n24343, pi0792, n_17486);
  not g38823 (n_17487, n24343);
  and g38824 (n24344, n_14387, n_17487);
  not g38825 (n_17488, n24333);
  and g38826 (n24345, n_17488, n24344);
  not g38827 (n_17489, n24255);
  not g38828 (n_17490, n24345);
  and g38829 (n24346, n_17489, n_17490);
  and g38830 (n24347, n_12411, n24346);
  and g38831 (n24348, n_11803, n_17412);
  and g38832 (n24349, pi1157, n_17415);
  not g38833 (n_17491, n24209);
  not g38834 (n_17492, n24349);
  and g38835 (n24350, n_17491, n_17492);
  not g38836 (n_17493, n24350);
  and g38837 (n24351, pi0787, n_17493);
  not g38838 (n_17494, n24348);
  not g38839 (n_17495, n24351);
  and g38840 (n24352, n_17494, n_17495);
  and g38841 (n24353, n_11819, n24352);
  and g38842 (n24354, pi0644, n24346);
  not g38843 (n_17496, n24353);
  and g38844 (n24355, pi0715, n_17496);
  not g38845 (n_17497, n24354);
  and g38846 (n24356, n_17497, n24355);
  not g38847 (n_17498, n24247);
  and g38848 (n24357, n_12392, n_17498);
  and g38849 (n24358, n17804, n24189);
  not g38850 (n_17499, n24357);
  not g38851 (n_17500, n24358);
  and g38852 (n24359, n_17499, n_17500);
  not g38853 (n_17501, n24359);
  and g38854 (n24360, pi0644, n_17501);
  and g38855 (n24361, n_11819, n24189);
  not g38856 (n_17502, n24361);
  and g38857 (n24362, n_12395, n_17502);
  not g38858 (n_17503, n24360);
  and g38859 (n24363, n_17503, n24362);
  not g38860 (n_17504, n24363);
  and g38861 (n24364, pi1160, n_17504);
  not g38862 (n_17505, n24356);
  and g38863 (n24365, n_17505, n24364);
  and g38864 (n24366, n_11819, n_17501);
  and g38865 (n24367, pi0644, n24189);
  not g38866 (n_17506, n24367);
  and g38867 (n24368, pi0715, n_17506);
  not g38868 (n_17507, n24366);
  and g38869 (n24369, n_17507, n24368);
  and g38870 (n24370, pi0644, n24352);
  and g38871 (n24371, n_11819, n24346);
  not g38872 (n_17508, n24370);
  and g38873 (n24372, n_12395, n_17508);
  not g38874 (n_17509, n24371);
  and g38875 (n24373, n_17509, n24372);
  not g38876 (n_17510, n24369);
  and g38877 (n24374, n_12405, n_17510);
  not g38878 (n_17511, n24373);
  and g38879 (n24375, n_17511, n24374);
  not g38880 (n_17512, n24365);
  not g38881 (n_17513, n24375);
  and g38882 (n24376, n_17512, n_17513);
  not g38883 (n_17514, n24376);
  and g38884 (n24377, pi0790, n_17514);
  not g38885 (n_17515, n24347);
  and g38886 (n24378, pi0832, n_17515);
  not g38887 (n_17516, n24377);
  and g38888 (n24379, n_17516, n24378);
  and g38889 (n24380, n_5742, po1038);
  and g38890 (n24381, n_5742, n_11751);
  not g38891 (n_17517, n24381);
  and g38892 (n24382, n16635, n_17517);
  and g38893 (n24383, n_161, n18076);
  not g38894 (n_17518, n16647);
  and g38895 (n24384, n2571, n_17518);
  not g38896 (n_17519, n24383);
  and g38897 (n24385, n_17519, n24384);
  not g38898 (n_17520, n24385);
  and g38899 (n24386, pi0176, n_17520);
  and g38900 (n24387, n_161, n18072);
  not g38901 (n_17521, n19899);
  not g38902 (n_17522, n24387);
  and g38903 (n24388, n_17521, n_17522);
  and g38904 (n24389, n_5742, n24388);
  not g38905 (n_17523, n24389);
  and g38906 (n24390, n_15329, n_17523);
  and g38907 (n24391, n_5742, n_11743);
  and g38908 (n24392, pi0704, n24391);
  not g38909 (n_17524, n24392);
  and g38910 (n24393, n2571, n_17524);
  not g38911 (n_17525, n24390);
  and g38912 (n24394, n_17525, n24393);
  not g38913 (n_17526, n24386);
  not g38914 (n_17527, n24394);
  and g38915 (n24395, n_17526, n_17527);
  not g38916 (n_17528, n24395);
  and g38917 (n24396, n_11749, n_17528);
  and g38918 (n24397, n_11753, n24381);
  and g38919 (n24398, pi0625, n24395);
  not g38920 (n_17529, n24397);
  and g38921 (n24399, pi1153, n_17529);
  not g38922 (n_17530, n24398);
  and g38923 (n24400, n_17530, n24399);
  and g38924 (n24401, n_11753, n24395);
  and g38925 (n24402, pi0625, n24381);
  not g38926 (n_17531, n24402);
  and g38927 (n24403, n_11757, n_17531);
  not g38928 (n_17532, n24401);
  and g38929 (n24404, n_17532, n24403);
  not g38930 (n_17533, n24400);
  not g38931 (n_17534, n24404);
  and g38932 (n24405, n_17533, n_17534);
  not g38933 (n_17535, n24405);
  and g38934 (n24406, pi0778, n_17535);
  not g38935 (n_17536, n24396);
  not g38936 (n_17537, n24406);
  and g38937 (n24407, n_17536, n_17537);
  not g38938 (n_17538, n24407);
  and g38939 (n24408, n_11773, n_17538);
  and g38940 (n24409, n17075, n_17517);
  not g38941 (n_17539, n24408);
  not g38942 (n_17540, n24409);
  and g38943 (n24410, n_17539, n_17540);
  and g38944 (n24411, n_11777, n24410);
  and g38945 (n24412, n16639, n24381);
  not g38946 (n_17541, n24411);
  not g38947 (n_17542, n24412);
  and g38948 (n24413, n_17541, n_17542);
  and g38949 (n24414, n_11780, n24413);
  not g38950 (n_17543, n24382);
  not g38951 (n_17544, n24414);
  and g38952 (n24415, n_17543, n_17544);
  and g38953 (n24416, n_11783, n24415);
  and g38954 (n24417, n16631, n24381);
  not g38955 (n_17545, n24416);
  not g38956 (n_17546, n24417);
  and g38957 (n24418, n_17545, n_17546);
  not g38958 (n_17547, n24418);
  and g38959 (n24419, n_11789, n_17547);
  and g38960 (n24420, pi0628, n24381);
  not g38961 (n_17548, n24419);
  not g38962 (n_17549, n24420);
  and g38963 (n24421, n_17548, n_17549);
  not g38964 (n_17550, n24421);
  and g38965 (n24422, n_11794, n_17550);
  and g38966 (n24423, pi0628, n_17547);
  and g38967 (n24424, n_11789, n24381);
  not g38968 (n_17551, n24423);
  not g38969 (n_17552, n24424);
  and g38970 (n24425, n_17551, n_17552);
  not g38971 (n_17553, n24425);
  and g38972 (n24426, pi1156, n_17553);
  not g38973 (n_17554, n24422);
  not g38974 (n_17555, n24426);
  and g38975 (n24427, n_17554, n_17555);
  not g38976 (n_17556, n24427);
  and g38977 (n24428, pi0792, n_17556);
  and g38978 (n24429, n_11787, n_17547);
  not g38979 (n_17557, n24428);
  not g38980 (n_17558, n24429);
  and g38981 (n24430, n_17557, n_17558);
  not g38982 (n_17559, n24430);
  and g38983 (n24431, n_11806, n_17559);
  and g38984 (n24432, pi0647, n24381);
  not g38985 (n_17560, n24431);
  not g38986 (n_17561, n24432);
  and g38987 (n24433, n_17560, n_17561);
  not g38988 (n_17562, n24433);
  and g38989 (n24434, n_11810, n_17562);
  and g38990 (n24435, pi0647, n_17559);
  and g38991 (n24436, n_11806, n24381);
  not g38992 (n_17563, n24435);
  not g38993 (n_17564, n24436);
  and g38994 (n24437, n_17563, n_17564);
  not g38995 (n_17565, n24437);
  and g38996 (n24438, pi1157, n_17565);
  not g38997 (n_17566, n24434);
  not g38998 (n_17567, n24438);
  and g38999 (n24439, n_17566, n_17567);
  not g39000 (n_17568, n24439);
  and g39001 (n24440, pi0787, n_17568);
  and g39002 (n24441, n_11803, n_17559);
  not g39003 (n_17569, n24440);
  not g39004 (n_17570, n24441);
  and g39005 (n24442, n_17569, n_17570);
  not g39006 (n_17571, n24442);
  and g39007 (n24443, n_11819, n_17571);
  not g39008 (n_17572, n24443);
  and g39009 (n24444, pi0715, n_17572);
  and g39010 (n24445, pi0176, n_11417);
  and g39011 (n24446, n_5742, n19439);
  and g39012 (n24447, n_13679, n_13671);
  and g39013 (n24448, pi0176, n24447);
  not g39014 (n_17573, n24446);
  not g39015 (n_17574, n24448);
  and g39016 (n24449, n_17573, n_17574);
  not g39017 (n_17575, n24449);
  and g39018 (n24450, n_15327, n_17575);
  not g39019 (n_17576, n24391);
  and g39020 (n24451, pi0742, n_17576);
  not g39021 (n_17577, n24450);
  not g39022 (n_17578, n24451);
  and g39023 (n24452, n_17577, n_17578);
  not g39024 (n_17579, n24452);
  and g39025 (n24453, n2571, n_17579);
  not g39026 (n_17580, n24445);
  not g39027 (n_17581, n24453);
  and g39028 (n24454, n_17580, n_17581);
  not g39029 (n_17582, n24454);
  and g39030 (n24455, n_11960, n_17582);
  and g39031 (n24456, n17117, n_17517);
  not g39032 (n_17583, n24455);
  not g39033 (n_17584, n24456);
  and g39034 (n24457, n_17583, n_17584);
  not g39035 (n_17585, n24457);
  and g39036 (n24458, n_11964, n_17585);
  and g39037 (n24459, n_11967, n_17517);
  and g39038 (n24460, pi0609, n24455);
  not g39039 (n_17586, n24459);
  not g39040 (n_17587, n24460);
  and g39041 (n24461, n_17586, n_17587);
  not g39042 (n_17588, n24461);
  and g39043 (n24462, pi1155, n_17588);
  and g39044 (n24463, n_11972, n_17517);
  and g39045 (n24464, n_11971, n24455);
  not g39046 (n_17589, n24463);
  not g39047 (n_17590, n24464);
  and g39048 (n24465, n_17589, n_17590);
  not g39049 (n_17591, n24465);
  and g39050 (n24466, n_11768, n_17591);
  not g39051 (n_17592, n24462);
  not g39052 (n_17593, n24466);
  and g39053 (n24467, n_17592, n_17593);
  not g39054 (n_17594, n24467);
  and g39055 (n24468, pi0785, n_17594);
  not g39056 (n_17595, n24458);
  not g39057 (n_17596, n24468);
  and g39058 (n24469, n_17595, n_17596);
  not g39059 (n_17597, n24469);
  and g39060 (n24470, n_11981, n_17597);
  and g39061 (n24471, n_11984, n24381);
  and g39062 (n24472, pi0618, n24469);
  not g39063 (n_17598, n24471);
  and g39064 (n24473, pi1154, n_17598);
  not g39065 (n_17599, n24472);
  and g39066 (n24474, n_17599, n24473);
  and g39067 (n24475, n_11984, n24469);
  and g39068 (n24476, pi0618, n24381);
  not g39069 (n_17600, n24476);
  and g39070 (n24477, n_11413, n_17600);
  not g39071 (n_17601, n24475);
  and g39072 (n24478, n_17601, n24477);
  not g39073 (n_17602, n24474);
  not g39074 (n_17603, n24478);
  and g39075 (n24479, n_17602, n_17603);
  not g39076 (n_17604, n24479);
  and g39077 (n24480, pi0781, n_17604);
  not g39078 (n_17605, n24470);
  not g39079 (n_17606, n24480);
  and g39080 (n24481, n_17605, n_17606);
  not g39081 (n_17607, n24481);
  and g39082 (n24482, n_12315, n_17607);
  and g39083 (n24483, n_11821, n24381);
  and g39084 (n24484, pi0619, n24481);
  not g39085 (n_17608, n24483);
  and g39086 (n24485, pi1159, n_17608);
  not g39087 (n_17609, n24484);
  and g39088 (n24486, n_17609, n24485);
  and g39089 (n24487, n_11821, n24481);
  and g39090 (n24488, pi0619, n24381);
  not g39091 (n_17610, n24488);
  and g39092 (n24489, n_11405, n_17610);
  not g39093 (n_17611, n24487);
  and g39094 (n24490, n_17611, n24489);
  not g39095 (n_17612, n24486);
  not g39096 (n_17613, n24490);
  and g39097 (n24491, n_17612, n_17613);
  not g39098 (n_17614, n24491);
  and g39099 (n24492, pi0789, n_17614);
  not g39100 (n_17615, n24482);
  not g39101 (n_17616, n24492);
  and g39102 (n24493, n_17615, n_17616);
  and g39103 (n24494, n_12524, n24493);
  and g39104 (n24495, n17969, n24381);
  not g39105 (n_17617, n24494);
  not g39106 (n_17618, n24495);
  and g39107 (n24496, n_17617, n_17618);
  not g39108 (n_17619, n24496);
  and g39109 (n24497, n_12368, n_17619);
  and g39110 (n24498, n17779, n24381);
  not g39111 (n_17620, n24497);
  not g39112 (n_17621, n24498);
  and g39113 (n24499, n_17620, n_17621);
  not g39114 (n_17622, n24499);
  and g39115 (n24500, n_12392, n_17622);
  and g39116 (n24501, n17804, n24381);
  not g39117 (n_17623, n24500);
  not g39118 (n_17624, n24501);
  and g39119 (n24502, n_17623, n_17624);
  not g39120 (n_17625, n24502);
  and g39121 (n24503, pi0644, n_17625);
  and g39122 (n24504, n_11819, n24381);
  not g39123 (n_17626, n24504);
  and g39124 (n24505, n_12395, n_17626);
  not g39125 (n_17627, n24503);
  and g39126 (n24506, n_17627, n24505);
  not g39127 (n_17628, n24506);
  and g39128 (n24507, pi1160, n_17628);
  not g39129 (n_17629, n24444);
  and g39130 (n24508, n_17629, n24507);
  and g39131 (n24509, pi0644, n_17571);
  not g39132 (n_17630, n24509);
  and g39133 (n24510, n_12395, n_17630);
  and g39134 (n24511, n_11819, n_17625);
  and g39135 (n24512, pi0644, n24381);
  not g39136 (n_17631, n24512);
  and g39137 (n24513, pi0715, n_17631);
  not g39138 (n_17632, n24511);
  and g39139 (n24514, n_17632, n24513);
  not g39140 (n_17633, n24514);
  and g39141 (n24515, n_12405, n_17633);
  not g39142 (n_17634, n24510);
  and g39143 (n24516, n_17634, n24515);
  not g39144 (n_17635, n24508);
  not g39145 (n_17636, n24516);
  and g39146 (n24517, n_17635, n_17636);
  not g39147 (n_17637, n24517);
  and g39148 (n24518, pi0790, n_17637);
  and g39149 (n24519, n17802, n24433);
  and g39150 (n24520, n_14548, n24499);
  and g39151 (n24521, n17801, n24437);
  not g39152 (n_17638, n24519);
  not g39153 (n_17639, n24520);
  and g39154 (n24522, n_17638, n_17639);
  not g39155 (n_17640, n24521);
  and g39156 (n24523, n_17640, n24522);
  not g39157 (n_17641, n24523);
  and g39158 (n24524, pi0787, n_17641);
  and g39159 (n24525, n17777, n24421);
  and g39160 (n24526, n_14557, n24496);
  and g39161 (n24527, n17776, n24425);
  not g39162 (n_17642, n24525);
  not g39163 (n_17643, n24527);
  and g39164 (n24528, n_17642, n_17643);
  not g39165 (n_17644, n24526);
  and g39166 (n24529, n_17644, n24528);
  not g39167 (n_17645, n24529);
  and g39168 (n24530, pi0792, n_17645);
  and g39169 (n24531, n17871, n24415);
  not g39170 (n_17646, n24493);
  and g39171 (n24532, n_12320, n_17646);
  and g39172 (n24533, pi0626, n_17517);
  not g39173 (n_17647, n24533);
  and g39174 (n24534, n16629, n_17647);
  not g39175 (n_17648, n24532);
  and g39176 (n24535, n_17648, n24534);
  and g39177 (n24536, pi0626, n_17646);
  and g39178 (n24537, n_12320, n_17517);
  not g39179 (n_17649, n24537);
  and g39180 (n24538, n16628, n_17649);
  not g39181 (n_17650, n24536);
  and g39182 (n24539, n_17650, n24538);
  not g39183 (n_17651, n24531);
  not g39184 (n_17652, n24535);
  and g39185 (n24540, n_17651, n_17652);
  not g39186 (n_17653, n24539);
  and g39187 (n24541, n_17653, n24540);
  not g39188 (n_17654, n24541);
  and g39189 (n24542, pi0788, n_17654);
  and g39190 (n24543, pi0609, n24407);
  and g39191 (n24544, n_5742, n_13718);
  and g39192 (n24545, pi0176, n19496);
  not g39193 (n_17655, n24544);
  and g39194 (n24546, n_15327, n_17655);
  not g39195 (n_17656, n24545);
  and g39196 (n24547, n_17656, n24546);
  and g39197 (n24548, n_5742, n19477);
  not g39198 (n_17657, n19468);
  and g39199 (n24549, n_17657, n_13711);
  not g39200 (n_17658, n24549);
  and g39201 (n24550, pi0176, n_17658);
  not g39202 (n_17659, n24550);
  and g39203 (n24551, pi0742, n_17659);
  not g39204 (n_17660, n24548);
  and g39205 (n24552, n_17660, n24551);
  not g39206 (n_17661, n24547);
  and g39207 (n24553, n_15329, n_17661);
  not g39208 (n_17662, n24552);
  and g39209 (n24554, n_17662, n24553);
  and g39210 (n24555, pi0704, n24452);
  not g39211 (n_17663, n24554);
  and g39212 (n24556, n2571, n_17663);
  not g39213 (n_17664, n24555);
  and g39214 (n24557, n_17664, n24556);
  not g39215 (n_17665, n24557);
  and g39216 (n24558, n_17580, n_17665);
  and g39217 (n24559, n_11753, n24558);
  and g39218 (n24560, pi0625, n24454);
  not g39219 (n_17666, n24560);
  and g39220 (n24561, n_11757, n_17666);
  not g39221 (n_17667, n24559);
  and g39222 (n24562, n_17667, n24561);
  and g39223 (n24563, n_11823, n_17533);
  not g39224 (n_17668, n24562);
  and g39225 (n24564, n_17668, n24563);
  and g39226 (n24565, n_11753, n24454);
  and g39227 (n24566, pi0625, n24558);
  not g39228 (n_17669, n24565);
  and g39229 (n24567, pi1153, n_17669);
  not g39230 (n_17670, n24566);
  and g39231 (n24568, n_17670, n24567);
  and g39232 (n24569, pi0608, n_17534);
  not g39233 (n_17671, n24568);
  and g39234 (n24570, n_17671, n24569);
  not g39235 (n_17672, n24564);
  not g39236 (n_17673, n24570);
  and g39237 (n24571, n_17672, n_17673);
  not g39238 (n_17674, n24571);
  and g39239 (n24572, pi0778, n_17674);
  and g39240 (n24573, n_11749, n24558);
  not g39241 (n_17675, n24572);
  not g39242 (n_17676, n24573);
  and g39243 (n24574, n_17675, n_17676);
  not g39244 (n_17677, n24574);
  and g39245 (n24575, n_11971, n_17677);
  not g39246 (n_17678, n24543);
  and g39247 (n24576, n_11768, n_17678);
  not g39248 (n_17679, n24575);
  and g39249 (n24577, n_17679, n24576);
  and g39250 (n24578, n_11767, n_17592);
  not g39251 (n_17680, n24577);
  and g39252 (n24579, n_17680, n24578);
  and g39253 (n24580, n_11971, n24407);
  and g39254 (n24581, pi0609, n_17677);
  not g39255 (n_17681, n24580);
  and g39256 (n24582, pi1155, n_17681);
  not g39257 (n_17682, n24581);
  and g39258 (n24583, n_17682, n24582);
  and g39259 (n24584, pi0660, n_17593);
  not g39260 (n_17683, n24583);
  and g39261 (n24585, n_17683, n24584);
  not g39262 (n_17684, n24579);
  not g39263 (n_17685, n24585);
  and g39264 (n24586, n_17684, n_17685);
  not g39265 (n_17686, n24586);
  and g39266 (n24587, pi0785, n_17686);
  and g39267 (n24588, n_11964, n_17677);
  not g39268 (n_17687, n24587);
  not g39269 (n_17688, n24588);
  and g39270 (n24589, n_17687, n_17688);
  not g39271 (n_17689, n24589);
  and g39272 (n24590, n_11984, n_17689);
  and g39273 (n24591, pi0618, n24410);
  not g39274 (n_17690, n24591);
  and g39275 (n24592, n_11413, n_17690);
  not g39276 (n_17691, n24590);
  and g39277 (n24593, n_17691, n24592);
  and g39278 (n24594, n_11412, n_17602);
  not g39279 (n_17692, n24593);
  and g39280 (n24595, n_17692, n24594);
  and g39281 (n24596, n_11984, n24410);
  and g39282 (n24597, pi0618, n_17689);
  not g39283 (n_17693, n24596);
  and g39284 (n24598, pi1154, n_17693);
  not g39285 (n_17694, n24597);
  and g39286 (n24599, n_17694, n24598);
  and g39287 (n24600, pi0627, n_17603);
  not g39288 (n_17695, n24599);
  and g39289 (n24601, n_17695, n24600);
  not g39290 (n_17696, n24595);
  not g39291 (n_17697, n24601);
  and g39292 (n24602, n_17696, n_17697);
  not g39293 (n_17698, n24602);
  and g39294 (n24603, pi0781, n_17698);
  and g39295 (n24604, n_11981, n_17689);
  not g39296 (n_17699, n24603);
  not g39297 (n_17700, n24604);
  and g39298 (n24605, n_17699, n_17700);
  and g39299 (n24606, n_12315, n24605);
  not g39300 (n_17701, n24413);
  and g39301 (n24607, pi0619, n_17701);
  not g39302 (n_17702, n24605);
  and g39303 (n24608, n_11821, n_17702);
  not g39304 (n_17703, n24607);
  and g39305 (n24609, n_11405, n_17703);
  not g39306 (n_17704, n24608);
  and g39307 (n24610, n_17704, n24609);
  and g39308 (n24611, n_11403, n_17612);
  not g39309 (n_17705, n24610);
  and g39310 (n24612, n_17705, n24611);
  and g39311 (n24613, pi0619, n_17702);
  and g39312 (n24614, n_11821, n_17701);
  not g39313 (n_17706, n24614);
  and g39314 (n24615, pi1159, n_17706);
  not g39315 (n_17707, n24613);
  and g39316 (n24616, n_17707, n24615);
  and g39317 (n24617, pi0648, n_17613);
  not g39318 (n_17708, n24616);
  and g39319 (n24618, n_17708, n24617);
  not g39320 (n_17709, n24612);
  and g39321 (n24619, pi0789, n_17709);
  not g39322 (n_17710, n24618);
  and g39323 (n24620, n_17710, n24619);
  not g39324 (n_17711, n24606);
  and g39325 (n24621, n17970, n_17711);
  not g39326 (n_17712, n24620);
  and g39327 (n24622, n_17712, n24621);
  not g39328 (n_17713, n24542);
  not g39329 (n_17714, n24622);
  and g39330 (n24623, n_17713, n_17714);
  not g39331 (n_17715, n24530);
  not g39332 (n_17716, n24623);
  and g39333 (n24624, n_17715, n_17716);
  and g39334 (n24625, n20364, n24529);
  not g39335 (n_17717, n24625);
  and g39336 (n24626, n_14387, n_17717);
  not g39337 (n_17718, n24624);
  and g39338 (n24627, n_17718, n24626);
  and g39339 (n24628, n_11819, n24515);
  and g39340 (n24629, pi0644, n24507);
  not g39341 (n_17719, n24628);
  and g39342 (n24630, pi0790, n_17719);
  not g39343 (n_17720, n24629);
  and g39344 (n24631, n_17720, n24630);
  not g39345 (n_17721, n24524);
  not g39346 (n_17722, n24627);
  and g39347 (n24632, n_17721, n_17722);
  not g39348 (n_17723, n24631);
  and g39349 (n24633, n_17723, n24632);
  not g39350 (n_17724, n24518);
  not g39351 (n_17725, n24633);
  and g39352 (n24634, n_17724, n_17725);
  not g39353 (n_17726, n24634);
  and g39354 (n24635, n_4226, n_17726);
  not g39355 (n_17727, n24380);
  and g39356 (n24636, n_12415, n_17727);
  not g39357 (n_17728, n24635);
  and g39358 (n24637, n_17728, n24636);
  not g39359 (n_17729, n24379);
  not g39360 (n_17730, n24637);
  and g39361 (po0333, n_17729, n_17730);
  and g39362 (n24639, n_6290, n_11751);
  not g39363 (n_17731, n24639);
  and g39364 (n24640, n16635, n_17731);
  and g39365 (n24641, pi0177, n_11417);
  and g39366 (n24642, n_6290, n18072);
  and g39367 (n24643, pi0177, n_12608);
  not g39368 (n_17732, n24643);
  and g39369 (n24644, n_161, n_17732);
  not g39370 (n_17733, n24642);
  and g39371 (n24645, n_17733, n24644);
  and g39372 (n24646, n_6290, n_11418);
  not g39373 (n_17734, n24646);
  and g39374 (n24647, n16647, n_17734);
  not g39375 (n_17735, n24647);
  and g39376 (n24648, n_15382, n_17735);
  not g39377 (n_17736, n24645);
  and g39378 (n24649, n_17736, n24648);
  and g39379 (n24650, n_6290, pi0686);
  and g39380 (n24651, n_11743, n24650);
  not g39381 (n_17737, n24651);
  and g39382 (n24652, n2571, n_17737);
  not g39383 (n_17738, n24649);
  and g39384 (n24653, n_17738, n24652);
  not g39385 (n_17739, n24641);
  not g39386 (n_17740, n24653);
  and g39387 (n24654, n_17739, n_17740);
  not g39388 (n_17741, n24654);
  and g39389 (n24655, n_11749, n_17741);
  and g39390 (n24656, n_11753, n24639);
  and g39391 (n24657, pi0625, n24654);
  not g39392 (n_17742, n24656);
  and g39393 (n24658, pi1153, n_17742);
  not g39394 (n_17743, n24657);
  and g39395 (n24659, n_17743, n24658);
  and g39396 (n24660, n_11753, n24654);
  and g39397 (n24661, pi0625, n24639);
  not g39398 (n_17744, n24661);
  and g39399 (n24662, n_11757, n_17744);
  not g39400 (n_17745, n24660);
  and g39401 (n24663, n_17745, n24662);
  not g39402 (n_17746, n24659);
  not g39403 (n_17747, n24663);
  and g39404 (n24664, n_17746, n_17747);
  not g39405 (n_17748, n24664);
  and g39406 (n24665, pi0778, n_17748);
  not g39407 (n_17749, n24655);
  not g39408 (n_17750, n24665);
  and g39409 (n24666, n_17749, n_17750);
  not g39410 (n_17751, n24666);
  and g39411 (n24667, n_11773, n_17751);
  and g39412 (n24668, n17075, n_17731);
  not g39413 (n_17752, n24667);
  not g39414 (n_17753, n24668);
  and g39415 (n24669, n_17752, n_17753);
  and g39416 (n24670, n_11777, n24669);
  and g39417 (n24671, n16639, n24639);
  not g39418 (n_17754, n24670);
  not g39419 (n_17755, n24671);
  and g39420 (n24672, n_17754, n_17755);
  and g39421 (n24673, n_11780, n24672);
  not g39422 (n_17756, n24640);
  not g39423 (n_17757, n24673);
  and g39424 (n24674, n_17756, n_17757);
  and g39425 (n24675, n_11783, n24674);
  and g39426 (n24676, n16631, n24639);
  not g39427 (n_17758, n24675);
  not g39428 (n_17759, n24676);
  and g39429 (n24677, n_17758, n_17759);
  and g39430 (n24678, n_11787, n24677);
  and g39431 (n24679, n_11789, n24639);
  not g39432 (n_17760, n24677);
  and g39433 (n24680, pi0628, n_17760);
  not g39434 (n_17761, n24679);
  and g39435 (n24681, pi1156, n_17761);
  not g39436 (n_17762, n24680);
  and g39437 (n24682, n_17762, n24681);
  and g39438 (n24683, pi0628, n24639);
  and g39439 (n24684, n_11789, n_17760);
  not g39440 (n_17763, n24683);
  and g39441 (n24685, n_11794, n_17763);
  not g39442 (n_17764, n24684);
  and g39443 (n24686, n_17764, n24685);
  not g39444 (n_17765, n24682);
  not g39445 (n_17766, n24686);
  and g39446 (n24687, n_17765, n_17766);
  not g39447 (n_17767, n24687);
  and g39448 (n24688, pi0792, n_17767);
  not g39449 (n_17768, n24678);
  not g39450 (n_17769, n24688);
  and g39451 (n24689, n_17768, n_17769);
  not g39452 (n_17770, n24689);
  and g39453 (n24690, n_11803, n_17770);
  and g39454 (n24691, n_11806, n24639);
  and g39455 (n24692, pi0647, n24689);
  not g39456 (n_17771, n24691);
  and g39457 (n24693, pi1157, n_17771);
  not g39458 (n_17772, n24692);
  and g39459 (n24694, n_17772, n24693);
  and g39460 (n24695, n_11806, n24689);
  and g39461 (n24696, pi0647, n24639);
  not g39462 (n_17773, n24696);
  and g39463 (n24697, n_11810, n_17773);
  not g39464 (n_17774, n24695);
  and g39465 (n24698, n_17774, n24697);
  not g39466 (n_17775, n24694);
  not g39467 (n_17776, n24698);
  and g39468 (n24699, n_17775, n_17776);
  not g39469 (n_17777, n24699);
  and g39470 (n24700, pi0787, n_17777);
  not g39471 (n_17778, n24690);
  not g39472 (n_17779, n24700);
  and g39473 (n24701, n_17778, n_17779);
  and g39474 (n24702, n_11819, n24701);
  and g39475 (n24703, n_11821, n24639);
  not g39476 (n_17780, n19439);
  and g39477 (n24704, n_15373, n_17780);
  not g39478 (n_17781, n24704);
  and g39479 (n24705, n_15396, n_17781);
  not g39480 (n_17782, n24705);
  and g39481 (n24706, n_6290, n_17782);
  and g39482 (n24707, n_6290, n_13679);
  not g39483 (n_17783, n24707);
  and g39484 (n24708, n_15373, n_17783);
  not g39485 (n_17784, n24447);
  and g39486 (n24709, n_17784, n24708);
  not g39487 (n_17785, n24706);
  not g39488 (n_17786, n24709);
  and g39489 (n24710, n_17785, n_17786);
  and g39490 (n24711, n2571, n24710);
  not g39491 (n_17787, n24711);
  and g39492 (n24712, n_17739, n_17787);
  not g39493 (n_17788, n24712);
  and g39494 (n24713, n_11960, n_17788);
  and g39495 (n24714, n17117, n_17731);
  not g39496 (n_17789, n24713);
  not g39497 (n_17790, n24714);
  and g39498 (n24715, n_17789, n_17790);
  not g39499 (n_17791, n24715);
  and g39500 (n24716, n_11964, n_17791);
  and g39501 (n24717, n_11967, n_17731);
  and g39502 (n24718, pi0609, n24713);
  not g39503 (n_17792, n24717);
  not g39504 (n_17793, n24718);
  and g39505 (n24719, n_17792, n_17793);
  not g39506 (n_17794, n24719);
  and g39507 (n24720, pi1155, n_17794);
  and g39508 (n24721, n_11972, n_17731);
  and g39509 (n24722, n_11971, n24713);
  not g39510 (n_17795, n24721);
  not g39511 (n_17796, n24722);
  and g39512 (n24723, n_17795, n_17796);
  not g39513 (n_17797, n24723);
  and g39514 (n24724, n_11768, n_17797);
  not g39515 (n_17798, n24720);
  not g39516 (n_17799, n24724);
  and g39517 (n24725, n_17798, n_17799);
  not g39518 (n_17800, n24725);
  and g39519 (n24726, pi0785, n_17800);
  not g39520 (n_17801, n24716);
  not g39521 (n_17802, n24726);
  and g39522 (n24727, n_17801, n_17802);
  not g39523 (n_17803, n24727);
  and g39524 (n24728, n_11981, n_17803);
  and g39525 (n24729, n_11984, n24639);
  and g39526 (n24730, pi0618, n24727);
  not g39527 (n_17804, n24729);
  and g39528 (n24731, pi1154, n_17804);
  not g39529 (n_17805, n24730);
  and g39530 (n24732, n_17805, n24731);
  and g39531 (n24733, n_11984, n24727);
  and g39532 (n24734, pi0618, n24639);
  not g39533 (n_17806, n24734);
  and g39534 (n24735, n_11413, n_17806);
  not g39535 (n_17807, n24733);
  and g39536 (n24736, n_17807, n24735);
  not g39537 (n_17808, n24732);
  not g39538 (n_17809, n24736);
  and g39539 (n24737, n_17808, n_17809);
  not g39540 (n_17810, n24737);
  and g39541 (n24738, pi0781, n_17810);
  not g39542 (n_17811, n24728);
  not g39543 (n_17812, n24738);
  and g39544 (n24739, n_17811, n_17812);
  and g39545 (n24740, pi0619, n24739);
  not g39546 (n_17813, n24703);
  and g39547 (n24741, pi1159, n_17813);
  not g39548 (n_17814, n24740);
  and g39549 (n24742, n_17814, n24741);
  and g39550 (n24743, n18176, n_17734);
  and g39551 (n24744, n_6290, n19475);
  and g39552 (n24745, pi0177, n19467);
  not g39553 (n_17815, n24745);
  and g39554 (n24746, n_161, n_17815);
  not g39555 (n_17816, n24744);
  and g39556 (n24747, n_17816, n24746);
  not g39557 (n_17817, n24743);
  and g39558 (n24748, pi0757, n_17817);
  not g39559 (n_17818, n24747);
  and g39560 (n24749, n_17818, n24748);
  and g39561 (n24750, n_6290, n_13714);
  and g39562 (n24751, pi0177, n19490);
  not g39563 (n_17819, n24751);
  and g39564 (n24752, pi0038, n_17819);
  not g39565 (n_17820, n24750);
  and g39566 (n24753, n_17820, n24752);
  not g39567 (n_17821, n19482);
  and g39568 (n24754, n_17821, n_13717);
  not g39569 (n_17822, n24754);
  and g39570 (n24755, n_6290, n_17822);
  and g39571 (n24756, pi0177, n19494);
  not g39572 (n_17823, n24755);
  and g39573 (n24757, n_161, n_17823);
  not g39574 (n_17824, n24756);
  and g39575 (n24758, n_17824, n24757);
  not g39576 (n_17825, n24753);
  and g39577 (n24759, n_15373, n_17825);
  not g39578 (n_17826, n24758);
  and g39579 (n24760, n_17826, n24759);
  not g39580 (n_17827, n24749);
  not g39581 (n_17828, n24760);
  and g39582 (n24761, n_17827, n_17828);
  not g39583 (n_17829, n24761);
  and g39584 (n24762, n_15382, n_17829);
  not g39585 (n_17830, n24710);
  and g39586 (n24763, pi0686, n_17830);
  not g39587 (n_17831, n24762);
  and g39588 (n24764, n2571, n_17831);
  not g39589 (n_17832, n24763);
  and g39590 (n24765, n_17832, n24764);
  not g39591 (n_17833, n24765);
  and g39592 (n24766, n_17739, n_17833);
  and g39593 (n24767, n_11753, n24766);
  and g39594 (n24768, pi0625, n24712);
  not g39595 (n_17834, n24768);
  and g39596 (n24769, n_11757, n_17834);
  not g39597 (n_17835, n24767);
  and g39598 (n24770, n_17835, n24769);
  and g39599 (n24771, n_11823, n_17746);
  not g39600 (n_17836, n24770);
  and g39601 (n24772, n_17836, n24771);
  and g39602 (n24773, n_11753, n24712);
  and g39603 (n24774, pi0625, n24766);
  not g39604 (n_17837, n24773);
  and g39605 (n24775, pi1153, n_17837);
  not g39606 (n_17838, n24774);
  and g39607 (n24776, n_17838, n24775);
  and g39608 (n24777, pi0608, n_17747);
  not g39609 (n_17839, n24776);
  and g39610 (n24778, n_17839, n24777);
  not g39611 (n_17840, n24772);
  not g39612 (n_17841, n24778);
  and g39613 (n24779, n_17840, n_17841);
  not g39614 (n_17842, n24779);
  and g39615 (n24780, pi0778, n_17842);
  and g39616 (n24781, n_11749, n24766);
  not g39617 (n_17843, n24780);
  not g39618 (n_17844, n24781);
  and g39619 (n24782, n_17843, n_17844);
  not g39620 (n_17845, n24782);
  and g39621 (n24783, n_11971, n_17845);
  and g39622 (n24784, pi0609, n24666);
  not g39623 (n_17846, n24784);
  and g39624 (n24785, n_11768, n_17846);
  not g39625 (n_17847, n24783);
  and g39626 (n24786, n_17847, n24785);
  and g39627 (n24787, n_11767, n_17798);
  not g39628 (n_17848, n24786);
  and g39629 (n24788, n_17848, n24787);
  and g39630 (n24789, n_11971, n24666);
  and g39631 (n24790, pi0609, n_17845);
  not g39632 (n_17849, n24789);
  and g39633 (n24791, pi1155, n_17849);
  not g39634 (n_17850, n24790);
  and g39635 (n24792, n_17850, n24791);
  and g39636 (n24793, pi0660, n_17799);
  not g39637 (n_17851, n24792);
  and g39638 (n24794, n_17851, n24793);
  not g39639 (n_17852, n24788);
  not g39640 (n_17853, n24794);
  and g39641 (n24795, n_17852, n_17853);
  not g39642 (n_17854, n24795);
  and g39643 (n24796, pi0785, n_17854);
  and g39644 (n24797, n_11964, n_17845);
  not g39645 (n_17855, n24796);
  not g39646 (n_17856, n24797);
  and g39647 (n24798, n_17855, n_17856);
  not g39648 (n_17857, n24798);
  and g39649 (n24799, n_11984, n_17857);
  and g39650 (n24800, pi0618, n24669);
  not g39651 (n_17858, n24800);
  and g39652 (n24801, n_11413, n_17858);
  not g39653 (n_17859, n24799);
  and g39654 (n24802, n_17859, n24801);
  and g39655 (n24803, n_11412, n_17808);
  not g39656 (n_17860, n24802);
  and g39657 (n24804, n_17860, n24803);
  and g39658 (n24805, n_11984, n24669);
  and g39659 (n24806, pi0618, n_17857);
  not g39660 (n_17861, n24805);
  and g39661 (n24807, pi1154, n_17861);
  not g39662 (n_17862, n24806);
  and g39663 (n24808, n_17862, n24807);
  and g39664 (n24809, pi0627, n_17809);
  not g39665 (n_17863, n24808);
  and g39666 (n24810, n_17863, n24809);
  not g39667 (n_17864, n24804);
  not g39668 (n_17865, n24810);
  and g39669 (n24811, n_17864, n_17865);
  not g39670 (n_17866, n24811);
  and g39671 (n24812, pi0781, n_17866);
  and g39672 (n24813, n_11981, n_17857);
  not g39673 (n_17867, n24812);
  not g39674 (n_17868, n24813);
  and g39675 (n24814, n_17867, n_17868);
  not g39676 (n_17869, n24814);
  and g39677 (n24815, n_11821, n_17869);
  not g39678 (n_17870, n24672);
  and g39679 (n24816, pi0619, n_17870);
  not g39680 (n_17871, n24816);
  and g39681 (n24817, n_11405, n_17871);
  not g39682 (n_17872, n24815);
  and g39683 (n24818, n_17872, n24817);
  not g39684 (n_17873, n24742);
  and g39685 (n24819, n_11403, n_17873);
  not g39686 (n_17874, n24818);
  and g39687 (n24820, n_17874, n24819);
  and g39688 (n24821, n_11821, n24739);
  and g39689 (n24822, pi0619, n24639);
  not g39690 (n_17875, n24822);
  and g39691 (n24823, n_11405, n_17875);
  not g39692 (n_17876, n24821);
  and g39693 (n24824, n_17876, n24823);
  and g39694 (n24825, pi0619, n_17869);
  and g39695 (n24826, n_11821, n_17870);
  not g39696 (n_17877, n24826);
  and g39697 (n24827, pi1159, n_17877);
  not g39698 (n_17878, n24825);
  and g39699 (n24828, n_17878, n24827);
  not g39700 (n_17879, n24824);
  and g39701 (n24829, pi0648, n_17879);
  not g39702 (n_17880, n24828);
  and g39703 (n24830, n_17880, n24829);
  not g39704 (n_17881, n24820);
  not g39705 (n_17882, n24830);
  and g39706 (n24831, n_17881, n_17882);
  not g39707 (n_17883, n24831);
  and g39708 (n24832, pi0789, n_17883);
  and g39709 (n24833, n_12315, n_17869);
  not g39710 (n_17884, n24832);
  not g39711 (n_17885, n24833);
  and g39712 (n24834, n_17884, n_17885);
  and g39713 (n24835, n_12318, n24834);
  and g39714 (n24836, n_12320, n24834);
  not g39715 (n_17886, n24674);
  and g39716 (n24837, pi0626, n_17886);
  not g39717 (n_17887, n24837);
  and g39718 (n24838, n_11395, n_17887);
  not g39719 (n_17888, n24836);
  and g39720 (n24839, n_17888, n24838);
  not g39721 (n_17889, n24739);
  and g39722 (n24840, n_12315, n_17889);
  and g39723 (n24841, n_17873, n_17879);
  not g39724 (n_17890, n24841);
  and g39725 (n24842, pi0789, n_17890);
  not g39726 (n_17891, n24840);
  not g39727 (n_17892, n24842);
  and g39728 (n24843, n_17891, n_17892);
  not g39729 (n_17893, n24843);
  and g39730 (n24844, n_12320, n_17893);
  and g39731 (n24845, pi0626, n_17731);
  not g39732 (n_17894, n24845);
  and g39733 (n24846, pi0641, n_17894);
  not g39734 (n_17895, n24844);
  and g39735 (n24847, n_17895, n24846);
  not g39736 (n_17896, n24847);
  and g39737 (n24848, n_11397, n_17896);
  not g39738 (n_17897, n24839);
  and g39739 (n24849, n_17897, n24848);
  and g39740 (n24850, pi0626, n24834);
  and g39741 (n24851, n_12320, n_17886);
  not g39742 (n_17898, n24851);
  and g39743 (n24852, pi0641, n_17898);
  not g39744 (n_17899, n24850);
  and g39745 (n24853, n_17899, n24852);
  and g39746 (n24854, pi0626, n_17893);
  and g39747 (n24855, n_12320, n_17731);
  not g39748 (n_17900, n24855);
  and g39749 (n24856, n_11395, n_17900);
  not g39750 (n_17901, n24854);
  and g39751 (n24857, n_17901, n24856);
  not g39752 (n_17902, n24857);
  and g39753 (n24858, pi1158, n_17902);
  not g39754 (n_17903, n24853);
  and g39755 (n24859, n_17903, n24858);
  not g39756 (n_17904, n24849);
  not g39757 (n_17905, n24859);
  and g39758 (n24860, n_17904, n_17905);
  not g39759 (n_17906, n24860);
  and g39760 (n24861, pi0788, n_17906);
  not g39761 (n_17907, n24835);
  not g39762 (n_17908, n24861);
  and g39763 (n24862, n_17907, n_17908);
  and g39764 (n24863, n_11789, n24862);
  and g39765 (n24864, n_12524, n24843);
  and g39766 (n24865, n17969, n24639);
  not g39767 (n_17909, n24864);
  not g39768 (n_17910, n24865);
  and g39769 (n24866, n_17909, n_17910);
  not g39770 (n_17911, n24866);
  and g39771 (n24867, pi0628, n_17911);
  not g39772 (n_17912, n24867);
  and g39773 (n24868, n_11794, n_17912);
  not g39774 (n_17913, n24863);
  and g39775 (n24869, n_17913, n24868);
  and g39776 (n24870, n_12354, n_17765);
  not g39777 (n_17914, n24869);
  and g39778 (n24871, n_17914, n24870);
  and g39779 (n24872, pi0628, n24862);
  and g39780 (n24873, n_11789, n_17911);
  not g39781 (n_17915, n24873);
  and g39782 (n24874, pi1156, n_17915);
  not g39783 (n_17916, n24872);
  and g39784 (n24875, n_17916, n24874);
  and g39785 (n24876, pi0629, n_17766);
  not g39786 (n_17917, n24875);
  and g39787 (n24877, n_17917, n24876);
  not g39788 (n_17918, n24871);
  not g39789 (n_17919, n24877);
  and g39790 (n24878, n_17918, n_17919);
  not g39791 (n_17920, n24878);
  and g39792 (n24879, pi0792, n_17920);
  and g39793 (n24880, n_11787, n24862);
  not g39794 (n_17921, n24879);
  not g39795 (n_17922, n24880);
  and g39796 (n24881, n_17921, n_17922);
  not g39797 (n_17923, n24881);
  and g39798 (n24882, n_11806, n_17923);
  and g39799 (n24883, n_12368, n_17911);
  and g39800 (n24884, n17779, n24639);
  not g39801 (n_17924, n24883);
  not g39802 (n_17925, n24884);
  and g39803 (n24885, n_17924, n_17925);
  not g39804 (n_17926, n24885);
  and g39805 (n24886, pi0647, n_17926);
  not g39806 (n_17927, n24886);
  and g39807 (n24887, n_11810, n_17927);
  not g39808 (n_17928, n24882);
  and g39809 (n24888, n_17928, n24887);
  and g39810 (n24889, n_12375, n_17775);
  not g39811 (n_17929, n24888);
  and g39812 (n24890, n_17929, n24889);
  and g39813 (n24891, pi0647, n_17923);
  and g39814 (n24892, n_11806, n_17926);
  not g39815 (n_17930, n24892);
  and g39816 (n24893, pi1157, n_17930);
  not g39817 (n_17931, n24891);
  and g39818 (n24894, n_17931, n24893);
  and g39819 (n24895, pi0630, n_17776);
  not g39820 (n_17932, n24894);
  and g39821 (n24896, n_17932, n24895);
  not g39822 (n_17933, n24890);
  not g39823 (n_17934, n24896);
  and g39824 (n24897, n_17933, n_17934);
  not g39825 (n_17935, n24897);
  and g39826 (n24898, pi0787, n_17935);
  and g39827 (n24899, n_11803, n_17923);
  not g39828 (n_17936, n24898);
  not g39829 (n_17937, n24899);
  and g39830 (n24900, n_17936, n_17937);
  not g39831 (n_17938, n24900);
  and g39832 (n24901, pi0644, n_17938);
  not g39833 (n_17939, n24702);
  and g39834 (n24902, pi0715, n_17939);
  not g39835 (n_17940, n24901);
  and g39836 (n24903, n_17940, n24902);
  and g39837 (n24904, n17804, n_17731);
  and g39838 (n24905, n_12392, n24885);
  not g39839 (n_17941, n24904);
  not g39840 (n_17942, n24905);
  and g39841 (n24906, n_17941, n_17942);
  and g39842 (n24907, pi0644, n24906);
  and g39843 (n24908, n_11819, n24639);
  not g39844 (n_17943, n24908);
  and g39845 (n24909, n_12395, n_17943);
  not g39846 (n_17944, n24907);
  and g39847 (n24910, n_17944, n24909);
  not g39848 (n_17945, n24910);
  and g39849 (n24911, pi1160, n_17945);
  not g39850 (n_17946, n24903);
  and g39851 (n24912, n_17946, n24911);
  and g39852 (n24913, n_11819, n_17938);
  and g39853 (n24914, pi0644, n24701);
  not g39854 (n_17947, n24914);
  and g39855 (n24915, n_12395, n_17947);
  not g39856 (n_17948, n24913);
  and g39857 (n24916, n_17948, n24915);
  and g39858 (n24917, n_11819, n24906);
  and g39859 (n24918, pi0644, n24639);
  not g39860 (n_17949, n24918);
  and g39861 (n24919, pi0715, n_17949);
  not g39862 (n_17950, n24917);
  and g39863 (n24920, n_17950, n24919);
  not g39864 (n_17951, n24920);
  and g39865 (n24921, n_12405, n_17951);
  not g39866 (n_17952, n24916);
  and g39867 (n24922, n_17952, n24921);
  not g39868 (n_17953, n24912);
  and g39869 (n24923, pi0790, n_17953);
  not g39870 (n_17954, n24922);
  and g39871 (n24924, n_17954, n24923);
  and g39872 (n24925, n_12411, n24900);
  not g39873 (n_17955, n24925);
  and g39874 (n24926, n_4226, n_17955);
  not g39875 (n_17956, n24924);
  and g39876 (n24927, n_17956, n24926);
  and g39877 (n24928, n_6290, po1038);
  not g39878 (n_17957, n24928);
  and g39879 (n24929, n_12415, n_17957);
  not g39880 (n_17958, n24927);
  and g39881 (n24930, n_17958, n24929);
  and g39882 (n24931, n_6290, n_12418);
  and g39883 (n24932, n_15382, n16645);
  not g39884 (n_17959, n24931);
  not g39885 (n_17960, n24932);
  and g39886 (n24933, n_17959, n_17960);
  and g39887 (n24934, n_11749, n24933);
  and g39888 (n24935, n_11753, n24932);
  not g39889 (n_17961, n24933);
  not g39890 (n_17962, n24935);
  and g39891 (n24936, n_17961, n_17962);
  not g39892 (n_17963, n24936);
  and g39893 (n24937, pi1153, n_17963);
  and g39894 (n24938, n_11757, n_17959);
  and g39895 (n24939, n_17962, n24938);
  not g39896 (n_17964, n24937);
  not g39897 (n_17965, n24939);
  and g39898 (n24940, n_17964, n_17965);
  not g39899 (n_17966, n24940);
  and g39900 (n24941, pi0778, n_17966);
  not g39901 (n_17967, n24934);
  not g39902 (n_17968, n24941);
  and g39903 (n24942, n_17967, n_17968);
  and g39904 (n24943, n_12429, n24942);
  and g39905 (n24944, n_12430, n24943);
  and g39906 (n24945, n_12431, n24944);
  and g39907 (n24946, n_12432, n24945);
  and g39908 (n24947, n_12436, n24946);
  and g39909 (n24948, n_11806, n24947);
  and g39910 (n24949, pi0647, n24931);
  not g39911 (n_17969, n24949);
  and g39912 (n24950, n_11810, n_17969);
  not g39913 (n_17970, n24948);
  and g39914 (n24951, n_17970, n24950);
  and g39915 (n24952, pi0630, n24951);
  and g39916 (n24953, n_15373, n17244);
  not g39917 (n_17971, n24953);
  and g39918 (n24954, n_17959, n_17971);
  not g39919 (n_17972, n24954);
  and g39920 (n24955, n_12448, n_17972);
  not g39921 (n_17973, n24955);
  and g39922 (n24956, n_11964, n_17973);
  and g39923 (n24957, n_12451, n_17972);
  not g39924 (n_17974, n24957);
  and g39925 (n24958, pi1155, n_17974);
  and g39926 (n24959, n_12453, n24955);
  not g39927 (n_17975, n24959);
  and g39928 (n24960, n_11768, n_17975);
  not g39929 (n_17976, n24958);
  not g39930 (n_17977, n24960);
  and g39931 (n24961, n_17976, n_17977);
  not g39932 (n_17978, n24961);
  and g39933 (n24962, pi0785, n_17978);
  not g39934 (n_17979, n24956);
  not g39935 (n_17980, n24962);
  and g39936 (n24963, n_17979, n_17980);
  not g39937 (n_17981, n24963);
  and g39938 (n24964, n_11981, n_17981);
  and g39939 (n24965, n_12461, n24963);
  not g39940 (n_17982, n24965);
  and g39941 (n24966, pi1154, n_17982);
  and g39942 (n24967, n_12463, n24963);
  not g39943 (n_17983, n24967);
  and g39944 (n24968, n_11413, n_17983);
  not g39945 (n_17984, n24966);
  not g39946 (n_17985, n24968);
  and g39947 (n24969, n_17984, n_17985);
  not g39948 (n_17986, n24969);
  and g39949 (n24970, pi0781, n_17986);
  not g39950 (n_17987, n24964);
  not g39951 (n_17988, n24970);
  and g39952 (n24971, n_17987, n_17988);
  not g39953 (n_17989, n24971);
  and g39954 (n24972, n_12315, n_17989);
  and g39955 (n24973, n_11821, n24931);
  and g39956 (n24974, pi0619, n24971);
  not g39957 (n_17990, n24973);
  and g39958 (n24975, pi1159, n_17990);
  not g39959 (n_17991, n24974);
  and g39960 (n24976, n_17991, n24975);
  and g39961 (n24977, n_11821, n24971);
  and g39962 (n24978, pi0619, n24931);
  not g39963 (n_17992, n24978);
  and g39964 (n24979, n_11405, n_17992);
  not g39965 (n_17993, n24977);
  and g39966 (n24980, n_17993, n24979);
  not g39967 (n_17994, n24976);
  not g39968 (n_17995, n24980);
  and g39969 (n24981, n_17994, n_17995);
  not g39970 (n_17996, n24981);
  and g39971 (n24982, pi0789, n_17996);
  not g39972 (n_17997, n24972);
  not g39973 (n_17998, n24982);
  and g39974 (n24983, n_17997, n_17998);
  and g39975 (n24984, n_12524, n24983);
  and g39976 (n24985, n17969, n24931);
  not g39977 (n_17999, n24984);
  not g39978 (n_18000, n24985);
  and g39979 (n24986, n_17999, n_18000);
  not g39980 (n_18001, n24986);
  and g39981 (n24987, n_12368, n_18001);
  and g39982 (n24988, n17779, n24931);
  not g39983 (n_18002, n24987);
  not g39984 (n_18003, n24988);
  and g39985 (n24989, n_18002, n_18003);
  and g39986 (n24990, n_14548, n24989);
  not g39987 (n_18004, n24947);
  and g39988 (n24991, pi0647, n_18004);
  and g39989 (n24992, n_11806, n_17959);
  not g39990 (n_18005, n24991);
  not g39991 (n_18006, n24992);
  and g39992 (n24993, n_18005, n_18006);
  not g39993 (n_18007, n24993);
  and g39994 (n24994, n17801, n_18007);
  not g39995 (n_18008, n24952);
  not g39996 (n_18009, n24994);
  and g39997 (n24995, n_18008, n_18009);
  not g39998 (n_18010, n24990);
  and g39999 (n24996, n_18010, n24995);
  not g40000 (n_18011, n24996);
  and g40001 (n24997, pi0787, n_18011);
  and g40002 (n24998, n17871, n24945);
  not g40003 (n_18012, n24983);
  and g40004 (n24999, n_12320, n_18012);
  and g40005 (n25000, pi0626, n_17959);
  not g40006 (n_18013, n25000);
  and g40007 (n25001, n16629, n_18013);
  not g40008 (n_18014, n24999);
  and g40009 (n25002, n_18014, n25001);
  and g40010 (n25003, pi0626, n_18012);
  and g40011 (n25004, n_12320, n_17959);
  not g40012 (n_18015, n25004);
  and g40013 (n25005, n16628, n_18015);
  not g40014 (n_18016, n25003);
  and g40015 (n25006, n_18016, n25005);
  not g40016 (n_18017, n24998);
  not g40017 (n_18018, n25002);
  and g40018 (n25007, n_18017, n_18018);
  not g40019 (n_18019, n25006);
  and g40020 (n25008, n_18019, n25007);
  not g40021 (n_18020, n25008);
  and g40022 (n25009, pi0788, n_18020);
  and g40023 (n25010, pi0618, n24943);
  and g40024 (n25011, pi0609, n24942);
  and g40025 (n25012, n_11866, n_17961);
  and g40026 (n25013, pi0625, n25012);
  not g40027 (n_18021, n25012);
  and g40028 (n25014, n24954, n_18021);
  not g40029 (n_18022, n25013);
  not g40030 (n_18023, n25014);
  and g40031 (n25015, n_18022, n_18023);
  not g40032 (n_18024, n25015);
  and g40033 (n25016, n24938, n_18024);
  and g40034 (n25017, n_11823, n_17964);
  not g40035 (n_18025, n25016);
  and g40036 (n25018, n_18025, n25017);
  and g40037 (n25019, pi1153, n24954);
  and g40038 (n25020, n_18022, n25019);
  and g40039 (n25021, pi0608, n_17965);
  not g40040 (n_18026, n25020);
  and g40041 (n25022, n_18026, n25021);
  not g40042 (n_18027, n25018);
  not g40043 (n_18028, n25022);
  and g40044 (n25023, n_18027, n_18028);
  not g40045 (n_18029, n25023);
  and g40046 (n25024, pi0778, n_18029);
  and g40047 (n25025, n_11749, n_18023);
  not g40048 (n_18030, n25024);
  not g40049 (n_18031, n25025);
  and g40050 (n25026, n_18030, n_18031);
  not g40051 (n_18032, n25026);
  and g40052 (n25027, n_11971, n_18032);
  not g40053 (n_18033, n25011);
  and g40054 (n25028, n_11768, n_18033);
  not g40055 (n_18034, n25027);
  and g40056 (n25029, n_18034, n25028);
  and g40057 (n25030, n_11767, n_17976);
  not g40058 (n_18035, n25029);
  and g40059 (n25031, n_18035, n25030);
  and g40060 (n25032, n_11971, n24942);
  and g40061 (n25033, pi0609, n_18032);
  not g40062 (n_18036, n25032);
  and g40063 (n25034, pi1155, n_18036);
  not g40064 (n_18037, n25033);
  and g40065 (n25035, n_18037, n25034);
  and g40066 (n25036, pi0660, n_17977);
  not g40067 (n_18038, n25035);
  and g40068 (n25037, n_18038, n25036);
  not g40069 (n_18039, n25031);
  not g40070 (n_18040, n25037);
  and g40071 (n25038, n_18039, n_18040);
  not g40072 (n_18041, n25038);
  and g40073 (n25039, pi0785, n_18041);
  and g40074 (n25040, n_11964, n_18032);
  not g40075 (n_18042, n25039);
  not g40076 (n_18043, n25040);
  and g40077 (n25041, n_18042, n_18043);
  not g40078 (n_18044, n25041);
  and g40079 (n25042, n_11984, n_18044);
  not g40080 (n_18045, n25010);
  and g40081 (n25043, n_11413, n_18045);
  not g40082 (n_18046, n25042);
  and g40083 (n25044, n_18046, n25043);
  and g40084 (n25045, n_11412, n_17984);
  not g40085 (n_18047, n25044);
  and g40086 (n25046, n_18047, n25045);
  and g40087 (n25047, n_11984, n24943);
  and g40088 (n25048, pi0618, n_18044);
  not g40089 (n_18048, n25047);
  and g40090 (n25049, pi1154, n_18048);
  not g40091 (n_18049, n25048);
  and g40092 (n25050, n_18049, n25049);
  and g40093 (n25051, pi0627, n_17985);
  not g40094 (n_18050, n25050);
  and g40095 (n25052, n_18050, n25051);
  not g40096 (n_18051, n25046);
  not g40097 (n_18052, n25052);
  and g40098 (n25053, n_18051, n_18052);
  not g40099 (n_18053, n25053);
  and g40100 (n25054, pi0781, n_18053);
  and g40101 (n25055, n_11981, n_18044);
  not g40102 (n_18054, n25054);
  not g40103 (n_18055, n25055);
  and g40104 (n25056, n_18054, n_18055);
  and g40105 (n25057, n_12315, n25056);
  not g40106 (n_18056, n25056);
  and g40107 (n25058, n_11821, n_18056);
  and g40108 (n25059, pi0619, n24944);
  not g40109 (n_18057, n25059);
  and g40110 (n25060, n_11405, n_18057);
  not g40111 (n_18058, n25058);
  and g40112 (n25061, n_18058, n25060);
  and g40113 (n25062, n_11403, n_17994);
  not g40114 (n_18059, n25061);
  and g40115 (n25063, n_18059, n25062);
  and g40116 (n25064, pi0619, n_18056);
  and g40117 (n25065, n_11821, n24944);
  not g40118 (n_18060, n25065);
  and g40119 (n25066, pi1159, n_18060);
  not g40120 (n_18061, n25064);
  and g40121 (n25067, n_18061, n25066);
  and g40122 (n25068, pi0648, n_17995);
  not g40123 (n_18062, n25067);
  and g40124 (n25069, n_18062, n25068);
  not g40125 (n_18063, n25063);
  and g40126 (n25070, pi0789, n_18063);
  not g40127 (n_18064, n25069);
  and g40128 (n25071, n_18064, n25070);
  not g40129 (n_18065, n25057);
  and g40130 (n25072, n17970, n_18065);
  not g40131 (n_18066, n25071);
  and g40132 (n25073, n_18066, n25072);
  not g40133 (n_18067, n25009);
  not g40134 (n_18068, n25073);
  and g40135 (n25074, n_18067, n_18068);
  not g40136 (n_18069, n25074);
  and g40137 (n25075, n_14638, n_18069);
  and g40138 (n25076, n17854, n_18001);
  and g40139 (n25077, n20851, n24946);
  not g40140 (n_18070, n25076);
  not g40141 (n_18071, n25077);
  and g40142 (n25078, n_18070, n_18071);
  not g40143 (n_18072, n25078);
  and g40144 (n25079, n_12354, n_18072);
  and g40145 (n25080, n20855, n24946);
  and g40146 (n25081, n17853, n_18001);
  not g40147 (n_18073, n25080);
  not g40148 (n_18074, n25081);
  and g40149 (n25082, n_18073, n_18074);
  not g40150 (n_18075, n25082);
  and g40151 (n25083, pi0629, n_18075);
  not g40152 (n_18076, n25079);
  not g40153 (n_18077, n25083);
  and g40154 (n25084, n_18076, n_18077);
  not g40155 (n_18078, n25084);
  and g40156 (n25085, pi0792, n_18078);
  not g40157 (n_18079, n25085);
  and g40158 (n25086, n_14387, n_18079);
  not g40159 (n_18080, n25075);
  and g40160 (n25087, n_18080, n25086);
  not g40161 (n_18081, n24997);
  not g40162 (n_18082, n25087);
  and g40163 (n25088, n_18081, n_18082);
  and g40164 (n25089, n_12411, n25088);
  and g40165 (n25090, n_11803, n_18004);
  and g40166 (n25091, pi1157, n_18007);
  not g40167 (n_18083, n24951);
  not g40168 (n_18084, n25091);
  and g40169 (n25092, n_18083, n_18084);
  not g40170 (n_18085, n25092);
  and g40171 (n25093, pi0787, n_18085);
  not g40172 (n_18086, n25090);
  not g40173 (n_18087, n25093);
  and g40174 (n25094, n_18086, n_18087);
  and g40175 (n25095, n_11819, n25094);
  and g40176 (n25096, pi0644, n25088);
  not g40177 (n_18088, n25095);
  and g40178 (n25097, pi0715, n_18088);
  not g40179 (n_18089, n25096);
  and g40180 (n25098, n_18089, n25097);
  not g40181 (n_18090, n24989);
  and g40182 (n25099, n_12392, n_18090);
  and g40183 (n25100, n17804, n24931);
  not g40184 (n_18091, n25099);
  not g40185 (n_18092, n25100);
  and g40186 (n25101, n_18091, n_18092);
  not g40187 (n_18093, n25101);
  and g40188 (n25102, pi0644, n_18093);
  and g40189 (n25103, n_11819, n24931);
  not g40190 (n_18094, n25103);
  and g40191 (n25104, n_12395, n_18094);
  not g40192 (n_18095, n25102);
  and g40193 (n25105, n_18095, n25104);
  not g40194 (n_18096, n25105);
  and g40195 (n25106, pi1160, n_18096);
  not g40196 (n_18097, n25098);
  and g40197 (n25107, n_18097, n25106);
  and g40198 (n25108, n_11819, n_18093);
  and g40199 (n25109, pi0644, n24931);
  not g40200 (n_18098, n25109);
  and g40201 (n25110, pi0715, n_18098);
  not g40202 (n_18099, n25108);
  and g40203 (n25111, n_18099, n25110);
  and g40204 (n25112, pi0644, n25094);
  and g40205 (n25113, n_11819, n25088);
  not g40206 (n_18100, n25112);
  and g40207 (n25114, n_12395, n_18100);
  not g40208 (n_18101, n25113);
  and g40209 (n25115, n_18101, n25114);
  not g40210 (n_18102, n25111);
  and g40211 (n25116, n_12405, n_18102);
  not g40212 (n_18103, n25115);
  and g40213 (n25117, n_18103, n25116);
  not g40214 (n_18104, n25107);
  not g40215 (n_18105, n25117);
  and g40216 (n25118, n_18104, n_18105);
  not g40217 (n_18106, n25118);
  and g40218 (n25119, pi0790, n_18106);
  not g40219 (n_18107, n25089);
  and g40220 (n25120, pi0832, n_18107);
  not g40221 (n_18108, n25119);
  and g40222 (n25121, n_18108, n25120);
  not g40223 (n_18109, n24930);
  not g40224 (n_18110, n25121);
  and g40225 (po0334, n_18109, n_18110);
  and g40226 (n25123, n_5708, n_12418);
  and g40227 (n25124, n_15444, n16645);
  not g40228 (n_18111, n25123);
  not g40229 (n_18112, n25124);
  and g40230 (n25125, n_18111, n_18112);
  not g40231 (n_18113, n25125);
  and g40232 (n25126, n_11749, n_18113);
  and g40233 (n25127, n_11753, n25124);
  not g40234 (n_18114, n25127);
  and g40235 (n25128, n_18113, n_18114);
  not g40236 (n_18115, n25128);
  and g40237 (n25129, pi1153, n_18115);
  and g40238 (n25130, n_11757, n_18111);
  and g40239 (n25131, n_18114, n25130);
  not g40240 (n_18116, n25131);
  and g40241 (n25132, pi0778, n_18116);
  not g40242 (n_18117, n25129);
  and g40243 (n25133, n_18117, n25132);
  not g40244 (n_18118, n25126);
  not g40245 (n_18119, n25133);
  and g40246 (n25134, n_18118, n_18119);
  not g40247 (n_18120, n25134);
  and g40248 (n25135, n_12429, n_18120);
  and g40249 (n25136, n_12430, n25135);
  and g40250 (n25137, n_12431, n25136);
  and g40251 (n25138, n_12432, n25137);
  and g40252 (n25139, n_12436, n25138);
  and g40253 (n25140, n_11806, n25139);
  and g40254 (n25141, pi0647, n25123);
  not g40255 (n_18121, n25141);
  and g40256 (n25142, n_11810, n_18121);
  not g40257 (n_18122, n25140);
  and g40258 (n25143, n_18122, n25142);
  and g40259 (n25144, pi0630, n25143);
  and g40260 (n25145, n_15442, n17244);
  not g40261 (n_18123, n25145);
  and g40262 (n25146, n_18111, n_18123);
  not g40263 (n_18124, n25146);
  and g40264 (n25147, n_12448, n_18124);
  not g40265 (n_18125, n25147);
  and g40266 (n25148, n_11964, n_18125);
  and g40267 (n25149, n17296, n25145);
  not g40268 (n_18126, n25149);
  and g40269 (n25150, n25147, n_18126);
  not g40270 (n_18127, n25150);
  and g40271 (n25151, pi1155, n_18127);
  and g40272 (n25152, n_11768, n_18111);
  and g40273 (n25153, n_18126, n25152);
  not g40274 (n_18128, n25151);
  not g40275 (n_18129, n25153);
  and g40276 (n25154, n_18128, n_18129);
  not g40277 (n_18130, n25154);
  and g40278 (n25155, pi0785, n_18130);
  not g40279 (n_18131, n25148);
  not g40280 (n_18132, n25155);
  and g40281 (n25156, n_18131, n_18132);
  not g40282 (n_18133, n25156);
  and g40283 (n25157, n_11981, n_18133);
  and g40284 (n25158, n_12461, n25156);
  not g40285 (n_18134, n25158);
  and g40286 (n25159, pi1154, n_18134);
  and g40287 (n25160, n_12463, n25156);
  not g40288 (n_18135, n25160);
  and g40289 (n25161, n_11413, n_18135);
  not g40290 (n_18136, n25159);
  not g40291 (n_18137, n25161);
  and g40292 (n25162, n_18136, n_18137);
  not g40293 (n_18138, n25162);
  and g40294 (n25163, pi0781, n_18138);
  not g40295 (n_18139, n25157);
  not g40296 (n_18140, n25163);
  and g40297 (n25164, n_18139, n_18140);
  not g40298 (n_18141, n25164);
  and g40299 (n25165, n_12315, n_18141);
  and g40300 (n25166, n_16503, n25164);
  not g40301 (n_18142, n25166);
  and g40302 (n25167, pi1159, n_18142);
  and g40303 (n25168, n_16505, n25164);
  not g40304 (n_18143, n25168);
  and g40305 (n25169, n_11405, n_18143);
  not g40306 (n_18144, n25167);
  not g40307 (n_18145, n25169);
  and g40308 (n25170, n_18144, n_18145);
  not g40309 (n_18146, n25170);
  and g40310 (n25171, pi0789, n_18146);
  not g40311 (n_18147, n25165);
  not g40312 (n_18148, n25171);
  and g40313 (n25172, n_18147, n_18148);
  and g40314 (n25173, n_12524, n25172);
  and g40315 (n25174, n17969, n25123);
  not g40316 (n_18149, n25173);
  not g40317 (n_18150, n25174);
  and g40318 (n25175, n_18149, n_18150);
  not g40319 (n_18151, n25175);
  and g40320 (n25176, n_12368, n_18151);
  and g40321 (n25177, n17779, n25123);
  not g40322 (n_18152, n25176);
  not g40323 (n_18153, n25177);
  and g40324 (n25178, n_18152, n_18153);
  and g40325 (n25179, n_14548, n25178);
  not g40326 (n_18154, n25139);
  and g40327 (n25180, pi0647, n_18154);
  and g40328 (n25181, n_11806, n_18111);
  not g40329 (n_18155, n25180);
  not g40330 (n_18156, n25181);
  and g40331 (n25182, n_18155, n_18156);
  not g40332 (n_18157, n25182);
  and g40333 (n25183, n17801, n_18157);
  not g40334 (n_18158, n25144);
  not g40335 (n_18159, n25183);
  and g40336 (n25184, n_18158, n_18159);
  not g40337 (n_18160, n25179);
  and g40338 (n25185, n_18160, n25184);
  not g40339 (n_18161, n25185);
  and g40340 (n25186, pi0787, n_18161);
  and g40341 (n25187, n17871, n25137);
  not g40342 (n_18162, n25172);
  and g40343 (n25188, n_12320, n_18162);
  and g40344 (n25189, pi0626, n_18111);
  not g40345 (n_18163, n25189);
  and g40346 (n25190, n16629, n_18163);
  not g40347 (n_18164, n25188);
  and g40348 (n25191, n_18164, n25190);
  and g40349 (n25192, pi0626, n_18162);
  and g40350 (n25193, n_12320, n_18111);
  not g40351 (n_18165, n25193);
  and g40352 (n25194, n16628, n_18165);
  not g40353 (n_18166, n25192);
  and g40354 (n25195, n_18166, n25194);
  not g40355 (n_18167, n25187);
  not g40356 (n_18168, n25191);
  and g40357 (n25196, n_18167, n_18168);
  not g40358 (n_18169, n25195);
  and g40359 (n25197, n_18169, n25196);
  not g40360 (n_18170, n25197);
  and g40361 (n25198, pi0788, n_18170);
  and g40362 (n25199, pi0618, n25135);
  and g40363 (n25200, n_11866, n_18113);
  and g40364 (n25201, pi0625, n25200);
  not g40365 (n_18171, n25200);
  and g40366 (n25202, n25146, n_18171);
  not g40367 (n_18172, n25201);
  not g40368 (n_18173, n25202);
  and g40369 (n25203, n_18172, n_18173);
  not g40370 (n_18174, n25203);
  and g40371 (n25204, n25130, n_18174);
  and g40372 (n25205, n_11823, n_18117);
  not g40373 (n_18175, n25204);
  and g40374 (n25206, n_18175, n25205);
  and g40375 (n25207, pi1153, n25146);
  and g40376 (n25208, n_18172, n25207);
  and g40377 (n25209, pi0608, n_18116);
  not g40378 (n_18176, n25208);
  and g40379 (n25210, n_18176, n25209);
  not g40380 (n_18177, n25206);
  not g40381 (n_18178, n25210);
  and g40382 (n25211, n_18177, n_18178);
  not g40383 (n_18179, n25211);
  and g40384 (n25212, pi0778, n_18179);
  and g40385 (n25213, n_11749, n_18173);
  not g40386 (n_18180, n25212);
  not g40387 (n_18181, n25213);
  and g40388 (n25214, n_18180, n_18181);
  not g40389 (n_18182, n25214);
  and g40390 (n25215, n_11971, n_18182);
  and g40391 (n25216, pi0609, n_18120);
  not g40392 (n_18183, n25216);
  and g40393 (n25217, n_11768, n_18183);
  not g40394 (n_18184, n25215);
  and g40395 (n25218, n_18184, n25217);
  and g40396 (n25219, n_11767, n_18128);
  not g40397 (n_18185, n25218);
  and g40398 (n25220, n_18185, n25219);
  and g40399 (n25221, pi0609, n_18182);
  and g40400 (n25222, n_11971, n_18120);
  not g40401 (n_18186, n25222);
  and g40402 (n25223, pi1155, n_18186);
  not g40403 (n_18187, n25221);
  and g40404 (n25224, n_18187, n25223);
  and g40405 (n25225, pi0660, n_18129);
  not g40406 (n_18188, n25224);
  and g40407 (n25226, n_18188, n25225);
  not g40408 (n_18189, n25220);
  not g40409 (n_18190, n25226);
  and g40410 (n25227, n_18189, n_18190);
  not g40411 (n_18191, n25227);
  and g40412 (n25228, pi0785, n_18191);
  and g40413 (n25229, n_11964, n_18182);
  not g40414 (n_18192, n25228);
  not g40415 (n_18193, n25229);
  and g40416 (n25230, n_18192, n_18193);
  not g40417 (n_18194, n25230);
  and g40418 (n25231, n_11984, n_18194);
  not g40419 (n_18195, n25199);
  and g40420 (n25232, n_11413, n_18195);
  not g40421 (n_18196, n25231);
  and g40422 (n25233, n_18196, n25232);
  and g40423 (n25234, n_11412, n_18136);
  not g40424 (n_18197, n25233);
  and g40425 (n25235, n_18197, n25234);
  and g40426 (n25236, n_11984, n25135);
  and g40427 (n25237, pi0618, n_18194);
  not g40428 (n_18198, n25236);
  and g40429 (n25238, pi1154, n_18198);
  not g40430 (n_18199, n25237);
  and g40431 (n25239, n_18199, n25238);
  and g40432 (n25240, pi0627, n_18137);
  not g40433 (n_18200, n25239);
  and g40434 (n25241, n_18200, n25240);
  not g40435 (n_18201, n25235);
  not g40436 (n_18202, n25241);
  and g40437 (n25242, n_18201, n_18202);
  not g40438 (n_18203, n25242);
  and g40439 (n25243, pi0781, n_18203);
  and g40440 (n25244, n_11981, n_18194);
  not g40441 (n_18204, n25243);
  not g40442 (n_18205, n25244);
  and g40443 (n25245, n_18204, n_18205);
  and g40444 (n25246, n_12315, n25245);
  not g40445 (n_18206, n25245);
  and g40446 (n25247, n_11821, n_18206);
  and g40447 (n25248, pi0619, n25136);
  not g40448 (n_18207, n25248);
  and g40449 (n25249, n_11405, n_18207);
  not g40450 (n_18208, n25247);
  and g40451 (n25250, n_18208, n25249);
  and g40452 (n25251, n_11403, n_18144);
  not g40453 (n_18209, n25250);
  and g40454 (n25252, n_18209, n25251);
  and g40455 (n25253, pi0619, n_18206);
  and g40456 (n25254, n_11821, n25136);
  not g40457 (n_18210, n25254);
  and g40458 (n25255, pi1159, n_18210);
  not g40459 (n_18211, n25253);
  and g40460 (n25256, n_18211, n25255);
  and g40461 (n25257, pi0648, n_18145);
  not g40462 (n_18212, n25256);
  and g40463 (n25258, n_18212, n25257);
  not g40464 (n_18213, n25252);
  and g40465 (n25259, pi0789, n_18213);
  not g40466 (n_18214, n25258);
  and g40467 (n25260, n_18214, n25259);
  not g40468 (n_18215, n25246);
  and g40469 (n25261, n17970, n_18215);
  not g40470 (n_18216, n25260);
  and g40471 (n25262, n_18216, n25261);
  not g40472 (n_18217, n25198);
  not g40473 (n_18218, n25262);
  and g40474 (n25263, n_18217, n_18218);
  not g40475 (n_18219, n25263);
  and g40476 (n25264, n_14638, n_18219);
  and g40477 (n25265, n17854, n_18151);
  and g40478 (n25266, n20851, n25138);
  not g40479 (n_18220, n25265);
  not g40480 (n_18221, n25266);
  and g40481 (n25267, n_18220, n_18221);
  not g40482 (n_18222, n25267);
  and g40483 (n25268, n_12354, n_18222);
  and g40484 (n25269, n20855, n25138);
  and g40485 (n25270, n17853, n_18151);
  not g40486 (n_18223, n25269);
  not g40487 (n_18224, n25270);
  and g40488 (n25271, n_18223, n_18224);
  not g40489 (n_18225, n25271);
  and g40490 (n25272, pi0629, n_18225);
  not g40491 (n_18226, n25268);
  not g40492 (n_18227, n25272);
  and g40493 (n25273, n_18226, n_18227);
  not g40494 (n_18228, n25273);
  and g40495 (n25274, pi0792, n_18228);
  not g40496 (n_18229, n25274);
  and g40497 (n25275, n_14387, n_18229);
  not g40498 (n_18230, n25264);
  and g40499 (n25276, n_18230, n25275);
  not g40500 (n_18231, n25186);
  not g40501 (n_18232, n25276);
  and g40502 (n25277, n_18231, n_18232);
  and g40503 (n25278, n_12411, n25277);
  and g40504 (n25279, n_11803, n_18154);
  and g40505 (n25280, pi1157, n_18157);
  not g40506 (n_18233, n25143);
  not g40507 (n_18234, n25280);
  and g40508 (n25281, n_18233, n_18234);
  not g40509 (n_18235, n25281);
  and g40510 (n25282, pi0787, n_18235);
  not g40511 (n_18236, n25279);
  not g40512 (n_18237, n25282);
  and g40513 (n25283, n_18236, n_18237);
  and g40514 (n25284, n_11819, n25283);
  and g40515 (n25285, pi0644, n25277);
  not g40516 (n_18238, n25284);
  and g40517 (n25286, pi0715, n_18238);
  not g40518 (n_18239, n25285);
  and g40519 (n25287, n_18239, n25286);
  not g40520 (n_18240, n25178);
  and g40521 (n25288, n_12392, n_18240);
  and g40522 (n25289, n17804, n25123);
  not g40523 (n_18241, n25288);
  not g40524 (n_18242, n25289);
  and g40525 (n25290, n_18241, n_18242);
  not g40526 (n_18243, n25290);
  and g40527 (n25291, pi0644, n_18243);
  and g40528 (n25292, n_11819, n25123);
  not g40529 (n_18244, n25292);
  and g40530 (n25293, n_12395, n_18244);
  not g40531 (n_18245, n25291);
  and g40532 (n25294, n_18245, n25293);
  not g40533 (n_18246, n25294);
  and g40534 (n25295, pi1160, n_18246);
  not g40535 (n_18247, n25287);
  and g40536 (n25296, n_18247, n25295);
  and g40537 (n25297, n_11819, n_18243);
  and g40538 (n25298, pi0644, n25123);
  not g40539 (n_18248, n25298);
  and g40540 (n25299, pi0715, n_18248);
  not g40541 (n_18249, n25297);
  and g40542 (n25300, n_18249, n25299);
  and g40543 (n25301, pi0644, n25283);
  and g40544 (n25302, n_11819, n25277);
  not g40545 (n_18250, n25301);
  and g40546 (n25303, n_12395, n_18250);
  not g40547 (n_18251, n25302);
  and g40548 (n25304, n_18251, n25303);
  not g40549 (n_18252, n25300);
  and g40550 (n25305, n_12405, n_18252);
  not g40551 (n_18253, n25304);
  and g40552 (n25306, n_18253, n25305);
  not g40553 (n_18254, n25296);
  not g40554 (n_18255, n25306);
  and g40555 (n25307, n_18254, n_18255);
  not g40556 (n_18256, n25307);
  and g40557 (n25308, pi0790, n_18256);
  not g40558 (n_18257, n25278);
  and g40559 (n25309, pi0832, n_18257);
  not g40560 (n_18258, n25308);
  and g40561 (n25310, n_18258, n25309);
  and g40562 (n25311, n_5708, po1038);
  and g40563 (n25312, n_5708, n_11751);
  not g40564 (n_18259, n25312);
  and g40565 (n25313, n16635, n_18259);
  and g40566 (n25314, n_15444, n2571);
  not g40567 (n_18260, n25314);
  and g40568 (n25315, n25312, n_18260);
  and g40569 (n25316, n_5708, n_11418);
  not g40570 (n_18261, n25316);
  and g40571 (n25317, n16647, n_18261);
  and g40572 (n25318, pi0178, n_12608);
  not g40573 (n_18262, n25318);
  and g40574 (n25319, n_161, n_18262);
  not g40575 (n_18263, n25319);
  and g40576 (n25320, n2571, n_18263);
  and g40577 (n25321, n_5708, n18072);
  not g40578 (n_18264, n25320);
  not g40579 (n_18265, n25321);
  and g40580 (n25322, n_18264, n_18265);
  not g40581 (n_18266, n25317);
  and g40582 (n25323, n_15444, n_18266);
  not g40583 (n_18267, n25322);
  and g40584 (n25324, n_18267, n25323);
  not g40585 (n_18268, n25315);
  not g40586 (n_18269, n25324);
  and g40587 (n25325, n_18268, n_18269);
  and g40588 (n25326, n_11749, n25325);
  and g40589 (n25327, n_11753, n25312);
  not g40590 (n_18270, n25325);
  and g40591 (n25328, pi0625, n_18270);
  not g40592 (n_18271, n25327);
  and g40593 (n25329, pi1153, n_18271);
  not g40594 (n_18272, n25328);
  and g40595 (n25330, n_18272, n25329);
  and g40596 (n25331, pi0625, n25312);
  and g40597 (n25332, n_11753, n_18270);
  not g40598 (n_18273, n25331);
  and g40599 (n25333, n_11757, n_18273);
  not g40600 (n_18274, n25332);
  and g40601 (n25334, n_18274, n25333);
  not g40602 (n_18275, n25330);
  not g40603 (n_18276, n25334);
  and g40604 (n25335, n_18275, n_18276);
  not g40605 (n_18277, n25335);
  and g40606 (n25336, pi0778, n_18277);
  not g40607 (n_18278, n25326);
  not g40608 (n_18279, n25336);
  and g40609 (n25337, n_18278, n_18279);
  not g40610 (n_18280, n25337);
  and g40611 (n25338, n_11773, n_18280);
  and g40612 (n25339, n17075, n_18259);
  not g40613 (n_18281, n25338);
  not g40614 (n_18282, n25339);
  and g40615 (n25340, n_18281, n_18282);
  and g40616 (n25341, n_11777, n25340);
  and g40617 (n25342, n16639, n25312);
  not g40618 (n_18283, n25341);
  not g40619 (n_18284, n25342);
  and g40620 (n25343, n_18283, n_18284);
  and g40621 (n25344, n_11780, n25343);
  not g40622 (n_18285, n25313);
  not g40623 (n_18286, n25344);
  and g40624 (n25345, n_18285, n_18286);
  and g40625 (n25346, n_11783, n25345);
  and g40626 (n25347, n16631, n25312);
  not g40627 (n_18287, n25346);
  not g40628 (n_18288, n25347);
  and g40629 (n25348, n_18287, n_18288);
  and g40630 (n25349, n_11787, n25348);
  not g40631 (n_18289, n25348);
  and g40632 (n25350, pi0628, n_18289);
  and g40633 (n25351, n_11789, n25312);
  not g40634 (n_18290, n25351);
  and g40635 (n25352, pi1156, n_18290);
  not g40636 (n_18291, n25350);
  and g40637 (n25353, n_18291, n25352);
  and g40638 (n25354, pi0628, n25312);
  and g40639 (n25355, n_11789, n_18289);
  not g40640 (n_18292, n25354);
  and g40641 (n25356, n_11794, n_18292);
  not g40642 (n_18293, n25355);
  and g40643 (n25357, n_18293, n25356);
  not g40644 (n_18294, n25353);
  not g40645 (n_18295, n25357);
  and g40646 (n25358, n_18294, n_18295);
  not g40647 (n_18296, n25358);
  and g40648 (n25359, pi0792, n_18296);
  not g40649 (n_18297, n25349);
  not g40650 (n_18298, n25359);
  and g40651 (n25360, n_18297, n_18298);
  not g40652 (n_18299, n25360);
  and g40653 (n25361, n_11806, n_18299);
  and g40654 (n25362, pi0647, n_18259);
  not g40655 (n_18300, n25361);
  not g40656 (n_18301, n25362);
  and g40657 (n25363, n_18300, n_18301);
  and g40658 (n25364, n_11810, n25363);
  and g40659 (n25365, pi0647, n_18299);
  and g40660 (n25366, n_11806, n_18259);
  not g40661 (n_18302, n25365);
  not g40662 (n_18303, n25366);
  and g40663 (n25367, n_18302, n_18303);
  and g40664 (n25368, pi1157, n25367);
  not g40665 (n_18304, n25364);
  not g40666 (n_18305, n25368);
  and g40667 (n25369, n_18304, n_18305);
  not g40668 (n_18306, n25369);
  and g40669 (n25370, pi0787, n_18306);
  and g40670 (n25371, n_11803, n25360);
  not g40671 (n_18307, n25370);
  not g40672 (n_18308, n25371);
  and g40673 (n25372, n_18307, n_18308);
  not g40674 (n_18309, n25372);
  and g40675 (n25373, n_11819, n_18309);
  not g40676 (n_18310, n25373);
  and g40677 (n25374, pi0715, n_18310);
  and g40678 (n25375, pi0178, n_11417);
  and g40679 (n25376, n_15442, n17280);
  not g40680 (n_18311, n25376);
  and g40681 (n25377, n_18261, n_18311);
  not g40682 (n_18312, n25377);
  and g40683 (n25378, pi0038, n_18312);
  and g40684 (n25379, n_5708, n17221);
  and g40685 (n25380, pi0178, n_14476);
  not g40686 (n_18313, n25380);
  and g40687 (n25381, n_15442, n_18313);
  not g40688 (n_18314, n25379);
  and g40689 (n25382, n_18314, n25381);
  and g40690 (n25383, n_5708, pi0760);
  and g40691 (n25384, n_11739, n25383);
  not g40692 (n_18315, n25382);
  not g40693 (n_18316, n25384);
  and g40694 (n25385, n_18315, n_18316);
  not g40695 (n_18317, n25385);
  and g40696 (n25386, n_161, n_18317);
  not g40697 (n_18318, n25378);
  not g40698 (n_18319, n25386);
  and g40699 (n25387, n_18318, n_18319);
  and g40700 (n25388, n2571, n25387);
  not g40701 (n_18320, n25375);
  not g40702 (n_18321, n25388);
  and g40703 (n25389, n_18320, n_18321);
  not g40704 (n_18322, n25389);
  and g40705 (n25390, n_11960, n_18322);
  and g40706 (n25391, n17117, n_18259);
  not g40707 (n_18323, n25390);
  not g40708 (n_18324, n25391);
  and g40709 (n25392, n_18323, n_18324);
  not g40710 (n_18325, n25392);
  and g40711 (n25393, n_11964, n_18325);
  and g40712 (n25394, n_11967, n_18259);
  and g40713 (n25395, pi0609, n25390);
  not g40714 (n_18326, n25394);
  not g40715 (n_18327, n25395);
  and g40716 (n25396, n_18326, n_18327);
  not g40717 (n_18328, n25396);
  and g40718 (n25397, pi1155, n_18328);
  and g40719 (n25398, n_11972, n_18259);
  and g40720 (n25399, n_11971, n25390);
  not g40721 (n_18329, n25398);
  not g40722 (n_18330, n25399);
  and g40723 (n25400, n_18329, n_18330);
  not g40724 (n_18331, n25400);
  and g40725 (n25401, n_11768, n_18331);
  not g40726 (n_18332, n25397);
  not g40727 (n_18333, n25401);
  and g40728 (n25402, n_18332, n_18333);
  not g40729 (n_18334, n25402);
  and g40730 (n25403, pi0785, n_18334);
  not g40731 (n_18335, n25393);
  not g40732 (n_18336, n25403);
  and g40733 (n25404, n_18335, n_18336);
  not g40734 (n_18337, n25404);
  and g40735 (n25405, n_11981, n_18337);
  and g40736 (n25406, n_11984, n25312);
  and g40737 (n25407, pi0618, n25404);
  not g40738 (n_18338, n25406);
  and g40739 (n25408, pi1154, n_18338);
  not g40740 (n_18339, n25407);
  and g40741 (n25409, n_18339, n25408);
  and g40742 (n25410, n_11984, n25404);
  and g40743 (n25411, pi0618, n25312);
  not g40744 (n_18340, n25411);
  and g40745 (n25412, n_11413, n_18340);
  not g40746 (n_18341, n25410);
  and g40747 (n25413, n_18341, n25412);
  not g40748 (n_18342, n25409);
  not g40749 (n_18343, n25413);
  and g40750 (n25414, n_18342, n_18343);
  not g40751 (n_18344, n25414);
  and g40752 (n25415, pi0781, n_18344);
  not g40753 (n_18345, n25405);
  not g40754 (n_18346, n25415);
  and g40755 (n25416, n_18345, n_18346);
  not g40756 (n_18347, n25416);
  and g40757 (n25417, n_12315, n_18347);
  and g40758 (n25418, n_11821, n25312);
  and g40759 (n25419, pi0619, n25416);
  not g40760 (n_18348, n25418);
  and g40761 (n25420, pi1159, n_18348);
  not g40762 (n_18349, n25419);
  and g40763 (n25421, n_18349, n25420);
  and g40764 (n25422, n_11821, n25416);
  and g40765 (n25423, pi0619, n25312);
  not g40766 (n_18350, n25423);
  and g40767 (n25424, n_11405, n_18350);
  not g40768 (n_18351, n25422);
  and g40769 (n25425, n_18351, n25424);
  not g40770 (n_18352, n25421);
  not g40771 (n_18353, n25425);
  and g40772 (n25426, n_18352, n_18353);
  not g40773 (n_18354, n25426);
  and g40774 (n25427, pi0789, n_18354);
  not g40775 (n_18355, n25417);
  not g40776 (n_18356, n25427);
  and g40777 (n25428, n_18355, n_18356);
  and g40778 (n25429, n_12524, n25428);
  and g40779 (n25430, n17969, n25312);
  not g40780 (n_18357, n25429);
  not g40781 (n_18358, n25430);
  and g40782 (n25431, n_18357, n_18358);
  not g40783 (n_18359, n25431);
  and g40784 (n25432, n_12368, n_18359);
  and g40785 (n25433, n17779, n25312);
  not g40786 (n_18360, n25432);
  not g40787 (n_18361, n25433);
  and g40788 (n25434, n_18360, n_18361);
  not g40789 (n_18362, n25434);
  and g40790 (n25435, n_12392, n_18362);
  and g40791 (n25436, n17804, n25312);
  not g40792 (n_18363, n25435);
  not g40793 (n_18364, n25436);
  and g40794 (n25437, n_18363, n_18364);
  not g40795 (n_18365, n25437);
  and g40796 (n25438, pi0644, n_18365);
  and g40797 (n25439, n_11819, n25312);
  not g40798 (n_18366, n25439);
  and g40799 (n25440, n_12395, n_18366);
  not g40800 (n_18367, n25438);
  and g40801 (n25441, n_18367, n25440);
  not g40802 (n_18368, n25441);
  and g40803 (n25442, pi1160, n_18368);
  not g40804 (n_18369, n25374);
  and g40805 (n25443, n_18369, n25442);
  and g40806 (n25444, pi0644, n_18309);
  not g40807 (n_18370, n25444);
  and g40808 (n25445, n_12395, n_18370);
  and g40809 (n25446, n_11819, n_18365);
  and g40810 (n25447, pi0644, n25312);
  not g40811 (n_18371, n25447);
  and g40812 (n25448, pi0715, n_18371);
  not g40813 (n_18372, n25446);
  and g40814 (n25449, n_18372, n25448);
  not g40815 (n_18373, n25449);
  and g40816 (n25450, n_12405, n_18373);
  not g40817 (n_18374, n25445);
  and g40818 (n25451, n_18374, n25450);
  not g40819 (n_18375, n25443);
  not g40820 (n_18376, n25451);
  and g40821 (n25452, n_18375, n_18376);
  not g40822 (n_18377, n25452);
  and g40823 (n25453, pi0790, n_18377);
  and g40824 (n25454, n_12354, n25353);
  and g40825 (n25455, n_14557, n25431);
  and g40826 (n25456, pi0629, n25357);
  not g40827 (n_18378, n25454);
  not g40828 (n_18379, n25456);
  and g40829 (n25457, n_18378, n_18379);
  not g40830 (n_18380, n25455);
  and g40831 (n25458, n_18380, n25457);
  not g40832 (n_18381, n25458);
  and g40833 (n25459, pi0792, n_18381);
  and g40834 (n25460, pi0609, n25337);
  and g40835 (n25461, pi0178, n_12240);
  and g40836 (n25462, n_5708, n_12230);
  not g40837 (n_18382, n25461);
  and g40838 (n25463, pi0760, n_18382);
  not g40839 (n_18383, n25462);
  and g40840 (n25464, n_18383, n25463);
  and g40841 (n25465, n_5708, n17629);
  and g40842 (n25466, pi0178, n17631);
  not g40843 (n_18384, n25466);
  and g40844 (n25467, n_15442, n_18384);
  not g40845 (n_18385, n25465);
  and g40846 (n25468, n_18385, n25467);
  not g40847 (n_18386, n25464);
  not g40848 (n_18387, n25468);
  and g40849 (n25469, n_18386, n_18387);
  not g40850 (n_18388, n25469);
  and g40851 (n25470, n_162, n_18388);
  and g40852 (n25471, pi0178, n17605);
  and g40853 (n25472, n_5708, n_12180);
  not g40854 (n_18389, n25472);
  and g40855 (n25473, n_15442, n_18389);
  not g40856 (n_18390, n25471);
  and g40857 (n25474, n_18390, n25473);
  and g40858 (n25475, n_5708, n17404);
  and g40859 (n25476, pi0178, n17485);
  not g40860 (n_18391, n25476);
  and g40861 (n25477, pi0760, n_18391);
  not g40862 (n_18392, n25475);
  and g40863 (n25478, n_18392, n25477);
  not g40864 (n_18393, n25474);
  and g40865 (n25479, pi0039, n_18393);
  not g40866 (n_18394, n25478);
  and g40867 (n25480, n_18394, n25479);
  not g40868 (n_18395, n25470);
  and g40869 (n25481, n_161, n_18395);
  not g40870 (n_18396, n25480);
  and g40871 (n25482, n_18396, n25481);
  and g40872 (n25483, n_15442, n_12250);
  not g40873 (n_18397, n25483);
  and g40874 (n25484, n19471, n_18397);
  not g40875 (n_18398, n25484);
  and g40876 (n25485, n_5708, n_18398);
  and g40877 (n25486, n_12120, n_18123);
  not g40878 (n_18399, n25486);
  and g40879 (n25487, pi0178, n_18399);
  and g40880 (n25488, n6284, n25487);
  not g40881 (n_18400, n25488);
  and g40882 (n25489, pi0038, n_18400);
  not g40883 (n_18401, n25485);
  and g40884 (n25490, n_18401, n25489);
  not g40885 (n_18402, n25490);
  and g40886 (n25491, n_15444, n_18402);
  not g40887 (n_18403, n25482);
  and g40888 (n25492, n_18403, n25491);
  not g40889 (n_18404, n25387);
  and g40890 (n25493, pi0688, n_18404);
  not g40891 (n_18405, n25492);
  and g40892 (n25494, n2571, n_18405);
  not g40893 (n_18406, n25493);
  and g40894 (n25495, n_18406, n25494);
  not g40895 (n_18407, n25495);
  and g40896 (n25496, n_18320, n_18407);
  and g40897 (n25497, n_11753, n25496);
  and g40898 (n25498, pi0625, n25389);
  not g40899 (n_18408, n25498);
  and g40900 (n25499, n_11757, n_18408);
  not g40901 (n_18409, n25497);
  and g40902 (n25500, n_18409, n25499);
  and g40903 (n25501, n_11823, n_18275);
  not g40904 (n_18410, n25500);
  and g40905 (n25502, n_18410, n25501);
  and g40906 (n25503, n_11753, n25389);
  and g40907 (n25504, pi0625, n25496);
  not g40908 (n_18411, n25503);
  and g40909 (n25505, pi1153, n_18411);
  not g40910 (n_18412, n25504);
  and g40911 (n25506, n_18412, n25505);
  and g40912 (n25507, pi0608, n_18276);
  not g40913 (n_18413, n25506);
  and g40914 (n25508, n_18413, n25507);
  not g40915 (n_18414, n25502);
  not g40916 (n_18415, n25508);
  and g40917 (n25509, n_18414, n_18415);
  not g40918 (n_18416, n25509);
  and g40919 (n25510, pi0778, n_18416);
  and g40920 (n25511, n_11749, n25496);
  not g40921 (n_18417, n25510);
  not g40922 (n_18418, n25511);
  and g40923 (n25512, n_18417, n_18418);
  not g40924 (n_18419, n25512);
  and g40925 (n25513, n_11971, n_18419);
  not g40926 (n_18420, n25460);
  and g40927 (n25514, n_11768, n_18420);
  not g40928 (n_18421, n25513);
  and g40929 (n25515, n_18421, n25514);
  and g40930 (n25516, n_11767, n_18332);
  not g40931 (n_18422, n25515);
  and g40932 (n25517, n_18422, n25516);
  and g40933 (n25518, n_11971, n25337);
  and g40934 (n25519, pi0609, n_18419);
  not g40935 (n_18423, n25518);
  and g40936 (n25520, pi1155, n_18423);
  not g40937 (n_18424, n25519);
  and g40938 (n25521, n_18424, n25520);
  and g40939 (n25522, pi0660, n_18333);
  not g40940 (n_18425, n25521);
  and g40941 (n25523, n_18425, n25522);
  not g40942 (n_18426, n25517);
  not g40943 (n_18427, n25523);
  and g40944 (n25524, n_18426, n_18427);
  not g40945 (n_18428, n25524);
  and g40946 (n25525, pi0785, n_18428);
  and g40947 (n25526, n_11964, n_18419);
  not g40948 (n_18429, n25525);
  not g40949 (n_18430, n25526);
  and g40950 (n25527, n_18429, n_18430);
  not g40951 (n_18431, n25527);
  and g40952 (n25528, n_11984, n_18431);
  and g40953 (n25529, pi0618, n25340);
  not g40954 (n_18432, n25529);
  and g40955 (n25530, n_11413, n_18432);
  not g40956 (n_18433, n25528);
  and g40957 (n25531, n_18433, n25530);
  and g40958 (n25532, n_11412, n_18342);
  not g40959 (n_18434, n25531);
  and g40960 (n25533, n_18434, n25532);
  and g40961 (n25534, n_11984, n25340);
  and g40962 (n25535, pi0618, n_18431);
  not g40963 (n_18435, n25534);
  and g40964 (n25536, pi1154, n_18435);
  not g40965 (n_18436, n25535);
  and g40966 (n25537, n_18436, n25536);
  and g40967 (n25538, pi0627, n_18343);
  not g40968 (n_18437, n25537);
  and g40969 (n25539, n_18437, n25538);
  not g40970 (n_18438, n25533);
  not g40971 (n_18439, n25539);
  and g40972 (n25540, n_18438, n_18439);
  not g40973 (n_18440, n25540);
  and g40974 (n25541, pi0781, n_18440);
  and g40975 (n25542, n_11981, n_18431);
  not g40976 (n_18441, n25541);
  not g40977 (n_18442, n25542);
  and g40978 (n25543, n_18441, n_18442);
  and g40979 (n25544, n_12315, n25543);
  not g40980 (n_18443, n25343);
  and g40981 (n25545, pi0619, n_18443);
  not g40982 (n_18444, n25543);
  and g40983 (n25546, n_11821, n_18444);
  not g40984 (n_18445, n25545);
  and g40985 (n25547, n_11405, n_18445);
  not g40986 (n_18446, n25546);
  and g40987 (n25548, n_18446, n25547);
  and g40988 (n25549, n_11403, n_18352);
  not g40989 (n_18447, n25548);
  and g40990 (n25550, n_18447, n25549);
  and g40991 (n25551, n_11821, n_18443);
  and g40992 (n25552, pi0619, n_18444);
  not g40993 (n_18448, n25551);
  and g40994 (n25553, pi1159, n_18448);
  not g40995 (n_18449, n25552);
  and g40996 (n25554, n_18449, n25553);
  and g40997 (n25555, pi0648, n_18353);
  not g40998 (n_18450, n25554);
  and g40999 (n25556, n_18450, n25555);
  not g41000 (n_18451, n25550);
  and g41001 (n25557, pi0789, n_18451);
  not g41002 (n_18452, n25556);
  and g41003 (n25558, n_18452, n25557);
  not g41004 (n_18453, n25544);
  and g41005 (n25559, n17970, n_18453);
  not g41006 (n_18454, n25558);
  and g41007 (n25560, n_18454, n25559);
  and g41008 (n25561, n17871, n25345);
  not g41009 (n_18455, n25428);
  and g41010 (n25562, n_12320, n_18455);
  and g41011 (n25563, pi0626, n_18259);
  not g41012 (n_18456, n25563);
  and g41013 (n25564, n16629, n_18456);
  not g41014 (n_18457, n25562);
  and g41015 (n25565, n_18457, n25564);
  and g41016 (n25566, pi0626, n_18455);
  and g41017 (n25567, n_12320, n_18259);
  not g41018 (n_18458, n25567);
  and g41019 (n25568, n16628, n_18458);
  not g41020 (n_18459, n25566);
  and g41021 (n25569, n_18459, n25568);
  not g41022 (n_18460, n25561);
  not g41023 (n_18461, n25565);
  and g41024 (n25570, n_18460, n_18461);
  not g41025 (n_18462, n25569);
  and g41026 (n25571, n_18462, n25570);
  not g41027 (n_18463, n25571);
  and g41028 (n25572, pi0788, n_18463);
  not g41029 (n_18464, n25572);
  and g41030 (n25573, n_14638, n_18464);
  not g41031 (n_18465, n25560);
  and g41032 (n25574, n_18465, n25573);
  not g41033 (n_18466, n25459);
  not g41034 (n_18467, n25574);
  and g41035 (n25575, n_18466, n_18467);
  not g41036 (n_18468, n25575);
  and g41037 (n25576, n_14387, n_18468);
  not g41038 (n_18469, n25363);
  and g41039 (n25577, n17802, n_18469);
  and g41040 (n25578, n_14548, n25434);
  not g41041 (n_18470, n25367);
  and g41042 (n25579, n17801, n_18470);
  not g41043 (n_18471, n25577);
  not g41044 (n_18472, n25579);
  and g41045 (n25580, n_18471, n_18472);
  not g41046 (n_18473, n25578);
  and g41047 (n25581, n_18473, n25580);
  not g41048 (n_18474, n25581);
  and g41049 (n25582, pi0787, n_18474);
  and g41050 (n25583, n_11819, n25450);
  and g41051 (n25584, pi0644, n25442);
  not g41052 (n_18475, n25583);
  and g41053 (n25585, pi0790, n_18475);
  not g41054 (n_18476, n25584);
  and g41055 (n25586, n_18476, n25585);
  not g41056 (n_18477, n25576);
  not g41057 (n_18478, n25582);
  and g41058 (n25587, n_18477, n_18478);
  not g41059 (n_18479, n25586);
  and g41060 (n25588, n_18479, n25587);
  not g41061 (n_18480, n25453);
  not g41062 (n_18481, n25588);
  and g41063 (n25589, n_18480, n_18481);
  not g41064 (n_18482, n25589);
  and g41065 (n25590, n_4226, n_18482);
  not g41066 (n_18483, n25311);
  and g41067 (n25591, n_12415, n_18483);
  not g41068 (n_18484, n25590);
  and g41069 (n25592, n_18484, n25591);
  not g41070 (n_18485, n25310);
  not g41071 (n_18486, n25592);
  and g41072 (po0335, n_18485, n_18486);
  and g41073 (n25594, n_7636, n_11751);
  not g41074 (n_18487, n25594);
  and g41075 (n25595, n16635, n_18487);
  and g41076 (n25596, n_15414, n2571);
  not g41077 (n_18488, n25596);
  and g41078 (n25597, n25594, n_18488);
  and g41079 (n25598, n_7636, n_11418);
  not g41080 (n_18489, n25598);
  and g41081 (n25599, n16647, n_18489);
  and g41082 (n25600, n_7636, n18072);
  and g41083 (n25601, pi0179, n_12608);
  not g41084 (n_18490, n25601);
  and g41085 (n25602, n_161, n_18490);
  not g41086 (n_18491, n25602);
  and g41087 (n25603, n2571, n_18491);
  not g41088 (n_18492, n25600);
  not g41089 (n_18493, n25603);
  and g41090 (n25604, n_18492, n_18493);
  not g41091 (n_18494, n25599);
  and g41092 (n25605, n_15414, n_18494);
  not g41093 (n_18495, n25604);
  and g41094 (n25606, n_18495, n25605);
  not g41095 (n_18496, n25597);
  not g41096 (n_18497, n25606);
  and g41097 (n25607, n_18496, n_18497);
  and g41098 (n25608, n_11749, n25607);
  and g41099 (n25609, n_11753, n25594);
  not g41100 (n_18498, n25607);
  and g41101 (n25610, pi0625, n_18498);
  not g41102 (n_18499, n25609);
  and g41103 (n25611, pi1153, n_18499);
  not g41104 (n_18500, n25610);
  and g41105 (n25612, n_18500, n25611);
  and g41106 (n25613, pi0625, n25594);
  and g41107 (n25614, n_11753, n_18498);
  not g41108 (n_18501, n25613);
  and g41109 (n25615, n_11757, n_18501);
  not g41110 (n_18502, n25614);
  and g41111 (n25616, n_18502, n25615);
  not g41112 (n_18503, n25612);
  not g41113 (n_18504, n25616);
  and g41114 (n25617, n_18503, n_18504);
  not g41115 (n_18505, n25617);
  and g41116 (n25618, pi0778, n_18505);
  not g41117 (n_18506, n25608);
  not g41118 (n_18507, n25618);
  and g41119 (n25619, n_18506, n_18507);
  not g41120 (n_18508, n25619);
  and g41121 (n25620, n_11773, n_18508);
  and g41122 (n25621, n17075, n_18487);
  not g41123 (n_18509, n25620);
  not g41124 (n_18510, n25621);
  and g41125 (n25622, n_18509, n_18510);
  and g41126 (n25623, n_11777, n25622);
  and g41127 (n25624, n16639, n25594);
  not g41128 (n_18511, n25623);
  not g41129 (n_18512, n25624);
  and g41130 (n25625, n_18511, n_18512);
  and g41131 (n25626, n_11780, n25625);
  not g41132 (n_18513, n25595);
  not g41133 (n_18514, n25626);
  and g41134 (n25627, n_18513, n_18514);
  and g41135 (n25628, n_11783, n25627);
  and g41136 (n25629, n16631, n25594);
  not g41137 (n_18515, n25628);
  not g41138 (n_18516, n25629);
  and g41139 (n25630, n_18515, n_18516);
  and g41140 (n25631, n_11787, n25630);
  and g41141 (n25632, n_11789, n25594);
  not g41142 (n_18517, n25630);
  and g41143 (n25633, pi0628, n_18517);
  not g41144 (n_18518, n25632);
  and g41145 (n25634, pi1156, n_18518);
  not g41146 (n_18519, n25633);
  and g41147 (n25635, n_18519, n25634);
  and g41148 (n25636, pi0628, n25594);
  and g41149 (n25637, n_11789, n_18517);
  not g41150 (n_18520, n25636);
  and g41151 (n25638, n_11794, n_18520);
  not g41152 (n_18521, n25637);
  and g41153 (n25639, n_18521, n25638);
  not g41154 (n_18522, n25635);
  not g41155 (n_18523, n25639);
  and g41156 (n25640, n_18522, n_18523);
  not g41157 (n_18524, n25640);
  and g41158 (n25641, pi0792, n_18524);
  not g41159 (n_18525, n25631);
  not g41160 (n_18526, n25641);
  and g41161 (n25642, n_18525, n_18526);
  not g41162 (n_18527, n25642);
  and g41163 (n25643, n_11803, n_18527);
  and g41164 (n25644, n_11806, n25594);
  and g41165 (n25645, pi0647, n25642);
  not g41166 (n_18528, n25644);
  and g41167 (n25646, pi1157, n_18528);
  not g41168 (n_18529, n25645);
  and g41169 (n25647, n_18529, n25646);
  and g41170 (n25648, n_11806, n25642);
  and g41171 (n25649, pi0647, n25594);
  not g41172 (n_18530, n25649);
  and g41173 (n25650, n_11810, n_18530);
  not g41174 (n_18531, n25648);
  and g41175 (n25651, n_18531, n25650);
  not g41176 (n_18532, n25647);
  not g41177 (n_18533, n25651);
  and g41178 (n25652, n_18532, n_18533);
  not g41179 (n_18534, n25652);
  and g41180 (n25653, pi0787, n_18534);
  not g41181 (n_18535, n25643);
  not g41182 (n_18536, n25653);
  and g41183 (n25654, n_18535, n_18536);
  and g41184 (n25655, n_11819, n25654);
  and g41185 (n25656, n_11984, n25594);
  and g41186 (n25657, pi0179, n_11417);
  and g41187 (n25658, n_15412, n_17784);
  not g41188 (n_18537, n25658);
  and g41189 (n25659, pi0179, n_18537);
  not g41193 (n_18538, n25659);
  not g41194 (n_18539, n25662);
  and g41195 (n25663, n_18538, n_18539);
  and g41196 (n25664, n_15425, n25663);
  not g41197 (n_18540, n25664);
  and g41198 (n25665, n2571, n_18540);
  not g41199 (n_18541, n25657);
  not g41200 (n_18542, n25665);
  and g41201 (n25666, n_18541, n_18542);
  not g41202 (n_18543, n25666);
  and g41203 (n25667, n_11960, n_18543);
  and g41204 (n25668, n17117, n_18487);
  not g41205 (n_18544, n25667);
  not g41206 (n_18545, n25668);
  and g41207 (n25669, n_18544, n_18545);
  not g41208 (n_18546, n25669);
  and g41209 (n25670, n_11964, n_18546);
  and g41210 (n25671, n_11967, n_18487);
  and g41211 (n25672, pi0609, n25667);
  not g41212 (n_18547, n25671);
  not g41213 (n_18548, n25672);
  and g41214 (n25673, n_18547, n_18548);
  not g41215 (n_18549, n25673);
  and g41216 (n25674, pi1155, n_18549);
  and g41217 (n25675, n_11972, n_18487);
  and g41218 (n25676, n_11971, n25667);
  not g41219 (n_18550, n25675);
  not g41220 (n_18551, n25676);
  and g41221 (n25677, n_18550, n_18551);
  not g41222 (n_18552, n25677);
  and g41223 (n25678, n_11768, n_18552);
  not g41224 (n_18553, n25674);
  not g41225 (n_18554, n25678);
  and g41226 (n25679, n_18553, n_18554);
  not g41227 (n_18555, n25679);
  and g41228 (n25680, pi0785, n_18555);
  not g41229 (n_18556, n25670);
  not g41230 (n_18557, n25680);
  and g41231 (n25681, n_18556, n_18557);
  and g41232 (n25682, pi0618, n25681);
  not g41233 (n_18558, n25656);
  and g41234 (n25683, pi1154, n_18558);
  not g41235 (n_18559, n25682);
  and g41236 (n25684, n_18559, n25683);
  and g41237 (n25685, n18176, n_18489);
  and g41238 (n25686, n_7636, n17404);
  and g41239 (n25687, pi0179, n17485);
  not g41240 (n_18560, n25687);
  and g41241 (n25688, pi0039, n_18560);
  not g41242 (n_18561, n25686);
  and g41243 (n25689, n_18561, n25688);
  and g41244 (n25690, n_7636, n17612);
  and g41245 (n25691, pi0179, n17625);
  not g41246 (n_18562, n25690);
  and g41247 (n25692, n_162, n_18562);
  not g41248 (n_18563, n25691);
  and g41249 (n25693, n_18563, n25692);
  not g41250 (n_18564, n25689);
  not g41251 (n_18565, n25693);
  and g41252 (n25694, n_18564, n_18565);
  not g41253 (n_18566, n25694);
  and g41254 (n25695, n_161, n_18566);
  not g41255 (n_18567, n25685);
  not g41256 (n_18568, n25695);
  and g41257 (n25696, n_18567, n_18568);
  not g41258 (n_18569, n25696);
  and g41259 (n25697, pi0741, n_18569);
  and g41260 (n25698, n_7636, n_13718);
  and g41261 (n25699, pi0179, n19496);
  not g41262 (n_18570, n25698);
  and g41263 (n25700, n_15412, n_18570);
  not g41264 (n_18571, n25699);
  and g41265 (n25701, n_18571, n25700);
  not g41266 (n_18572, n25701);
  and g41267 (n25702, n_15414, n_18572);
  not g41268 (n_18573, n25697);
  and g41269 (n25703, n_18573, n25702);
  and g41270 (n25704, pi0724, n25664);
  not g41271 (n_18574, n25704);
  and g41272 (n25705, n2571, n_18574);
  not g41273 (n_18575, n25703);
  and g41274 (n25706, n_18575, n25705);
  not g41275 (n_18576, n25706);
  and g41276 (n25707, n_18541, n_18576);
  and g41277 (n25708, n_11753, n25707);
  and g41278 (n25709, pi0625, n25666);
  not g41279 (n_18577, n25709);
  and g41280 (n25710, n_11757, n_18577);
  not g41281 (n_18578, n25708);
  and g41282 (n25711, n_18578, n25710);
  and g41283 (n25712, n_11823, n_18503);
  not g41284 (n_18579, n25711);
  and g41285 (n25713, n_18579, n25712);
  and g41286 (n25714, n_11753, n25666);
  and g41287 (n25715, pi0625, n25707);
  not g41288 (n_18580, n25714);
  and g41289 (n25716, pi1153, n_18580);
  not g41290 (n_18581, n25715);
  and g41291 (n25717, n_18581, n25716);
  and g41292 (n25718, pi0608, n_18504);
  not g41293 (n_18582, n25717);
  and g41294 (n25719, n_18582, n25718);
  not g41295 (n_18583, n25713);
  not g41296 (n_18584, n25719);
  and g41297 (n25720, n_18583, n_18584);
  not g41298 (n_18585, n25720);
  and g41299 (n25721, pi0778, n_18585);
  and g41300 (n25722, n_11749, n25707);
  not g41301 (n_18586, n25721);
  not g41302 (n_18587, n25722);
  and g41303 (n25723, n_18586, n_18587);
  not g41304 (n_18588, n25723);
  and g41305 (n25724, n_11971, n_18588);
  and g41306 (n25725, pi0609, n25619);
  not g41307 (n_18589, n25725);
  and g41308 (n25726, n_11768, n_18589);
  not g41309 (n_18590, n25724);
  and g41310 (n25727, n_18590, n25726);
  and g41311 (n25728, n_11767, n_18553);
  not g41312 (n_18591, n25727);
  and g41313 (n25729, n_18591, n25728);
  and g41314 (n25730, n_11971, n25619);
  and g41315 (n25731, pi0609, n_18588);
  not g41316 (n_18592, n25730);
  and g41317 (n25732, pi1155, n_18592);
  not g41318 (n_18593, n25731);
  and g41319 (n25733, n_18593, n25732);
  and g41320 (n25734, pi0660, n_18554);
  not g41321 (n_18594, n25733);
  and g41322 (n25735, n_18594, n25734);
  not g41323 (n_18595, n25729);
  not g41324 (n_18596, n25735);
  and g41325 (n25736, n_18595, n_18596);
  not g41326 (n_18597, n25736);
  and g41327 (n25737, pi0785, n_18597);
  and g41328 (n25738, n_11964, n_18588);
  not g41329 (n_18598, n25737);
  not g41330 (n_18599, n25738);
  and g41331 (n25739, n_18598, n_18599);
  not g41332 (n_18600, n25739);
  and g41333 (n25740, n_11984, n_18600);
  and g41334 (n25741, pi0618, n25622);
  not g41335 (n_18601, n25741);
  and g41336 (n25742, n_11413, n_18601);
  not g41337 (n_18602, n25740);
  and g41338 (n25743, n_18602, n25742);
  not g41339 (n_18603, n25684);
  and g41340 (n25744, n_11412, n_18603);
  not g41341 (n_18604, n25743);
  and g41342 (n25745, n_18604, n25744);
  and g41343 (n25746, n_11984, n25681);
  and g41344 (n25747, pi0618, n25594);
  not g41345 (n_18605, n25747);
  and g41346 (n25748, n_11413, n_18605);
  not g41347 (n_18606, n25746);
  and g41348 (n25749, n_18606, n25748);
  and g41349 (n25750, n_11984, n25622);
  and g41350 (n25751, pi0618, n_18600);
  not g41351 (n_18607, n25750);
  and g41352 (n25752, pi1154, n_18607);
  not g41353 (n_18608, n25751);
  and g41354 (n25753, n_18608, n25752);
  not g41355 (n_18609, n25749);
  and g41356 (n25754, pi0627, n_18609);
  not g41357 (n_18610, n25753);
  and g41358 (n25755, n_18610, n25754);
  not g41359 (n_18611, n25745);
  not g41360 (n_18612, n25755);
  and g41361 (n25756, n_18611, n_18612);
  not g41362 (n_18613, n25756);
  and g41363 (n25757, pi0781, n_18613);
  and g41364 (n25758, n_11981, n_18600);
  not g41365 (n_18614, n25757);
  not g41366 (n_18615, n25758);
  and g41367 (n25759, n_18614, n_18615);
  not g41368 (n_18616, n25759);
  and g41369 (n25760, n_11821, n_18616);
  not g41370 (n_18617, n25625);
  and g41371 (n25761, pi0619, n_18617);
  not g41372 (n_18618, n25761);
  and g41373 (n25762, n_11405, n_18618);
  not g41374 (n_18619, n25760);
  and g41375 (n25763, n_18619, n25762);
  and g41376 (n25764, n_11821, n25594);
  not g41377 (n_18620, n25681);
  and g41378 (n25765, n_11981, n_18620);
  and g41379 (n25766, n_18603, n_18609);
  not g41380 (n_18621, n25766);
  and g41381 (n25767, pi0781, n_18621);
  not g41382 (n_18622, n25765);
  not g41383 (n_18623, n25767);
  and g41384 (n25768, n_18622, n_18623);
  and g41385 (n25769, pi0619, n25768);
  not g41386 (n_18624, n25764);
  and g41387 (n25770, pi1159, n_18624);
  not g41388 (n_18625, n25769);
  and g41389 (n25771, n_18625, n25770);
  not g41390 (n_18626, n25771);
  and g41391 (n25772, n_11403, n_18626);
  not g41392 (n_18627, n25763);
  and g41393 (n25773, n_18627, n25772);
  and g41394 (n25774, pi0619, n_18616);
  and g41395 (n25775, n_11821, n_18617);
  not g41396 (n_18628, n25775);
  and g41397 (n25776, pi1159, n_18628);
  not g41398 (n_18629, n25774);
  and g41399 (n25777, n_18629, n25776);
  and g41400 (n25778, n_11821, n25768);
  and g41401 (n25779, pi0619, n25594);
  not g41402 (n_18630, n25779);
  and g41403 (n25780, n_11405, n_18630);
  not g41404 (n_18631, n25778);
  and g41405 (n25781, n_18631, n25780);
  not g41406 (n_18632, n25781);
  and g41407 (n25782, pi0648, n_18632);
  not g41408 (n_18633, n25777);
  and g41409 (n25783, n_18633, n25782);
  not g41410 (n_18634, n25773);
  not g41411 (n_18635, n25783);
  and g41412 (n25784, n_18634, n_18635);
  not g41413 (n_18636, n25784);
  and g41414 (n25785, pi0789, n_18636);
  and g41415 (n25786, n_12315, n_18616);
  not g41416 (n_18637, n25785);
  not g41417 (n_18638, n25786);
  and g41418 (n25787, n_18637, n_18638);
  and g41419 (n25788, n_12318, n25787);
  and g41420 (n25789, n_12320, n25787);
  not g41421 (n_18639, n25627);
  and g41422 (n25790, pi0626, n_18639);
  not g41423 (n_18640, n25790);
  and g41424 (n25791, n_11395, n_18640);
  not g41425 (n_18641, n25789);
  and g41426 (n25792, n_18641, n25791);
  not g41427 (n_18642, n25768);
  and g41428 (n25793, n_12315, n_18642);
  and g41429 (n25794, n_18626, n_18632);
  not g41430 (n_18643, n25794);
  and g41431 (n25795, pi0789, n_18643);
  not g41432 (n_18644, n25793);
  not g41433 (n_18645, n25795);
  and g41434 (n25796, n_18644, n_18645);
  not g41435 (n_18646, n25796);
  and g41436 (n25797, n_12320, n_18646);
  and g41437 (n25798, pi0626, n_18487);
  not g41438 (n_18647, n25798);
  and g41439 (n25799, pi0641, n_18647);
  not g41440 (n_18648, n25797);
  and g41441 (n25800, n_18648, n25799);
  not g41442 (n_18649, n25800);
  and g41443 (n25801, n_11397, n_18649);
  not g41444 (n_18650, n25792);
  and g41445 (n25802, n_18650, n25801);
  and g41446 (n25803, pi0626, n25787);
  and g41447 (n25804, n_12320, n_18639);
  not g41448 (n_18651, n25804);
  and g41449 (n25805, pi0641, n_18651);
  not g41450 (n_18652, n25803);
  and g41451 (n25806, n_18652, n25805);
  and g41452 (n25807, pi0626, n_18646);
  and g41453 (n25808, n_12320, n_18487);
  not g41454 (n_18653, n25808);
  and g41455 (n25809, n_11395, n_18653);
  not g41456 (n_18654, n25807);
  and g41457 (n25810, n_18654, n25809);
  not g41458 (n_18655, n25810);
  and g41459 (n25811, pi1158, n_18655);
  not g41460 (n_18656, n25806);
  and g41461 (n25812, n_18656, n25811);
  not g41462 (n_18657, n25802);
  not g41463 (n_18658, n25812);
  and g41464 (n25813, n_18657, n_18658);
  not g41465 (n_18659, n25813);
  and g41466 (n25814, pi0788, n_18659);
  not g41467 (n_18660, n25788);
  not g41468 (n_18661, n25814);
  and g41469 (n25815, n_18660, n_18661);
  and g41470 (n25816, n_11789, n25815);
  and g41471 (n25817, n_12524, n25796);
  and g41472 (n25818, n17969, n25594);
  not g41473 (n_18662, n25817);
  not g41474 (n_18663, n25818);
  and g41475 (n25819, n_18662, n_18663);
  not g41476 (n_18664, n25819);
  and g41477 (n25820, pi0628, n_18664);
  not g41478 (n_18665, n25820);
  and g41479 (n25821, n_11794, n_18665);
  not g41480 (n_18666, n25816);
  and g41481 (n25822, n_18666, n25821);
  and g41482 (n25823, n_12354, n_18522);
  not g41483 (n_18667, n25822);
  and g41484 (n25824, n_18667, n25823);
  and g41485 (n25825, pi0628, n25815);
  and g41486 (n25826, n_11789, n_18664);
  not g41487 (n_18668, n25826);
  and g41488 (n25827, pi1156, n_18668);
  not g41489 (n_18669, n25825);
  and g41490 (n25828, n_18669, n25827);
  and g41491 (n25829, pi0629, n_18523);
  not g41492 (n_18670, n25828);
  and g41493 (n25830, n_18670, n25829);
  not g41494 (n_18671, n25824);
  not g41495 (n_18672, n25830);
  and g41496 (n25831, n_18671, n_18672);
  not g41497 (n_18673, n25831);
  and g41498 (n25832, pi0792, n_18673);
  and g41499 (n25833, n_11787, n25815);
  not g41500 (n_18674, n25832);
  not g41501 (n_18675, n25833);
  and g41502 (n25834, n_18674, n_18675);
  not g41503 (n_18676, n25834);
  and g41504 (n25835, n_11806, n_18676);
  and g41505 (n25836, n_12368, n_18664);
  and g41506 (n25837, n17779, n25594);
  not g41507 (n_18677, n25836);
  not g41508 (n_18678, n25837);
  and g41509 (n25838, n_18677, n_18678);
  not g41510 (n_18679, n25838);
  and g41511 (n25839, pi0647, n_18679);
  not g41512 (n_18680, n25839);
  and g41513 (n25840, n_11810, n_18680);
  not g41514 (n_18681, n25835);
  and g41515 (n25841, n_18681, n25840);
  and g41516 (n25842, n_12375, n_18532);
  not g41517 (n_18682, n25841);
  and g41518 (n25843, n_18682, n25842);
  and g41519 (n25844, pi0647, n_18676);
  and g41520 (n25845, n_11806, n_18679);
  not g41521 (n_18683, n25845);
  and g41522 (n25846, pi1157, n_18683);
  not g41523 (n_18684, n25844);
  and g41524 (n25847, n_18684, n25846);
  and g41525 (n25848, pi0630, n_18533);
  not g41526 (n_18685, n25847);
  and g41527 (n25849, n_18685, n25848);
  not g41528 (n_18686, n25843);
  not g41529 (n_18687, n25849);
  and g41530 (n25850, n_18686, n_18687);
  not g41531 (n_18688, n25850);
  and g41532 (n25851, pi0787, n_18688);
  and g41533 (n25852, n_11803, n_18676);
  not g41534 (n_18689, n25851);
  not g41535 (n_18690, n25852);
  and g41536 (n25853, n_18689, n_18690);
  not g41537 (n_18691, n25853);
  and g41538 (n25854, pi0644, n_18691);
  not g41539 (n_18692, n25655);
  and g41540 (n25855, pi0715, n_18692);
  not g41541 (n_18693, n25854);
  and g41542 (n25856, n_18693, n25855);
  and g41543 (n25857, n17804, n_18487);
  and g41544 (n25858, n_12392, n25838);
  not g41545 (n_18694, n25857);
  not g41546 (n_18695, n25858);
  and g41547 (n25859, n_18694, n_18695);
  and g41548 (n25860, pi0644, n25859);
  and g41549 (n25861, n_11819, n25594);
  not g41550 (n_18696, n25861);
  and g41551 (n25862, n_12395, n_18696);
  not g41552 (n_18697, n25860);
  and g41553 (n25863, n_18697, n25862);
  not g41554 (n_18698, n25863);
  and g41555 (n25864, pi1160, n_18698);
  not g41556 (n_18699, n25856);
  and g41557 (n25865, n_18699, n25864);
  and g41558 (n25866, n_11819, n_18691);
  and g41559 (n25867, pi0644, n25654);
  not g41560 (n_18700, n25867);
  and g41561 (n25868, n_12395, n_18700);
  not g41562 (n_18701, n25866);
  and g41563 (n25869, n_18701, n25868);
  and g41564 (n25870, n_11819, n25859);
  and g41565 (n25871, pi0644, n25594);
  not g41566 (n_18702, n25871);
  and g41567 (n25872, pi0715, n_18702);
  not g41568 (n_18703, n25870);
  and g41569 (n25873, n_18703, n25872);
  not g41570 (n_18704, n25873);
  and g41571 (n25874, n_12405, n_18704);
  not g41572 (n_18705, n25869);
  and g41573 (n25875, n_18705, n25874);
  not g41574 (n_18706, n25865);
  and g41575 (n25876, pi0790, n_18706);
  not g41576 (n_18707, n25875);
  and g41577 (n25877, n_18707, n25876);
  and g41578 (n25878, n_12411, n25853);
  not g41579 (n_18708, n25878);
  and g41580 (n25879, n_4226, n_18708);
  not g41581 (n_18709, n25877);
  and g41582 (n25880, n_18709, n25879);
  and g41583 (n25881, n_7636, po1038);
  not g41584 (n_18710, n25881);
  and g41585 (n25882, n_12415, n_18710);
  not g41586 (n_18711, n25880);
  and g41587 (n25883, n_18711, n25882);
  and g41588 (n25884, n_7636, n_12418);
  and g41589 (n25885, n_15414, n16645);
  not g41590 (n_18712, n25884);
  not g41591 (n_18713, n25885);
  and g41592 (n25886, n_18712, n_18713);
  and g41593 (n25887, n_11749, n25886);
  and g41594 (n25888, n_11753, n25885);
  not g41595 (n_18714, n25886);
  not g41596 (n_18715, n25888);
  and g41597 (n25889, n_18714, n_18715);
  not g41598 (n_18716, n25889);
  and g41599 (n25890, pi1153, n_18716);
  and g41600 (n25891, n_11757, n_18712);
  and g41601 (n25892, n_18715, n25891);
  not g41602 (n_18717, n25890);
  not g41603 (n_18718, n25892);
  and g41604 (n25893, n_18717, n_18718);
  not g41605 (n_18719, n25893);
  and g41606 (n25894, pi0778, n_18719);
  not g41607 (n_18720, n25887);
  not g41608 (n_18721, n25894);
  and g41609 (n25895, n_18720, n_18721);
  and g41610 (n25896, n_12429, n25895);
  and g41611 (n25897, n_12430, n25896);
  and g41612 (n25898, n_12431, n25897);
  and g41613 (n25899, n_12432, n25898);
  and g41614 (n25900, n_12436, n25899);
  and g41615 (n25901, n_11806, n25900);
  and g41616 (n25902, pi0647, n25884);
  not g41617 (n_18722, n25902);
  and g41618 (n25903, n_11810, n_18722);
  not g41619 (n_18723, n25901);
  and g41620 (n25904, n_18723, n25903);
  and g41621 (n25905, pi0630, n25904);
  and g41622 (n25906, n_15412, n17244);
  not g41623 (n_18724, n25906);
  and g41624 (n25907, n_18712, n_18724);
  not g41625 (n_18725, n25907);
  and g41626 (n25908, n_12448, n_18725);
  not g41627 (n_18726, n25908);
  and g41628 (n25909, n_11964, n_18726);
  and g41629 (n25910, n_12451, n_18725);
  not g41630 (n_18727, n25910);
  and g41631 (n25911, pi1155, n_18727);
  and g41632 (n25912, n_12453, n25908);
  not g41633 (n_18728, n25912);
  and g41634 (n25913, n_11768, n_18728);
  not g41635 (n_18729, n25911);
  not g41636 (n_18730, n25913);
  and g41637 (n25914, n_18729, n_18730);
  not g41638 (n_18731, n25914);
  and g41639 (n25915, pi0785, n_18731);
  not g41640 (n_18732, n25909);
  not g41641 (n_18733, n25915);
  and g41642 (n25916, n_18732, n_18733);
  not g41643 (n_18734, n25916);
  and g41644 (n25917, n_11981, n_18734);
  and g41645 (n25918, n_12461, n25916);
  not g41646 (n_18735, n25918);
  and g41647 (n25919, pi1154, n_18735);
  and g41648 (n25920, n_12463, n25916);
  not g41649 (n_18736, n25920);
  and g41650 (n25921, n_11413, n_18736);
  not g41651 (n_18737, n25919);
  not g41652 (n_18738, n25921);
  and g41653 (n25922, n_18737, n_18738);
  not g41654 (n_18739, n25922);
  and g41655 (n25923, pi0781, n_18739);
  not g41656 (n_18740, n25917);
  not g41657 (n_18741, n25923);
  and g41658 (n25924, n_18740, n_18741);
  not g41659 (n_18742, n25924);
  and g41660 (n25925, n_12315, n_18742);
  and g41661 (n25926, n_11821, n25884);
  and g41662 (n25927, pi0619, n25924);
  not g41663 (n_18743, n25926);
  and g41664 (n25928, pi1159, n_18743);
  not g41665 (n_18744, n25927);
  and g41666 (n25929, n_18744, n25928);
  and g41667 (n25930, n_11821, n25924);
  and g41668 (n25931, pi0619, n25884);
  not g41669 (n_18745, n25931);
  and g41670 (n25932, n_11405, n_18745);
  not g41671 (n_18746, n25930);
  and g41672 (n25933, n_18746, n25932);
  not g41673 (n_18747, n25929);
  not g41674 (n_18748, n25933);
  and g41675 (n25934, n_18747, n_18748);
  not g41676 (n_18749, n25934);
  and g41677 (n25935, pi0789, n_18749);
  not g41678 (n_18750, n25925);
  not g41679 (n_18751, n25935);
  and g41680 (n25936, n_18750, n_18751);
  and g41681 (n25937, n_12524, n25936);
  and g41682 (n25938, n17969, n25884);
  not g41683 (n_18752, n25937);
  not g41684 (n_18753, n25938);
  and g41685 (n25939, n_18752, n_18753);
  not g41686 (n_18754, n25939);
  and g41687 (n25940, n_12368, n_18754);
  and g41688 (n25941, n17779, n25884);
  not g41689 (n_18755, n25940);
  not g41690 (n_18756, n25941);
  and g41691 (n25942, n_18755, n_18756);
  and g41692 (n25943, n_14548, n25942);
  not g41693 (n_18757, n25900);
  and g41694 (n25944, pi0647, n_18757);
  and g41695 (n25945, n_11806, n_18712);
  not g41696 (n_18758, n25944);
  not g41697 (n_18759, n25945);
  and g41698 (n25946, n_18758, n_18759);
  not g41699 (n_18760, n25946);
  and g41700 (n25947, n17801, n_18760);
  not g41701 (n_18761, n25905);
  not g41702 (n_18762, n25947);
  and g41703 (n25948, n_18761, n_18762);
  not g41704 (n_18763, n25943);
  and g41705 (n25949, n_18763, n25948);
  not g41706 (n_18764, n25949);
  and g41707 (n25950, pi0787, n_18764);
  and g41708 (n25951, n17871, n25898);
  not g41709 (n_18765, n25936);
  and g41710 (n25952, n_12320, n_18765);
  and g41711 (n25953, pi0626, n_18712);
  not g41712 (n_18766, n25953);
  and g41713 (n25954, n16629, n_18766);
  not g41714 (n_18767, n25952);
  and g41715 (n25955, n_18767, n25954);
  and g41716 (n25956, pi0626, n_18765);
  and g41717 (n25957, n_12320, n_18712);
  not g41718 (n_18768, n25957);
  and g41719 (n25958, n16628, n_18768);
  not g41720 (n_18769, n25956);
  and g41721 (n25959, n_18769, n25958);
  not g41722 (n_18770, n25951);
  not g41723 (n_18771, n25955);
  and g41724 (n25960, n_18770, n_18771);
  not g41725 (n_18772, n25959);
  and g41726 (n25961, n_18772, n25960);
  not g41727 (n_18773, n25961);
  and g41728 (n25962, pi0788, n_18773);
  and g41729 (n25963, pi0618, n25896);
  and g41730 (n25964, pi0609, n25895);
  and g41731 (n25965, n_11866, n_18714);
  and g41732 (n25966, pi0625, n25965);
  not g41733 (n_18774, n25965);
  and g41734 (n25967, n25907, n_18774);
  not g41735 (n_18775, n25966);
  not g41736 (n_18776, n25967);
  and g41737 (n25968, n_18775, n_18776);
  not g41738 (n_18777, n25968);
  and g41739 (n25969, n25891, n_18777);
  and g41740 (n25970, n_11823, n_18717);
  not g41741 (n_18778, n25969);
  and g41742 (n25971, n_18778, n25970);
  and g41743 (n25972, pi1153, n25907);
  and g41744 (n25973, n_18775, n25972);
  and g41745 (n25974, pi0608, n_18718);
  not g41746 (n_18779, n25973);
  and g41747 (n25975, n_18779, n25974);
  not g41748 (n_18780, n25971);
  not g41749 (n_18781, n25975);
  and g41750 (n25976, n_18780, n_18781);
  not g41751 (n_18782, n25976);
  and g41752 (n25977, pi0778, n_18782);
  and g41753 (n25978, n_11749, n_18776);
  not g41754 (n_18783, n25977);
  not g41755 (n_18784, n25978);
  and g41756 (n25979, n_18783, n_18784);
  not g41757 (n_18785, n25979);
  and g41758 (n25980, n_11971, n_18785);
  not g41759 (n_18786, n25964);
  and g41760 (n25981, n_11768, n_18786);
  not g41761 (n_18787, n25980);
  and g41762 (n25982, n_18787, n25981);
  and g41763 (n25983, n_11767, n_18729);
  not g41764 (n_18788, n25982);
  and g41765 (n25984, n_18788, n25983);
  and g41766 (n25985, n_11971, n25895);
  and g41767 (n25986, pi0609, n_18785);
  not g41768 (n_18789, n25985);
  and g41769 (n25987, pi1155, n_18789);
  not g41770 (n_18790, n25986);
  and g41771 (n25988, n_18790, n25987);
  and g41772 (n25989, pi0660, n_18730);
  not g41773 (n_18791, n25988);
  and g41774 (n25990, n_18791, n25989);
  not g41775 (n_18792, n25984);
  not g41776 (n_18793, n25990);
  and g41777 (n25991, n_18792, n_18793);
  not g41778 (n_18794, n25991);
  and g41779 (n25992, pi0785, n_18794);
  and g41780 (n25993, n_11964, n_18785);
  not g41781 (n_18795, n25992);
  not g41782 (n_18796, n25993);
  and g41783 (n25994, n_18795, n_18796);
  not g41784 (n_18797, n25994);
  and g41785 (n25995, n_11984, n_18797);
  not g41786 (n_18798, n25963);
  and g41787 (n25996, n_11413, n_18798);
  not g41788 (n_18799, n25995);
  and g41789 (n25997, n_18799, n25996);
  and g41790 (n25998, n_11412, n_18737);
  not g41791 (n_18800, n25997);
  and g41792 (n25999, n_18800, n25998);
  and g41793 (n26000, n_11984, n25896);
  and g41794 (n26001, pi0618, n_18797);
  not g41795 (n_18801, n26000);
  and g41796 (n26002, pi1154, n_18801);
  not g41797 (n_18802, n26001);
  and g41798 (n26003, n_18802, n26002);
  and g41799 (n26004, pi0627, n_18738);
  not g41800 (n_18803, n26003);
  and g41801 (n26005, n_18803, n26004);
  not g41802 (n_18804, n25999);
  not g41803 (n_18805, n26005);
  and g41804 (n26006, n_18804, n_18805);
  not g41805 (n_18806, n26006);
  and g41806 (n26007, pi0781, n_18806);
  and g41807 (n26008, n_11981, n_18797);
  not g41808 (n_18807, n26007);
  not g41809 (n_18808, n26008);
  and g41810 (n26009, n_18807, n_18808);
  and g41811 (n26010, n_12315, n26009);
  not g41812 (n_18809, n26009);
  and g41813 (n26011, n_11821, n_18809);
  and g41814 (n26012, pi0619, n25897);
  not g41815 (n_18810, n26012);
  and g41816 (n26013, n_11405, n_18810);
  not g41817 (n_18811, n26011);
  and g41818 (n26014, n_18811, n26013);
  and g41819 (n26015, n_11403, n_18747);
  not g41820 (n_18812, n26014);
  and g41821 (n26016, n_18812, n26015);
  and g41822 (n26017, pi0619, n_18809);
  and g41823 (n26018, n_11821, n25897);
  not g41824 (n_18813, n26018);
  and g41825 (n26019, pi1159, n_18813);
  not g41826 (n_18814, n26017);
  and g41827 (n26020, n_18814, n26019);
  and g41828 (n26021, pi0648, n_18748);
  not g41829 (n_18815, n26020);
  and g41830 (n26022, n_18815, n26021);
  not g41831 (n_18816, n26016);
  and g41832 (n26023, pi0789, n_18816);
  not g41833 (n_18817, n26022);
  and g41834 (n26024, n_18817, n26023);
  not g41835 (n_18818, n26010);
  and g41836 (n26025, n17970, n_18818);
  not g41837 (n_18819, n26024);
  and g41838 (n26026, n_18819, n26025);
  not g41839 (n_18820, n25962);
  not g41840 (n_18821, n26026);
  and g41841 (n26027, n_18820, n_18821);
  not g41842 (n_18822, n26027);
  and g41843 (n26028, n_14638, n_18822);
  and g41844 (n26029, n17854, n_18754);
  and g41845 (n26030, n20851, n25899);
  not g41846 (n_18823, n26029);
  not g41847 (n_18824, n26030);
  and g41848 (n26031, n_18823, n_18824);
  not g41849 (n_18825, n26031);
  and g41850 (n26032, n_12354, n_18825);
  and g41851 (n26033, n20855, n25899);
  and g41852 (n26034, n17853, n_18754);
  not g41853 (n_18826, n26033);
  not g41854 (n_18827, n26034);
  and g41855 (n26035, n_18826, n_18827);
  not g41856 (n_18828, n26035);
  and g41857 (n26036, pi0629, n_18828);
  not g41858 (n_18829, n26032);
  not g41859 (n_18830, n26036);
  and g41860 (n26037, n_18829, n_18830);
  not g41861 (n_18831, n26037);
  and g41862 (n26038, pi0792, n_18831);
  not g41863 (n_18832, n26038);
  and g41864 (n26039, n_14387, n_18832);
  not g41865 (n_18833, n26028);
  and g41866 (n26040, n_18833, n26039);
  not g41867 (n_18834, n25950);
  not g41868 (n_18835, n26040);
  and g41869 (n26041, n_18834, n_18835);
  and g41870 (n26042, n_12411, n26041);
  and g41871 (n26043, n_11803, n_18757);
  and g41872 (n26044, pi1157, n_18760);
  not g41873 (n_18836, n25904);
  not g41874 (n_18837, n26044);
  and g41875 (n26045, n_18836, n_18837);
  not g41876 (n_18838, n26045);
  and g41877 (n26046, pi0787, n_18838);
  not g41878 (n_18839, n26043);
  not g41879 (n_18840, n26046);
  and g41880 (n26047, n_18839, n_18840);
  and g41881 (n26048, n_11819, n26047);
  and g41882 (n26049, pi0644, n26041);
  not g41883 (n_18841, n26048);
  and g41884 (n26050, pi0715, n_18841);
  not g41885 (n_18842, n26049);
  and g41886 (n26051, n_18842, n26050);
  not g41887 (n_18843, n25942);
  and g41888 (n26052, n_12392, n_18843);
  and g41889 (n26053, n17804, n25884);
  not g41890 (n_18844, n26052);
  not g41891 (n_18845, n26053);
  and g41892 (n26054, n_18844, n_18845);
  not g41893 (n_18846, n26054);
  and g41894 (n26055, pi0644, n_18846);
  and g41895 (n26056, n_11819, n25884);
  not g41896 (n_18847, n26056);
  and g41897 (n26057, n_12395, n_18847);
  not g41898 (n_18848, n26055);
  and g41899 (n26058, n_18848, n26057);
  not g41900 (n_18849, n26058);
  and g41901 (n26059, pi1160, n_18849);
  not g41902 (n_18850, n26051);
  and g41903 (n26060, n_18850, n26059);
  and g41904 (n26061, n_11819, n_18846);
  and g41905 (n26062, pi0644, n25884);
  not g41906 (n_18851, n26062);
  and g41907 (n26063, pi0715, n_18851);
  not g41908 (n_18852, n26061);
  and g41909 (n26064, n_18852, n26063);
  and g41910 (n26065, pi0644, n26047);
  and g41911 (n26066, n_11819, n26041);
  not g41912 (n_18853, n26065);
  and g41913 (n26067, n_12395, n_18853);
  not g41914 (n_18854, n26066);
  and g41915 (n26068, n_18854, n26067);
  not g41916 (n_18855, n26064);
  and g41917 (n26069, n_12405, n_18855);
  not g41918 (n_18856, n26068);
  and g41919 (n26070, n_18856, n26069);
  not g41920 (n_18857, n26060);
  not g41921 (n_18858, n26070);
  and g41922 (n26071, n_18857, n_18858);
  not g41923 (n_18859, n26071);
  and g41924 (n26072, pi0790, n_18859);
  not g41925 (n_18860, n26042);
  and g41926 (n26073, pi0832, n_18860);
  not g41927 (n_18861, n26072);
  and g41928 (n26074, n_18861, n26073);
  not g41929 (n_18862, n25883);
  not g41930 (n_18863, n26074);
  and g41931 (po0336, n_18862, n_18863);
  and g41932 (n26076, n_6015, n_12418);
  and g41933 (n26077, n_15518, n16645);
  not g41934 (n_18864, n26076);
  not g41935 (n_18865, n26077);
  and g41936 (n26078, n_18864, n_18865);
  not g41937 (n_18866, n26078);
  and g41938 (n26079, n_11749, n_18866);
  and g41939 (n26080, n_11753, n26077);
  not g41940 (n_18867, n26080);
  and g41941 (n26081, n_18866, n_18867);
  not g41942 (n_18868, n26081);
  and g41943 (n26082, pi1153, n_18868);
  and g41944 (n26083, n_11757, n_18864);
  and g41945 (n26084, n_18867, n26083);
  not g41946 (n_18869, n26084);
  and g41947 (n26085, pi0778, n_18869);
  not g41948 (n_18870, n26082);
  and g41949 (n26086, n_18870, n26085);
  not g41950 (n_18871, n26079);
  not g41951 (n_18872, n26086);
  and g41952 (n26087, n_18871, n_18872);
  not g41953 (n_18873, n26087);
  and g41954 (n26088, n_12429, n_18873);
  and g41955 (n26089, n_12430, n26088);
  and g41956 (n26090, n_12431, n26089);
  and g41957 (n26091, n_12432, n26090);
  and g41958 (n26092, n_12436, n26091);
  and g41959 (n26093, n_11806, n26092);
  and g41960 (n26094, pi0647, n26076);
  not g41961 (n_18874, n26094);
  and g41962 (n26095, n_11810, n_18874);
  not g41963 (n_18875, n26093);
  and g41964 (n26096, n_18875, n26095);
  and g41965 (n26097, pi0630, n26096);
  and g41966 (n26098, n_15488, n17244);
  not g41967 (n_18876, n26098);
  and g41968 (n26099, n_18864, n_18876);
  not g41969 (n_18877, n26099);
  and g41970 (n26100, n_12448, n_18877);
  not g41971 (n_18878, n26100);
  and g41972 (n26101, n_11964, n_18878);
  and g41973 (n26102, n17296, n26098);
  not g41974 (n_18879, n26102);
  and g41975 (n26103, n26100, n_18879);
  not g41976 (n_18880, n26103);
  and g41977 (n26104, pi1155, n_18880);
  and g41978 (n26105, n_11768, n_18864);
  and g41979 (n26106, n_18879, n26105);
  not g41980 (n_18881, n26104);
  not g41981 (n_18882, n26106);
  and g41982 (n26107, n_18881, n_18882);
  not g41983 (n_18883, n26107);
  and g41984 (n26108, pi0785, n_18883);
  not g41985 (n_18884, n26101);
  not g41986 (n_18885, n26108);
  and g41987 (n26109, n_18884, n_18885);
  not g41988 (n_18886, n26109);
  and g41989 (n26110, n_11981, n_18886);
  and g41990 (n26111, n_12461, n26109);
  not g41991 (n_18887, n26111);
  and g41992 (n26112, pi1154, n_18887);
  and g41993 (n26113, n_12463, n26109);
  not g41994 (n_18888, n26113);
  and g41995 (n26114, n_11413, n_18888);
  not g41996 (n_18889, n26112);
  not g41997 (n_18890, n26114);
  and g41998 (n26115, n_18889, n_18890);
  not g41999 (n_18891, n26115);
  and g42000 (n26116, pi0781, n_18891);
  not g42001 (n_18892, n26110);
  not g42002 (n_18893, n26116);
  and g42003 (n26117, n_18892, n_18893);
  not g42004 (n_18894, n26117);
  and g42005 (n26118, n_12315, n_18894);
  and g42006 (n26119, n_16503, n26117);
  not g42007 (n_18895, n26119);
  and g42008 (n26120, pi1159, n_18895);
  and g42009 (n26121, n_16505, n26117);
  not g42010 (n_18896, n26121);
  and g42011 (n26122, n_11405, n_18896);
  not g42012 (n_18897, n26120);
  not g42013 (n_18898, n26122);
  and g42014 (n26123, n_18897, n_18898);
  not g42015 (n_18899, n26123);
  and g42016 (n26124, pi0789, n_18899);
  not g42017 (n_18900, n26118);
  not g42018 (n_18901, n26124);
  and g42019 (n26125, n_18900, n_18901);
  and g42020 (n26126, n_12524, n26125);
  and g42021 (n26127, n17969, n26076);
  not g42022 (n_18902, n26126);
  not g42023 (n_18903, n26127);
  and g42024 (n26128, n_18902, n_18903);
  not g42025 (n_18904, n26128);
  and g42026 (n26129, n_12368, n_18904);
  and g42027 (n26130, n17779, n26076);
  not g42028 (n_18905, n26129);
  not g42029 (n_18906, n26130);
  and g42030 (n26131, n_18905, n_18906);
  and g42031 (n26132, n_14548, n26131);
  not g42032 (n_18907, n26092);
  and g42033 (n26133, pi0647, n_18907);
  and g42034 (n26134, n_11806, n_18864);
  not g42035 (n_18908, n26133);
  not g42036 (n_18909, n26134);
  and g42037 (n26135, n_18908, n_18909);
  not g42038 (n_18910, n26135);
  and g42039 (n26136, n17801, n_18910);
  not g42040 (n_18911, n26097);
  not g42041 (n_18912, n26136);
  and g42042 (n26137, n_18911, n_18912);
  not g42043 (n_18913, n26132);
  and g42044 (n26138, n_18913, n26137);
  not g42045 (n_18914, n26138);
  and g42046 (n26139, pi0787, n_18914);
  and g42047 (n26140, n17871, n26090);
  not g42048 (n_18915, n26125);
  and g42049 (n26141, n_12320, n_18915);
  and g42050 (n26142, pi0626, n_18864);
  not g42051 (n_18916, n26142);
  and g42052 (n26143, n16629, n_18916);
  not g42053 (n_18917, n26141);
  and g42054 (n26144, n_18917, n26143);
  and g42055 (n26145, pi0626, n_18915);
  and g42056 (n26146, n_12320, n_18864);
  not g42057 (n_18918, n26146);
  and g42058 (n26147, n16628, n_18918);
  not g42059 (n_18919, n26145);
  and g42060 (n26148, n_18919, n26147);
  not g42061 (n_18920, n26140);
  not g42062 (n_18921, n26144);
  and g42063 (n26149, n_18920, n_18921);
  not g42064 (n_18922, n26148);
  and g42065 (n26150, n_18922, n26149);
  not g42066 (n_18923, n26150);
  and g42067 (n26151, pi0788, n_18923);
  and g42068 (n26152, pi0618, n26088);
  and g42069 (n26153, n_11866, n_18866);
  and g42070 (n26154, pi0625, n26153);
  not g42071 (n_18924, n26153);
  and g42072 (n26155, n26099, n_18924);
  not g42073 (n_18925, n26154);
  not g42074 (n_18926, n26155);
  and g42075 (n26156, n_18925, n_18926);
  not g42076 (n_18927, n26156);
  and g42077 (n26157, n26083, n_18927);
  and g42078 (n26158, n_11823, n_18870);
  not g42079 (n_18928, n26157);
  and g42080 (n26159, n_18928, n26158);
  and g42081 (n26160, pi1153, n26099);
  and g42082 (n26161, n_18925, n26160);
  and g42083 (n26162, pi0608, n_18869);
  not g42084 (n_18929, n26161);
  and g42085 (n26163, n_18929, n26162);
  not g42086 (n_18930, n26159);
  not g42087 (n_18931, n26163);
  and g42088 (n26164, n_18930, n_18931);
  not g42089 (n_18932, n26164);
  and g42090 (n26165, pi0778, n_18932);
  and g42091 (n26166, n_11749, n_18926);
  not g42092 (n_18933, n26165);
  not g42093 (n_18934, n26166);
  and g42094 (n26167, n_18933, n_18934);
  not g42095 (n_18935, n26167);
  and g42096 (n26168, n_11971, n_18935);
  and g42097 (n26169, pi0609, n_18873);
  not g42098 (n_18936, n26169);
  and g42099 (n26170, n_11768, n_18936);
  not g42100 (n_18937, n26168);
  and g42101 (n26171, n_18937, n26170);
  and g42102 (n26172, n_11767, n_18881);
  not g42103 (n_18938, n26171);
  and g42104 (n26173, n_18938, n26172);
  and g42105 (n26174, pi0609, n_18935);
  and g42106 (n26175, n_11971, n_18873);
  not g42107 (n_18939, n26175);
  and g42108 (n26176, pi1155, n_18939);
  not g42109 (n_18940, n26174);
  and g42110 (n26177, n_18940, n26176);
  and g42111 (n26178, pi0660, n_18882);
  not g42112 (n_18941, n26177);
  and g42113 (n26179, n_18941, n26178);
  not g42114 (n_18942, n26173);
  not g42115 (n_18943, n26179);
  and g42116 (n26180, n_18942, n_18943);
  not g42117 (n_18944, n26180);
  and g42118 (n26181, pi0785, n_18944);
  and g42119 (n26182, n_11964, n_18935);
  not g42120 (n_18945, n26181);
  not g42121 (n_18946, n26182);
  and g42122 (n26183, n_18945, n_18946);
  not g42123 (n_18947, n26183);
  and g42124 (n26184, n_11984, n_18947);
  not g42125 (n_18948, n26152);
  and g42126 (n26185, n_11413, n_18948);
  not g42127 (n_18949, n26184);
  and g42128 (n26186, n_18949, n26185);
  and g42129 (n26187, n_11412, n_18889);
  not g42130 (n_18950, n26186);
  and g42131 (n26188, n_18950, n26187);
  and g42132 (n26189, n_11984, n26088);
  and g42133 (n26190, pi0618, n_18947);
  not g42134 (n_18951, n26189);
  and g42135 (n26191, pi1154, n_18951);
  not g42136 (n_18952, n26190);
  and g42137 (n26192, n_18952, n26191);
  and g42138 (n26193, pi0627, n_18890);
  not g42139 (n_18953, n26192);
  and g42140 (n26194, n_18953, n26193);
  not g42141 (n_18954, n26188);
  not g42142 (n_18955, n26194);
  and g42143 (n26195, n_18954, n_18955);
  not g42144 (n_18956, n26195);
  and g42145 (n26196, pi0781, n_18956);
  and g42146 (n26197, n_11981, n_18947);
  not g42147 (n_18957, n26196);
  not g42148 (n_18958, n26197);
  and g42149 (n26198, n_18957, n_18958);
  and g42150 (n26199, n_12315, n26198);
  not g42151 (n_18959, n26198);
  and g42152 (n26200, n_11821, n_18959);
  and g42153 (n26201, pi0619, n26089);
  not g42154 (n_18960, n26201);
  and g42155 (n26202, n_11405, n_18960);
  not g42156 (n_18961, n26200);
  and g42157 (n26203, n_18961, n26202);
  and g42158 (n26204, n_11403, n_18897);
  not g42159 (n_18962, n26203);
  and g42160 (n26205, n_18962, n26204);
  and g42161 (n26206, pi0619, n_18959);
  and g42162 (n26207, n_11821, n26089);
  not g42163 (n_18963, n26207);
  and g42164 (n26208, pi1159, n_18963);
  not g42165 (n_18964, n26206);
  and g42166 (n26209, n_18964, n26208);
  and g42167 (n26210, pi0648, n_18898);
  not g42168 (n_18965, n26209);
  and g42169 (n26211, n_18965, n26210);
  not g42170 (n_18966, n26205);
  and g42171 (n26212, pi0789, n_18966);
  not g42172 (n_18967, n26211);
  and g42173 (n26213, n_18967, n26212);
  not g42174 (n_18968, n26199);
  and g42175 (n26214, n17970, n_18968);
  not g42176 (n_18969, n26213);
  and g42177 (n26215, n_18969, n26214);
  not g42178 (n_18970, n26151);
  not g42179 (n_18971, n26215);
  and g42180 (n26216, n_18970, n_18971);
  not g42181 (n_18972, n26216);
  and g42182 (n26217, n_14638, n_18972);
  and g42183 (n26218, n17854, n_18904);
  and g42184 (n26219, n20851, n26091);
  not g42185 (n_18973, n26218);
  not g42186 (n_18974, n26219);
  and g42187 (n26220, n_18973, n_18974);
  not g42188 (n_18975, n26220);
  and g42189 (n26221, n_12354, n_18975);
  and g42190 (n26222, n20855, n26091);
  and g42191 (n26223, n17853, n_18904);
  not g42192 (n_18976, n26222);
  not g42193 (n_18977, n26223);
  and g42194 (n26224, n_18976, n_18977);
  not g42195 (n_18978, n26224);
  and g42196 (n26225, pi0629, n_18978);
  not g42197 (n_18979, n26221);
  not g42198 (n_18980, n26225);
  and g42199 (n26226, n_18979, n_18980);
  not g42200 (n_18981, n26226);
  and g42201 (n26227, pi0792, n_18981);
  not g42202 (n_18982, n26227);
  and g42203 (n26228, n_14387, n_18982);
  not g42204 (n_18983, n26217);
  and g42205 (n26229, n_18983, n26228);
  not g42206 (n_18984, n26139);
  not g42207 (n_18985, n26229);
  and g42208 (n26230, n_18984, n_18985);
  and g42209 (n26231, n_12411, n26230);
  and g42210 (n26232, n_11803, n_18907);
  and g42211 (n26233, pi1157, n_18910);
  not g42212 (n_18986, n26096);
  not g42213 (n_18987, n26233);
  and g42214 (n26234, n_18986, n_18987);
  not g42215 (n_18988, n26234);
  and g42216 (n26235, pi0787, n_18988);
  not g42217 (n_18989, n26232);
  not g42218 (n_18990, n26235);
  and g42219 (n26236, n_18989, n_18990);
  and g42220 (n26237, n_11819, n26236);
  and g42221 (n26238, pi0644, n26230);
  not g42222 (n_18991, n26237);
  and g42223 (n26239, pi0715, n_18991);
  not g42224 (n_18992, n26238);
  and g42225 (n26240, n_18992, n26239);
  not g42226 (n_18993, n26131);
  and g42227 (n26241, n_12392, n_18993);
  and g42228 (n26242, n17804, n26076);
  not g42229 (n_18994, n26241);
  not g42230 (n_18995, n26242);
  and g42231 (n26243, n_18994, n_18995);
  not g42232 (n_18996, n26243);
  and g42233 (n26244, pi0644, n_18996);
  and g42234 (n26245, n_11819, n26076);
  not g42235 (n_18997, n26245);
  and g42236 (n26246, n_12395, n_18997);
  not g42237 (n_18998, n26244);
  and g42238 (n26247, n_18998, n26246);
  not g42239 (n_18999, n26247);
  and g42240 (n26248, pi1160, n_18999);
  not g42241 (n_19000, n26240);
  and g42242 (n26249, n_19000, n26248);
  and g42243 (n26250, n_11819, n_18996);
  and g42244 (n26251, pi0644, n26076);
  not g42245 (n_19001, n26251);
  and g42246 (n26252, pi0715, n_19001);
  not g42247 (n_19002, n26250);
  and g42248 (n26253, n_19002, n26252);
  and g42249 (n26254, pi0644, n26236);
  and g42250 (n26255, n_11819, n26230);
  not g42251 (n_19003, n26254);
  and g42252 (n26256, n_12395, n_19003);
  not g42253 (n_19004, n26255);
  and g42254 (n26257, n_19004, n26256);
  not g42255 (n_19005, n26253);
  and g42256 (n26258, n_12405, n_19005);
  not g42257 (n_19006, n26257);
  and g42258 (n26259, n_19006, n26258);
  not g42259 (n_19007, n26249);
  not g42260 (n_19008, n26259);
  and g42261 (n26260, n_19007, n_19008);
  not g42262 (n_19009, n26260);
  and g42263 (n26261, pi0790, n_19009);
  not g42264 (n_19010, n26231);
  and g42265 (n26262, pi0832, n_19010);
  not g42266 (n_19011, n26261);
  and g42267 (n26263, n_19011, n26262);
  and g42268 (n26264, n_6015, po1038);
  and g42269 (n26265, n_6015, n_11751);
  not g42270 (n_19012, n26265);
  and g42271 (n26266, n16635, n_19012);
  and g42272 (n26267, n_15518, n2571);
  not g42273 (n_19013, n26267);
  and g42274 (n26268, n26265, n_19013);
  and g42275 (n26269, n_6015, n_11418);
  not g42276 (n_19014, n26269);
  and g42277 (n26270, n16647, n_19014);
  and g42278 (n26271, pi0180, n_12608);
  not g42279 (n_19015, n26271);
  and g42280 (n26272, n_161, n_19015);
  not g42281 (n_19016, n26272);
  and g42282 (n26273, n2571, n_19016);
  and g42283 (n26274, n_6015, n18072);
  not g42284 (n_19017, n26273);
  not g42285 (n_19018, n26274);
  and g42286 (n26275, n_19017, n_19018);
  not g42287 (n_19019, n26270);
  and g42288 (n26276, n_15518, n_19019);
  not g42289 (n_19020, n26275);
  and g42290 (n26277, n_19020, n26276);
  not g42291 (n_19021, n26268);
  not g42292 (n_19022, n26277);
  and g42293 (n26278, n_19021, n_19022);
  and g42294 (n26279, n_11749, n26278);
  and g42295 (n26280, n_11753, n26265);
  not g42296 (n_19023, n26278);
  and g42297 (n26281, pi0625, n_19023);
  not g42298 (n_19024, n26280);
  and g42299 (n26282, pi1153, n_19024);
  not g42300 (n_19025, n26281);
  and g42301 (n26283, n_19025, n26282);
  and g42302 (n26284, pi0625, n26265);
  and g42303 (n26285, n_11753, n_19023);
  not g42304 (n_19026, n26284);
  and g42305 (n26286, n_11757, n_19026);
  not g42306 (n_19027, n26285);
  and g42307 (n26287, n_19027, n26286);
  not g42308 (n_19028, n26283);
  not g42309 (n_19029, n26287);
  and g42310 (n26288, n_19028, n_19029);
  not g42311 (n_19030, n26288);
  and g42312 (n26289, pi0778, n_19030);
  not g42313 (n_19031, n26279);
  not g42314 (n_19032, n26289);
  and g42315 (n26290, n_19031, n_19032);
  not g42316 (n_19033, n26290);
  and g42317 (n26291, n_11773, n_19033);
  and g42318 (n26292, n17075, n_19012);
  not g42319 (n_19034, n26291);
  not g42320 (n_19035, n26292);
  and g42321 (n26293, n_19034, n_19035);
  and g42322 (n26294, n_11777, n26293);
  and g42323 (n26295, n16639, n26265);
  not g42324 (n_19036, n26294);
  not g42325 (n_19037, n26295);
  and g42326 (n26296, n_19036, n_19037);
  and g42327 (n26297, n_11780, n26296);
  not g42328 (n_19038, n26266);
  not g42329 (n_19039, n26297);
  and g42330 (n26298, n_19038, n_19039);
  and g42331 (n26299, n_11783, n26298);
  and g42332 (n26300, n16631, n26265);
  not g42333 (n_19040, n26299);
  not g42334 (n_19041, n26300);
  and g42335 (n26301, n_19040, n_19041);
  and g42336 (n26302, n_11787, n26301);
  not g42337 (n_19042, n26301);
  and g42338 (n26303, pi0628, n_19042);
  and g42339 (n26304, n_11789, n26265);
  not g42340 (n_19043, n26304);
  and g42341 (n26305, pi1156, n_19043);
  not g42342 (n_19044, n26303);
  and g42343 (n26306, n_19044, n26305);
  and g42344 (n26307, pi0628, n26265);
  and g42345 (n26308, n_11789, n_19042);
  not g42346 (n_19045, n26307);
  and g42347 (n26309, n_11794, n_19045);
  not g42348 (n_19046, n26308);
  and g42349 (n26310, n_19046, n26309);
  not g42350 (n_19047, n26306);
  not g42351 (n_19048, n26310);
  and g42352 (n26311, n_19047, n_19048);
  not g42353 (n_19049, n26311);
  and g42354 (n26312, pi0792, n_19049);
  not g42355 (n_19050, n26302);
  not g42356 (n_19051, n26312);
  and g42357 (n26313, n_19050, n_19051);
  not g42358 (n_19052, n26313);
  and g42359 (n26314, n_11806, n_19052);
  and g42360 (n26315, pi0647, n_19012);
  not g42361 (n_19053, n26314);
  not g42362 (n_19054, n26315);
  and g42363 (n26316, n_19053, n_19054);
  and g42364 (n26317, n_11810, n26316);
  and g42365 (n26318, pi0647, n_19052);
  and g42366 (n26319, n_11806, n_19012);
  not g42367 (n_19055, n26318);
  not g42368 (n_19056, n26319);
  and g42369 (n26320, n_19055, n_19056);
  and g42370 (n26321, pi1157, n26320);
  not g42371 (n_19057, n26317);
  not g42372 (n_19058, n26321);
  and g42373 (n26322, n_19057, n_19058);
  not g42374 (n_19059, n26322);
  and g42375 (n26323, pi0787, n_19059);
  and g42376 (n26324, n_11803, n26313);
  not g42377 (n_19060, n26323);
  not g42378 (n_19061, n26324);
  and g42379 (n26325, n_19060, n_19061);
  not g42380 (n_19062, n26325);
  and g42381 (n26326, n_11819, n_19062);
  not g42382 (n_19063, n26326);
  and g42383 (n26327, pi0715, n_19063);
  and g42384 (n26328, pi0180, n_11417);
  and g42385 (n26329, pi0180, pi0753);
  and g42386 (n26330, pi0753, n17046);
  and g42387 (n26331, pi0180, n17273);
  not g42388 (n_19064, n26330);
  not g42389 (n_19065, n26331);
  and g42390 (n26332, n_19064, n_19065);
  not g42391 (n_19066, n26332);
  and g42392 (n26333, pi0039, n_19066);
  and g42393 (n26334, pi0180, n_11923);
  not g42394 (n_19067, n26334);
  and g42395 (n26335, n_15494, n_19067);
  not g42396 (n_19068, n26335);
  and g42397 (n26336, n_162, n_19068);
  and g42398 (n26337, n_6015, n_15488);
  and g42399 (n26338, n17221, n26337);
  not g42407 (n_19073, n26341);
  and g42408 (n26342, n_161, n_19073);
  and g42409 (n26343, n_15488, n17280);
  and g42410 (n26344, pi0038, n_19014);
  not g42411 (n_19074, n26343);
  and g42412 (n26345, n_19074, n26344);
  not g42413 (n_19075, n26342);
  not g42414 (n_19076, n26345);
  and g42415 (n26346, n_19075, n_19076);
  not g42416 (n_19077, n26346);
  and g42417 (n26347, n2571, n_19077);
  not g42418 (n_19078, n26328);
  not g42419 (n_19079, n26347);
  and g42420 (n26348, n_19078, n_19079);
  not g42421 (n_19080, n26348);
  and g42422 (n26349, n_11960, n_19080);
  and g42423 (n26350, n17117, n_19012);
  not g42424 (n_19081, n26349);
  not g42425 (n_19082, n26350);
  and g42426 (n26351, n_19081, n_19082);
  not g42427 (n_19083, n26351);
  and g42428 (n26352, n_11964, n_19083);
  and g42429 (n26353, n_11967, n_19012);
  and g42430 (n26354, pi0609, n26349);
  not g42431 (n_19084, n26353);
  not g42432 (n_19085, n26354);
  and g42433 (n26355, n_19084, n_19085);
  not g42434 (n_19086, n26355);
  and g42435 (n26356, pi1155, n_19086);
  and g42436 (n26357, n_11972, n_19012);
  and g42437 (n26358, n_11971, n26349);
  not g42438 (n_19087, n26357);
  not g42439 (n_19088, n26358);
  and g42440 (n26359, n_19087, n_19088);
  not g42441 (n_19089, n26359);
  and g42442 (n26360, n_11768, n_19089);
  not g42443 (n_19090, n26356);
  not g42444 (n_19091, n26360);
  and g42445 (n26361, n_19090, n_19091);
  not g42446 (n_19092, n26361);
  and g42447 (n26362, pi0785, n_19092);
  not g42448 (n_19093, n26352);
  not g42449 (n_19094, n26362);
  and g42450 (n26363, n_19093, n_19094);
  not g42451 (n_19095, n26363);
  and g42452 (n26364, n_11981, n_19095);
  and g42453 (n26365, n_11984, n26265);
  and g42454 (n26366, pi0618, n26363);
  not g42455 (n_19096, n26365);
  and g42456 (n26367, pi1154, n_19096);
  not g42457 (n_19097, n26366);
  and g42458 (n26368, n_19097, n26367);
  and g42459 (n26369, n_11984, n26363);
  and g42460 (n26370, pi0618, n26265);
  not g42461 (n_19098, n26370);
  and g42462 (n26371, n_11413, n_19098);
  not g42463 (n_19099, n26369);
  and g42464 (n26372, n_19099, n26371);
  not g42465 (n_19100, n26368);
  not g42466 (n_19101, n26372);
  and g42467 (n26373, n_19100, n_19101);
  not g42468 (n_19102, n26373);
  and g42469 (n26374, pi0781, n_19102);
  not g42470 (n_19103, n26364);
  not g42471 (n_19104, n26374);
  and g42472 (n26375, n_19103, n_19104);
  not g42473 (n_19105, n26375);
  and g42474 (n26376, n_12315, n_19105);
  and g42475 (n26377, n_11821, n26265);
  and g42476 (n26378, pi0619, n26375);
  not g42477 (n_19106, n26377);
  and g42478 (n26379, pi1159, n_19106);
  not g42479 (n_19107, n26378);
  and g42480 (n26380, n_19107, n26379);
  and g42481 (n26381, n_11821, n26375);
  and g42482 (n26382, pi0619, n26265);
  not g42483 (n_19108, n26382);
  and g42484 (n26383, n_11405, n_19108);
  not g42485 (n_19109, n26381);
  and g42486 (n26384, n_19109, n26383);
  not g42487 (n_19110, n26380);
  not g42488 (n_19111, n26384);
  and g42489 (n26385, n_19110, n_19111);
  not g42490 (n_19112, n26385);
  and g42491 (n26386, pi0789, n_19112);
  not g42492 (n_19113, n26376);
  not g42493 (n_19114, n26386);
  and g42494 (n26387, n_19113, n_19114);
  and g42495 (n26388, n_12524, n26387);
  and g42496 (n26389, n17969, n26265);
  not g42497 (n_19115, n26388);
  not g42498 (n_19116, n26389);
  and g42499 (n26390, n_19115, n_19116);
  not g42500 (n_19117, n26390);
  and g42501 (n26391, n_12368, n_19117);
  and g42502 (n26392, n17779, n26265);
  not g42503 (n_19118, n26391);
  not g42504 (n_19119, n26392);
  and g42505 (n26393, n_19118, n_19119);
  not g42506 (n_19120, n26393);
  and g42507 (n26394, n_12392, n_19120);
  and g42508 (n26395, n17804, n26265);
  not g42509 (n_19121, n26394);
  not g42510 (n_19122, n26395);
  and g42511 (n26396, n_19121, n_19122);
  not g42512 (n_19123, n26396);
  and g42513 (n26397, pi0644, n_19123);
  and g42514 (n26398, n_11819, n26265);
  not g42515 (n_19124, n26398);
  and g42516 (n26399, n_12395, n_19124);
  not g42517 (n_19125, n26397);
  and g42518 (n26400, n_19125, n26399);
  not g42519 (n_19126, n26400);
  and g42520 (n26401, pi1160, n_19126);
  not g42521 (n_19127, n26327);
  and g42522 (n26402, n_19127, n26401);
  and g42523 (n26403, pi0644, n_19062);
  not g42524 (n_19128, n26403);
  and g42525 (n26404, n_12395, n_19128);
  and g42526 (n26405, n_11819, n_19123);
  and g42527 (n26406, pi0644, n26265);
  not g42528 (n_19129, n26406);
  and g42529 (n26407, pi0715, n_19129);
  not g42530 (n_19130, n26405);
  and g42531 (n26408, n_19130, n26407);
  not g42532 (n_19131, n26408);
  and g42533 (n26409, n_12405, n_19131);
  not g42534 (n_19132, n26404);
  and g42535 (n26410, n_19132, n26409);
  not g42536 (n_19133, n26402);
  not g42537 (n_19134, n26410);
  and g42538 (n26411, n_19133, n_19134);
  not g42539 (n_19135, n26411);
  and g42540 (n26412, pi0790, n_19135);
  and g42541 (n26413, n_12354, n26306);
  and g42542 (n26414, n_14557, n26390);
  and g42543 (n26415, pi0629, n26310);
  not g42544 (n_19136, n26413);
  not g42545 (n_19137, n26415);
  and g42546 (n26416, n_19136, n_19137);
  not g42547 (n_19138, n26414);
  and g42548 (n26417, n_19138, n26416);
  not g42549 (n_19139, n26417);
  and g42550 (n26418, pi0792, n_19139);
  and g42551 (n26419, pi0609, n26290);
  and g42552 (n26420, pi0180, n_12240);
  and g42553 (n26421, n_6015, n_12230);
  not g42554 (n_19140, n26420);
  and g42555 (n26422, pi0753, n_19140);
  not g42556 (n_19141, n26421);
  and g42557 (n26423, n_19141, n26422);
  and g42558 (n26424, n_6015, n17629);
  and g42559 (n26425, pi0180, n17631);
  not g42560 (n_19142, n26425);
  and g42561 (n26426, n_15488, n_19142);
  not g42562 (n_19143, n26424);
  and g42563 (n26427, n_19143, n26426);
  not g42564 (n_19144, n26423);
  not g42565 (n_19145, n26427);
  and g42566 (n26428, n_19144, n_19145);
  not g42567 (n_19146, n26428);
  and g42568 (n26429, n_162, n_19146);
  and g42569 (n26430, pi0180, n17605);
  and g42570 (n26431, n_6015, n_12180);
  not g42571 (n_19147, n26431);
  and g42572 (n26432, n_15488, n_19147);
  not g42573 (n_19148, n26430);
  and g42574 (n26433, n_19148, n26432);
  and g42575 (n26434, n_6015, n17404);
  and g42576 (n26435, pi0180, n17485);
  not g42577 (n_19149, n26435);
  and g42578 (n26436, pi0753, n_19149);
  not g42579 (n_19150, n26434);
  and g42580 (n26437, n_19150, n26436);
  not g42581 (n_19151, n26433);
  and g42582 (n26438, pi0039, n_19151);
  not g42583 (n_19152, n26437);
  and g42584 (n26439, n_19152, n26438);
  not g42585 (n_19153, n26429);
  and g42586 (n26440, n_161, n_19153);
  not g42587 (n_19154, n26439);
  and g42588 (n26441, n_19154, n26440);
  and g42589 (n26442, n_12120, n_18876);
  not g42590 (n_19155, n26442);
  and g42591 (n26443, pi0180, n_19155);
  and g42592 (n26444, n6284, n26443);
  and g42593 (n26445, n_15488, n_12250);
  not g42594 (n_19156, n26445);
  and g42595 (n26446, n19471, n_19156);
  not g42596 (n_19157, n26446);
  and g42597 (n26447, n_6015, n_19157);
  not g42598 (n_19158, n26444);
  and g42599 (n26448, pi0038, n_19158);
  not g42600 (n_19159, n26447);
  and g42601 (n26449, n_19159, n26448);
  not g42602 (n_19160, n26449);
  and g42603 (n26450, n_15518, n_19160);
  not g42604 (n_19161, n26441);
  and g42605 (n26451, n_19161, n26450);
  and g42606 (n26452, pi0702, n26346);
  not g42607 (n_19162, n26451);
  and g42608 (n26453, n2571, n_19162);
  not g42609 (n_19163, n26452);
  and g42610 (n26454, n_19163, n26453);
  not g42611 (n_19164, n26454);
  and g42612 (n26455, n_19078, n_19164);
  and g42613 (n26456, n_11753, n26455);
  and g42614 (n26457, pi0625, n26348);
  not g42615 (n_19165, n26457);
  and g42616 (n26458, n_11757, n_19165);
  not g42617 (n_19166, n26456);
  and g42618 (n26459, n_19166, n26458);
  and g42619 (n26460, n_11823, n_19028);
  not g42620 (n_19167, n26459);
  and g42621 (n26461, n_19167, n26460);
  and g42622 (n26462, n_11753, n26348);
  and g42623 (n26463, pi0625, n26455);
  not g42624 (n_19168, n26462);
  and g42625 (n26464, pi1153, n_19168);
  not g42626 (n_19169, n26463);
  and g42627 (n26465, n_19169, n26464);
  and g42628 (n26466, pi0608, n_19029);
  not g42629 (n_19170, n26465);
  and g42630 (n26467, n_19170, n26466);
  not g42631 (n_19171, n26461);
  not g42632 (n_19172, n26467);
  and g42633 (n26468, n_19171, n_19172);
  not g42634 (n_19173, n26468);
  and g42635 (n26469, pi0778, n_19173);
  and g42636 (n26470, n_11749, n26455);
  not g42637 (n_19174, n26469);
  not g42638 (n_19175, n26470);
  and g42639 (n26471, n_19174, n_19175);
  not g42640 (n_19176, n26471);
  and g42641 (n26472, n_11971, n_19176);
  not g42642 (n_19177, n26419);
  and g42643 (n26473, n_11768, n_19177);
  not g42644 (n_19178, n26472);
  and g42645 (n26474, n_19178, n26473);
  and g42646 (n26475, n_11767, n_19090);
  not g42647 (n_19179, n26474);
  and g42648 (n26476, n_19179, n26475);
  and g42649 (n26477, n_11971, n26290);
  and g42650 (n26478, pi0609, n_19176);
  not g42651 (n_19180, n26477);
  and g42652 (n26479, pi1155, n_19180);
  not g42653 (n_19181, n26478);
  and g42654 (n26480, n_19181, n26479);
  and g42655 (n26481, pi0660, n_19091);
  not g42656 (n_19182, n26480);
  and g42657 (n26482, n_19182, n26481);
  not g42658 (n_19183, n26476);
  not g42659 (n_19184, n26482);
  and g42660 (n26483, n_19183, n_19184);
  not g42661 (n_19185, n26483);
  and g42662 (n26484, pi0785, n_19185);
  and g42663 (n26485, n_11964, n_19176);
  not g42664 (n_19186, n26484);
  not g42665 (n_19187, n26485);
  and g42666 (n26486, n_19186, n_19187);
  not g42667 (n_19188, n26486);
  and g42668 (n26487, n_11984, n_19188);
  and g42669 (n26488, pi0618, n26293);
  not g42670 (n_19189, n26488);
  and g42671 (n26489, n_11413, n_19189);
  not g42672 (n_19190, n26487);
  and g42673 (n26490, n_19190, n26489);
  and g42674 (n26491, n_11412, n_19100);
  not g42675 (n_19191, n26490);
  and g42676 (n26492, n_19191, n26491);
  and g42677 (n26493, n_11984, n26293);
  and g42678 (n26494, pi0618, n_19188);
  not g42679 (n_19192, n26493);
  and g42680 (n26495, pi1154, n_19192);
  not g42681 (n_19193, n26494);
  and g42682 (n26496, n_19193, n26495);
  and g42683 (n26497, pi0627, n_19101);
  not g42684 (n_19194, n26496);
  and g42685 (n26498, n_19194, n26497);
  not g42686 (n_19195, n26492);
  not g42687 (n_19196, n26498);
  and g42688 (n26499, n_19195, n_19196);
  not g42689 (n_19197, n26499);
  and g42690 (n26500, pi0781, n_19197);
  and g42691 (n26501, n_11981, n_19188);
  not g42692 (n_19198, n26500);
  not g42693 (n_19199, n26501);
  and g42694 (n26502, n_19198, n_19199);
  and g42695 (n26503, n_12315, n26502);
  not g42696 (n_19200, n26296);
  and g42697 (n26504, pi0619, n_19200);
  not g42698 (n_19201, n26502);
  and g42699 (n26505, n_11821, n_19201);
  not g42700 (n_19202, n26504);
  and g42701 (n26506, n_11405, n_19202);
  not g42702 (n_19203, n26505);
  and g42703 (n26507, n_19203, n26506);
  and g42704 (n26508, n_11403, n_19110);
  not g42705 (n_19204, n26507);
  and g42706 (n26509, n_19204, n26508);
  and g42707 (n26510, n_11821, n_19200);
  and g42708 (n26511, pi0619, n_19201);
  not g42709 (n_19205, n26510);
  and g42710 (n26512, pi1159, n_19205);
  not g42711 (n_19206, n26511);
  and g42712 (n26513, n_19206, n26512);
  and g42713 (n26514, pi0648, n_19111);
  not g42714 (n_19207, n26513);
  and g42715 (n26515, n_19207, n26514);
  not g42716 (n_19208, n26509);
  and g42717 (n26516, pi0789, n_19208);
  not g42718 (n_19209, n26515);
  and g42719 (n26517, n_19209, n26516);
  not g42720 (n_19210, n26503);
  and g42721 (n26518, n17970, n_19210);
  not g42722 (n_19211, n26517);
  and g42723 (n26519, n_19211, n26518);
  and g42724 (n26520, n17871, n26298);
  not g42725 (n_19212, n26387);
  and g42726 (n26521, n_12320, n_19212);
  and g42727 (n26522, pi0626, n_19012);
  not g42728 (n_19213, n26522);
  and g42729 (n26523, n16629, n_19213);
  not g42730 (n_19214, n26521);
  and g42731 (n26524, n_19214, n26523);
  and g42732 (n26525, pi0626, n_19212);
  and g42733 (n26526, n_12320, n_19012);
  not g42734 (n_19215, n26526);
  and g42735 (n26527, n16628, n_19215);
  not g42736 (n_19216, n26525);
  and g42737 (n26528, n_19216, n26527);
  not g42738 (n_19217, n26520);
  not g42739 (n_19218, n26524);
  and g42740 (n26529, n_19217, n_19218);
  not g42741 (n_19219, n26528);
  and g42742 (n26530, n_19219, n26529);
  not g42743 (n_19220, n26530);
  and g42744 (n26531, pi0788, n_19220);
  not g42745 (n_19221, n26531);
  and g42746 (n26532, n_14638, n_19221);
  not g42747 (n_19222, n26519);
  and g42748 (n26533, n_19222, n26532);
  not g42749 (n_19223, n26418);
  not g42750 (n_19224, n26533);
  and g42751 (n26534, n_19223, n_19224);
  not g42752 (n_19225, n26534);
  and g42753 (n26535, n_14387, n_19225);
  not g42754 (n_19226, n26316);
  and g42755 (n26536, n17802, n_19226);
  and g42756 (n26537, n_14548, n26393);
  not g42757 (n_19227, n26320);
  and g42758 (n26538, n17801, n_19227);
  not g42759 (n_19228, n26536);
  not g42760 (n_19229, n26538);
  and g42761 (n26539, n_19228, n_19229);
  not g42762 (n_19230, n26537);
  and g42763 (n26540, n_19230, n26539);
  not g42764 (n_19231, n26540);
  and g42765 (n26541, pi0787, n_19231);
  and g42766 (n26542, n_11819, n26409);
  and g42767 (n26543, pi0644, n26401);
  not g42768 (n_19232, n26542);
  and g42769 (n26544, pi0790, n_19232);
  not g42770 (n_19233, n26543);
  and g42771 (n26545, n_19233, n26544);
  not g42772 (n_19234, n26535);
  not g42773 (n_19235, n26541);
  and g42774 (n26546, n_19234, n_19235);
  not g42775 (n_19236, n26545);
  and g42776 (n26547, n_19236, n26546);
  not g42777 (n_19237, n26412);
  not g42778 (n_19238, n26547);
  and g42779 (n26548, n_19237, n_19238);
  not g42780 (n_19239, n26548);
  and g42781 (n26549, n_4226, n_19239);
  not g42782 (n_19240, n26264);
  and g42783 (n26550, n_12415, n_19240);
  not g42784 (n_19241, n26549);
  and g42785 (n26551, n_19241, n26550);
  not g42786 (n_19242, n26263);
  not g42787 (n_19243, n26551);
  and g42788 (po0337, n_19242, n_19243);
  and g42789 (n26553, n_6429, n_12418);
  and g42790 (n26554, n_15563, n16645);
  not g42791 (n_19244, n26553);
  not g42792 (n_19245, n26554);
  and g42793 (n26555, n_19244, n_19245);
  not g42794 (n_19246, n26555);
  and g42795 (n26556, n_11749, n_19246);
  and g42796 (n26557, n_11753, n26554);
  not g42797 (n_19247, n26557);
  and g42798 (n26558, n_19246, n_19247);
  not g42799 (n_19248, n26558);
  and g42800 (n26559, pi1153, n_19248);
  and g42801 (n26560, n_11757, n_19244);
  and g42802 (n26561, n_19247, n26560);
  not g42803 (n_19249, n26561);
  and g42804 (n26562, pi0778, n_19249);
  not g42805 (n_19250, n26559);
  and g42806 (n26563, n_19250, n26562);
  not g42807 (n_19251, n26556);
  not g42808 (n_19252, n26563);
  and g42809 (n26564, n_19251, n_19252);
  not g42810 (n_19253, n26564);
  and g42811 (n26565, n_12429, n_19253);
  and g42812 (n26566, n_12430, n26565);
  and g42813 (n26567, n_12431, n26566);
  and g42814 (n26568, n_12432, n26567);
  and g42815 (n26569, n_12436, n26568);
  and g42816 (n26570, n_11806, n26569);
  and g42817 (n26571, pi0647, n26553);
  not g42818 (n_19254, n26571);
  and g42819 (n26572, n_11810, n_19254);
  not g42820 (n_19255, n26570);
  and g42821 (n26573, n_19255, n26572);
  and g42822 (n26574, pi0630, n26573);
  and g42823 (n26575, n_15533, n17244);
  not g42824 (n_19256, n26575);
  and g42825 (n26576, n_19244, n_19256);
  not g42826 (n_19257, n26576);
  and g42827 (n26577, n_12448, n_19257);
  not g42828 (n_19258, n26577);
  and g42829 (n26578, n_11964, n_19258);
  and g42830 (n26579, n17296, n26575);
  not g42831 (n_19259, n26579);
  and g42832 (n26580, n26577, n_19259);
  not g42833 (n_19260, n26580);
  and g42834 (n26581, pi1155, n_19260);
  and g42835 (n26582, n_11768, n_19244);
  and g42836 (n26583, n_19259, n26582);
  not g42837 (n_19261, n26581);
  not g42838 (n_19262, n26583);
  and g42839 (n26584, n_19261, n_19262);
  not g42840 (n_19263, n26584);
  and g42841 (n26585, pi0785, n_19263);
  not g42842 (n_19264, n26578);
  not g42843 (n_19265, n26585);
  and g42844 (n26586, n_19264, n_19265);
  not g42845 (n_19266, n26586);
  and g42846 (n26587, n_11981, n_19266);
  and g42847 (n26588, n_12461, n26586);
  not g42848 (n_19267, n26588);
  and g42849 (n26589, pi1154, n_19267);
  and g42850 (n26590, n_12463, n26586);
  not g42851 (n_19268, n26590);
  and g42852 (n26591, n_11413, n_19268);
  not g42853 (n_19269, n26589);
  not g42854 (n_19270, n26591);
  and g42855 (n26592, n_19269, n_19270);
  not g42856 (n_19271, n26592);
  and g42857 (n26593, pi0781, n_19271);
  not g42858 (n_19272, n26587);
  not g42859 (n_19273, n26593);
  and g42860 (n26594, n_19272, n_19273);
  not g42861 (n_19274, n26594);
  and g42862 (n26595, n_12315, n_19274);
  and g42863 (n26596, n_16503, n26594);
  not g42864 (n_19275, n26596);
  and g42865 (n26597, pi1159, n_19275);
  and g42866 (n26598, n_16505, n26594);
  not g42867 (n_19276, n26598);
  and g42868 (n26599, n_11405, n_19276);
  not g42869 (n_19277, n26597);
  not g42870 (n_19278, n26599);
  and g42871 (n26600, n_19277, n_19278);
  not g42872 (n_19279, n26600);
  and g42873 (n26601, pi0789, n_19279);
  not g42874 (n_19280, n26595);
  not g42875 (n_19281, n26601);
  and g42876 (n26602, n_19280, n_19281);
  and g42877 (n26603, n_12524, n26602);
  and g42878 (n26604, n17969, n26553);
  not g42879 (n_19282, n26603);
  not g42880 (n_19283, n26604);
  and g42881 (n26605, n_19282, n_19283);
  not g42882 (n_19284, n26605);
  and g42883 (n26606, n_12368, n_19284);
  and g42884 (n26607, n17779, n26553);
  not g42885 (n_19285, n26606);
  not g42886 (n_19286, n26607);
  and g42887 (n26608, n_19285, n_19286);
  and g42888 (n26609, n_14548, n26608);
  not g42889 (n_19287, n26569);
  and g42890 (n26610, pi0647, n_19287);
  and g42891 (n26611, n_11806, n_19244);
  not g42892 (n_19288, n26610);
  not g42893 (n_19289, n26611);
  and g42894 (n26612, n_19288, n_19289);
  not g42895 (n_19290, n26612);
  and g42896 (n26613, n17801, n_19290);
  not g42897 (n_19291, n26574);
  not g42898 (n_19292, n26613);
  and g42899 (n26614, n_19291, n_19292);
  not g42900 (n_19293, n26609);
  and g42901 (n26615, n_19293, n26614);
  not g42902 (n_19294, n26615);
  and g42903 (n26616, pi0787, n_19294);
  and g42904 (n26617, n17871, n26567);
  not g42905 (n_19295, n26602);
  and g42906 (n26618, n_12320, n_19295);
  and g42907 (n26619, pi0626, n_19244);
  not g42908 (n_19296, n26619);
  and g42909 (n26620, n16629, n_19296);
  not g42910 (n_19297, n26618);
  and g42911 (n26621, n_19297, n26620);
  and g42912 (n26622, pi0626, n_19295);
  and g42913 (n26623, n_12320, n_19244);
  not g42914 (n_19298, n26623);
  and g42915 (n26624, n16628, n_19298);
  not g42916 (n_19299, n26622);
  and g42917 (n26625, n_19299, n26624);
  not g42918 (n_19300, n26617);
  not g42919 (n_19301, n26621);
  and g42920 (n26626, n_19300, n_19301);
  not g42921 (n_19302, n26625);
  and g42922 (n26627, n_19302, n26626);
  not g42923 (n_19303, n26627);
  and g42924 (n26628, pi0788, n_19303);
  and g42925 (n26629, pi0618, n26565);
  and g42926 (n26630, n_11866, n_19246);
  and g42927 (n26631, pi0625, n26630);
  not g42928 (n_19304, n26630);
  and g42929 (n26632, n26576, n_19304);
  not g42930 (n_19305, n26631);
  not g42931 (n_19306, n26632);
  and g42932 (n26633, n_19305, n_19306);
  not g42933 (n_19307, n26633);
  and g42934 (n26634, n26560, n_19307);
  and g42935 (n26635, n_11823, n_19250);
  not g42936 (n_19308, n26634);
  and g42937 (n26636, n_19308, n26635);
  and g42938 (n26637, pi1153, n26576);
  and g42939 (n26638, n_19305, n26637);
  and g42940 (n26639, pi0608, n_19249);
  not g42941 (n_19309, n26638);
  and g42942 (n26640, n_19309, n26639);
  not g42943 (n_19310, n26636);
  not g42944 (n_19311, n26640);
  and g42945 (n26641, n_19310, n_19311);
  not g42946 (n_19312, n26641);
  and g42947 (n26642, pi0778, n_19312);
  and g42948 (n26643, n_11749, n_19306);
  not g42949 (n_19313, n26642);
  not g42950 (n_19314, n26643);
  and g42951 (n26644, n_19313, n_19314);
  not g42952 (n_19315, n26644);
  and g42953 (n26645, n_11971, n_19315);
  and g42954 (n26646, pi0609, n_19253);
  not g42955 (n_19316, n26646);
  and g42956 (n26647, n_11768, n_19316);
  not g42957 (n_19317, n26645);
  and g42958 (n26648, n_19317, n26647);
  and g42959 (n26649, n_11767, n_19261);
  not g42960 (n_19318, n26648);
  and g42961 (n26650, n_19318, n26649);
  and g42962 (n26651, pi0609, n_19315);
  and g42963 (n26652, n_11971, n_19253);
  not g42964 (n_19319, n26652);
  and g42965 (n26653, pi1155, n_19319);
  not g42966 (n_19320, n26651);
  and g42967 (n26654, n_19320, n26653);
  and g42968 (n26655, pi0660, n_19262);
  not g42969 (n_19321, n26654);
  and g42970 (n26656, n_19321, n26655);
  not g42971 (n_19322, n26650);
  not g42972 (n_19323, n26656);
  and g42973 (n26657, n_19322, n_19323);
  not g42974 (n_19324, n26657);
  and g42975 (n26658, pi0785, n_19324);
  and g42976 (n26659, n_11964, n_19315);
  not g42977 (n_19325, n26658);
  not g42978 (n_19326, n26659);
  and g42979 (n26660, n_19325, n_19326);
  not g42980 (n_19327, n26660);
  and g42981 (n26661, n_11984, n_19327);
  not g42982 (n_19328, n26629);
  and g42983 (n26662, n_11413, n_19328);
  not g42984 (n_19329, n26661);
  and g42985 (n26663, n_19329, n26662);
  and g42986 (n26664, n_11412, n_19269);
  not g42987 (n_19330, n26663);
  and g42988 (n26665, n_19330, n26664);
  and g42989 (n26666, n_11984, n26565);
  and g42990 (n26667, pi0618, n_19327);
  not g42991 (n_19331, n26666);
  and g42992 (n26668, pi1154, n_19331);
  not g42993 (n_19332, n26667);
  and g42994 (n26669, n_19332, n26668);
  and g42995 (n26670, pi0627, n_19270);
  not g42996 (n_19333, n26669);
  and g42997 (n26671, n_19333, n26670);
  not g42998 (n_19334, n26665);
  not g42999 (n_19335, n26671);
  and g43000 (n26672, n_19334, n_19335);
  not g43001 (n_19336, n26672);
  and g43002 (n26673, pi0781, n_19336);
  and g43003 (n26674, n_11981, n_19327);
  not g43004 (n_19337, n26673);
  not g43005 (n_19338, n26674);
  and g43006 (n26675, n_19337, n_19338);
  and g43007 (n26676, n_12315, n26675);
  not g43008 (n_19339, n26675);
  and g43009 (n26677, n_11821, n_19339);
  and g43010 (n26678, pi0619, n26566);
  not g43011 (n_19340, n26678);
  and g43012 (n26679, n_11405, n_19340);
  not g43013 (n_19341, n26677);
  and g43014 (n26680, n_19341, n26679);
  and g43015 (n26681, n_11403, n_19277);
  not g43016 (n_19342, n26680);
  and g43017 (n26682, n_19342, n26681);
  and g43018 (n26683, pi0619, n_19339);
  and g43019 (n26684, n_11821, n26566);
  not g43020 (n_19343, n26684);
  and g43021 (n26685, pi1159, n_19343);
  not g43022 (n_19344, n26683);
  and g43023 (n26686, n_19344, n26685);
  and g43024 (n26687, pi0648, n_19278);
  not g43025 (n_19345, n26686);
  and g43026 (n26688, n_19345, n26687);
  not g43027 (n_19346, n26682);
  and g43028 (n26689, pi0789, n_19346);
  not g43029 (n_19347, n26688);
  and g43030 (n26690, n_19347, n26689);
  not g43031 (n_19348, n26676);
  and g43032 (n26691, n17970, n_19348);
  not g43033 (n_19349, n26690);
  and g43034 (n26692, n_19349, n26691);
  not g43035 (n_19350, n26628);
  not g43036 (n_19351, n26692);
  and g43037 (n26693, n_19350, n_19351);
  not g43038 (n_19352, n26693);
  and g43039 (n26694, n_14638, n_19352);
  and g43040 (n26695, n17854, n_19284);
  and g43041 (n26696, n20851, n26568);
  not g43042 (n_19353, n26695);
  not g43043 (n_19354, n26696);
  and g43044 (n26697, n_19353, n_19354);
  not g43045 (n_19355, n26697);
  and g43046 (n26698, n_12354, n_19355);
  and g43047 (n26699, n20855, n26568);
  and g43048 (n26700, n17853, n_19284);
  not g43049 (n_19356, n26699);
  not g43050 (n_19357, n26700);
  and g43051 (n26701, n_19356, n_19357);
  not g43052 (n_19358, n26701);
  and g43053 (n26702, pi0629, n_19358);
  not g43054 (n_19359, n26698);
  not g43055 (n_19360, n26702);
  and g43056 (n26703, n_19359, n_19360);
  not g43057 (n_19361, n26703);
  and g43058 (n26704, pi0792, n_19361);
  not g43059 (n_19362, n26704);
  and g43060 (n26705, n_14387, n_19362);
  not g43061 (n_19363, n26694);
  and g43062 (n26706, n_19363, n26705);
  not g43063 (n_19364, n26616);
  not g43064 (n_19365, n26706);
  and g43065 (n26707, n_19364, n_19365);
  and g43066 (n26708, n_12411, n26707);
  and g43067 (n26709, n_11803, n_19287);
  and g43068 (n26710, pi1157, n_19290);
  not g43069 (n_19366, n26573);
  not g43070 (n_19367, n26710);
  and g43071 (n26711, n_19366, n_19367);
  not g43072 (n_19368, n26711);
  and g43073 (n26712, pi0787, n_19368);
  not g43074 (n_19369, n26709);
  not g43075 (n_19370, n26712);
  and g43076 (n26713, n_19369, n_19370);
  and g43077 (n26714, n_11819, n26713);
  and g43078 (n26715, pi0644, n26707);
  not g43079 (n_19371, n26714);
  and g43080 (n26716, pi0715, n_19371);
  not g43081 (n_19372, n26715);
  and g43082 (n26717, n_19372, n26716);
  not g43083 (n_19373, n26608);
  and g43084 (n26718, n_12392, n_19373);
  and g43085 (n26719, n17804, n26553);
  not g43086 (n_19374, n26718);
  not g43087 (n_19375, n26719);
  and g43088 (n26720, n_19374, n_19375);
  not g43089 (n_19376, n26720);
  and g43090 (n26721, pi0644, n_19376);
  and g43091 (n26722, n_11819, n26553);
  not g43092 (n_19377, n26722);
  and g43093 (n26723, n_12395, n_19377);
  not g43094 (n_19378, n26721);
  and g43095 (n26724, n_19378, n26723);
  not g43096 (n_19379, n26724);
  and g43097 (n26725, pi1160, n_19379);
  not g43098 (n_19380, n26717);
  and g43099 (n26726, n_19380, n26725);
  and g43100 (n26727, n_11819, n_19376);
  and g43101 (n26728, pi0644, n26553);
  not g43102 (n_19381, n26728);
  and g43103 (n26729, pi0715, n_19381);
  not g43104 (n_19382, n26727);
  and g43105 (n26730, n_19382, n26729);
  and g43106 (n26731, pi0644, n26713);
  and g43107 (n26732, n_11819, n26707);
  not g43108 (n_19383, n26731);
  and g43109 (n26733, n_12395, n_19383);
  not g43110 (n_19384, n26732);
  and g43111 (n26734, n_19384, n26733);
  not g43112 (n_19385, n26730);
  and g43113 (n26735, n_12405, n_19385);
  not g43114 (n_19386, n26734);
  and g43115 (n26736, n_19386, n26735);
  not g43116 (n_19387, n26726);
  not g43117 (n_19388, n26736);
  and g43118 (n26737, n_19387, n_19388);
  not g43119 (n_19389, n26737);
  and g43120 (n26738, pi0790, n_19389);
  not g43121 (n_19390, n26708);
  and g43122 (n26739, pi0832, n_19390);
  not g43123 (n_19391, n26738);
  and g43124 (n26740, n_19391, n26739);
  and g43125 (n26741, n_6429, po1038);
  and g43126 (n26742, n_6429, n_11751);
  not g43127 (n_19392, n26742);
  and g43128 (n26743, n16635, n_19392);
  and g43129 (n26744, n_15563, n2571);
  not g43130 (n_19393, n26744);
  and g43131 (n26745, n26742, n_19393);
  and g43132 (n26746, n_6429, n_11418);
  not g43133 (n_19394, n26746);
  and g43134 (n26747, n16647, n_19394);
  and g43135 (n26748, pi0181, n_12608);
  not g43136 (n_19395, n26748);
  and g43137 (n26749, n_161, n_19395);
  not g43138 (n_19396, n26749);
  and g43139 (n26750, n2571, n_19396);
  and g43140 (n26751, n_6429, n18072);
  not g43141 (n_19397, n26750);
  not g43142 (n_19398, n26751);
  and g43143 (n26752, n_19397, n_19398);
  not g43144 (n_19399, n26747);
  and g43145 (n26753, n_15563, n_19399);
  not g43146 (n_19400, n26752);
  and g43147 (n26754, n_19400, n26753);
  not g43148 (n_19401, n26745);
  not g43149 (n_19402, n26754);
  and g43150 (n26755, n_19401, n_19402);
  and g43151 (n26756, n_11749, n26755);
  and g43152 (n26757, n_11753, n26742);
  not g43153 (n_19403, n26755);
  and g43154 (n26758, pi0625, n_19403);
  not g43155 (n_19404, n26757);
  and g43156 (n26759, pi1153, n_19404);
  not g43157 (n_19405, n26758);
  and g43158 (n26760, n_19405, n26759);
  and g43159 (n26761, pi0625, n26742);
  and g43160 (n26762, n_11753, n_19403);
  not g43161 (n_19406, n26761);
  and g43162 (n26763, n_11757, n_19406);
  not g43163 (n_19407, n26762);
  and g43164 (n26764, n_19407, n26763);
  not g43165 (n_19408, n26760);
  not g43166 (n_19409, n26764);
  and g43167 (n26765, n_19408, n_19409);
  not g43168 (n_19410, n26765);
  and g43169 (n26766, pi0778, n_19410);
  not g43170 (n_19411, n26756);
  not g43171 (n_19412, n26766);
  and g43172 (n26767, n_19411, n_19412);
  not g43173 (n_19413, n26767);
  and g43174 (n26768, n_11773, n_19413);
  and g43175 (n26769, n17075, n_19392);
  not g43176 (n_19414, n26768);
  not g43177 (n_19415, n26769);
  and g43178 (n26770, n_19414, n_19415);
  and g43179 (n26771, n_11777, n26770);
  and g43180 (n26772, n16639, n26742);
  not g43181 (n_19416, n26771);
  not g43182 (n_19417, n26772);
  and g43183 (n26773, n_19416, n_19417);
  and g43184 (n26774, n_11780, n26773);
  not g43185 (n_19418, n26743);
  not g43186 (n_19419, n26774);
  and g43187 (n26775, n_19418, n_19419);
  and g43188 (n26776, n_11783, n26775);
  and g43189 (n26777, n16631, n26742);
  not g43190 (n_19420, n26776);
  not g43191 (n_19421, n26777);
  and g43192 (n26778, n_19420, n_19421);
  and g43193 (n26779, n_11787, n26778);
  not g43194 (n_19422, n26778);
  and g43195 (n26780, pi0628, n_19422);
  and g43196 (n26781, n_11789, n26742);
  not g43197 (n_19423, n26781);
  and g43198 (n26782, pi1156, n_19423);
  not g43199 (n_19424, n26780);
  and g43200 (n26783, n_19424, n26782);
  and g43201 (n26784, pi0628, n26742);
  and g43202 (n26785, n_11789, n_19422);
  not g43203 (n_19425, n26784);
  and g43204 (n26786, n_11794, n_19425);
  not g43205 (n_19426, n26785);
  and g43206 (n26787, n_19426, n26786);
  not g43207 (n_19427, n26783);
  not g43208 (n_19428, n26787);
  and g43209 (n26788, n_19427, n_19428);
  not g43210 (n_19429, n26788);
  and g43211 (n26789, pi0792, n_19429);
  not g43212 (n_19430, n26779);
  not g43213 (n_19431, n26789);
  and g43214 (n26790, n_19430, n_19431);
  not g43215 (n_19432, n26790);
  and g43216 (n26791, n_11806, n_19432);
  and g43217 (n26792, pi0647, n_19392);
  not g43218 (n_19433, n26791);
  not g43219 (n_19434, n26792);
  and g43220 (n26793, n_19433, n_19434);
  and g43221 (n26794, n_11810, n26793);
  and g43222 (n26795, pi0647, n_19432);
  and g43223 (n26796, n_11806, n_19392);
  not g43224 (n_19435, n26795);
  not g43225 (n_19436, n26796);
  and g43226 (n26797, n_19435, n_19436);
  and g43227 (n26798, pi1157, n26797);
  not g43228 (n_19437, n26794);
  not g43229 (n_19438, n26798);
  and g43230 (n26799, n_19437, n_19438);
  not g43231 (n_19439, n26799);
  and g43232 (n26800, pi0787, n_19439);
  and g43233 (n26801, n_11803, n26790);
  not g43234 (n_19440, n26800);
  not g43235 (n_19441, n26801);
  and g43236 (n26802, n_19440, n_19441);
  not g43237 (n_19442, n26802);
  and g43238 (n26803, n_11819, n_19442);
  not g43239 (n_19443, n26803);
  and g43240 (n26804, pi0715, n_19443);
  and g43241 (n26805, pi0181, n_11417);
  and g43242 (n26806, pi0181, pi0754);
  and g43243 (n26807, pi0754, n17046);
  and g43244 (n26808, pi0181, n17273);
  not g43245 (n_19444, n26807);
  not g43246 (n_19445, n26808);
  and g43247 (n26809, n_19444, n_19445);
  not g43248 (n_19446, n26809);
  and g43249 (n26810, pi0039, n_19446);
  and g43250 (n26811, pi0181, n_11923);
  not g43251 (n_19447, n26811);
  and g43252 (n26812, n_15539, n_19447);
  not g43253 (n_19448, n26812);
  and g43254 (n26813, n_162, n_19448);
  and g43255 (n26814, n_6429, n_15533);
  and g43256 (n26815, n17221, n26814);
  not g43264 (n_19453, n26818);
  and g43265 (n26819, n_161, n_19453);
  and g43266 (n26820, n_15533, n17280);
  and g43267 (n26821, pi0038, n_19394);
  not g43268 (n_19454, n26820);
  and g43269 (n26822, n_19454, n26821);
  not g43270 (n_19455, n26819);
  not g43271 (n_19456, n26822);
  and g43272 (n26823, n_19455, n_19456);
  not g43273 (n_19457, n26823);
  and g43274 (n26824, n2571, n_19457);
  not g43275 (n_19458, n26805);
  not g43276 (n_19459, n26824);
  and g43277 (n26825, n_19458, n_19459);
  not g43278 (n_19460, n26825);
  and g43279 (n26826, n_11960, n_19460);
  and g43280 (n26827, n17117, n_19392);
  not g43281 (n_19461, n26826);
  not g43282 (n_19462, n26827);
  and g43283 (n26828, n_19461, n_19462);
  not g43284 (n_19463, n26828);
  and g43285 (n26829, n_11964, n_19463);
  and g43286 (n26830, n_11967, n_19392);
  and g43287 (n26831, pi0609, n26826);
  not g43288 (n_19464, n26830);
  not g43289 (n_19465, n26831);
  and g43290 (n26832, n_19464, n_19465);
  not g43291 (n_19466, n26832);
  and g43292 (n26833, pi1155, n_19466);
  and g43293 (n26834, n_11972, n_19392);
  and g43294 (n26835, n_11971, n26826);
  not g43295 (n_19467, n26834);
  not g43296 (n_19468, n26835);
  and g43297 (n26836, n_19467, n_19468);
  not g43298 (n_19469, n26836);
  and g43299 (n26837, n_11768, n_19469);
  not g43300 (n_19470, n26833);
  not g43301 (n_19471, n26837);
  and g43302 (n26838, n_19470, n_19471);
  not g43303 (n_19472, n26838);
  and g43304 (n26839, pi0785, n_19472);
  not g43305 (n_19473, n26829);
  not g43306 (n_19474, n26839);
  and g43307 (n26840, n_19473, n_19474);
  not g43308 (n_19475, n26840);
  and g43309 (n26841, n_11981, n_19475);
  and g43310 (n26842, n_11984, n26742);
  and g43311 (n26843, pi0618, n26840);
  not g43312 (n_19476, n26842);
  and g43313 (n26844, pi1154, n_19476);
  not g43314 (n_19477, n26843);
  and g43315 (n26845, n_19477, n26844);
  and g43316 (n26846, n_11984, n26840);
  and g43317 (n26847, pi0618, n26742);
  not g43318 (n_19478, n26847);
  and g43319 (n26848, n_11413, n_19478);
  not g43320 (n_19479, n26846);
  and g43321 (n26849, n_19479, n26848);
  not g43322 (n_19480, n26845);
  not g43323 (n_19481, n26849);
  and g43324 (n26850, n_19480, n_19481);
  not g43325 (n_19482, n26850);
  and g43326 (n26851, pi0781, n_19482);
  not g43327 (n_19483, n26841);
  not g43328 (n_19484, n26851);
  and g43329 (n26852, n_19483, n_19484);
  not g43330 (n_19485, n26852);
  and g43331 (n26853, n_12315, n_19485);
  and g43332 (n26854, n_11821, n26742);
  and g43333 (n26855, pi0619, n26852);
  not g43334 (n_19486, n26854);
  and g43335 (n26856, pi1159, n_19486);
  not g43336 (n_19487, n26855);
  and g43337 (n26857, n_19487, n26856);
  and g43338 (n26858, n_11821, n26852);
  and g43339 (n26859, pi0619, n26742);
  not g43340 (n_19488, n26859);
  and g43341 (n26860, n_11405, n_19488);
  not g43342 (n_19489, n26858);
  and g43343 (n26861, n_19489, n26860);
  not g43344 (n_19490, n26857);
  not g43345 (n_19491, n26861);
  and g43346 (n26862, n_19490, n_19491);
  not g43347 (n_19492, n26862);
  and g43348 (n26863, pi0789, n_19492);
  not g43349 (n_19493, n26853);
  not g43350 (n_19494, n26863);
  and g43351 (n26864, n_19493, n_19494);
  and g43352 (n26865, n_12524, n26864);
  and g43353 (n26866, n17969, n26742);
  not g43354 (n_19495, n26865);
  not g43355 (n_19496, n26866);
  and g43356 (n26867, n_19495, n_19496);
  not g43357 (n_19497, n26867);
  and g43358 (n26868, n_12368, n_19497);
  and g43359 (n26869, n17779, n26742);
  not g43360 (n_19498, n26868);
  not g43361 (n_19499, n26869);
  and g43362 (n26870, n_19498, n_19499);
  not g43363 (n_19500, n26870);
  and g43364 (n26871, n_12392, n_19500);
  and g43365 (n26872, n17804, n26742);
  not g43366 (n_19501, n26871);
  not g43367 (n_19502, n26872);
  and g43368 (n26873, n_19501, n_19502);
  not g43369 (n_19503, n26873);
  and g43370 (n26874, pi0644, n_19503);
  and g43371 (n26875, n_11819, n26742);
  not g43372 (n_19504, n26875);
  and g43373 (n26876, n_12395, n_19504);
  not g43374 (n_19505, n26874);
  and g43375 (n26877, n_19505, n26876);
  not g43376 (n_19506, n26877);
  and g43377 (n26878, pi1160, n_19506);
  not g43378 (n_19507, n26804);
  and g43379 (n26879, n_19507, n26878);
  and g43380 (n26880, pi0644, n_19442);
  not g43381 (n_19508, n26880);
  and g43382 (n26881, n_12395, n_19508);
  and g43383 (n26882, n_11819, n_19503);
  and g43384 (n26883, pi0644, n26742);
  not g43385 (n_19509, n26883);
  and g43386 (n26884, pi0715, n_19509);
  not g43387 (n_19510, n26882);
  and g43388 (n26885, n_19510, n26884);
  not g43389 (n_19511, n26885);
  and g43390 (n26886, n_12405, n_19511);
  not g43391 (n_19512, n26881);
  and g43392 (n26887, n_19512, n26886);
  not g43393 (n_19513, n26879);
  not g43394 (n_19514, n26887);
  and g43395 (n26888, n_19513, n_19514);
  not g43396 (n_19515, n26888);
  and g43397 (n26889, pi0790, n_19515);
  and g43398 (n26890, n_12354, n26783);
  and g43399 (n26891, n_14557, n26867);
  and g43400 (n26892, pi0629, n26787);
  not g43401 (n_19516, n26890);
  not g43402 (n_19517, n26892);
  and g43403 (n26893, n_19516, n_19517);
  not g43404 (n_19518, n26891);
  and g43405 (n26894, n_19518, n26893);
  not g43406 (n_19519, n26894);
  and g43407 (n26895, pi0792, n_19519);
  and g43408 (n26896, pi0609, n26767);
  and g43409 (n26897, pi0181, n_12240);
  and g43410 (n26898, n_6429, n_12230);
  not g43411 (n_19520, n26897);
  and g43412 (n26899, pi0754, n_19520);
  not g43413 (n_19521, n26898);
  and g43414 (n26900, n_19521, n26899);
  and g43415 (n26901, n_6429, n17629);
  and g43416 (n26902, pi0181, n17631);
  not g43417 (n_19522, n26902);
  and g43418 (n26903, n_15533, n_19522);
  not g43419 (n_19523, n26901);
  and g43420 (n26904, n_19523, n26903);
  not g43421 (n_19524, n26900);
  not g43422 (n_19525, n26904);
  and g43423 (n26905, n_19524, n_19525);
  not g43424 (n_19526, n26905);
  and g43425 (n26906, n_162, n_19526);
  and g43426 (n26907, pi0181, n17605);
  and g43427 (n26908, n_6429, n_12180);
  not g43428 (n_19527, n26908);
  and g43429 (n26909, n_15533, n_19527);
  not g43430 (n_19528, n26907);
  and g43431 (n26910, n_19528, n26909);
  and g43432 (n26911, n_6429, n17404);
  and g43433 (n26912, pi0181, n17485);
  not g43434 (n_19529, n26912);
  and g43435 (n26913, pi0754, n_19529);
  not g43436 (n_19530, n26911);
  and g43437 (n26914, n_19530, n26913);
  not g43438 (n_19531, n26910);
  and g43439 (n26915, pi0039, n_19531);
  not g43440 (n_19532, n26914);
  and g43441 (n26916, n_19532, n26915);
  not g43442 (n_19533, n26906);
  and g43443 (n26917, n_161, n_19533);
  not g43444 (n_19534, n26916);
  and g43445 (n26918, n_19534, n26917);
  and g43446 (n26919, n_12120, n_19256);
  not g43447 (n_19535, n26919);
  and g43448 (n26920, pi0181, n_19535);
  and g43449 (n26921, n6284, n26920);
  and g43450 (n26922, n_15533, n_12250);
  not g43451 (n_19536, n26922);
  and g43452 (n26923, n19471, n_19536);
  not g43453 (n_19537, n26923);
  and g43454 (n26924, n_6429, n_19537);
  not g43455 (n_19538, n26921);
  and g43456 (n26925, pi0038, n_19538);
  not g43457 (n_19539, n26924);
  and g43458 (n26926, n_19539, n26925);
  not g43459 (n_19540, n26926);
  and g43460 (n26927, n_15563, n_19540);
  not g43461 (n_19541, n26918);
  and g43462 (n26928, n_19541, n26927);
  and g43463 (n26929, pi0709, n26823);
  not g43464 (n_19542, n26928);
  and g43465 (n26930, n2571, n_19542);
  not g43466 (n_19543, n26929);
  and g43467 (n26931, n_19543, n26930);
  not g43468 (n_19544, n26931);
  and g43469 (n26932, n_19458, n_19544);
  and g43470 (n26933, n_11753, n26932);
  and g43471 (n26934, pi0625, n26825);
  not g43472 (n_19545, n26934);
  and g43473 (n26935, n_11757, n_19545);
  not g43474 (n_19546, n26933);
  and g43475 (n26936, n_19546, n26935);
  and g43476 (n26937, n_11823, n_19408);
  not g43477 (n_19547, n26936);
  and g43478 (n26938, n_19547, n26937);
  and g43479 (n26939, n_11753, n26825);
  and g43480 (n26940, pi0625, n26932);
  not g43481 (n_19548, n26939);
  and g43482 (n26941, pi1153, n_19548);
  not g43483 (n_19549, n26940);
  and g43484 (n26942, n_19549, n26941);
  and g43485 (n26943, pi0608, n_19409);
  not g43486 (n_19550, n26942);
  and g43487 (n26944, n_19550, n26943);
  not g43488 (n_19551, n26938);
  not g43489 (n_19552, n26944);
  and g43490 (n26945, n_19551, n_19552);
  not g43491 (n_19553, n26945);
  and g43492 (n26946, pi0778, n_19553);
  and g43493 (n26947, n_11749, n26932);
  not g43494 (n_19554, n26946);
  not g43495 (n_19555, n26947);
  and g43496 (n26948, n_19554, n_19555);
  not g43497 (n_19556, n26948);
  and g43498 (n26949, n_11971, n_19556);
  not g43499 (n_19557, n26896);
  and g43500 (n26950, n_11768, n_19557);
  not g43501 (n_19558, n26949);
  and g43502 (n26951, n_19558, n26950);
  and g43503 (n26952, n_11767, n_19470);
  not g43504 (n_19559, n26951);
  and g43505 (n26953, n_19559, n26952);
  and g43506 (n26954, n_11971, n26767);
  and g43507 (n26955, pi0609, n_19556);
  not g43508 (n_19560, n26954);
  and g43509 (n26956, pi1155, n_19560);
  not g43510 (n_19561, n26955);
  and g43511 (n26957, n_19561, n26956);
  and g43512 (n26958, pi0660, n_19471);
  not g43513 (n_19562, n26957);
  and g43514 (n26959, n_19562, n26958);
  not g43515 (n_19563, n26953);
  not g43516 (n_19564, n26959);
  and g43517 (n26960, n_19563, n_19564);
  not g43518 (n_19565, n26960);
  and g43519 (n26961, pi0785, n_19565);
  and g43520 (n26962, n_11964, n_19556);
  not g43521 (n_19566, n26961);
  not g43522 (n_19567, n26962);
  and g43523 (n26963, n_19566, n_19567);
  not g43524 (n_19568, n26963);
  and g43525 (n26964, n_11984, n_19568);
  and g43526 (n26965, pi0618, n26770);
  not g43527 (n_19569, n26965);
  and g43528 (n26966, n_11413, n_19569);
  not g43529 (n_19570, n26964);
  and g43530 (n26967, n_19570, n26966);
  and g43531 (n26968, n_11412, n_19480);
  not g43532 (n_19571, n26967);
  and g43533 (n26969, n_19571, n26968);
  and g43534 (n26970, n_11984, n26770);
  and g43535 (n26971, pi0618, n_19568);
  not g43536 (n_19572, n26970);
  and g43537 (n26972, pi1154, n_19572);
  not g43538 (n_19573, n26971);
  and g43539 (n26973, n_19573, n26972);
  and g43540 (n26974, pi0627, n_19481);
  not g43541 (n_19574, n26973);
  and g43542 (n26975, n_19574, n26974);
  not g43543 (n_19575, n26969);
  not g43544 (n_19576, n26975);
  and g43545 (n26976, n_19575, n_19576);
  not g43546 (n_19577, n26976);
  and g43547 (n26977, pi0781, n_19577);
  and g43548 (n26978, n_11981, n_19568);
  not g43549 (n_19578, n26977);
  not g43550 (n_19579, n26978);
  and g43551 (n26979, n_19578, n_19579);
  and g43552 (n26980, n_12315, n26979);
  not g43553 (n_19580, n26773);
  and g43554 (n26981, pi0619, n_19580);
  not g43555 (n_19581, n26979);
  and g43556 (n26982, n_11821, n_19581);
  not g43557 (n_19582, n26981);
  and g43558 (n26983, n_11405, n_19582);
  not g43559 (n_19583, n26982);
  and g43560 (n26984, n_19583, n26983);
  and g43561 (n26985, n_11403, n_19490);
  not g43562 (n_19584, n26984);
  and g43563 (n26986, n_19584, n26985);
  and g43564 (n26987, n_11821, n_19580);
  and g43565 (n26988, pi0619, n_19581);
  not g43566 (n_19585, n26987);
  and g43567 (n26989, pi1159, n_19585);
  not g43568 (n_19586, n26988);
  and g43569 (n26990, n_19586, n26989);
  and g43570 (n26991, pi0648, n_19491);
  not g43571 (n_19587, n26990);
  and g43572 (n26992, n_19587, n26991);
  not g43573 (n_19588, n26986);
  and g43574 (n26993, pi0789, n_19588);
  not g43575 (n_19589, n26992);
  and g43576 (n26994, n_19589, n26993);
  not g43577 (n_19590, n26980);
  and g43578 (n26995, n17970, n_19590);
  not g43579 (n_19591, n26994);
  and g43580 (n26996, n_19591, n26995);
  and g43581 (n26997, n17871, n26775);
  not g43582 (n_19592, n26864);
  and g43583 (n26998, n_12320, n_19592);
  and g43584 (n26999, pi0626, n_19392);
  not g43585 (n_19593, n26999);
  and g43586 (n27000, n16629, n_19593);
  not g43587 (n_19594, n26998);
  and g43588 (n27001, n_19594, n27000);
  and g43589 (n27002, pi0626, n_19592);
  and g43590 (n27003, n_12320, n_19392);
  not g43591 (n_19595, n27003);
  and g43592 (n27004, n16628, n_19595);
  not g43593 (n_19596, n27002);
  and g43594 (n27005, n_19596, n27004);
  not g43595 (n_19597, n26997);
  not g43596 (n_19598, n27001);
  and g43597 (n27006, n_19597, n_19598);
  not g43598 (n_19599, n27005);
  and g43599 (n27007, n_19599, n27006);
  not g43600 (n_19600, n27007);
  and g43601 (n27008, pi0788, n_19600);
  not g43602 (n_19601, n27008);
  and g43603 (n27009, n_14638, n_19601);
  not g43604 (n_19602, n26996);
  and g43605 (n27010, n_19602, n27009);
  not g43606 (n_19603, n26895);
  not g43607 (n_19604, n27010);
  and g43608 (n27011, n_19603, n_19604);
  not g43609 (n_19605, n27011);
  and g43610 (n27012, n_14387, n_19605);
  not g43611 (n_19606, n26793);
  and g43612 (n27013, n17802, n_19606);
  and g43613 (n27014, n_14548, n26870);
  not g43614 (n_19607, n26797);
  and g43615 (n27015, n17801, n_19607);
  not g43616 (n_19608, n27013);
  not g43617 (n_19609, n27015);
  and g43618 (n27016, n_19608, n_19609);
  not g43619 (n_19610, n27014);
  and g43620 (n27017, n_19610, n27016);
  not g43621 (n_19611, n27017);
  and g43622 (n27018, pi0787, n_19611);
  and g43623 (n27019, n_11819, n26886);
  and g43624 (n27020, pi0644, n26878);
  not g43625 (n_19612, n27019);
  and g43626 (n27021, pi0790, n_19612);
  not g43627 (n_19613, n27020);
  and g43628 (n27022, n_19613, n27021);
  not g43629 (n_19614, n27012);
  not g43630 (n_19615, n27018);
  and g43631 (n27023, n_19614, n_19615);
  not g43632 (n_19616, n27022);
  and g43633 (n27024, n_19616, n27023);
  not g43634 (n_19617, n26889);
  not g43635 (n_19618, n27024);
  and g43636 (n27025, n_19617, n_19618);
  not g43637 (n_19619, n27025);
  and g43638 (n27026, n_4226, n_19619);
  not g43639 (n_19620, n26741);
  and g43640 (n27027, n_12415, n_19620);
  not g43641 (n_19621, n27026);
  and g43642 (n27028, n_19621, n27027);
  not g43643 (n_19622, n26740);
  not g43644 (n_19623, n27028);
  and g43645 (po0338, n_19622, n_19623);
  and g43646 (n27030, n_7715, n_12418);
  and g43647 (n27031, n_15580, n16645);
  not g43648 (n_19624, n27030);
  not g43649 (n_19625, n27031);
  and g43650 (n27032, n_19624, n_19625);
  not g43651 (n_19626, n27032);
  and g43652 (n27033, n_11749, n_19626);
  and g43653 (n27034, n_11753, n27031);
  not g43654 (n_19627, n27034);
  and g43655 (n27035, n_19626, n_19627);
  not g43656 (n_19628, n27035);
  and g43657 (n27036, pi1153, n_19628);
  and g43658 (n27037, n_11757, n_19624);
  and g43659 (n27038, n_19627, n27037);
  not g43660 (n_19629, n27038);
  and g43661 (n27039, pi0778, n_19629);
  not g43662 (n_19630, n27036);
  and g43663 (n27040, n_19630, n27039);
  not g43664 (n_19631, n27033);
  not g43665 (n_19632, n27040);
  and g43666 (n27041, n_19631, n_19632);
  not g43667 (n_19633, n27041);
  and g43668 (n27042, n_12429, n_19633);
  and g43669 (n27043, n_12430, n27042);
  and g43670 (n27044, n_12431, n27043);
  and g43671 (n27045, n_12432, n27044);
  and g43672 (n27046, n_12436, n27045);
  and g43673 (n27047, n_11806, n27046);
  and g43674 (n27048, pi0647, n27030);
  not g43675 (n_19634, n27048);
  and g43676 (n27049, n_11810, n_19634);
  not g43677 (n_19635, n27047);
  and g43678 (n27050, n_19635, n27049);
  and g43679 (n27051, pi0630, n27050);
  and g43680 (n27052, n_15578, n17244);
  not g43681 (n_19636, n27052);
  and g43682 (n27053, n_19624, n_19636);
  not g43683 (n_19637, n27053);
  and g43684 (n27054, n_12448, n_19637);
  not g43685 (n_19638, n27054);
  and g43686 (n27055, n_11964, n_19638);
  and g43687 (n27056, n17296, n27052);
  not g43688 (n_19639, n27056);
  and g43689 (n27057, n27054, n_19639);
  not g43690 (n_19640, n27057);
  and g43691 (n27058, pi1155, n_19640);
  and g43692 (n27059, n_11768, n_19624);
  and g43693 (n27060, n_19639, n27059);
  not g43694 (n_19641, n27058);
  not g43695 (n_19642, n27060);
  and g43696 (n27061, n_19641, n_19642);
  not g43697 (n_19643, n27061);
  and g43698 (n27062, pi0785, n_19643);
  not g43699 (n_19644, n27055);
  not g43700 (n_19645, n27062);
  and g43701 (n27063, n_19644, n_19645);
  not g43702 (n_19646, n27063);
  and g43703 (n27064, n_11981, n_19646);
  and g43704 (n27065, n_12461, n27063);
  not g43705 (n_19647, n27065);
  and g43706 (n27066, pi1154, n_19647);
  and g43707 (n27067, n_12463, n27063);
  not g43708 (n_19648, n27067);
  and g43709 (n27068, n_11413, n_19648);
  not g43710 (n_19649, n27066);
  not g43711 (n_19650, n27068);
  and g43712 (n27069, n_19649, n_19650);
  not g43713 (n_19651, n27069);
  and g43714 (n27070, pi0781, n_19651);
  not g43715 (n_19652, n27064);
  not g43716 (n_19653, n27070);
  and g43717 (n27071, n_19652, n_19653);
  not g43718 (n_19654, n27071);
  and g43719 (n27072, n_12315, n_19654);
  and g43720 (n27073, n_16503, n27071);
  not g43721 (n_19655, n27073);
  and g43722 (n27074, pi1159, n_19655);
  and g43723 (n27075, n_16505, n27071);
  not g43724 (n_19656, n27075);
  and g43725 (n27076, n_11405, n_19656);
  not g43726 (n_19657, n27074);
  not g43727 (n_19658, n27076);
  and g43728 (n27077, n_19657, n_19658);
  not g43729 (n_19659, n27077);
  and g43730 (n27078, pi0789, n_19659);
  not g43731 (n_19660, n27072);
  not g43732 (n_19661, n27078);
  and g43733 (n27079, n_19660, n_19661);
  and g43734 (n27080, n_12524, n27079);
  and g43735 (n27081, n17969, n27030);
  not g43736 (n_19662, n27080);
  not g43737 (n_19663, n27081);
  and g43738 (n27082, n_19662, n_19663);
  not g43739 (n_19664, n27082);
  and g43740 (n27083, n_12368, n_19664);
  and g43741 (n27084, n17779, n27030);
  not g43742 (n_19665, n27083);
  not g43743 (n_19666, n27084);
  and g43744 (n27085, n_19665, n_19666);
  and g43745 (n27086, n_14548, n27085);
  not g43746 (n_19667, n27046);
  and g43747 (n27087, pi0647, n_19667);
  and g43748 (n27088, n_11806, n_19624);
  not g43749 (n_19668, n27087);
  not g43750 (n_19669, n27088);
  and g43751 (n27089, n_19668, n_19669);
  not g43752 (n_19670, n27089);
  and g43753 (n27090, n17801, n_19670);
  not g43754 (n_19671, n27051);
  not g43755 (n_19672, n27090);
  and g43756 (n27091, n_19671, n_19672);
  not g43757 (n_19673, n27086);
  and g43758 (n27092, n_19673, n27091);
  not g43759 (n_19674, n27092);
  and g43760 (n27093, pi0787, n_19674);
  and g43761 (n27094, n17871, n27044);
  not g43762 (n_19675, n27079);
  and g43763 (n27095, n_12320, n_19675);
  and g43764 (n27096, pi0626, n_19624);
  not g43765 (n_19676, n27096);
  and g43766 (n27097, n16629, n_19676);
  not g43767 (n_19677, n27095);
  and g43768 (n27098, n_19677, n27097);
  and g43769 (n27099, pi0626, n_19675);
  and g43770 (n27100, n_12320, n_19624);
  not g43771 (n_19678, n27100);
  and g43772 (n27101, n16628, n_19678);
  not g43773 (n_19679, n27099);
  and g43774 (n27102, n_19679, n27101);
  not g43775 (n_19680, n27094);
  not g43776 (n_19681, n27098);
  and g43777 (n27103, n_19680, n_19681);
  not g43778 (n_19682, n27102);
  and g43779 (n27104, n_19682, n27103);
  not g43780 (n_19683, n27104);
  and g43781 (n27105, pi0788, n_19683);
  and g43782 (n27106, pi0618, n27042);
  and g43783 (n27107, n_11866, n_19626);
  and g43784 (n27108, pi0625, n27107);
  not g43785 (n_19684, n27107);
  and g43786 (n27109, n27053, n_19684);
  not g43787 (n_19685, n27108);
  not g43788 (n_19686, n27109);
  and g43789 (n27110, n_19685, n_19686);
  not g43790 (n_19687, n27110);
  and g43791 (n27111, n27037, n_19687);
  and g43792 (n27112, n_11823, n_19630);
  not g43793 (n_19688, n27111);
  and g43794 (n27113, n_19688, n27112);
  and g43795 (n27114, pi1153, n27053);
  and g43796 (n27115, n_19685, n27114);
  and g43797 (n27116, pi0608, n_19629);
  not g43798 (n_19689, n27115);
  and g43799 (n27117, n_19689, n27116);
  not g43800 (n_19690, n27113);
  not g43801 (n_19691, n27117);
  and g43802 (n27118, n_19690, n_19691);
  not g43803 (n_19692, n27118);
  and g43804 (n27119, pi0778, n_19692);
  and g43805 (n27120, n_11749, n_19686);
  not g43806 (n_19693, n27119);
  not g43807 (n_19694, n27120);
  and g43808 (n27121, n_19693, n_19694);
  not g43809 (n_19695, n27121);
  and g43810 (n27122, n_11971, n_19695);
  and g43811 (n27123, pi0609, n_19633);
  not g43812 (n_19696, n27123);
  and g43813 (n27124, n_11768, n_19696);
  not g43814 (n_19697, n27122);
  and g43815 (n27125, n_19697, n27124);
  and g43816 (n27126, n_11767, n_19641);
  not g43817 (n_19698, n27125);
  and g43818 (n27127, n_19698, n27126);
  and g43819 (n27128, pi0609, n_19695);
  and g43820 (n27129, n_11971, n_19633);
  not g43821 (n_19699, n27129);
  and g43822 (n27130, pi1155, n_19699);
  not g43823 (n_19700, n27128);
  and g43824 (n27131, n_19700, n27130);
  and g43825 (n27132, pi0660, n_19642);
  not g43826 (n_19701, n27131);
  and g43827 (n27133, n_19701, n27132);
  not g43828 (n_19702, n27127);
  not g43829 (n_19703, n27133);
  and g43830 (n27134, n_19702, n_19703);
  not g43831 (n_19704, n27134);
  and g43832 (n27135, pi0785, n_19704);
  and g43833 (n27136, n_11964, n_19695);
  not g43834 (n_19705, n27135);
  not g43835 (n_19706, n27136);
  and g43836 (n27137, n_19705, n_19706);
  not g43837 (n_19707, n27137);
  and g43838 (n27138, n_11984, n_19707);
  not g43839 (n_19708, n27106);
  and g43840 (n27139, n_11413, n_19708);
  not g43841 (n_19709, n27138);
  and g43842 (n27140, n_19709, n27139);
  and g43843 (n27141, n_11412, n_19649);
  not g43844 (n_19710, n27140);
  and g43845 (n27142, n_19710, n27141);
  and g43846 (n27143, n_11984, n27042);
  and g43847 (n27144, pi0618, n_19707);
  not g43848 (n_19711, n27143);
  and g43849 (n27145, pi1154, n_19711);
  not g43850 (n_19712, n27144);
  and g43851 (n27146, n_19712, n27145);
  and g43852 (n27147, pi0627, n_19650);
  not g43853 (n_19713, n27146);
  and g43854 (n27148, n_19713, n27147);
  not g43855 (n_19714, n27142);
  not g43856 (n_19715, n27148);
  and g43857 (n27149, n_19714, n_19715);
  not g43858 (n_19716, n27149);
  and g43859 (n27150, pi0781, n_19716);
  and g43860 (n27151, n_11981, n_19707);
  not g43861 (n_19717, n27150);
  not g43862 (n_19718, n27151);
  and g43863 (n27152, n_19717, n_19718);
  and g43864 (n27153, n_12315, n27152);
  not g43865 (n_19719, n27152);
  and g43866 (n27154, n_11821, n_19719);
  and g43867 (n27155, pi0619, n27043);
  not g43868 (n_19720, n27155);
  and g43869 (n27156, n_11405, n_19720);
  not g43870 (n_19721, n27154);
  and g43871 (n27157, n_19721, n27156);
  and g43872 (n27158, n_11403, n_19657);
  not g43873 (n_19722, n27157);
  and g43874 (n27159, n_19722, n27158);
  and g43875 (n27160, pi0619, n_19719);
  and g43876 (n27161, n_11821, n27043);
  not g43877 (n_19723, n27161);
  and g43878 (n27162, pi1159, n_19723);
  not g43879 (n_19724, n27160);
  and g43880 (n27163, n_19724, n27162);
  and g43881 (n27164, pi0648, n_19658);
  not g43882 (n_19725, n27163);
  and g43883 (n27165, n_19725, n27164);
  not g43884 (n_19726, n27159);
  and g43885 (n27166, pi0789, n_19726);
  not g43886 (n_19727, n27165);
  and g43887 (n27167, n_19727, n27166);
  not g43888 (n_19728, n27153);
  and g43889 (n27168, n17970, n_19728);
  not g43890 (n_19729, n27167);
  and g43891 (n27169, n_19729, n27168);
  not g43892 (n_19730, n27105);
  not g43893 (n_19731, n27169);
  and g43894 (n27170, n_19730, n_19731);
  not g43895 (n_19732, n27170);
  and g43896 (n27171, n_14638, n_19732);
  and g43897 (n27172, n17854, n_19664);
  and g43898 (n27173, n20851, n27045);
  not g43899 (n_19733, n27172);
  not g43900 (n_19734, n27173);
  and g43901 (n27174, n_19733, n_19734);
  not g43902 (n_19735, n27174);
  and g43903 (n27175, n_12354, n_19735);
  and g43904 (n27176, n20855, n27045);
  and g43905 (n27177, n17853, n_19664);
  not g43906 (n_19736, n27176);
  not g43907 (n_19737, n27177);
  and g43908 (n27178, n_19736, n_19737);
  not g43909 (n_19738, n27178);
  and g43910 (n27179, pi0629, n_19738);
  not g43911 (n_19739, n27175);
  not g43912 (n_19740, n27179);
  and g43913 (n27180, n_19739, n_19740);
  not g43914 (n_19741, n27180);
  and g43915 (n27181, pi0792, n_19741);
  not g43916 (n_19742, n27181);
  and g43917 (n27182, n_14387, n_19742);
  not g43918 (n_19743, n27171);
  and g43919 (n27183, n_19743, n27182);
  not g43920 (n_19744, n27093);
  not g43921 (n_19745, n27183);
  and g43922 (n27184, n_19744, n_19745);
  and g43923 (n27185, n_12411, n27184);
  and g43924 (n27186, n_11803, n_19667);
  and g43925 (n27187, pi1157, n_19670);
  not g43926 (n_19746, n27050);
  not g43927 (n_19747, n27187);
  and g43928 (n27188, n_19746, n_19747);
  not g43929 (n_19748, n27188);
  and g43930 (n27189, pi0787, n_19748);
  not g43931 (n_19749, n27186);
  not g43932 (n_19750, n27189);
  and g43933 (n27190, n_19749, n_19750);
  and g43934 (n27191, n_11819, n27190);
  and g43935 (n27192, pi0644, n27184);
  not g43936 (n_19751, n27191);
  and g43937 (n27193, pi0715, n_19751);
  not g43938 (n_19752, n27192);
  and g43939 (n27194, n_19752, n27193);
  not g43940 (n_19753, n27085);
  and g43941 (n27195, n_12392, n_19753);
  and g43942 (n27196, n17804, n27030);
  not g43943 (n_19754, n27195);
  not g43944 (n_19755, n27196);
  and g43945 (n27197, n_19754, n_19755);
  not g43946 (n_19756, n27197);
  and g43947 (n27198, pi0644, n_19756);
  and g43948 (n27199, n_11819, n27030);
  not g43949 (n_19757, n27199);
  and g43950 (n27200, n_12395, n_19757);
  not g43951 (n_19758, n27198);
  and g43952 (n27201, n_19758, n27200);
  not g43953 (n_19759, n27201);
  and g43954 (n27202, pi1160, n_19759);
  not g43955 (n_19760, n27194);
  and g43956 (n27203, n_19760, n27202);
  and g43957 (n27204, n_11819, n_19756);
  and g43958 (n27205, pi0644, n27030);
  not g43959 (n_19761, n27205);
  and g43960 (n27206, pi0715, n_19761);
  not g43961 (n_19762, n27204);
  and g43962 (n27207, n_19762, n27206);
  and g43963 (n27208, pi0644, n27190);
  and g43964 (n27209, n_11819, n27184);
  not g43965 (n_19763, n27208);
  and g43966 (n27210, n_12395, n_19763);
  not g43967 (n_19764, n27209);
  and g43968 (n27211, n_19764, n27210);
  not g43969 (n_19765, n27207);
  and g43970 (n27212, n_12405, n_19765);
  not g43971 (n_19766, n27211);
  and g43972 (n27213, n_19766, n27212);
  not g43973 (n_19767, n27203);
  not g43974 (n_19768, n27213);
  and g43975 (n27214, n_19767, n_19768);
  not g43976 (n_19769, n27214);
  and g43977 (n27215, pi0790, n_19769);
  not g43978 (n_19770, n27185);
  and g43979 (n27216, pi0832, n_19770);
  not g43980 (n_19771, n27215);
  and g43981 (n27217, n_19771, n27216);
  and g43982 (n27218, n_7715, po1038);
  and g43983 (n27219, n_7715, n_11751);
  not g43984 (n_19772, n27219);
  and g43985 (n27220, n16635, n_19772);
  and g43986 (n27221, n_15580, n2571);
  not g43987 (n_19773, n27221);
  and g43988 (n27222, n27219, n_19773);
  and g43989 (n27223, n_7715, n_11418);
  not g43990 (n_19774, n27223);
  and g43991 (n27224, n16647, n_19774);
  and g43992 (n27225, pi0182, n_12608);
  not g43993 (n_19775, n27225);
  and g43994 (n27226, n_161, n_19775);
  not g43995 (n_19776, n27226);
  and g43996 (n27227, n2571, n_19776);
  and g43997 (n27228, n_7715, n18072);
  not g43998 (n_19777, n27227);
  not g43999 (n_19778, n27228);
  and g44000 (n27229, n_19777, n_19778);
  not g44001 (n_19779, n27224);
  and g44002 (n27230, n_15580, n_19779);
  not g44003 (n_19780, n27229);
  and g44004 (n27231, n_19780, n27230);
  not g44005 (n_19781, n27222);
  not g44006 (n_19782, n27231);
  and g44007 (n27232, n_19781, n_19782);
  and g44008 (n27233, n_11749, n27232);
  and g44009 (n27234, n_11753, n27219);
  not g44010 (n_19783, n27232);
  and g44011 (n27235, pi0625, n_19783);
  not g44012 (n_19784, n27234);
  and g44013 (n27236, pi1153, n_19784);
  not g44014 (n_19785, n27235);
  and g44015 (n27237, n_19785, n27236);
  and g44016 (n27238, pi0625, n27219);
  and g44017 (n27239, n_11753, n_19783);
  not g44018 (n_19786, n27238);
  and g44019 (n27240, n_11757, n_19786);
  not g44020 (n_19787, n27239);
  and g44021 (n27241, n_19787, n27240);
  not g44022 (n_19788, n27237);
  not g44023 (n_19789, n27241);
  and g44024 (n27242, n_19788, n_19789);
  not g44025 (n_19790, n27242);
  and g44026 (n27243, pi0778, n_19790);
  not g44027 (n_19791, n27233);
  not g44028 (n_19792, n27243);
  and g44029 (n27244, n_19791, n_19792);
  not g44030 (n_19793, n27244);
  and g44031 (n27245, n_11773, n_19793);
  and g44032 (n27246, n17075, n_19772);
  not g44033 (n_19794, n27245);
  not g44034 (n_19795, n27246);
  and g44035 (n27247, n_19794, n_19795);
  and g44036 (n27248, n_11777, n27247);
  and g44037 (n27249, n16639, n27219);
  not g44038 (n_19796, n27248);
  not g44039 (n_19797, n27249);
  and g44040 (n27250, n_19796, n_19797);
  and g44041 (n27251, n_11780, n27250);
  not g44042 (n_19798, n27220);
  not g44043 (n_19799, n27251);
  and g44044 (n27252, n_19798, n_19799);
  and g44045 (n27253, n_11783, n27252);
  and g44046 (n27254, n16631, n27219);
  not g44047 (n_19800, n27253);
  not g44048 (n_19801, n27254);
  and g44049 (n27255, n_19800, n_19801);
  and g44050 (n27256, n_11787, n27255);
  not g44051 (n_19802, n27255);
  and g44052 (n27257, pi0628, n_19802);
  and g44053 (n27258, n_11789, n27219);
  not g44054 (n_19803, n27258);
  and g44055 (n27259, pi1156, n_19803);
  not g44056 (n_19804, n27257);
  and g44057 (n27260, n_19804, n27259);
  and g44058 (n27261, pi0628, n27219);
  and g44059 (n27262, n_11789, n_19802);
  not g44060 (n_19805, n27261);
  and g44061 (n27263, n_11794, n_19805);
  not g44062 (n_19806, n27262);
  and g44063 (n27264, n_19806, n27263);
  not g44064 (n_19807, n27260);
  not g44065 (n_19808, n27264);
  and g44066 (n27265, n_19807, n_19808);
  not g44067 (n_19809, n27265);
  and g44068 (n27266, pi0792, n_19809);
  not g44069 (n_19810, n27256);
  not g44070 (n_19811, n27266);
  and g44071 (n27267, n_19810, n_19811);
  not g44072 (n_19812, n27267);
  and g44073 (n27268, n_11806, n_19812);
  and g44074 (n27269, pi0647, n_19772);
  not g44075 (n_19813, n27268);
  not g44076 (n_19814, n27269);
  and g44077 (n27270, n_19813, n_19814);
  and g44078 (n27271, n_11810, n27270);
  and g44079 (n27272, pi0647, n_19812);
  and g44080 (n27273, n_11806, n_19772);
  not g44081 (n_19815, n27272);
  not g44082 (n_19816, n27273);
  and g44083 (n27274, n_19815, n_19816);
  and g44084 (n27275, pi1157, n27274);
  not g44085 (n_19817, n27271);
  not g44086 (n_19818, n27275);
  and g44087 (n27276, n_19817, n_19818);
  not g44088 (n_19819, n27276);
  and g44089 (n27277, pi0787, n_19819);
  and g44090 (n27278, n_11803, n27267);
  not g44091 (n_19820, n27277);
  not g44092 (n_19821, n27278);
  and g44093 (n27279, n_19820, n_19821);
  not g44094 (n_19822, n27279);
  and g44095 (n27280, n_11819, n_19822);
  not g44096 (n_19823, n27280);
  and g44097 (n27281, pi0715, n_19823);
  and g44098 (n27282, pi0182, n_11417);
  and g44099 (n27283, n_15578, n17280);
  not g44100 (n_19824, n27283);
  and g44101 (n27284, n_19774, n_19824);
  not g44102 (n_19825, n27284);
  and g44103 (n27285, pi0038, n_19825);
  and g44104 (n27286, n_7715, n17221);
  and g44105 (n27287, pi0182, n_14476);
  not g44106 (n_19826, n27287);
  and g44107 (n27288, n_15578, n_19826);
  not g44108 (n_19827, n27286);
  and g44109 (n27289, n_19827, n27288);
  and g44110 (n27290, n_7715, pi0756);
  and g44111 (n27291, n_11739, n27290);
  not g44112 (n_19828, n27289);
  not g44113 (n_19829, n27291);
  and g44114 (n27292, n_19828, n_19829);
  not g44115 (n_19830, n27292);
  and g44116 (n27293, n_161, n_19830);
  not g44117 (n_19831, n27285);
  not g44118 (n_19832, n27293);
  and g44119 (n27294, n_19831, n_19832);
  and g44120 (n27295, n2571, n27294);
  not g44121 (n_19833, n27282);
  not g44122 (n_19834, n27295);
  and g44123 (n27296, n_19833, n_19834);
  not g44124 (n_19835, n27296);
  and g44125 (n27297, n_11960, n_19835);
  and g44126 (n27298, n17117, n_19772);
  not g44127 (n_19836, n27297);
  not g44128 (n_19837, n27298);
  and g44129 (n27299, n_19836, n_19837);
  not g44130 (n_19838, n27299);
  and g44131 (n27300, n_11964, n_19838);
  and g44132 (n27301, n_11967, n_19772);
  and g44133 (n27302, pi0609, n27297);
  not g44134 (n_19839, n27301);
  not g44135 (n_19840, n27302);
  and g44136 (n27303, n_19839, n_19840);
  not g44137 (n_19841, n27303);
  and g44138 (n27304, pi1155, n_19841);
  and g44139 (n27305, n_11972, n_19772);
  and g44140 (n27306, n_11971, n27297);
  not g44141 (n_19842, n27305);
  not g44142 (n_19843, n27306);
  and g44143 (n27307, n_19842, n_19843);
  not g44144 (n_19844, n27307);
  and g44145 (n27308, n_11768, n_19844);
  not g44146 (n_19845, n27304);
  not g44147 (n_19846, n27308);
  and g44148 (n27309, n_19845, n_19846);
  not g44149 (n_19847, n27309);
  and g44150 (n27310, pi0785, n_19847);
  not g44151 (n_19848, n27300);
  not g44152 (n_19849, n27310);
  and g44153 (n27311, n_19848, n_19849);
  not g44154 (n_19850, n27311);
  and g44155 (n27312, n_11981, n_19850);
  and g44156 (n27313, n_11984, n27219);
  and g44157 (n27314, pi0618, n27311);
  not g44158 (n_19851, n27313);
  and g44159 (n27315, pi1154, n_19851);
  not g44160 (n_19852, n27314);
  and g44161 (n27316, n_19852, n27315);
  and g44162 (n27317, n_11984, n27311);
  and g44163 (n27318, pi0618, n27219);
  not g44164 (n_19853, n27318);
  and g44165 (n27319, n_11413, n_19853);
  not g44166 (n_19854, n27317);
  and g44167 (n27320, n_19854, n27319);
  not g44168 (n_19855, n27316);
  not g44169 (n_19856, n27320);
  and g44170 (n27321, n_19855, n_19856);
  not g44171 (n_19857, n27321);
  and g44172 (n27322, pi0781, n_19857);
  not g44173 (n_19858, n27312);
  not g44174 (n_19859, n27322);
  and g44175 (n27323, n_19858, n_19859);
  not g44176 (n_19860, n27323);
  and g44177 (n27324, n_12315, n_19860);
  and g44178 (n27325, n_11821, n27219);
  and g44179 (n27326, pi0619, n27323);
  not g44180 (n_19861, n27325);
  and g44181 (n27327, pi1159, n_19861);
  not g44182 (n_19862, n27326);
  and g44183 (n27328, n_19862, n27327);
  and g44184 (n27329, n_11821, n27323);
  and g44185 (n27330, pi0619, n27219);
  not g44186 (n_19863, n27330);
  and g44187 (n27331, n_11405, n_19863);
  not g44188 (n_19864, n27329);
  and g44189 (n27332, n_19864, n27331);
  not g44190 (n_19865, n27328);
  not g44191 (n_19866, n27332);
  and g44192 (n27333, n_19865, n_19866);
  not g44193 (n_19867, n27333);
  and g44194 (n27334, pi0789, n_19867);
  not g44195 (n_19868, n27324);
  not g44196 (n_19869, n27334);
  and g44197 (n27335, n_19868, n_19869);
  and g44198 (n27336, n_12524, n27335);
  and g44199 (n27337, n17969, n27219);
  not g44200 (n_19870, n27336);
  not g44201 (n_19871, n27337);
  and g44202 (n27338, n_19870, n_19871);
  not g44203 (n_19872, n27338);
  and g44204 (n27339, n_12368, n_19872);
  and g44205 (n27340, n17779, n27219);
  not g44206 (n_19873, n27339);
  not g44207 (n_19874, n27340);
  and g44208 (n27341, n_19873, n_19874);
  not g44209 (n_19875, n27341);
  and g44210 (n27342, n_12392, n_19875);
  and g44211 (n27343, n17804, n27219);
  not g44212 (n_19876, n27342);
  not g44213 (n_19877, n27343);
  and g44214 (n27344, n_19876, n_19877);
  not g44215 (n_19878, n27344);
  and g44216 (n27345, pi0644, n_19878);
  and g44217 (n27346, n_11819, n27219);
  not g44218 (n_19879, n27346);
  and g44219 (n27347, n_12395, n_19879);
  not g44220 (n_19880, n27345);
  and g44221 (n27348, n_19880, n27347);
  not g44222 (n_19881, n27348);
  and g44223 (n27349, pi1160, n_19881);
  not g44224 (n_19882, n27281);
  and g44225 (n27350, n_19882, n27349);
  and g44226 (n27351, pi0644, n_19822);
  not g44227 (n_19883, n27351);
  and g44228 (n27352, n_12395, n_19883);
  and g44229 (n27353, n_11819, n_19878);
  and g44230 (n27354, pi0644, n27219);
  not g44231 (n_19884, n27354);
  and g44232 (n27355, pi0715, n_19884);
  not g44233 (n_19885, n27353);
  and g44234 (n27356, n_19885, n27355);
  not g44235 (n_19886, n27356);
  and g44236 (n27357, n_12405, n_19886);
  not g44237 (n_19887, n27352);
  and g44238 (n27358, n_19887, n27357);
  not g44239 (n_19888, n27350);
  not g44240 (n_19889, n27358);
  and g44241 (n27359, n_19888, n_19889);
  not g44242 (n_19890, n27359);
  and g44243 (n27360, pi0790, n_19890);
  and g44244 (n27361, n_12354, n27260);
  and g44245 (n27362, n_14557, n27338);
  and g44246 (n27363, pi0629, n27264);
  not g44247 (n_19891, n27361);
  not g44248 (n_19892, n27363);
  and g44249 (n27364, n_19891, n_19892);
  not g44250 (n_19893, n27362);
  and g44251 (n27365, n_19893, n27364);
  not g44252 (n_19894, n27365);
  and g44253 (n27366, pi0792, n_19894);
  and g44254 (n27367, pi0609, n27244);
  and g44255 (n27368, pi0182, n_12240);
  and g44256 (n27369, n_7715, n_12230);
  not g44257 (n_19895, n27368);
  and g44258 (n27370, pi0756, n_19895);
  not g44259 (n_19896, n27369);
  and g44260 (n27371, n_19896, n27370);
  and g44261 (n27372, n_7715, n17629);
  and g44262 (n27373, pi0182, n17631);
  not g44263 (n_19897, n27373);
  and g44264 (n27374, n_15578, n_19897);
  not g44265 (n_19898, n27372);
  and g44266 (n27375, n_19898, n27374);
  not g44267 (n_19899, n27371);
  not g44268 (n_19900, n27375);
  and g44269 (n27376, n_19899, n_19900);
  not g44270 (n_19901, n27376);
  and g44271 (n27377, n_162, n_19901);
  and g44272 (n27378, pi0182, n17605);
  and g44273 (n27379, n_7715, n_12180);
  not g44274 (n_19902, n27379);
  and g44275 (n27380, n_15578, n_19902);
  not g44276 (n_19903, n27378);
  and g44277 (n27381, n_19903, n27380);
  and g44278 (n27382, n_7715, n17404);
  and g44279 (n27383, pi0182, n17485);
  not g44280 (n_19904, n27383);
  and g44281 (n27384, pi0756, n_19904);
  not g44282 (n_19905, n27382);
  and g44283 (n27385, n_19905, n27384);
  not g44284 (n_19906, n27381);
  and g44285 (n27386, pi0039, n_19906);
  not g44286 (n_19907, n27385);
  and g44287 (n27387, n_19907, n27386);
  not g44288 (n_19908, n27377);
  and g44289 (n27388, n_161, n_19908);
  not g44290 (n_19909, n27387);
  and g44291 (n27389, n_19909, n27388);
  and g44292 (n27390, n_15578, n_12250);
  not g44293 (n_19910, n27390);
  and g44294 (n27391, n19471, n_19910);
  not g44295 (n_19911, n27391);
  and g44296 (n27392, n_7715, n_19911);
  and g44297 (n27393, n_12120, n_19636);
  not g44298 (n_19912, n27393);
  and g44299 (n27394, pi0182, n_19912);
  and g44300 (n27395, n6284, n27394);
  not g44301 (n_19913, n27395);
  and g44302 (n27396, pi0038, n_19913);
  not g44303 (n_19914, n27392);
  and g44304 (n27397, n_19914, n27396);
  not g44305 (n_19915, n27397);
  and g44306 (n27398, n_15580, n_19915);
  not g44307 (n_19916, n27389);
  and g44308 (n27399, n_19916, n27398);
  not g44309 (n_19917, n27294);
  and g44310 (n27400, pi0734, n_19917);
  not g44311 (n_19918, n27399);
  and g44312 (n27401, n2571, n_19918);
  not g44313 (n_19919, n27400);
  and g44314 (n27402, n_19919, n27401);
  not g44315 (n_19920, n27402);
  and g44316 (n27403, n_19833, n_19920);
  and g44317 (n27404, n_11753, n27403);
  and g44318 (n27405, pi0625, n27296);
  not g44319 (n_19921, n27405);
  and g44320 (n27406, n_11757, n_19921);
  not g44321 (n_19922, n27404);
  and g44322 (n27407, n_19922, n27406);
  and g44323 (n27408, n_11823, n_19788);
  not g44324 (n_19923, n27407);
  and g44325 (n27409, n_19923, n27408);
  and g44326 (n27410, n_11753, n27296);
  and g44327 (n27411, pi0625, n27403);
  not g44328 (n_19924, n27410);
  and g44329 (n27412, pi1153, n_19924);
  not g44330 (n_19925, n27411);
  and g44331 (n27413, n_19925, n27412);
  and g44332 (n27414, pi0608, n_19789);
  not g44333 (n_19926, n27413);
  and g44334 (n27415, n_19926, n27414);
  not g44335 (n_19927, n27409);
  not g44336 (n_19928, n27415);
  and g44337 (n27416, n_19927, n_19928);
  not g44338 (n_19929, n27416);
  and g44339 (n27417, pi0778, n_19929);
  and g44340 (n27418, n_11749, n27403);
  not g44341 (n_19930, n27417);
  not g44342 (n_19931, n27418);
  and g44343 (n27419, n_19930, n_19931);
  not g44344 (n_19932, n27419);
  and g44345 (n27420, n_11971, n_19932);
  not g44346 (n_19933, n27367);
  and g44347 (n27421, n_11768, n_19933);
  not g44348 (n_19934, n27420);
  and g44349 (n27422, n_19934, n27421);
  and g44350 (n27423, n_11767, n_19845);
  not g44351 (n_19935, n27422);
  and g44352 (n27424, n_19935, n27423);
  and g44353 (n27425, n_11971, n27244);
  and g44354 (n27426, pi0609, n_19932);
  not g44355 (n_19936, n27425);
  and g44356 (n27427, pi1155, n_19936);
  not g44357 (n_19937, n27426);
  and g44358 (n27428, n_19937, n27427);
  and g44359 (n27429, pi0660, n_19846);
  not g44360 (n_19938, n27428);
  and g44361 (n27430, n_19938, n27429);
  not g44362 (n_19939, n27424);
  not g44363 (n_19940, n27430);
  and g44364 (n27431, n_19939, n_19940);
  not g44365 (n_19941, n27431);
  and g44366 (n27432, pi0785, n_19941);
  and g44367 (n27433, n_11964, n_19932);
  not g44368 (n_19942, n27432);
  not g44369 (n_19943, n27433);
  and g44370 (n27434, n_19942, n_19943);
  not g44371 (n_19944, n27434);
  and g44372 (n27435, n_11984, n_19944);
  and g44373 (n27436, pi0618, n27247);
  not g44374 (n_19945, n27436);
  and g44375 (n27437, n_11413, n_19945);
  not g44376 (n_19946, n27435);
  and g44377 (n27438, n_19946, n27437);
  and g44378 (n27439, n_11412, n_19855);
  not g44379 (n_19947, n27438);
  and g44380 (n27440, n_19947, n27439);
  and g44381 (n27441, n_11984, n27247);
  and g44382 (n27442, pi0618, n_19944);
  not g44383 (n_19948, n27441);
  and g44384 (n27443, pi1154, n_19948);
  not g44385 (n_19949, n27442);
  and g44386 (n27444, n_19949, n27443);
  and g44387 (n27445, pi0627, n_19856);
  not g44388 (n_19950, n27444);
  and g44389 (n27446, n_19950, n27445);
  not g44390 (n_19951, n27440);
  not g44391 (n_19952, n27446);
  and g44392 (n27447, n_19951, n_19952);
  not g44393 (n_19953, n27447);
  and g44394 (n27448, pi0781, n_19953);
  and g44395 (n27449, n_11981, n_19944);
  not g44396 (n_19954, n27448);
  not g44397 (n_19955, n27449);
  and g44398 (n27450, n_19954, n_19955);
  and g44399 (n27451, n_12315, n27450);
  not g44400 (n_19956, n27250);
  and g44401 (n27452, pi0619, n_19956);
  not g44402 (n_19957, n27450);
  and g44403 (n27453, n_11821, n_19957);
  not g44404 (n_19958, n27452);
  and g44405 (n27454, n_11405, n_19958);
  not g44406 (n_19959, n27453);
  and g44407 (n27455, n_19959, n27454);
  and g44408 (n27456, n_11403, n_19865);
  not g44409 (n_19960, n27455);
  and g44410 (n27457, n_19960, n27456);
  and g44411 (n27458, n_11821, n_19956);
  and g44412 (n27459, pi0619, n_19957);
  not g44413 (n_19961, n27458);
  and g44414 (n27460, pi1159, n_19961);
  not g44415 (n_19962, n27459);
  and g44416 (n27461, n_19962, n27460);
  and g44417 (n27462, pi0648, n_19866);
  not g44418 (n_19963, n27461);
  and g44419 (n27463, n_19963, n27462);
  not g44420 (n_19964, n27457);
  and g44421 (n27464, pi0789, n_19964);
  not g44422 (n_19965, n27463);
  and g44423 (n27465, n_19965, n27464);
  not g44424 (n_19966, n27451);
  and g44425 (n27466, n17970, n_19966);
  not g44426 (n_19967, n27465);
  and g44427 (n27467, n_19967, n27466);
  and g44428 (n27468, n17871, n27252);
  not g44429 (n_19968, n27335);
  and g44430 (n27469, n_12320, n_19968);
  and g44431 (n27470, pi0626, n_19772);
  not g44432 (n_19969, n27470);
  and g44433 (n27471, n16629, n_19969);
  not g44434 (n_19970, n27469);
  and g44435 (n27472, n_19970, n27471);
  and g44436 (n27473, pi0626, n_19968);
  and g44437 (n27474, n_12320, n_19772);
  not g44438 (n_19971, n27474);
  and g44439 (n27475, n16628, n_19971);
  not g44440 (n_19972, n27473);
  and g44441 (n27476, n_19972, n27475);
  not g44442 (n_19973, n27468);
  not g44443 (n_19974, n27472);
  and g44444 (n27477, n_19973, n_19974);
  not g44445 (n_19975, n27476);
  and g44446 (n27478, n_19975, n27477);
  not g44447 (n_19976, n27478);
  and g44448 (n27479, pi0788, n_19976);
  not g44449 (n_19977, n27479);
  and g44450 (n27480, n_14638, n_19977);
  not g44451 (n_19978, n27467);
  and g44452 (n27481, n_19978, n27480);
  not g44453 (n_19979, n27366);
  not g44454 (n_19980, n27481);
  and g44455 (n27482, n_19979, n_19980);
  not g44456 (n_19981, n27482);
  and g44457 (n27483, n_14387, n_19981);
  not g44458 (n_19982, n27270);
  and g44459 (n27484, n17802, n_19982);
  and g44460 (n27485, n_14548, n27341);
  not g44461 (n_19983, n27274);
  and g44462 (n27486, n17801, n_19983);
  not g44463 (n_19984, n27484);
  not g44464 (n_19985, n27486);
  and g44465 (n27487, n_19984, n_19985);
  not g44466 (n_19986, n27485);
  and g44467 (n27488, n_19986, n27487);
  not g44468 (n_19987, n27488);
  and g44469 (n27489, pi0787, n_19987);
  and g44470 (n27490, n_11819, n27357);
  and g44471 (n27491, pi0644, n27349);
  not g44472 (n_19988, n27490);
  and g44473 (n27492, pi0790, n_19988);
  not g44474 (n_19989, n27491);
  and g44475 (n27493, n_19989, n27492);
  not g44476 (n_19990, n27483);
  not g44477 (n_19991, n27489);
  and g44478 (n27494, n_19990, n_19991);
  not g44479 (n_19992, n27493);
  and g44480 (n27495, n_19992, n27494);
  not g44481 (n_19993, n27360);
  not g44482 (n_19994, n27495);
  and g44483 (n27496, n_19993, n_19994);
  not g44484 (n_19995, n27496);
  and g44485 (n27497, n_4226, n_19995);
  not g44486 (n_19996, n27218);
  and g44487 (n27498, n_12415, n_19996);
  not g44488 (n_19997, n27497);
  and g44489 (n27499, n_19997, n27498);
  not g44490 (n_19998, n27217);
  not g44491 (n_19999, n27499);
  and g44492 (po0339, n_19998, n_19999);
  and g44493 (n27501, n_5709, n_12418);
  and g44494 (n27502, n_15036, n16645);
  not g44495 (n_20000, n27501);
  not g44496 (n_20001, n27502);
  and g44497 (n27503, n_20000, n_20001);
  not g44498 (n_20002, n27503);
  and g44499 (n27504, n_11749, n_20002);
  and g44500 (n27505, n_11753, n27502);
  not g44501 (n_20003, n27505);
  and g44502 (n27506, n_20002, n_20003);
  not g44503 (n_20004, n27506);
  and g44504 (n27507, pi1153, n_20004);
  and g44505 (n27508, n_11757, n_20000);
  and g44506 (n27509, n_20003, n27508);
  not g44507 (n_20005, n27509);
  and g44508 (n27510, pi0778, n_20005);
  not g44509 (n_20006, n27507);
  and g44510 (n27511, n_20006, n27510);
  not g44511 (n_20007, n27504);
  not g44512 (n_20008, n27511);
  and g44513 (n27512, n_20007, n_20008);
  not g44514 (n_20009, n27512);
  and g44515 (n27513, n_12429, n_20009);
  and g44516 (n27514, n_12430, n27513);
  and g44517 (n27515, n_12431, n27514);
  and g44518 (n27516, n_12432, n27515);
  and g44519 (n27517, n_12436, n27516);
  and g44520 (n27518, n_11806, n27517);
  and g44521 (n27519, pi0647, n27501);
  not g44522 (n_20010, n27519);
  and g44523 (n27520, n_11810, n_20010);
  not g44524 (n_20011, n27518);
  and g44525 (n27521, n_20011, n27520);
  and g44526 (n27522, pi0630, n27521);
  and g44527 (n27523, n_15034, n17244);
  not g44528 (n_20012, n27523);
  and g44529 (n27524, n_20000, n_20012);
  not g44530 (n_20013, n27524);
  and g44531 (n27525, n_12448, n_20013);
  not g44532 (n_20014, n27525);
  and g44533 (n27526, n_11964, n_20014);
  and g44534 (n27527, n17296, n27523);
  not g44535 (n_20015, n27527);
  and g44536 (n27528, n27525, n_20015);
  not g44537 (n_20016, n27528);
  and g44538 (n27529, pi1155, n_20016);
  and g44539 (n27530, n_11768, n_20000);
  and g44540 (n27531, n_20015, n27530);
  not g44541 (n_20017, n27529);
  not g44542 (n_20018, n27531);
  and g44543 (n27532, n_20017, n_20018);
  not g44544 (n_20019, n27532);
  and g44545 (n27533, pi0785, n_20019);
  not g44546 (n_20020, n27526);
  not g44547 (n_20021, n27533);
  and g44548 (n27534, n_20020, n_20021);
  not g44549 (n_20022, n27534);
  and g44550 (n27535, n_11981, n_20022);
  and g44551 (n27536, n_12461, n27534);
  not g44552 (n_20023, n27536);
  and g44553 (n27537, pi1154, n_20023);
  and g44554 (n27538, n_12463, n27534);
  not g44555 (n_20024, n27538);
  and g44556 (n27539, n_11413, n_20024);
  not g44557 (n_20025, n27537);
  not g44558 (n_20026, n27539);
  and g44559 (n27540, n_20025, n_20026);
  not g44560 (n_20027, n27540);
  and g44561 (n27541, pi0781, n_20027);
  not g44562 (n_20028, n27535);
  not g44563 (n_20029, n27541);
  and g44564 (n27542, n_20028, n_20029);
  not g44565 (n_20030, n27542);
  and g44566 (n27543, n_12315, n_20030);
  and g44567 (n27544, n_16503, n27542);
  not g44568 (n_20031, n27544);
  and g44569 (n27545, pi1159, n_20031);
  and g44570 (n27546, n_16505, n27542);
  not g44571 (n_20032, n27546);
  and g44572 (n27547, n_11405, n_20032);
  not g44573 (n_20033, n27545);
  not g44574 (n_20034, n27547);
  and g44575 (n27548, n_20033, n_20034);
  not g44576 (n_20035, n27548);
  and g44577 (n27549, pi0789, n_20035);
  not g44578 (n_20036, n27543);
  not g44579 (n_20037, n27549);
  and g44580 (n27550, n_20036, n_20037);
  and g44581 (n27551, n_12524, n27550);
  and g44582 (n27552, n17969, n27501);
  not g44583 (n_20038, n27551);
  not g44584 (n_20039, n27552);
  and g44585 (n27553, n_20038, n_20039);
  not g44586 (n_20040, n27553);
  and g44587 (n27554, n_12368, n_20040);
  and g44588 (n27555, n17779, n27501);
  not g44589 (n_20041, n27554);
  not g44590 (n_20042, n27555);
  and g44591 (n27556, n_20041, n_20042);
  and g44592 (n27557, n_14548, n27556);
  not g44593 (n_20043, n27517);
  and g44594 (n27558, pi0647, n_20043);
  and g44595 (n27559, n_11806, n_20000);
  not g44596 (n_20044, n27558);
  not g44597 (n_20045, n27559);
  and g44598 (n27560, n_20044, n_20045);
  not g44599 (n_20046, n27560);
  and g44600 (n27561, n17801, n_20046);
  not g44601 (n_20047, n27522);
  not g44602 (n_20048, n27561);
  and g44603 (n27562, n_20047, n_20048);
  not g44604 (n_20049, n27557);
  and g44605 (n27563, n_20049, n27562);
  not g44606 (n_20050, n27563);
  and g44607 (n27564, pi0787, n_20050);
  and g44608 (n27565, n17871, n27515);
  not g44609 (n_20051, n27550);
  and g44610 (n27566, n_12320, n_20051);
  and g44611 (n27567, pi0626, n_20000);
  not g44612 (n_20052, n27567);
  and g44613 (n27568, n16629, n_20052);
  not g44614 (n_20053, n27566);
  and g44615 (n27569, n_20053, n27568);
  and g44616 (n27570, pi0626, n_20051);
  and g44617 (n27571, n_12320, n_20000);
  not g44618 (n_20054, n27571);
  and g44619 (n27572, n16628, n_20054);
  not g44620 (n_20055, n27570);
  and g44621 (n27573, n_20055, n27572);
  not g44622 (n_20056, n27565);
  not g44623 (n_20057, n27569);
  and g44624 (n27574, n_20056, n_20057);
  not g44625 (n_20058, n27573);
  and g44626 (n27575, n_20058, n27574);
  not g44627 (n_20059, n27575);
  and g44628 (n27576, pi0788, n_20059);
  and g44629 (n27577, pi0618, n27513);
  and g44630 (n27578, n_11866, n_20002);
  and g44631 (n27579, pi0625, n27578);
  not g44632 (n_20060, n27578);
  and g44633 (n27580, n27524, n_20060);
  not g44634 (n_20061, n27579);
  not g44635 (n_20062, n27580);
  and g44636 (n27581, n_20061, n_20062);
  not g44637 (n_20063, n27581);
  and g44638 (n27582, n27508, n_20063);
  and g44639 (n27583, n_11823, n_20006);
  not g44640 (n_20064, n27582);
  and g44641 (n27584, n_20064, n27583);
  and g44642 (n27585, pi1153, n27524);
  and g44643 (n27586, n_20061, n27585);
  and g44644 (n27587, pi0608, n_20005);
  not g44645 (n_20065, n27586);
  and g44646 (n27588, n_20065, n27587);
  not g44647 (n_20066, n27584);
  not g44648 (n_20067, n27588);
  and g44649 (n27589, n_20066, n_20067);
  not g44650 (n_20068, n27589);
  and g44651 (n27590, pi0778, n_20068);
  and g44652 (n27591, n_11749, n_20062);
  not g44653 (n_20069, n27590);
  not g44654 (n_20070, n27591);
  and g44655 (n27592, n_20069, n_20070);
  not g44656 (n_20071, n27592);
  and g44657 (n27593, n_11971, n_20071);
  and g44658 (n27594, pi0609, n_20009);
  not g44659 (n_20072, n27594);
  and g44660 (n27595, n_11768, n_20072);
  not g44661 (n_20073, n27593);
  and g44662 (n27596, n_20073, n27595);
  and g44663 (n27597, n_11767, n_20017);
  not g44664 (n_20074, n27596);
  and g44665 (n27598, n_20074, n27597);
  and g44666 (n27599, pi0609, n_20071);
  and g44667 (n27600, n_11971, n_20009);
  not g44668 (n_20075, n27600);
  and g44669 (n27601, pi1155, n_20075);
  not g44670 (n_20076, n27599);
  and g44671 (n27602, n_20076, n27601);
  and g44672 (n27603, pi0660, n_20018);
  not g44673 (n_20077, n27602);
  and g44674 (n27604, n_20077, n27603);
  not g44675 (n_20078, n27598);
  not g44676 (n_20079, n27604);
  and g44677 (n27605, n_20078, n_20079);
  not g44678 (n_20080, n27605);
  and g44679 (n27606, pi0785, n_20080);
  and g44680 (n27607, n_11964, n_20071);
  not g44681 (n_20081, n27606);
  not g44682 (n_20082, n27607);
  and g44683 (n27608, n_20081, n_20082);
  not g44684 (n_20083, n27608);
  and g44685 (n27609, n_11984, n_20083);
  not g44686 (n_20084, n27577);
  and g44687 (n27610, n_11413, n_20084);
  not g44688 (n_20085, n27609);
  and g44689 (n27611, n_20085, n27610);
  and g44690 (n27612, n_11412, n_20025);
  not g44691 (n_20086, n27611);
  and g44692 (n27613, n_20086, n27612);
  and g44693 (n27614, n_11984, n27513);
  and g44694 (n27615, pi0618, n_20083);
  not g44695 (n_20087, n27614);
  and g44696 (n27616, pi1154, n_20087);
  not g44697 (n_20088, n27615);
  and g44698 (n27617, n_20088, n27616);
  and g44699 (n27618, pi0627, n_20026);
  not g44700 (n_20089, n27617);
  and g44701 (n27619, n_20089, n27618);
  not g44702 (n_20090, n27613);
  not g44703 (n_20091, n27619);
  and g44704 (n27620, n_20090, n_20091);
  not g44705 (n_20092, n27620);
  and g44706 (n27621, pi0781, n_20092);
  and g44707 (n27622, n_11981, n_20083);
  not g44708 (n_20093, n27621);
  not g44709 (n_20094, n27622);
  and g44710 (n27623, n_20093, n_20094);
  and g44711 (n27624, n_12315, n27623);
  not g44712 (n_20095, n27623);
  and g44713 (n27625, n_11821, n_20095);
  and g44714 (n27626, pi0619, n27514);
  not g44715 (n_20096, n27626);
  and g44716 (n27627, n_11405, n_20096);
  not g44717 (n_20097, n27625);
  and g44718 (n27628, n_20097, n27627);
  and g44719 (n27629, n_11403, n_20033);
  not g44720 (n_20098, n27628);
  and g44721 (n27630, n_20098, n27629);
  and g44722 (n27631, pi0619, n_20095);
  and g44723 (n27632, n_11821, n27514);
  not g44724 (n_20099, n27632);
  and g44725 (n27633, pi1159, n_20099);
  not g44726 (n_20100, n27631);
  and g44727 (n27634, n_20100, n27633);
  and g44728 (n27635, pi0648, n_20034);
  not g44729 (n_20101, n27634);
  and g44730 (n27636, n_20101, n27635);
  not g44731 (n_20102, n27630);
  and g44732 (n27637, pi0789, n_20102);
  not g44733 (n_20103, n27636);
  and g44734 (n27638, n_20103, n27637);
  not g44735 (n_20104, n27624);
  and g44736 (n27639, n17970, n_20104);
  not g44737 (n_20105, n27638);
  and g44738 (n27640, n_20105, n27639);
  not g44739 (n_20106, n27576);
  not g44740 (n_20107, n27640);
  and g44741 (n27641, n_20106, n_20107);
  not g44742 (n_20108, n27641);
  and g44743 (n27642, n_14638, n_20108);
  and g44744 (n27643, n17854, n_20040);
  and g44745 (n27644, n20851, n27516);
  not g44746 (n_20109, n27643);
  not g44747 (n_20110, n27644);
  and g44748 (n27645, n_20109, n_20110);
  not g44749 (n_20111, n27645);
  and g44750 (n27646, n_12354, n_20111);
  and g44751 (n27647, n20855, n27516);
  and g44752 (n27648, n17853, n_20040);
  not g44753 (n_20112, n27647);
  not g44754 (n_20113, n27648);
  and g44755 (n27649, n_20112, n_20113);
  not g44756 (n_20114, n27649);
  and g44757 (n27650, pi0629, n_20114);
  not g44758 (n_20115, n27646);
  not g44759 (n_20116, n27650);
  and g44760 (n27651, n_20115, n_20116);
  not g44761 (n_20117, n27651);
  and g44762 (n27652, pi0792, n_20117);
  not g44763 (n_20118, n27652);
  and g44764 (n27653, n_14387, n_20118);
  not g44765 (n_20119, n27642);
  and g44766 (n27654, n_20119, n27653);
  not g44767 (n_20120, n27564);
  not g44768 (n_20121, n27654);
  and g44769 (n27655, n_20120, n_20121);
  and g44770 (n27656, n_12411, n27655);
  and g44771 (n27657, n_11803, n_20043);
  and g44772 (n27658, pi1157, n_20046);
  not g44773 (n_20122, n27521);
  not g44774 (n_20123, n27658);
  and g44775 (n27659, n_20122, n_20123);
  not g44776 (n_20124, n27659);
  and g44777 (n27660, pi0787, n_20124);
  not g44778 (n_20125, n27657);
  not g44779 (n_20126, n27660);
  and g44780 (n27661, n_20125, n_20126);
  and g44781 (n27662, n_11819, n27661);
  and g44782 (n27663, pi0644, n27655);
  not g44783 (n_20127, n27662);
  and g44784 (n27664, pi0715, n_20127);
  not g44785 (n_20128, n27663);
  and g44786 (n27665, n_20128, n27664);
  not g44787 (n_20129, n27556);
  and g44788 (n27666, n_12392, n_20129);
  and g44789 (n27667, n17804, n27501);
  not g44790 (n_20130, n27666);
  not g44791 (n_20131, n27667);
  and g44792 (n27668, n_20130, n_20131);
  not g44793 (n_20132, n27668);
  and g44794 (n27669, pi0644, n_20132);
  and g44795 (n27670, n_11819, n27501);
  not g44796 (n_20133, n27670);
  and g44797 (n27671, n_12395, n_20133);
  not g44798 (n_20134, n27669);
  and g44799 (n27672, n_20134, n27671);
  not g44800 (n_20135, n27672);
  and g44801 (n27673, pi1160, n_20135);
  not g44802 (n_20136, n27665);
  and g44803 (n27674, n_20136, n27673);
  and g44804 (n27675, n_11819, n_20132);
  and g44805 (n27676, pi0644, n27501);
  not g44806 (n_20137, n27676);
  and g44807 (n27677, pi0715, n_20137);
  not g44808 (n_20138, n27675);
  and g44809 (n27678, n_20138, n27677);
  and g44810 (n27679, pi0644, n27661);
  and g44811 (n27680, n_11819, n27655);
  not g44812 (n_20139, n27679);
  and g44813 (n27681, n_12395, n_20139);
  not g44814 (n_20140, n27680);
  and g44815 (n27682, n_20140, n27681);
  not g44816 (n_20141, n27678);
  and g44817 (n27683, n_12405, n_20141);
  not g44818 (n_20142, n27682);
  and g44819 (n27684, n_20142, n27683);
  not g44820 (n_20143, n27674);
  not g44821 (n_20144, n27684);
  and g44822 (n27685, n_20143, n_20144);
  not g44823 (n_20145, n27685);
  and g44824 (n27686, pi0790, n_20145);
  not g44825 (n_20146, n27656);
  and g44826 (n27687, pi0832, n_20146);
  not g44827 (n_20147, n27686);
  and g44828 (n27688, n_20147, n27687);
  and g44829 (n27689, n_5709, po1038);
  and g44830 (n27690, n_5709, n_11751);
  not g44831 (n_20148, n27690);
  and g44832 (n27691, n16635, n_20148);
  and g44833 (n27692, n_15036, n2571);
  not g44834 (n_20149, n27692);
  and g44835 (n27693, n27690, n_20149);
  and g44836 (n27694, n_5709, n_11418);
  not g44837 (n_20150, n27694);
  and g44838 (n27695, n16647, n_20150);
  and g44839 (n27696, pi0183, n_12608);
  not g44840 (n_20151, n27696);
  and g44841 (n27697, n_161, n_20151);
  not g44842 (n_20152, n27697);
  and g44843 (n27698, n2571, n_20152);
  and g44844 (n27699, n_5709, n18072);
  not g44845 (n_20153, n27698);
  not g44846 (n_20154, n27699);
  and g44847 (n27700, n_20153, n_20154);
  not g44848 (n_20155, n27695);
  and g44849 (n27701, n_15036, n_20155);
  not g44850 (n_20156, n27700);
  and g44851 (n27702, n_20156, n27701);
  not g44852 (n_20157, n27693);
  not g44853 (n_20158, n27702);
  and g44854 (n27703, n_20157, n_20158);
  and g44855 (n27704, n_11749, n27703);
  and g44856 (n27705, n_11753, n27690);
  not g44857 (n_20159, n27703);
  and g44858 (n27706, pi0625, n_20159);
  not g44859 (n_20160, n27705);
  and g44860 (n27707, pi1153, n_20160);
  not g44861 (n_20161, n27706);
  and g44862 (n27708, n_20161, n27707);
  and g44863 (n27709, pi0625, n27690);
  and g44864 (n27710, n_11753, n_20159);
  not g44865 (n_20162, n27709);
  and g44866 (n27711, n_11757, n_20162);
  not g44867 (n_20163, n27710);
  and g44868 (n27712, n_20163, n27711);
  not g44869 (n_20164, n27708);
  not g44870 (n_20165, n27712);
  and g44871 (n27713, n_20164, n_20165);
  not g44872 (n_20166, n27713);
  and g44873 (n27714, pi0778, n_20166);
  not g44874 (n_20167, n27704);
  not g44875 (n_20168, n27714);
  and g44876 (n27715, n_20167, n_20168);
  not g44877 (n_20169, n27715);
  and g44878 (n27716, n_11773, n_20169);
  and g44879 (n27717, n17075, n_20148);
  not g44880 (n_20170, n27716);
  not g44881 (n_20171, n27717);
  and g44882 (n27718, n_20170, n_20171);
  and g44883 (n27719, n_11777, n27718);
  and g44884 (n27720, n16639, n27690);
  not g44885 (n_20172, n27719);
  not g44886 (n_20173, n27720);
  and g44887 (n27721, n_20172, n_20173);
  and g44888 (n27722, n_11780, n27721);
  not g44889 (n_20174, n27691);
  not g44890 (n_20175, n27722);
  and g44891 (n27723, n_20174, n_20175);
  and g44892 (n27724, n_11783, n27723);
  and g44893 (n27725, n16631, n27690);
  not g44894 (n_20176, n27724);
  not g44895 (n_20177, n27725);
  and g44896 (n27726, n_20176, n_20177);
  and g44897 (n27727, n_11787, n27726);
  not g44898 (n_20178, n27726);
  and g44899 (n27728, pi0628, n_20178);
  and g44900 (n27729, n_11789, n27690);
  not g44901 (n_20179, n27729);
  and g44902 (n27730, pi1156, n_20179);
  not g44903 (n_20180, n27728);
  and g44904 (n27731, n_20180, n27730);
  and g44905 (n27732, pi0628, n27690);
  and g44906 (n27733, n_11789, n_20178);
  not g44907 (n_20181, n27732);
  and g44908 (n27734, n_11794, n_20181);
  not g44909 (n_20182, n27733);
  and g44910 (n27735, n_20182, n27734);
  not g44911 (n_20183, n27731);
  not g44912 (n_20184, n27735);
  and g44913 (n27736, n_20183, n_20184);
  not g44914 (n_20185, n27736);
  and g44915 (n27737, pi0792, n_20185);
  not g44916 (n_20186, n27727);
  not g44917 (n_20187, n27737);
  and g44918 (n27738, n_20186, n_20187);
  not g44919 (n_20188, n27738);
  and g44920 (n27739, n_11806, n_20188);
  and g44921 (n27740, pi0647, n_20148);
  not g44922 (n_20189, n27739);
  not g44923 (n_20190, n27740);
  and g44924 (n27741, n_20189, n_20190);
  and g44925 (n27742, n_11810, n27741);
  and g44926 (n27743, pi0647, n_20188);
  and g44927 (n27744, n_11806, n_20148);
  not g44928 (n_20191, n27743);
  not g44929 (n_20192, n27744);
  and g44930 (n27745, n_20191, n_20192);
  and g44931 (n27746, pi1157, n27745);
  not g44932 (n_20193, n27742);
  not g44933 (n_20194, n27746);
  and g44934 (n27747, n_20193, n_20194);
  not g44935 (n_20195, n27747);
  and g44936 (n27748, pi0787, n_20195);
  and g44937 (n27749, n_11803, n27738);
  not g44938 (n_20196, n27748);
  not g44939 (n_20197, n27749);
  and g44940 (n27750, n_20196, n_20197);
  not g44941 (n_20198, n27750);
  and g44942 (n27751, n_11819, n_20198);
  not g44943 (n_20199, n27751);
  and g44944 (n27752, pi0715, n_20199);
  and g44945 (n27753, pi0183, n_11417);
  and g44946 (n27754, n_15034, n17280);
  not g44947 (n_20200, n27754);
  and g44948 (n27755, n_20150, n_20200);
  not g44949 (n_20201, n27755);
  and g44950 (n27756, pi0038, n_20201);
  and g44951 (n27757, n_5709, n17221);
  and g44952 (n27758, pi0183, n_14476);
  not g44953 (n_20202, n27758);
  and g44954 (n27759, n_15034, n_20202);
  not g44955 (n_20203, n27757);
  and g44956 (n27760, n_20203, n27759);
  and g44957 (n27761, n_5709, pi0755);
  and g44958 (n27762, n_11739, n27761);
  not g44959 (n_20204, n27760);
  not g44960 (n_20205, n27762);
  and g44961 (n27763, n_20204, n_20205);
  not g44962 (n_20206, n27763);
  and g44963 (n27764, n_161, n_20206);
  not g44964 (n_20207, n27756);
  not g44965 (n_20208, n27764);
  and g44966 (n27765, n_20207, n_20208);
  and g44967 (n27766, n2571, n27765);
  not g44968 (n_20209, n27753);
  not g44969 (n_20210, n27766);
  and g44970 (n27767, n_20209, n_20210);
  not g44971 (n_20211, n27767);
  and g44972 (n27768, n_11960, n_20211);
  and g44973 (n27769, n17117, n_20148);
  not g44974 (n_20212, n27768);
  not g44975 (n_20213, n27769);
  and g44976 (n27770, n_20212, n_20213);
  not g44977 (n_20214, n27770);
  and g44978 (n27771, n_11964, n_20214);
  and g44979 (n27772, n_11967, n_20148);
  and g44980 (n27773, pi0609, n27768);
  not g44981 (n_20215, n27772);
  not g44982 (n_20216, n27773);
  and g44983 (n27774, n_20215, n_20216);
  not g44984 (n_20217, n27774);
  and g44985 (n27775, pi1155, n_20217);
  and g44986 (n27776, n_11972, n_20148);
  and g44987 (n27777, n_11971, n27768);
  not g44988 (n_20218, n27776);
  not g44989 (n_20219, n27777);
  and g44990 (n27778, n_20218, n_20219);
  not g44991 (n_20220, n27778);
  and g44992 (n27779, n_11768, n_20220);
  not g44993 (n_20221, n27775);
  not g44994 (n_20222, n27779);
  and g44995 (n27780, n_20221, n_20222);
  not g44996 (n_20223, n27780);
  and g44997 (n27781, pi0785, n_20223);
  not g44998 (n_20224, n27771);
  not g44999 (n_20225, n27781);
  and g45000 (n27782, n_20224, n_20225);
  not g45001 (n_20226, n27782);
  and g45002 (n27783, n_11981, n_20226);
  and g45003 (n27784, n_11984, n27690);
  and g45004 (n27785, pi0618, n27782);
  not g45005 (n_20227, n27784);
  and g45006 (n27786, pi1154, n_20227);
  not g45007 (n_20228, n27785);
  and g45008 (n27787, n_20228, n27786);
  and g45009 (n27788, n_11984, n27782);
  and g45010 (n27789, pi0618, n27690);
  not g45011 (n_20229, n27789);
  and g45012 (n27790, n_11413, n_20229);
  not g45013 (n_20230, n27788);
  and g45014 (n27791, n_20230, n27790);
  not g45015 (n_20231, n27787);
  not g45016 (n_20232, n27791);
  and g45017 (n27792, n_20231, n_20232);
  not g45018 (n_20233, n27792);
  and g45019 (n27793, pi0781, n_20233);
  not g45020 (n_20234, n27783);
  not g45021 (n_20235, n27793);
  and g45022 (n27794, n_20234, n_20235);
  not g45023 (n_20236, n27794);
  and g45024 (n27795, n_12315, n_20236);
  and g45025 (n27796, n_11821, n27690);
  and g45026 (n27797, pi0619, n27794);
  not g45027 (n_20237, n27796);
  and g45028 (n27798, pi1159, n_20237);
  not g45029 (n_20238, n27797);
  and g45030 (n27799, n_20238, n27798);
  and g45031 (n27800, n_11821, n27794);
  and g45032 (n27801, pi0619, n27690);
  not g45033 (n_20239, n27801);
  and g45034 (n27802, n_11405, n_20239);
  not g45035 (n_20240, n27800);
  and g45036 (n27803, n_20240, n27802);
  not g45037 (n_20241, n27799);
  not g45038 (n_20242, n27803);
  and g45039 (n27804, n_20241, n_20242);
  not g45040 (n_20243, n27804);
  and g45041 (n27805, pi0789, n_20243);
  not g45042 (n_20244, n27795);
  not g45043 (n_20245, n27805);
  and g45044 (n27806, n_20244, n_20245);
  and g45045 (n27807, n_12524, n27806);
  and g45046 (n27808, n17969, n27690);
  not g45047 (n_20246, n27807);
  not g45048 (n_20247, n27808);
  and g45049 (n27809, n_20246, n_20247);
  not g45050 (n_20248, n27809);
  and g45051 (n27810, n_12368, n_20248);
  and g45052 (n27811, n17779, n27690);
  not g45053 (n_20249, n27810);
  not g45054 (n_20250, n27811);
  and g45055 (n27812, n_20249, n_20250);
  not g45056 (n_20251, n27812);
  and g45057 (n27813, n_12392, n_20251);
  and g45058 (n27814, n17804, n27690);
  not g45059 (n_20252, n27813);
  not g45060 (n_20253, n27814);
  and g45061 (n27815, n_20252, n_20253);
  not g45062 (n_20254, n27815);
  and g45063 (n27816, pi0644, n_20254);
  and g45064 (n27817, n_11819, n27690);
  not g45065 (n_20255, n27817);
  and g45066 (n27818, n_12395, n_20255);
  not g45067 (n_20256, n27816);
  and g45068 (n27819, n_20256, n27818);
  not g45069 (n_20257, n27819);
  and g45070 (n27820, pi1160, n_20257);
  not g45071 (n_20258, n27752);
  and g45072 (n27821, n_20258, n27820);
  and g45073 (n27822, pi0644, n_20198);
  not g45074 (n_20259, n27822);
  and g45075 (n27823, n_12395, n_20259);
  and g45076 (n27824, n_11819, n_20254);
  and g45077 (n27825, pi0644, n27690);
  not g45078 (n_20260, n27825);
  and g45079 (n27826, pi0715, n_20260);
  not g45080 (n_20261, n27824);
  and g45081 (n27827, n_20261, n27826);
  not g45082 (n_20262, n27827);
  and g45083 (n27828, n_12405, n_20262);
  not g45084 (n_20263, n27823);
  and g45085 (n27829, n_20263, n27828);
  not g45086 (n_20264, n27821);
  not g45087 (n_20265, n27829);
  and g45088 (n27830, n_20264, n_20265);
  not g45089 (n_20266, n27830);
  and g45090 (n27831, pi0790, n_20266);
  and g45091 (n27832, n_12354, n27731);
  and g45092 (n27833, n_14557, n27809);
  and g45093 (n27834, pi0629, n27735);
  not g45094 (n_20267, n27832);
  not g45095 (n_20268, n27834);
  and g45096 (n27835, n_20267, n_20268);
  not g45097 (n_20269, n27833);
  and g45098 (n27836, n_20269, n27835);
  not g45099 (n_20270, n27836);
  and g45100 (n27837, pi0792, n_20270);
  and g45101 (n27838, pi0609, n27715);
  and g45102 (n27839, pi0183, n_12240);
  and g45103 (n27840, n_5709, n_12230);
  not g45104 (n_20271, n27839);
  and g45105 (n27841, pi0755, n_20271);
  not g45106 (n_20272, n27840);
  and g45107 (n27842, n_20272, n27841);
  and g45108 (n27843, n_5709, n17629);
  and g45109 (n27844, pi0183, n17631);
  not g45110 (n_20273, n27844);
  and g45111 (n27845, n_15034, n_20273);
  not g45112 (n_20274, n27843);
  and g45113 (n27846, n_20274, n27845);
  not g45114 (n_20275, n27842);
  not g45115 (n_20276, n27846);
  and g45116 (n27847, n_20275, n_20276);
  not g45117 (n_20277, n27847);
  and g45118 (n27848, n_162, n_20277);
  and g45119 (n27849, pi0183, n17605);
  and g45120 (n27850, n_5709, n_12180);
  not g45121 (n_20278, n27850);
  and g45122 (n27851, n_15034, n_20278);
  not g45123 (n_20279, n27849);
  and g45124 (n27852, n_20279, n27851);
  and g45125 (n27853, n_5709, n17404);
  and g45126 (n27854, pi0183, n17485);
  not g45127 (n_20280, n27854);
  and g45128 (n27855, pi0755, n_20280);
  not g45129 (n_20281, n27853);
  and g45130 (n27856, n_20281, n27855);
  not g45131 (n_20282, n27852);
  and g45132 (n27857, pi0039, n_20282);
  not g45133 (n_20283, n27856);
  and g45134 (n27858, n_20283, n27857);
  not g45135 (n_20284, n27848);
  and g45136 (n27859, n_161, n_20284);
  not g45137 (n_20285, n27858);
  and g45138 (n27860, n_20285, n27859);
  and g45139 (n27861, n_15034, n_12250);
  not g45140 (n_20286, n27861);
  and g45141 (n27862, n19471, n_20286);
  not g45142 (n_20287, n27862);
  and g45143 (n27863, n_5709, n_20287);
  and g45144 (n27864, n_12120, n_20012);
  not g45145 (n_20288, n27864);
  and g45146 (n27865, pi0183, n_20288);
  and g45147 (n27866, n6284, n27865);
  not g45148 (n_20289, n27866);
  and g45149 (n27867, pi0038, n_20289);
  not g45150 (n_20290, n27863);
  and g45151 (n27868, n_20290, n27867);
  not g45152 (n_20291, n27868);
  and g45153 (n27869, n_15036, n_20291);
  not g45154 (n_20292, n27860);
  and g45155 (n27870, n_20292, n27869);
  not g45156 (n_20293, n27765);
  and g45157 (n27871, pi0725, n_20293);
  not g45158 (n_20294, n27870);
  and g45159 (n27872, n2571, n_20294);
  not g45160 (n_20295, n27871);
  and g45161 (n27873, n_20295, n27872);
  not g45162 (n_20296, n27873);
  and g45163 (n27874, n_20209, n_20296);
  and g45164 (n27875, n_11753, n27874);
  and g45165 (n27876, pi0625, n27767);
  not g45166 (n_20297, n27876);
  and g45167 (n27877, n_11757, n_20297);
  not g45168 (n_20298, n27875);
  and g45169 (n27878, n_20298, n27877);
  and g45170 (n27879, n_11823, n_20164);
  not g45171 (n_20299, n27878);
  and g45172 (n27880, n_20299, n27879);
  and g45173 (n27881, n_11753, n27767);
  and g45174 (n27882, pi0625, n27874);
  not g45175 (n_20300, n27881);
  and g45176 (n27883, pi1153, n_20300);
  not g45177 (n_20301, n27882);
  and g45178 (n27884, n_20301, n27883);
  and g45179 (n27885, pi0608, n_20165);
  not g45180 (n_20302, n27884);
  and g45181 (n27886, n_20302, n27885);
  not g45182 (n_20303, n27880);
  not g45183 (n_20304, n27886);
  and g45184 (n27887, n_20303, n_20304);
  not g45185 (n_20305, n27887);
  and g45186 (n27888, pi0778, n_20305);
  and g45187 (n27889, n_11749, n27874);
  not g45188 (n_20306, n27888);
  not g45189 (n_20307, n27889);
  and g45190 (n27890, n_20306, n_20307);
  not g45191 (n_20308, n27890);
  and g45192 (n27891, n_11971, n_20308);
  not g45193 (n_20309, n27838);
  and g45194 (n27892, n_11768, n_20309);
  not g45195 (n_20310, n27891);
  and g45196 (n27893, n_20310, n27892);
  and g45197 (n27894, n_11767, n_20221);
  not g45198 (n_20311, n27893);
  and g45199 (n27895, n_20311, n27894);
  and g45200 (n27896, n_11971, n27715);
  and g45201 (n27897, pi0609, n_20308);
  not g45202 (n_20312, n27896);
  and g45203 (n27898, pi1155, n_20312);
  not g45204 (n_20313, n27897);
  and g45205 (n27899, n_20313, n27898);
  and g45206 (n27900, pi0660, n_20222);
  not g45207 (n_20314, n27899);
  and g45208 (n27901, n_20314, n27900);
  not g45209 (n_20315, n27895);
  not g45210 (n_20316, n27901);
  and g45211 (n27902, n_20315, n_20316);
  not g45212 (n_20317, n27902);
  and g45213 (n27903, pi0785, n_20317);
  and g45214 (n27904, n_11964, n_20308);
  not g45215 (n_20318, n27903);
  not g45216 (n_20319, n27904);
  and g45217 (n27905, n_20318, n_20319);
  not g45218 (n_20320, n27905);
  and g45219 (n27906, n_11984, n_20320);
  and g45220 (n27907, pi0618, n27718);
  not g45221 (n_20321, n27907);
  and g45222 (n27908, n_11413, n_20321);
  not g45223 (n_20322, n27906);
  and g45224 (n27909, n_20322, n27908);
  and g45225 (n27910, n_11412, n_20231);
  not g45226 (n_20323, n27909);
  and g45227 (n27911, n_20323, n27910);
  and g45228 (n27912, n_11984, n27718);
  and g45229 (n27913, pi0618, n_20320);
  not g45230 (n_20324, n27912);
  and g45231 (n27914, pi1154, n_20324);
  not g45232 (n_20325, n27913);
  and g45233 (n27915, n_20325, n27914);
  and g45234 (n27916, pi0627, n_20232);
  not g45235 (n_20326, n27915);
  and g45236 (n27917, n_20326, n27916);
  not g45237 (n_20327, n27911);
  not g45238 (n_20328, n27917);
  and g45239 (n27918, n_20327, n_20328);
  not g45240 (n_20329, n27918);
  and g45241 (n27919, pi0781, n_20329);
  and g45242 (n27920, n_11981, n_20320);
  not g45243 (n_20330, n27919);
  not g45244 (n_20331, n27920);
  and g45245 (n27921, n_20330, n_20331);
  and g45246 (n27922, n_12315, n27921);
  not g45247 (n_20332, n27721);
  and g45248 (n27923, pi0619, n_20332);
  not g45249 (n_20333, n27921);
  and g45250 (n27924, n_11821, n_20333);
  not g45251 (n_20334, n27923);
  and g45252 (n27925, n_11405, n_20334);
  not g45253 (n_20335, n27924);
  and g45254 (n27926, n_20335, n27925);
  and g45255 (n27927, n_11403, n_20241);
  not g45256 (n_20336, n27926);
  and g45257 (n27928, n_20336, n27927);
  and g45258 (n27929, n_11821, n_20332);
  and g45259 (n27930, pi0619, n_20333);
  not g45260 (n_20337, n27929);
  and g45261 (n27931, pi1159, n_20337);
  not g45262 (n_20338, n27930);
  and g45263 (n27932, n_20338, n27931);
  and g45264 (n27933, pi0648, n_20242);
  not g45265 (n_20339, n27932);
  and g45266 (n27934, n_20339, n27933);
  not g45267 (n_20340, n27928);
  and g45268 (n27935, pi0789, n_20340);
  not g45269 (n_20341, n27934);
  and g45270 (n27936, n_20341, n27935);
  not g45271 (n_20342, n27922);
  and g45272 (n27937, n17970, n_20342);
  not g45273 (n_20343, n27936);
  and g45274 (n27938, n_20343, n27937);
  and g45275 (n27939, n17871, n27723);
  not g45276 (n_20344, n27806);
  and g45277 (n27940, n_12320, n_20344);
  and g45278 (n27941, pi0626, n_20148);
  not g45279 (n_20345, n27941);
  and g45280 (n27942, n16629, n_20345);
  not g45281 (n_20346, n27940);
  and g45282 (n27943, n_20346, n27942);
  and g45283 (n27944, pi0626, n_20344);
  and g45284 (n27945, n_12320, n_20148);
  not g45285 (n_20347, n27945);
  and g45286 (n27946, n16628, n_20347);
  not g45287 (n_20348, n27944);
  and g45288 (n27947, n_20348, n27946);
  not g45289 (n_20349, n27939);
  not g45290 (n_20350, n27943);
  and g45291 (n27948, n_20349, n_20350);
  not g45292 (n_20351, n27947);
  and g45293 (n27949, n_20351, n27948);
  not g45294 (n_20352, n27949);
  and g45295 (n27950, pi0788, n_20352);
  not g45296 (n_20353, n27950);
  and g45297 (n27951, n_14638, n_20353);
  not g45298 (n_20354, n27938);
  and g45299 (n27952, n_20354, n27951);
  not g45300 (n_20355, n27837);
  not g45301 (n_20356, n27952);
  and g45302 (n27953, n_20355, n_20356);
  not g45303 (n_20357, n27953);
  and g45304 (n27954, n_14387, n_20357);
  not g45305 (n_20358, n27741);
  and g45306 (n27955, n17802, n_20358);
  and g45307 (n27956, n_14548, n27812);
  not g45308 (n_20359, n27745);
  and g45309 (n27957, n17801, n_20359);
  not g45310 (n_20360, n27955);
  not g45311 (n_20361, n27957);
  and g45312 (n27958, n_20360, n_20361);
  not g45313 (n_20362, n27956);
  and g45314 (n27959, n_20362, n27958);
  not g45315 (n_20363, n27959);
  and g45316 (n27960, pi0787, n_20363);
  and g45317 (n27961, n_11819, n27828);
  and g45318 (n27962, pi0644, n27820);
  not g45319 (n_20364, n27961);
  and g45320 (n27963, pi0790, n_20364);
  not g45321 (n_20365, n27962);
  and g45322 (n27964, n_20365, n27963);
  not g45323 (n_20366, n27954);
  not g45324 (n_20367, n27960);
  and g45325 (n27965, n_20366, n_20367);
  not g45326 (n_20368, n27964);
  and g45327 (n27966, n_20368, n27965);
  not g45328 (n_20369, n27831);
  not g45329 (n_20370, n27966);
  and g45330 (n27967, n_20369, n_20370);
  not g45331 (n_20371, n27967);
  and g45332 (n27968, n_4226, n_20371);
  not g45333 (n_20372, n27689);
  and g45334 (n27969, n_12415, n_20372);
  not g45335 (n_20373, n27968);
  and g45336 (n27970, n_20373, n27969);
  not g45337 (n_20374, n27688);
  not g45338 (n_20375, n27970);
  and g45339 (po0340, n_20374, n_20375);
  and g45340 (n27972, n_7617, n_12418);
  and g45341 (n27973, n_15732, n16645);
  not g45342 (n_20376, n27972);
  not g45343 (n_20377, n27973);
  and g45344 (n27974, n_20376, n_20377);
  not g45345 (n_20378, n27974);
  and g45346 (n27975, n_11749, n_20378);
  and g45347 (n27976, n_11753, n27973);
  not g45348 (n_20379, n27976);
  and g45349 (n27977, n_20378, n_20379);
  not g45350 (n_20380, n27977);
  and g45351 (n27978, pi1153, n_20380);
  and g45352 (n27979, n_11757, n_20376);
  and g45353 (n27980, n_20379, n27979);
  not g45354 (n_20381, n27980);
  and g45355 (n27981, pi0778, n_20381);
  not g45356 (n_20382, n27978);
  and g45357 (n27982, n_20382, n27981);
  not g45358 (n_20383, n27975);
  not g45359 (n_20384, n27982);
  and g45360 (n27983, n_20383, n_20384);
  not g45361 (n_20385, n27983);
  and g45362 (n27984, n_12429, n_20385);
  and g45363 (n27985, n_12430, n27984);
  and g45364 (n27986, n_12431, n27985);
  and g45365 (n27987, n_12432, n27986);
  and g45366 (n27988, n_12436, n27987);
  and g45367 (n27989, n_11806, n27988);
  and g45368 (n27990, pi0647, n27972);
  not g45369 (n_20386, n27990);
  and g45370 (n27991, n_11810, n_20386);
  not g45371 (n_20387, n27989);
  and g45372 (n27992, n_20387, n27991);
  and g45373 (n27993, pi0630, n27992);
  and g45374 (n27994, n_15730, n17244);
  not g45375 (n_20388, n27994);
  and g45376 (n27995, n_20376, n_20388);
  not g45377 (n_20389, n27995);
  and g45378 (n27996, n_12448, n_20389);
  not g45379 (n_20390, n27996);
  and g45380 (n27997, n_11964, n_20390);
  and g45381 (n27998, n17296, n27994);
  not g45382 (n_20391, n27998);
  and g45383 (n27999, n27996, n_20391);
  not g45384 (n_20392, n27999);
  and g45385 (n28000, pi1155, n_20392);
  and g45386 (n28001, n_11768, n_20376);
  and g45387 (n28002, n_20391, n28001);
  not g45388 (n_20393, n28000);
  not g45389 (n_20394, n28002);
  and g45390 (n28003, n_20393, n_20394);
  not g45391 (n_20395, n28003);
  and g45392 (n28004, pi0785, n_20395);
  not g45393 (n_20396, n27997);
  not g45394 (n_20397, n28004);
  and g45395 (n28005, n_20396, n_20397);
  not g45396 (n_20398, n28005);
  and g45397 (n28006, n_11981, n_20398);
  and g45398 (n28007, n_12461, n28005);
  not g45399 (n_20399, n28007);
  and g45400 (n28008, pi1154, n_20399);
  and g45401 (n28009, n_12463, n28005);
  not g45402 (n_20400, n28009);
  and g45403 (n28010, n_11413, n_20400);
  not g45404 (n_20401, n28008);
  not g45405 (n_20402, n28010);
  and g45406 (n28011, n_20401, n_20402);
  not g45407 (n_20403, n28011);
  and g45408 (n28012, pi0781, n_20403);
  not g45409 (n_20404, n28006);
  not g45410 (n_20405, n28012);
  and g45411 (n28013, n_20404, n_20405);
  not g45412 (n_20406, n28013);
  and g45413 (n28014, n_12315, n_20406);
  and g45414 (n28015, n_16503, n28013);
  not g45415 (n_20407, n28015);
  and g45416 (n28016, pi1159, n_20407);
  and g45417 (n28017, n_16505, n28013);
  not g45418 (n_20408, n28017);
  and g45419 (n28018, n_11405, n_20408);
  not g45420 (n_20409, n28016);
  not g45421 (n_20410, n28018);
  and g45422 (n28019, n_20409, n_20410);
  not g45423 (n_20411, n28019);
  and g45424 (n28020, pi0789, n_20411);
  not g45425 (n_20412, n28014);
  not g45426 (n_20413, n28020);
  and g45427 (n28021, n_20412, n_20413);
  and g45428 (n28022, n_12524, n28021);
  and g45429 (n28023, n17969, n27972);
  not g45430 (n_20414, n28022);
  not g45431 (n_20415, n28023);
  and g45432 (n28024, n_20414, n_20415);
  not g45433 (n_20416, n28024);
  and g45434 (n28025, n_12368, n_20416);
  and g45435 (n28026, n17779, n27972);
  not g45436 (n_20417, n28025);
  not g45437 (n_20418, n28026);
  and g45438 (n28027, n_20417, n_20418);
  and g45439 (n28028, n_14548, n28027);
  not g45440 (n_20419, n27988);
  and g45441 (n28029, pi0647, n_20419);
  and g45442 (n28030, n_11806, n_20376);
  not g45443 (n_20420, n28029);
  not g45444 (n_20421, n28030);
  and g45445 (n28031, n_20420, n_20421);
  not g45446 (n_20422, n28031);
  and g45447 (n28032, n17801, n_20422);
  not g45448 (n_20423, n27993);
  not g45449 (n_20424, n28032);
  and g45450 (n28033, n_20423, n_20424);
  not g45451 (n_20425, n28028);
  and g45452 (n28034, n_20425, n28033);
  not g45453 (n_20426, n28034);
  and g45454 (n28035, pi0787, n_20426);
  and g45455 (n28036, n17871, n27986);
  not g45456 (n_20427, n28021);
  and g45457 (n28037, n_12320, n_20427);
  and g45458 (n28038, pi0626, n_20376);
  not g45459 (n_20428, n28038);
  and g45460 (n28039, n16629, n_20428);
  not g45461 (n_20429, n28037);
  and g45462 (n28040, n_20429, n28039);
  and g45463 (n28041, pi0626, n_20427);
  and g45464 (n28042, n_12320, n_20376);
  not g45465 (n_20430, n28042);
  and g45466 (n28043, n16628, n_20430);
  not g45467 (n_20431, n28041);
  and g45468 (n28044, n_20431, n28043);
  not g45469 (n_20432, n28036);
  not g45470 (n_20433, n28040);
  and g45471 (n28045, n_20432, n_20433);
  not g45472 (n_20434, n28044);
  and g45473 (n28046, n_20434, n28045);
  not g45474 (n_20435, n28046);
  and g45475 (n28047, pi0788, n_20435);
  and g45476 (n28048, pi0618, n27984);
  and g45477 (n28049, n_11866, n_20378);
  and g45478 (n28050, pi0625, n28049);
  not g45479 (n_20436, n28049);
  and g45480 (n28051, n27995, n_20436);
  not g45481 (n_20437, n28050);
  not g45482 (n_20438, n28051);
  and g45483 (n28052, n_20437, n_20438);
  not g45484 (n_20439, n28052);
  and g45485 (n28053, n27979, n_20439);
  and g45486 (n28054, n_11823, n_20382);
  not g45487 (n_20440, n28053);
  and g45488 (n28055, n_20440, n28054);
  and g45489 (n28056, pi1153, n27995);
  and g45490 (n28057, n_20437, n28056);
  and g45491 (n28058, pi0608, n_20381);
  not g45492 (n_20441, n28057);
  and g45493 (n28059, n_20441, n28058);
  not g45494 (n_20442, n28055);
  not g45495 (n_20443, n28059);
  and g45496 (n28060, n_20442, n_20443);
  not g45497 (n_20444, n28060);
  and g45498 (n28061, pi0778, n_20444);
  and g45499 (n28062, n_11749, n_20438);
  not g45500 (n_20445, n28061);
  not g45501 (n_20446, n28062);
  and g45502 (n28063, n_20445, n_20446);
  not g45503 (n_20447, n28063);
  and g45504 (n28064, n_11971, n_20447);
  and g45505 (n28065, pi0609, n_20385);
  not g45506 (n_20448, n28065);
  and g45507 (n28066, n_11768, n_20448);
  not g45508 (n_20449, n28064);
  and g45509 (n28067, n_20449, n28066);
  and g45510 (n28068, n_11767, n_20393);
  not g45511 (n_20450, n28067);
  and g45512 (n28069, n_20450, n28068);
  and g45513 (n28070, pi0609, n_20447);
  and g45514 (n28071, n_11971, n_20385);
  not g45515 (n_20451, n28071);
  and g45516 (n28072, pi1155, n_20451);
  not g45517 (n_20452, n28070);
  and g45518 (n28073, n_20452, n28072);
  and g45519 (n28074, pi0660, n_20394);
  not g45520 (n_20453, n28073);
  and g45521 (n28075, n_20453, n28074);
  not g45522 (n_20454, n28069);
  not g45523 (n_20455, n28075);
  and g45524 (n28076, n_20454, n_20455);
  not g45525 (n_20456, n28076);
  and g45526 (n28077, pi0785, n_20456);
  and g45527 (n28078, n_11964, n_20447);
  not g45528 (n_20457, n28077);
  not g45529 (n_20458, n28078);
  and g45530 (n28079, n_20457, n_20458);
  not g45531 (n_20459, n28079);
  and g45532 (n28080, n_11984, n_20459);
  not g45533 (n_20460, n28048);
  and g45534 (n28081, n_11413, n_20460);
  not g45535 (n_20461, n28080);
  and g45536 (n28082, n_20461, n28081);
  and g45537 (n28083, n_11412, n_20401);
  not g45538 (n_20462, n28082);
  and g45539 (n28084, n_20462, n28083);
  and g45540 (n28085, n_11984, n27984);
  and g45541 (n28086, pi0618, n_20459);
  not g45542 (n_20463, n28085);
  and g45543 (n28087, pi1154, n_20463);
  not g45544 (n_20464, n28086);
  and g45545 (n28088, n_20464, n28087);
  and g45546 (n28089, pi0627, n_20402);
  not g45547 (n_20465, n28088);
  and g45548 (n28090, n_20465, n28089);
  not g45549 (n_20466, n28084);
  not g45550 (n_20467, n28090);
  and g45551 (n28091, n_20466, n_20467);
  not g45552 (n_20468, n28091);
  and g45553 (n28092, pi0781, n_20468);
  and g45554 (n28093, n_11981, n_20459);
  not g45555 (n_20469, n28092);
  not g45556 (n_20470, n28093);
  and g45557 (n28094, n_20469, n_20470);
  and g45558 (n28095, n_12315, n28094);
  not g45559 (n_20471, n28094);
  and g45560 (n28096, n_11821, n_20471);
  and g45561 (n28097, pi0619, n27985);
  not g45562 (n_20472, n28097);
  and g45563 (n28098, n_11405, n_20472);
  not g45564 (n_20473, n28096);
  and g45565 (n28099, n_20473, n28098);
  and g45566 (n28100, n_11403, n_20409);
  not g45567 (n_20474, n28099);
  and g45568 (n28101, n_20474, n28100);
  and g45569 (n28102, pi0619, n_20471);
  and g45570 (n28103, n_11821, n27985);
  not g45571 (n_20475, n28103);
  and g45572 (n28104, pi1159, n_20475);
  not g45573 (n_20476, n28102);
  and g45574 (n28105, n_20476, n28104);
  and g45575 (n28106, pi0648, n_20410);
  not g45576 (n_20477, n28105);
  and g45577 (n28107, n_20477, n28106);
  not g45578 (n_20478, n28101);
  and g45579 (n28108, pi0789, n_20478);
  not g45580 (n_20479, n28107);
  and g45581 (n28109, n_20479, n28108);
  not g45582 (n_20480, n28095);
  and g45583 (n28110, n17970, n_20480);
  not g45584 (n_20481, n28109);
  and g45585 (n28111, n_20481, n28110);
  not g45586 (n_20482, n28047);
  not g45587 (n_20483, n28111);
  and g45588 (n28112, n_20482, n_20483);
  not g45589 (n_20484, n28112);
  and g45590 (n28113, n_14638, n_20484);
  and g45591 (n28114, n17854, n_20416);
  and g45592 (n28115, n20851, n27987);
  not g45593 (n_20485, n28114);
  not g45594 (n_20486, n28115);
  and g45595 (n28116, n_20485, n_20486);
  not g45596 (n_20487, n28116);
  and g45597 (n28117, n_12354, n_20487);
  and g45598 (n28118, n20855, n27987);
  and g45599 (n28119, n17853, n_20416);
  not g45600 (n_20488, n28118);
  not g45601 (n_20489, n28119);
  and g45602 (n28120, n_20488, n_20489);
  not g45603 (n_20490, n28120);
  and g45604 (n28121, pi0629, n_20490);
  not g45605 (n_20491, n28117);
  not g45606 (n_20492, n28121);
  and g45607 (n28122, n_20491, n_20492);
  not g45608 (n_20493, n28122);
  and g45609 (n28123, pi0792, n_20493);
  not g45610 (n_20494, n28123);
  and g45611 (n28124, n_14387, n_20494);
  not g45612 (n_20495, n28113);
  and g45613 (n28125, n_20495, n28124);
  not g45614 (n_20496, n28035);
  not g45615 (n_20497, n28125);
  and g45616 (n28126, n_20496, n_20497);
  and g45617 (n28127, n_12411, n28126);
  and g45618 (n28128, n_11803, n_20419);
  and g45619 (n28129, pi1157, n_20422);
  not g45620 (n_20498, n27992);
  not g45621 (n_20499, n28129);
  and g45622 (n28130, n_20498, n_20499);
  not g45623 (n_20500, n28130);
  and g45624 (n28131, pi0787, n_20500);
  not g45625 (n_20501, n28128);
  not g45626 (n_20502, n28131);
  and g45627 (n28132, n_20501, n_20502);
  and g45628 (n28133, n_11819, n28132);
  and g45629 (n28134, pi0644, n28126);
  not g45630 (n_20503, n28133);
  and g45631 (n28135, pi0715, n_20503);
  not g45632 (n_20504, n28134);
  and g45633 (n28136, n_20504, n28135);
  not g45634 (n_20505, n28027);
  and g45635 (n28137, n_12392, n_20505);
  and g45636 (n28138, n17804, n27972);
  not g45637 (n_20506, n28137);
  not g45638 (n_20507, n28138);
  and g45639 (n28139, n_20506, n_20507);
  not g45640 (n_20508, n28139);
  and g45641 (n28140, pi0644, n_20508);
  and g45642 (n28141, n_11819, n27972);
  not g45643 (n_20509, n28141);
  and g45644 (n28142, n_12395, n_20509);
  not g45645 (n_20510, n28140);
  and g45646 (n28143, n_20510, n28142);
  not g45647 (n_20511, n28143);
  and g45648 (n28144, pi1160, n_20511);
  not g45649 (n_20512, n28136);
  and g45650 (n28145, n_20512, n28144);
  and g45651 (n28146, n_11819, n_20508);
  and g45652 (n28147, pi0644, n27972);
  not g45653 (n_20513, n28147);
  and g45654 (n28148, pi0715, n_20513);
  not g45655 (n_20514, n28146);
  and g45656 (n28149, n_20514, n28148);
  and g45657 (n28150, pi0644, n28132);
  and g45658 (n28151, n_11819, n28126);
  not g45659 (n_20515, n28150);
  and g45660 (n28152, n_12395, n_20515);
  not g45661 (n_20516, n28151);
  and g45662 (n28153, n_20516, n28152);
  not g45663 (n_20517, n28149);
  and g45664 (n28154, n_12405, n_20517);
  not g45665 (n_20518, n28153);
  and g45666 (n28155, n_20518, n28154);
  not g45667 (n_20519, n28145);
  not g45668 (n_20520, n28155);
  and g45669 (n28156, n_20519, n_20520);
  not g45670 (n_20521, n28156);
  and g45671 (n28157, pi0790, n_20521);
  not g45672 (n_20522, n28127);
  and g45673 (n28158, pi0832, n_20522);
  not g45674 (n_20523, n28157);
  and g45675 (n28159, n_20523, n28158);
  and g45676 (n28160, n_7617, po1038);
  and g45677 (n28161, n_7617, n_11751);
  not g45678 (n_20524, n28161);
  and g45679 (n28162, n16635, n_20524);
  and g45680 (n28163, n_15732, n2571);
  not g45681 (n_20525, n28163);
  and g45682 (n28164, n28161, n_20525);
  and g45683 (n28165, n_7617, n_11418);
  not g45684 (n_20526, n28165);
  and g45685 (n28166, n16647, n_20526);
  and g45686 (n28167, pi0184, n_12608);
  not g45687 (n_20527, n28167);
  and g45688 (n28168, n_161, n_20527);
  not g45689 (n_20528, n28168);
  and g45690 (n28169, n2571, n_20528);
  and g45691 (n28170, n_7617, n18072);
  not g45692 (n_20529, n28169);
  not g45693 (n_20530, n28170);
  and g45694 (n28171, n_20529, n_20530);
  not g45695 (n_20531, n28166);
  and g45696 (n28172, n_15732, n_20531);
  not g45697 (n_20532, n28171);
  and g45698 (n28173, n_20532, n28172);
  not g45699 (n_20533, n28164);
  not g45700 (n_20534, n28173);
  and g45701 (n28174, n_20533, n_20534);
  and g45702 (n28175, n_11749, n28174);
  and g45703 (n28176, n_11753, n28161);
  not g45704 (n_20535, n28174);
  and g45705 (n28177, pi0625, n_20535);
  not g45706 (n_20536, n28176);
  and g45707 (n28178, pi1153, n_20536);
  not g45708 (n_20537, n28177);
  and g45709 (n28179, n_20537, n28178);
  and g45710 (n28180, pi0625, n28161);
  and g45711 (n28181, n_11753, n_20535);
  not g45712 (n_20538, n28180);
  and g45713 (n28182, n_11757, n_20538);
  not g45714 (n_20539, n28181);
  and g45715 (n28183, n_20539, n28182);
  not g45716 (n_20540, n28179);
  not g45717 (n_20541, n28183);
  and g45718 (n28184, n_20540, n_20541);
  not g45719 (n_20542, n28184);
  and g45720 (n28185, pi0778, n_20542);
  not g45721 (n_20543, n28175);
  not g45722 (n_20544, n28185);
  and g45723 (n28186, n_20543, n_20544);
  not g45724 (n_20545, n28186);
  and g45725 (n28187, n_11773, n_20545);
  and g45726 (n28188, n17075, n_20524);
  not g45727 (n_20546, n28187);
  not g45728 (n_20547, n28188);
  and g45729 (n28189, n_20546, n_20547);
  and g45730 (n28190, n_11777, n28189);
  and g45731 (n28191, n16639, n28161);
  not g45732 (n_20548, n28190);
  not g45733 (n_20549, n28191);
  and g45734 (n28192, n_20548, n_20549);
  and g45735 (n28193, n_11780, n28192);
  not g45736 (n_20550, n28162);
  not g45737 (n_20551, n28193);
  and g45738 (n28194, n_20550, n_20551);
  and g45739 (n28195, n_11783, n28194);
  and g45740 (n28196, n16631, n28161);
  not g45741 (n_20552, n28195);
  not g45742 (n_20553, n28196);
  and g45743 (n28197, n_20552, n_20553);
  and g45744 (n28198, n_11787, n28197);
  not g45745 (n_20554, n28197);
  and g45746 (n28199, pi0628, n_20554);
  and g45747 (n28200, n_11789, n28161);
  not g45748 (n_20555, n28200);
  and g45749 (n28201, pi1156, n_20555);
  not g45750 (n_20556, n28199);
  and g45751 (n28202, n_20556, n28201);
  and g45752 (n28203, pi0628, n28161);
  and g45753 (n28204, n_11789, n_20554);
  not g45754 (n_20557, n28203);
  and g45755 (n28205, n_11794, n_20557);
  not g45756 (n_20558, n28204);
  and g45757 (n28206, n_20558, n28205);
  not g45758 (n_20559, n28202);
  not g45759 (n_20560, n28206);
  and g45760 (n28207, n_20559, n_20560);
  not g45761 (n_20561, n28207);
  and g45762 (n28208, pi0792, n_20561);
  not g45763 (n_20562, n28198);
  not g45764 (n_20563, n28208);
  and g45765 (n28209, n_20562, n_20563);
  not g45766 (n_20564, n28209);
  and g45767 (n28210, n_11806, n_20564);
  and g45768 (n28211, pi0647, n_20524);
  not g45769 (n_20565, n28210);
  not g45770 (n_20566, n28211);
  and g45771 (n28212, n_20565, n_20566);
  and g45772 (n28213, n_11810, n28212);
  and g45773 (n28214, pi0647, n_20564);
  and g45774 (n28215, n_11806, n_20524);
  not g45775 (n_20567, n28214);
  not g45776 (n_20568, n28215);
  and g45777 (n28216, n_20567, n_20568);
  and g45778 (n28217, pi1157, n28216);
  not g45779 (n_20569, n28213);
  not g45780 (n_20570, n28217);
  and g45781 (n28218, n_20569, n_20570);
  not g45782 (n_20571, n28218);
  and g45783 (n28219, pi0787, n_20571);
  and g45784 (n28220, n_11803, n28209);
  not g45785 (n_20572, n28219);
  not g45786 (n_20573, n28220);
  and g45787 (n28221, n_20572, n_20573);
  not g45788 (n_20574, n28221);
  and g45789 (n28222, n_11819, n_20574);
  not g45790 (n_20575, n28222);
  and g45791 (n28223, pi0715, n_20575);
  and g45792 (n28224, pi0184, n_11417);
  and g45793 (n28225, n_15730, n17280);
  not g45794 (n_20576, n28225);
  and g45795 (n28226, n_20526, n_20576);
  not g45796 (n_20577, n28226);
  and g45797 (n28227, pi0038, n_20577);
  and g45798 (n28228, n_7617, n17221);
  and g45799 (n28229, pi0184, n_14476);
  not g45800 (n_20578, n28229);
  and g45801 (n28230, n_15730, n_20578);
  not g45802 (n_20579, n28228);
  and g45803 (n28231, n_20579, n28230);
  and g45804 (n28232, n_7617, pi0777);
  and g45805 (n28233, n_11739, n28232);
  not g45806 (n_20580, n28231);
  not g45807 (n_20581, n28233);
  and g45808 (n28234, n_20580, n_20581);
  not g45809 (n_20582, n28234);
  and g45810 (n28235, n_161, n_20582);
  not g45811 (n_20583, n28227);
  not g45812 (n_20584, n28235);
  and g45813 (n28236, n_20583, n_20584);
  and g45814 (n28237, n2571, n28236);
  not g45815 (n_20585, n28224);
  not g45816 (n_20586, n28237);
  and g45817 (n28238, n_20585, n_20586);
  not g45818 (n_20587, n28238);
  and g45819 (n28239, n_11960, n_20587);
  and g45820 (n28240, n17117, n_20524);
  not g45821 (n_20588, n28239);
  not g45822 (n_20589, n28240);
  and g45823 (n28241, n_20588, n_20589);
  not g45824 (n_20590, n28241);
  and g45825 (n28242, n_11964, n_20590);
  and g45826 (n28243, n_11967, n_20524);
  and g45827 (n28244, pi0609, n28239);
  not g45828 (n_20591, n28243);
  not g45829 (n_20592, n28244);
  and g45830 (n28245, n_20591, n_20592);
  not g45831 (n_20593, n28245);
  and g45832 (n28246, pi1155, n_20593);
  and g45833 (n28247, n_11972, n_20524);
  and g45834 (n28248, n_11971, n28239);
  not g45835 (n_20594, n28247);
  not g45836 (n_20595, n28248);
  and g45837 (n28249, n_20594, n_20595);
  not g45838 (n_20596, n28249);
  and g45839 (n28250, n_11768, n_20596);
  not g45840 (n_20597, n28246);
  not g45841 (n_20598, n28250);
  and g45842 (n28251, n_20597, n_20598);
  not g45843 (n_20599, n28251);
  and g45844 (n28252, pi0785, n_20599);
  not g45845 (n_20600, n28242);
  not g45846 (n_20601, n28252);
  and g45847 (n28253, n_20600, n_20601);
  not g45848 (n_20602, n28253);
  and g45849 (n28254, n_11981, n_20602);
  and g45850 (n28255, n_11984, n28161);
  and g45851 (n28256, pi0618, n28253);
  not g45852 (n_20603, n28255);
  and g45853 (n28257, pi1154, n_20603);
  not g45854 (n_20604, n28256);
  and g45855 (n28258, n_20604, n28257);
  and g45856 (n28259, n_11984, n28253);
  and g45857 (n28260, pi0618, n28161);
  not g45858 (n_20605, n28260);
  and g45859 (n28261, n_11413, n_20605);
  not g45860 (n_20606, n28259);
  and g45861 (n28262, n_20606, n28261);
  not g45862 (n_20607, n28258);
  not g45863 (n_20608, n28262);
  and g45864 (n28263, n_20607, n_20608);
  not g45865 (n_20609, n28263);
  and g45866 (n28264, pi0781, n_20609);
  not g45867 (n_20610, n28254);
  not g45868 (n_20611, n28264);
  and g45869 (n28265, n_20610, n_20611);
  not g45870 (n_20612, n28265);
  and g45871 (n28266, n_12315, n_20612);
  and g45872 (n28267, n_11821, n28161);
  and g45873 (n28268, pi0619, n28265);
  not g45874 (n_20613, n28267);
  and g45875 (n28269, pi1159, n_20613);
  not g45876 (n_20614, n28268);
  and g45877 (n28270, n_20614, n28269);
  and g45878 (n28271, n_11821, n28265);
  and g45879 (n28272, pi0619, n28161);
  not g45880 (n_20615, n28272);
  and g45881 (n28273, n_11405, n_20615);
  not g45882 (n_20616, n28271);
  and g45883 (n28274, n_20616, n28273);
  not g45884 (n_20617, n28270);
  not g45885 (n_20618, n28274);
  and g45886 (n28275, n_20617, n_20618);
  not g45887 (n_20619, n28275);
  and g45888 (n28276, pi0789, n_20619);
  not g45889 (n_20620, n28266);
  not g45890 (n_20621, n28276);
  and g45891 (n28277, n_20620, n_20621);
  and g45892 (n28278, n_12524, n28277);
  and g45893 (n28279, n17969, n28161);
  not g45894 (n_20622, n28278);
  not g45895 (n_20623, n28279);
  and g45896 (n28280, n_20622, n_20623);
  not g45897 (n_20624, n28280);
  and g45898 (n28281, n_12368, n_20624);
  and g45899 (n28282, n17779, n28161);
  not g45900 (n_20625, n28281);
  not g45901 (n_20626, n28282);
  and g45902 (n28283, n_20625, n_20626);
  not g45903 (n_20627, n28283);
  and g45904 (n28284, n_12392, n_20627);
  and g45905 (n28285, n17804, n28161);
  not g45906 (n_20628, n28284);
  not g45907 (n_20629, n28285);
  and g45908 (n28286, n_20628, n_20629);
  not g45909 (n_20630, n28286);
  and g45910 (n28287, pi0644, n_20630);
  and g45911 (n28288, n_11819, n28161);
  not g45912 (n_20631, n28288);
  and g45913 (n28289, n_12395, n_20631);
  not g45914 (n_20632, n28287);
  and g45915 (n28290, n_20632, n28289);
  not g45916 (n_20633, n28290);
  and g45917 (n28291, pi1160, n_20633);
  not g45918 (n_20634, n28223);
  and g45919 (n28292, n_20634, n28291);
  and g45920 (n28293, pi0644, n_20574);
  not g45921 (n_20635, n28293);
  and g45922 (n28294, n_12395, n_20635);
  and g45923 (n28295, n_11819, n_20630);
  and g45924 (n28296, pi0644, n28161);
  not g45925 (n_20636, n28296);
  and g45926 (n28297, pi0715, n_20636);
  not g45927 (n_20637, n28295);
  and g45928 (n28298, n_20637, n28297);
  not g45929 (n_20638, n28298);
  and g45930 (n28299, n_12405, n_20638);
  not g45931 (n_20639, n28294);
  and g45932 (n28300, n_20639, n28299);
  not g45933 (n_20640, n28292);
  not g45934 (n_20641, n28300);
  and g45935 (n28301, n_20640, n_20641);
  not g45936 (n_20642, n28301);
  and g45937 (n28302, pi0790, n_20642);
  and g45938 (n28303, n_12354, n28202);
  and g45939 (n28304, n_14557, n28280);
  and g45940 (n28305, pi0629, n28206);
  not g45941 (n_20643, n28303);
  not g45942 (n_20644, n28305);
  and g45943 (n28306, n_20643, n_20644);
  not g45944 (n_20645, n28304);
  and g45945 (n28307, n_20645, n28306);
  not g45946 (n_20646, n28307);
  and g45947 (n28308, pi0792, n_20646);
  and g45948 (n28309, pi0609, n28186);
  and g45949 (n28310, pi0184, n_12240);
  and g45950 (n28311, n_7617, n_12230);
  not g45951 (n_20647, n28310);
  and g45952 (n28312, pi0777, n_20647);
  not g45953 (n_20648, n28311);
  and g45954 (n28313, n_20648, n28312);
  and g45955 (n28314, n_7617, n17629);
  and g45956 (n28315, pi0184, n17631);
  not g45957 (n_20649, n28315);
  and g45958 (n28316, n_15730, n_20649);
  not g45959 (n_20650, n28314);
  and g45960 (n28317, n_20650, n28316);
  not g45961 (n_20651, n28313);
  not g45962 (n_20652, n28317);
  and g45963 (n28318, n_20651, n_20652);
  not g45964 (n_20653, n28318);
  and g45965 (n28319, n_162, n_20653);
  and g45966 (n28320, pi0184, n17605);
  and g45967 (n28321, n_7617, n_12180);
  not g45968 (n_20654, n28321);
  and g45969 (n28322, n_15730, n_20654);
  not g45970 (n_20655, n28320);
  and g45971 (n28323, n_20655, n28322);
  and g45972 (n28324, n_7617, n17404);
  and g45973 (n28325, pi0184, n17485);
  not g45974 (n_20656, n28325);
  and g45975 (n28326, pi0777, n_20656);
  not g45976 (n_20657, n28324);
  and g45977 (n28327, n_20657, n28326);
  not g45978 (n_20658, n28323);
  and g45979 (n28328, pi0039, n_20658);
  not g45980 (n_20659, n28327);
  and g45981 (n28329, n_20659, n28328);
  not g45982 (n_20660, n28319);
  and g45983 (n28330, n_161, n_20660);
  not g45984 (n_20661, n28329);
  and g45985 (n28331, n_20661, n28330);
  and g45986 (n28332, n_15730, n_12250);
  not g45987 (n_20662, n28332);
  and g45988 (n28333, n19471, n_20662);
  not g45989 (n_20663, n28333);
  and g45990 (n28334, n_7617, n_20663);
  and g45991 (n28335, n_12120, n_20388);
  not g45992 (n_20664, n28335);
  and g45993 (n28336, pi0184, n_20664);
  and g45994 (n28337, n6284, n28336);
  not g45995 (n_20665, n28337);
  and g45996 (n28338, pi0038, n_20665);
  not g45997 (n_20666, n28334);
  and g45998 (n28339, n_20666, n28338);
  not g45999 (n_20667, n28339);
  and g46000 (n28340, n_15732, n_20667);
  not g46001 (n_20668, n28331);
  and g46002 (n28341, n_20668, n28340);
  not g46003 (n_20669, n28236);
  and g46004 (n28342, pi0737, n_20669);
  not g46005 (n_20670, n28341);
  and g46006 (n28343, n2571, n_20670);
  not g46007 (n_20671, n28342);
  and g46008 (n28344, n_20671, n28343);
  not g46009 (n_20672, n28344);
  and g46010 (n28345, n_20585, n_20672);
  and g46011 (n28346, n_11753, n28345);
  and g46012 (n28347, pi0625, n28238);
  not g46013 (n_20673, n28347);
  and g46014 (n28348, n_11757, n_20673);
  not g46015 (n_20674, n28346);
  and g46016 (n28349, n_20674, n28348);
  and g46017 (n28350, n_11823, n_20540);
  not g46018 (n_20675, n28349);
  and g46019 (n28351, n_20675, n28350);
  and g46020 (n28352, n_11753, n28238);
  and g46021 (n28353, pi0625, n28345);
  not g46022 (n_20676, n28352);
  and g46023 (n28354, pi1153, n_20676);
  not g46024 (n_20677, n28353);
  and g46025 (n28355, n_20677, n28354);
  and g46026 (n28356, pi0608, n_20541);
  not g46027 (n_20678, n28355);
  and g46028 (n28357, n_20678, n28356);
  not g46029 (n_20679, n28351);
  not g46030 (n_20680, n28357);
  and g46031 (n28358, n_20679, n_20680);
  not g46032 (n_20681, n28358);
  and g46033 (n28359, pi0778, n_20681);
  and g46034 (n28360, n_11749, n28345);
  not g46035 (n_20682, n28359);
  not g46036 (n_20683, n28360);
  and g46037 (n28361, n_20682, n_20683);
  not g46038 (n_20684, n28361);
  and g46039 (n28362, n_11971, n_20684);
  not g46040 (n_20685, n28309);
  and g46041 (n28363, n_11768, n_20685);
  not g46042 (n_20686, n28362);
  and g46043 (n28364, n_20686, n28363);
  and g46044 (n28365, n_11767, n_20597);
  not g46045 (n_20687, n28364);
  and g46046 (n28366, n_20687, n28365);
  and g46047 (n28367, n_11971, n28186);
  and g46048 (n28368, pi0609, n_20684);
  not g46049 (n_20688, n28367);
  and g46050 (n28369, pi1155, n_20688);
  not g46051 (n_20689, n28368);
  and g46052 (n28370, n_20689, n28369);
  and g46053 (n28371, pi0660, n_20598);
  not g46054 (n_20690, n28370);
  and g46055 (n28372, n_20690, n28371);
  not g46056 (n_20691, n28366);
  not g46057 (n_20692, n28372);
  and g46058 (n28373, n_20691, n_20692);
  not g46059 (n_20693, n28373);
  and g46060 (n28374, pi0785, n_20693);
  and g46061 (n28375, n_11964, n_20684);
  not g46062 (n_20694, n28374);
  not g46063 (n_20695, n28375);
  and g46064 (n28376, n_20694, n_20695);
  not g46065 (n_20696, n28376);
  and g46066 (n28377, n_11984, n_20696);
  and g46067 (n28378, pi0618, n28189);
  not g46068 (n_20697, n28378);
  and g46069 (n28379, n_11413, n_20697);
  not g46070 (n_20698, n28377);
  and g46071 (n28380, n_20698, n28379);
  and g46072 (n28381, n_11412, n_20607);
  not g46073 (n_20699, n28380);
  and g46074 (n28382, n_20699, n28381);
  and g46075 (n28383, n_11984, n28189);
  and g46076 (n28384, pi0618, n_20696);
  not g46077 (n_20700, n28383);
  and g46078 (n28385, pi1154, n_20700);
  not g46079 (n_20701, n28384);
  and g46080 (n28386, n_20701, n28385);
  and g46081 (n28387, pi0627, n_20608);
  not g46082 (n_20702, n28386);
  and g46083 (n28388, n_20702, n28387);
  not g46084 (n_20703, n28382);
  not g46085 (n_20704, n28388);
  and g46086 (n28389, n_20703, n_20704);
  not g46087 (n_20705, n28389);
  and g46088 (n28390, pi0781, n_20705);
  and g46089 (n28391, n_11981, n_20696);
  not g46090 (n_20706, n28390);
  not g46091 (n_20707, n28391);
  and g46092 (n28392, n_20706, n_20707);
  and g46093 (n28393, n_12315, n28392);
  not g46094 (n_20708, n28192);
  and g46095 (n28394, pi0619, n_20708);
  not g46096 (n_20709, n28392);
  and g46097 (n28395, n_11821, n_20709);
  not g46098 (n_20710, n28394);
  and g46099 (n28396, n_11405, n_20710);
  not g46100 (n_20711, n28395);
  and g46101 (n28397, n_20711, n28396);
  and g46102 (n28398, n_11403, n_20617);
  not g46103 (n_20712, n28397);
  and g46104 (n28399, n_20712, n28398);
  and g46105 (n28400, n_11821, n_20708);
  and g46106 (n28401, pi0619, n_20709);
  not g46107 (n_20713, n28400);
  and g46108 (n28402, pi1159, n_20713);
  not g46109 (n_20714, n28401);
  and g46110 (n28403, n_20714, n28402);
  and g46111 (n28404, pi0648, n_20618);
  not g46112 (n_20715, n28403);
  and g46113 (n28405, n_20715, n28404);
  not g46114 (n_20716, n28399);
  and g46115 (n28406, pi0789, n_20716);
  not g46116 (n_20717, n28405);
  and g46117 (n28407, n_20717, n28406);
  not g46118 (n_20718, n28393);
  and g46119 (n28408, n17970, n_20718);
  not g46120 (n_20719, n28407);
  and g46121 (n28409, n_20719, n28408);
  and g46122 (n28410, n17871, n28194);
  not g46123 (n_20720, n28277);
  and g46124 (n28411, n_12320, n_20720);
  and g46125 (n28412, pi0626, n_20524);
  not g46126 (n_20721, n28412);
  and g46127 (n28413, n16629, n_20721);
  not g46128 (n_20722, n28411);
  and g46129 (n28414, n_20722, n28413);
  and g46130 (n28415, pi0626, n_20720);
  and g46131 (n28416, n_12320, n_20524);
  not g46132 (n_20723, n28416);
  and g46133 (n28417, n16628, n_20723);
  not g46134 (n_20724, n28415);
  and g46135 (n28418, n_20724, n28417);
  not g46136 (n_20725, n28410);
  not g46137 (n_20726, n28414);
  and g46138 (n28419, n_20725, n_20726);
  not g46139 (n_20727, n28418);
  and g46140 (n28420, n_20727, n28419);
  not g46141 (n_20728, n28420);
  and g46142 (n28421, pi0788, n_20728);
  not g46143 (n_20729, n28421);
  and g46144 (n28422, n_14638, n_20729);
  not g46145 (n_20730, n28409);
  and g46146 (n28423, n_20730, n28422);
  not g46147 (n_20731, n28308);
  not g46148 (n_20732, n28423);
  and g46149 (n28424, n_20731, n_20732);
  not g46150 (n_20733, n28424);
  and g46151 (n28425, n_14387, n_20733);
  not g46152 (n_20734, n28212);
  and g46153 (n28426, n17802, n_20734);
  and g46154 (n28427, n_14548, n28283);
  not g46155 (n_20735, n28216);
  and g46156 (n28428, n17801, n_20735);
  not g46157 (n_20736, n28426);
  not g46158 (n_20737, n28428);
  and g46159 (n28429, n_20736, n_20737);
  not g46160 (n_20738, n28427);
  and g46161 (n28430, n_20738, n28429);
  not g46162 (n_20739, n28430);
  and g46163 (n28431, pi0787, n_20739);
  and g46164 (n28432, n_11819, n28299);
  and g46165 (n28433, pi0644, n28291);
  not g46166 (n_20740, n28432);
  and g46167 (n28434, pi0790, n_20740);
  not g46168 (n_20741, n28433);
  and g46169 (n28435, n_20741, n28434);
  not g46170 (n_20742, n28425);
  not g46171 (n_20743, n28431);
  and g46172 (n28436, n_20742, n_20743);
  not g46173 (n_20744, n28435);
  and g46174 (n28437, n_20744, n28436);
  not g46175 (n_20745, n28302);
  not g46176 (n_20746, n28437);
  and g46177 (n28438, n_20745, n_20746);
  not g46178 (n_20747, n28438);
  and g46179 (n28439, n_4226, n_20747);
  not g46180 (n_20748, n28160);
  and g46181 (n28440, n_12415, n_20748);
  not g46182 (n_20749, n28439);
  and g46183 (n28441, n_20749, n28440);
  not g46184 (n_20750, n28159);
  not g46185 (n_20751, n28441);
  and g46186 (po0341, n_20750, n_20751);
  and g46187 (n28443, n_9132, n_12418);
  and g46188 (n28444, n_15110, n16645);
  not g46189 (n_20752, n28443);
  not g46190 (n_20753, n28444);
  and g46191 (n28445, n_20752, n_20753);
  not g46192 (n_20754, n28445);
  and g46193 (n28446, n_11749, n_20754);
  and g46194 (n28447, n_11753, n28444);
  not g46195 (n_20755, n28447);
  and g46196 (n28448, n_20754, n_20755);
  not g46197 (n_20756, n28448);
  and g46198 (n28449, pi1153, n_20756);
  and g46199 (n28450, n_11757, n_20752);
  and g46200 (n28451, n_20755, n28450);
  not g46201 (n_20757, n28451);
  and g46202 (n28452, pi0778, n_20757);
  not g46203 (n_20758, n28449);
  and g46204 (n28453, n_20758, n28452);
  not g46205 (n_20759, n28446);
  not g46206 (n_20760, n28453);
  and g46207 (n28454, n_20759, n_20760);
  not g46208 (n_20761, n28454);
  and g46209 (n28455, n_12429, n_20761);
  and g46210 (n28456, n_12430, n28455);
  and g46211 (n28457, n_12431, n28456);
  and g46212 (n28458, n_12432, n28457);
  and g46213 (n28459, n_12436, n28458);
  and g46214 (n28460, n_11806, n28459);
  and g46215 (n28461, pi0647, n28443);
  not g46216 (n_20762, n28461);
  and g46217 (n28462, n_11810, n_20762);
  not g46218 (n_20763, n28460);
  and g46219 (n28463, n_20763, n28462);
  and g46220 (n28464, pi0630, n28463);
  and g46221 (n28465, n_15080, n17244);
  not g46222 (n_20764, n28465);
  and g46223 (n28466, n_20752, n_20764);
  not g46224 (n_20765, n28466);
  and g46225 (n28467, n_12448, n_20765);
  not g46226 (n_20766, n28467);
  and g46227 (n28468, n_11964, n_20766);
  and g46228 (n28469, n17296, n28465);
  not g46229 (n_20767, n28469);
  and g46230 (n28470, n28467, n_20767);
  not g46231 (n_20768, n28470);
  and g46232 (n28471, pi1155, n_20768);
  and g46233 (n28472, n_11768, n_20752);
  and g46234 (n28473, n_20767, n28472);
  not g46235 (n_20769, n28471);
  not g46236 (n_20770, n28473);
  and g46237 (n28474, n_20769, n_20770);
  not g46238 (n_20771, n28474);
  and g46239 (n28475, pi0785, n_20771);
  not g46240 (n_20772, n28468);
  not g46241 (n_20773, n28475);
  and g46242 (n28476, n_20772, n_20773);
  not g46243 (n_20774, n28476);
  and g46244 (n28477, n_11981, n_20774);
  and g46245 (n28478, n_12461, n28476);
  not g46246 (n_20775, n28478);
  and g46247 (n28479, pi1154, n_20775);
  and g46248 (n28480, n_12463, n28476);
  not g46249 (n_20776, n28480);
  and g46250 (n28481, n_11413, n_20776);
  not g46251 (n_20777, n28479);
  not g46252 (n_20778, n28481);
  and g46253 (n28482, n_20777, n_20778);
  not g46254 (n_20779, n28482);
  and g46255 (n28483, pi0781, n_20779);
  not g46256 (n_20780, n28477);
  not g46257 (n_20781, n28483);
  and g46258 (n28484, n_20780, n_20781);
  not g46259 (n_20782, n28484);
  and g46260 (n28485, n_12315, n_20782);
  and g46261 (n28486, n_16503, n28484);
  not g46262 (n_20783, n28486);
  and g46263 (n28487, pi1159, n_20783);
  and g46264 (n28488, n_16505, n28484);
  not g46265 (n_20784, n28488);
  and g46266 (n28489, n_11405, n_20784);
  not g46267 (n_20785, n28487);
  not g46268 (n_20786, n28489);
  and g46269 (n28490, n_20785, n_20786);
  not g46270 (n_20787, n28490);
  and g46271 (n28491, pi0789, n_20787);
  not g46272 (n_20788, n28485);
  not g46273 (n_20789, n28491);
  and g46274 (n28492, n_20788, n_20789);
  and g46275 (n28493, n_12524, n28492);
  and g46276 (n28494, n17969, n28443);
  not g46277 (n_20790, n28493);
  not g46278 (n_20791, n28494);
  and g46279 (n28495, n_20790, n_20791);
  not g46280 (n_20792, n28495);
  and g46281 (n28496, n_12368, n_20792);
  and g46282 (n28497, n17779, n28443);
  not g46283 (n_20793, n28496);
  not g46284 (n_20794, n28497);
  and g46285 (n28498, n_20793, n_20794);
  and g46286 (n28499, n_14548, n28498);
  not g46287 (n_20795, n28459);
  and g46288 (n28500, pi0647, n_20795);
  and g46289 (n28501, n_11806, n_20752);
  not g46290 (n_20796, n28500);
  not g46291 (n_20797, n28501);
  and g46292 (n28502, n_20796, n_20797);
  not g46293 (n_20798, n28502);
  and g46294 (n28503, n17801, n_20798);
  not g46295 (n_20799, n28464);
  not g46296 (n_20800, n28503);
  and g46297 (n28504, n_20799, n_20800);
  not g46298 (n_20801, n28499);
  and g46299 (n28505, n_20801, n28504);
  not g46300 (n_20802, n28505);
  and g46301 (n28506, pi0787, n_20802);
  and g46302 (n28507, n17871, n28457);
  not g46303 (n_20803, n28492);
  and g46304 (n28508, n_12320, n_20803);
  and g46305 (n28509, pi0626, n_20752);
  not g46306 (n_20804, n28509);
  and g46307 (n28510, n16629, n_20804);
  not g46308 (n_20805, n28508);
  and g46309 (n28511, n_20805, n28510);
  and g46310 (n28512, pi0626, n_20803);
  and g46311 (n28513, n_12320, n_20752);
  not g46312 (n_20806, n28513);
  and g46313 (n28514, n16628, n_20806);
  not g46314 (n_20807, n28512);
  and g46315 (n28515, n_20807, n28514);
  not g46316 (n_20808, n28507);
  not g46317 (n_20809, n28511);
  and g46318 (n28516, n_20808, n_20809);
  not g46319 (n_20810, n28515);
  and g46320 (n28517, n_20810, n28516);
  not g46321 (n_20811, n28517);
  and g46322 (n28518, pi0788, n_20811);
  and g46323 (n28519, pi0618, n28455);
  and g46324 (n28520, n_11866, n_20754);
  and g46325 (n28521, pi0625, n28520);
  not g46326 (n_20812, n28520);
  and g46327 (n28522, n28466, n_20812);
  not g46328 (n_20813, n28521);
  not g46329 (n_20814, n28522);
  and g46330 (n28523, n_20813, n_20814);
  not g46331 (n_20815, n28523);
  and g46332 (n28524, n28450, n_20815);
  and g46333 (n28525, n_11823, n_20758);
  not g46334 (n_20816, n28524);
  and g46335 (n28526, n_20816, n28525);
  and g46336 (n28527, pi1153, n28466);
  and g46337 (n28528, n_20813, n28527);
  and g46338 (n28529, pi0608, n_20757);
  not g46339 (n_20817, n28528);
  and g46340 (n28530, n_20817, n28529);
  not g46341 (n_20818, n28526);
  not g46342 (n_20819, n28530);
  and g46343 (n28531, n_20818, n_20819);
  not g46344 (n_20820, n28531);
  and g46345 (n28532, pi0778, n_20820);
  and g46346 (n28533, n_11749, n_20814);
  not g46347 (n_20821, n28532);
  not g46348 (n_20822, n28533);
  and g46349 (n28534, n_20821, n_20822);
  not g46350 (n_20823, n28534);
  and g46351 (n28535, n_11971, n_20823);
  and g46352 (n28536, pi0609, n_20761);
  not g46353 (n_20824, n28536);
  and g46354 (n28537, n_11768, n_20824);
  not g46355 (n_20825, n28535);
  and g46356 (n28538, n_20825, n28537);
  and g46357 (n28539, n_11767, n_20769);
  not g46358 (n_20826, n28538);
  and g46359 (n28540, n_20826, n28539);
  and g46360 (n28541, pi0609, n_20823);
  and g46361 (n28542, n_11971, n_20761);
  not g46362 (n_20827, n28542);
  and g46363 (n28543, pi1155, n_20827);
  not g46364 (n_20828, n28541);
  and g46365 (n28544, n_20828, n28543);
  and g46366 (n28545, pi0660, n_20770);
  not g46367 (n_20829, n28544);
  and g46368 (n28546, n_20829, n28545);
  not g46369 (n_20830, n28540);
  not g46370 (n_20831, n28546);
  and g46371 (n28547, n_20830, n_20831);
  not g46372 (n_20832, n28547);
  and g46373 (n28548, pi0785, n_20832);
  and g46374 (n28549, n_11964, n_20823);
  not g46375 (n_20833, n28548);
  not g46376 (n_20834, n28549);
  and g46377 (n28550, n_20833, n_20834);
  not g46378 (n_20835, n28550);
  and g46379 (n28551, n_11984, n_20835);
  not g46380 (n_20836, n28519);
  and g46381 (n28552, n_11413, n_20836);
  not g46382 (n_20837, n28551);
  and g46383 (n28553, n_20837, n28552);
  and g46384 (n28554, n_11412, n_20777);
  not g46385 (n_20838, n28553);
  and g46386 (n28555, n_20838, n28554);
  and g46387 (n28556, n_11984, n28455);
  and g46388 (n28557, pi0618, n_20835);
  not g46389 (n_20839, n28556);
  and g46390 (n28558, pi1154, n_20839);
  not g46391 (n_20840, n28557);
  and g46392 (n28559, n_20840, n28558);
  and g46393 (n28560, pi0627, n_20778);
  not g46394 (n_20841, n28559);
  and g46395 (n28561, n_20841, n28560);
  not g46396 (n_20842, n28555);
  not g46397 (n_20843, n28561);
  and g46398 (n28562, n_20842, n_20843);
  not g46399 (n_20844, n28562);
  and g46400 (n28563, pi0781, n_20844);
  and g46401 (n28564, n_11981, n_20835);
  not g46402 (n_20845, n28563);
  not g46403 (n_20846, n28564);
  and g46404 (n28565, n_20845, n_20846);
  and g46405 (n28566, n_12315, n28565);
  not g46406 (n_20847, n28565);
  and g46407 (n28567, n_11821, n_20847);
  and g46408 (n28568, pi0619, n28456);
  not g46409 (n_20848, n28568);
  and g46410 (n28569, n_11405, n_20848);
  not g46411 (n_20849, n28567);
  and g46412 (n28570, n_20849, n28569);
  and g46413 (n28571, n_11403, n_20785);
  not g46414 (n_20850, n28570);
  and g46415 (n28572, n_20850, n28571);
  and g46416 (n28573, pi0619, n_20847);
  and g46417 (n28574, n_11821, n28456);
  not g46418 (n_20851, n28574);
  and g46419 (n28575, pi1159, n_20851);
  not g46420 (n_20852, n28573);
  and g46421 (n28576, n_20852, n28575);
  and g46422 (n28577, pi0648, n_20786);
  not g46423 (n_20853, n28576);
  and g46424 (n28578, n_20853, n28577);
  not g46425 (n_20854, n28572);
  and g46426 (n28579, pi0789, n_20854);
  not g46427 (n_20855, n28578);
  and g46428 (n28580, n_20855, n28579);
  not g46429 (n_20856, n28566);
  and g46430 (n28581, n17970, n_20856);
  not g46431 (n_20857, n28580);
  and g46432 (n28582, n_20857, n28581);
  not g46433 (n_20858, n28518);
  not g46434 (n_20859, n28582);
  and g46435 (n28583, n_20858, n_20859);
  not g46436 (n_20860, n28583);
  and g46437 (n28584, n_14638, n_20860);
  and g46438 (n28585, n17854, n_20792);
  and g46439 (n28586, n20851, n28458);
  not g46440 (n_20861, n28585);
  not g46441 (n_20862, n28586);
  and g46442 (n28587, n_20861, n_20862);
  not g46443 (n_20863, n28587);
  and g46444 (n28588, n_12354, n_20863);
  and g46445 (n28589, n20855, n28458);
  and g46446 (n28590, n17853, n_20792);
  not g46447 (n_20864, n28589);
  not g46448 (n_20865, n28590);
  and g46449 (n28591, n_20864, n_20865);
  not g46450 (n_20866, n28591);
  and g46451 (n28592, pi0629, n_20866);
  not g46452 (n_20867, n28588);
  not g46453 (n_20868, n28592);
  and g46454 (n28593, n_20867, n_20868);
  not g46455 (n_20869, n28593);
  and g46456 (n28594, pi0792, n_20869);
  not g46457 (n_20870, n28594);
  and g46458 (n28595, n_14387, n_20870);
  not g46459 (n_20871, n28584);
  and g46460 (n28596, n_20871, n28595);
  not g46461 (n_20872, n28506);
  not g46462 (n_20873, n28596);
  and g46463 (n28597, n_20872, n_20873);
  and g46464 (n28598, n_12411, n28597);
  and g46465 (n28599, n_11803, n_20795);
  and g46466 (n28600, pi1157, n_20798);
  not g46467 (n_20874, n28463);
  not g46468 (n_20875, n28600);
  and g46469 (n28601, n_20874, n_20875);
  not g46470 (n_20876, n28601);
  and g46471 (n28602, pi0787, n_20876);
  not g46472 (n_20877, n28599);
  not g46473 (n_20878, n28602);
  and g46474 (n28603, n_20877, n_20878);
  and g46475 (n28604, n_11819, n28603);
  and g46476 (n28605, pi0644, n28597);
  not g46477 (n_20879, n28604);
  and g46478 (n28606, pi0715, n_20879);
  not g46479 (n_20880, n28605);
  and g46480 (n28607, n_20880, n28606);
  not g46481 (n_20881, n28498);
  and g46482 (n28608, n_12392, n_20881);
  and g46483 (n28609, n17804, n28443);
  not g46484 (n_20882, n28608);
  not g46485 (n_20883, n28609);
  and g46486 (n28610, n_20882, n_20883);
  not g46487 (n_20884, n28610);
  and g46488 (n28611, pi0644, n_20884);
  and g46489 (n28612, n_11819, n28443);
  not g46490 (n_20885, n28612);
  and g46491 (n28613, n_12395, n_20885);
  not g46492 (n_20886, n28611);
  and g46493 (n28614, n_20886, n28613);
  not g46494 (n_20887, n28614);
  and g46495 (n28615, pi1160, n_20887);
  not g46496 (n_20888, n28607);
  and g46497 (n28616, n_20888, n28615);
  and g46498 (n28617, n_11819, n_20884);
  and g46499 (n28618, pi0644, n28443);
  not g46500 (n_20889, n28618);
  and g46501 (n28619, pi0715, n_20889);
  not g46502 (n_20890, n28617);
  and g46503 (n28620, n_20890, n28619);
  and g46504 (n28621, pi0644, n28603);
  and g46505 (n28622, n_11819, n28597);
  not g46506 (n_20891, n28621);
  and g46507 (n28623, n_12395, n_20891);
  not g46508 (n_20892, n28622);
  and g46509 (n28624, n_20892, n28623);
  not g46510 (n_20893, n28620);
  and g46511 (n28625, n_12405, n_20893);
  not g46512 (n_20894, n28624);
  and g46513 (n28626, n_20894, n28625);
  not g46514 (n_20895, n28616);
  not g46515 (n_20896, n28626);
  and g46516 (n28627, n_20895, n_20896);
  not g46517 (n_20897, n28627);
  and g46518 (n28628, pi0790, n_20897);
  not g46519 (n_20898, n28598);
  and g46520 (n28629, pi0832, n_20898);
  not g46521 (n_20899, n28628);
  and g46522 (n28630, n_20899, n28629);
  and g46523 (n28631, n_9132, po1038);
  and g46524 (n28632, n_9132, n_11751);
  not g46525 (n_20900, n28632);
  and g46526 (n28633, n16635, n_20900);
  and g46527 (n28634, n_15110, n2571);
  not g46528 (n_20901, n28634);
  and g46529 (n28635, n28632, n_20901);
  and g46530 (n28636, n_9132, n_11418);
  not g46531 (n_20902, n28636);
  and g46532 (n28637, n16647, n_20902);
  and g46533 (n28638, pi0185, n_12608);
  not g46534 (n_20903, n28638);
  and g46535 (n28639, n_161, n_20903);
  not g46536 (n_20904, n28639);
  and g46537 (n28640, n2571, n_20904);
  and g46538 (n28641, n_9132, n18072);
  not g46539 (n_20905, n28640);
  not g46540 (n_20906, n28641);
  and g46541 (n28642, n_20905, n_20906);
  not g46542 (n_20907, n28637);
  and g46543 (n28643, n_15110, n_20907);
  not g46544 (n_20908, n28642);
  and g46545 (n28644, n_20908, n28643);
  not g46546 (n_20909, n28635);
  not g46547 (n_20910, n28644);
  and g46548 (n28645, n_20909, n_20910);
  and g46549 (n28646, n_11749, n28645);
  and g46550 (n28647, n_11753, n28632);
  not g46551 (n_20911, n28645);
  and g46552 (n28648, pi0625, n_20911);
  not g46553 (n_20912, n28647);
  and g46554 (n28649, pi1153, n_20912);
  not g46555 (n_20913, n28648);
  and g46556 (n28650, n_20913, n28649);
  and g46557 (n28651, pi0625, n28632);
  and g46558 (n28652, n_11753, n_20911);
  not g46559 (n_20914, n28651);
  and g46560 (n28653, n_11757, n_20914);
  not g46561 (n_20915, n28652);
  and g46562 (n28654, n_20915, n28653);
  not g46563 (n_20916, n28650);
  not g46564 (n_20917, n28654);
  and g46565 (n28655, n_20916, n_20917);
  not g46566 (n_20918, n28655);
  and g46567 (n28656, pi0778, n_20918);
  not g46568 (n_20919, n28646);
  not g46569 (n_20920, n28656);
  and g46570 (n28657, n_20919, n_20920);
  not g46571 (n_20921, n28657);
  and g46572 (n28658, n_11773, n_20921);
  and g46573 (n28659, n17075, n_20900);
  not g46574 (n_20922, n28658);
  not g46575 (n_20923, n28659);
  and g46576 (n28660, n_20922, n_20923);
  and g46577 (n28661, n_11777, n28660);
  and g46578 (n28662, n16639, n28632);
  not g46579 (n_20924, n28661);
  not g46580 (n_20925, n28662);
  and g46581 (n28663, n_20924, n_20925);
  and g46582 (n28664, n_11780, n28663);
  not g46583 (n_20926, n28633);
  not g46584 (n_20927, n28664);
  and g46585 (n28665, n_20926, n_20927);
  and g46586 (n28666, n_11783, n28665);
  and g46587 (n28667, n16631, n28632);
  not g46588 (n_20928, n28666);
  not g46589 (n_20929, n28667);
  and g46590 (n28668, n_20928, n_20929);
  and g46591 (n28669, n_11787, n28668);
  not g46592 (n_20930, n28668);
  and g46593 (n28670, pi0628, n_20930);
  and g46594 (n28671, n_11789, n28632);
  not g46595 (n_20931, n28671);
  and g46596 (n28672, pi1156, n_20931);
  not g46597 (n_20932, n28670);
  and g46598 (n28673, n_20932, n28672);
  and g46599 (n28674, pi0628, n28632);
  and g46600 (n28675, n_11789, n_20930);
  not g46601 (n_20933, n28674);
  and g46602 (n28676, n_11794, n_20933);
  not g46603 (n_20934, n28675);
  and g46604 (n28677, n_20934, n28676);
  not g46605 (n_20935, n28673);
  not g46606 (n_20936, n28677);
  and g46607 (n28678, n_20935, n_20936);
  not g46608 (n_20937, n28678);
  and g46609 (n28679, pi0792, n_20937);
  not g46610 (n_20938, n28669);
  not g46611 (n_20939, n28679);
  and g46612 (n28680, n_20938, n_20939);
  not g46613 (n_20940, n28680);
  and g46614 (n28681, n_11806, n_20940);
  and g46615 (n28682, pi0647, n_20900);
  not g46616 (n_20941, n28681);
  not g46617 (n_20942, n28682);
  and g46618 (n28683, n_20941, n_20942);
  and g46619 (n28684, n_11810, n28683);
  and g46620 (n28685, pi0647, n_20940);
  and g46621 (n28686, n_11806, n_20900);
  not g46622 (n_20943, n28685);
  not g46623 (n_20944, n28686);
  and g46624 (n28687, n_20943, n_20944);
  and g46625 (n28688, pi1157, n28687);
  not g46626 (n_20945, n28684);
  not g46627 (n_20946, n28688);
  and g46628 (n28689, n_20945, n_20946);
  not g46629 (n_20947, n28689);
  and g46630 (n28690, pi0787, n_20947);
  and g46631 (n28691, n_11803, n28680);
  not g46632 (n_20948, n28690);
  not g46633 (n_20949, n28691);
  and g46634 (n28692, n_20948, n_20949);
  not g46635 (n_20950, n28692);
  and g46636 (n28693, n_11819, n_20950);
  not g46637 (n_20951, n28693);
  and g46638 (n28694, pi0715, n_20951);
  and g46639 (n28695, pi0185, n_11417);
  and g46640 (n28696, pi0185, pi0751);
  and g46641 (n28697, pi0751, n17046);
  and g46642 (n28698, pi0185, n17273);
  not g46643 (n_20952, n28697);
  not g46644 (n_20953, n28698);
  and g46645 (n28699, n_20952, n_20953);
  not g46646 (n_20954, n28699);
  and g46647 (n28700, pi0039, n_20954);
  and g46648 (n28701, pi0185, n_11923);
  not g46649 (n_20955, n28701);
  and g46650 (n28702, n_15086, n_20955);
  not g46651 (n_20956, n28702);
  and g46652 (n28703, n_162, n_20956);
  and g46653 (n28704, n_9132, n_15080);
  and g46654 (n28705, n17221, n28704);
  not g46662 (n_20961, n28708);
  and g46663 (n28709, n_161, n_20961);
  and g46664 (n28710, n_15080, n17280);
  and g46665 (n28711, pi0038, n_20902);
  not g46666 (n_20962, n28710);
  and g46667 (n28712, n_20962, n28711);
  not g46668 (n_20963, n28709);
  not g46669 (n_20964, n28712);
  and g46670 (n28713, n_20963, n_20964);
  not g46671 (n_20965, n28713);
  and g46672 (n28714, n2571, n_20965);
  not g46673 (n_20966, n28695);
  not g46674 (n_20967, n28714);
  and g46675 (n28715, n_20966, n_20967);
  not g46676 (n_20968, n28715);
  and g46677 (n28716, n_11960, n_20968);
  and g46678 (n28717, n17117, n_20900);
  not g46679 (n_20969, n28716);
  not g46680 (n_20970, n28717);
  and g46681 (n28718, n_20969, n_20970);
  not g46682 (n_20971, n28718);
  and g46683 (n28719, n_11964, n_20971);
  and g46684 (n28720, n_11967, n_20900);
  and g46685 (n28721, pi0609, n28716);
  not g46686 (n_20972, n28720);
  not g46687 (n_20973, n28721);
  and g46688 (n28722, n_20972, n_20973);
  not g46689 (n_20974, n28722);
  and g46690 (n28723, pi1155, n_20974);
  and g46691 (n28724, n_11972, n_20900);
  and g46692 (n28725, n_11971, n28716);
  not g46693 (n_20975, n28724);
  not g46694 (n_20976, n28725);
  and g46695 (n28726, n_20975, n_20976);
  not g46696 (n_20977, n28726);
  and g46697 (n28727, n_11768, n_20977);
  not g46698 (n_20978, n28723);
  not g46699 (n_20979, n28727);
  and g46700 (n28728, n_20978, n_20979);
  not g46701 (n_20980, n28728);
  and g46702 (n28729, pi0785, n_20980);
  not g46703 (n_20981, n28719);
  not g46704 (n_20982, n28729);
  and g46705 (n28730, n_20981, n_20982);
  not g46706 (n_20983, n28730);
  and g46707 (n28731, n_11981, n_20983);
  and g46708 (n28732, n_11984, n28632);
  and g46709 (n28733, pi0618, n28730);
  not g46710 (n_20984, n28732);
  and g46711 (n28734, pi1154, n_20984);
  not g46712 (n_20985, n28733);
  and g46713 (n28735, n_20985, n28734);
  and g46714 (n28736, n_11984, n28730);
  and g46715 (n28737, pi0618, n28632);
  not g46716 (n_20986, n28737);
  and g46717 (n28738, n_11413, n_20986);
  not g46718 (n_20987, n28736);
  and g46719 (n28739, n_20987, n28738);
  not g46720 (n_20988, n28735);
  not g46721 (n_20989, n28739);
  and g46722 (n28740, n_20988, n_20989);
  not g46723 (n_20990, n28740);
  and g46724 (n28741, pi0781, n_20990);
  not g46725 (n_20991, n28731);
  not g46726 (n_20992, n28741);
  and g46727 (n28742, n_20991, n_20992);
  not g46728 (n_20993, n28742);
  and g46729 (n28743, n_12315, n_20993);
  and g46730 (n28744, n_11821, n28632);
  and g46731 (n28745, pi0619, n28742);
  not g46732 (n_20994, n28744);
  and g46733 (n28746, pi1159, n_20994);
  not g46734 (n_20995, n28745);
  and g46735 (n28747, n_20995, n28746);
  and g46736 (n28748, n_11821, n28742);
  and g46737 (n28749, pi0619, n28632);
  not g46738 (n_20996, n28749);
  and g46739 (n28750, n_11405, n_20996);
  not g46740 (n_20997, n28748);
  and g46741 (n28751, n_20997, n28750);
  not g46742 (n_20998, n28747);
  not g46743 (n_20999, n28751);
  and g46744 (n28752, n_20998, n_20999);
  not g46745 (n_21000, n28752);
  and g46746 (n28753, pi0789, n_21000);
  not g46747 (n_21001, n28743);
  not g46748 (n_21002, n28753);
  and g46749 (n28754, n_21001, n_21002);
  and g46750 (n28755, n_12524, n28754);
  and g46751 (n28756, n17969, n28632);
  not g46752 (n_21003, n28755);
  not g46753 (n_21004, n28756);
  and g46754 (n28757, n_21003, n_21004);
  not g46755 (n_21005, n28757);
  and g46756 (n28758, n_12368, n_21005);
  and g46757 (n28759, n17779, n28632);
  not g46758 (n_21006, n28758);
  not g46759 (n_21007, n28759);
  and g46760 (n28760, n_21006, n_21007);
  not g46761 (n_21008, n28760);
  and g46762 (n28761, n_12392, n_21008);
  and g46763 (n28762, n17804, n28632);
  not g46764 (n_21009, n28761);
  not g46765 (n_21010, n28762);
  and g46766 (n28763, n_21009, n_21010);
  not g46767 (n_21011, n28763);
  and g46768 (n28764, pi0644, n_21011);
  and g46769 (n28765, n_11819, n28632);
  not g46770 (n_21012, n28765);
  and g46771 (n28766, n_12395, n_21012);
  not g46772 (n_21013, n28764);
  and g46773 (n28767, n_21013, n28766);
  not g46774 (n_21014, n28767);
  and g46775 (n28768, pi1160, n_21014);
  not g46776 (n_21015, n28694);
  and g46777 (n28769, n_21015, n28768);
  and g46778 (n28770, pi0644, n_20950);
  not g46779 (n_21016, n28770);
  and g46780 (n28771, n_12395, n_21016);
  and g46781 (n28772, n_11819, n_21011);
  and g46782 (n28773, pi0644, n28632);
  not g46783 (n_21017, n28773);
  and g46784 (n28774, pi0715, n_21017);
  not g46785 (n_21018, n28772);
  and g46786 (n28775, n_21018, n28774);
  not g46787 (n_21019, n28775);
  and g46788 (n28776, n_12405, n_21019);
  not g46789 (n_21020, n28771);
  and g46790 (n28777, n_21020, n28776);
  not g46791 (n_21021, n28769);
  not g46792 (n_21022, n28777);
  and g46793 (n28778, n_21021, n_21022);
  not g46794 (n_21023, n28778);
  and g46795 (n28779, pi0790, n_21023);
  and g46796 (n28780, n_12354, n28673);
  and g46797 (n28781, n_14557, n28757);
  and g46798 (n28782, pi0629, n28677);
  not g46799 (n_21024, n28780);
  not g46800 (n_21025, n28782);
  and g46801 (n28783, n_21024, n_21025);
  not g46802 (n_21026, n28781);
  and g46803 (n28784, n_21026, n28783);
  not g46804 (n_21027, n28784);
  and g46805 (n28785, pi0792, n_21027);
  and g46806 (n28786, pi0609, n28657);
  and g46807 (n28787, pi0185, n_12240);
  and g46808 (n28788, n_9132, n_12230);
  not g46809 (n_21028, n28787);
  and g46810 (n28789, pi0751, n_21028);
  not g46811 (n_21029, n28788);
  and g46812 (n28790, n_21029, n28789);
  and g46813 (n28791, n_9132, n17629);
  and g46814 (n28792, pi0185, n17631);
  not g46815 (n_21030, n28792);
  and g46816 (n28793, n_15080, n_21030);
  not g46817 (n_21031, n28791);
  and g46818 (n28794, n_21031, n28793);
  not g46819 (n_21032, n28790);
  not g46820 (n_21033, n28794);
  and g46821 (n28795, n_21032, n_21033);
  not g46822 (n_21034, n28795);
  and g46823 (n28796, n_162, n_21034);
  and g46824 (n28797, pi0185, n17605);
  and g46825 (n28798, n_9132, n_12180);
  not g46826 (n_21035, n28798);
  and g46827 (n28799, n_15080, n_21035);
  not g46828 (n_21036, n28797);
  and g46829 (n28800, n_21036, n28799);
  and g46830 (n28801, n_9132, n17404);
  and g46831 (n28802, pi0185, n17485);
  not g46832 (n_21037, n28802);
  and g46833 (n28803, pi0751, n_21037);
  not g46834 (n_21038, n28801);
  and g46835 (n28804, n_21038, n28803);
  not g46836 (n_21039, n28800);
  and g46837 (n28805, pi0039, n_21039);
  not g46838 (n_21040, n28804);
  and g46839 (n28806, n_21040, n28805);
  not g46840 (n_21041, n28796);
  and g46841 (n28807, n_161, n_21041);
  not g46842 (n_21042, n28806);
  and g46843 (n28808, n_21042, n28807);
  and g46844 (n28809, n_12120, n_20764);
  not g46845 (n_21043, n28809);
  and g46846 (n28810, pi0185, n_21043);
  and g46847 (n28811, n6284, n28810);
  and g46848 (n28812, n_15080, n_12250);
  not g46849 (n_21044, n28812);
  and g46850 (n28813, n19471, n_21044);
  not g46851 (n_21045, n28813);
  and g46852 (n28814, n_9132, n_21045);
  not g46853 (n_21046, n28811);
  and g46854 (n28815, pi0038, n_21046);
  not g46855 (n_21047, n28814);
  and g46856 (n28816, n_21047, n28815);
  not g46857 (n_21048, n28816);
  and g46858 (n28817, n_15110, n_21048);
  not g46859 (n_21049, n28808);
  and g46860 (n28818, n_21049, n28817);
  and g46861 (n28819, pi0701, n28713);
  not g46862 (n_21050, n28818);
  and g46863 (n28820, n2571, n_21050);
  not g46864 (n_21051, n28819);
  and g46865 (n28821, n_21051, n28820);
  not g46866 (n_21052, n28821);
  and g46867 (n28822, n_20966, n_21052);
  and g46868 (n28823, n_11753, n28822);
  and g46869 (n28824, pi0625, n28715);
  not g46870 (n_21053, n28824);
  and g46871 (n28825, n_11757, n_21053);
  not g46872 (n_21054, n28823);
  and g46873 (n28826, n_21054, n28825);
  and g46874 (n28827, n_11823, n_20916);
  not g46875 (n_21055, n28826);
  and g46876 (n28828, n_21055, n28827);
  and g46877 (n28829, n_11753, n28715);
  and g46878 (n28830, pi0625, n28822);
  not g46879 (n_21056, n28829);
  and g46880 (n28831, pi1153, n_21056);
  not g46881 (n_21057, n28830);
  and g46882 (n28832, n_21057, n28831);
  and g46883 (n28833, pi0608, n_20917);
  not g46884 (n_21058, n28832);
  and g46885 (n28834, n_21058, n28833);
  not g46886 (n_21059, n28828);
  not g46887 (n_21060, n28834);
  and g46888 (n28835, n_21059, n_21060);
  not g46889 (n_21061, n28835);
  and g46890 (n28836, pi0778, n_21061);
  and g46891 (n28837, n_11749, n28822);
  not g46892 (n_21062, n28836);
  not g46893 (n_21063, n28837);
  and g46894 (n28838, n_21062, n_21063);
  not g46895 (n_21064, n28838);
  and g46896 (n28839, n_11971, n_21064);
  not g46897 (n_21065, n28786);
  and g46898 (n28840, n_11768, n_21065);
  not g46899 (n_21066, n28839);
  and g46900 (n28841, n_21066, n28840);
  and g46901 (n28842, n_11767, n_20978);
  not g46902 (n_21067, n28841);
  and g46903 (n28843, n_21067, n28842);
  and g46904 (n28844, n_11971, n28657);
  and g46905 (n28845, pi0609, n_21064);
  not g46906 (n_21068, n28844);
  and g46907 (n28846, pi1155, n_21068);
  not g46908 (n_21069, n28845);
  and g46909 (n28847, n_21069, n28846);
  and g46910 (n28848, pi0660, n_20979);
  not g46911 (n_21070, n28847);
  and g46912 (n28849, n_21070, n28848);
  not g46913 (n_21071, n28843);
  not g46914 (n_21072, n28849);
  and g46915 (n28850, n_21071, n_21072);
  not g46916 (n_21073, n28850);
  and g46917 (n28851, pi0785, n_21073);
  and g46918 (n28852, n_11964, n_21064);
  not g46919 (n_21074, n28851);
  not g46920 (n_21075, n28852);
  and g46921 (n28853, n_21074, n_21075);
  not g46922 (n_21076, n28853);
  and g46923 (n28854, n_11984, n_21076);
  and g46924 (n28855, pi0618, n28660);
  not g46925 (n_21077, n28855);
  and g46926 (n28856, n_11413, n_21077);
  not g46927 (n_21078, n28854);
  and g46928 (n28857, n_21078, n28856);
  and g46929 (n28858, n_11412, n_20988);
  not g46930 (n_21079, n28857);
  and g46931 (n28859, n_21079, n28858);
  and g46932 (n28860, n_11984, n28660);
  and g46933 (n28861, pi0618, n_21076);
  not g46934 (n_21080, n28860);
  and g46935 (n28862, pi1154, n_21080);
  not g46936 (n_21081, n28861);
  and g46937 (n28863, n_21081, n28862);
  and g46938 (n28864, pi0627, n_20989);
  not g46939 (n_21082, n28863);
  and g46940 (n28865, n_21082, n28864);
  not g46941 (n_21083, n28859);
  not g46942 (n_21084, n28865);
  and g46943 (n28866, n_21083, n_21084);
  not g46944 (n_21085, n28866);
  and g46945 (n28867, pi0781, n_21085);
  and g46946 (n28868, n_11981, n_21076);
  not g46947 (n_21086, n28867);
  not g46948 (n_21087, n28868);
  and g46949 (n28869, n_21086, n_21087);
  and g46950 (n28870, n_12315, n28869);
  not g46951 (n_21088, n28663);
  and g46952 (n28871, pi0619, n_21088);
  not g46953 (n_21089, n28869);
  and g46954 (n28872, n_11821, n_21089);
  not g46955 (n_21090, n28871);
  and g46956 (n28873, n_11405, n_21090);
  not g46957 (n_21091, n28872);
  and g46958 (n28874, n_21091, n28873);
  and g46959 (n28875, n_11403, n_20998);
  not g46960 (n_21092, n28874);
  and g46961 (n28876, n_21092, n28875);
  and g46962 (n28877, n_11821, n_21088);
  and g46963 (n28878, pi0619, n_21089);
  not g46964 (n_21093, n28877);
  and g46965 (n28879, pi1159, n_21093);
  not g46966 (n_21094, n28878);
  and g46967 (n28880, n_21094, n28879);
  and g46968 (n28881, pi0648, n_20999);
  not g46969 (n_21095, n28880);
  and g46970 (n28882, n_21095, n28881);
  not g46971 (n_21096, n28876);
  and g46972 (n28883, pi0789, n_21096);
  not g46973 (n_21097, n28882);
  and g46974 (n28884, n_21097, n28883);
  not g46975 (n_21098, n28870);
  and g46976 (n28885, n17970, n_21098);
  not g46977 (n_21099, n28884);
  and g46978 (n28886, n_21099, n28885);
  and g46979 (n28887, n17871, n28665);
  not g46980 (n_21100, n28754);
  and g46981 (n28888, n_12320, n_21100);
  and g46982 (n28889, pi0626, n_20900);
  not g46983 (n_21101, n28889);
  and g46984 (n28890, n16629, n_21101);
  not g46985 (n_21102, n28888);
  and g46986 (n28891, n_21102, n28890);
  and g46987 (n28892, pi0626, n_21100);
  and g46988 (n28893, n_12320, n_20900);
  not g46989 (n_21103, n28893);
  and g46990 (n28894, n16628, n_21103);
  not g46991 (n_21104, n28892);
  and g46992 (n28895, n_21104, n28894);
  not g46993 (n_21105, n28887);
  not g46994 (n_21106, n28891);
  and g46995 (n28896, n_21105, n_21106);
  not g46996 (n_21107, n28895);
  and g46997 (n28897, n_21107, n28896);
  not g46998 (n_21108, n28897);
  and g46999 (n28898, pi0788, n_21108);
  not g47000 (n_21109, n28898);
  and g47001 (n28899, n_14638, n_21109);
  not g47002 (n_21110, n28886);
  and g47003 (n28900, n_21110, n28899);
  not g47004 (n_21111, n28785);
  not g47005 (n_21112, n28900);
  and g47006 (n28901, n_21111, n_21112);
  not g47007 (n_21113, n28901);
  and g47008 (n28902, n_14387, n_21113);
  not g47009 (n_21114, n28683);
  and g47010 (n28903, n17802, n_21114);
  and g47011 (n28904, n_14548, n28760);
  not g47012 (n_21115, n28687);
  and g47013 (n28905, n17801, n_21115);
  not g47014 (n_21116, n28903);
  not g47015 (n_21117, n28905);
  and g47016 (n28906, n_21116, n_21117);
  not g47017 (n_21118, n28904);
  and g47018 (n28907, n_21118, n28906);
  not g47019 (n_21119, n28907);
  and g47020 (n28908, pi0787, n_21119);
  and g47021 (n28909, n_11819, n28776);
  and g47022 (n28910, pi0644, n28768);
  not g47023 (n_21120, n28909);
  and g47024 (n28911, pi0790, n_21120);
  not g47025 (n_21121, n28910);
  and g47026 (n28912, n_21121, n28911);
  not g47027 (n_21122, n28902);
  not g47028 (n_21123, n28908);
  and g47029 (n28913, n_21122, n_21123);
  not g47030 (n_21124, n28912);
  and g47031 (n28914, n_21124, n28913);
  not g47032 (n_21125, n28779);
  not g47033 (n_21126, n28914);
  and g47034 (n28915, n_21125, n_21126);
  not g47035 (n_21127, n28915);
  and g47036 (n28916, n_4226, n_21127);
  not g47037 (n_21128, n28631);
  and g47038 (n28917, n_12415, n_21128);
  not g47039 (n_21129, n28916);
  and g47040 (n28918, n_21129, n28917);
  not g47041 (n_21130, n28630);
  not g47042 (n_21131, n28918);
  and g47043 (po0342, n_21130, n_21131);
  and g47044 (n28920, n_5726, n_11751);
  not g47045 (n_21132, n28920);
  and g47046 (n28921, n16635, n_21132);
  and g47047 (n28922, pi0186, n_11417);
  and g47048 (n28923, n_5726, n_11743);
  and g47049 (n28924, n_15798, n28923);
  and g47050 (n28925, n_5726, n_11418);
  not g47051 (n_21133, n28925);
  and g47052 (n28926, n16647, n_21133);
  and g47053 (n28927, n_5726, n18072);
  and g47054 (n28928, pi0186, n_12608);
  not g47055 (n_21134, n28928);
  and g47056 (n28929, n_161, n_21134);
  not g47057 (n_21135, n28927);
  and g47058 (n28930, n_21135, n28929);
  not g47059 (n_21136, n28926);
  and g47060 (n28931, pi0703, n_21136);
  not g47061 (n_21137, n28930);
  and g47062 (n28932, n_21137, n28931);
  not g47063 (n_21138, n28924);
  and g47064 (n28933, n2571, n_21138);
  not g47065 (n_21139, n28932);
  and g47066 (n28934, n_21139, n28933);
  not g47067 (n_21140, n28922);
  not g47068 (n_21141, n28934);
  and g47069 (n28935, n_21140, n_21141);
  not g47070 (n_21142, n28935);
  and g47071 (n28936, n_11749, n_21142);
  and g47072 (n28937, n_11753, n28920);
  and g47073 (n28938, pi0625, n28935);
  not g47074 (n_21143, n28937);
  and g47075 (n28939, pi1153, n_21143);
  not g47076 (n_21144, n28938);
  and g47077 (n28940, n_21144, n28939);
  and g47078 (n28941, n_11753, n28935);
  and g47079 (n28942, pi0625, n28920);
  not g47080 (n_21145, n28942);
  and g47081 (n28943, n_11757, n_21145);
  not g47082 (n_21146, n28941);
  and g47083 (n28944, n_21146, n28943);
  not g47084 (n_21147, n28940);
  not g47085 (n_21148, n28944);
  and g47086 (n28945, n_21147, n_21148);
  not g47087 (n_21149, n28945);
  and g47088 (n28946, pi0778, n_21149);
  not g47089 (n_21150, n28936);
  not g47090 (n_21151, n28946);
  and g47091 (n28947, n_21150, n_21151);
  not g47092 (n_21152, n28947);
  and g47093 (n28948, n_11773, n_21152);
  and g47094 (n28949, n17075, n_21132);
  not g47095 (n_21153, n28948);
  not g47096 (n_21154, n28949);
  and g47097 (n28950, n_21153, n_21154);
  and g47098 (n28951, n_11777, n28950);
  and g47099 (n28952, n16639, n28920);
  not g47100 (n_21155, n28951);
  not g47101 (n_21156, n28952);
  and g47102 (n28953, n_21155, n_21156);
  and g47103 (n28954, n_11780, n28953);
  not g47104 (n_21157, n28921);
  not g47105 (n_21158, n28954);
  and g47106 (n28955, n_21157, n_21158);
  and g47107 (n28956, n_11783, n28955);
  and g47108 (n28957, n16631, n28920);
  not g47109 (n_21159, n28956);
  not g47110 (n_21160, n28957);
  and g47111 (n28958, n_21159, n_21160);
  and g47112 (n28959, n_11787, n28958);
  and g47113 (n28960, n_11789, n28920);
  not g47114 (n_21161, n28958);
  and g47115 (n28961, pi0628, n_21161);
  not g47116 (n_21162, n28960);
  and g47117 (n28962, pi1156, n_21162);
  not g47118 (n_21163, n28961);
  and g47119 (n28963, n_21163, n28962);
  and g47120 (n28964, pi0628, n28920);
  and g47121 (n28965, n_11789, n_21161);
  not g47122 (n_21164, n28964);
  and g47123 (n28966, n_11794, n_21164);
  not g47124 (n_21165, n28965);
  and g47125 (n28967, n_21165, n28966);
  not g47126 (n_21166, n28963);
  not g47127 (n_21167, n28967);
  and g47128 (n28968, n_21166, n_21167);
  not g47129 (n_21168, n28968);
  and g47130 (n28969, pi0792, n_21168);
  not g47131 (n_21169, n28959);
  not g47132 (n_21170, n28969);
  and g47133 (n28970, n_21169, n_21170);
  not g47134 (n_21171, n28970);
  and g47135 (n28971, n_11803, n_21171);
  and g47136 (n28972, n_11806, n28920);
  and g47137 (n28973, pi0647, n28970);
  not g47138 (n_21172, n28972);
  and g47139 (n28974, pi1157, n_21172);
  not g47140 (n_21173, n28973);
  and g47141 (n28975, n_21173, n28974);
  and g47142 (n28976, n_11806, n28970);
  and g47143 (n28977, pi0647, n28920);
  not g47144 (n_21174, n28977);
  and g47145 (n28978, n_11810, n_21174);
  not g47146 (n_21175, n28976);
  and g47147 (n28979, n_21175, n28978);
  not g47148 (n_21176, n28975);
  not g47149 (n_21177, n28979);
  and g47150 (n28980, n_21176, n_21177);
  not g47151 (n_21178, n28980);
  and g47152 (n28981, pi0787, n_21178);
  not g47153 (n_21179, n28971);
  not g47154 (n_21180, n28981);
  and g47155 (n28982, n_21179, n_21180);
  and g47156 (n28983, n_11819, n28982);
  and g47157 (n28984, n_11984, n28920);
  not g47158 (n_21181, n28923);
  and g47159 (n28985, pi0752, n_21181);
  and g47160 (n28986, pi0186, n_13671);
  and g47161 (n28987, n_5726, n_15776);
  and g47162 (n28988, n19439, n28987);
  not g47163 (n_21182, n28986);
  not g47164 (n_21183, n28988);
  and g47165 (n28989, n_21182, n_21183);
  not g47166 (n_21184, n28989);
  and g47167 (n28990, n_13679, n_21184);
  not g47168 (n_21185, n28985);
  not g47169 (n_21186, n28990);
  and g47170 (n28991, n_21185, n_21186);
  not g47171 (n_21187, n28991);
  and g47172 (n28992, n2571, n_21187);
  not g47173 (n_21188, n28992);
  and g47174 (n28993, n_21140, n_21188);
  not g47175 (n_21189, n28993);
  and g47176 (n28994, n_11960, n_21189);
  and g47177 (n28995, n17117, n_21132);
  not g47178 (n_21190, n28994);
  not g47179 (n_21191, n28995);
  and g47180 (n28996, n_21190, n_21191);
  not g47181 (n_21192, n28996);
  and g47182 (n28997, n_11964, n_21192);
  and g47183 (n28998, n_11967, n_21132);
  and g47184 (n28999, pi0609, n28994);
  not g47185 (n_21193, n28998);
  not g47186 (n_21194, n28999);
  and g47187 (n29000, n_21193, n_21194);
  not g47188 (n_21195, n29000);
  and g47189 (n29001, pi1155, n_21195);
  and g47190 (n29002, n_11972, n_21132);
  and g47191 (n29003, n_11971, n28994);
  not g47192 (n_21196, n29002);
  not g47193 (n_21197, n29003);
  and g47194 (n29004, n_21196, n_21197);
  not g47195 (n_21198, n29004);
  and g47196 (n29005, n_11768, n_21198);
  not g47197 (n_21199, n29001);
  not g47198 (n_21200, n29005);
  and g47199 (n29006, n_21199, n_21200);
  not g47200 (n_21201, n29006);
  and g47201 (n29007, pi0785, n_21201);
  not g47202 (n_21202, n28997);
  not g47203 (n_21203, n29007);
  and g47204 (n29008, n_21202, n_21203);
  and g47205 (n29009, pi0618, n29008);
  not g47206 (n_21204, n28984);
  and g47207 (n29010, pi1154, n_21204);
  not g47208 (n_21205, n29009);
  and g47209 (n29011, n_21205, n29010);
  and g47210 (n29012, pi0186, n19468);
  and g47211 (n29013, n_5726, n19477);
  and g47217 (n29017, n_5726, n_13718);
  and g47218 (n29018, pi0186, n19496);
  not g47219 (n_21208, n29017);
  and g47220 (n29019, n_15776, n_21208);
  not g47221 (n_21209, n29018);
  and g47222 (n29020, n_21209, n29019);
  not g47223 (n_21210, n29020);
  and g47224 (n29021, pi0703, n_21210);
  not g47225 (n_21211, n29016);
  and g47226 (n29022, n_21211, n29021);
  and g47227 (n29023, n_15798, n28991);
  not g47228 (n_21212, n29022);
  and g47229 (n29024, n2571, n_21212);
  not g47230 (n_21213, n29023);
  and g47231 (n29025, n_21213, n29024);
  not g47232 (n_21214, n29025);
  and g47233 (n29026, n_21140, n_21214);
  and g47234 (n29027, n_11753, n29026);
  and g47235 (n29028, pi0625, n28993);
  not g47236 (n_21215, n29028);
  and g47237 (n29029, n_11757, n_21215);
  not g47238 (n_21216, n29027);
  and g47239 (n29030, n_21216, n29029);
  and g47240 (n29031, n_11823, n_21147);
  not g47241 (n_21217, n29030);
  and g47242 (n29032, n_21217, n29031);
  and g47243 (n29033, n_11753, n28993);
  and g47244 (n29034, pi0625, n29026);
  not g47245 (n_21218, n29033);
  and g47246 (n29035, pi1153, n_21218);
  not g47247 (n_21219, n29034);
  and g47248 (n29036, n_21219, n29035);
  and g47249 (n29037, pi0608, n_21148);
  not g47250 (n_21220, n29036);
  and g47251 (n29038, n_21220, n29037);
  not g47252 (n_21221, n29032);
  not g47253 (n_21222, n29038);
  and g47254 (n29039, n_21221, n_21222);
  not g47255 (n_21223, n29039);
  and g47256 (n29040, pi0778, n_21223);
  and g47257 (n29041, n_11749, n29026);
  not g47258 (n_21224, n29040);
  not g47259 (n_21225, n29041);
  and g47260 (n29042, n_21224, n_21225);
  not g47261 (n_21226, n29042);
  and g47262 (n29043, n_11971, n_21226);
  and g47263 (n29044, pi0609, n28947);
  not g47264 (n_21227, n29044);
  and g47265 (n29045, n_11768, n_21227);
  not g47266 (n_21228, n29043);
  and g47267 (n29046, n_21228, n29045);
  and g47268 (n29047, n_11767, n_21199);
  not g47269 (n_21229, n29046);
  and g47270 (n29048, n_21229, n29047);
  and g47271 (n29049, n_11971, n28947);
  and g47272 (n29050, pi0609, n_21226);
  not g47273 (n_21230, n29049);
  and g47274 (n29051, pi1155, n_21230);
  not g47275 (n_21231, n29050);
  and g47276 (n29052, n_21231, n29051);
  and g47277 (n29053, pi0660, n_21200);
  not g47278 (n_21232, n29052);
  and g47279 (n29054, n_21232, n29053);
  not g47280 (n_21233, n29048);
  not g47281 (n_21234, n29054);
  and g47282 (n29055, n_21233, n_21234);
  not g47283 (n_21235, n29055);
  and g47284 (n29056, pi0785, n_21235);
  and g47285 (n29057, n_11964, n_21226);
  not g47286 (n_21236, n29056);
  not g47287 (n_21237, n29057);
  and g47288 (n29058, n_21236, n_21237);
  not g47289 (n_21238, n29058);
  and g47290 (n29059, n_11984, n_21238);
  and g47291 (n29060, pi0618, n28950);
  not g47292 (n_21239, n29060);
  and g47293 (n29061, n_11413, n_21239);
  not g47294 (n_21240, n29059);
  and g47295 (n29062, n_21240, n29061);
  not g47296 (n_21241, n29011);
  and g47297 (n29063, n_11412, n_21241);
  not g47298 (n_21242, n29062);
  and g47299 (n29064, n_21242, n29063);
  and g47300 (n29065, n_11984, n29008);
  and g47301 (n29066, pi0618, n28920);
  not g47302 (n_21243, n29066);
  and g47303 (n29067, n_11413, n_21243);
  not g47304 (n_21244, n29065);
  and g47305 (n29068, n_21244, n29067);
  and g47306 (n29069, n_11984, n28950);
  and g47307 (n29070, pi0618, n_21238);
  not g47308 (n_21245, n29069);
  and g47309 (n29071, pi1154, n_21245);
  not g47310 (n_21246, n29070);
  and g47311 (n29072, n_21246, n29071);
  not g47312 (n_21247, n29068);
  and g47313 (n29073, pi0627, n_21247);
  not g47314 (n_21248, n29072);
  and g47315 (n29074, n_21248, n29073);
  not g47316 (n_21249, n29064);
  not g47317 (n_21250, n29074);
  and g47318 (n29075, n_21249, n_21250);
  not g47319 (n_21251, n29075);
  and g47320 (n29076, pi0781, n_21251);
  and g47321 (n29077, n_11981, n_21238);
  not g47322 (n_21252, n29076);
  not g47323 (n_21253, n29077);
  and g47324 (n29078, n_21252, n_21253);
  not g47325 (n_21254, n29078);
  and g47326 (n29079, n_11821, n_21254);
  not g47327 (n_21255, n28953);
  and g47328 (n29080, pi0619, n_21255);
  not g47329 (n_21256, n29080);
  and g47330 (n29081, n_11405, n_21256);
  not g47331 (n_21257, n29079);
  and g47332 (n29082, n_21257, n29081);
  and g47333 (n29083, n_11821, n28920);
  not g47334 (n_21258, n29008);
  and g47335 (n29084, n_11981, n_21258);
  and g47336 (n29085, n_21241, n_21247);
  not g47337 (n_21259, n29085);
  and g47338 (n29086, pi0781, n_21259);
  not g47339 (n_21260, n29084);
  not g47340 (n_21261, n29086);
  and g47341 (n29087, n_21260, n_21261);
  and g47342 (n29088, pi0619, n29087);
  not g47343 (n_21262, n29083);
  and g47344 (n29089, pi1159, n_21262);
  not g47345 (n_21263, n29088);
  and g47346 (n29090, n_21263, n29089);
  not g47347 (n_21264, n29090);
  and g47348 (n29091, n_11403, n_21264);
  not g47349 (n_21265, n29082);
  and g47350 (n29092, n_21265, n29091);
  and g47351 (n29093, pi0619, n_21254);
  and g47352 (n29094, n_11821, n_21255);
  not g47353 (n_21266, n29094);
  and g47354 (n29095, pi1159, n_21266);
  not g47355 (n_21267, n29093);
  and g47356 (n29096, n_21267, n29095);
  and g47357 (n29097, n_11821, n29087);
  and g47358 (n29098, pi0619, n28920);
  not g47359 (n_21268, n29098);
  and g47360 (n29099, n_11405, n_21268);
  not g47361 (n_21269, n29097);
  and g47362 (n29100, n_21269, n29099);
  not g47363 (n_21270, n29100);
  and g47364 (n29101, pi0648, n_21270);
  not g47365 (n_21271, n29096);
  and g47366 (n29102, n_21271, n29101);
  not g47367 (n_21272, n29092);
  not g47368 (n_21273, n29102);
  and g47369 (n29103, n_21272, n_21273);
  not g47370 (n_21274, n29103);
  and g47371 (n29104, pi0789, n_21274);
  and g47372 (n29105, n_12315, n_21254);
  not g47373 (n_21275, n29104);
  not g47374 (n_21276, n29105);
  and g47375 (n29106, n_21275, n_21276);
  and g47376 (n29107, n_12318, n29106);
  and g47377 (n29108, n_12320, n29106);
  not g47378 (n_21277, n28955);
  and g47379 (n29109, pi0626, n_21277);
  not g47380 (n_21278, n29109);
  and g47381 (n29110, n_11395, n_21278);
  not g47382 (n_21279, n29108);
  and g47383 (n29111, n_21279, n29110);
  not g47384 (n_21280, n29087);
  and g47385 (n29112, n_12315, n_21280);
  and g47386 (n29113, n_21264, n_21270);
  not g47387 (n_21281, n29113);
  and g47388 (n29114, pi0789, n_21281);
  not g47389 (n_21282, n29112);
  not g47390 (n_21283, n29114);
  and g47391 (n29115, n_21282, n_21283);
  not g47392 (n_21284, n29115);
  and g47393 (n29116, n_12320, n_21284);
  and g47394 (n29117, pi0626, n_21132);
  not g47395 (n_21285, n29117);
  and g47396 (n29118, pi0641, n_21285);
  not g47397 (n_21286, n29116);
  and g47398 (n29119, n_21286, n29118);
  not g47399 (n_21287, n29119);
  and g47400 (n29120, n_11397, n_21287);
  not g47401 (n_21288, n29111);
  and g47402 (n29121, n_21288, n29120);
  and g47403 (n29122, pi0626, n29106);
  and g47404 (n29123, n_12320, n_21277);
  not g47405 (n_21289, n29123);
  and g47406 (n29124, pi0641, n_21289);
  not g47407 (n_21290, n29122);
  and g47408 (n29125, n_21290, n29124);
  and g47409 (n29126, pi0626, n_21284);
  and g47410 (n29127, n_12320, n_21132);
  not g47411 (n_21291, n29127);
  and g47412 (n29128, n_11395, n_21291);
  not g47413 (n_21292, n29126);
  and g47414 (n29129, n_21292, n29128);
  not g47415 (n_21293, n29129);
  and g47416 (n29130, pi1158, n_21293);
  not g47417 (n_21294, n29125);
  and g47418 (n29131, n_21294, n29130);
  not g47419 (n_21295, n29121);
  not g47420 (n_21296, n29131);
  and g47421 (n29132, n_21295, n_21296);
  not g47422 (n_21297, n29132);
  and g47423 (n29133, pi0788, n_21297);
  not g47424 (n_21298, n29107);
  not g47425 (n_21299, n29133);
  and g47426 (n29134, n_21298, n_21299);
  and g47427 (n29135, n_11789, n29134);
  and g47428 (n29136, n_12524, n29115);
  and g47429 (n29137, n17969, n28920);
  not g47430 (n_21300, n29136);
  not g47431 (n_21301, n29137);
  and g47432 (n29138, n_21300, n_21301);
  not g47433 (n_21302, n29138);
  and g47434 (n29139, pi0628, n_21302);
  not g47435 (n_21303, n29139);
  and g47436 (n29140, n_11794, n_21303);
  not g47437 (n_21304, n29135);
  and g47438 (n29141, n_21304, n29140);
  and g47439 (n29142, n_12354, n_21166);
  not g47440 (n_21305, n29141);
  and g47441 (n29143, n_21305, n29142);
  and g47442 (n29144, pi0628, n29134);
  and g47443 (n29145, n_11789, n_21302);
  not g47444 (n_21306, n29145);
  and g47445 (n29146, pi1156, n_21306);
  not g47446 (n_21307, n29144);
  and g47447 (n29147, n_21307, n29146);
  and g47448 (n29148, pi0629, n_21167);
  not g47449 (n_21308, n29147);
  and g47450 (n29149, n_21308, n29148);
  not g47451 (n_21309, n29143);
  not g47452 (n_21310, n29149);
  and g47453 (n29150, n_21309, n_21310);
  not g47454 (n_21311, n29150);
  and g47455 (n29151, pi0792, n_21311);
  and g47456 (n29152, n_11787, n29134);
  not g47457 (n_21312, n29151);
  not g47458 (n_21313, n29152);
  and g47459 (n29153, n_21312, n_21313);
  not g47460 (n_21314, n29153);
  and g47461 (n29154, n_11806, n_21314);
  and g47462 (n29155, n_12368, n_21302);
  and g47463 (n29156, n17779, n28920);
  not g47464 (n_21315, n29155);
  not g47465 (n_21316, n29156);
  and g47466 (n29157, n_21315, n_21316);
  not g47467 (n_21317, n29157);
  and g47468 (n29158, pi0647, n_21317);
  not g47469 (n_21318, n29158);
  and g47470 (n29159, n_11810, n_21318);
  not g47471 (n_21319, n29154);
  and g47472 (n29160, n_21319, n29159);
  and g47473 (n29161, n_12375, n_21176);
  not g47474 (n_21320, n29160);
  and g47475 (n29162, n_21320, n29161);
  and g47476 (n29163, pi0647, n_21314);
  and g47477 (n29164, n_11806, n_21317);
  not g47478 (n_21321, n29164);
  and g47479 (n29165, pi1157, n_21321);
  not g47480 (n_21322, n29163);
  and g47481 (n29166, n_21322, n29165);
  and g47482 (n29167, pi0630, n_21177);
  not g47483 (n_21323, n29166);
  and g47484 (n29168, n_21323, n29167);
  not g47485 (n_21324, n29162);
  not g47486 (n_21325, n29168);
  and g47487 (n29169, n_21324, n_21325);
  not g47488 (n_21326, n29169);
  and g47489 (n29170, pi0787, n_21326);
  and g47490 (n29171, n_11803, n_21314);
  not g47491 (n_21327, n29170);
  not g47492 (n_21328, n29171);
  and g47493 (n29172, n_21327, n_21328);
  not g47494 (n_21329, n29172);
  and g47495 (n29173, pi0644, n_21329);
  not g47496 (n_21330, n28983);
  and g47497 (n29174, pi0715, n_21330);
  not g47498 (n_21331, n29173);
  and g47499 (n29175, n_21331, n29174);
  and g47500 (n29176, n17804, n_21132);
  and g47501 (n29177, n_12392, n29157);
  not g47502 (n_21332, n29176);
  not g47503 (n_21333, n29177);
  and g47504 (n29178, n_21332, n_21333);
  and g47505 (n29179, pi0644, n29178);
  and g47506 (n29180, n_11819, n28920);
  not g47507 (n_21334, n29180);
  and g47508 (n29181, n_12395, n_21334);
  not g47509 (n_21335, n29179);
  and g47510 (n29182, n_21335, n29181);
  not g47511 (n_21336, n29182);
  and g47512 (n29183, pi1160, n_21336);
  not g47513 (n_21337, n29175);
  and g47514 (n29184, n_21337, n29183);
  and g47515 (n29185, n_11819, n_21329);
  and g47516 (n29186, pi0644, n28982);
  not g47517 (n_21338, n29186);
  and g47518 (n29187, n_12395, n_21338);
  not g47519 (n_21339, n29185);
  and g47520 (n29188, n_21339, n29187);
  and g47521 (n29189, n_11819, n29178);
  and g47522 (n29190, pi0644, n28920);
  not g47523 (n_21340, n29190);
  and g47524 (n29191, pi0715, n_21340);
  not g47525 (n_21341, n29189);
  and g47526 (n29192, n_21341, n29191);
  not g47527 (n_21342, n29192);
  and g47528 (n29193, n_12405, n_21342);
  not g47529 (n_21343, n29188);
  and g47530 (n29194, n_21343, n29193);
  not g47531 (n_21344, n29184);
  and g47532 (n29195, pi0790, n_21344);
  not g47533 (n_21345, n29194);
  and g47534 (n29196, n_21345, n29195);
  and g47535 (n29197, n_12411, n29172);
  not g47536 (n_21346, n29197);
  and g47537 (n29198, n_4226, n_21346);
  not g47538 (n_21347, n29196);
  and g47539 (n29199, n_21347, n29198);
  and g47540 (n29200, n_5726, po1038);
  not g47541 (n_21348, n29200);
  and g47542 (n29201, n_12415, n_21348);
  not g47543 (n_21349, n29199);
  and g47544 (n29202, n_21349, n29201);
  and g47545 (n29203, n_5726, n_12418);
  and g47546 (n29204, pi0703, n16645);
  not g47547 (n_21350, n29203);
  not g47548 (n_21351, n29204);
  and g47549 (n29205, n_21350, n_21351);
  and g47550 (n29206, n_11749, n29205);
  and g47551 (n29207, n_11753, n29204);
  not g47552 (n_21352, n29205);
  not g47553 (n_21353, n29207);
  and g47554 (n29208, n_21352, n_21353);
  not g47555 (n_21354, n29208);
  and g47556 (n29209, pi1153, n_21354);
  and g47557 (n29210, n_11757, n_21350);
  and g47558 (n29211, n_21353, n29210);
  not g47559 (n_21355, n29209);
  not g47560 (n_21356, n29211);
  and g47561 (n29212, n_21355, n_21356);
  not g47562 (n_21357, n29212);
  and g47563 (n29213, pi0778, n_21357);
  not g47564 (n_21358, n29206);
  not g47565 (n_21359, n29213);
  and g47566 (n29214, n_21358, n_21359);
  and g47567 (n29215, n_12429, n29214);
  and g47568 (n29216, n_12430, n29215);
  and g47569 (n29217, n_12431, n29216);
  and g47570 (n29218, n_12432, n29217);
  and g47571 (n29219, n_12436, n29218);
  and g47572 (n29220, n_11806, n29219);
  and g47573 (n29221, pi0647, n29203);
  not g47574 (n_21360, n29221);
  and g47575 (n29222, n_11810, n_21360);
  not g47576 (n_21361, n29220);
  and g47577 (n29223, n_21361, n29222);
  and g47578 (n29224, pi0630, n29223);
  and g47579 (n29225, n_15776, n17244);
  not g47580 (n_21362, n29225);
  and g47581 (n29226, n_21350, n_21362);
  not g47582 (n_21363, n29226);
  and g47583 (n29227, n_12448, n_21363);
  not g47584 (n_21364, n29227);
  and g47585 (n29228, n_11964, n_21364);
  and g47586 (n29229, n_12451, n_21363);
  not g47587 (n_21365, n29229);
  and g47588 (n29230, pi1155, n_21365);
  and g47589 (n29231, n_12453, n29227);
  not g47590 (n_21366, n29231);
  and g47591 (n29232, n_11768, n_21366);
  not g47592 (n_21367, n29230);
  not g47593 (n_21368, n29232);
  and g47594 (n29233, n_21367, n_21368);
  not g47595 (n_21369, n29233);
  and g47596 (n29234, pi0785, n_21369);
  not g47597 (n_21370, n29228);
  not g47598 (n_21371, n29234);
  and g47599 (n29235, n_21370, n_21371);
  not g47600 (n_21372, n29235);
  and g47601 (n29236, n_11981, n_21372);
  and g47602 (n29237, n_12461, n29235);
  not g47603 (n_21373, n29237);
  and g47604 (n29238, pi1154, n_21373);
  and g47605 (n29239, n_12463, n29235);
  not g47606 (n_21374, n29239);
  and g47607 (n29240, n_11413, n_21374);
  not g47608 (n_21375, n29238);
  not g47609 (n_21376, n29240);
  and g47610 (n29241, n_21375, n_21376);
  not g47611 (n_21377, n29241);
  and g47612 (n29242, pi0781, n_21377);
  not g47613 (n_21378, n29236);
  not g47614 (n_21379, n29242);
  and g47615 (n29243, n_21378, n_21379);
  not g47616 (n_21380, n29243);
  and g47617 (n29244, n_12315, n_21380);
  and g47618 (n29245, n_11821, n29203);
  and g47619 (n29246, pi0619, n29243);
  not g47620 (n_21381, n29245);
  and g47621 (n29247, pi1159, n_21381);
  not g47622 (n_21382, n29246);
  and g47623 (n29248, n_21382, n29247);
  and g47624 (n29249, n_11821, n29243);
  and g47625 (n29250, pi0619, n29203);
  not g47626 (n_21383, n29250);
  and g47627 (n29251, n_11405, n_21383);
  not g47628 (n_21384, n29249);
  and g47629 (n29252, n_21384, n29251);
  not g47630 (n_21385, n29248);
  not g47631 (n_21386, n29252);
  and g47632 (n29253, n_21385, n_21386);
  not g47633 (n_21387, n29253);
  and g47634 (n29254, pi0789, n_21387);
  not g47635 (n_21388, n29244);
  not g47636 (n_21389, n29254);
  and g47637 (n29255, n_21388, n_21389);
  and g47638 (n29256, n_12524, n29255);
  and g47639 (n29257, n17969, n29203);
  not g47640 (n_21390, n29256);
  not g47641 (n_21391, n29257);
  and g47642 (n29258, n_21390, n_21391);
  not g47643 (n_21392, n29258);
  and g47644 (n29259, n_12368, n_21392);
  and g47645 (n29260, n17779, n29203);
  not g47646 (n_21393, n29259);
  not g47647 (n_21394, n29260);
  and g47648 (n29261, n_21393, n_21394);
  and g47649 (n29262, n_14548, n29261);
  not g47650 (n_21395, n29219);
  and g47651 (n29263, pi0647, n_21395);
  and g47652 (n29264, n_11806, n_21350);
  not g47653 (n_21396, n29263);
  not g47654 (n_21397, n29264);
  and g47655 (n29265, n_21396, n_21397);
  not g47656 (n_21398, n29265);
  and g47657 (n29266, n17801, n_21398);
  not g47658 (n_21399, n29224);
  not g47659 (n_21400, n29266);
  and g47660 (n29267, n_21399, n_21400);
  not g47661 (n_21401, n29262);
  and g47662 (n29268, n_21401, n29267);
  not g47663 (n_21402, n29268);
  and g47664 (n29269, pi0787, n_21402);
  and g47665 (n29270, n17871, n29217);
  not g47666 (n_21403, n29255);
  and g47667 (n29271, n_12320, n_21403);
  and g47668 (n29272, pi0626, n_21350);
  not g47669 (n_21404, n29272);
  and g47670 (n29273, n16629, n_21404);
  not g47671 (n_21405, n29271);
  and g47672 (n29274, n_21405, n29273);
  and g47673 (n29275, pi0626, n_21403);
  and g47674 (n29276, n_12320, n_21350);
  not g47675 (n_21406, n29276);
  and g47676 (n29277, n16628, n_21406);
  not g47677 (n_21407, n29275);
  and g47678 (n29278, n_21407, n29277);
  not g47679 (n_21408, n29270);
  not g47680 (n_21409, n29274);
  and g47681 (n29279, n_21408, n_21409);
  not g47682 (n_21410, n29278);
  and g47683 (n29280, n_21410, n29279);
  not g47684 (n_21411, n29280);
  and g47685 (n29281, pi0788, n_21411);
  and g47686 (n29282, pi0618, n29215);
  and g47687 (n29283, pi0609, n29214);
  and g47688 (n29284, n_11866, n_21352);
  and g47689 (n29285, pi0625, n29284);
  not g47690 (n_21412, n29284);
  and g47691 (n29286, n29226, n_21412);
  not g47692 (n_21413, n29285);
  not g47693 (n_21414, n29286);
  and g47694 (n29287, n_21413, n_21414);
  not g47695 (n_21415, n29287);
  and g47696 (n29288, n29210, n_21415);
  and g47697 (n29289, n_11823, n_21355);
  not g47698 (n_21416, n29288);
  and g47699 (n29290, n_21416, n29289);
  and g47700 (n29291, pi1153, n29226);
  and g47701 (n29292, n_21413, n29291);
  and g47702 (n29293, pi0608, n_21356);
  not g47703 (n_21417, n29292);
  and g47704 (n29294, n_21417, n29293);
  not g47705 (n_21418, n29290);
  not g47706 (n_21419, n29294);
  and g47707 (n29295, n_21418, n_21419);
  not g47708 (n_21420, n29295);
  and g47709 (n29296, pi0778, n_21420);
  and g47710 (n29297, n_11749, n_21414);
  not g47711 (n_21421, n29296);
  not g47712 (n_21422, n29297);
  and g47713 (n29298, n_21421, n_21422);
  not g47714 (n_21423, n29298);
  and g47715 (n29299, n_11971, n_21423);
  not g47716 (n_21424, n29283);
  and g47717 (n29300, n_11768, n_21424);
  not g47718 (n_21425, n29299);
  and g47719 (n29301, n_21425, n29300);
  and g47720 (n29302, n_11767, n_21367);
  not g47721 (n_21426, n29301);
  and g47722 (n29303, n_21426, n29302);
  and g47723 (n29304, n_11971, n29214);
  and g47724 (n29305, pi0609, n_21423);
  not g47725 (n_21427, n29304);
  and g47726 (n29306, pi1155, n_21427);
  not g47727 (n_21428, n29305);
  and g47728 (n29307, n_21428, n29306);
  and g47729 (n29308, pi0660, n_21368);
  not g47730 (n_21429, n29307);
  and g47731 (n29309, n_21429, n29308);
  not g47732 (n_21430, n29303);
  not g47733 (n_21431, n29309);
  and g47734 (n29310, n_21430, n_21431);
  not g47735 (n_21432, n29310);
  and g47736 (n29311, pi0785, n_21432);
  and g47737 (n29312, n_11964, n_21423);
  not g47738 (n_21433, n29311);
  not g47739 (n_21434, n29312);
  and g47740 (n29313, n_21433, n_21434);
  not g47741 (n_21435, n29313);
  and g47742 (n29314, n_11984, n_21435);
  not g47743 (n_21436, n29282);
  and g47744 (n29315, n_11413, n_21436);
  not g47745 (n_21437, n29314);
  and g47746 (n29316, n_21437, n29315);
  and g47747 (n29317, n_11412, n_21375);
  not g47748 (n_21438, n29316);
  and g47749 (n29318, n_21438, n29317);
  and g47750 (n29319, n_11984, n29215);
  and g47751 (n29320, pi0618, n_21435);
  not g47752 (n_21439, n29319);
  and g47753 (n29321, pi1154, n_21439);
  not g47754 (n_21440, n29320);
  and g47755 (n29322, n_21440, n29321);
  and g47756 (n29323, pi0627, n_21376);
  not g47757 (n_21441, n29322);
  and g47758 (n29324, n_21441, n29323);
  not g47759 (n_21442, n29318);
  not g47760 (n_21443, n29324);
  and g47761 (n29325, n_21442, n_21443);
  not g47762 (n_21444, n29325);
  and g47763 (n29326, pi0781, n_21444);
  and g47764 (n29327, n_11981, n_21435);
  not g47765 (n_21445, n29326);
  not g47766 (n_21446, n29327);
  and g47767 (n29328, n_21445, n_21446);
  and g47768 (n29329, n_12315, n29328);
  not g47769 (n_21447, n29328);
  and g47770 (n29330, n_11821, n_21447);
  and g47771 (n29331, pi0619, n29216);
  not g47772 (n_21448, n29331);
  and g47773 (n29332, n_11405, n_21448);
  not g47774 (n_21449, n29330);
  and g47775 (n29333, n_21449, n29332);
  and g47776 (n29334, n_11403, n_21385);
  not g47777 (n_21450, n29333);
  and g47778 (n29335, n_21450, n29334);
  and g47779 (n29336, pi0619, n_21447);
  and g47780 (n29337, n_11821, n29216);
  not g47781 (n_21451, n29337);
  and g47782 (n29338, pi1159, n_21451);
  not g47783 (n_21452, n29336);
  and g47784 (n29339, n_21452, n29338);
  and g47785 (n29340, pi0648, n_21386);
  not g47786 (n_21453, n29339);
  and g47787 (n29341, n_21453, n29340);
  not g47788 (n_21454, n29335);
  and g47789 (n29342, pi0789, n_21454);
  not g47790 (n_21455, n29341);
  and g47791 (n29343, n_21455, n29342);
  not g47792 (n_21456, n29329);
  and g47793 (n29344, n17970, n_21456);
  not g47794 (n_21457, n29343);
  and g47795 (n29345, n_21457, n29344);
  not g47796 (n_21458, n29281);
  not g47797 (n_21459, n29345);
  and g47798 (n29346, n_21458, n_21459);
  not g47799 (n_21460, n29346);
  and g47800 (n29347, n_14638, n_21460);
  and g47801 (n29348, n17854, n_21392);
  and g47802 (n29349, n20851, n29218);
  not g47803 (n_21461, n29348);
  not g47804 (n_21462, n29349);
  and g47805 (n29350, n_21461, n_21462);
  not g47806 (n_21463, n29350);
  and g47807 (n29351, n_12354, n_21463);
  and g47808 (n29352, n20855, n29218);
  and g47809 (n29353, n17853, n_21392);
  not g47810 (n_21464, n29352);
  not g47811 (n_21465, n29353);
  and g47812 (n29354, n_21464, n_21465);
  not g47813 (n_21466, n29354);
  and g47814 (n29355, pi0629, n_21466);
  not g47815 (n_21467, n29351);
  not g47816 (n_21468, n29355);
  and g47817 (n29356, n_21467, n_21468);
  not g47818 (n_21469, n29356);
  and g47819 (n29357, pi0792, n_21469);
  not g47820 (n_21470, n29357);
  and g47821 (n29358, n_14387, n_21470);
  not g47822 (n_21471, n29347);
  and g47823 (n29359, n_21471, n29358);
  not g47824 (n_21472, n29269);
  not g47825 (n_21473, n29359);
  and g47826 (n29360, n_21472, n_21473);
  and g47827 (n29361, n_12411, n29360);
  and g47828 (n29362, n_11803, n_21395);
  and g47829 (n29363, pi1157, n_21398);
  not g47830 (n_21474, n29223);
  not g47831 (n_21475, n29363);
  and g47832 (n29364, n_21474, n_21475);
  not g47833 (n_21476, n29364);
  and g47834 (n29365, pi0787, n_21476);
  not g47835 (n_21477, n29362);
  not g47836 (n_21478, n29365);
  and g47837 (n29366, n_21477, n_21478);
  and g47838 (n29367, n_11819, n29366);
  and g47839 (n29368, pi0644, n29360);
  not g47840 (n_21479, n29367);
  and g47841 (n29369, pi0715, n_21479);
  not g47842 (n_21480, n29368);
  and g47843 (n29370, n_21480, n29369);
  not g47844 (n_21481, n29261);
  and g47845 (n29371, n_12392, n_21481);
  and g47846 (n29372, n17804, n29203);
  not g47847 (n_21482, n29371);
  not g47848 (n_21483, n29372);
  and g47849 (n29373, n_21482, n_21483);
  not g47850 (n_21484, n29373);
  and g47851 (n29374, pi0644, n_21484);
  and g47852 (n29375, n_11819, n29203);
  not g47853 (n_21485, n29375);
  and g47854 (n29376, n_12395, n_21485);
  not g47855 (n_21486, n29374);
  and g47856 (n29377, n_21486, n29376);
  not g47857 (n_21487, n29377);
  and g47858 (n29378, pi1160, n_21487);
  not g47859 (n_21488, n29370);
  and g47860 (n29379, n_21488, n29378);
  and g47861 (n29380, n_11819, n_21484);
  and g47862 (n29381, pi0644, n29203);
  not g47863 (n_21489, n29381);
  and g47864 (n29382, pi0715, n_21489);
  not g47865 (n_21490, n29380);
  and g47866 (n29383, n_21490, n29382);
  and g47867 (n29384, pi0644, n29366);
  and g47868 (n29385, n_11819, n29360);
  not g47869 (n_21491, n29384);
  and g47870 (n29386, n_12395, n_21491);
  not g47871 (n_21492, n29385);
  and g47872 (n29387, n_21492, n29386);
  not g47873 (n_21493, n29383);
  and g47874 (n29388, n_12405, n_21493);
  not g47875 (n_21494, n29387);
  and g47876 (n29389, n_21494, n29388);
  not g47877 (n_21495, n29379);
  not g47878 (n_21496, n29389);
  and g47879 (n29390, n_21495, n_21496);
  not g47880 (n_21497, n29390);
  and g47881 (n29391, pi0790, n_21497);
  not g47882 (n_21498, n29361);
  and g47883 (n29392, pi0832, n_21498);
  not g47884 (n_21499, n29391);
  and g47885 (n29393, n_21499, n29392);
  not g47886 (n_21500, n29202);
  not g47887 (n_21501, n29393);
  and g47888 (po0343, n_21500, n_21501);
  and g47889 (n29395, n_7627, n_11751);
  not g47890 (n_21502, n29395);
  and g47891 (n29396, n16635, n_21502);
  and g47892 (n29397, pi0187, n_11417);
  and g47893 (n29398, n_7627, n_14917);
  and g47894 (n29399, n_11743, n29398);
  and g47895 (n29400, n_7627, n_11418);
  not g47896 (n_21503, n29400);
  and g47897 (n29401, n16647, n_21503);
  and g47898 (n29402, n_7627, n18072);
  and g47899 (n29403, pi0187, n_12608);
  not g47900 (n_21504, n29403);
  and g47901 (n29404, n_161, n_21504);
  not g47902 (n_21505, n29402);
  and g47903 (n29405, n_21505, n29404);
  not g47904 (n_21506, n29401);
  and g47905 (n29406, pi0726, n_21506);
  not g47906 (n_21507, n29405);
  and g47907 (n29407, n_21507, n29406);
  not g47908 (n_21508, n29399);
  and g47909 (n29408, n2571, n_21508);
  not g47910 (n_21509, n29407);
  and g47911 (n29409, n_21509, n29408);
  not g47912 (n_21510, n29397);
  not g47913 (n_21511, n29409);
  and g47914 (n29410, n_21510, n_21511);
  not g47915 (n_21512, n29410);
  and g47916 (n29411, n_11749, n_21512);
  and g47917 (n29412, n_11753, n29395);
  and g47918 (n29413, pi0625, n29410);
  not g47919 (n_21513, n29412);
  and g47920 (n29414, pi1153, n_21513);
  not g47921 (n_21514, n29413);
  and g47922 (n29415, n_21514, n29414);
  and g47923 (n29416, n_11753, n29410);
  and g47924 (n29417, pi0625, n29395);
  not g47925 (n_21515, n29417);
  and g47926 (n29418, n_11757, n_21515);
  not g47927 (n_21516, n29416);
  and g47928 (n29419, n_21516, n29418);
  not g47929 (n_21517, n29415);
  not g47930 (n_21518, n29419);
  and g47931 (n29420, n_21517, n_21518);
  not g47932 (n_21519, n29420);
  and g47933 (n29421, pi0778, n_21519);
  not g47934 (n_21520, n29411);
  not g47935 (n_21521, n29421);
  and g47936 (n29422, n_21520, n_21521);
  not g47937 (n_21522, n29422);
  and g47938 (n29423, n_11773, n_21522);
  and g47939 (n29424, n17075, n_21502);
  not g47940 (n_21523, n29423);
  not g47941 (n_21524, n29424);
  and g47942 (n29425, n_21523, n_21524);
  and g47943 (n29426, n_11777, n29425);
  and g47944 (n29427, n16639, n29395);
  not g47945 (n_21525, n29426);
  not g47946 (n_21526, n29427);
  and g47947 (n29428, n_21525, n_21526);
  and g47948 (n29429, n_11780, n29428);
  not g47949 (n_21527, n29396);
  not g47950 (n_21528, n29429);
  and g47951 (n29430, n_21527, n_21528);
  and g47952 (n29431, n_11783, n29430);
  and g47953 (n29432, n16631, n29395);
  not g47954 (n_21529, n29431);
  not g47955 (n_21530, n29432);
  and g47956 (n29433, n_21529, n_21530);
  and g47957 (n29434, n_11787, n29433);
  and g47958 (n29435, n_11789, n29395);
  not g47959 (n_21531, n29433);
  and g47960 (n29436, pi0628, n_21531);
  not g47961 (n_21532, n29435);
  and g47962 (n29437, pi1156, n_21532);
  not g47963 (n_21533, n29436);
  and g47964 (n29438, n_21533, n29437);
  and g47965 (n29439, pi0628, n29395);
  and g47966 (n29440, n_11789, n_21531);
  not g47967 (n_21534, n29439);
  and g47968 (n29441, n_11794, n_21534);
  not g47969 (n_21535, n29440);
  and g47970 (n29442, n_21535, n29441);
  not g47971 (n_21536, n29438);
  not g47972 (n_21537, n29442);
  and g47973 (n29443, n_21536, n_21537);
  not g47974 (n_21538, n29443);
  and g47975 (n29444, pi0792, n_21538);
  not g47976 (n_21539, n29434);
  not g47977 (n_21540, n29444);
  and g47978 (n29445, n_21539, n_21540);
  not g47979 (n_21541, n29445);
  and g47980 (n29446, n_11803, n_21541);
  and g47981 (n29447, n_11806, n29395);
  and g47982 (n29448, pi0647, n29445);
  not g47983 (n_21542, n29447);
  and g47984 (n29449, pi1157, n_21542);
  not g47985 (n_21543, n29448);
  and g47986 (n29450, n_21543, n29449);
  and g47987 (n29451, n_11806, n29445);
  and g47988 (n29452, pi0647, n29395);
  not g47989 (n_21544, n29452);
  and g47990 (n29453, n_11810, n_21544);
  not g47991 (n_21545, n29451);
  and g47992 (n29454, n_21545, n29453);
  not g47993 (n_21546, n29450);
  not g47994 (n_21547, n29454);
  and g47995 (n29455, n_21546, n_21547);
  not g47996 (n_21548, n29455);
  and g47997 (n29456, pi0787, n_21548);
  not g47998 (n_21549, n29446);
  not g47999 (n_21550, n29456);
  and g48000 (n29457, n_21549, n_21550);
  and g48001 (n29458, n_11819, n29457);
  and g48002 (n29459, n_11984, n29395);
  and g48003 (n29460, n_14875, n_17780);
  not g48004 (n_21551, n29460);
  and g48005 (n29461, n_14900, n_21551);
  not g48006 (n_21552, n29461);
  and g48007 (n29462, n_7627, n_21552);
  and g48008 (n29463, n_7627, n_13679);
  not g48009 (n_21553, n29463);
  and g48010 (n29464, n_14875, n_21553);
  and g48011 (n29465, n_17784, n29464);
  not g48012 (n_21554, n29462);
  not g48013 (n_21555, n29465);
  and g48014 (n29466, n_21554, n_21555);
  and g48015 (n29467, n2571, n29466);
  not g48016 (n_21556, n29467);
  and g48017 (n29468, n_21510, n_21556);
  not g48018 (n_21557, n29468);
  and g48019 (n29469, n_11960, n_21557);
  and g48020 (n29470, n17117, n_21502);
  not g48021 (n_21558, n29469);
  not g48022 (n_21559, n29470);
  and g48023 (n29471, n_21558, n_21559);
  not g48024 (n_21560, n29471);
  and g48025 (n29472, n_11964, n_21560);
  and g48026 (n29473, n_11967, n_21502);
  and g48027 (n29474, pi0609, n29469);
  not g48028 (n_21561, n29473);
  not g48029 (n_21562, n29474);
  and g48030 (n29475, n_21561, n_21562);
  not g48031 (n_21563, n29475);
  and g48032 (n29476, pi1155, n_21563);
  and g48033 (n29477, n_11972, n_21502);
  and g48034 (n29478, n_11971, n29469);
  not g48035 (n_21564, n29477);
  not g48036 (n_21565, n29478);
  and g48037 (n29479, n_21564, n_21565);
  not g48038 (n_21566, n29479);
  and g48039 (n29480, n_11768, n_21566);
  not g48040 (n_21567, n29476);
  not g48041 (n_21568, n29480);
  and g48042 (n29481, n_21567, n_21568);
  not g48043 (n_21569, n29481);
  and g48044 (n29482, pi0785, n_21569);
  not g48045 (n_21570, n29472);
  not g48046 (n_21571, n29482);
  and g48047 (n29483, n_21570, n_21571);
  and g48048 (n29484, pi0618, n29483);
  not g48049 (n_21572, n29459);
  and g48050 (n29485, pi1154, n_21572);
  not g48051 (n_21573, n29484);
  and g48052 (n29486, n_21573, n29485);
  and g48053 (n29487, pi0187, n19468);
  and g48054 (n29488, n_7627, n19477);
  and g48060 (n29492, n_7627, n_13718);
  and g48061 (n29493, pi0187, n19496);
  not g48062 (n_21576, n29492);
  and g48063 (n29494, n_14875, n_21576);
  not g48064 (n_21577, n29493);
  and g48065 (n29495, n_21577, n29494);
  not g48066 (n_21578, n29495);
  and g48067 (n29496, pi0726, n_21578);
  not g48068 (n_21579, n29491);
  and g48069 (n29497, n_21579, n29496);
  not g48070 (n_21580, n29466);
  and g48071 (n29498, n_14917, n_21580);
  not g48072 (n_21581, n29497);
  and g48073 (n29499, n2571, n_21581);
  not g48074 (n_21582, n29498);
  and g48075 (n29500, n_21582, n29499);
  not g48076 (n_21583, n29500);
  and g48077 (n29501, n_21510, n_21583);
  and g48078 (n29502, n_11753, n29501);
  and g48079 (n29503, pi0625, n29468);
  not g48080 (n_21584, n29503);
  and g48081 (n29504, n_11757, n_21584);
  not g48082 (n_21585, n29502);
  and g48083 (n29505, n_21585, n29504);
  and g48084 (n29506, n_11823, n_21517);
  not g48085 (n_21586, n29505);
  and g48086 (n29507, n_21586, n29506);
  and g48087 (n29508, n_11753, n29468);
  and g48088 (n29509, pi0625, n29501);
  not g48089 (n_21587, n29508);
  and g48090 (n29510, pi1153, n_21587);
  not g48091 (n_21588, n29509);
  and g48092 (n29511, n_21588, n29510);
  and g48093 (n29512, pi0608, n_21518);
  not g48094 (n_21589, n29511);
  and g48095 (n29513, n_21589, n29512);
  not g48096 (n_21590, n29507);
  not g48097 (n_21591, n29513);
  and g48098 (n29514, n_21590, n_21591);
  not g48099 (n_21592, n29514);
  and g48100 (n29515, pi0778, n_21592);
  and g48101 (n29516, n_11749, n29501);
  not g48102 (n_21593, n29515);
  not g48103 (n_21594, n29516);
  and g48104 (n29517, n_21593, n_21594);
  not g48105 (n_21595, n29517);
  and g48106 (n29518, n_11971, n_21595);
  and g48107 (n29519, pi0609, n29422);
  not g48108 (n_21596, n29519);
  and g48109 (n29520, n_11768, n_21596);
  not g48110 (n_21597, n29518);
  and g48111 (n29521, n_21597, n29520);
  and g48112 (n29522, n_11767, n_21567);
  not g48113 (n_21598, n29521);
  and g48114 (n29523, n_21598, n29522);
  and g48115 (n29524, n_11971, n29422);
  and g48116 (n29525, pi0609, n_21595);
  not g48117 (n_21599, n29524);
  and g48118 (n29526, pi1155, n_21599);
  not g48119 (n_21600, n29525);
  and g48120 (n29527, n_21600, n29526);
  and g48121 (n29528, pi0660, n_21568);
  not g48122 (n_21601, n29527);
  and g48123 (n29529, n_21601, n29528);
  not g48124 (n_21602, n29523);
  not g48125 (n_21603, n29529);
  and g48126 (n29530, n_21602, n_21603);
  not g48127 (n_21604, n29530);
  and g48128 (n29531, pi0785, n_21604);
  and g48129 (n29532, n_11964, n_21595);
  not g48130 (n_21605, n29531);
  not g48131 (n_21606, n29532);
  and g48132 (n29533, n_21605, n_21606);
  not g48133 (n_21607, n29533);
  and g48134 (n29534, n_11984, n_21607);
  and g48135 (n29535, pi0618, n29425);
  not g48136 (n_21608, n29535);
  and g48137 (n29536, n_11413, n_21608);
  not g48138 (n_21609, n29534);
  and g48139 (n29537, n_21609, n29536);
  not g48140 (n_21610, n29486);
  and g48141 (n29538, n_11412, n_21610);
  not g48142 (n_21611, n29537);
  and g48143 (n29539, n_21611, n29538);
  and g48144 (n29540, n_11984, n29483);
  and g48145 (n29541, pi0618, n29395);
  not g48146 (n_21612, n29541);
  and g48147 (n29542, n_11413, n_21612);
  not g48148 (n_21613, n29540);
  and g48149 (n29543, n_21613, n29542);
  and g48150 (n29544, n_11984, n29425);
  and g48151 (n29545, pi0618, n_21607);
  not g48152 (n_21614, n29544);
  and g48153 (n29546, pi1154, n_21614);
  not g48154 (n_21615, n29545);
  and g48155 (n29547, n_21615, n29546);
  not g48156 (n_21616, n29543);
  and g48157 (n29548, pi0627, n_21616);
  not g48158 (n_21617, n29547);
  and g48159 (n29549, n_21617, n29548);
  not g48160 (n_21618, n29539);
  not g48161 (n_21619, n29549);
  and g48162 (n29550, n_21618, n_21619);
  not g48163 (n_21620, n29550);
  and g48164 (n29551, pi0781, n_21620);
  and g48165 (n29552, n_11981, n_21607);
  not g48166 (n_21621, n29551);
  not g48167 (n_21622, n29552);
  and g48168 (n29553, n_21621, n_21622);
  not g48169 (n_21623, n29553);
  and g48170 (n29554, n_11821, n_21623);
  not g48171 (n_21624, n29428);
  and g48172 (n29555, pi0619, n_21624);
  not g48173 (n_21625, n29555);
  and g48174 (n29556, n_11405, n_21625);
  not g48175 (n_21626, n29554);
  and g48176 (n29557, n_21626, n29556);
  and g48177 (n29558, n_11821, n29395);
  not g48178 (n_21627, n29483);
  and g48179 (n29559, n_11981, n_21627);
  and g48180 (n29560, n_21610, n_21616);
  not g48181 (n_21628, n29560);
  and g48182 (n29561, pi0781, n_21628);
  not g48183 (n_21629, n29559);
  not g48184 (n_21630, n29561);
  and g48185 (n29562, n_21629, n_21630);
  and g48186 (n29563, pi0619, n29562);
  not g48187 (n_21631, n29558);
  and g48188 (n29564, pi1159, n_21631);
  not g48189 (n_21632, n29563);
  and g48190 (n29565, n_21632, n29564);
  not g48191 (n_21633, n29565);
  and g48192 (n29566, n_11403, n_21633);
  not g48193 (n_21634, n29557);
  and g48194 (n29567, n_21634, n29566);
  and g48195 (n29568, pi0619, n_21623);
  and g48196 (n29569, n_11821, n_21624);
  not g48197 (n_21635, n29569);
  and g48198 (n29570, pi1159, n_21635);
  not g48199 (n_21636, n29568);
  and g48200 (n29571, n_21636, n29570);
  and g48201 (n29572, n_11821, n29562);
  and g48202 (n29573, pi0619, n29395);
  not g48203 (n_21637, n29573);
  and g48204 (n29574, n_11405, n_21637);
  not g48205 (n_21638, n29572);
  and g48206 (n29575, n_21638, n29574);
  not g48207 (n_21639, n29575);
  and g48208 (n29576, pi0648, n_21639);
  not g48209 (n_21640, n29571);
  and g48210 (n29577, n_21640, n29576);
  not g48211 (n_21641, n29567);
  not g48212 (n_21642, n29577);
  and g48213 (n29578, n_21641, n_21642);
  not g48214 (n_21643, n29578);
  and g48215 (n29579, pi0789, n_21643);
  and g48216 (n29580, n_12315, n_21623);
  not g48217 (n_21644, n29579);
  not g48218 (n_21645, n29580);
  and g48219 (n29581, n_21644, n_21645);
  and g48220 (n29582, n_12318, n29581);
  and g48221 (n29583, n_12320, n29581);
  not g48222 (n_21646, n29430);
  and g48223 (n29584, pi0626, n_21646);
  not g48224 (n_21647, n29584);
  and g48225 (n29585, n_11395, n_21647);
  not g48226 (n_21648, n29583);
  and g48227 (n29586, n_21648, n29585);
  not g48228 (n_21649, n29562);
  and g48229 (n29587, n_12315, n_21649);
  and g48230 (n29588, n_21633, n_21639);
  not g48231 (n_21650, n29588);
  and g48232 (n29589, pi0789, n_21650);
  not g48233 (n_21651, n29587);
  not g48234 (n_21652, n29589);
  and g48235 (n29590, n_21651, n_21652);
  not g48236 (n_21653, n29590);
  and g48237 (n29591, n_12320, n_21653);
  and g48238 (n29592, pi0626, n_21502);
  not g48239 (n_21654, n29592);
  and g48240 (n29593, pi0641, n_21654);
  not g48241 (n_21655, n29591);
  and g48242 (n29594, n_21655, n29593);
  not g48243 (n_21656, n29594);
  and g48244 (n29595, n_11397, n_21656);
  not g48245 (n_21657, n29586);
  and g48246 (n29596, n_21657, n29595);
  and g48247 (n29597, pi0626, n29581);
  and g48248 (n29598, n_12320, n_21646);
  not g48249 (n_21658, n29598);
  and g48250 (n29599, pi0641, n_21658);
  not g48251 (n_21659, n29597);
  and g48252 (n29600, n_21659, n29599);
  and g48253 (n29601, pi0626, n_21653);
  and g48254 (n29602, n_12320, n_21502);
  not g48255 (n_21660, n29602);
  and g48256 (n29603, n_11395, n_21660);
  not g48257 (n_21661, n29601);
  and g48258 (n29604, n_21661, n29603);
  not g48259 (n_21662, n29604);
  and g48260 (n29605, pi1158, n_21662);
  not g48261 (n_21663, n29600);
  and g48262 (n29606, n_21663, n29605);
  not g48263 (n_21664, n29596);
  not g48264 (n_21665, n29606);
  and g48265 (n29607, n_21664, n_21665);
  not g48266 (n_21666, n29607);
  and g48267 (n29608, pi0788, n_21666);
  not g48268 (n_21667, n29582);
  not g48269 (n_21668, n29608);
  and g48270 (n29609, n_21667, n_21668);
  and g48271 (n29610, n_11789, n29609);
  and g48272 (n29611, n_12524, n29590);
  and g48273 (n29612, n17969, n29395);
  not g48274 (n_21669, n29611);
  not g48275 (n_21670, n29612);
  and g48276 (n29613, n_21669, n_21670);
  not g48277 (n_21671, n29613);
  and g48278 (n29614, pi0628, n_21671);
  not g48279 (n_21672, n29614);
  and g48280 (n29615, n_11794, n_21672);
  not g48281 (n_21673, n29610);
  and g48282 (n29616, n_21673, n29615);
  and g48283 (n29617, n_12354, n_21536);
  not g48284 (n_21674, n29616);
  and g48285 (n29618, n_21674, n29617);
  and g48286 (n29619, pi0628, n29609);
  and g48287 (n29620, n_11789, n_21671);
  not g48288 (n_21675, n29620);
  and g48289 (n29621, pi1156, n_21675);
  not g48290 (n_21676, n29619);
  and g48291 (n29622, n_21676, n29621);
  and g48292 (n29623, pi0629, n_21537);
  not g48293 (n_21677, n29622);
  and g48294 (n29624, n_21677, n29623);
  not g48295 (n_21678, n29618);
  not g48296 (n_21679, n29624);
  and g48297 (n29625, n_21678, n_21679);
  not g48298 (n_21680, n29625);
  and g48299 (n29626, pi0792, n_21680);
  and g48300 (n29627, n_11787, n29609);
  not g48301 (n_21681, n29626);
  not g48302 (n_21682, n29627);
  and g48303 (n29628, n_21681, n_21682);
  not g48304 (n_21683, n29628);
  and g48305 (n29629, n_11806, n_21683);
  and g48306 (n29630, n_12368, n_21671);
  and g48307 (n29631, n17779, n29395);
  not g48308 (n_21684, n29630);
  not g48309 (n_21685, n29631);
  and g48310 (n29632, n_21684, n_21685);
  not g48311 (n_21686, n29632);
  and g48312 (n29633, pi0647, n_21686);
  not g48313 (n_21687, n29633);
  and g48314 (n29634, n_11810, n_21687);
  not g48315 (n_21688, n29629);
  and g48316 (n29635, n_21688, n29634);
  and g48317 (n29636, n_12375, n_21546);
  not g48318 (n_21689, n29635);
  and g48319 (n29637, n_21689, n29636);
  and g48320 (n29638, pi0647, n_21683);
  and g48321 (n29639, n_11806, n_21686);
  not g48322 (n_21690, n29639);
  and g48323 (n29640, pi1157, n_21690);
  not g48324 (n_21691, n29638);
  and g48325 (n29641, n_21691, n29640);
  and g48326 (n29642, pi0630, n_21547);
  not g48327 (n_21692, n29641);
  and g48328 (n29643, n_21692, n29642);
  not g48329 (n_21693, n29637);
  not g48330 (n_21694, n29643);
  and g48331 (n29644, n_21693, n_21694);
  not g48332 (n_21695, n29644);
  and g48333 (n29645, pi0787, n_21695);
  and g48334 (n29646, n_11803, n_21683);
  not g48335 (n_21696, n29645);
  not g48336 (n_21697, n29646);
  and g48337 (n29647, n_21696, n_21697);
  not g48338 (n_21698, n29647);
  and g48339 (n29648, pi0644, n_21698);
  not g48340 (n_21699, n29458);
  and g48341 (n29649, pi0715, n_21699);
  not g48342 (n_21700, n29648);
  and g48343 (n29650, n_21700, n29649);
  and g48344 (n29651, n17804, n_21502);
  and g48345 (n29652, n_12392, n29632);
  not g48346 (n_21701, n29651);
  not g48347 (n_21702, n29652);
  and g48348 (n29653, n_21701, n_21702);
  and g48349 (n29654, pi0644, n29653);
  and g48350 (n29655, n_11819, n29395);
  not g48351 (n_21703, n29655);
  and g48352 (n29656, n_12395, n_21703);
  not g48353 (n_21704, n29654);
  and g48354 (n29657, n_21704, n29656);
  not g48355 (n_21705, n29657);
  and g48356 (n29658, pi1160, n_21705);
  not g48357 (n_21706, n29650);
  and g48358 (n29659, n_21706, n29658);
  and g48359 (n29660, n_11819, n_21698);
  and g48360 (n29661, pi0644, n29457);
  not g48361 (n_21707, n29661);
  and g48362 (n29662, n_12395, n_21707);
  not g48363 (n_21708, n29660);
  and g48364 (n29663, n_21708, n29662);
  and g48365 (n29664, n_11819, n29653);
  and g48366 (n29665, pi0644, n29395);
  not g48367 (n_21709, n29665);
  and g48368 (n29666, pi0715, n_21709);
  not g48369 (n_21710, n29664);
  and g48370 (n29667, n_21710, n29666);
  not g48371 (n_21711, n29667);
  and g48372 (n29668, n_12405, n_21711);
  not g48373 (n_21712, n29663);
  and g48374 (n29669, n_21712, n29668);
  not g48375 (n_21713, n29659);
  and g48376 (n29670, pi0790, n_21713);
  not g48377 (n_21714, n29669);
  and g48378 (n29671, n_21714, n29670);
  and g48379 (n29672, n_12411, n29647);
  not g48380 (n_21715, n29672);
  and g48381 (n29673, n_4226, n_21715);
  not g48382 (n_21716, n29671);
  and g48383 (n29674, n_21716, n29673);
  and g48384 (n29675, n_7627, po1038);
  not g48385 (n_21717, n29675);
  and g48386 (n29676, n_12415, n_21717);
  not g48387 (n_21718, n29674);
  and g48388 (n29677, n_21718, n29676);
  and g48389 (n29678, n_7627, n_12418);
  and g48390 (n29679, pi0726, n16645);
  not g48391 (n_21719, n29678);
  not g48392 (n_21720, n29679);
  and g48393 (n29680, n_21719, n_21720);
  and g48394 (n29681, n_11749, n29680);
  and g48395 (n29682, n_11753, n29679);
  not g48396 (n_21721, n29680);
  not g48397 (n_21722, n29682);
  and g48398 (n29683, n_21721, n_21722);
  not g48399 (n_21723, n29683);
  and g48400 (n29684, pi1153, n_21723);
  and g48401 (n29685, n_11757, n_21719);
  and g48402 (n29686, n_21722, n29685);
  not g48403 (n_21724, n29684);
  not g48404 (n_21725, n29686);
  and g48405 (n29687, n_21724, n_21725);
  not g48406 (n_21726, n29687);
  and g48407 (n29688, pi0778, n_21726);
  not g48408 (n_21727, n29681);
  not g48409 (n_21728, n29688);
  and g48410 (n29689, n_21727, n_21728);
  and g48411 (n29690, n_12429, n29689);
  and g48412 (n29691, n_12430, n29690);
  and g48413 (n29692, n_12431, n29691);
  and g48414 (n29693, n_12432, n29692);
  and g48415 (n29694, n_12436, n29693);
  and g48416 (n29695, n_11806, n29694);
  and g48417 (n29696, pi0647, n29678);
  not g48418 (n_21729, n29696);
  and g48419 (n29697, n_11810, n_21729);
  not g48420 (n_21730, n29695);
  and g48421 (n29698, n_21730, n29697);
  and g48422 (n29699, pi0630, n29698);
  and g48423 (n29700, n_14875, n17244);
  not g48424 (n_21731, n29700);
  and g48425 (n29701, n_21719, n_21731);
  not g48426 (n_21732, n29701);
  and g48427 (n29702, n_12448, n_21732);
  not g48428 (n_21733, n29702);
  and g48429 (n29703, n_11964, n_21733);
  and g48430 (n29704, n_12451, n_21732);
  not g48431 (n_21734, n29704);
  and g48432 (n29705, pi1155, n_21734);
  and g48433 (n29706, n_12453, n29702);
  not g48434 (n_21735, n29706);
  and g48435 (n29707, n_11768, n_21735);
  not g48436 (n_21736, n29705);
  not g48437 (n_21737, n29707);
  and g48438 (n29708, n_21736, n_21737);
  not g48439 (n_21738, n29708);
  and g48440 (n29709, pi0785, n_21738);
  not g48441 (n_21739, n29703);
  not g48442 (n_21740, n29709);
  and g48443 (n29710, n_21739, n_21740);
  not g48444 (n_21741, n29710);
  and g48445 (n29711, n_11981, n_21741);
  and g48446 (n29712, n_12461, n29710);
  not g48447 (n_21742, n29712);
  and g48448 (n29713, pi1154, n_21742);
  and g48449 (n29714, n_12463, n29710);
  not g48450 (n_21743, n29714);
  and g48451 (n29715, n_11413, n_21743);
  not g48452 (n_21744, n29713);
  not g48453 (n_21745, n29715);
  and g48454 (n29716, n_21744, n_21745);
  not g48455 (n_21746, n29716);
  and g48456 (n29717, pi0781, n_21746);
  not g48457 (n_21747, n29711);
  not g48458 (n_21748, n29717);
  and g48459 (n29718, n_21747, n_21748);
  not g48460 (n_21749, n29718);
  and g48461 (n29719, n_12315, n_21749);
  and g48462 (n29720, n_11821, n29678);
  and g48463 (n29721, pi0619, n29718);
  not g48464 (n_21750, n29720);
  and g48465 (n29722, pi1159, n_21750);
  not g48466 (n_21751, n29721);
  and g48467 (n29723, n_21751, n29722);
  and g48468 (n29724, n_11821, n29718);
  and g48469 (n29725, pi0619, n29678);
  not g48470 (n_21752, n29725);
  and g48471 (n29726, n_11405, n_21752);
  not g48472 (n_21753, n29724);
  and g48473 (n29727, n_21753, n29726);
  not g48474 (n_21754, n29723);
  not g48475 (n_21755, n29727);
  and g48476 (n29728, n_21754, n_21755);
  not g48477 (n_21756, n29728);
  and g48478 (n29729, pi0789, n_21756);
  not g48479 (n_21757, n29719);
  not g48480 (n_21758, n29729);
  and g48481 (n29730, n_21757, n_21758);
  and g48482 (n29731, n_12524, n29730);
  and g48483 (n29732, n17969, n29678);
  not g48484 (n_21759, n29731);
  not g48485 (n_21760, n29732);
  and g48486 (n29733, n_21759, n_21760);
  not g48487 (n_21761, n29733);
  and g48488 (n29734, n_12368, n_21761);
  and g48489 (n29735, n17779, n29678);
  not g48490 (n_21762, n29734);
  not g48491 (n_21763, n29735);
  and g48492 (n29736, n_21762, n_21763);
  and g48493 (n29737, n_14548, n29736);
  not g48494 (n_21764, n29694);
  and g48495 (n29738, pi0647, n_21764);
  and g48496 (n29739, n_11806, n_21719);
  not g48497 (n_21765, n29738);
  not g48498 (n_21766, n29739);
  and g48499 (n29740, n_21765, n_21766);
  not g48500 (n_21767, n29740);
  and g48501 (n29741, n17801, n_21767);
  not g48502 (n_21768, n29699);
  not g48503 (n_21769, n29741);
  and g48504 (n29742, n_21768, n_21769);
  not g48505 (n_21770, n29737);
  and g48506 (n29743, n_21770, n29742);
  not g48507 (n_21771, n29743);
  and g48508 (n29744, pi0787, n_21771);
  and g48509 (n29745, n17871, n29692);
  not g48510 (n_21772, n29730);
  and g48511 (n29746, n_12320, n_21772);
  and g48512 (n29747, pi0626, n_21719);
  not g48513 (n_21773, n29747);
  and g48514 (n29748, n16629, n_21773);
  not g48515 (n_21774, n29746);
  and g48516 (n29749, n_21774, n29748);
  and g48517 (n29750, pi0626, n_21772);
  and g48518 (n29751, n_12320, n_21719);
  not g48519 (n_21775, n29751);
  and g48520 (n29752, n16628, n_21775);
  not g48521 (n_21776, n29750);
  and g48522 (n29753, n_21776, n29752);
  not g48523 (n_21777, n29745);
  not g48524 (n_21778, n29749);
  and g48525 (n29754, n_21777, n_21778);
  not g48526 (n_21779, n29753);
  and g48527 (n29755, n_21779, n29754);
  not g48528 (n_21780, n29755);
  and g48529 (n29756, pi0788, n_21780);
  and g48530 (n29757, pi0618, n29690);
  and g48531 (n29758, pi0609, n29689);
  and g48532 (n29759, n_11866, n_21721);
  and g48533 (n29760, pi0625, n29759);
  not g48534 (n_21781, n29759);
  and g48535 (n29761, n29701, n_21781);
  not g48536 (n_21782, n29760);
  not g48537 (n_21783, n29761);
  and g48538 (n29762, n_21782, n_21783);
  not g48539 (n_21784, n29762);
  and g48540 (n29763, n29685, n_21784);
  and g48541 (n29764, n_11823, n_21724);
  not g48542 (n_21785, n29763);
  and g48543 (n29765, n_21785, n29764);
  and g48544 (n29766, pi1153, n29701);
  and g48545 (n29767, n_21782, n29766);
  and g48546 (n29768, pi0608, n_21725);
  not g48547 (n_21786, n29767);
  and g48548 (n29769, n_21786, n29768);
  not g48549 (n_21787, n29765);
  not g48550 (n_21788, n29769);
  and g48551 (n29770, n_21787, n_21788);
  not g48552 (n_21789, n29770);
  and g48553 (n29771, pi0778, n_21789);
  and g48554 (n29772, n_11749, n_21783);
  not g48555 (n_21790, n29771);
  not g48556 (n_21791, n29772);
  and g48557 (n29773, n_21790, n_21791);
  not g48558 (n_21792, n29773);
  and g48559 (n29774, n_11971, n_21792);
  not g48560 (n_21793, n29758);
  and g48561 (n29775, n_11768, n_21793);
  not g48562 (n_21794, n29774);
  and g48563 (n29776, n_21794, n29775);
  and g48564 (n29777, n_11767, n_21736);
  not g48565 (n_21795, n29776);
  and g48566 (n29778, n_21795, n29777);
  and g48567 (n29779, n_11971, n29689);
  and g48568 (n29780, pi0609, n_21792);
  not g48569 (n_21796, n29779);
  and g48570 (n29781, pi1155, n_21796);
  not g48571 (n_21797, n29780);
  and g48572 (n29782, n_21797, n29781);
  and g48573 (n29783, pi0660, n_21737);
  not g48574 (n_21798, n29782);
  and g48575 (n29784, n_21798, n29783);
  not g48576 (n_21799, n29778);
  not g48577 (n_21800, n29784);
  and g48578 (n29785, n_21799, n_21800);
  not g48579 (n_21801, n29785);
  and g48580 (n29786, pi0785, n_21801);
  and g48581 (n29787, n_11964, n_21792);
  not g48582 (n_21802, n29786);
  not g48583 (n_21803, n29787);
  and g48584 (n29788, n_21802, n_21803);
  not g48585 (n_21804, n29788);
  and g48586 (n29789, n_11984, n_21804);
  not g48587 (n_21805, n29757);
  and g48588 (n29790, n_11413, n_21805);
  not g48589 (n_21806, n29789);
  and g48590 (n29791, n_21806, n29790);
  and g48591 (n29792, n_11412, n_21744);
  not g48592 (n_21807, n29791);
  and g48593 (n29793, n_21807, n29792);
  and g48594 (n29794, n_11984, n29690);
  and g48595 (n29795, pi0618, n_21804);
  not g48596 (n_21808, n29794);
  and g48597 (n29796, pi1154, n_21808);
  not g48598 (n_21809, n29795);
  and g48599 (n29797, n_21809, n29796);
  and g48600 (n29798, pi0627, n_21745);
  not g48601 (n_21810, n29797);
  and g48602 (n29799, n_21810, n29798);
  not g48603 (n_21811, n29793);
  not g48604 (n_21812, n29799);
  and g48605 (n29800, n_21811, n_21812);
  not g48606 (n_21813, n29800);
  and g48607 (n29801, pi0781, n_21813);
  and g48608 (n29802, n_11981, n_21804);
  not g48609 (n_21814, n29801);
  not g48610 (n_21815, n29802);
  and g48611 (n29803, n_21814, n_21815);
  and g48612 (n29804, n_12315, n29803);
  not g48613 (n_21816, n29803);
  and g48614 (n29805, n_11821, n_21816);
  and g48615 (n29806, pi0619, n29691);
  not g48616 (n_21817, n29806);
  and g48617 (n29807, n_11405, n_21817);
  not g48618 (n_21818, n29805);
  and g48619 (n29808, n_21818, n29807);
  and g48620 (n29809, n_11403, n_21754);
  not g48621 (n_21819, n29808);
  and g48622 (n29810, n_21819, n29809);
  and g48623 (n29811, pi0619, n_21816);
  and g48624 (n29812, n_11821, n29691);
  not g48625 (n_21820, n29812);
  and g48626 (n29813, pi1159, n_21820);
  not g48627 (n_21821, n29811);
  and g48628 (n29814, n_21821, n29813);
  and g48629 (n29815, pi0648, n_21755);
  not g48630 (n_21822, n29814);
  and g48631 (n29816, n_21822, n29815);
  not g48632 (n_21823, n29810);
  and g48633 (n29817, pi0789, n_21823);
  not g48634 (n_21824, n29816);
  and g48635 (n29818, n_21824, n29817);
  not g48636 (n_21825, n29804);
  and g48637 (n29819, n17970, n_21825);
  not g48638 (n_21826, n29818);
  and g48639 (n29820, n_21826, n29819);
  not g48640 (n_21827, n29756);
  not g48641 (n_21828, n29820);
  and g48642 (n29821, n_21827, n_21828);
  not g48643 (n_21829, n29821);
  and g48644 (n29822, n_14638, n_21829);
  and g48645 (n29823, n17854, n_21761);
  and g48646 (n29824, n20851, n29693);
  not g48647 (n_21830, n29823);
  not g48648 (n_21831, n29824);
  and g48649 (n29825, n_21830, n_21831);
  not g48650 (n_21832, n29825);
  and g48651 (n29826, n_12354, n_21832);
  and g48652 (n29827, n20855, n29693);
  and g48653 (n29828, n17853, n_21761);
  not g48654 (n_21833, n29827);
  not g48655 (n_21834, n29828);
  and g48656 (n29829, n_21833, n_21834);
  not g48657 (n_21835, n29829);
  and g48658 (n29830, pi0629, n_21835);
  not g48659 (n_21836, n29826);
  not g48660 (n_21837, n29830);
  and g48661 (n29831, n_21836, n_21837);
  not g48662 (n_21838, n29831);
  and g48663 (n29832, pi0792, n_21838);
  not g48664 (n_21839, n29832);
  and g48665 (n29833, n_14387, n_21839);
  not g48666 (n_21840, n29822);
  and g48667 (n29834, n_21840, n29833);
  not g48668 (n_21841, n29744);
  not g48669 (n_21842, n29834);
  and g48670 (n29835, n_21841, n_21842);
  and g48671 (n29836, n_12411, n29835);
  and g48672 (n29837, n_11803, n_21764);
  and g48673 (n29838, pi1157, n_21767);
  not g48674 (n_21843, n29698);
  not g48675 (n_21844, n29838);
  and g48676 (n29839, n_21843, n_21844);
  not g48677 (n_21845, n29839);
  and g48678 (n29840, pi0787, n_21845);
  not g48679 (n_21846, n29837);
  not g48680 (n_21847, n29840);
  and g48681 (n29841, n_21846, n_21847);
  and g48682 (n29842, n_11819, n29841);
  and g48683 (n29843, pi0644, n29835);
  not g48684 (n_21848, n29842);
  and g48685 (n29844, pi0715, n_21848);
  not g48686 (n_21849, n29843);
  and g48687 (n29845, n_21849, n29844);
  not g48688 (n_21850, n29736);
  and g48689 (n29846, n_12392, n_21850);
  and g48690 (n29847, n17804, n29678);
  not g48691 (n_21851, n29846);
  not g48692 (n_21852, n29847);
  and g48693 (n29848, n_21851, n_21852);
  not g48694 (n_21853, n29848);
  and g48695 (n29849, pi0644, n_21853);
  and g48696 (n29850, n_11819, n29678);
  not g48697 (n_21854, n29850);
  and g48698 (n29851, n_12395, n_21854);
  not g48699 (n_21855, n29849);
  and g48700 (n29852, n_21855, n29851);
  not g48701 (n_21856, n29852);
  and g48702 (n29853, pi1160, n_21856);
  not g48703 (n_21857, n29845);
  and g48704 (n29854, n_21857, n29853);
  and g48705 (n29855, n_11819, n_21853);
  and g48706 (n29856, pi0644, n29678);
  not g48707 (n_21858, n29856);
  and g48708 (n29857, pi0715, n_21858);
  not g48709 (n_21859, n29855);
  and g48710 (n29858, n_21859, n29857);
  and g48711 (n29859, pi0644, n29841);
  and g48712 (n29860, n_11819, n29835);
  not g48713 (n_21860, n29859);
  and g48714 (n29861, n_12395, n_21860);
  not g48715 (n_21861, n29860);
  and g48716 (n29862, n_21861, n29861);
  not g48717 (n_21862, n29858);
  and g48718 (n29863, n_12405, n_21862);
  not g48719 (n_21863, n29862);
  and g48720 (n29864, n_21863, n29863);
  not g48721 (n_21864, n29854);
  not g48722 (n_21865, n29864);
  and g48723 (n29865, n_21864, n_21865);
  not g48724 (n_21866, n29865);
  and g48725 (n29866, pi0790, n_21866);
  not g48726 (n_21867, n29836);
  and g48727 (n29867, pi0832, n_21867);
  not g48728 (n_21868, n29866);
  and g48729 (n29868, n_21868, n29867);
  not g48730 (n_21869, n29677);
  not g48731 (n_21870, n29868);
  and g48732 (po0344, n_21869, n_21870);
  and g48733 (n29870, n_6272, n_11751);
  not g48734 (n_21871, n29870);
  and g48735 (n29871, n16635, n_21871);
  and g48736 (n29872, pi0188, n_11417);
  and g48737 (n29873, n_6272, n_15924);
  and g48738 (n29874, n_11743, n29873);
  and g48739 (n29875, n_6272, n_11418);
  not g48740 (n_21872, n29875);
  and g48741 (n29876, n16647, n_21872);
  and g48742 (n29877, n_6272, n18072);
  and g48743 (n29878, pi0188, n_12608);
  not g48744 (n_21873, n29878);
  and g48745 (n29879, n_161, n_21873);
  not g48746 (n_21874, n29877);
  and g48747 (n29880, n_21874, n29879);
  not g48748 (n_21875, n29876);
  and g48749 (n29881, pi0705, n_21875);
  not g48750 (n_21876, n29880);
  and g48751 (n29882, n_21876, n29881);
  not g48752 (n_21877, n29874);
  and g48753 (n29883, n2571, n_21877);
  not g48754 (n_21878, n29882);
  and g48755 (n29884, n_21878, n29883);
  not g48756 (n_21879, n29872);
  not g48757 (n_21880, n29884);
  and g48758 (n29885, n_21879, n_21880);
  not g48759 (n_21881, n29885);
  and g48760 (n29886, n_11749, n_21881);
  and g48761 (n29887, n_11753, n29870);
  and g48762 (n29888, pi0625, n29885);
  not g48763 (n_21882, n29887);
  and g48764 (n29889, pi1153, n_21882);
  not g48765 (n_21883, n29888);
  and g48766 (n29890, n_21883, n29889);
  and g48767 (n29891, n_11753, n29885);
  and g48768 (n29892, pi0625, n29870);
  not g48769 (n_21884, n29892);
  and g48770 (n29893, n_11757, n_21884);
  not g48771 (n_21885, n29891);
  and g48772 (n29894, n_21885, n29893);
  not g48773 (n_21886, n29890);
  not g48774 (n_21887, n29894);
  and g48775 (n29895, n_21886, n_21887);
  not g48776 (n_21888, n29895);
  and g48777 (n29896, pi0778, n_21888);
  not g48778 (n_21889, n29886);
  not g48779 (n_21890, n29896);
  and g48780 (n29897, n_21889, n_21890);
  not g48781 (n_21891, n29897);
  and g48782 (n29898, n_11773, n_21891);
  and g48783 (n29899, n17075, n_21871);
  not g48784 (n_21892, n29898);
  not g48785 (n_21893, n29899);
  and g48786 (n29900, n_21892, n_21893);
  and g48787 (n29901, n_11777, n29900);
  and g48788 (n29902, n16639, n29870);
  not g48789 (n_21894, n29901);
  not g48790 (n_21895, n29902);
  and g48791 (n29903, n_21894, n_21895);
  and g48792 (n29904, n_11780, n29903);
  not g48793 (n_21896, n29871);
  not g48794 (n_21897, n29904);
  and g48795 (n29905, n_21896, n_21897);
  and g48796 (n29906, n_11783, n29905);
  and g48797 (n29907, n16631, n29870);
  not g48798 (n_21898, n29906);
  not g48799 (n_21899, n29907);
  and g48800 (n29908, n_21898, n_21899);
  and g48801 (n29909, n_11787, n29908);
  and g48802 (n29910, n_11789, n29870);
  not g48803 (n_21900, n29908);
  and g48804 (n29911, pi0628, n_21900);
  not g48805 (n_21901, n29910);
  and g48806 (n29912, pi1156, n_21901);
  not g48807 (n_21902, n29911);
  and g48808 (n29913, n_21902, n29912);
  and g48809 (n29914, pi0628, n29870);
  and g48810 (n29915, n_11789, n_21900);
  not g48811 (n_21903, n29914);
  and g48812 (n29916, n_11794, n_21903);
  not g48813 (n_21904, n29915);
  and g48814 (n29917, n_21904, n29916);
  not g48815 (n_21905, n29913);
  not g48816 (n_21906, n29917);
  and g48817 (n29918, n_21905, n_21906);
  not g48818 (n_21907, n29918);
  and g48819 (n29919, pi0792, n_21907);
  not g48820 (n_21908, n29909);
  not g48821 (n_21909, n29919);
  and g48822 (n29920, n_21908, n_21909);
  not g48823 (n_21910, n29920);
  and g48824 (n29921, n_11803, n_21910);
  and g48825 (n29922, n_11806, n29870);
  and g48826 (n29923, pi0647, n29920);
  not g48827 (n_21911, n29922);
  and g48828 (n29924, pi1157, n_21911);
  not g48829 (n_21912, n29923);
  and g48830 (n29925, n_21912, n29924);
  and g48831 (n29926, n_11806, n29920);
  and g48832 (n29927, pi0647, n29870);
  not g48833 (n_21913, n29927);
  and g48834 (n29928, n_11810, n_21913);
  not g48835 (n_21914, n29926);
  and g48836 (n29929, n_21914, n29928);
  not g48837 (n_21915, n29925);
  not g48838 (n_21916, n29929);
  and g48839 (n29930, n_21915, n_21916);
  not g48840 (n_21917, n29930);
  and g48841 (n29931, pi0787, n_21917);
  not g48842 (n_21918, n29921);
  not g48843 (n_21919, n29931);
  and g48844 (n29932, n_21918, n_21919);
  and g48845 (n29933, n_11819, n29932);
  and g48846 (n29934, n_11984, n29870);
  and g48847 (n29935, n_15911, n_17780);
  not g48848 (n_21920, n22313);
  not g48849 (n_21921, n29935);
  and g48850 (n29936, n_21920, n_21921);
  not g48851 (n_21922, n29936);
  and g48852 (n29937, n_6272, n_21922);
  and g48853 (n29938, n_6272, n_13679);
  not g48854 (n_21923, n29938);
  and g48855 (n29939, n_15911, n_21923);
  and g48856 (n29940, n_17784, n29939);
  not g48857 (n_21924, n29937);
  not g48858 (n_21925, n29940);
  and g48859 (n29941, n_21924, n_21925);
  and g48860 (n29942, n2571, n29941);
  not g48861 (n_21926, n29942);
  and g48862 (n29943, n_21879, n_21926);
  not g48863 (n_21927, n29943);
  and g48864 (n29944, n_11960, n_21927);
  and g48865 (n29945, n17117, n_21871);
  not g48866 (n_21928, n29944);
  not g48867 (n_21929, n29945);
  and g48868 (n29946, n_21928, n_21929);
  not g48869 (n_21930, n29946);
  and g48870 (n29947, n_11964, n_21930);
  and g48871 (n29948, n_11967, n_21871);
  and g48872 (n29949, pi0609, n29944);
  not g48873 (n_21931, n29948);
  not g48874 (n_21932, n29949);
  and g48875 (n29950, n_21931, n_21932);
  not g48876 (n_21933, n29950);
  and g48877 (n29951, pi1155, n_21933);
  and g48878 (n29952, n_11972, n_21871);
  and g48879 (n29953, n_11971, n29944);
  not g48880 (n_21934, n29952);
  not g48881 (n_21935, n29953);
  and g48882 (n29954, n_21934, n_21935);
  not g48883 (n_21936, n29954);
  and g48884 (n29955, n_11768, n_21936);
  not g48885 (n_21937, n29951);
  not g48886 (n_21938, n29955);
  and g48887 (n29956, n_21937, n_21938);
  not g48888 (n_21939, n29956);
  and g48889 (n29957, pi0785, n_21939);
  not g48890 (n_21940, n29947);
  not g48891 (n_21941, n29957);
  and g48892 (n29958, n_21940, n_21941);
  and g48893 (n29959, pi0618, n29958);
  not g48894 (n_21942, n29934);
  and g48895 (n29960, pi1154, n_21942);
  not g48896 (n_21943, n29959);
  and g48897 (n29961, n_21943, n29960);
  and g48898 (n29962, pi0188, n19468);
  and g48899 (n29963, n_6272, n19477);
  and g48905 (n29967, n_6272, n_13718);
  and g48906 (n29968, pi0188, n19496);
  not g48907 (n_21946, n29967);
  and g48908 (n29969, n_15911, n_21946);
  not g48909 (n_21947, n29968);
  and g48910 (n29970, n_21947, n29969);
  not g48911 (n_21948, n29970);
  and g48912 (n29971, pi0705, n_21948);
  not g48913 (n_21949, n29966);
  and g48914 (n29972, n_21949, n29971);
  not g48915 (n_21950, n29941);
  and g48916 (n29973, n_15924, n_21950);
  not g48917 (n_21951, n29972);
  and g48918 (n29974, n2571, n_21951);
  not g48919 (n_21952, n29973);
  and g48920 (n29975, n_21952, n29974);
  not g48921 (n_21953, n29975);
  and g48922 (n29976, n_21879, n_21953);
  and g48923 (n29977, n_11753, n29976);
  and g48924 (n29978, pi0625, n29943);
  not g48925 (n_21954, n29978);
  and g48926 (n29979, n_11757, n_21954);
  not g48927 (n_21955, n29977);
  and g48928 (n29980, n_21955, n29979);
  and g48929 (n29981, n_11823, n_21886);
  not g48930 (n_21956, n29980);
  and g48931 (n29982, n_21956, n29981);
  and g48932 (n29983, n_11753, n29943);
  and g48933 (n29984, pi0625, n29976);
  not g48934 (n_21957, n29983);
  and g48935 (n29985, pi1153, n_21957);
  not g48936 (n_21958, n29984);
  and g48937 (n29986, n_21958, n29985);
  and g48938 (n29987, pi0608, n_21887);
  not g48939 (n_21959, n29986);
  and g48940 (n29988, n_21959, n29987);
  not g48941 (n_21960, n29982);
  not g48942 (n_21961, n29988);
  and g48943 (n29989, n_21960, n_21961);
  not g48944 (n_21962, n29989);
  and g48945 (n29990, pi0778, n_21962);
  and g48946 (n29991, n_11749, n29976);
  not g48947 (n_21963, n29990);
  not g48948 (n_21964, n29991);
  and g48949 (n29992, n_21963, n_21964);
  not g48950 (n_21965, n29992);
  and g48951 (n29993, n_11971, n_21965);
  and g48952 (n29994, pi0609, n29897);
  not g48953 (n_21966, n29994);
  and g48954 (n29995, n_11768, n_21966);
  not g48955 (n_21967, n29993);
  and g48956 (n29996, n_21967, n29995);
  and g48957 (n29997, n_11767, n_21937);
  not g48958 (n_21968, n29996);
  and g48959 (n29998, n_21968, n29997);
  and g48960 (n29999, n_11971, n29897);
  and g48961 (n30000, pi0609, n_21965);
  not g48962 (n_21969, n29999);
  and g48963 (n30001, pi1155, n_21969);
  not g48964 (n_21970, n30000);
  and g48965 (n30002, n_21970, n30001);
  and g48966 (n30003, pi0660, n_21938);
  not g48967 (n_21971, n30002);
  and g48968 (n30004, n_21971, n30003);
  not g48969 (n_21972, n29998);
  not g48970 (n_21973, n30004);
  and g48971 (n30005, n_21972, n_21973);
  not g48972 (n_21974, n30005);
  and g48973 (n30006, pi0785, n_21974);
  and g48974 (n30007, n_11964, n_21965);
  not g48975 (n_21975, n30006);
  not g48976 (n_21976, n30007);
  and g48977 (n30008, n_21975, n_21976);
  not g48978 (n_21977, n30008);
  and g48979 (n30009, n_11984, n_21977);
  and g48980 (n30010, pi0618, n29900);
  not g48981 (n_21978, n30010);
  and g48982 (n30011, n_11413, n_21978);
  not g48983 (n_21979, n30009);
  and g48984 (n30012, n_21979, n30011);
  not g48985 (n_21980, n29961);
  and g48986 (n30013, n_11412, n_21980);
  not g48987 (n_21981, n30012);
  and g48988 (n30014, n_21981, n30013);
  and g48989 (n30015, n_11984, n29958);
  and g48990 (n30016, pi0618, n29870);
  not g48991 (n_21982, n30016);
  and g48992 (n30017, n_11413, n_21982);
  not g48993 (n_21983, n30015);
  and g48994 (n30018, n_21983, n30017);
  and g48995 (n30019, n_11984, n29900);
  and g48996 (n30020, pi0618, n_21977);
  not g48997 (n_21984, n30019);
  and g48998 (n30021, pi1154, n_21984);
  not g48999 (n_21985, n30020);
  and g49000 (n30022, n_21985, n30021);
  not g49001 (n_21986, n30018);
  and g49002 (n30023, pi0627, n_21986);
  not g49003 (n_21987, n30022);
  and g49004 (n30024, n_21987, n30023);
  not g49005 (n_21988, n30014);
  not g49006 (n_21989, n30024);
  and g49007 (n30025, n_21988, n_21989);
  not g49008 (n_21990, n30025);
  and g49009 (n30026, pi0781, n_21990);
  and g49010 (n30027, n_11981, n_21977);
  not g49011 (n_21991, n30026);
  not g49012 (n_21992, n30027);
  and g49013 (n30028, n_21991, n_21992);
  not g49014 (n_21993, n30028);
  and g49015 (n30029, n_11821, n_21993);
  not g49016 (n_21994, n29903);
  and g49017 (n30030, pi0619, n_21994);
  not g49018 (n_21995, n30030);
  and g49019 (n30031, n_11405, n_21995);
  not g49020 (n_21996, n30029);
  and g49021 (n30032, n_21996, n30031);
  and g49022 (n30033, n_11821, n29870);
  not g49023 (n_21997, n29958);
  and g49024 (n30034, n_11981, n_21997);
  and g49025 (n30035, n_21980, n_21986);
  not g49026 (n_21998, n30035);
  and g49027 (n30036, pi0781, n_21998);
  not g49028 (n_21999, n30034);
  not g49029 (n_22000, n30036);
  and g49030 (n30037, n_21999, n_22000);
  and g49031 (n30038, pi0619, n30037);
  not g49032 (n_22001, n30033);
  and g49033 (n30039, pi1159, n_22001);
  not g49034 (n_22002, n30038);
  and g49035 (n30040, n_22002, n30039);
  not g49036 (n_22003, n30040);
  and g49037 (n30041, n_11403, n_22003);
  not g49038 (n_22004, n30032);
  and g49039 (n30042, n_22004, n30041);
  and g49040 (n30043, pi0619, n_21993);
  and g49041 (n30044, n_11821, n_21994);
  not g49042 (n_22005, n30044);
  and g49043 (n30045, pi1159, n_22005);
  not g49044 (n_22006, n30043);
  and g49045 (n30046, n_22006, n30045);
  and g49046 (n30047, n_11821, n30037);
  and g49047 (n30048, pi0619, n29870);
  not g49048 (n_22007, n30048);
  and g49049 (n30049, n_11405, n_22007);
  not g49050 (n_22008, n30047);
  and g49051 (n30050, n_22008, n30049);
  not g49052 (n_22009, n30050);
  and g49053 (n30051, pi0648, n_22009);
  not g49054 (n_22010, n30046);
  and g49055 (n30052, n_22010, n30051);
  not g49056 (n_22011, n30042);
  not g49057 (n_22012, n30052);
  and g49058 (n30053, n_22011, n_22012);
  not g49059 (n_22013, n30053);
  and g49060 (n30054, pi0789, n_22013);
  and g49061 (n30055, n_12315, n_21993);
  not g49062 (n_22014, n30054);
  not g49063 (n_22015, n30055);
  and g49064 (n30056, n_22014, n_22015);
  and g49065 (n30057, n_12318, n30056);
  and g49066 (n30058, n_12320, n30056);
  not g49067 (n_22016, n29905);
  and g49068 (n30059, pi0626, n_22016);
  not g49069 (n_22017, n30059);
  and g49070 (n30060, n_11395, n_22017);
  not g49071 (n_22018, n30058);
  and g49072 (n30061, n_22018, n30060);
  not g49073 (n_22019, n30037);
  and g49074 (n30062, n_12315, n_22019);
  and g49075 (n30063, n_22003, n_22009);
  not g49076 (n_22020, n30063);
  and g49077 (n30064, pi0789, n_22020);
  not g49078 (n_22021, n30062);
  not g49079 (n_22022, n30064);
  and g49080 (n30065, n_22021, n_22022);
  not g49081 (n_22023, n30065);
  and g49082 (n30066, n_12320, n_22023);
  and g49083 (n30067, pi0626, n_21871);
  not g49084 (n_22024, n30067);
  and g49085 (n30068, pi0641, n_22024);
  not g49086 (n_22025, n30066);
  and g49087 (n30069, n_22025, n30068);
  not g49088 (n_22026, n30069);
  and g49089 (n30070, n_11397, n_22026);
  not g49090 (n_22027, n30061);
  and g49091 (n30071, n_22027, n30070);
  and g49092 (n30072, pi0626, n30056);
  and g49093 (n30073, n_12320, n_22016);
  not g49094 (n_22028, n30073);
  and g49095 (n30074, pi0641, n_22028);
  not g49096 (n_22029, n30072);
  and g49097 (n30075, n_22029, n30074);
  and g49098 (n30076, pi0626, n_22023);
  and g49099 (n30077, n_12320, n_21871);
  not g49100 (n_22030, n30077);
  and g49101 (n30078, n_11395, n_22030);
  not g49102 (n_22031, n30076);
  and g49103 (n30079, n_22031, n30078);
  not g49104 (n_22032, n30079);
  and g49105 (n30080, pi1158, n_22032);
  not g49106 (n_22033, n30075);
  and g49107 (n30081, n_22033, n30080);
  not g49108 (n_22034, n30071);
  not g49109 (n_22035, n30081);
  and g49110 (n30082, n_22034, n_22035);
  not g49111 (n_22036, n30082);
  and g49112 (n30083, pi0788, n_22036);
  not g49113 (n_22037, n30057);
  not g49114 (n_22038, n30083);
  and g49115 (n30084, n_22037, n_22038);
  and g49116 (n30085, n_11789, n30084);
  and g49117 (n30086, n_12524, n30065);
  and g49118 (n30087, n17969, n29870);
  not g49119 (n_22039, n30086);
  not g49120 (n_22040, n30087);
  and g49121 (n30088, n_22039, n_22040);
  not g49122 (n_22041, n30088);
  and g49123 (n30089, pi0628, n_22041);
  not g49124 (n_22042, n30089);
  and g49125 (n30090, n_11794, n_22042);
  not g49126 (n_22043, n30085);
  and g49127 (n30091, n_22043, n30090);
  and g49128 (n30092, n_12354, n_21905);
  not g49129 (n_22044, n30091);
  and g49130 (n30093, n_22044, n30092);
  and g49131 (n30094, pi0628, n30084);
  and g49132 (n30095, n_11789, n_22041);
  not g49133 (n_22045, n30095);
  and g49134 (n30096, pi1156, n_22045);
  not g49135 (n_22046, n30094);
  and g49136 (n30097, n_22046, n30096);
  and g49137 (n30098, pi0629, n_21906);
  not g49138 (n_22047, n30097);
  and g49139 (n30099, n_22047, n30098);
  not g49140 (n_22048, n30093);
  not g49141 (n_22049, n30099);
  and g49142 (n30100, n_22048, n_22049);
  not g49143 (n_22050, n30100);
  and g49144 (n30101, pi0792, n_22050);
  and g49145 (n30102, n_11787, n30084);
  not g49146 (n_22051, n30101);
  not g49147 (n_22052, n30102);
  and g49148 (n30103, n_22051, n_22052);
  not g49149 (n_22053, n30103);
  and g49150 (n30104, n_11806, n_22053);
  and g49151 (n30105, n_12368, n_22041);
  and g49152 (n30106, n17779, n29870);
  not g49153 (n_22054, n30105);
  not g49154 (n_22055, n30106);
  and g49155 (n30107, n_22054, n_22055);
  not g49156 (n_22056, n30107);
  and g49157 (n30108, pi0647, n_22056);
  not g49158 (n_22057, n30108);
  and g49159 (n30109, n_11810, n_22057);
  not g49160 (n_22058, n30104);
  and g49161 (n30110, n_22058, n30109);
  and g49162 (n30111, n_12375, n_21915);
  not g49163 (n_22059, n30110);
  and g49164 (n30112, n_22059, n30111);
  and g49165 (n30113, pi0647, n_22053);
  and g49166 (n30114, n_11806, n_22056);
  not g49167 (n_22060, n30114);
  and g49168 (n30115, pi1157, n_22060);
  not g49169 (n_22061, n30113);
  and g49170 (n30116, n_22061, n30115);
  and g49171 (n30117, pi0630, n_21916);
  not g49172 (n_22062, n30116);
  and g49173 (n30118, n_22062, n30117);
  not g49174 (n_22063, n30112);
  not g49175 (n_22064, n30118);
  and g49176 (n30119, n_22063, n_22064);
  not g49177 (n_22065, n30119);
  and g49178 (n30120, pi0787, n_22065);
  and g49179 (n30121, n_11803, n_22053);
  not g49180 (n_22066, n30120);
  not g49181 (n_22067, n30121);
  and g49182 (n30122, n_22066, n_22067);
  not g49183 (n_22068, n30122);
  and g49184 (n30123, pi0644, n_22068);
  not g49185 (n_22069, n29933);
  and g49186 (n30124, pi0715, n_22069);
  not g49187 (n_22070, n30123);
  and g49188 (n30125, n_22070, n30124);
  and g49189 (n30126, n17804, n_21871);
  and g49190 (n30127, n_12392, n30107);
  not g49191 (n_22071, n30126);
  not g49192 (n_22072, n30127);
  and g49193 (n30128, n_22071, n_22072);
  and g49194 (n30129, pi0644, n30128);
  and g49195 (n30130, n_11819, n29870);
  not g49196 (n_22073, n30130);
  and g49197 (n30131, n_12395, n_22073);
  not g49198 (n_22074, n30129);
  and g49199 (n30132, n_22074, n30131);
  not g49200 (n_22075, n30132);
  and g49201 (n30133, pi1160, n_22075);
  not g49202 (n_22076, n30125);
  and g49203 (n30134, n_22076, n30133);
  and g49204 (n30135, n_11819, n_22068);
  and g49205 (n30136, pi0644, n29932);
  not g49206 (n_22077, n30136);
  and g49207 (n30137, n_12395, n_22077);
  not g49208 (n_22078, n30135);
  and g49209 (n30138, n_22078, n30137);
  and g49210 (n30139, n_11819, n30128);
  and g49211 (n30140, pi0644, n29870);
  not g49212 (n_22079, n30140);
  and g49213 (n30141, pi0715, n_22079);
  not g49214 (n_22080, n30139);
  and g49215 (n30142, n_22080, n30141);
  not g49216 (n_22081, n30142);
  and g49217 (n30143, n_12405, n_22081);
  not g49218 (n_22082, n30138);
  and g49219 (n30144, n_22082, n30143);
  not g49220 (n_22083, n30134);
  and g49221 (n30145, pi0790, n_22083);
  not g49222 (n_22084, n30144);
  and g49223 (n30146, n_22084, n30145);
  and g49224 (n30147, n_12411, n30122);
  not g49225 (n_22085, n30147);
  and g49226 (n30148, n_4226, n_22085);
  not g49227 (n_22086, n30146);
  and g49228 (n30149, n_22086, n30148);
  and g49229 (n30150, n_6272, po1038);
  not g49230 (n_22087, n30150);
  and g49231 (n30151, n_12415, n_22087);
  not g49232 (n_22088, n30149);
  and g49233 (n30152, n_22088, n30151);
  and g49234 (n30153, n_6272, n_12418);
  and g49235 (n30154, pi0705, n16645);
  not g49236 (n_22089, n30153);
  not g49237 (n_22090, n30154);
  and g49238 (n30155, n_22089, n_22090);
  and g49239 (n30156, n_11749, n30155);
  and g49240 (n30157, n_11753, n30154);
  not g49241 (n_22091, n30155);
  not g49242 (n_22092, n30157);
  and g49243 (n30158, n_22091, n_22092);
  not g49244 (n_22093, n30158);
  and g49245 (n30159, pi1153, n_22093);
  and g49246 (n30160, n_11757, n_22089);
  and g49247 (n30161, n_22092, n30160);
  not g49248 (n_22094, n30159);
  not g49249 (n_22095, n30161);
  and g49250 (n30162, n_22094, n_22095);
  not g49251 (n_22096, n30162);
  and g49252 (n30163, pi0778, n_22096);
  not g49253 (n_22097, n30156);
  not g49254 (n_22098, n30163);
  and g49255 (n30164, n_22097, n_22098);
  and g49256 (n30165, n_12429, n30164);
  and g49257 (n30166, n_12430, n30165);
  and g49258 (n30167, n_12431, n30166);
  and g49259 (n30168, n_12432, n30167);
  and g49260 (n30169, n_12436, n30168);
  and g49261 (n30170, n_11806, n30169);
  and g49262 (n30171, pi0647, n30153);
  not g49263 (n_22099, n30171);
  and g49264 (n30172, n_11810, n_22099);
  not g49265 (n_22100, n30170);
  and g49266 (n30173, n_22100, n30172);
  and g49267 (n30174, pi0630, n30173);
  and g49268 (n30175, n_15911, n17244);
  not g49269 (n_22101, n30175);
  and g49270 (n30176, n_22089, n_22101);
  not g49271 (n_22102, n30176);
  and g49272 (n30177, n_12448, n_22102);
  not g49273 (n_22103, n30177);
  and g49274 (n30178, n_11964, n_22103);
  and g49275 (n30179, n_12451, n_22102);
  not g49276 (n_22104, n30179);
  and g49277 (n30180, pi1155, n_22104);
  and g49278 (n30181, n_12453, n30177);
  not g49279 (n_22105, n30181);
  and g49280 (n30182, n_11768, n_22105);
  not g49281 (n_22106, n30180);
  not g49282 (n_22107, n30182);
  and g49283 (n30183, n_22106, n_22107);
  not g49284 (n_22108, n30183);
  and g49285 (n30184, pi0785, n_22108);
  not g49286 (n_22109, n30178);
  not g49287 (n_22110, n30184);
  and g49288 (n30185, n_22109, n_22110);
  not g49289 (n_22111, n30185);
  and g49290 (n30186, n_11981, n_22111);
  and g49291 (n30187, n_12461, n30185);
  not g49292 (n_22112, n30187);
  and g49293 (n30188, pi1154, n_22112);
  and g49294 (n30189, n_12463, n30185);
  not g49295 (n_22113, n30189);
  and g49296 (n30190, n_11413, n_22113);
  not g49297 (n_22114, n30188);
  not g49298 (n_22115, n30190);
  and g49299 (n30191, n_22114, n_22115);
  not g49300 (n_22116, n30191);
  and g49301 (n30192, pi0781, n_22116);
  not g49302 (n_22117, n30186);
  not g49303 (n_22118, n30192);
  and g49304 (n30193, n_22117, n_22118);
  not g49305 (n_22119, n30193);
  and g49306 (n30194, n_12315, n_22119);
  and g49307 (n30195, n_11821, n30153);
  and g49308 (n30196, pi0619, n30193);
  not g49309 (n_22120, n30195);
  and g49310 (n30197, pi1159, n_22120);
  not g49311 (n_22121, n30196);
  and g49312 (n30198, n_22121, n30197);
  and g49313 (n30199, n_11821, n30193);
  and g49314 (n30200, pi0619, n30153);
  not g49315 (n_22122, n30200);
  and g49316 (n30201, n_11405, n_22122);
  not g49317 (n_22123, n30199);
  and g49318 (n30202, n_22123, n30201);
  not g49319 (n_22124, n30198);
  not g49320 (n_22125, n30202);
  and g49321 (n30203, n_22124, n_22125);
  not g49322 (n_22126, n30203);
  and g49323 (n30204, pi0789, n_22126);
  not g49324 (n_22127, n30194);
  not g49325 (n_22128, n30204);
  and g49326 (n30205, n_22127, n_22128);
  and g49327 (n30206, n_12524, n30205);
  and g49328 (n30207, n17969, n30153);
  not g49329 (n_22129, n30206);
  not g49330 (n_22130, n30207);
  and g49331 (n30208, n_22129, n_22130);
  not g49332 (n_22131, n30208);
  and g49333 (n30209, n_12368, n_22131);
  and g49334 (n30210, n17779, n30153);
  not g49335 (n_22132, n30209);
  not g49336 (n_22133, n30210);
  and g49337 (n30211, n_22132, n_22133);
  and g49338 (n30212, n_14548, n30211);
  not g49339 (n_22134, n30169);
  and g49340 (n30213, pi0647, n_22134);
  and g49341 (n30214, n_11806, n_22089);
  not g49342 (n_22135, n30213);
  not g49343 (n_22136, n30214);
  and g49344 (n30215, n_22135, n_22136);
  not g49345 (n_22137, n30215);
  and g49346 (n30216, n17801, n_22137);
  not g49347 (n_22138, n30174);
  not g49348 (n_22139, n30216);
  and g49349 (n30217, n_22138, n_22139);
  not g49350 (n_22140, n30212);
  and g49351 (n30218, n_22140, n30217);
  not g49352 (n_22141, n30218);
  and g49353 (n30219, pi0787, n_22141);
  and g49354 (n30220, n17871, n30167);
  not g49355 (n_22142, n30205);
  and g49356 (n30221, n_12320, n_22142);
  and g49357 (n30222, pi0626, n_22089);
  not g49358 (n_22143, n30222);
  and g49359 (n30223, n16629, n_22143);
  not g49360 (n_22144, n30221);
  and g49361 (n30224, n_22144, n30223);
  and g49362 (n30225, pi0626, n_22142);
  and g49363 (n30226, n_12320, n_22089);
  not g49364 (n_22145, n30226);
  and g49365 (n30227, n16628, n_22145);
  not g49366 (n_22146, n30225);
  and g49367 (n30228, n_22146, n30227);
  not g49368 (n_22147, n30220);
  not g49369 (n_22148, n30224);
  and g49370 (n30229, n_22147, n_22148);
  not g49371 (n_22149, n30228);
  and g49372 (n30230, n_22149, n30229);
  not g49373 (n_22150, n30230);
  and g49374 (n30231, pi0788, n_22150);
  and g49375 (n30232, pi0618, n30165);
  and g49376 (n30233, pi0609, n30164);
  and g49377 (n30234, n_11866, n_22091);
  and g49378 (n30235, pi0625, n30234);
  not g49379 (n_22151, n30234);
  and g49380 (n30236, n30176, n_22151);
  not g49381 (n_22152, n30235);
  not g49382 (n_22153, n30236);
  and g49383 (n30237, n_22152, n_22153);
  not g49384 (n_22154, n30237);
  and g49385 (n30238, n30160, n_22154);
  and g49386 (n30239, n_11823, n_22094);
  not g49387 (n_22155, n30238);
  and g49388 (n30240, n_22155, n30239);
  and g49389 (n30241, pi1153, n30176);
  and g49390 (n30242, n_22152, n30241);
  and g49391 (n30243, pi0608, n_22095);
  not g49392 (n_22156, n30242);
  and g49393 (n30244, n_22156, n30243);
  not g49394 (n_22157, n30240);
  not g49395 (n_22158, n30244);
  and g49396 (n30245, n_22157, n_22158);
  not g49397 (n_22159, n30245);
  and g49398 (n30246, pi0778, n_22159);
  and g49399 (n30247, n_11749, n_22153);
  not g49400 (n_22160, n30246);
  not g49401 (n_22161, n30247);
  and g49402 (n30248, n_22160, n_22161);
  not g49403 (n_22162, n30248);
  and g49404 (n30249, n_11971, n_22162);
  not g49405 (n_22163, n30233);
  and g49406 (n30250, n_11768, n_22163);
  not g49407 (n_22164, n30249);
  and g49408 (n30251, n_22164, n30250);
  and g49409 (n30252, n_11767, n_22106);
  not g49410 (n_22165, n30251);
  and g49411 (n30253, n_22165, n30252);
  and g49412 (n30254, n_11971, n30164);
  and g49413 (n30255, pi0609, n_22162);
  not g49414 (n_22166, n30254);
  and g49415 (n30256, pi1155, n_22166);
  not g49416 (n_22167, n30255);
  and g49417 (n30257, n_22167, n30256);
  and g49418 (n30258, pi0660, n_22107);
  not g49419 (n_22168, n30257);
  and g49420 (n30259, n_22168, n30258);
  not g49421 (n_22169, n30253);
  not g49422 (n_22170, n30259);
  and g49423 (n30260, n_22169, n_22170);
  not g49424 (n_22171, n30260);
  and g49425 (n30261, pi0785, n_22171);
  and g49426 (n30262, n_11964, n_22162);
  not g49427 (n_22172, n30261);
  not g49428 (n_22173, n30262);
  and g49429 (n30263, n_22172, n_22173);
  not g49430 (n_22174, n30263);
  and g49431 (n30264, n_11984, n_22174);
  not g49432 (n_22175, n30232);
  and g49433 (n30265, n_11413, n_22175);
  not g49434 (n_22176, n30264);
  and g49435 (n30266, n_22176, n30265);
  and g49436 (n30267, n_11412, n_22114);
  not g49437 (n_22177, n30266);
  and g49438 (n30268, n_22177, n30267);
  and g49439 (n30269, n_11984, n30165);
  and g49440 (n30270, pi0618, n_22174);
  not g49441 (n_22178, n30269);
  and g49442 (n30271, pi1154, n_22178);
  not g49443 (n_22179, n30270);
  and g49444 (n30272, n_22179, n30271);
  and g49445 (n30273, pi0627, n_22115);
  not g49446 (n_22180, n30272);
  and g49447 (n30274, n_22180, n30273);
  not g49448 (n_22181, n30268);
  not g49449 (n_22182, n30274);
  and g49450 (n30275, n_22181, n_22182);
  not g49451 (n_22183, n30275);
  and g49452 (n30276, pi0781, n_22183);
  and g49453 (n30277, n_11981, n_22174);
  not g49454 (n_22184, n30276);
  not g49455 (n_22185, n30277);
  and g49456 (n30278, n_22184, n_22185);
  and g49457 (n30279, n_12315, n30278);
  not g49458 (n_22186, n30278);
  and g49459 (n30280, n_11821, n_22186);
  and g49460 (n30281, pi0619, n30166);
  not g49461 (n_22187, n30281);
  and g49462 (n30282, n_11405, n_22187);
  not g49463 (n_22188, n30280);
  and g49464 (n30283, n_22188, n30282);
  and g49465 (n30284, n_11403, n_22124);
  not g49466 (n_22189, n30283);
  and g49467 (n30285, n_22189, n30284);
  and g49468 (n30286, pi0619, n_22186);
  and g49469 (n30287, n_11821, n30166);
  not g49470 (n_22190, n30287);
  and g49471 (n30288, pi1159, n_22190);
  not g49472 (n_22191, n30286);
  and g49473 (n30289, n_22191, n30288);
  and g49474 (n30290, pi0648, n_22125);
  not g49475 (n_22192, n30289);
  and g49476 (n30291, n_22192, n30290);
  not g49477 (n_22193, n30285);
  and g49478 (n30292, pi0789, n_22193);
  not g49479 (n_22194, n30291);
  and g49480 (n30293, n_22194, n30292);
  not g49481 (n_22195, n30279);
  and g49482 (n30294, n17970, n_22195);
  not g49483 (n_22196, n30293);
  and g49484 (n30295, n_22196, n30294);
  not g49485 (n_22197, n30231);
  not g49486 (n_22198, n30295);
  and g49487 (n30296, n_22197, n_22198);
  not g49488 (n_22199, n30296);
  and g49489 (n30297, n_14638, n_22199);
  and g49490 (n30298, n17854, n_22131);
  and g49491 (n30299, n20851, n30168);
  not g49492 (n_22200, n30298);
  not g49493 (n_22201, n30299);
  and g49494 (n30300, n_22200, n_22201);
  not g49495 (n_22202, n30300);
  and g49496 (n30301, n_12354, n_22202);
  and g49497 (n30302, n20855, n30168);
  and g49498 (n30303, n17853, n_22131);
  not g49499 (n_22203, n30302);
  not g49500 (n_22204, n30303);
  and g49501 (n30304, n_22203, n_22204);
  not g49502 (n_22205, n30304);
  and g49503 (n30305, pi0629, n_22205);
  not g49504 (n_22206, n30301);
  not g49505 (n_22207, n30305);
  and g49506 (n30306, n_22206, n_22207);
  not g49507 (n_22208, n30306);
  and g49508 (n30307, pi0792, n_22208);
  not g49509 (n_22209, n30307);
  and g49510 (n30308, n_14387, n_22209);
  not g49511 (n_22210, n30297);
  and g49512 (n30309, n_22210, n30308);
  not g49513 (n_22211, n30219);
  not g49514 (n_22212, n30309);
  and g49515 (n30310, n_22211, n_22212);
  and g49516 (n30311, n_12411, n30310);
  and g49517 (n30312, n_11803, n_22134);
  and g49518 (n30313, pi1157, n_22137);
  not g49519 (n_22213, n30173);
  not g49520 (n_22214, n30313);
  and g49521 (n30314, n_22213, n_22214);
  not g49522 (n_22215, n30314);
  and g49523 (n30315, pi0787, n_22215);
  not g49524 (n_22216, n30312);
  not g49525 (n_22217, n30315);
  and g49526 (n30316, n_22216, n_22217);
  and g49527 (n30317, n_11819, n30316);
  and g49528 (n30318, pi0644, n30310);
  not g49529 (n_22218, n30317);
  and g49530 (n30319, pi0715, n_22218);
  not g49531 (n_22219, n30318);
  and g49532 (n30320, n_22219, n30319);
  not g49533 (n_22220, n30211);
  and g49534 (n30321, n_12392, n_22220);
  and g49535 (n30322, n17804, n30153);
  not g49536 (n_22221, n30321);
  not g49537 (n_22222, n30322);
  and g49538 (n30323, n_22221, n_22222);
  not g49539 (n_22223, n30323);
  and g49540 (n30324, pi0644, n_22223);
  and g49541 (n30325, n_11819, n30153);
  not g49542 (n_22224, n30325);
  and g49543 (n30326, n_12395, n_22224);
  not g49544 (n_22225, n30324);
  and g49545 (n30327, n_22225, n30326);
  not g49546 (n_22226, n30327);
  and g49547 (n30328, pi1160, n_22226);
  not g49548 (n_22227, n30320);
  and g49549 (n30329, n_22227, n30328);
  and g49550 (n30330, n_11819, n_22223);
  and g49551 (n30331, pi0644, n30153);
  not g49552 (n_22228, n30331);
  and g49553 (n30332, pi0715, n_22228);
  not g49554 (n_22229, n30330);
  and g49555 (n30333, n_22229, n30332);
  and g49556 (n30334, pi0644, n30316);
  and g49557 (n30335, n_11819, n30310);
  not g49558 (n_22230, n30334);
  and g49559 (n30336, n_12395, n_22230);
  not g49560 (n_22231, n30335);
  and g49561 (n30337, n_22231, n30336);
  not g49562 (n_22232, n30333);
  and g49563 (n30338, n_12405, n_22232);
  not g49564 (n_22233, n30337);
  and g49565 (n30339, n_22233, n30338);
  not g49566 (n_22234, n30329);
  not g49567 (n_22235, n30339);
  and g49568 (n30340, n_22234, n_22235);
  not g49569 (n_22236, n30340);
  and g49570 (n30341, pi0790, n_22236);
  not g49571 (n_22237, n30311);
  and g49572 (n30342, pi0832, n_22237);
  not g49573 (n_22238, n30341);
  and g49574 (n30343, n_22238, n30342);
  not g49575 (n_22239, n30152);
  not g49576 (n_22240, n30343);
  and g49577 (po0345, n_22239, n_22240);
  and g49578 (n30345, pi0189, n_11751);
  not g49579 (n_22241, n30345);
  and g49580 (n30346, n16635, n_22241);
  and g49581 (n30347, n17075, n_22241);
  and g49582 (n30348, pi0727, n2571);
  not g49583 (n_22242, n30348);
  and g49584 (n30349, n_22241, n_22242);
  and g49585 (n30350, n_301, n_11418);
  not g49586 (n_22243, n30350);
  and g49587 (n30351, n19899, n_22243);
  and g49588 (n30352, n_301, n18076);
  and g49589 (n30353, pi0189, n_14037);
  not g49590 (n_22244, n30352);
  and g49591 (n30354, n_161, n_22244);
  not g49592 (n_22245, n30353);
  and g49593 (n30355, n_22245, n30354);
  not g49594 (n_22246, n30351);
  and g49595 (n30356, n30348, n_22246);
  not g49596 (n_22247, n30355);
  and g49597 (n30357, n_22247, n30356);
  not g49598 (n_22248, n30349);
  not g49599 (n_22249, n30357);
  and g49600 (n30358, n_22248, n_22249);
  and g49601 (n30359, n_11749, n30358);
  and g49602 (n30360, n_11753, n_22241);
  not g49603 (n_22250, n30358);
  and g49604 (n30361, pi0625, n_22250);
  not g49605 (n_22251, n30360);
  and g49606 (n30362, pi1153, n_22251);
  not g49607 (n_22252, n30361);
  and g49608 (n30363, n_22252, n30362);
  and g49609 (n30364, n_11753, n_22250);
  and g49610 (n30365, pi0625, n_22241);
  not g49611 (n_22253, n30365);
  and g49612 (n30366, n_11757, n_22253);
  not g49613 (n_22254, n30364);
  and g49614 (n30367, n_22254, n30366);
  not g49615 (n_22255, n30363);
  not g49616 (n_22256, n30367);
  and g49617 (n30368, n_22255, n_22256);
  not g49618 (n_22257, n30368);
  and g49619 (n30369, pi0778, n_22257);
  not g49620 (n_22258, n30359);
  not g49621 (n_22259, n30369);
  and g49622 (n30370, n_22258, n_22259);
  and g49623 (n30371, n_11773, n30370);
  not g49624 (n_22260, n30347);
  not g49625 (n_22261, n30371);
  and g49626 (n30372, n_22260, n_22261);
  and g49627 (n30373, n_11777, n30372);
  and g49628 (n30374, n16639, n30345);
  not g49629 (n_22262, n30373);
  not g49630 (n_22263, n30374);
  and g49631 (n30375, n_22262, n_22263);
  and g49632 (n30376, n_11780, n30375);
  not g49633 (n_22264, n30346);
  not g49634 (n_22265, n30376);
  and g49635 (n30377, n_22264, n_22265);
  and g49636 (n30378, n_11783, n30377);
  and g49637 (n30379, n16631, n30345);
  not g49638 (n_22266, n30378);
  not g49639 (n_22267, n30379);
  and g49640 (n30380, n_22266, n_22267);
  not g49641 (n_22268, n30380);
  and g49642 (n30381, n_11787, n_22268);
  and g49643 (n30382, n_11789, n_22241);
  and g49644 (n30383, pi0628, n30380);
  not g49645 (n_22269, n30382);
  and g49646 (n30384, pi1156, n_22269);
  not g49647 (n_22270, n30383);
  and g49648 (n30385, n_22270, n30384);
  and g49649 (n30386, pi0628, n_22241);
  and g49650 (n30387, n_11789, n30380);
  not g49651 (n_22271, n30386);
  and g49652 (n30388, n_11794, n_22271);
  not g49653 (n_22272, n30387);
  and g49654 (n30389, n_22272, n30388);
  not g49655 (n_22273, n30385);
  not g49656 (n_22274, n30389);
  and g49657 (n30390, n_22273, n_22274);
  not g49658 (n_22275, n30390);
  and g49659 (n30391, pi0792, n_22275);
  not g49660 (n_22276, n30381);
  not g49661 (n_22277, n30391);
  and g49662 (n30392, n_22276, n_22277);
  not g49663 (n_22278, n30392);
  and g49664 (n30393, n_11803, n_22278);
  and g49665 (n30394, n_11806, n_22241);
  and g49666 (n30395, pi0647, n30392);
  not g49667 (n_22279, n30394);
  and g49668 (n30396, pi1157, n_22279);
  not g49669 (n_22280, n30395);
  and g49670 (n30397, n_22280, n30396);
  and g49671 (n30398, pi0647, n_22241);
  and g49672 (n30399, n_11806, n30392);
  not g49673 (n_22281, n30398);
  and g49674 (n30400, n_11810, n_22281);
  not g49675 (n_22282, n30399);
  and g49676 (n30401, n_22282, n30400);
  not g49677 (n_22283, n30397);
  not g49678 (n_22284, n30401);
  and g49679 (n30402, n_22283, n_22284);
  not g49680 (n_22285, n30402);
  and g49681 (n30403, pi0787, n_22285);
  not g49682 (n_22286, n30393);
  not g49683 (n_22287, n30403);
  and g49684 (n30404, n_22286, n_22287);
  and g49685 (n30405, n_11819, n30404);
  and g49686 (n30406, n_11821, n_22241);
  and g49687 (n30407, n17117, n_22241);
  and g49688 (n30408, pi0189, n_11417);
  and g49689 (n30409, pi0772, n17219);
  not g49690 (n_22288, n22241);
  not g49691 (n_22289, n30409);
  and g49692 (n30410, n_22288, n_22289);
  not g49693 (n_22290, n30410);
  and g49694 (n30411, pi0039, n_22290);
  and g49695 (n30412, n_15864, n16958);
  and g49696 (n30413, pi0772, n17139);
  not g49697 (n_22291, n30412);
  and g49698 (n30414, n_162, n_22291);
  not g49699 (n_22292, n30413);
  and g49700 (n30415, n_22292, n30414);
  not g49701 (n_22293, n30411);
  not g49702 (n_22294, n30415);
  and g49703 (n30416, n_22293, n_22294);
  not g49704 (n_22295, n30416);
  and g49705 (n30417, pi0189, n_22295);
  and g49706 (n30418, n_301, pi0772);
  and g49707 (n30419, n17275, n30418);
  not g49708 (n_22296, n30417);
  not g49709 (n_22297, n30419);
  and g49710 (n30420, n_22296, n_22297);
  not g49711 (n_22298, n30420);
  and g49712 (n30421, n_161, n_22298);
  and g49713 (n30422, pi0772, n17168);
  not g49714 (n_22299, n30422);
  and g49715 (n30423, n16641, n_22299);
  and g49716 (n30424, pi0038, n_22243);
  not g49717 (n_22300, n30423);
  and g49718 (n30425, n_22300, n30424);
  not g49719 (n_22301, n30421);
  not g49720 (n_22302, n30425);
  and g49721 (n30426, n_22301, n_22302);
  not g49722 (n_22303, n30426);
  and g49723 (n30427, n2571, n_22303);
  not g49724 (n_22304, n30408);
  not g49725 (n_22305, n30427);
  and g49726 (n30428, n_22304, n_22305);
  and g49727 (n30429, n_11960, n30428);
  not g49728 (n_22306, n30407);
  not g49729 (n_22307, n30429);
  and g49730 (n30430, n_22306, n_22307);
  and g49731 (n30431, n_11964, n30430);
  and g49732 (n30432, n_11971, n_22241);
  not g49733 (n_22308, n30430);
  and g49734 (n30433, pi0609, n_22308);
  not g49735 (n_22309, n30432);
  and g49736 (n30434, pi1155, n_22309);
  not g49737 (n_22310, n30433);
  and g49738 (n30435, n_22310, n30434);
  and g49739 (n30436, n_11971, n_22308);
  and g49740 (n30437, pi0609, n_22241);
  not g49741 (n_22311, n30437);
  and g49742 (n30438, n_11768, n_22311);
  not g49743 (n_22312, n30436);
  and g49744 (n30439, n_22312, n30438);
  not g49745 (n_22313, n30435);
  not g49746 (n_22314, n30439);
  and g49747 (n30440, n_22313, n_22314);
  not g49748 (n_22315, n30440);
  and g49749 (n30441, pi0785, n_22315);
  not g49750 (n_22316, n30431);
  not g49751 (n_22317, n30441);
  and g49752 (n30442, n_22316, n_22317);
  not g49753 (n_22318, n30442);
  and g49754 (n30443, n_11981, n_22318);
  and g49755 (n30444, n_11984, n_22241);
  and g49756 (n30445, pi0618, n30442);
  not g49757 (n_22319, n30444);
  and g49758 (n30446, pi1154, n_22319);
  not g49759 (n_22320, n30445);
  and g49760 (n30447, n_22320, n30446);
  and g49761 (n30448, pi0618, n_22241);
  and g49762 (n30449, n_11984, n30442);
  not g49763 (n_22321, n30448);
  and g49764 (n30450, n_11413, n_22321);
  not g49765 (n_22322, n30449);
  and g49766 (n30451, n_22322, n30450);
  not g49767 (n_22323, n30447);
  not g49768 (n_22324, n30451);
  and g49769 (n30452, n_22323, n_22324);
  not g49770 (n_22325, n30452);
  and g49771 (n30453, pi0781, n_22325);
  not g49772 (n_22326, n30443);
  not g49773 (n_22327, n30453);
  and g49774 (n30454, n_22326, n_22327);
  and g49775 (n30455, pi0619, n30454);
  not g49776 (n_22328, n30406);
  and g49777 (n30456, pi1159, n_22328);
  not g49778 (n_22329, n30455);
  and g49779 (n30457, n_22329, n30456);
  and g49780 (n30458, n_15870, n30426);
  and g49781 (n30459, n_301, n_13720);
  and g49782 (n30460, pi0189, n17546);
  not g49783 (n_22330, n30460);
  and g49784 (n30461, pi0772, n_22330);
  not g49785 (n_22331, n30459);
  and g49786 (n30462, n_22331, n30461);
  and g49787 (n30463, pi0189, n_13705);
  and g49788 (n30464, n_301, n_13702);
  not g49789 (n_22332, n30464);
  and g49790 (n30465, n_15864, n_22332);
  not g49791 (n_22333, n30463);
  and g49792 (n30466, n_22333, n30465);
  not g49793 (n_22334, n30462);
  and g49794 (n30467, pi0039, n_22334);
  not g49795 (n_22335, n30466);
  and g49796 (n30468, n_22335, n30467);
  and g49797 (n30469, n_301, n17631);
  and g49798 (n30470, pi0189, n17629);
  not g49799 (n_22336, n30469);
  and g49800 (n30471, pi0772, n_22336);
  not g49801 (n_22337, n30470);
  and g49802 (n30472, n_22337, n30471);
  and g49803 (n30473, n_301, n_12240);
  and g49804 (n30474, pi0189, n_12230);
  not g49805 (n_22338, n30473);
  and g49806 (n30475, n_15864, n_22338);
  not g49807 (n_22339, n30474);
  and g49808 (n30476, n_22339, n30475);
  not g49809 (n_22340, n30472);
  and g49810 (n30477, n_162, n_22340);
  not g49811 (n_22341, n30476);
  and g49812 (n30478, n_22341, n30477);
  not g49813 (n_22342, n30478);
  and g49814 (n30479, n_161, n_22342);
  not g49815 (n_22343, n30468);
  and g49816 (n30480, n_22343, n30479);
  not g49821 (n_22345, n30483);
  and g49822 (n30484, n2571, n_22345);
  not g49823 (n_22346, n30458);
  and g49824 (n30485, n_22346, n30484);
  not g49825 (n_22347, n30485);
  and g49826 (n30486, n_22304, n_22347);
  and g49827 (n30487, n_11753, n30486);
  and g49828 (n30488, pi0625, n30428);
  not g49829 (n_22348, n30488);
  and g49830 (n30489, n_11757, n_22348);
  not g49831 (n_22349, n30487);
  and g49832 (n30490, n_22349, n30489);
  and g49833 (n30491, n_11823, n_22255);
  not g49834 (n_22350, n30490);
  and g49835 (n30492, n_22350, n30491);
  and g49836 (n30493, n_11753, n30428);
  and g49837 (n30494, pi0625, n30486);
  not g49838 (n_22351, n30493);
  and g49839 (n30495, pi1153, n_22351);
  not g49840 (n_22352, n30494);
  and g49841 (n30496, n_22352, n30495);
  and g49842 (n30497, pi0608, n_22256);
  not g49843 (n_22353, n30496);
  and g49844 (n30498, n_22353, n30497);
  not g49845 (n_22354, n30492);
  not g49846 (n_22355, n30498);
  and g49847 (n30499, n_22354, n_22355);
  not g49848 (n_22356, n30499);
  and g49849 (n30500, pi0778, n_22356);
  and g49850 (n30501, n_11749, n30486);
  not g49851 (n_22357, n30500);
  not g49852 (n_22358, n30501);
  and g49853 (n30502, n_22357, n_22358);
  not g49854 (n_22359, n30502);
  and g49855 (n30503, n_11971, n_22359);
  and g49856 (n30504, pi0609, n30370);
  not g49857 (n_22360, n30504);
  and g49858 (n30505, n_11768, n_22360);
  not g49859 (n_22361, n30503);
  and g49860 (n30506, n_22361, n30505);
  and g49861 (n30507, n_11767, n_22313);
  not g49862 (n_22362, n30506);
  and g49863 (n30508, n_22362, n30507);
  and g49864 (n30509, n_11971, n30370);
  and g49865 (n30510, pi0609, n_22359);
  not g49866 (n_22363, n30509);
  and g49867 (n30511, pi1155, n_22363);
  not g49868 (n_22364, n30510);
  and g49869 (n30512, n_22364, n30511);
  and g49870 (n30513, pi0660, n_22314);
  not g49871 (n_22365, n30512);
  and g49872 (n30514, n_22365, n30513);
  not g49873 (n_22366, n30508);
  not g49874 (n_22367, n30514);
  and g49875 (n30515, n_22366, n_22367);
  not g49876 (n_22368, n30515);
  and g49877 (n30516, pi0785, n_22368);
  and g49878 (n30517, n_11964, n_22359);
  not g49879 (n_22369, n30516);
  not g49880 (n_22370, n30517);
  and g49881 (n30518, n_22369, n_22370);
  not g49882 (n_22371, n30518);
  and g49883 (n30519, n_11984, n_22371);
  not g49884 (n_22372, n30372);
  and g49885 (n30520, pi0618, n_22372);
  not g49886 (n_22373, n30520);
  and g49887 (n30521, n_11413, n_22373);
  not g49888 (n_22374, n30519);
  and g49889 (n30522, n_22374, n30521);
  and g49890 (n30523, n_11412, n_22323);
  not g49891 (n_22375, n30522);
  and g49892 (n30524, n_22375, n30523);
  and g49893 (n30525, pi0618, n_22371);
  and g49894 (n30526, n_11984, n_22372);
  not g49895 (n_22376, n30526);
  and g49896 (n30527, pi1154, n_22376);
  not g49897 (n_22377, n30525);
  and g49898 (n30528, n_22377, n30527);
  and g49899 (n30529, pi0627, n_22324);
  not g49900 (n_22378, n30528);
  and g49901 (n30530, n_22378, n30529);
  not g49902 (n_22379, n30524);
  not g49903 (n_22380, n30530);
  and g49904 (n30531, n_22379, n_22380);
  not g49905 (n_22381, n30531);
  and g49906 (n30532, pi0781, n_22381);
  and g49907 (n30533, n_11981, n_22371);
  not g49908 (n_22382, n30532);
  not g49909 (n_22383, n30533);
  and g49910 (n30534, n_22382, n_22383);
  not g49911 (n_22384, n30534);
  and g49912 (n30535, n_11821, n_22384);
  and g49913 (n30536, pi0619, n30375);
  not g49914 (n_22385, n30536);
  and g49915 (n30537, n_11405, n_22385);
  not g49916 (n_22386, n30535);
  and g49917 (n30538, n_22386, n30537);
  not g49918 (n_22387, n30457);
  and g49919 (n30539, n_11403, n_22387);
  not g49920 (n_22388, n30538);
  and g49921 (n30540, n_22388, n30539);
  and g49922 (n30541, pi0619, n_22241);
  and g49923 (n30542, n_11821, n30454);
  not g49924 (n_22389, n30541);
  and g49925 (n30543, n_11405, n_22389);
  not g49926 (n_22390, n30542);
  and g49927 (n30544, n_22390, n30543);
  and g49928 (n30545, n_11821, n30375);
  and g49929 (n30546, pi0619, n_22384);
  not g49930 (n_22391, n30545);
  and g49931 (n30547, pi1159, n_22391);
  not g49932 (n_22392, n30546);
  and g49933 (n30548, n_22392, n30547);
  not g49934 (n_22393, n30544);
  and g49935 (n30549, pi0648, n_22393);
  not g49936 (n_22394, n30548);
  and g49937 (n30550, n_22394, n30549);
  not g49938 (n_22395, n30540);
  not g49939 (n_22396, n30550);
  and g49940 (n30551, n_22395, n_22396);
  not g49941 (n_22397, n30551);
  and g49942 (n30552, pi0789, n_22397);
  and g49943 (n30553, n_12315, n_22384);
  not g49944 (n_22398, n30552);
  not g49945 (n_22399, n30553);
  and g49946 (n30554, n_22398, n_22399);
  and g49947 (n30555, n_12318, n30554);
  and g49948 (n30556, n_12320, n30554);
  and g49949 (n30557, pi0626, n30377);
  not g49950 (n_22400, n30557);
  and g49951 (n30558, n_11395, n_22400);
  not g49952 (n_22401, n30556);
  and g49953 (n30559, n_22401, n30558);
  not g49954 (n_22402, n30454);
  and g49955 (n30560, n_12315, n_22402);
  and g49956 (n30561, n_22387, n_22393);
  not g49957 (n_22403, n30561);
  and g49958 (n30562, pi0789, n_22403);
  not g49959 (n_22404, n30560);
  not g49960 (n_22405, n30562);
  and g49961 (n30563, n_22404, n_22405);
  not g49962 (n_22406, n30563);
  and g49963 (n30564, n_12320, n_22406);
  and g49964 (n30565, pi0626, n30345);
  not g49965 (n_22407, n30565);
  and g49966 (n30566, pi0641, n_22407);
  not g49967 (n_22408, n30564);
  and g49968 (n30567, n_22408, n30566);
  not g49969 (n_22409, n30567);
  and g49970 (n30568, n_11397, n_22409);
  not g49971 (n_22410, n30559);
  and g49972 (n30569, n_22410, n30568);
  and g49973 (n30570, pi0626, n30554);
  and g49974 (n30571, n_12320, n30377);
  not g49975 (n_22411, n30571);
  and g49976 (n30572, pi0641, n_22411);
  not g49977 (n_22412, n30570);
  and g49978 (n30573, n_22412, n30572);
  and g49979 (n30574, pi0626, n_22406);
  and g49980 (n30575, n_12320, n30345);
  not g49981 (n_22413, n30575);
  and g49982 (n30576, n_11395, n_22413);
  not g49983 (n_22414, n30574);
  and g49984 (n30577, n_22414, n30576);
  not g49985 (n_22415, n30577);
  and g49986 (n30578, pi1158, n_22415);
  not g49987 (n_22416, n30573);
  and g49988 (n30579, n_22416, n30578);
  not g49989 (n_22417, n30569);
  not g49990 (n_22418, n30579);
  and g49991 (n30580, n_22417, n_22418);
  not g49992 (n_22419, n30580);
  and g49993 (n30581, pi0788, n_22419);
  not g49994 (n_22420, n30555);
  not g49995 (n_22421, n30581);
  and g49996 (n30582, n_22420, n_22421);
  and g49997 (n30583, n_11789, n30582);
  and g49998 (n30584, n_12524, n_22406);
  and g49999 (n30585, n17969, n30345);
  not g50000 (n_22422, n30584);
  not g50001 (n_22423, n30585);
  and g50002 (n30586, n_22422, n_22423);
  and g50003 (n30587, pi0628, n30586);
  not g50004 (n_22424, n30587);
  and g50005 (n30588, n_11794, n_22424);
  not g50006 (n_22425, n30583);
  and g50007 (n30589, n_22425, n30588);
  and g50008 (n30590, n_12354, n_22273);
  not g50009 (n_22426, n30589);
  and g50010 (n30591, n_22426, n30590);
  and g50011 (n30592, pi0628, n30582);
  and g50012 (n30593, n_11789, n30586);
  not g50013 (n_22427, n30593);
  and g50014 (n30594, pi1156, n_22427);
  not g50015 (n_22428, n30592);
  and g50016 (n30595, n_22428, n30594);
  and g50017 (n30596, pi0629, n_22274);
  not g50018 (n_22429, n30595);
  and g50019 (n30597, n_22429, n30596);
  not g50020 (n_22430, n30591);
  not g50021 (n_22431, n30597);
  and g50022 (n30598, n_22430, n_22431);
  not g50023 (n_22432, n30598);
  and g50024 (n30599, pi0792, n_22432);
  and g50025 (n30600, n_11787, n30582);
  not g50026 (n_22433, n30599);
  not g50027 (n_22434, n30600);
  and g50028 (n30601, n_22433, n_22434);
  not g50029 (n_22435, n30601);
  and g50030 (n30602, n_11806, n_22435);
  not g50031 (n_22436, n30586);
  and g50032 (n30603, n_12368, n_22436);
  and g50033 (n30604, n17779, n30345);
  not g50034 (n_22437, n30603);
  not g50035 (n_22438, n30604);
  and g50036 (n30605, n_22437, n_22438);
  and g50037 (n30606, pi0647, n30605);
  not g50038 (n_22439, n30606);
  and g50039 (n30607, n_11810, n_22439);
  not g50040 (n_22440, n30602);
  and g50041 (n30608, n_22440, n30607);
  and g50042 (n30609, n_12375, n_22283);
  not g50043 (n_22441, n30608);
  and g50044 (n30610, n_22441, n30609);
  and g50045 (n30611, pi0647, n_22435);
  and g50046 (n30612, n_11806, n30605);
  not g50047 (n_22442, n30612);
  and g50048 (n30613, pi1157, n_22442);
  not g50049 (n_22443, n30611);
  and g50050 (n30614, n_22443, n30613);
  and g50051 (n30615, pi0630, n_22284);
  not g50052 (n_22444, n30614);
  and g50053 (n30616, n_22444, n30615);
  not g50054 (n_22445, n30610);
  not g50055 (n_22446, n30616);
  and g50056 (n30617, n_22445, n_22446);
  not g50057 (n_22447, n30617);
  and g50058 (n30618, pi0787, n_22447);
  and g50059 (n30619, n_11803, n_22435);
  not g50060 (n_22448, n30618);
  not g50061 (n_22449, n30619);
  and g50062 (n30620, n_22448, n_22449);
  not g50063 (n_22450, n30620);
  and g50064 (n30621, pi0644, n_22450);
  not g50065 (n_22451, n30405);
  and g50066 (n30622, pi0715, n_22451);
  not g50067 (n_22452, n30621);
  and g50068 (n30623, n_22452, n30622);
  and g50069 (n30624, n17804, n_22241);
  and g50070 (n30625, n_12392, n30605);
  not g50071 (n_22453, n30624);
  not g50072 (n_22454, n30625);
  and g50073 (n30626, n_22453, n_22454);
  not g50074 (n_22455, n30626);
  and g50075 (n30627, pi0644, n_22455);
  and g50076 (n30628, n_11819, n_22241);
  not g50077 (n_22456, n30628);
  and g50078 (n30629, n_12395, n_22456);
  not g50079 (n_22457, n30627);
  and g50080 (n30630, n_22457, n30629);
  not g50081 (n_22458, n30630);
  and g50082 (n30631, pi1160, n_22458);
  not g50083 (n_22459, n30623);
  and g50084 (n30632, n_22459, n30631);
  and g50085 (n30633, n_11819, n_22450);
  and g50086 (n30634, pi0644, n30404);
  not g50087 (n_22460, n30634);
  and g50088 (n30635, n_12395, n_22460);
  not g50089 (n_22461, n30633);
  and g50090 (n30636, n_22461, n30635);
  and g50091 (n30637, n_11819, n_22455);
  and g50092 (n30638, pi0644, n_22241);
  not g50093 (n_22462, n30638);
  and g50094 (n30639, pi0715, n_22462);
  not g50095 (n_22463, n30637);
  and g50096 (n30640, n_22463, n30639);
  not g50097 (n_22464, n30640);
  and g50098 (n30641, n_12405, n_22464);
  not g50099 (n_22465, n30636);
  and g50100 (n30642, n_22465, n30641);
  not g50101 (n_22466, n30632);
  and g50102 (n30643, pi0790, n_22466);
  not g50103 (n_22467, n30642);
  and g50104 (n30644, n_22467, n30643);
  and g50105 (n30645, n_12411, n30620);
  not g50106 (n_22468, n30645);
  and g50107 (n30646, n6305, n_22468);
  not g50108 (n_22469, n30644);
  and g50109 (n30647, n_22469, n30646);
  and g50110 (n30648, n_301, n_3232);
  not g50111 (n_22470, n30648);
  and g50112 (n30649, n_796, n_22470);
  not g50113 (n_22471, n30647);
  and g50114 (n30650, n_22471, n30649);
  and g50115 (n30651, pi0057, pi0189);
  not g50116 (n_22472, n30651);
  and g50117 (n30652, n_12415, n_22472);
  not g50118 (n_22473, n30650);
  and g50119 (n30653, n_22473, n30652);
  and g50120 (n30654, pi0189, n_12418);
  and g50121 (n30655, pi0772, n17244);
  and g50122 (n30656, n17291, n30655);
  not g50123 (n_22474, n30654);
  and g50124 (n30657, pi1155, n_22474);
  not g50125 (n_22475, n30656);
  and g50126 (n30658, n_22475, n30657);
  and g50127 (n30659, pi0727, n16645);
  not g50128 (n_22476, n30659);
  and g50129 (n30660, n_22474, n_22476);
  and g50130 (n30661, n_11749, n30660);
  and g50131 (n30662, pi0625, n30659);
  not g50132 (n_22477, n30660);
  not g50133 (n_22478, n30662);
  and g50134 (n30663, n_22477, n_22478);
  not g50135 (n_22479, n30663);
  and g50136 (n30664, n_11757, n_22479);
  and g50137 (n30665, pi1153, n_22474);
  and g50138 (n30666, n_22478, n30665);
  not g50139 (n_22480, n30664);
  not g50140 (n_22481, n30666);
  and g50141 (n30667, n_22480, n_22481);
  not g50142 (n_22482, n30667);
  and g50143 (n30668, pi0778, n_22482);
  not g50144 (n_22483, n30661);
  not g50145 (n_22484, n30668);
  and g50146 (n30669, n_22483, n_22484);
  and g50147 (n30670, pi0609, n30669);
  not g50148 (n_22485, n30655);
  and g50149 (n30671, n_22474, n_22485);
  and g50150 (n30672, pi0727, n17469);
  not g50151 (n_22486, n30672);
  and g50152 (n30673, n30671, n_22486);
  and g50153 (n30674, pi0625, n30672);
  not g50154 (n_22487, n30673);
  not g50155 (n_22488, n30674);
  and g50156 (n30675, n_22487, n_22488);
  not g50157 (n_22489, n30675);
  and g50158 (n30676, n_11757, n_22489);
  and g50159 (n30677, n_11823, n_22481);
  not g50160 (n_22490, n30676);
  and g50161 (n30678, n_22490, n30677);
  and g50162 (n30679, pi1153, n30671);
  and g50163 (n30680, n_22488, n30679);
  and g50164 (n30681, pi0608, n_22480);
  not g50165 (n_22491, n30680);
  and g50166 (n30682, n_22491, n30681);
  not g50167 (n_22492, n30678);
  not g50168 (n_22493, n30682);
  and g50169 (n30683, n_22492, n_22493);
  not g50170 (n_22494, n30683);
  and g50171 (n30684, pi0778, n_22494);
  and g50172 (n30685, n_11749, n_22487);
  not g50173 (n_22495, n30684);
  not g50174 (n_22496, n30685);
  and g50175 (n30686, n_22495, n_22496);
  not g50176 (n_22497, n30686);
  and g50177 (n30687, n_11971, n_22497);
  not g50178 (n_22498, n30670);
  and g50179 (n30688, n_11768, n_22498);
  not g50180 (n_22499, n30687);
  and g50181 (n30689, n_22499, n30688);
  not g50182 (n_22500, n30658);
  and g50183 (n30690, n_11767, n_22500);
  not g50184 (n_22501, n30689);
  and g50185 (n30691, n_22501, n30690);
  and g50186 (n30692, n17296, n30655);
  and g50187 (n30693, n_11768, n_22474);
  not g50188 (n_22502, n30692);
  and g50189 (n30694, n_22502, n30693);
  and g50190 (n30695, n_11971, n30669);
  and g50191 (n30696, pi0609, n_22497);
  not g50192 (n_22503, n30695);
  and g50193 (n30697, pi1155, n_22503);
  not g50194 (n_22504, n30696);
  and g50195 (n30698, n_22504, n30697);
  not g50196 (n_22505, n30694);
  and g50197 (n30699, pi0660, n_22505);
  not g50198 (n_22506, n30698);
  and g50199 (n30700, n_22506, n30699);
  not g50200 (n_22507, n30691);
  not g50201 (n_22508, n30700);
  and g50202 (n30701, n_22507, n_22508);
  not g50203 (n_22509, n30701);
  and g50204 (n30702, pi0785, n_22509);
  and g50205 (n30703, n_11964, n_22497);
  not g50206 (n_22510, n30702);
  not g50207 (n_22511, n30703);
  and g50208 (n30704, n_22510, n_22511);
  not g50209 (n_22512, n30704);
  and g50210 (n30705, n_11981, n_22512);
  and g50211 (n30706, n_14288, n30655);
  and g50212 (n30707, n20319, n30706);
  and g50213 (n30708, n_11413, n_22474);
  not g50214 (n_22513, n30707);
  and g50215 (n30709, n_22513, n30708);
  and g50216 (n30710, n_11773, n30669);
  not g50217 (n_22514, n30710);
  and g50218 (n30711, n_22474, n_22514);
  not g50219 (n_22515, n30711);
  and g50220 (n30712, n_11984, n_22515);
  and g50221 (n30713, pi0618, n_22512);
  not g50222 (n_22516, n30712);
  and g50223 (n30714, pi1154, n_22516);
  not g50224 (n_22517, n30713);
  and g50225 (n30715, n_22517, n30714);
  not g50226 (n_22518, n30709);
  and g50227 (n30716, pi0627, n_22518);
  not g50228 (n_22519, n30715);
  and g50229 (n30717, n_22519, n30716);
  and g50230 (n30718, n20270, n30706);
  and g50231 (n30719, pi1154, n_22474);
  not g50232 (n_22520, n30718);
  and g50233 (n30720, n_22520, n30719);
  and g50234 (n30721, pi0618, n_22515);
  and g50235 (n30722, n_11984, n_22512);
  not g50236 (n_22521, n30721);
  and g50237 (n30723, n_11413, n_22521);
  not g50238 (n_22522, n30722);
  and g50239 (n30724, n_22522, n30723);
  not g50240 (n_22523, n30720);
  and g50241 (n30725, n_11412, n_22523);
  not g50242 (n_22524, n30724);
  and g50243 (n30726, n_22524, n30725);
  not g50244 (n_22525, n30717);
  not g50245 (n_22526, n30726);
  and g50246 (n30727, n_22525, n_22526);
  not g50247 (n_22527, n30727);
  and g50248 (n30728, pi0781, n_22527);
  not g50249 (n_22528, n30705);
  and g50250 (n30729, n_16916, n_22528);
  not g50251 (n_22529, n30728);
  and g50252 (n30730, n_22529, n30729);
  and g50253 (n30731, n_14295, n30706);
  and g50254 (n30732, n20345, n30731);
  not g50255 (n_22530, n30732);
  and g50256 (n30733, n16633, n_22530);
  and g50257 (n30734, n19150, n30669);
  not g50258 (n_22531, n30734);
  and g50259 (n30735, n_16919, n_22531);
  and g50260 (n30736, n20335, n30731);
  not g50261 (n_22532, n30736);
  and g50262 (n30737, n16632, n_22532);
  not g50263 (n_22533, n30733);
  not g50264 (n_22534, n30737);
  and g50265 (n30738, n_22533, n_22534);
  not g50266 (n_22535, n30735);
  and g50267 (n30739, n_22535, n30738);
  and g50268 (n30740, pi0789, n_22474);
  not g50269 (n_22536, n30739);
  and g50270 (n30741, n_22536, n30740);
  not g50271 (n_22537, n30741);
  and g50272 (n30742, n17970, n_22537);
  not g50273 (n_22538, n30730);
  and g50274 (n30743, n_22538, n30742);
  and g50275 (n30744, n_11780, n30734);
  not g50276 (n_22539, n30744);
  and g50277 (n30745, n_22474, n_22539);
  not g50278 (n_22540, n30745);
  and g50279 (n30746, n17865, n_22540);
  and g50280 (n30747, n20237, n30706);
  and g50281 (n30748, n_12320, n30747);
  not g50282 (n_22541, n30748);
  and g50283 (n30749, n_22474, n_22541);
  not g50284 (n_22542, n30749);
  and g50285 (n30750, n_11397, n_22542);
  not g50286 (n_22543, n30750);
  and g50287 (n30751, pi0641, n_22543);
  not g50288 (n_22544, n30746);
  and g50289 (n30752, n_22544, n30751);
  and g50290 (n30753, pi0626, n30747);
  not g50291 (n_22545, n30753);
  and g50292 (n30754, n_22474, n_22545);
  not g50293 (n_22546, n30754);
  and g50294 (n30755, pi1158, n_22546);
  and g50295 (n30756, n17866, n_22540);
  not g50296 (n_22547, n30755);
  and g50297 (n30757, n_11395, n_22547);
  not g50298 (n_22548, n30756);
  and g50299 (n30758, n_22548, n30757);
  not g50300 (n_22549, n30752);
  and g50301 (n30759, pi0788, n_22549);
  not g50302 (n_22550, n30758);
  and g50303 (n30760, n_22550, n30759);
  not g50304 (n_22551, n30760);
  and g50305 (n30761, n_14638, n_22551);
  not g50306 (n_22552, n30743);
  and g50307 (n30762, n_22552, n30761);
  and g50308 (n30763, n_12524, n30747);
  and g50309 (n30764, n_12354, n30763);
  not g50310 (n_22553, n30764);
  and g50311 (n30765, pi0628, n_22553);
  and g50312 (n30766, n19151, n30669);
  not g50313 (n_22554, n30766);
  and g50314 (n30767, pi0629, n_22554);
  not g50315 (n_22555, n30765);
  not g50316 (n_22556, n30767);
  and g50317 (n30768, n_22555, n_22556);
  not g50318 (n_22557, n30768);
  and g50319 (n30769, n_11794, n_22557);
  not g50320 (n_22558, n30763);
  and g50321 (n30770, n_11789, n_22558);
  not g50322 (n_22559, n30770);
  and g50323 (n30771, pi0629, n_22559);
  and g50324 (n30772, pi0628, n30766);
  not g50325 (n_22560, n30771);
  and g50326 (n30773, pi1156, n_22560);
  not g50327 (n_22561, n30772);
  and g50328 (n30774, n_22561, n30773);
  not g50329 (n_22562, n30769);
  not g50330 (n_22563, n30774);
  and g50331 (n30775, n_22562, n_22563);
  and g50332 (n30776, pi0792, n_22474);
  not g50333 (n_22564, n30775);
  and g50334 (n30777, n_22564, n30776);
  not g50335 (n_22565, n30762);
  not g50336 (n_22566, n30777);
  and g50337 (n30778, n_22565, n_22566);
  not g50338 (n_22567, n30778);
  and g50339 (n30779, n_14387, n_22567);
  and g50340 (n30780, n_12368, n30763);
  and g50341 (n30781, n_12375, n30780);
  not g50342 (n_22568, n30781);
  and g50343 (n30782, pi0647, n_22568);
  and g50344 (n30783, n_13453, n30766);
  not g50345 (n_22569, n30783);
  and g50346 (n30784, pi0630, n_22569);
  not g50347 (n_22570, n30782);
  not g50348 (n_22571, n30784);
  and g50349 (n30785, n_22570, n_22571);
  not g50350 (n_22572, n30785);
  and g50351 (n30786, n_11810, n_22572);
  and g50352 (n30787, pi0630, n30780);
  and g50353 (n30788, n_12375, n_22569);
  not g50354 (n_22573, n30788);
  and g50355 (n30789, pi0647, n_22573);
  not g50356 (n_22574, n30787);
  and g50357 (n30790, pi1157, n_22574);
  not g50358 (n_22575, n30789);
  and g50359 (n30791, n_22575, n30790);
  not g50360 (n_22576, n30786);
  not g50361 (n_22577, n30791);
  and g50362 (n30792, n_22576, n_22577);
  and g50363 (n30793, pi0787, n_22474);
  not g50364 (n_22578, n30792);
  and g50365 (n30794, n_22578, n30793);
  not g50366 (n_22579, n30779);
  not g50367 (n_22580, n30794);
  and g50368 (n30795, n_22579, n_22580);
  and g50369 (n30796, n_12411, n30795);
  and g50370 (n30797, n_12524, n23684);
  and g50371 (n30798, n30747, n30797);
  and g50372 (n30799, pi0644, n30798);
  and g50373 (n30800, n_12395, n_22474);
  not g50374 (n_22581, n30799);
  and g50375 (n30801, n_22581, n30800);
  and g50376 (n30802, n_13598, n30783);
  not g50377 (n_22582, n30802);
  and g50378 (n30803, n_22474, n_22582);
  not g50379 (n_22583, n30803);
  and g50380 (n30804, n_11819, n_22583);
  and g50381 (n30805, pi0644, n30795);
  not g50382 (n_22584, n30804);
  and g50383 (n30806, pi0715, n_22584);
  not g50384 (n_22585, n30805);
  and g50385 (n30807, n_22585, n30806);
  not g50386 (n_22586, n30801);
  and g50387 (n30808, pi1160, n_22586);
  not g50388 (n_22587, n30807);
  and g50389 (n30809, n_22587, n30808);
  and g50390 (n30810, n_11819, n30798);
  and g50391 (n30811, pi0715, n_22474);
  not g50392 (n_22588, n30810);
  and g50393 (n30812, n_22588, n30811);
  and g50394 (n30813, n_11819, n30795);
  and g50395 (n30814, pi0644, n_22583);
  not g50396 (n_22589, n30814);
  and g50397 (n30815, n_12395, n_22589);
  not g50398 (n_22590, n30813);
  and g50399 (n30816, n_22590, n30815);
  not g50400 (n_22591, n30812);
  and g50401 (n30817, n_12405, n_22591);
  not g50402 (n_22592, n30816);
  and g50403 (n30818, n_22592, n30817);
  not g50404 (n_22593, n30809);
  not g50405 (n_22594, n30818);
  and g50406 (n30819, n_22593, n_22594);
  not g50407 (n_22595, n30819);
  and g50408 (n30820, pi0790, n_22595);
  not g50409 (n_22596, n30796);
  and g50410 (n30821, pi0832, n_22596);
  not g50411 (n_22597, n30820);
  and g50412 (n30822, n_22597, n30821);
  not g50413 (n_22598, n30653);
  not g50414 (n_22599, n30822);
  and g50415 (po0346, n_22598, n_22599);
  and g50416 (n30824, n_9199, n_12418);
  and g50417 (n30825, pi0699, n16645);
  not g50418 (n_22600, n30824);
  not g50419 (n_22601, n30825);
  and g50420 (n30826, n_22600, n_22601);
  not g50421 (n_22602, n30826);
  and g50422 (n30827, n_11749, n_22602);
  and g50423 (n30828, n_11753, n30825);
  not g50424 (n_22603, n30828);
  and g50425 (n30829, n_22602, n_22603);
  not g50426 (n_22604, n30829);
  and g50427 (n30830, pi1153, n_22604);
  and g50428 (n30831, n_11757, n_22600);
  and g50429 (n30832, n_22603, n30831);
  not g50430 (n_22605, n30832);
  and g50431 (n30833, pi0778, n_22605);
  not g50432 (n_22606, n30830);
  and g50433 (n30834, n_22606, n30833);
  not g50434 (n_22607, n30827);
  not g50435 (n_22608, n30834);
  and g50436 (n30835, n_22607, n_22608);
  not g50437 (n_22609, n30835);
  and g50438 (n30836, n_12429, n_22609);
  and g50439 (n30837, n_12430, n30836);
  and g50440 (n30838, n_12431, n30837);
  and g50441 (n30839, n_12432, n30838);
  and g50442 (n30840, n_12436, n30839);
  and g50443 (n30841, n_11806, n30840);
  and g50444 (n30842, pi0647, n30824);
  not g50445 (n_22610, n30842);
  and g50446 (n30843, n_11810, n_22610);
  not g50447 (n_22611, n30841);
  and g50448 (n30844, n_22611, n30843);
  and g50449 (n30845, pi0630, n30844);
  and g50450 (n30846, pi0763, n17244);
  not g50451 (n_22612, n30846);
  and g50452 (n30847, n_22600, n_22612);
  not g50453 (n_22613, n30847);
  and g50454 (n30848, n_12448, n_22613);
  not g50455 (n_22614, n30848);
  and g50456 (n30849, n_11964, n_22614);
  and g50457 (n30850, n17296, n30846);
  not g50458 (n_22615, n30850);
  and g50459 (n30851, n30848, n_22615);
  not g50460 (n_22616, n30851);
  and g50461 (n30852, pi1155, n_22616);
  and g50462 (n30853, n_11768, n_22600);
  and g50463 (n30854, n_22615, n30853);
  not g50464 (n_22617, n30852);
  not g50465 (n_22618, n30854);
  and g50466 (n30855, n_22617, n_22618);
  not g50467 (n_22619, n30855);
  and g50468 (n30856, pi0785, n_22619);
  not g50469 (n_22620, n30849);
  not g50470 (n_22621, n30856);
  and g50471 (n30857, n_22620, n_22621);
  not g50472 (n_22622, n30857);
  and g50473 (n30858, n_11981, n_22622);
  and g50474 (n30859, n_12461, n30857);
  not g50475 (n_22623, n30859);
  and g50476 (n30860, pi1154, n_22623);
  and g50477 (n30861, n_12463, n30857);
  not g50478 (n_22624, n30861);
  and g50479 (n30862, n_11413, n_22624);
  not g50480 (n_22625, n30860);
  not g50481 (n_22626, n30862);
  and g50482 (n30863, n_22625, n_22626);
  not g50483 (n_22627, n30863);
  and g50484 (n30864, pi0781, n_22627);
  not g50485 (n_22628, n30858);
  not g50486 (n_22629, n30864);
  and g50487 (n30865, n_22628, n_22629);
  not g50488 (n_22630, n30865);
  and g50489 (n30866, n_12315, n_22630);
  and g50490 (n30867, n_16503, n30865);
  not g50491 (n_22631, n30867);
  and g50492 (n30868, pi1159, n_22631);
  and g50493 (n30869, n_16505, n30865);
  not g50494 (n_22632, n30869);
  and g50495 (n30870, n_11405, n_22632);
  not g50496 (n_22633, n30868);
  not g50497 (n_22634, n30870);
  and g50498 (n30871, n_22633, n_22634);
  not g50499 (n_22635, n30871);
  and g50500 (n30872, pi0789, n_22635);
  not g50501 (n_22636, n30866);
  not g50502 (n_22637, n30872);
  and g50503 (n30873, n_22636, n_22637);
  and g50504 (n30874, n_12524, n30873);
  and g50505 (n30875, n17969, n30824);
  not g50506 (n_22638, n30874);
  not g50507 (n_22639, n30875);
  and g50508 (n30876, n_22638, n_22639);
  not g50509 (n_22640, n30876);
  and g50510 (n30877, n_12368, n_22640);
  and g50511 (n30878, n17779, n30824);
  not g50512 (n_22641, n30877);
  not g50513 (n_22642, n30878);
  and g50514 (n30879, n_22641, n_22642);
  and g50515 (n30880, n_14548, n30879);
  not g50516 (n_22643, n30840);
  and g50517 (n30881, pi0647, n_22643);
  and g50518 (n30882, n_11806, n_22600);
  not g50519 (n_22644, n30881);
  not g50520 (n_22645, n30882);
  and g50521 (n30883, n_22644, n_22645);
  not g50522 (n_22646, n30883);
  and g50523 (n30884, n17801, n_22646);
  not g50524 (n_22647, n30845);
  not g50525 (n_22648, n30884);
  and g50526 (n30885, n_22647, n_22648);
  not g50527 (n_22649, n30880);
  and g50528 (n30886, n_22649, n30885);
  not g50529 (n_22650, n30886);
  and g50530 (n30887, pi0787, n_22650);
  and g50531 (n30888, n17871, n30838);
  not g50532 (n_22651, n30873);
  and g50533 (n30889, n_12320, n_22651);
  and g50534 (n30890, pi0626, n_22600);
  not g50535 (n_22652, n30890);
  and g50536 (n30891, n16629, n_22652);
  not g50537 (n_22653, n30889);
  and g50538 (n30892, n_22653, n30891);
  and g50539 (n30893, pi0626, n_22651);
  and g50540 (n30894, n_12320, n_22600);
  not g50541 (n_22654, n30894);
  and g50542 (n30895, n16628, n_22654);
  not g50543 (n_22655, n30893);
  and g50544 (n30896, n_22655, n30895);
  not g50545 (n_22656, n30888);
  not g50546 (n_22657, n30892);
  and g50547 (n30897, n_22656, n_22657);
  not g50548 (n_22658, n30896);
  and g50549 (n30898, n_22658, n30897);
  not g50550 (n_22659, n30898);
  and g50551 (n30899, pi0788, n_22659);
  and g50552 (n30900, pi0618, n30836);
  and g50553 (n30901, n_11866, n_22602);
  and g50554 (n30902, pi0625, n30901);
  not g50555 (n_22660, n30901);
  and g50556 (n30903, n30847, n_22660);
  not g50557 (n_22661, n30902);
  not g50558 (n_22662, n30903);
  and g50559 (n30904, n_22661, n_22662);
  not g50560 (n_22663, n30904);
  and g50561 (n30905, n30831, n_22663);
  and g50562 (n30906, n_11823, n_22606);
  not g50563 (n_22664, n30905);
  and g50564 (n30907, n_22664, n30906);
  and g50565 (n30908, pi1153, n30847);
  and g50566 (n30909, n_22661, n30908);
  and g50567 (n30910, pi0608, n_22605);
  not g50568 (n_22665, n30909);
  and g50569 (n30911, n_22665, n30910);
  not g50570 (n_22666, n30907);
  not g50571 (n_22667, n30911);
  and g50572 (n30912, n_22666, n_22667);
  not g50573 (n_22668, n30912);
  and g50574 (n30913, pi0778, n_22668);
  and g50575 (n30914, n_11749, n_22662);
  not g50576 (n_22669, n30913);
  not g50577 (n_22670, n30914);
  and g50578 (n30915, n_22669, n_22670);
  not g50579 (n_22671, n30915);
  and g50580 (n30916, n_11971, n_22671);
  and g50581 (n30917, pi0609, n_22609);
  not g50582 (n_22672, n30917);
  and g50583 (n30918, n_11768, n_22672);
  not g50584 (n_22673, n30916);
  and g50585 (n30919, n_22673, n30918);
  and g50586 (n30920, n_11767, n_22617);
  not g50587 (n_22674, n30919);
  and g50588 (n30921, n_22674, n30920);
  and g50589 (n30922, pi0609, n_22671);
  and g50590 (n30923, n_11971, n_22609);
  not g50591 (n_22675, n30923);
  and g50592 (n30924, pi1155, n_22675);
  not g50593 (n_22676, n30922);
  and g50594 (n30925, n_22676, n30924);
  and g50595 (n30926, pi0660, n_22618);
  not g50596 (n_22677, n30925);
  and g50597 (n30927, n_22677, n30926);
  not g50598 (n_22678, n30921);
  not g50599 (n_22679, n30927);
  and g50600 (n30928, n_22678, n_22679);
  not g50601 (n_22680, n30928);
  and g50602 (n30929, pi0785, n_22680);
  and g50603 (n30930, n_11964, n_22671);
  not g50604 (n_22681, n30929);
  not g50605 (n_22682, n30930);
  and g50606 (n30931, n_22681, n_22682);
  not g50607 (n_22683, n30931);
  and g50608 (n30932, n_11984, n_22683);
  not g50609 (n_22684, n30900);
  and g50610 (n30933, n_11413, n_22684);
  not g50611 (n_22685, n30932);
  and g50612 (n30934, n_22685, n30933);
  and g50613 (n30935, n_11412, n_22625);
  not g50614 (n_22686, n30934);
  and g50615 (n30936, n_22686, n30935);
  and g50616 (n30937, n_11984, n30836);
  and g50617 (n30938, pi0618, n_22683);
  not g50618 (n_22687, n30937);
  and g50619 (n30939, pi1154, n_22687);
  not g50620 (n_22688, n30938);
  and g50621 (n30940, n_22688, n30939);
  and g50622 (n30941, pi0627, n_22626);
  not g50623 (n_22689, n30940);
  and g50624 (n30942, n_22689, n30941);
  not g50625 (n_22690, n30936);
  not g50626 (n_22691, n30942);
  and g50627 (n30943, n_22690, n_22691);
  not g50628 (n_22692, n30943);
  and g50629 (n30944, pi0781, n_22692);
  and g50630 (n30945, n_11981, n_22683);
  not g50631 (n_22693, n30944);
  not g50632 (n_22694, n30945);
  and g50633 (n30946, n_22693, n_22694);
  and g50634 (n30947, n_12315, n30946);
  not g50635 (n_22695, n30946);
  and g50636 (n30948, n_11821, n_22695);
  and g50637 (n30949, pi0619, n30837);
  not g50638 (n_22696, n30949);
  and g50639 (n30950, n_11405, n_22696);
  not g50640 (n_22697, n30948);
  and g50641 (n30951, n_22697, n30950);
  and g50642 (n30952, n_11403, n_22633);
  not g50643 (n_22698, n30951);
  and g50644 (n30953, n_22698, n30952);
  and g50645 (n30954, pi0619, n_22695);
  and g50646 (n30955, n_11821, n30837);
  not g50647 (n_22699, n30955);
  and g50648 (n30956, pi1159, n_22699);
  not g50649 (n_22700, n30954);
  and g50650 (n30957, n_22700, n30956);
  and g50651 (n30958, pi0648, n_22634);
  not g50652 (n_22701, n30957);
  and g50653 (n30959, n_22701, n30958);
  not g50654 (n_22702, n30953);
  and g50655 (n30960, pi0789, n_22702);
  not g50656 (n_22703, n30959);
  and g50657 (n30961, n_22703, n30960);
  not g50658 (n_22704, n30947);
  and g50659 (n30962, n17970, n_22704);
  not g50660 (n_22705, n30961);
  and g50661 (n30963, n_22705, n30962);
  not g50662 (n_22706, n30899);
  not g50663 (n_22707, n30963);
  and g50664 (n30964, n_22706, n_22707);
  not g50665 (n_22708, n30964);
  and g50666 (n30965, n_14638, n_22708);
  and g50667 (n30966, n17854, n_22640);
  and g50668 (n30967, n20851, n30839);
  not g50669 (n_22709, n30966);
  not g50670 (n_22710, n30967);
  and g50671 (n30968, n_22709, n_22710);
  not g50672 (n_22711, n30968);
  and g50673 (n30969, n_12354, n_22711);
  and g50674 (n30970, n20855, n30839);
  and g50675 (n30971, n17853, n_22640);
  not g50676 (n_22712, n30970);
  not g50677 (n_22713, n30971);
  and g50678 (n30972, n_22712, n_22713);
  not g50679 (n_22714, n30972);
  and g50680 (n30973, pi0629, n_22714);
  not g50681 (n_22715, n30969);
  not g50682 (n_22716, n30973);
  and g50683 (n30974, n_22715, n_22716);
  not g50684 (n_22717, n30974);
  and g50685 (n30975, pi0792, n_22717);
  not g50686 (n_22718, n30975);
  and g50687 (n30976, n_14387, n_22718);
  not g50688 (n_22719, n30965);
  and g50689 (n30977, n_22719, n30976);
  not g50690 (n_22720, n30887);
  not g50691 (n_22721, n30977);
  and g50692 (n30978, n_22720, n_22721);
  and g50693 (n30979, n_12411, n30978);
  and g50694 (n30980, n_11803, n_22643);
  and g50695 (n30981, pi1157, n_22646);
  not g50696 (n_22722, n30844);
  not g50697 (n_22723, n30981);
  and g50698 (n30982, n_22722, n_22723);
  not g50699 (n_22724, n30982);
  and g50700 (n30983, pi0787, n_22724);
  not g50701 (n_22725, n30980);
  not g50702 (n_22726, n30983);
  and g50703 (n30984, n_22725, n_22726);
  and g50704 (n30985, n_11819, n30984);
  and g50705 (n30986, pi0644, n30978);
  not g50706 (n_22727, n30985);
  and g50707 (n30987, pi0715, n_22727);
  not g50708 (n_22728, n30986);
  and g50709 (n30988, n_22728, n30987);
  not g50710 (n_22729, n30879);
  and g50711 (n30989, n_12392, n_22729);
  and g50712 (n30990, n17804, n30824);
  not g50713 (n_22730, n30989);
  not g50714 (n_22731, n30990);
  and g50715 (n30991, n_22730, n_22731);
  not g50716 (n_22732, n30991);
  and g50717 (n30992, pi0644, n_22732);
  and g50718 (n30993, n_11819, n30824);
  not g50719 (n_22733, n30993);
  and g50720 (n30994, n_12395, n_22733);
  not g50721 (n_22734, n30992);
  and g50722 (n30995, n_22734, n30994);
  not g50723 (n_22735, n30995);
  and g50724 (n30996, pi1160, n_22735);
  not g50725 (n_22736, n30988);
  and g50726 (n30997, n_22736, n30996);
  and g50727 (n30998, n_11819, n_22732);
  and g50728 (n30999, pi0644, n30824);
  not g50729 (n_22737, n30999);
  and g50730 (n31000, pi0715, n_22737);
  not g50731 (n_22738, n30998);
  and g50732 (n31001, n_22738, n31000);
  and g50733 (n31002, pi0644, n30984);
  and g50734 (n31003, n_11819, n30978);
  not g50735 (n_22739, n31002);
  and g50736 (n31004, n_12395, n_22739);
  not g50737 (n_22740, n31003);
  and g50738 (n31005, n_22740, n31004);
  not g50739 (n_22741, n31001);
  and g50740 (n31006, n_12405, n_22741);
  not g50741 (n_22742, n31005);
  and g50742 (n31007, n_22742, n31006);
  not g50743 (n_22743, n30997);
  not g50744 (n_22744, n31007);
  and g50745 (n31008, n_22743, n_22744);
  not g50746 (n_22745, n31008);
  and g50747 (n31009, pi0790, n_22745);
  not g50748 (n_22746, n30979);
  and g50749 (n31010, pi0832, n_22746);
  not g50750 (n_22747, n31009);
  and g50751 (n31011, n_22747, n31010);
  and g50752 (n31012, n_9199, po1038);
  and g50753 (n31013, n_9199, n_11751);
  not g50754 (n_22748, n31013);
  and g50755 (n31014, n16635, n_22748);
  and g50756 (n31015, pi0190, n_11417);
  and g50757 (n31016, n_9199, n_11418);
  not g50758 (n_22749, n31016);
  and g50759 (n31017, n16647, n_22749);
  and g50760 (n31018, n_9199, n18072);
  and g50761 (n31019, pi0190, n_12608);
  not g50762 (n_22750, n31019);
  and g50763 (n31020, n_161, n_22750);
  not g50764 (n_22751, n31018);
  and g50765 (n31021, n_22751, n31020);
  not g50766 (n_22752, n31017);
  and g50767 (n31022, pi0699, n_22752);
  not g50768 (n_22753, n31021);
  and g50769 (n31023, n_22753, n31022);
  and g50770 (n31024, n_9199, n_15996);
  and g50771 (n31025, n_11743, n31024);
  not g50772 (n_22754, n31025);
  and g50773 (n31026, n2571, n_22754);
  not g50774 (n_22755, n31023);
  and g50775 (n31027, n_22755, n31026);
  not g50776 (n_22756, n31015);
  not g50777 (n_22757, n31027);
  and g50778 (n31028, n_22756, n_22757);
  not g50779 (n_22758, n31028);
  and g50780 (n31029, n_11749, n_22758);
  and g50781 (n31030, n_11753, n31013);
  and g50782 (n31031, pi0625, n31028);
  not g50783 (n_22759, n31030);
  and g50784 (n31032, pi1153, n_22759);
  not g50785 (n_22760, n31031);
  and g50786 (n31033, n_22760, n31032);
  and g50787 (n31034, n_11753, n31028);
  and g50788 (n31035, pi0625, n31013);
  not g50789 (n_22761, n31035);
  and g50790 (n31036, n_11757, n_22761);
  not g50791 (n_22762, n31034);
  and g50792 (n31037, n_22762, n31036);
  not g50793 (n_22763, n31033);
  not g50794 (n_22764, n31037);
  and g50795 (n31038, n_22763, n_22764);
  not g50796 (n_22765, n31038);
  and g50797 (n31039, pi0778, n_22765);
  not g50798 (n_22766, n31029);
  not g50799 (n_22767, n31039);
  and g50800 (n31040, n_22766, n_22767);
  not g50801 (n_22768, n31040);
  and g50802 (n31041, n_11773, n_22768);
  and g50803 (n31042, n17075, n_22748);
  not g50804 (n_22769, n31041);
  not g50805 (n_22770, n31042);
  and g50806 (n31043, n_22769, n_22770);
  and g50807 (n31044, n_11777, n31043);
  and g50808 (n31045, n16639, n31013);
  not g50809 (n_22771, n31044);
  not g50810 (n_22772, n31045);
  and g50811 (n31046, n_22771, n_22772);
  and g50812 (n31047, n_11780, n31046);
  not g50813 (n_22773, n31014);
  not g50814 (n_22774, n31047);
  and g50815 (n31048, n_22773, n_22774);
  and g50816 (n31049, n_11783, n31048);
  and g50817 (n31050, n16631, n31013);
  not g50818 (n_22775, n31049);
  not g50819 (n_22776, n31050);
  and g50820 (n31051, n_22775, n_22776);
  not g50821 (n_22777, n31051);
  and g50822 (n31052, n_11789, n_22777);
  and g50823 (n31053, pi0628, n31013);
  not g50824 (n_22778, n31052);
  not g50825 (n_22779, n31053);
  and g50826 (n31054, n_22778, n_22779);
  not g50827 (n_22780, n31054);
  and g50828 (n31055, n_11794, n_22780);
  and g50829 (n31056, pi0628, n_22777);
  and g50830 (n31057, n_11789, n31013);
  not g50831 (n_22781, n31056);
  not g50832 (n_22782, n31057);
  and g50833 (n31058, n_22781, n_22782);
  not g50834 (n_22783, n31058);
  and g50835 (n31059, pi1156, n_22783);
  not g50836 (n_22784, n31055);
  not g50837 (n_22785, n31059);
  and g50838 (n31060, n_22784, n_22785);
  not g50839 (n_22786, n31060);
  and g50840 (n31061, pi0792, n_22786);
  and g50841 (n31062, n_11787, n_22777);
  not g50842 (n_22787, n31061);
  not g50843 (n_22788, n31062);
  and g50844 (n31063, n_22787, n_22788);
  not g50845 (n_22789, n31063);
  and g50846 (n31064, n_11806, n_22789);
  and g50847 (n31065, pi0647, n31013);
  not g50848 (n_22790, n31064);
  not g50849 (n_22791, n31065);
  and g50850 (n31066, n_22790, n_22791);
  not g50851 (n_22792, n31066);
  and g50852 (n31067, n_11810, n_22792);
  and g50853 (n31068, pi0647, n_22789);
  and g50854 (n31069, n_11806, n31013);
  not g50855 (n_22793, n31068);
  not g50856 (n_22794, n31069);
  and g50857 (n31070, n_22793, n_22794);
  not g50858 (n_22795, n31070);
  and g50859 (n31071, pi1157, n_22795);
  not g50860 (n_22796, n31067);
  not g50861 (n_22797, n31071);
  and g50862 (n31072, n_22796, n_22797);
  not g50863 (n_22798, n31072);
  and g50864 (n31073, pi0787, n_22798);
  and g50865 (n31074, n_11803, n_22789);
  not g50866 (n_22799, n31073);
  not g50867 (n_22800, n31074);
  and g50868 (n31075, n_22799, n_22800);
  not g50869 (n_22801, n31075);
  and g50870 (n31076, n_11819, n_22801);
  not g50871 (n_22802, n31076);
  and g50872 (n31077, pi0715, n_22802);
  and g50873 (n31078, n_15951, n17046);
  and g50874 (n31079, pi0190, n17273);
  not g50875 (n_22803, n31078);
  not g50876 (n_22804, n31079);
  and g50877 (n31080, n_22803, n_22804);
  not g50878 (n_22805, n31080);
  and g50879 (n31081, pi0039, n_22805);
  and g50880 (n31082, pi0763, n_11950);
  not g50881 (n_22806, n31082);
  and g50882 (n31083, pi0190, n_22806);
  and g50883 (n31084, n_9199, pi0763);
  and g50884 (n31085, n17221, n31084);
  not g50891 (n_22810, n31088);
  and g50892 (n31089, n_161, n_22810);
  and g50893 (n31090, pi0763, n17280);
  and g50894 (n31091, pi0038, n_22749);
  not g50895 (n_22811, n31090);
  and g50896 (n31092, n_22811, n31091);
  not g50897 (n_22812, n31089);
  not g50898 (n_22813, n31092);
  and g50899 (n31093, n_22812, n_22813);
  not g50900 (n_22814, n31093);
  and g50901 (n31094, n2571, n_22814);
  not g50902 (n_22815, n31094);
  and g50903 (n31095, n_22756, n_22815);
  not g50904 (n_22816, n31095);
  and g50905 (n31096, n_11960, n_22816);
  and g50906 (n31097, n17117, n_22748);
  not g50907 (n_22817, n31096);
  not g50908 (n_22818, n31097);
  and g50909 (n31098, n_22817, n_22818);
  not g50910 (n_22819, n31098);
  and g50911 (n31099, n_11964, n_22819);
  and g50912 (n31100, n_11967, n_22748);
  and g50913 (n31101, pi0609, n31096);
  not g50914 (n_22820, n31100);
  not g50915 (n_22821, n31101);
  and g50916 (n31102, n_22820, n_22821);
  not g50917 (n_22822, n31102);
  and g50918 (n31103, pi1155, n_22822);
  and g50919 (n31104, n_11972, n_22748);
  and g50920 (n31105, n_11971, n31096);
  not g50921 (n_22823, n31104);
  not g50922 (n_22824, n31105);
  and g50923 (n31106, n_22823, n_22824);
  not g50924 (n_22825, n31106);
  and g50925 (n31107, n_11768, n_22825);
  not g50926 (n_22826, n31103);
  not g50927 (n_22827, n31107);
  and g50928 (n31108, n_22826, n_22827);
  not g50929 (n_22828, n31108);
  and g50930 (n31109, pi0785, n_22828);
  not g50931 (n_22829, n31099);
  not g50932 (n_22830, n31109);
  and g50933 (n31110, n_22829, n_22830);
  not g50934 (n_22831, n31110);
  and g50935 (n31111, n_11981, n_22831);
  and g50936 (n31112, n_11984, n31013);
  and g50937 (n31113, pi0618, n31110);
  not g50938 (n_22832, n31112);
  and g50939 (n31114, pi1154, n_22832);
  not g50940 (n_22833, n31113);
  and g50941 (n31115, n_22833, n31114);
  and g50942 (n31116, n_11984, n31110);
  and g50943 (n31117, pi0618, n31013);
  not g50944 (n_22834, n31117);
  and g50945 (n31118, n_11413, n_22834);
  not g50946 (n_22835, n31116);
  and g50947 (n31119, n_22835, n31118);
  not g50948 (n_22836, n31115);
  not g50949 (n_22837, n31119);
  and g50950 (n31120, n_22836, n_22837);
  not g50951 (n_22838, n31120);
  and g50952 (n31121, pi0781, n_22838);
  not g50953 (n_22839, n31111);
  not g50954 (n_22840, n31121);
  and g50955 (n31122, n_22839, n_22840);
  not g50956 (n_22841, n31122);
  and g50957 (n31123, n_12315, n_22841);
  and g50958 (n31124, n_11821, n31013);
  and g50959 (n31125, pi0619, n31122);
  not g50960 (n_22842, n31124);
  and g50961 (n31126, pi1159, n_22842);
  not g50962 (n_22843, n31125);
  and g50963 (n31127, n_22843, n31126);
  and g50964 (n31128, n_11821, n31122);
  and g50965 (n31129, pi0619, n31013);
  not g50966 (n_22844, n31129);
  and g50967 (n31130, n_11405, n_22844);
  not g50968 (n_22845, n31128);
  and g50969 (n31131, n_22845, n31130);
  not g50970 (n_22846, n31127);
  not g50971 (n_22847, n31131);
  and g50972 (n31132, n_22846, n_22847);
  not g50973 (n_22848, n31132);
  and g50974 (n31133, pi0789, n_22848);
  not g50975 (n_22849, n31123);
  not g50976 (n_22850, n31133);
  and g50977 (n31134, n_22849, n_22850);
  and g50978 (n31135, n_12524, n31134);
  and g50979 (n31136, n17969, n31013);
  not g50980 (n_22851, n31135);
  not g50981 (n_22852, n31136);
  and g50982 (n31137, n_22851, n_22852);
  not g50983 (n_22853, n31137);
  and g50984 (n31138, n_12368, n_22853);
  and g50985 (n31139, n17779, n31013);
  not g50986 (n_22854, n31138);
  not g50987 (n_22855, n31139);
  and g50988 (n31140, n_22854, n_22855);
  not g50989 (n_22856, n31140);
  and g50990 (n31141, n_12392, n_22856);
  and g50991 (n31142, n17804, n31013);
  not g50992 (n_22857, n31141);
  not g50993 (n_22858, n31142);
  and g50994 (n31143, n_22857, n_22858);
  not g50995 (n_22859, n31143);
  and g50996 (n31144, pi0644, n_22859);
  and g50997 (n31145, n_11819, n31013);
  not g50998 (n_22860, n31145);
  and g50999 (n31146, n_12395, n_22860);
  not g51000 (n_22861, n31144);
  and g51001 (n31147, n_22861, n31146);
  not g51002 (n_22862, n31147);
  and g51003 (n31148, pi1160, n_22862);
  not g51004 (n_22863, n31077);
  and g51005 (n31149, n_22863, n31148);
  and g51006 (n31150, pi0644, n_22801);
  not g51007 (n_22864, n31150);
  and g51008 (n31151, n_12395, n_22864);
  and g51009 (n31152, n_11819, n_22859);
  and g51010 (n31153, pi0644, n31013);
  not g51011 (n_22865, n31153);
  and g51012 (n31154, pi0715, n_22865);
  not g51013 (n_22866, n31152);
  and g51014 (n31155, n_22866, n31154);
  not g51015 (n_22867, n31155);
  and g51016 (n31156, n_12405, n_22867);
  not g51017 (n_22868, n31151);
  and g51018 (n31157, n_22868, n31156);
  not g51019 (n_22869, n31149);
  not g51020 (n_22870, n31157);
  and g51021 (n31158, n_22869, n_22870);
  not g51022 (n_22871, n31158);
  and g51023 (n31159, pi0790, n_22871);
  and g51024 (n31160, n17777, n31054);
  and g51025 (n31161, n_14557, n31137);
  and g51026 (n31162, n17776, n31058);
  not g51027 (n_22872, n31160);
  not g51028 (n_22873, n31162);
  and g51029 (n31163, n_22872, n_22873);
  not g51030 (n_22874, n31161);
  and g51031 (n31164, n_22874, n31163);
  not g51032 (n_22875, n31164);
  and g51033 (n31165, pi0792, n_22875);
  and g51034 (n31166, pi0609, n31040);
  and g51035 (n31167, n_15996, n31093);
  and g51036 (n31168, n_15951, n24055);
  not g51037 (n_22876, n31168);
  and g51038 (n31169, n_12250, n_22876);
  not g51039 (n_22877, n31169);
  and g51040 (n31170, n_162, n_22877);
  not g51041 (n_22878, n31170);
  and g51042 (n31171, n_9199, n_22878);
  and g51043 (n31172, n_12120, n_22612);
  not g51044 (n_22879, n31172);
  and g51045 (n31173, pi0190, n_22879);
  and g51046 (n31174, n6284, n31173);
  not g51047 (n_22880, n31174);
  and g51048 (n31175, pi0038, n_22880);
  not g51049 (n_22881, n31171);
  and g51050 (n31176, n_22881, n31175);
  and g51051 (n31177, n_9199, n_12694);
  and g51052 (n31178, pi0190, n_12695);
  not g51053 (n_22882, n31178);
  and g51054 (n31179, pi0763, n_22882);
  not g51055 (n_22883, n31177);
  and g51056 (n31180, n_22883, n31179);
  and g51057 (n31181, n_9199, n17612);
  and g51058 (n31182, pi0190, n17625);
  not g51059 (n_22884, n31181);
  and g51060 (n31183, n_15951, n_22884);
  not g51061 (n_22885, n31182);
  and g51062 (n31184, n_22885, n31183);
  not g51063 (n_22886, n31180);
  and g51064 (n31185, n_162, n_22886);
  not g51065 (n_22887, n31184);
  and g51066 (n31186, n_22887, n31185);
  and g51067 (n31187, pi0190, n17605);
  and g51068 (n31188, n_9199, n_12180);
  not g51069 (n_22888, n31188);
  and g51070 (n31189, pi0763, n_22888);
  not g51071 (n_22889, n31187);
  and g51072 (n31190, n_22889, n31189);
  and g51073 (n31191, n_9199, n17404);
  and g51074 (n31192, pi0190, n17485);
  not g51075 (n_22890, n31192);
  and g51076 (n31193, n_15951, n_22890);
  not g51077 (n_22891, n31191);
  and g51078 (n31194, n_22891, n31193);
  not g51079 (n_22892, n31190);
  and g51080 (n31195, pi0039, n_22892);
  not g51081 (n_22893, n31194);
  and g51082 (n31196, n_22893, n31195);
  not g51083 (n_22894, n31186);
  and g51084 (n31197, n_161, n_22894);
  not g51085 (n_22895, n31196);
  and g51086 (n31198, n_22895, n31197);
  not g51087 (n_22896, n31176);
  and g51088 (n31199, pi0699, n_22896);
  not g51089 (n_22897, n31198);
  and g51090 (n31200, n_22897, n31199);
  not g51091 (n_22898, n31200);
  and g51092 (n31201, n2571, n_22898);
  not g51093 (n_22899, n31167);
  and g51094 (n31202, n_22899, n31201);
  not g51095 (n_22900, n31202);
  and g51096 (n31203, n_22756, n_22900);
  and g51097 (n31204, n_11753, n31203);
  and g51098 (n31205, pi0625, n31095);
  not g51099 (n_22901, n31205);
  and g51100 (n31206, n_11757, n_22901);
  not g51101 (n_22902, n31204);
  and g51102 (n31207, n_22902, n31206);
  and g51103 (n31208, n_11823, n_22763);
  not g51104 (n_22903, n31207);
  and g51105 (n31209, n_22903, n31208);
  and g51106 (n31210, n_11753, n31095);
  and g51107 (n31211, pi0625, n31203);
  not g51108 (n_22904, n31210);
  and g51109 (n31212, pi1153, n_22904);
  not g51110 (n_22905, n31211);
  and g51111 (n31213, n_22905, n31212);
  and g51112 (n31214, pi0608, n_22764);
  not g51113 (n_22906, n31213);
  and g51114 (n31215, n_22906, n31214);
  not g51115 (n_22907, n31209);
  not g51116 (n_22908, n31215);
  and g51117 (n31216, n_22907, n_22908);
  not g51118 (n_22909, n31216);
  and g51119 (n31217, pi0778, n_22909);
  and g51120 (n31218, n_11749, n31203);
  not g51121 (n_22910, n31217);
  not g51122 (n_22911, n31218);
  and g51123 (n31219, n_22910, n_22911);
  not g51124 (n_22912, n31219);
  and g51125 (n31220, n_11971, n_22912);
  not g51126 (n_22913, n31166);
  and g51127 (n31221, n_11768, n_22913);
  not g51128 (n_22914, n31220);
  and g51129 (n31222, n_22914, n31221);
  and g51130 (n31223, n_11767, n_22826);
  not g51131 (n_22915, n31222);
  and g51132 (n31224, n_22915, n31223);
  and g51133 (n31225, n_11971, n31040);
  and g51134 (n31226, pi0609, n_22912);
  not g51135 (n_22916, n31225);
  and g51136 (n31227, pi1155, n_22916);
  not g51137 (n_22917, n31226);
  and g51138 (n31228, n_22917, n31227);
  and g51139 (n31229, pi0660, n_22827);
  not g51140 (n_22918, n31228);
  and g51141 (n31230, n_22918, n31229);
  not g51142 (n_22919, n31224);
  not g51143 (n_22920, n31230);
  and g51144 (n31231, n_22919, n_22920);
  not g51145 (n_22921, n31231);
  and g51146 (n31232, pi0785, n_22921);
  and g51147 (n31233, n_11964, n_22912);
  not g51148 (n_22922, n31232);
  not g51149 (n_22923, n31233);
  and g51150 (n31234, n_22922, n_22923);
  not g51151 (n_22924, n31234);
  and g51152 (n31235, n_11984, n_22924);
  and g51153 (n31236, pi0618, n31043);
  not g51154 (n_22925, n31236);
  and g51155 (n31237, n_11413, n_22925);
  not g51156 (n_22926, n31235);
  and g51157 (n31238, n_22926, n31237);
  and g51158 (n31239, n_11412, n_22836);
  not g51159 (n_22927, n31238);
  and g51160 (n31240, n_22927, n31239);
  and g51161 (n31241, n_11984, n31043);
  and g51162 (n31242, pi0618, n_22924);
  not g51163 (n_22928, n31241);
  and g51164 (n31243, pi1154, n_22928);
  not g51165 (n_22929, n31242);
  and g51166 (n31244, n_22929, n31243);
  and g51167 (n31245, pi0627, n_22837);
  not g51168 (n_22930, n31244);
  and g51169 (n31246, n_22930, n31245);
  not g51170 (n_22931, n31240);
  not g51171 (n_22932, n31246);
  and g51172 (n31247, n_22931, n_22932);
  not g51173 (n_22933, n31247);
  and g51174 (n31248, pi0781, n_22933);
  and g51175 (n31249, n_11981, n_22924);
  not g51176 (n_22934, n31248);
  not g51177 (n_22935, n31249);
  and g51178 (n31250, n_22934, n_22935);
  and g51179 (n31251, n_12315, n31250);
  not g51180 (n_22936, n31046);
  and g51181 (n31252, pi0619, n_22936);
  not g51182 (n_22937, n31250);
  and g51183 (n31253, n_11821, n_22937);
  not g51184 (n_22938, n31252);
  and g51185 (n31254, n_11405, n_22938);
  not g51186 (n_22939, n31253);
  and g51187 (n31255, n_22939, n31254);
  and g51188 (n31256, n_11403, n_22846);
  not g51189 (n_22940, n31255);
  and g51190 (n31257, n_22940, n31256);
  and g51191 (n31258, n_11821, n_22936);
  and g51192 (n31259, pi0619, n_22937);
  not g51193 (n_22941, n31258);
  and g51194 (n31260, pi1159, n_22941);
  not g51195 (n_22942, n31259);
  and g51196 (n31261, n_22942, n31260);
  and g51197 (n31262, pi0648, n_22847);
  not g51198 (n_22943, n31261);
  and g51199 (n31263, n_22943, n31262);
  not g51200 (n_22944, n31257);
  and g51201 (n31264, pi0789, n_22944);
  not g51202 (n_22945, n31263);
  and g51203 (n31265, n_22945, n31264);
  not g51204 (n_22946, n31251);
  and g51205 (n31266, n17970, n_22946);
  not g51206 (n_22947, n31265);
  and g51207 (n31267, n_22947, n31266);
  and g51208 (n31268, n17871, n31048);
  not g51209 (n_22948, n31134);
  and g51210 (n31269, n_12320, n_22948);
  and g51211 (n31270, pi0626, n_22748);
  not g51212 (n_22949, n31270);
  and g51213 (n31271, n16629, n_22949);
  not g51214 (n_22950, n31269);
  and g51215 (n31272, n_22950, n31271);
  and g51216 (n31273, pi0626, n_22948);
  and g51217 (n31274, n_12320, n_22748);
  not g51218 (n_22951, n31274);
  and g51219 (n31275, n16628, n_22951);
  not g51220 (n_22952, n31273);
  and g51221 (n31276, n_22952, n31275);
  not g51222 (n_22953, n31268);
  not g51223 (n_22954, n31272);
  and g51224 (n31277, n_22953, n_22954);
  not g51225 (n_22955, n31276);
  and g51226 (n31278, n_22955, n31277);
  not g51227 (n_22956, n31278);
  and g51228 (n31279, pi0788, n_22956);
  not g51229 (n_22957, n31279);
  and g51230 (n31280, n_14638, n_22957);
  not g51231 (n_22958, n31267);
  and g51232 (n31281, n_22958, n31280);
  not g51233 (n_22959, n31165);
  not g51234 (n_22960, n31281);
  and g51235 (n31282, n_22959, n_22960);
  not g51236 (n_22961, n31282);
  and g51237 (n31283, n_14387, n_22961);
  and g51238 (n31284, n17802, n31066);
  and g51239 (n31285, n_14548, n31140);
  and g51240 (n31286, n17801, n31070);
  not g51241 (n_22962, n31284);
  not g51242 (n_22963, n31285);
  and g51243 (n31287, n_22962, n_22963);
  not g51244 (n_22964, n31286);
  and g51245 (n31288, n_22964, n31287);
  not g51246 (n_22965, n31288);
  and g51247 (n31289, pi0787, n_22965);
  and g51248 (n31290, n_11819, n31156);
  and g51249 (n31291, pi0644, n31148);
  not g51250 (n_22966, n31290);
  and g51251 (n31292, pi0790, n_22966);
  not g51252 (n_22967, n31291);
  and g51253 (n31293, n_22967, n31292);
  not g51254 (n_22968, n31283);
  not g51255 (n_22969, n31289);
  and g51256 (n31294, n_22968, n_22969);
  not g51257 (n_22970, n31293);
  and g51258 (n31295, n_22970, n31294);
  not g51259 (n_22971, n31159);
  not g51260 (n_22972, n31295);
  and g51261 (n31296, n_22971, n_22972);
  not g51262 (n_22973, n31296);
  and g51263 (n31297, n_4226, n_22973);
  not g51264 (n_22974, n31012);
  and g51265 (n31298, n_12415, n_22974);
  not g51266 (n_22975, n31297);
  and g51267 (n31299, n_22975, n31298);
  not g51268 (n_22976, n31011);
  not g51269 (n_22977, n31299);
  and g51270 (po0347, n_22976, n_22977);
  and g51271 (n31301, n_10720, n_12418);
  and g51272 (n31302, pi0729, n16645);
  not g51273 (n_22978, n31301);
  not g51274 (n_22979, n31302);
  and g51275 (n31303, n_22978, n_22979);
  not g51276 (n_22980, n31303);
  and g51277 (n31304, n_11749, n_22980);
  and g51278 (n31305, n_11753, n31302);
  not g51279 (n_22981, n31305);
  and g51280 (n31306, n_22980, n_22981);
  not g51281 (n_22982, n31306);
  and g51282 (n31307, pi1153, n_22982);
  and g51283 (n31308, n_11757, n_22978);
  and g51284 (n31309, n_22981, n31308);
  not g51285 (n_22983, n31309);
  and g51286 (n31310, pi0778, n_22983);
  not g51287 (n_22984, n31307);
  and g51288 (n31311, n_22984, n31310);
  not g51289 (n_22985, n31304);
  not g51290 (n_22986, n31311);
  and g51291 (n31312, n_22985, n_22986);
  not g51292 (n_22987, n31312);
  and g51293 (n31313, n_12429, n_22987);
  and g51294 (n31314, n_12430, n31313);
  and g51295 (n31315, n_12431, n31314);
  and g51296 (n31316, n_12432, n31315);
  and g51297 (n31317, n_12436, n31316);
  and g51298 (n31318, n_11806, n31317);
  and g51299 (n31319, pi0647, n31301);
  not g51300 (n_22988, n31319);
  and g51301 (n31320, n_11810, n_22988);
  not g51302 (n_22989, n31318);
  and g51303 (n31321, n_22989, n31320);
  and g51304 (n31322, pi0630, n31321);
  and g51305 (n31323, pi0746, n17244);
  not g51306 (n_22990, n31323);
  and g51307 (n31324, n_22978, n_22990);
  not g51308 (n_22991, n31324);
  and g51309 (n31325, n_12448, n_22991);
  not g51310 (n_22992, n31325);
  and g51311 (n31326, n_11964, n_22992);
  and g51312 (n31327, n17296, n31323);
  not g51313 (n_22993, n31327);
  and g51314 (n31328, n31325, n_22993);
  not g51315 (n_22994, n31328);
  and g51316 (n31329, pi1155, n_22994);
  and g51317 (n31330, n_11768, n_22978);
  and g51318 (n31331, n_22993, n31330);
  not g51319 (n_22995, n31329);
  not g51320 (n_22996, n31331);
  and g51321 (n31332, n_22995, n_22996);
  not g51322 (n_22997, n31332);
  and g51323 (n31333, pi0785, n_22997);
  not g51324 (n_22998, n31326);
  not g51325 (n_22999, n31333);
  and g51326 (n31334, n_22998, n_22999);
  not g51327 (n_23000, n31334);
  and g51328 (n31335, n_11981, n_23000);
  and g51329 (n31336, n_12461, n31334);
  not g51330 (n_23001, n31336);
  and g51331 (n31337, pi1154, n_23001);
  and g51332 (n31338, n_12463, n31334);
  not g51333 (n_23002, n31338);
  and g51334 (n31339, n_11413, n_23002);
  not g51335 (n_23003, n31337);
  not g51336 (n_23004, n31339);
  and g51337 (n31340, n_23003, n_23004);
  not g51338 (n_23005, n31340);
  and g51339 (n31341, pi0781, n_23005);
  not g51340 (n_23006, n31335);
  not g51341 (n_23007, n31341);
  and g51342 (n31342, n_23006, n_23007);
  not g51343 (n_23008, n31342);
  and g51344 (n31343, n_12315, n_23008);
  and g51345 (n31344, n_16503, n31342);
  not g51346 (n_23009, n31344);
  and g51347 (n31345, pi1159, n_23009);
  and g51348 (n31346, n_16505, n31342);
  not g51349 (n_23010, n31346);
  and g51350 (n31347, n_11405, n_23010);
  not g51351 (n_23011, n31345);
  not g51352 (n_23012, n31347);
  and g51353 (n31348, n_23011, n_23012);
  not g51354 (n_23013, n31348);
  and g51355 (n31349, pi0789, n_23013);
  not g51356 (n_23014, n31343);
  not g51357 (n_23015, n31349);
  and g51358 (n31350, n_23014, n_23015);
  and g51359 (n31351, n_12524, n31350);
  and g51360 (n31352, n17969, n31301);
  not g51361 (n_23016, n31351);
  not g51362 (n_23017, n31352);
  and g51363 (n31353, n_23016, n_23017);
  not g51364 (n_23018, n31353);
  and g51365 (n31354, n_12368, n_23018);
  and g51366 (n31355, n17779, n31301);
  not g51367 (n_23019, n31354);
  not g51368 (n_23020, n31355);
  and g51369 (n31356, n_23019, n_23020);
  and g51370 (n31357, n_14548, n31356);
  not g51371 (n_23021, n31317);
  and g51372 (n31358, pi0647, n_23021);
  and g51373 (n31359, n_11806, n_22978);
  not g51374 (n_23022, n31358);
  not g51375 (n_23023, n31359);
  and g51376 (n31360, n_23022, n_23023);
  not g51377 (n_23024, n31360);
  and g51378 (n31361, n17801, n_23024);
  not g51379 (n_23025, n31322);
  not g51380 (n_23026, n31361);
  and g51381 (n31362, n_23025, n_23026);
  not g51382 (n_23027, n31357);
  and g51383 (n31363, n_23027, n31362);
  not g51384 (n_23028, n31363);
  and g51385 (n31364, pi0787, n_23028);
  and g51386 (n31365, n17871, n31315);
  not g51387 (n_23029, n31350);
  and g51388 (n31366, n_12320, n_23029);
  and g51389 (n31367, pi0626, n_22978);
  not g51390 (n_23030, n31367);
  and g51391 (n31368, n16629, n_23030);
  not g51392 (n_23031, n31366);
  and g51393 (n31369, n_23031, n31368);
  and g51394 (n31370, pi0626, n_23029);
  and g51395 (n31371, n_12320, n_22978);
  not g51396 (n_23032, n31371);
  and g51397 (n31372, n16628, n_23032);
  not g51398 (n_23033, n31370);
  and g51399 (n31373, n_23033, n31372);
  not g51400 (n_23034, n31365);
  not g51401 (n_23035, n31369);
  and g51402 (n31374, n_23034, n_23035);
  not g51403 (n_23036, n31373);
  and g51404 (n31375, n_23036, n31374);
  not g51405 (n_23037, n31375);
  and g51406 (n31376, pi0788, n_23037);
  and g51407 (n31377, pi0618, n31313);
  and g51408 (n31378, n_11866, n_22980);
  and g51409 (n31379, pi0625, n31378);
  not g51410 (n_23038, n31378);
  and g51411 (n31380, n31324, n_23038);
  not g51412 (n_23039, n31379);
  not g51413 (n_23040, n31380);
  and g51414 (n31381, n_23039, n_23040);
  not g51415 (n_23041, n31381);
  and g51416 (n31382, n31308, n_23041);
  and g51417 (n31383, n_11823, n_22984);
  not g51418 (n_23042, n31382);
  and g51419 (n31384, n_23042, n31383);
  and g51420 (n31385, pi1153, n31324);
  and g51421 (n31386, n_23039, n31385);
  and g51422 (n31387, pi0608, n_22983);
  not g51423 (n_23043, n31386);
  and g51424 (n31388, n_23043, n31387);
  not g51425 (n_23044, n31384);
  not g51426 (n_23045, n31388);
  and g51427 (n31389, n_23044, n_23045);
  not g51428 (n_23046, n31389);
  and g51429 (n31390, pi0778, n_23046);
  and g51430 (n31391, n_11749, n_23040);
  not g51431 (n_23047, n31390);
  not g51432 (n_23048, n31391);
  and g51433 (n31392, n_23047, n_23048);
  not g51434 (n_23049, n31392);
  and g51435 (n31393, n_11971, n_23049);
  and g51436 (n31394, pi0609, n_22987);
  not g51437 (n_23050, n31394);
  and g51438 (n31395, n_11768, n_23050);
  not g51439 (n_23051, n31393);
  and g51440 (n31396, n_23051, n31395);
  and g51441 (n31397, n_11767, n_22995);
  not g51442 (n_23052, n31396);
  and g51443 (n31398, n_23052, n31397);
  and g51444 (n31399, pi0609, n_23049);
  and g51445 (n31400, n_11971, n_22987);
  not g51446 (n_23053, n31400);
  and g51447 (n31401, pi1155, n_23053);
  not g51448 (n_23054, n31399);
  and g51449 (n31402, n_23054, n31401);
  and g51450 (n31403, pi0660, n_22996);
  not g51451 (n_23055, n31402);
  and g51452 (n31404, n_23055, n31403);
  not g51453 (n_23056, n31398);
  not g51454 (n_23057, n31404);
  and g51455 (n31405, n_23056, n_23057);
  not g51456 (n_23058, n31405);
  and g51457 (n31406, pi0785, n_23058);
  and g51458 (n31407, n_11964, n_23049);
  not g51459 (n_23059, n31406);
  not g51460 (n_23060, n31407);
  and g51461 (n31408, n_23059, n_23060);
  not g51462 (n_23061, n31408);
  and g51463 (n31409, n_11984, n_23061);
  not g51464 (n_23062, n31377);
  and g51465 (n31410, n_11413, n_23062);
  not g51466 (n_23063, n31409);
  and g51467 (n31411, n_23063, n31410);
  and g51468 (n31412, n_11412, n_23003);
  not g51469 (n_23064, n31411);
  and g51470 (n31413, n_23064, n31412);
  and g51471 (n31414, n_11984, n31313);
  and g51472 (n31415, pi0618, n_23061);
  not g51473 (n_23065, n31414);
  and g51474 (n31416, pi1154, n_23065);
  not g51475 (n_23066, n31415);
  and g51476 (n31417, n_23066, n31416);
  and g51477 (n31418, pi0627, n_23004);
  not g51478 (n_23067, n31417);
  and g51479 (n31419, n_23067, n31418);
  not g51480 (n_23068, n31413);
  not g51481 (n_23069, n31419);
  and g51482 (n31420, n_23068, n_23069);
  not g51483 (n_23070, n31420);
  and g51484 (n31421, pi0781, n_23070);
  and g51485 (n31422, n_11981, n_23061);
  not g51486 (n_23071, n31421);
  not g51487 (n_23072, n31422);
  and g51488 (n31423, n_23071, n_23072);
  and g51489 (n31424, n_12315, n31423);
  not g51490 (n_23073, n31423);
  and g51491 (n31425, n_11821, n_23073);
  and g51492 (n31426, pi0619, n31314);
  not g51493 (n_23074, n31426);
  and g51494 (n31427, n_11405, n_23074);
  not g51495 (n_23075, n31425);
  and g51496 (n31428, n_23075, n31427);
  and g51497 (n31429, n_11403, n_23011);
  not g51498 (n_23076, n31428);
  and g51499 (n31430, n_23076, n31429);
  and g51500 (n31431, pi0619, n_23073);
  and g51501 (n31432, n_11821, n31314);
  not g51502 (n_23077, n31432);
  and g51503 (n31433, pi1159, n_23077);
  not g51504 (n_23078, n31431);
  and g51505 (n31434, n_23078, n31433);
  and g51506 (n31435, pi0648, n_23012);
  not g51507 (n_23079, n31434);
  and g51508 (n31436, n_23079, n31435);
  not g51509 (n_23080, n31430);
  and g51510 (n31437, pi0789, n_23080);
  not g51511 (n_23081, n31436);
  and g51512 (n31438, n_23081, n31437);
  not g51513 (n_23082, n31424);
  and g51514 (n31439, n17970, n_23082);
  not g51515 (n_23083, n31438);
  and g51516 (n31440, n_23083, n31439);
  not g51517 (n_23084, n31376);
  not g51518 (n_23085, n31440);
  and g51519 (n31441, n_23084, n_23085);
  not g51520 (n_23086, n31441);
  and g51521 (n31442, n_14638, n_23086);
  and g51522 (n31443, n17854, n_23018);
  and g51523 (n31444, n20851, n31316);
  not g51524 (n_23087, n31443);
  not g51525 (n_23088, n31444);
  and g51526 (n31445, n_23087, n_23088);
  not g51527 (n_23089, n31445);
  and g51528 (n31446, n_12354, n_23089);
  and g51529 (n31447, n20855, n31316);
  and g51530 (n31448, n17853, n_23018);
  not g51531 (n_23090, n31447);
  not g51532 (n_23091, n31448);
  and g51533 (n31449, n_23090, n_23091);
  not g51534 (n_23092, n31449);
  and g51535 (n31450, pi0629, n_23092);
  not g51536 (n_23093, n31446);
  not g51537 (n_23094, n31450);
  and g51538 (n31451, n_23093, n_23094);
  not g51539 (n_23095, n31451);
  and g51540 (n31452, pi0792, n_23095);
  not g51541 (n_23096, n31452);
  and g51542 (n31453, n_14387, n_23096);
  not g51543 (n_23097, n31442);
  and g51544 (n31454, n_23097, n31453);
  not g51545 (n_23098, n31364);
  not g51546 (n_23099, n31454);
  and g51547 (n31455, n_23098, n_23099);
  and g51548 (n31456, n_12411, n31455);
  and g51549 (n31457, n_11803, n_23021);
  and g51550 (n31458, pi1157, n_23024);
  not g51551 (n_23100, n31321);
  not g51552 (n_23101, n31458);
  and g51553 (n31459, n_23100, n_23101);
  not g51554 (n_23102, n31459);
  and g51555 (n31460, pi0787, n_23102);
  not g51556 (n_23103, n31457);
  not g51557 (n_23104, n31460);
  and g51558 (n31461, n_23103, n_23104);
  and g51559 (n31462, n_11819, n31461);
  and g51560 (n31463, pi0644, n31455);
  not g51561 (n_23105, n31462);
  and g51562 (n31464, pi0715, n_23105);
  not g51563 (n_23106, n31463);
  and g51564 (n31465, n_23106, n31464);
  not g51565 (n_23107, n31356);
  and g51566 (n31466, n_12392, n_23107);
  and g51567 (n31467, n17804, n31301);
  not g51568 (n_23108, n31466);
  not g51569 (n_23109, n31467);
  and g51570 (n31468, n_23108, n_23109);
  not g51571 (n_23110, n31468);
  and g51572 (n31469, pi0644, n_23110);
  and g51573 (n31470, n_11819, n31301);
  not g51574 (n_23111, n31470);
  and g51575 (n31471, n_12395, n_23111);
  not g51576 (n_23112, n31469);
  and g51577 (n31472, n_23112, n31471);
  not g51578 (n_23113, n31472);
  and g51579 (n31473, pi1160, n_23113);
  not g51580 (n_23114, n31465);
  and g51581 (n31474, n_23114, n31473);
  and g51582 (n31475, n_11819, n_23110);
  and g51583 (n31476, pi0644, n31301);
  not g51584 (n_23115, n31476);
  and g51585 (n31477, pi0715, n_23115);
  not g51586 (n_23116, n31475);
  and g51587 (n31478, n_23116, n31477);
  and g51588 (n31479, pi0644, n31461);
  and g51589 (n31480, n_11819, n31455);
  not g51590 (n_23117, n31479);
  and g51591 (n31481, n_12395, n_23117);
  not g51592 (n_23118, n31480);
  and g51593 (n31482, n_23118, n31481);
  not g51594 (n_23119, n31478);
  and g51595 (n31483, n_12405, n_23119);
  not g51596 (n_23120, n31482);
  and g51597 (n31484, n_23120, n31483);
  not g51598 (n_23121, n31474);
  not g51599 (n_23122, n31484);
  and g51600 (n31485, n_23121, n_23122);
  not g51601 (n_23123, n31485);
  and g51602 (n31486, pi0790, n_23123);
  not g51603 (n_23124, n31456);
  and g51604 (n31487, pi0832, n_23124);
  not g51605 (n_23125, n31486);
  and g51606 (n31488, n_23125, n31487);
  and g51607 (n31489, n_10720, po1038);
  and g51608 (n31490, n_10720, n_11751);
  not g51609 (n_23126, n31490);
  and g51610 (n31491, n16635, n_23126);
  and g51611 (n31492, pi0191, n_11417);
  and g51612 (n31493, n_10720, n_11418);
  not g51613 (n_23127, n31493);
  and g51614 (n31494, n16647, n_23127);
  and g51615 (n31495, n_10720, n18072);
  and g51616 (n31496, pi0191, n_12608);
  not g51617 (n_23128, n31496);
  and g51618 (n31497, n_161, n_23128);
  not g51619 (n_23129, n31495);
  and g51620 (n31498, n_23129, n31497);
  not g51621 (n_23130, n31494);
  and g51622 (n31499, pi0729, n_23130);
  not g51623 (n_23131, n31498);
  and g51624 (n31500, n_23131, n31499);
  and g51625 (n31501, n_10720, n_16056);
  and g51626 (n31502, n_11743, n31501);
  not g51627 (n_23132, n31502);
  and g51628 (n31503, n2571, n_23132);
  not g51629 (n_23133, n31500);
  and g51630 (n31504, n_23133, n31503);
  not g51631 (n_23134, n31492);
  not g51632 (n_23135, n31504);
  and g51633 (n31505, n_23134, n_23135);
  not g51634 (n_23136, n31505);
  and g51635 (n31506, n_11749, n_23136);
  and g51636 (n31507, n_11753, n31490);
  and g51637 (n31508, pi0625, n31505);
  not g51638 (n_23137, n31507);
  and g51639 (n31509, pi1153, n_23137);
  not g51640 (n_23138, n31508);
  and g51641 (n31510, n_23138, n31509);
  and g51642 (n31511, n_11753, n31505);
  and g51643 (n31512, pi0625, n31490);
  not g51644 (n_23139, n31512);
  and g51645 (n31513, n_11757, n_23139);
  not g51646 (n_23140, n31511);
  and g51647 (n31514, n_23140, n31513);
  not g51648 (n_23141, n31510);
  not g51649 (n_23142, n31514);
  and g51650 (n31515, n_23141, n_23142);
  not g51651 (n_23143, n31515);
  and g51652 (n31516, pi0778, n_23143);
  not g51653 (n_23144, n31506);
  not g51654 (n_23145, n31516);
  and g51655 (n31517, n_23144, n_23145);
  not g51656 (n_23146, n31517);
  and g51657 (n31518, n_11773, n_23146);
  and g51658 (n31519, n17075, n_23126);
  not g51659 (n_23147, n31518);
  not g51660 (n_23148, n31519);
  and g51661 (n31520, n_23147, n_23148);
  and g51662 (n31521, n_11777, n31520);
  and g51663 (n31522, n16639, n31490);
  not g51664 (n_23149, n31521);
  not g51665 (n_23150, n31522);
  and g51666 (n31523, n_23149, n_23150);
  and g51667 (n31524, n_11780, n31523);
  not g51668 (n_23151, n31491);
  not g51669 (n_23152, n31524);
  and g51670 (n31525, n_23151, n_23152);
  and g51671 (n31526, n_11783, n31525);
  and g51672 (n31527, n16631, n31490);
  not g51673 (n_23153, n31526);
  not g51674 (n_23154, n31527);
  and g51675 (n31528, n_23153, n_23154);
  not g51676 (n_23155, n31528);
  and g51677 (n31529, n_11789, n_23155);
  and g51678 (n31530, pi0628, n31490);
  not g51679 (n_23156, n31529);
  not g51680 (n_23157, n31530);
  and g51681 (n31531, n_23156, n_23157);
  not g51682 (n_23158, n31531);
  and g51683 (n31532, n_11794, n_23158);
  and g51684 (n31533, pi0628, n_23155);
  and g51685 (n31534, n_11789, n31490);
  not g51686 (n_23159, n31533);
  not g51687 (n_23160, n31534);
  and g51688 (n31535, n_23159, n_23160);
  not g51689 (n_23161, n31535);
  and g51690 (n31536, pi1156, n_23161);
  not g51691 (n_23162, n31532);
  not g51692 (n_23163, n31536);
  and g51693 (n31537, n_23162, n_23163);
  not g51694 (n_23164, n31537);
  and g51695 (n31538, pi0792, n_23164);
  and g51696 (n31539, n_11787, n_23155);
  not g51697 (n_23165, n31538);
  not g51698 (n_23166, n31539);
  and g51699 (n31540, n_23165, n_23166);
  not g51700 (n_23167, n31540);
  and g51701 (n31541, n_11806, n_23167);
  and g51702 (n31542, pi0647, n31490);
  not g51703 (n_23168, n31541);
  not g51704 (n_23169, n31542);
  and g51705 (n31543, n_23168, n_23169);
  not g51706 (n_23170, n31543);
  and g51707 (n31544, n_11810, n_23170);
  and g51708 (n31545, pi0647, n_23167);
  and g51709 (n31546, n_11806, n31490);
  not g51710 (n_23171, n31545);
  not g51711 (n_23172, n31546);
  and g51712 (n31547, n_23171, n_23172);
  not g51713 (n_23173, n31547);
  and g51714 (n31548, pi1157, n_23173);
  not g51715 (n_23174, n31544);
  not g51716 (n_23175, n31548);
  and g51717 (n31549, n_23174, n_23175);
  not g51718 (n_23176, n31549);
  and g51719 (n31550, pi0787, n_23176);
  and g51720 (n31551, n_11803, n_23167);
  not g51721 (n_23177, n31550);
  not g51722 (n_23178, n31551);
  and g51723 (n31552, n_23177, n_23178);
  not g51724 (n_23179, n31552);
  and g51725 (n31553, n_11819, n_23179);
  not g51726 (n_23180, n31553);
  and g51727 (n31554, pi0715, n_23180);
  and g51728 (n31555, n_16011, n17046);
  and g51729 (n31556, pi0191, n17273);
  not g51730 (n_23181, n31555);
  not g51731 (n_23182, n31556);
  and g51732 (n31557, n_23181, n_23182);
  not g51733 (n_23183, n31557);
  and g51734 (n31558, pi0039, n_23183);
  and g51735 (n31559, pi0746, n_11950);
  not g51736 (n_23184, n31559);
  and g51737 (n31560, pi0191, n_23184);
  and g51738 (n31561, n_10720, pi0746);
  and g51739 (n31562, n17221, n31561);
  not g51746 (n_23188, n31565);
  and g51747 (n31566, n_161, n_23188);
  and g51748 (n31567, pi0746, n17280);
  and g51749 (n31568, pi0038, n_23127);
  not g51750 (n_23189, n31567);
  and g51751 (n31569, n_23189, n31568);
  not g51752 (n_23190, n31566);
  not g51753 (n_23191, n31569);
  and g51754 (n31570, n_23190, n_23191);
  not g51755 (n_23192, n31570);
  and g51756 (n31571, n2571, n_23192);
  not g51757 (n_23193, n31571);
  and g51758 (n31572, n_23134, n_23193);
  not g51759 (n_23194, n31572);
  and g51760 (n31573, n_11960, n_23194);
  and g51761 (n31574, n17117, n_23126);
  not g51762 (n_23195, n31573);
  not g51763 (n_23196, n31574);
  and g51764 (n31575, n_23195, n_23196);
  not g51765 (n_23197, n31575);
  and g51766 (n31576, n_11964, n_23197);
  and g51767 (n31577, n_11967, n_23126);
  and g51768 (n31578, pi0609, n31573);
  not g51769 (n_23198, n31577);
  not g51770 (n_23199, n31578);
  and g51771 (n31579, n_23198, n_23199);
  not g51772 (n_23200, n31579);
  and g51773 (n31580, pi1155, n_23200);
  and g51774 (n31581, n_11972, n_23126);
  and g51775 (n31582, n_11971, n31573);
  not g51776 (n_23201, n31581);
  not g51777 (n_23202, n31582);
  and g51778 (n31583, n_23201, n_23202);
  not g51779 (n_23203, n31583);
  and g51780 (n31584, n_11768, n_23203);
  not g51781 (n_23204, n31580);
  not g51782 (n_23205, n31584);
  and g51783 (n31585, n_23204, n_23205);
  not g51784 (n_23206, n31585);
  and g51785 (n31586, pi0785, n_23206);
  not g51786 (n_23207, n31576);
  not g51787 (n_23208, n31586);
  and g51788 (n31587, n_23207, n_23208);
  not g51789 (n_23209, n31587);
  and g51790 (n31588, n_11981, n_23209);
  and g51791 (n31589, n_11984, n31490);
  and g51792 (n31590, pi0618, n31587);
  not g51793 (n_23210, n31589);
  and g51794 (n31591, pi1154, n_23210);
  not g51795 (n_23211, n31590);
  and g51796 (n31592, n_23211, n31591);
  and g51797 (n31593, n_11984, n31587);
  and g51798 (n31594, pi0618, n31490);
  not g51799 (n_23212, n31594);
  and g51800 (n31595, n_11413, n_23212);
  not g51801 (n_23213, n31593);
  and g51802 (n31596, n_23213, n31595);
  not g51803 (n_23214, n31592);
  not g51804 (n_23215, n31596);
  and g51805 (n31597, n_23214, n_23215);
  not g51806 (n_23216, n31597);
  and g51807 (n31598, pi0781, n_23216);
  not g51808 (n_23217, n31588);
  not g51809 (n_23218, n31598);
  and g51810 (n31599, n_23217, n_23218);
  not g51811 (n_23219, n31599);
  and g51812 (n31600, n_12315, n_23219);
  and g51813 (n31601, n_11821, n31490);
  and g51814 (n31602, pi0619, n31599);
  not g51815 (n_23220, n31601);
  and g51816 (n31603, pi1159, n_23220);
  not g51817 (n_23221, n31602);
  and g51818 (n31604, n_23221, n31603);
  and g51819 (n31605, n_11821, n31599);
  and g51820 (n31606, pi0619, n31490);
  not g51821 (n_23222, n31606);
  and g51822 (n31607, n_11405, n_23222);
  not g51823 (n_23223, n31605);
  and g51824 (n31608, n_23223, n31607);
  not g51825 (n_23224, n31604);
  not g51826 (n_23225, n31608);
  and g51827 (n31609, n_23224, n_23225);
  not g51828 (n_23226, n31609);
  and g51829 (n31610, pi0789, n_23226);
  not g51830 (n_23227, n31600);
  not g51831 (n_23228, n31610);
  and g51832 (n31611, n_23227, n_23228);
  and g51833 (n31612, n_12524, n31611);
  and g51834 (n31613, n17969, n31490);
  not g51835 (n_23229, n31612);
  not g51836 (n_23230, n31613);
  and g51837 (n31614, n_23229, n_23230);
  not g51838 (n_23231, n31614);
  and g51839 (n31615, n_12368, n_23231);
  and g51840 (n31616, n17779, n31490);
  not g51841 (n_23232, n31615);
  not g51842 (n_23233, n31616);
  and g51843 (n31617, n_23232, n_23233);
  not g51844 (n_23234, n31617);
  and g51845 (n31618, n_12392, n_23234);
  and g51846 (n31619, n17804, n31490);
  not g51847 (n_23235, n31618);
  not g51848 (n_23236, n31619);
  and g51849 (n31620, n_23235, n_23236);
  not g51850 (n_23237, n31620);
  and g51851 (n31621, pi0644, n_23237);
  and g51852 (n31622, n_11819, n31490);
  not g51853 (n_23238, n31622);
  and g51854 (n31623, n_12395, n_23238);
  not g51855 (n_23239, n31621);
  and g51856 (n31624, n_23239, n31623);
  not g51857 (n_23240, n31624);
  and g51858 (n31625, pi1160, n_23240);
  not g51859 (n_23241, n31554);
  and g51860 (n31626, n_23241, n31625);
  and g51861 (n31627, pi0644, n_23179);
  not g51862 (n_23242, n31627);
  and g51863 (n31628, n_12395, n_23242);
  and g51864 (n31629, n_11819, n_23237);
  and g51865 (n31630, pi0644, n31490);
  not g51866 (n_23243, n31630);
  and g51867 (n31631, pi0715, n_23243);
  not g51868 (n_23244, n31629);
  and g51869 (n31632, n_23244, n31631);
  not g51870 (n_23245, n31632);
  and g51871 (n31633, n_12405, n_23245);
  not g51872 (n_23246, n31628);
  and g51873 (n31634, n_23246, n31633);
  not g51874 (n_23247, n31626);
  not g51875 (n_23248, n31634);
  and g51876 (n31635, n_23247, n_23248);
  not g51877 (n_23249, n31635);
  and g51878 (n31636, pi0790, n_23249);
  and g51879 (n31637, n17777, n31531);
  and g51880 (n31638, n_14557, n31614);
  and g51881 (n31639, n17776, n31535);
  not g51882 (n_23250, n31637);
  not g51883 (n_23251, n31639);
  and g51884 (n31640, n_23250, n_23251);
  not g51885 (n_23252, n31638);
  and g51886 (n31641, n_23252, n31640);
  not g51887 (n_23253, n31641);
  and g51888 (n31642, pi0792, n_23253);
  and g51889 (n31643, pi0609, n31517);
  and g51890 (n31644, n_16056, n31570);
  and g51891 (n31645, n_16011, n24055);
  not g51892 (n_23254, n31645);
  and g51893 (n31646, n_12250, n_23254);
  not g51894 (n_23255, n31646);
  and g51895 (n31647, n_162, n_23255);
  not g51896 (n_23256, n31647);
  and g51897 (n31648, n_10720, n_23256);
  and g51898 (n31649, n_12120, n_22990);
  not g51899 (n_23257, n31649);
  and g51900 (n31650, pi0191, n_23257);
  and g51901 (n31651, n6284, n31650);
  not g51902 (n_23258, n31651);
  and g51903 (n31652, pi0038, n_23258);
  not g51904 (n_23259, n31648);
  and g51905 (n31653, n_23259, n31652);
  and g51906 (n31654, n_10720, n_12694);
  and g51907 (n31655, pi0191, n_12695);
  not g51908 (n_23260, n31655);
  and g51909 (n31656, pi0746, n_23260);
  not g51910 (n_23261, n31654);
  and g51911 (n31657, n_23261, n31656);
  and g51912 (n31658, n_10720, n17612);
  and g51913 (n31659, pi0191, n17625);
  not g51914 (n_23262, n31658);
  and g51915 (n31660, n_16011, n_23262);
  not g51916 (n_23263, n31659);
  and g51917 (n31661, n_23263, n31660);
  not g51918 (n_23264, n31657);
  and g51919 (n31662, n_162, n_23264);
  not g51920 (n_23265, n31661);
  and g51921 (n31663, n_23265, n31662);
  and g51922 (n31664, pi0191, n17605);
  and g51923 (n31665, n_10720, n_12180);
  not g51924 (n_23266, n31665);
  and g51925 (n31666, pi0746, n_23266);
  not g51926 (n_23267, n31664);
  and g51927 (n31667, n_23267, n31666);
  and g51928 (n31668, n_10720, n17404);
  and g51929 (n31669, pi0191, n17485);
  not g51930 (n_23268, n31669);
  and g51931 (n31670, n_16011, n_23268);
  not g51932 (n_23269, n31668);
  and g51933 (n31671, n_23269, n31670);
  not g51934 (n_23270, n31667);
  and g51935 (n31672, pi0039, n_23270);
  not g51936 (n_23271, n31671);
  and g51937 (n31673, n_23271, n31672);
  not g51938 (n_23272, n31663);
  and g51939 (n31674, n_161, n_23272);
  not g51940 (n_23273, n31673);
  and g51941 (n31675, n_23273, n31674);
  not g51942 (n_23274, n31653);
  and g51943 (n31676, pi0729, n_23274);
  not g51944 (n_23275, n31675);
  and g51945 (n31677, n_23275, n31676);
  not g51946 (n_23276, n31677);
  and g51947 (n31678, n2571, n_23276);
  not g51948 (n_23277, n31644);
  and g51949 (n31679, n_23277, n31678);
  not g51950 (n_23278, n31679);
  and g51951 (n31680, n_23134, n_23278);
  and g51952 (n31681, n_11753, n31680);
  and g51953 (n31682, pi0625, n31572);
  not g51954 (n_23279, n31682);
  and g51955 (n31683, n_11757, n_23279);
  not g51956 (n_23280, n31681);
  and g51957 (n31684, n_23280, n31683);
  and g51958 (n31685, n_11823, n_23141);
  not g51959 (n_23281, n31684);
  and g51960 (n31686, n_23281, n31685);
  and g51961 (n31687, n_11753, n31572);
  and g51962 (n31688, pi0625, n31680);
  not g51963 (n_23282, n31687);
  and g51964 (n31689, pi1153, n_23282);
  not g51965 (n_23283, n31688);
  and g51966 (n31690, n_23283, n31689);
  and g51967 (n31691, pi0608, n_23142);
  not g51968 (n_23284, n31690);
  and g51969 (n31692, n_23284, n31691);
  not g51970 (n_23285, n31686);
  not g51971 (n_23286, n31692);
  and g51972 (n31693, n_23285, n_23286);
  not g51973 (n_23287, n31693);
  and g51974 (n31694, pi0778, n_23287);
  and g51975 (n31695, n_11749, n31680);
  not g51976 (n_23288, n31694);
  not g51977 (n_23289, n31695);
  and g51978 (n31696, n_23288, n_23289);
  not g51979 (n_23290, n31696);
  and g51980 (n31697, n_11971, n_23290);
  not g51981 (n_23291, n31643);
  and g51982 (n31698, n_11768, n_23291);
  not g51983 (n_23292, n31697);
  and g51984 (n31699, n_23292, n31698);
  and g51985 (n31700, n_11767, n_23204);
  not g51986 (n_23293, n31699);
  and g51987 (n31701, n_23293, n31700);
  and g51988 (n31702, n_11971, n31517);
  and g51989 (n31703, pi0609, n_23290);
  not g51990 (n_23294, n31702);
  and g51991 (n31704, pi1155, n_23294);
  not g51992 (n_23295, n31703);
  and g51993 (n31705, n_23295, n31704);
  and g51994 (n31706, pi0660, n_23205);
  not g51995 (n_23296, n31705);
  and g51996 (n31707, n_23296, n31706);
  not g51997 (n_23297, n31701);
  not g51998 (n_23298, n31707);
  and g51999 (n31708, n_23297, n_23298);
  not g52000 (n_23299, n31708);
  and g52001 (n31709, pi0785, n_23299);
  and g52002 (n31710, n_11964, n_23290);
  not g52003 (n_23300, n31709);
  not g52004 (n_23301, n31710);
  and g52005 (n31711, n_23300, n_23301);
  not g52006 (n_23302, n31711);
  and g52007 (n31712, n_11984, n_23302);
  and g52008 (n31713, pi0618, n31520);
  not g52009 (n_23303, n31713);
  and g52010 (n31714, n_11413, n_23303);
  not g52011 (n_23304, n31712);
  and g52012 (n31715, n_23304, n31714);
  and g52013 (n31716, n_11412, n_23214);
  not g52014 (n_23305, n31715);
  and g52015 (n31717, n_23305, n31716);
  and g52016 (n31718, n_11984, n31520);
  and g52017 (n31719, pi0618, n_23302);
  not g52018 (n_23306, n31718);
  and g52019 (n31720, pi1154, n_23306);
  not g52020 (n_23307, n31719);
  and g52021 (n31721, n_23307, n31720);
  and g52022 (n31722, pi0627, n_23215);
  not g52023 (n_23308, n31721);
  and g52024 (n31723, n_23308, n31722);
  not g52025 (n_23309, n31717);
  not g52026 (n_23310, n31723);
  and g52027 (n31724, n_23309, n_23310);
  not g52028 (n_23311, n31724);
  and g52029 (n31725, pi0781, n_23311);
  and g52030 (n31726, n_11981, n_23302);
  not g52031 (n_23312, n31725);
  not g52032 (n_23313, n31726);
  and g52033 (n31727, n_23312, n_23313);
  and g52034 (n31728, n_12315, n31727);
  not g52035 (n_23314, n31523);
  and g52036 (n31729, pi0619, n_23314);
  not g52037 (n_23315, n31727);
  and g52038 (n31730, n_11821, n_23315);
  not g52039 (n_23316, n31729);
  and g52040 (n31731, n_11405, n_23316);
  not g52041 (n_23317, n31730);
  and g52042 (n31732, n_23317, n31731);
  and g52043 (n31733, n_11403, n_23224);
  not g52044 (n_23318, n31732);
  and g52045 (n31734, n_23318, n31733);
  and g52046 (n31735, n_11821, n_23314);
  and g52047 (n31736, pi0619, n_23315);
  not g52048 (n_23319, n31735);
  and g52049 (n31737, pi1159, n_23319);
  not g52050 (n_23320, n31736);
  and g52051 (n31738, n_23320, n31737);
  and g52052 (n31739, pi0648, n_23225);
  not g52053 (n_23321, n31738);
  and g52054 (n31740, n_23321, n31739);
  not g52055 (n_23322, n31734);
  and g52056 (n31741, pi0789, n_23322);
  not g52057 (n_23323, n31740);
  and g52058 (n31742, n_23323, n31741);
  not g52059 (n_23324, n31728);
  and g52060 (n31743, n17970, n_23324);
  not g52061 (n_23325, n31742);
  and g52062 (n31744, n_23325, n31743);
  and g52063 (n31745, n17871, n31525);
  not g52064 (n_23326, n31611);
  and g52065 (n31746, n_12320, n_23326);
  and g52066 (n31747, pi0626, n_23126);
  not g52067 (n_23327, n31747);
  and g52068 (n31748, n16629, n_23327);
  not g52069 (n_23328, n31746);
  and g52070 (n31749, n_23328, n31748);
  and g52071 (n31750, pi0626, n_23326);
  and g52072 (n31751, n_12320, n_23126);
  not g52073 (n_23329, n31751);
  and g52074 (n31752, n16628, n_23329);
  not g52075 (n_23330, n31750);
  and g52076 (n31753, n_23330, n31752);
  not g52077 (n_23331, n31745);
  not g52078 (n_23332, n31749);
  and g52079 (n31754, n_23331, n_23332);
  not g52080 (n_23333, n31753);
  and g52081 (n31755, n_23333, n31754);
  not g52082 (n_23334, n31755);
  and g52083 (n31756, pi0788, n_23334);
  not g52084 (n_23335, n31756);
  and g52085 (n31757, n_14638, n_23335);
  not g52086 (n_23336, n31744);
  and g52087 (n31758, n_23336, n31757);
  not g52088 (n_23337, n31642);
  not g52089 (n_23338, n31758);
  and g52090 (n31759, n_23337, n_23338);
  not g52091 (n_23339, n31759);
  and g52092 (n31760, n_14387, n_23339);
  and g52093 (n31761, n17802, n31543);
  and g52094 (n31762, n_14548, n31617);
  and g52095 (n31763, n17801, n31547);
  not g52096 (n_23340, n31761);
  not g52097 (n_23341, n31762);
  and g52098 (n31764, n_23340, n_23341);
  not g52099 (n_23342, n31763);
  and g52100 (n31765, n_23342, n31764);
  not g52101 (n_23343, n31765);
  and g52102 (n31766, pi0787, n_23343);
  and g52103 (n31767, n_11819, n31633);
  and g52104 (n31768, pi0644, n31625);
  not g52105 (n_23344, n31767);
  and g52106 (n31769, pi0790, n_23344);
  not g52107 (n_23345, n31768);
  and g52108 (n31770, n_23345, n31769);
  not g52109 (n_23346, n31760);
  not g52110 (n_23347, n31766);
  and g52111 (n31771, n_23346, n_23347);
  not g52112 (n_23348, n31770);
  and g52113 (n31772, n_23348, n31771);
  not g52114 (n_23349, n31636);
  not g52115 (n_23350, n31772);
  and g52116 (n31773, n_23349, n_23350);
  not g52117 (n_23351, n31773);
  and g52118 (n31774, n_4226, n_23351);
  not g52119 (n_23352, n31489);
  and g52120 (n31775, n_12415, n_23352);
  not g52121 (n_23353, n31774);
  and g52122 (n31776, n_23353, n31775);
  not g52123 (n_23354, n31488);
  not g52124 (n_23355, n31776);
  and g52125 (po0348, n_23354, n_23355);
  and g52126 (n31778, n_11043, n_12418);
  and g52127 (n31779, pi0691, n16645);
  not g52128 (n_23356, n31778);
  not g52129 (n_23357, n31779);
  and g52130 (n31780, n_23356, n_23357);
  not g52131 (n_23358, n31780);
  and g52132 (n31781, n_11749, n_23358);
  and g52133 (n31782, n_11753, n31779);
  not g52134 (n_23359, n31782);
  and g52135 (n31783, n_23358, n_23359);
  not g52136 (n_23360, n31783);
  and g52137 (n31784, pi1153, n_23360);
  and g52138 (n31785, n_11757, n_23356);
  and g52139 (n31786, n_23359, n31785);
  not g52140 (n_23361, n31786);
  and g52141 (n31787, pi0778, n_23361);
  not g52142 (n_23362, n31784);
  and g52143 (n31788, n_23362, n31787);
  not g52144 (n_23363, n31781);
  not g52145 (n_23364, n31788);
  and g52146 (n31789, n_23363, n_23364);
  not g52147 (n_23365, n31789);
  and g52148 (n31790, n_12429, n_23365);
  and g52149 (n31791, n_12430, n31790);
  and g52150 (n31792, n_12431, n31791);
  and g52151 (n31793, n_12432, n31792);
  and g52152 (n31794, n_12436, n31793);
  and g52153 (n31795, n_11806, n31794);
  and g52154 (n31796, pi0647, n31778);
  not g52155 (n_23366, n31796);
  and g52156 (n31797, n_11810, n_23366);
  not g52157 (n_23367, n31795);
  and g52158 (n31798, n_23367, n31797);
  and g52159 (n31799, pi0630, n31798);
  and g52160 (n31800, pi0764, n17244);
  not g52161 (n_23368, n31800);
  and g52162 (n31801, n_23356, n_23368);
  not g52163 (n_23369, n31801);
  and g52164 (n31802, n_12448, n_23369);
  not g52165 (n_23370, n31802);
  and g52166 (n31803, n_11964, n_23370);
  and g52167 (n31804, n17296, n31800);
  not g52168 (n_23371, n31804);
  and g52169 (n31805, n31802, n_23371);
  not g52170 (n_23372, n31805);
  and g52171 (n31806, pi1155, n_23372);
  and g52172 (n31807, n_11768, n_23356);
  and g52173 (n31808, n_23371, n31807);
  not g52174 (n_23373, n31806);
  not g52175 (n_23374, n31808);
  and g52176 (n31809, n_23373, n_23374);
  not g52177 (n_23375, n31809);
  and g52178 (n31810, pi0785, n_23375);
  not g52179 (n_23376, n31803);
  not g52180 (n_23377, n31810);
  and g52181 (n31811, n_23376, n_23377);
  not g52182 (n_23378, n31811);
  and g52183 (n31812, n_11981, n_23378);
  and g52184 (n31813, n_12461, n31811);
  not g52185 (n_23379, n31813);
  and g52186 (n31814, pi1154, n_23379);
  and g52187 (n31815, n_12463, n31811);
  not g52188 (n_23380, n31815);
  and g52189 (n31816, n_11413, n_23380);
  not g52190 (n_23381, n31814);
  not g52191 (n_23382, n31816);
  and g52192 (n31817, n_23381, n_23382);
  not g52193 (n_23383, n31817);
  and g52194 (n31818, pi0781, n_23383);
  not g52195 (n_23384, n31812);
  not g52196 (n_23385, n31818);
  and g52197 (n31819, n_23384, n_23385);
  not g52198 (n_23386, n31819);
  and g52199 (n31820, n_12315, n_23386);
  and g52200 (n31821, n_16503, n31819);
  not g52201 (n_23387, n31821);
  and g52202 (n31822, pi1159, n_23387);
  and g52203 (n31823, n_16505, n31819);
  not g52204 (n_23388, n31823);
  and g52205 (n31824, n_11405, n_23388);
  not g52206 (n_23389, n31822);
  not g52207 (n_23390, n31824);
  and g52208 (n31825, n_23389, n_23390);
  not g52209 (n_23391, n31825);
  and g52210 (n31826, pi0789, n_23391);
  not g52211 (n_23392, n31820);
  not g52212 (n_23393, n31826);
  and g52213 (n31827, n_23392, n_23393);
  and g52214 (n31828, n_12524, n31827);
  and g52215 (n31829, n17969, n31778);
  not g52216 (n_23394, n31828);
  not g52217 (n_23395, n31829);
  and g52218 (n31830, n_23394, n_23395);
  not g52219 (n_23396, n31830);
  and g52220 (n31831, n_12368, n_23396);
  and g52221 (n31832, n17779, n31778);
  not g52222 (n_23397, n31831);
  not g52223 (n_23398, n31832);
  and g52224 (n31833, n_23397, n_23398);
  and g52225 (n31834, n_14548, n31833);
  not g52226 (n_23399, n31794);
  and g52227 (n31835, pi0647, n_23399);
  and g52228 (n31836, n_11806, n_23356);
  not g52229 (n_23400, n31835);
  not g52230 (n_23401, n31836);
  and g52231 (n31837, n_23400, n_23401);
  not g52232 (n_23402, n31837);
  and g52233 (n31838, n17801, n_23402);
  not g52234 (n_23403, n31799);
  not g52235 (n_23404, n31838);
  and g52236 (n31839, n_23403, n_23404);
  not g52237 (n_23405, n31834);
  and g52238 (n31840, n_23405, n31839);
  not g52239 (n_23406, n31840);
  and g52240 (n31841, pi0787, n_23406);
  and g52241 (n31842, n17871, n31792);
  not g52242 (n_23407, n31827);
  and g52243 (n31843, n_12320, n_23407);
  and g52244 (n31844, pi0626, n_23356);
  not g52245 (n_23408, n31844);
  and g52246 (n31845, n16629, n_23408);
  not g52247 (n_23409, n31843);
  and g52248 (n31846, n_23409, n31845);
  and g52249 (n31847, pi0626, n_23407);
  and g52250 (n31848, n_12320, n_23356);
  not g52251 (n_23410, n31848);
  and g52252 (n31849, n16628, n_23410);
  not g52253 (n_23411, n31847);
  and g52254 (n31850, n_23411, n31849);
  not g52255 (n_23412, n31842);
  not g52256 (n_23413, n31846);
  and g52257 (n31851, n_23412, n_23413);
  not g52258 (n_23414, n31850);
  and g52259 (n31852, n_23414, n31851);
  not g52260 (n_23415, n31852);
  and g52261 (n31853, pi0788, n_23415);
  and g52262 (n31854, pi0618, n31790);
  and g52263 (n31855, n_11866, n_23358);
  and g52264 (n31856, pi0625, n31855);
  not g52265 (n_23416, n31855);
  and g52266 (n31857, n31801, n_23416);
  not g52267 (n_23417, n31856);
  not g52268 (n_23418, n31857);
  and g52269 (n31858, n_23417, n_23418);
  not g52270 (n_23419, n31858);
  and g52271 (n31859, n31785, n_23419);
  and g52272 (n31860, n_11823, n_23362);
  not g52273 (n_23420, n31859);
  and g52274 (n31861, n_23420, n31860);
  and g52275 (n31862, pi1153, n31801);
  and g52276 (n31863, n_23417, n31862);
  and g52277 (n31864, pi0608, n_23361);
  not g52278 (n_23421, n31863);
  and g52279 (n31865, n_23421, n31864);
  not g52280 (n_23422, n31861);
  not g52281 (n_23423, n31865);
  and g52282 (n31866, n_23422, n_23423);
  not g52283 (n_23424, n31866);
  and g52284 (n31867, pi0778, n_23424);
  and g52285 (n31868, n_11749, n_23418);
  not g52286 (n_23425, n31867);
  not g52287 (n_23426, n31868);
  and g52288 (n31869, n_23425, n_23426);
  not g52289 (n_23427, n31869);
  and g52290 (n31870, n_11971, n_23427);
  and g52291 (n31871, pi0609, n_23365);
  not g52292 (n_23428, n31871);
  and g52293 (n31872, n_11768, n_23428);
  not g52294 (n_23429, n31870);
  and g52295 (n31873, n_23429, n31872);
  and g52296 (n31874, n_11767, n_23373);
  not g52297 (n_23430, n31873);
  and g52298 (n31875, n_23430, n31874);
  and g52299 (n31876, pi0609, n_23427);
  and g52300 (n31877, n_11971, n_23365);
  not g52301 (n_23431, n31877);
  and g52302 (n31878, pi1155, n_23431);
  not g52303 (n_23432, n31876);
  and g52304 (n31879, n_23432, n31878);
  and g52305 (n31880, pi0660, n_23374);
  not g52306 (n_23433, n31879);
  and g52307 (n31881, n_23433, n31880);
  not g52308 (n_23434, n31875);
  not g52309 (n_23435, n31881);
  and g52310 (n31882, n_23434, n_23435);
  not g52311 (n_23436, n31882);
  and g52312 (n31883, pi0785, n_23436);
  and g52313 (n31884, n_11964, n_23427);
  not g52314 (n_23437, n31883);
  not g52315 (n_23438, n31884);
  and g52316 (n31885, n_23437, n_23438);
  not g52317 (n_23439, n31885);
  and g52318 (n31886, n_11984, n_23439);
  not g52319 (n_23440, n31854);
  and g52320 (n31887, n_11413, n_23440);
  not g52321 (n_23441, n31886);
  and g52322 (n31888, n_23441, n31887);
  and g52323 (n31889, n_11412, n_23381);
  not g52324 (n_23442, n31888);
  and g52325 (n31890, n_23442, n31889);
  and g52326 (n31891, n_11984, n31790);
  and g52327 (n31892, pi0618, n_23439);
  not g52328 (n_23443, n31891);
  and g52329 (n31893, pi1154, n_23443);
  not g52330 (n_23444, n31892);
  and g52331 (n31894, n_23444, n31893);
  and g52332 (n31895, pi0627, n_23382);
  not g52333 (n_23445, n31894);
  and g52334 (n31896, n_23445, n31895);
  not g52335 (n_23446, n31890);
  not g52336 (n_23447, n31896);
  and g52337 (n31897, n_23446, n_23447);
  not g52338 (n_23448, n31897);
  and g52339 (n31898, pi0781, n_23448);
  and g52340 (n31899, n_11981, n_23439);
  not g52341 (n_23449, n31898);
  not g52342 (n_23450, n31899);
  and g52343 (n31900, n_23449, n_23450);
  and g52344 (n31901, n_12315, n31900);
  not g52345 (n_23451, n31900);
  and g52346 (n31902, n_11821, n_23451);
  and g52347 (n31903, pi0619, n31791);
  not g52348 (n_23452, n31903);
  and g52349 (n31904, n_11405, n_23452);
  not g52350 (n_23453, n31902);
  and g52351 (n31905, n_23453, n31904);
  and g52352 (n31906, n_11403, n_23389);
  not g52353 (n_23454, n31905);
  and g52354 (n31907, n_23454, n31906);
  and g52355 (n31908, pi0619, n_23451);
  and g52356 (n31909, n_11821, n31791);
  not g52357 (n_23455, n31909);
  and g52358 (n31910, pi1159, n_23455);
  not g52359 (n_23456, n31908);
  and g52360 (n31911, n_23456, n31910);
  and g52361 (n31912, pi0648, n_23390);
  not g52362 (n_23457, n31911);
  and g52363 (n31913, n_23457, n31912);
  not g52364 (n_23458, n31907);
  and g52365 (n31914, pi0789, n_23458);
  not g52366 (n_23459, n31913);
  and g52367 (n31915, n_23459, n31914);
  not g52368 (n_23460, n31901);
  and g52369 (n31916, n17970, n_23460);
  not g52370 (n_23461, n31915);
  and g52371 (n31917, n_23461, n31916);
  not g52372 (n_23462, n31853);
  not g52373 (n_23463, n31917);
  and g52374 (n31918, n_23462, n_23463);
  not g52375 (n_23464, n31918);
  and g52376 (n31919, n_14638, n_23464);
  and g52377 (n31920, n17854, n_23396);
  and g52378 (n31921, n20851, n31793);
  not g52379 (n_23465, n31920);
  not g52380 (n_23466, n31921);
  and g52381 (n31922, n_23465, n_23466);
  not g52382 (n_23467, n31922);
  and g52383 (n31923, n_12354, n_23467);
  and g52384 (n31924, n20855, n31793);
  and g52385 (n31925, n17853, n_23396);
  not g52386 (n_23468, n31924);
  not g52387 (n_23469, n31925);
  and g52388 (n31926, n_23468, n_23469);
  not g52389 (n_23470, n31926);
  and g52390 (n31927, pi0629, n_23470);
  not g52391 (n_23471, n31923);
  not g52392 (n_23472, n31927);
  and g52393 (n31928, n_23471, n_23472);
  not g52394 (n_23473, n31928);
  and g52395 (n31929, pi0792, n_23473);
  not g52396 (n_23474, n31929);
  and g52397 (n31930, n_14387, n_23474);
  not g52398 (n_23475, n31919);
  and g52399 (n31931, n_23475, n31930);
  not g52400 (n_23476, n31841);
  not g52401 (n_23477, n31931);
  and g52402 (n31932, n_23476, n_23477);
  and g52403 (n31933, n_12411, n31932);
  and g52404 (n31934, n_11803, n_23399);
  and g52405 (n31935, pi1157, n_23402);
  not g52406 (n_23478, n31798);
  not g52407 (n_23479, n31935);
  and g52408 (n31936, n_23478, n_23479);
  not g52409 (n_23480, n31936);
  and g52410 (n31937, pi0787, n_23480);
  not g52411 (n_23481, n31934);
  not g52412 (n_23482, n31937);
  and g52413 (n31938, n_23481, n_23482);
  and g52414 (n31939, n_11819, n31938);
  and g52415 (n31940, pi0644, n31932);
  not g52416 (n_23483, n31939);
  and g52417 (n31941, pi0715, n_23483);
  not g52418 (n_23484, n31940);
  and g52419 (n31942, n_23484, n31941);
  not g52420 (n_23485, n31833);
  and g52421 (n31943, n_12392, n_23485);
  and g52422 (n31944, n17804, n31778);
  not g52423 (n_23486, n31943);
  not g52424 (n_23487, n31944);
  and g52425 (n31945, n_23486, n_23487);
  not g52426 (n_23488, n31945);
  and g52427 (n31946, pi0644, n_23488);
  and g52428 (n31947, n_11819, n31778);
  not g52429 (n_23489, n31947);
  and g52430 (n31948, n_12395, n_23489);
  not g52431 (n_23490, n31946);
  and g52432 (n31949, n_23490, n31948);
  not g52433 (n_23491, n31949);
  and g52434 (n31950, pi1160, n_23491);
  not g52435 (n_23492, n31942);
  and g52436 (n31951, n_23492, n31950);
  and g52437 (n31952, n_11819, n_23488);
  and g52438 (n31953, pi0644, n31778);
  not g52439 (n_23493, n31953);
  and g52440 (n31954, pi0715, n_23493);
  not g52441 (n_23494, n31952);
  and g52442 (n31955, n_23494, n31954);
  and g52443 (n31956, pi0644, n31938);
  and g52444 (n31957, n_11819, n31932);
  not g52445 (n_23495, n31956);
  and g52446 (n31958, n_12395, n_23495);
  not g52447 (n_23496, n31957);
  and g52448 (n31959, n_23496, n31958);
  not g52449 (n_23497, n31955);
  and g52450 (n31960, n_12405, n_23497);
  not g52451 (n_23498, n31959);
  and g52452 (n31961, n_23498, n31960);
  not g52453 (n_23499, n31951);
  not g52454 (n_23500, n31961);
  and g52455 (n31962, n_23499, n_23500);
  not g52456 (n_23501, n31962);
  and g52457 (n31963, pi0790, n_23501);
  not g52458 (n_23502, n31933);
  and g52459 (n31964, pi0832, n_23502);
  not g52460 (n_23503, n31963);
  and g52461 (n31965, n_23503, n31964);
  and g52462 (n31966, n_11043, po1038);
  and g52463 (n31967, n_11043, n_11751);
  not g52464 (n_23504, n31967);
  and g52465 (n31968, n16635, n_23504);
  and g52466 (n31969, pi0192, n_11417);
  and g52467 (n31970, n_11043, n_11418);
  not g52468 (n_23505, n31970);
  and g52469 (n31971, n16647, n_23505);
  and g52470 (n31972, n_11043, n18072);
  and g52471 (n31973, pi0192, n_12608);
  not g52472 (n_23506, n31973);
  and g52473 (n31974, n_161, n_23506);
  not g52474 (n_23507, n31972);
  and g52475 (n31975, n_23507, n31974);
  not g52476 (n_23508, n31971);
  and g52477 (n31976, pi0691, n_23508);
  not g52478 (n_23509, n31975);
  and g52479 (n31977, n_23509, n31976);
  and g52480 (n31978, n_11043, n_16177);
  and g52481 (n31979, n_11743, n31978);
  not g52482 (n_23510, n31979);
  and g52483 (n31980, n2571, n_23510);
  not g52484 (n_23511, n31977);
  and g52485 (n31981, n_23511, n31980);
  not g52486 (n_23512, n31969);
  not g52487 (n_23513, n31981);
  and g52488 (n31982, n_23512, n_23513);
  not g52489 (n_23514, n31982);
  and g52490 (n31983, n_11749, n_23514);
  and g52491 (n31984, n_11753, n31967);
  and g52492 (n31985, pi0625, n31982);
  not g52493 (n_23515, n31984);
  and g52494 (n31986, pi1153, n_23515);
  not g52495 (n_23516, n31985);
  and g52496 (n31987, n_23516, n31986);
  and g52497 (n31988, n_11753, n31982);
  and g52498 (n31989, pi0625, n31967);
  not g52499 (n_23517, n31989);
  and g52500 (n31990, n_11757, n_23517);
  not g52501 (n_23518, n31988);
  and g52502 (n31991, n_23518, n31990);
  not g52503 (n_23519, n31987);
  not g52504 (n_23520, n31991);
  and g52505 (n31992, n_23519, n_23520);
  not g52506 (n_23521, n31992);
  and g52507 (n31993, pi0778, n_23521);
  not g52508 (n_23522, n31983);
  not g52509 (n_23523, n31993);
  and g52510 (n31994, n_23522, n_23523);
  not g52511 (n_23524, n31994);
  and g52512 (n31995, n_11773, n_23524);
  and g52513 (n31996, n17075, n_23504);
  not g52514 (n_23525, n31995);
  not g52515 (n_23526, n31996);
  and g52516 (n31997, n_23525, n_23526);
  and g52517 (n31998, n_11777, n31997);
  and g52518 (n31999, n16639, n31967);
  not g52519 (n_23527, n31998);
  not g52520 (n_23528, n31999);
  and g52521 (n32000, n_23527, n_23528);
  and g52522 (n32001, n_11780, n32000);
  not g52523 (n_23529, n31968);
  not g52524 (n_23530, n32001);
  and g52525 (n32002, n_23529, n_23530);
  and g52526 (n32003, n_11783, n32002);
  and g52527 (n32004, n16631, n31967);
  not g52528 (n_23531, n32003);
  not g52529 (n_23532, n32004);
  and g52530 (n32005, n_23531, n_23532);
  not g52531 (n_23533, n32005);
  and g52532 (n32006, n_11789, n_23533);
  and g52533 (n32007, pi0628, n31967);
  not g52534 (n_23534, n32006);
  not g52535 (n_23535, n32007);
  and g52536 (n32008, n_23534, n_23535);
  not g52537 (n_23536, n32008);
  and g52538 (n32009, n_11794, n_23536);
  and g52539 (n32010, pi0628, n_23533);
  and g52540 (n32011, n_11789, n31967);
  not g52541 (n_23537, n32010);
  not g52542 (n_23538, n32011);
  and g52543 (n32012, n_23537, n_23538);
  not g52544 (n_23539, n32012);
  and g52545 (n32013, pi1156, n_23539);
  not g52546 (n_23540, n32009);
  not g52547 (n_23541, n32013);
  and g52548 (n32014, n_23540, n_23541);
  not g52549 (n_23542, n32014);
  and g52550 (n32015, pi0792, n_23542);
  and g52551 (n32016, n_11787, n_23533);
  not g52552 (n_23543, n32015);
  not g52553 (n_23544, n32016);
  and g52554 (n32017, n_23543, n_23544);
  not g52555 (n_23545, n32017);
  and g52556 (n32018, n_11806, n_23545);
  and g52557 (n32019, pi0647, n31967);
  not g52558 (n_23546, n32018);
  not g52559 (n_23547, n32019);
  and g52560 (n32020, n_23546, n_23547);
  not g52561 (n_23548, n32020);
  and g52562 (n32021, n_11810, n_23548);
  and g52563 (n32022, pi0647, n_23545);
  and g52564 (n32023, n_11806, n31967);
  not g52565 (n_23549, n32022);
  not g52566 (n_23550, n32023);
  and g52567 (n32024, n_23549, n_23550);
  not g52568 (n_23551, n32024);
  and g52569 (n32025, pi1157, n_23551);
  not g52570 (n_23552, n32021);
  not g52571 (n_23553, n32025);
  and g52572 (n32026, n_23552, n_23553);
  not g52573 (n_23554, n32026);
  and g52574 (n32027, pi0787, n_23554);
  and g52575 (n32028, n_11803, n_23545);
  not g52576 (n_23555, n32027);
  not g52577 (n_23556, n32028);
  and g52578 (n32029, n_23555, n_23556);
  not g52579 (n_23557, n32029);
  and g52580 (n32030, n_11819, n_23557);
  not g52581 (n_23558, n32030);
  and g52582 (n32031, pi0715, n_23558);
  and g52583 (n32032, n_16132, n17046);
  and g52584 (n32033, pi0192, n17273);
  not g52585 (n_23559, n32032);
  not g52586 (n_23560, n32033);
  and g52587 (n32034, n_23559, n_23560);
  not g52588 (n_23561, n32034);
  and g52589 (n32035, pi0039, n_23561);
  and g52590 (n32036, pi0764, n_11950);
  not g52591 (n_23562, n32036);
  and g52592 (n32037, pi0192, n_23562);
  and g52593 (n32038, n_11043, pi0764);
  and g52594 (n32039, n17221, n32038);
  not g52601 (n_23566, n32042);
  and g52602 (n32043, n_161, n_23566);
  and g52603 (n32044, pi0764, n17280);
  and g52604 (n32045, pi0038, n_23505);
  not g52605 (n_23567, n32044);
  and g52606 (n32046, n_23567, n32045);
  not g52607 (n_23568, n32043);
  not g52608 (n_23569, n32046);
  and g52609 (n32047, n_23568, n_23569);
  not g52610 (n_23570, n32047);
  and g52611 (n32048, n2571, n_23570);
  not g52612 (n_23571, n32048);
  and g52613 (n32049, n_23512, n_23571);
  not g52614 (n_23572, n32049);
  and g52615 (n32050, n_11960, n_23572);
  and g52616 (n32051, n17117, n_23504);
  not g52617 (n_23573, n32050);
  not g52618 (n_23574, n32051);
  and g52619 (n32052, n_23573, n_23574);
  not g52620 (n_23575, n32052);
  and g52621 (n32053, n_11964, n_23575);
  and g52622 (n32054, n_11967, n_23504);
  and g52623 (n32055, pi0609, n32050);
  not g52624 (n_23576, n32054);
  not g52625 (n_23577, n32055);
  and g52626 (n32056, n_23576, n_23577);
  not g52627 (n_23578, n32056);
  and g52628 (n32057, pi1155, n_23578);
  and g52629 (n32058, n_11972, n_23504);
  and g52630 (n32059, n_11971, n32050);
  not g52631 (n_23579, n32058);
  not g52632 (n_23580, n32059);
  and g52633 (n32060, n_23579, n_23580);
  not g52634 (n_23581, n32060);
  and g52635 (n32061, n_11768, n_23581);
  not g52636 (n_23582, n32057);
  not g52637 (n_23583, n32061);
  and g52638 (n32062, n_23582, n_23583);
  not g52639 (n_23584, n32062);
  and g52640 (n32063, pi0785, n_23584);
  not g52641 (n_23585, n32053);
  not g52642 (n_23586, n32063);
  and g52643 (n32064, n_23585, n_23586);
  not g52644 (n_23587, n32064);
  and g52645 (n32065, n_11981, n_23587);
  and g52646 (n32066, n_11984, n31967);
  and g52647 (n32067, pi0618, n32064);
  not g52648 (n_23588, n32066);
  and g52649 (n32068, pi1154, n_23588);
  not g52650 (n_23589, n32067);
  and g52651 (n32069, n_23589, n32068);
  and g52652 (n32070, n_11984, n32064);
  and g52653 (n32071, pi0618, n31967);
  not g52654 (n_23590, n32071);
  and g52655 (n32072, n_11413, n_23590);
  not g52656 (n_23591, n32070);
  and g52657 (n32073, n_23591, n32072);
  not g52658 (n_23592, n32069);
  not g52659 (n_23593, n32073);
  and g52660 (n32074, n_23592, n_23593);
  not g52661 (n_23594, n32074);
  and g52662 (n32075, pi0781, n_23594);
  not g52663 (n_23595, n32065);
  not g52664 (n_23596, n32075);
  and g52665 (n32076, n_23595, n_23596);
  not g52666 (n_23597, n32076);
  and g52667 (n32077, n_12315, n_23597);
  and g52668 (n32078, n_11821, n31967);
  and g52669 (n32079, pi0619, n32076);
  not g52670 (n_23598, n32078);
  and g52671 (n32080, pi1159, n_23598);
  not g52672 (n_23599, n32079);
  and g52673 (n32081, n_23599, n32080);
  and g52674 (n32082, n_11821, n32076);
  and g52675 (n32083, pi0619, n31967);
  not g52676 (n_23600, n32083);
  and g52677 (n32084, n_11405, n_23600);
  not g52678 (n_23601, n32082);
  and g52679 (n32085, n_23601, n32084);
  not g52680 (n_23602, n32081);
  not g52681 (n_23603, n32085);
  and g52682 (n32086, n_23602, n_23603);
  not g52683 (n_23604, n32086);
  and g52684 (n32087, pi0789, n_23604);
  not g52685 (n_23605, n32077);
  not g52686 (n_23606, n32087);
  and g52687 (n32088, n_23605, n_23606);
  and g52688 (n32089, n_12524, n32088);
  and g52689 (n32090, n17969, n31967);
  not g52690 (n_23607, n32089);
  not g52691 (n_23608, n32090);
  and g52692 (n32091, n_23607, n_23608);
  not g52693 (n_23609, n32091);
  and g52694 (n32092, n_12368, n_23609);
  and g52695 (n32093, n17779, n31967);
  not g52696 (n_23610, n32092);
  not g52697 (n_23611, n32093);
  and g52698 (n32094, n_23610, n_23611);
  not g52699 (n_23612, n32094);
  and g52700 (n32095, n_12392, n_23612);
  and g52701 (n32096, n17804, n31967);
  not g52702 (n_23613, n32095);
  not g52703 (n_23614, n32096);
  and g52704 (n32097, n_23613, n_23614);
  not g52705 (n_23615, n32097);
  and g52706 (n32098, pi0644, n_23615);
  and g52707 (n32099, n_11819, n31967);
  not g52708 (n_23616, n32099);
  and g52709 (n32100, n_12395, n_23616);
  not g52710 (n_23617, n32098);
  and g52711 (n32101, n_23617, n32100);
  not g52712 (n_23618, n32101);
  and g52713 (n32102, pi1160, n_23618);
  not g52714 (n_23619, n32031);
  and g52715 (n32103, n_23619, n32102);
  and g52716 (n32104, pi0644, n_23557);
  not g52717 (n_23620, n32104);
  and g52718 (n32105, n_12395, n_23620);
  and g52719 (n32106, n_11819, n_23615);
  and g52720 (n32107, pi0644, n31967);
  not g52721 (n_23621, n32107);
  and g52722 (n32108, pi0715, n_23621);
  not g52723 (n_23622, n32106);
  and g52724 (n32109, n_23622, n32108);
  not g52725 (n_23623, n32109);
  and g52726 (n32110, n_12405, n_23623);
  not g52727 (n_23624, n32105);
  and g52728 (n32111, n_23624, n32110);
  not g52729 (n_23625, n32103);
  not g52730 (n_23626, n32111);
  and g52731 (n32112, n_23625, n_23626);
  not g52732 (n_23627, n32112);
  and g52733 (n32113, pi0790, n_23627);
  and g52734 (n32114, n17777, n32008);
  and g52735 (n32115, n_14557, n32091);
  and g52736 (n32116, n17776, n32012);
  not g52737 (n_23628, n32114);
  not g52738 (n_23629, n32116);
  and g52739 (n32117, n_23628, n_23629);
  not g52740 (n_23630, n32115);
  and g52741 (n32118, n_23630, n32117);
  not g52742 (n_23631, n32118);
  and g52743 (n32119, pi0792, n_23631);
  and g52744 (n32120, pi0609, n31994);
  and g52745 (n32121, n_16177, n32047);
  and g52746 (n32122, n_16132, n24055);
  not g52747 (n_23632, n32122);
  and g52748 (n32123, n_12250, n_23632);
  not g52749 (n_23633, n32123);
  and g52750 (n32124, n_162, n_23633);
  not g52751 (n_23634, n32124);
  and g52752 (n32125, n_11043, n_23634);
  and g52753 (n32126, n_12120, n_23368);
  not g52754 (n_23635, n32126);
  and g52755 (n32127, pi0192, n_23635);
  and g52756 (n32128, n6284, n32127);
  not g52757 (n_23636, n32128);
  and g52758 (n32129, pi0038, n_23636);
  not g52759 (n_23637, n32125);
  and g52760 (n32130, n_23637, n32129);
  and g52761 (n32131, n_11043, n_12694);
  and g52762 (n32132, pi0192, n_12695);
  not g52763 (n_23638, n32132);
  and g52764 (n32133, pi0764, n_23638);
  not g52765 (n_23639, n32131);
  and g52766 (n32134, n_23639, n32133);
  and g52767 (n32135, n_11043, n17612);
  and g52768 (n32136, pi0192, n17625);
  not g52769 (n_23640, n32135);
  and g52770 (n32137, n_16132, n_23640);
  not g52771 (n_23641, n32136);
  and g52772 (n32138, n_23641, n32137);
  not g52773 (n_23642, n32134);
  and g52774 (n32139, n_162, n_23642);
  not g52775 (n_23643, n32138);
  and g52776 (n32140, n_23643, n32139);
  and g52777 (n32141, pi0192, n17605);
  and g52778 (n32142, n_11043, n_12180);
  not g52779 (n_23644, n32142);
  and g52780 (n32143, pi0764, n_23644);
  not g52781 (n_23645, n32141);
  and g52782 (n32144, n_23645, n32143);
  and g52783 (n32145, n_11043, n17404);
  and g52784 (n32146, pi0192, n17485);
  not g52785 (n_23646, n32146);
  and g52786 (n32147, n_16132, n_23646);
  not g52787 (n_23647, n32145);
  and g52788 (n32148, n_23647, n32147);
  not g52789 (n_23648, n32144);
  and g52790 (n32149, pi0039, n_23648);
  not g52791 (n_23649, n32148);
  and g52792 (n32150, n_23649, n32149);
  not g52793 (n_23650, n32140);
  and g52794 (n32151, n_161, n_23650);
  not g52795 (n_23651, n32150);
  and g52796 (n32152, n_23651, n32151);
  not g52797 (n_23652, n32130);
  and g52798 (n32153, pi0691, n_23652);
  not g52799 (n_23653, n32152);
  and g52800 (n32154, n_23653, n32153);
  not g52801 (n_23654, n32154);
  and g52802 (n32155, n2571, n_23654);
  not g52803 (n_23655, n32121);
  and g52804 (n32156, n_23655, n32155);
  not g52805 (n_23656, n32156);
  and g52806 (n32157, n_23512, n_23656);
  and g52807 (n32158, n_11753, n32157);
  and g52808 (n32159, pi0625, n32049);
  not g52809 (n_23657, n32159);
  and g52810 (n32160, n_11757, n_23657);
  not g52811 (n_23658, n32158);
  and g52812 (n32161, n_23658, n32160);
  and g52813 (n32162, n_11823, n_23519);
  not g52814 (n_23659, n32161);
  and g52815 (n32163, n_23659, n32162);
  and g52816 (n32164, n_11753, n32049);
  and g52817 (n32165, pi0625, n32157);
  not g52818 (n_23660, n32164);
  and g52819 (n32166, pi1153, n_23660);
  not g52820 (n_23661, n32165);
  and g52821 (n32167, n_23661, n32166);
  and g52822 (n32168, pi0608, n_23520);
  not g52823 (n_23662, n32167);
  and g52824 (n32169, n_23662, n32168);
  not g52825 (n_23663, n32163);
  not g52826 (n_23664, n32169);
  and g52827 (n32170, n_23663, n_23664);
  not g52828 (n_23665, n32170);
  and g52829 (n32171, pi0778, n_23665);
  and g52830 (n32172, n_11749, n32157);
  not g52831 (n_23666, n32171);
  not g52832 (n_23667, n32172);
  and g52833 (n32173, n_23666, n_23667);
  not g52834 (n_23668, n32173);
  and g52835 (n32174, n_11971, n_23668);
  not g52836 (n_23669, n32120);
  and g52837 (n32175, n_11768, n_23669);
  not g52838 (n_23670, n32174);
  and g52839 (n32176, n_23670, n32175);
  and g52840 (n32177, n_11767, n_23582);
  not g52841 (n_23671, n32176);
  and g52842 (n32178, n_23671, n32177);
  and g52843 (n32179, n_11971, n31994);
  and g52844 (n32180, pi0609, n_23668);
  not g52845 (n_23672, n32179);
  and g52846 (n32181, pi1155, n_23672);
  not g52847 (n_23673, n32180);
  and g52848 (n32182, n_23673, n32181);
  and g52849 (n32183, pi0660, n_23583);
  not g52850 (n_23674, n32182);
  and g52851 (n32184, n_23674, n32183);
  not g52852 (n_23675, n32178);
  not g52853 (n_23676, n32184);
  and g52854 (n32185, n_23675, n_23676);
  not g52855 (n_23677, n32185);
  and g52856 (n32186, pi0785, n_23677);
  and g52857 (n32187, n_11964, n_23668);
  not g52858 (n_23678, n32186);
  not g52859 (n_23679, n32187);
  and g52860 (n32188, n_23678, n_23679);
  not g52861 (n_23680, n32188);
  and g52862 (n32189, n_11984, n_23680);
  and g52863 (n32190, pi0618, n31997);
  not g52864 (n_23681, n32190);
  and g52865 (n32191, n_11413, n_23681);
  not g52866 (n_23682, n32189);
  and g52867 (n32192, n_23682, n32191);
  and g52868 (n32193, n_11412, n_23592);
  not g52869 (n_23683, n32192);
  and g52870 (n32194, n_23683, n32193);
  and g52871 (n32195, n_11984, n31997);
  and g52872 (n32196, pi0618, n_23680);
  not g52873 (n_23684, n32195);
  and g52874 (n32197, pi1154, n_23684);
  not g52875 (n_23685, n32196);
  and g52876 (n32198, n_23685, n32197);
  and g52877 (n32199, pi0627, n_23593);
  not g52878 (n_23686, n32198);
  and g52879 (n32200, n_23686, n32199);
  not g52880 (n_23687, n32194);
  not g52881 (n_23688, n32200);
  and g52882 (n32201, n_23687, n_23688);
  not g52883 (n_23689, n32201);
  and g52884 (n32202, pi0781, n_23689);
  and g52885 (n32203, n_11981, n_23680);
  not g52886 (n_23690, n32202);
  not g52887 (n_23691, n32203);
  and g52888 (n32204, n_23690, n_23691);
  and g52889 (n32205, n_12315, n32204);
  not g52890 (n_23692, n32000);
  and g52891 (n32206, pi0619, n_23692);
  not g52892 (n_23693, n32204);
  and g52893 (n32207, n_11821, n_23693);
  not g52894 (n_23694, n32206);
  and g52895 (n32208, n_11405, n_23694);
  not g52896 (n_23695, n32207);
  and g52897 (n32209, n_23695, n32208);
  and g52898 (n32210, n_11403, n_23602);
  not g52899 (n_23696, n32209);
  and g52900 (n32211, n_23696, n32210);
  and g52901 (n32212, n_11821, n_23692);
  and g52902 (n32213, pi0619, n_23693);
  not g52903 (n_23697, n32212);
  and g52904 (n32214, pi1159, n_23697);
  not g52905 (n_23698, n32213);
  and g52906 (n32215, n_23698, n32214);
  and g52907 (n32216, pi0648, n_23603);
  not g52908 (n_23699, n32215);
  and g52909 (n32217, n_23699, n32216);
  not g52910 (n_23700, n32211);
  and g52911 (n32218, pi0789, n_23700);
  not g52912 (n_23701, n32217);
  and g52913 (n32219, n_23701, n32218);
  not g52914 (n_23702, n32205);
  and g52915 (n32220, n17970, n_23702);
  not g52916 (n_23703, n32219);
  and g52917 (n32221, n_23703, n32220);
  and g52918 (n32222, n17871, n32002);
  not g52919 (n_23704, n32088);
  and g52920 (n32223, n_12320, n_23704);
  and g52921 (n32224, pi0626, n_23504);
  not g52922 (n_23705, n32224);
  and g52923 (n32225, n16629, n_23705);
  not g52924 (n_23706, n32223);
  and g52925 (n32226, n_23706, n32225);
  and g52926 (n32227, pi0626, n_23704);
  and g52927 (n32228, n_12320, n_23504);
  not g52928 (n_23707, n32228);
  and g52929 (n32229, n16628, n_23707);
  not g52930 (n_23708, n32227);
  and g52931 (n32230, n_23708, n32229);
  not g52932 (n_23709, n32222);
  not g52933 (n_23710, n32226);
  and g52934 (n32231, n_23709, n_23710);
  not g52935 (n_23711, n32230);
  and g52936 (n32232, n_23711, n32231);
  not g52937 (n_23712, n32232);
  and g52938 (n32233, pi0788, n_23712);
  not g52939 (n_23713, n32233);
  and g52940 (n32234, n_14638, n_23713);
  not g52941 (n_23714, n32221);
  and g52942 (n32235, n_23714, n32234);
  not g52943 (n_23715, n32119);
  not g52944 (n_23716, n32235);
  and g52945 (n32236, n_23715, n_23716);
  not g52946 (n_23717, n32236);
  and g52947 (n32237, n_14387, n_23717);
  and g52948 (n32238, n17802, n32020);
  and g52949 (n32239, n_14548, n32094);
  and g52950 (n32240, n17801, n32024);
  not g52951 (n_23718, n32238);
  not g52952 (n_23719, n32239);
  and g52953 (n32241, n_23718, n_23719);
  not g52954 (n_23720, n32240);
  and g52955 (n32242, n_23720, n32241);
  not g52956 (n_23721, n32242);
  and g52957 (n32243, pi0787, n_23721);
  and g52958 (n32244, n_11819, n32110);
  and g52959 (n32245, pi0644, n32102);
  not g52960 (n_23722, n32244);
  and g52961 (n32246, pi0790, n_23722);
  not g52962 (n_23723, n32245);
  and g52963 (n32247, n_23723, n32246);
  not g52964 (n_23724, n32237);
  not g52965 (n_23725, n32243);
  and g52966 (n32248, n_23724, n_23725);
  not g52967 (n_23726, n32247);
  and g52968 (n32249, n_23726, n32248);
  not g52969 (n_23727, n32113);
  not g52970 (n_23728, n32249);
  and g52971 (n32250, n_23727, n_23728);
  not g52972 (n_23729, n32250);
  and g52973 (n32251, n_4226, n_23729);
  not g52974 (n_23730, n31966);
  and g52975 (n32252, n_12415, n_23730);
  not g52976 (n_23731, n32251);
  and g52977 (n32253, n_23731, n32252);
  not g52978 (n_23732, n31965);
  not g52979 (n_23733, n32253);
  and g52980 (po0349, n_23732, n_23733);
  and g52981 (n32255, n_5790, n_12418);
  and g52982 (n32256, pi0690, n16645);
  not g52983 (n_23734, n32255);
  not g52984 (n_23735, n32256);
  and g52985 (n32257, n_23734, n_23735);
  not g52986 (n_23736, n32257);
  and g52987 (n32258, n_11749, n_23736);
  and g52988 (n32259, n_11753, n32256);
  not g52989 (n_23737, n32259);
  and g52990 (n32260, n_23736, n_23737);
  not g52991 (n_23738, n32260);
  and g52992 (n32261, pi1153, n_23738);
  and g52993 (n32262, n_11757, n_23734);
  and g52994 (n32263, n_23737, n32262);
  not g52995 (n_23739, n32263);
  and g52996 (n32264, pi0778, n_23739);
  not g52997 (n_23740, n32261);
  and g52998 (n32265, n_23740, n32264);
  not g52999 (n_23741, n32258);
  not g53000 (n_23742, n32265);
  and g53001 (n32266, n_23741, n_23742);
  not g53002 (n_23743, n32266);
  and g53003 (n32267, n_12429, n_23743);
  and g53004 (n32268, n_12430, n32267);
  and g53005 (n32269, n_12431, n32268);
  and g53006 (n32270, n_12432, n32269);
  and g53007 (n32271, n_12436, n32270);
  and g53008 (n32272, n_11806, n32271);
  and g53009 (n32273, pi0647, n32255);
  not g53010 (n_23744, n32273);
  and g53011 (n32274, n_11810, n_23744);
  not g53012 (n_23745, n32272);
  and g53013 (n32275, n_23745, n32274);
  and g53014 (n32276, pi0630, n32275);
  and g53015 (n32277, pi0739, n17244);
  not g53016 (n_23746, n32277);
  and g53017 (n32278, n_23734, n_23746);
  not g53018 (n_23747, n32278);
  and g53019 (n32279, n_12448, n_23747);
  not g53020 (n_23748, n32279);
  and g53021 (n32280, n_11964, n_23748);
  and g53022 (n32281, n17296, n32277);
  not g53023 (n_23749, n32281);
  and g53024 (n32282, n32279, n_23749);
  not g53025 (n_23750, n32282);
  and g53026 (n32283, pi1155, n_23750);
  and g53027 (n32284, n_11768, n_23734);
  and g53028 (n32285, n_23749, n32284);
  not g53029 (n_23751, n32283);
  not g53030 (n_23752, n32285);
  and g53031 (n32286, n_23751, n_23752);
  not g53032 (n_23753, n32286);
  and g53033 (n32287, pi0785, n_23753);
  not g53034 (n_23754, n32280);
  not g53035 (n_23755, n32287);
  and g53036 (n32288, n_23754, n_23755);
  not g53037 (n_23756, n32288);
  and g53038 (n32289, n_11981, n_23756);
  and g53039 (n32290, n_12461, n32288);
  not g53040 (n_23757, n32290);
  and g53041 (n32291, pi1154, n_23757);
  and g53042 (n32292, n_12463, n32288);
  not g53043 (n_23758, n32292);
  and g53044 (n32293, n_11413, n_23758);
  not g53045 (n_23759, n32291);
  not g53046 (n_23760, n32293);
  and g53047 (n32294, n_23759, n_23760);
  not g53048 (n_23761, n32294);
  and g53049 (n32295, pi0781, n_23761);
  not g53050 (n_23762, n32289);
  not g53051 (n_23763, n32295);
  and g53052 (n32296, n_23762, n_23763);
  not g53053 (n_23764, n32296);
  and g53054 (n32297, n_12315, n_23764);
  and g53055 (n32298, n_16503, n32296);
  not g53056 (n_23765, n32298);
  and g53057 (n32299, pi1159, n_23765);
  and g53058 (n32300, n_16505, n32296);
  not g53059 (n_23766, n32300);
  and g53060 (n32301, n_11405, n_23766);
  not g53061 (n_23767, n32299);
  not g53062 (n_23768, n32301);
  and g53063 (n32302, n_23767, n_23768);
  not g53064 (n_23769, n32302);
  and g53065 (n32303, pi0789, n_23769);
  not g53066 (n_23770, n32297);
  not g53067 (n_23771, n32303);
  and g53068 (n32304, n_23770, n_23771);
  and g53069 (n32305, n_12524, n32304);
  and g53070 (n32306, n17969, n32255);
  not g53071 (n_23772, n32305);
  not g53072 (n_23773, n32306);
  and g53073 (n32307, n_23772, n_23773);
  not g53074 (n_23774, n32307);
  and g53075 (n32308, n_12368, n_23774);
  and g53076 (n32309, n17779, n32255);
  not g53077 (n_23775, n32308);
  not g53078 (n_23776, n32309);
  and g53079 (n32310, n_23775, n_23776);
  and g53080 (n32311, n_14548, n32310);
  not g53081 (n_23777, n32271);
  and g53082 (n32312, pi0647, n_23777);
  and g53083 (n32313, n_11806, n_23734);
  not g53084 (n_23778, n32312);
  not g53085 (n_23779, n32313);
  and g53086 (n32314, n_23778, n_23779);
  not g53087 (n_23780, n32314);
  and g53088 (n32315, n17801, n_23780);
  not g53089 (n_23781, n32276);
  not g53090 (n_23782, n32315);
  and g53091 (n32316, n_23781, n_23782);
  not g53092 (n_23783, n32311);
  and g53093 (n32317, n_23783, n32316);
  not g53094 (n_23784, n32317);
  and g53095 (n32318, pi0787, n_23784);
  and g53096 (n32319, n17871, n32269);
  not g53097 (n_23785, n32304);
  and g53098 (n32320, n_12320, n_23785);
  and g53099 (n32321, pi0626, n_23734);
  not g53100 (n_23786, n32321);
  and g53101 (n32322, n16629, n_23786);
  not g53102 (n_23787, n32320);
  and g53103 (n32323, n_23787, n32322);
  and g53104 (n32324, pi0626, n_23785);
  and g53105 (n32325, n_12320, n_23734);
  not g53106 (n_23788, n32325);
  and g53107 (n32326, n16628, n_23788);
  not g53108 (n_23789, n32324);
  and g53109 (n32327, n_23789, n32326);
  not g53110 (n_23790, n32319);
  not g53111 (n_23791, n32323);
  and g53112 (n32328, n_23790, n_23791);
  not g53113 (n_23792, n32327);
  and g53114 (n32329, n_23792, n32328);
  not g53115 (n_23793, n32329);
  and g53116 (n32330, pi0788, n_23793);
  and g53117 (n32331, pi0618, n32267);
  and g53118 (n32332, n_11866, n_23736);
  and g53119 (n32333, pi0625, n32332);
  not g53120 (n_23794, n32332);
  and g53121 (n32334, n32278, n_23794);
  not g53122 (n_23795, n32333);
  not g53123 (n_23796, n32334);
  and g53124 (n32335, n_23795, n_23796);
  not g53125 (n_23797, n32335);
  and g53126 (n32336, n32262, n_23797);
  and g53127 (n32337, n_11823, n_23740);
  not g53128 (n_23798, n32336);
  and g53129 (n32338, n_23798, n32337);
  and g53130 (n32339, pi1153, n32278);
  and g53131 (n32340, n_23795, n32339);
  and g53132 (n32341, pi0608, n_23739);
  not g53133 (n_23799, n32340);
  and g53134 (n32342, n_23799, n32341);
  not g53135 (n_23800, n32338);
  not g53136 (n_23801, n32342);
  and g53137 (n32343, n_23800, n_23801);
  not g53138 (n_23802, n32343);
  and g53139 (n32344, pi0778, n_23802);
  and g53140 (n32345, n_11749, n_23796);
  not g53141 (n_23803, n32344);
  not g53142 (n_23804, n32345);
  and g53143 (n32346, n_23803, n_23804);
  not g53144 (n_23805, n32346);
  and g53145 (n32347, n_11971, n_23805);
  and g53146 (n32348, pi0609, n_23743);
  not g53147 (n_23806, n32348);
  and g53148 (n32349, n_11768, n_23806);
  not g53149 (n_23807, n32347);
  and g53150 (n32350, n_23807, n32349);
  and g53151 (n32351, n_11767, n_23751);
  not g53152 (n_23808, n32350);
  and g53153 (n32352, n_23808, n32351);
  and g53154 (n32353, pi0609, n_23805);
  and g53155 (n32354, n_11971, n_23743);
  not g53156 (n_23809, n32354);
  and g53157 (n32355, pi1155, n_23809);
  not g53158 (n_23810, n32353);
  and g53159 (n32356, n_23810, n32355);
  and g53160 (n32357, pi0660, n_23752);
  not g53161 (n_23811, n32356);
  and g53162 (n32358, n_23811, n32357);
  not g53163 (n_23812, n32352);
  not g53164 (n_23813, n32358);
  and g53165 (n32359, n_23812, n_23813);
  not g53166 (n_23814, n32359);
  and g53167 (n32360, pi0785, n_23814);
  and g53168 (n32361, n_11964, n_23805);
  not g53169 (n_23815, n32360);
  not g53170 (n_23816, n32361);
  and g53171 (n32362, n_23815, n_23816);
  not g53172 (n_23817, n32362);
  and g53173 (n32363, n_11984, n_23817);
  not g53174 (n_23818, n32331);
  and g53175 (n32364, n_11413, n_23818);
  not g53176 (n_23819, n32363);
  and g53177 (n32365, n_23819, n32364);
  and g53178 (n32366, n_11412, n_23759);
  not g53179 (n_23820, n32365);
  and g53180 (n32367, n_23820, n32366);
  and g53181 (n32368, n_11984, n32267);
  and g53182 (n32369, pi0618, n_23817);
  not g53183 (n_23821, n32368);
  and g53184 (n32370, pi1154, n_23821);
  not g53185 (n_23822, n32369);
  and g53186 (n32371, n_23822, n32370);
  and g53187 (n32372, pi0627, n_23760);
  not g53188 (n_23823, n32371);
  and g53189 (n32373, n_23823, n32372);
  not g53190 (n_23824, n32367);
  not g53191 (n_23825, n32373);
  and g53192 (n32374, n_23824, n_23825);
  not g53193 (n_23826, n32374);
  and g53194 (n32375, pi0781, n_23826);
  and g53195 (n32376, n_11981, n_23817);
  not g53196 (n_23827, n32375);
  not g53197 (n_23828, n32376);
  and g53198 (n32377, n_23827, n_23828);
  and g53199 (n32378, n_12315, n32377);
  not g53200 (n_23829, n32377);
  and g53201 (n32379, n_11821, n_23829);
  and g53202 (n32380, pi0619, n32268);
  not g53203 (n_23830, n32380);
  and g53204 (n32381, n_11405, n_23830);
  not g53205 (n_23831, n32379);
  and g53206 (n32382, n_23831, n32381);
  and g53207 (n32383, n_11403, n_23767);
  not g53208 (n_23832, n32382);
  and g53209 (n32384, n_23832, n32383);
  and g53210 (n32385, pi0619, n_23829);
  and g53211 (n32386, n_11821, n32268);
  not g53212 (n_23833, n32386);
  and g53213 (n32387, pi1159, n_23833);
  not g53214 (n_23834, n32385);
  and g53215 (n32388, n_23834, n32387);
  and g53216 (n32389, pi0648, n_23768);
  not g53217 (n_23835, n32388);
  and g53218 (n32390, n_23835, n32389);
  not g53219 (n_23836, n32384);
  and g53220 (n32391, pi0789, n_23836);
  not g53221 (n_23837, n32390);
  and g53222 (n32392, n_23837, n32391);
  not g53223 (n_23838, n32378);
  and g53224 (n32393, n17970, n_23838);
  not g53225 (n_23839, n32392);
  and g53226 (n32394, n_23839, n32393);
  not g53227 (n_23840, n32330);
  not g53228 (n_23841, n32394);
  and g53229 (n32395, n_23840, n_23841);
  not g53230 (n_23842, n32395);
  and g53231 (n32396, n_14638, n_23842);
  and g53232 (n32397, n17854, n_23774);
  and g53233 (n32398, n20851, n32270);
  not g53234 (n_23843, n32397);
  not g53235 (n_23844, n32398);
  and g53236 (n32399, n_23843, n_23844);
  not g53237 (n_23845, n32399);
  and g53238 (n32400, n_12354, n_23845);
  and g53239 (n32401, n20855, n32270);
  and g53240 (n32402, n17853, n_23774);
  not g53241 (n_23846, n32401);
  not g53242 (n_23847, n32402);
  and g53243 (n32403, n_23846, n_23847);
  not g53244 (n_23848, n32403);
  and g53245 (n32404, pi0629, n_23848);
  not g53246 (n_23849, n32400);
  not g53247 (n_23850, n32404);
  and g53248 (n32405, n_23849, n_23850);
  not g53249 (n_23851, n32405);
  and g53250 (n32406, pi0792, n_23851);
  not g53251 (n_23852, n32406);
  and g53252 (n32407, n_14387, n_23852);
  not g53253 (n_23853, n32396);
  and g53254 (n32408, n_23853, n32407);
  not g53255 (n_23854, n32318);
  not g53256 (n_23855, n32408);
  and g53257 (n32409, n_23854, n_23855);
  and g53258 (n32410, n_12411, n32409);
  and g53259 (n32411, n_11803, n_23777);
  and g53260 (n32412, pi1157, n_23780);
  not g53261 (n_23856, n32275);
  not g53262 (n_23857, n32412);
  and g53263 (n32413, n_23856, n_23857);
  not g53264 (n_23858, n32413);
  and g53265 (n32414, pi0787, n_23858);
  not g53266 (n_23859, n32411);
  not g53267 (n_23860, n32414);
  and g53268 (n32415, n_23859, n_23860);
  and g53269 (n32416, n_11819, n32415);
  and g53270 (n32417, pi0644, n32409);
  not g53271 (n_23861, n32416);
  and g53272 (n32418, pi0715, n_23861);
  not g53273 (n_23862, n32417);
  and g53274 (n32419, n_23862, n32418);
  not g53275 (n_23863, n32310);
  and g53276 (n32420, n_12392, n_23863);
  and g53277 (n32421, n17804, n32255);
  not g53278 (n_23864, n32420);
  not g53279 (n_23865, n32421);
  and g53280 (n32422, n_23864, n_23865);
  not g53281 (n_23866, n32422);
  and g53282 (n32423, pi0644, n_23866);
  and g53283 (n32424, n_11819, n32255);
  not g53284 (n_23867, n32424);
  and g53285 (n32425, n_12395, n_23867);
  not g53286 (n_23868, n32423);
  and g53287 (n32426, n_23868, n32425);
  not g53288 (n_23869, n32426);
  and g53289 (n32427, pi1160, n_23869);
  not g53290 (n_23870, n32419);
  and g53291 (n32428, n_23870, n32427);
  and g53292 (n32429, n_11819, n_23866);
  and g53293 (n32430, pi0644, n32255);
  not g53294 (n_23871, n32430);
  and g53295 (n32431, pi0715, n_23871);
  not g53296 (n_23872, n32429);
  and g53297 (n32432, n_23872, n32431);
  and g53298 (n32433, pi0644, n32415);
  and g53299 (n32434, n_11819, n32409);
  not g53300 (n_23873, n32433);
  and g53301 (n32435, n_12395, n_23873);
  not g53302 (n_23874, n32434);
  and g53303 (n32436, n_23874, n32435);
  not g53304 (n_23875, n32432);
  and g53305 (n32437, n_12405, n_23875);
  not g53306 (n_23876, n32436);
  and g53307 (n32438, n_23876, n32437);
  not g53308 (n_23877, n32428);
  not g53309 (n_23878, n32438);
  and g53310 (n32439, n_23877, n_23878);
  not g53311 (n_23879, n32439);
  and g53312 (n32440, pi0790, n_23879);
  not g53313 (n_23880, n32410);
  and g53314 (n32441, pi0832, n_23880);
  not g53315 (n_23881, n32440);
  and g53316 (n32442, n_23881, n32441);
  and g53317 (n32443, n_5790, po1038);
  and g53318 (n32444, n_5790, n_11751);
  not g53319 (n_23882, n32444);
  and g53320 (n32445, n16635, n_23882);
  and g53321 (n32446, pi0690, n2571);
  not g53322 (n_23883, n32446);
  and g53323 (n32447, n32444, n_23883);
  and g53324 (n32448, n_5790, n_11418);
  not g53325 (n_23884, n32448);
  and g53326 (n32449, n16647, n_23884);
  and g53327 (n32450, pi0193, n_12608);
  not g53328 (n_23885, n32450);
  and g53329 (n32451, n_161, n_23885);
  not g53330 (n_23886, n32451);
  and g53331 (n32452, n2571, n_23886);
  and g53332 (n32453, n_5790, n18072);
  not g53333 (n_23887, n32452);
  not g53334 (n_23888, n32453);
  and g53335 (n32454, n_23887, n_23888);
  not g53336 (n_23889, n32449);
  and g53337 (n32455, pi0690, n_23889);
  not g53338 (n_23890, n32454);
  and g53339 (n32456, n_23890, n32455);
  not g53340 (n_23891, n32447);
  not g53341 (n_23892, n32456);
  and g53342 (n32457, n_23891, n_23892);
  and g53343 (n32458, n_11749, n32457);
  and g53344 (n32459, n_11753, n32444);
  not g53345 (n_23893, n32457);
  and g53346 (n32460, pi0625, n_23893);
  not g53347 (n_23894, n32459);
  and g53348 (n32461, pi1153, n_23894);
  not g53349 (n_23895, n32460);
  and g53350 (n32462, n_23895, n32461);
  and g53351 (n32463, pi0625, n32444);
  and g53352 (n32464, n_11753, n_23893);
  not g53353 (n_23896, n32463);
  and g53354 (n32465, n_11757, n_23896);
  not g53355 (n_23897, n32464);
  and g53356 (n32466, n_23897, n32465);
  not g53357 (n_23898, n32462);
  not g53358 (n_23899, n32466);
  and g53359 (n32467, n_23898, n_23899);
  not g53360 (n_23900, n32467);
  and g53361 (n32468, pi0778, n_23900);
  not g53362 (n_23901, n32458);
  not g53363 (n_23902, n32468);
  and g53364 (n32469, n_23901, n_23902);
  not g53365 (n_23903, n32469);
  and g53366 (n32470, n_11773, n_23903);
  and g53367 (n32471, n17075, n_23882);
  not g53368 (n_23904, n32470);
  not g53369 (n_23905, n32471);
  and g53370 (n32472, n_23904, n_23905);
  and g53371 (n32473, n_11777, n32472);
  and g53372 (n32474, n16639, n32444);
  not g53373 (n_23906, n32473);
  not g53374 (n_23907, n32474);
  and g53375 (n32475, n_23906, n_23907);
  and g53376 (n32476, n_11780, n32475);
  not g53377 (n_23908, n32445);
  not g53378 (n_23909, n32476);
  and g53379 (n32477, n_23908, n_23909);
  and g53380 (n32478, n_11783, n32477);
  and g53381 (n32479, n16631, n32444);
  not g53382 (n_23910, n32478);
  not g53383 (n_23911, n32479);
  and g53384 (n32480, n_23910, n_23911);
  and g53385 (n32481, n_11787, n32480);
  not g53386 (n_23912, n32480);
  and g53387 (n32482, pi0628, n_23912);
  and g53388 (n32483, n_11789, n32444);
  not g53389 (n_23913, n32483);
  and g53390 (n32484, pi1156, n_23913);
  not g53391 (n_23914, n32482);
  and g53392 (n32485, n_23914, n32484);
  and g53393 (n32486, pi0628, n32444);
  and g53394 (n32487, n_11789, n_23912);
  not g53395 (n_23915, n32486);
  and g53396 (n32488, n_11794, n_23915);
  not g53397 (n_23916, n32487);
  and g53398 (n32489, n_23916, n32488);
  not g53399 (n_23917, n32485);
  not g53400 (n_23918, n32489);
  and g53401 (n32490, n_23917, n_23918);
  not g53402 (n_23919, n32490);
  and g53403 (n32491, pi0792, n_23919);
  not g53404 (n_23920, n32481);
  not g53405 (n_23921, n32491);
  and g53406 (n32492, n_23920, n_23921);
  not g53407 (n_23922, n32492);
  and g53408 (n32493, n_11806, n_23922);
  and g53409 (n32494, pi0647, n_23882);
  not g53410 (n_23923, n32493);
  not g53411 (n_23924, n32494);
  and g53412 (n32495, n_23923, n_23924);
  and g53413 (n32496, n_11810, n32495);
  and g53414 (n32497, pi0647, n_23922);
  and g53415 (n32498, n_11806, n_23882);
  not g53416 (n_23925, n32497);
  not g53417 (n_23926, n32498);
  and g53418 (n32499, n_23925, n_23926);
  and g53419 (n32500, pi1157, n32499);
  not g53420 (n_23927, n32496);
  not g53421 (n_23928, n32500);
  and g53422 (n32501, n_23927, n_23928);
  not g53423 (n_23929, n32501);
  and g53424 (n32502, pi0787, n_23929);
  and g53425 (n32503, n_11803, n32492);
  not g53426 (n_23930, n32502);
  not g53427 (n_23931, n32503);
  and g53428 (n32504, n_23930, n_23931);
  not g53429 (n_23932, n32504);
  and g53430 (n32505, n_11819, n_23932);
  not g53431 (n_23933, n32505);
  and g53432 (n32506, pi0715, n_23933);
  and g53433 (n32507, pi0193, n_11417);
  and g53434 (n32508, pi0739, n17280);
  not g53435 (n_23934, n32508);
  and g53436 (n32509, n_23884, n_23934);
  not g53437 (n_23935, n32509);
  and g53438 (n32510, pi0038, n_23935);
  and g53439 (n32511, n_5790, n17221);
  and g53440 (n32512, pi0193, n_14476);
  not g53441 (n_23936, n32512);
  and g53442 (n32513, pi0739, n_23936);
  not g53443 (n_23937, n32511);
  and g53444 (n32514, n_23937, n32513);
  and g53445 (n32515, n_5790, n_16204);
  and g53446 (n32516, n_11739, n32515);
  not g53447 (n_23938, n32514);
  not g53448 (n_23939, n32516);
  and g53449 (n32517, n_23938, n_23939);
  not g53450 (n_23940, n32517);
  and g53451 (n32518, n_161, n_23940);
  not g53452 (n_23941, n32510);
  not g53453 (n_23942, n32518);
  and g53454 (n32519, n_23941, n_23942);
  and g53455 (n32520, n2571, n32519);
  not g53456 (n_23943, n32507);
  not g53457 (n_23944, n32520);
  and g53458 (n32521, n_23943, n_23944);
  not g53459 (n_23945, n32521);
  and g53460 (n32522, n_11960, n_23945);
  and g53461 (n32523, n17117, n_23882);
  not g53462 (n_23946, n32522);
  not g53463 (n_23947, n32523);
  and g53464 (n32524, n_23946, n_23947);
  not g53465 (n_23948, n32524);
  and g53466 (n32525, n_11964, n_23948);
  and g53467 (n32526, n_11967, n_23882);
  and g53468 (n32527, pi0609, n32522);
  not g53469 (n_23949, n32526);
  not g53470 (n_23950, n32527);
  and g53471 (n32528, n_23949, n_23950);
  not g53472 (n_23951, n32528);
  and g53473 (n32529, pi1155, n_23951);
  and g53474 (n32530, n_11972, n_23882);
  and g53475 (n32531, n_11971, n32522);
  not g53476 (n_23952, n32530);
  not g53477 (n_23953, n32531);
  and g53478 (n32532, n_23952, n_23953);
  not g53479 (n_23954, n32532);
  and g53480 (n32533, n_11768, n_23954);
  not g53481 (n_23955, n32529);
  not g53482 (n_23956, n32533);
  and g53483 (n32534, n_23955, n_23956);
  not g53484 (n_23957, n32534);
  and g53485 (n32535, pi0785, n_23957);
  not g53486 (n_23958, n32525);
  not g53487 (n_23959, n32535);
  and g53488 (n32536, n_23958, n_23959);
  not g53489 (n_23960, n32536);
  and g53490 (n32537, n_11981, n_23960);
  and g53491 (n32538, n_11984, n32444);
  and g53492 (n32539, pi0618, n32536);
  not g53493 (n_23961, n32538);
  and g53494 (n32540, pi1154, n_23961);
  not g53495 (n_23962, n32539);
  and g53496 (n32541, n_23962, n32540);
  and g53497 (n32542, n_11984, n32536);
  and g53498 (n32543, pi0618, n32444);
  not g53499 (n_23963, n32543);
  and g53500 (n32544, n_11413, n_23963);
  not g53501 (n_23964, n32542);
  and g53502 (n32545, n_23964, n32544);
  not g53503 (n_23965, n32541);
  not g53504 (n_23966, n32545);
  and g53505 (n32546, n_23965, n_23966);
  not g53506 (n_23967, n32546);
  and g53507 (n32547, pi0781, n_23967);
  not g53508 (n_23968, n32537);
  not g53509 (n_23969, n32547);
  and g53510 (n32548, n_23968, n_23969);
  not g53511 (n_23970, n32548);
  and g53512 (n32549, n_12315, n_23970);
  and g53513 (n32550, n_11821, n32444);
  and g53514 (n32551, pi0619, n32548);
  not g53515 (n_23971, n32550);
  and g53516 (n32552, pi1159, n_23971);
  not g53517 (n_23972, n32551);
  and g53518 (n32553, n_23972, n32552);
  and g53519 (n32554, n_11821, n32548);
  and g53520 (n32555, pi0619, n32444);
  not g53521 (n_23973, n32555);
  and g53522 (n32556, n_11405, n_23973);
  not g53523 (n_23974, n32554);
  and g53524 (n32557, n_23974, n32556);
  not g53525 (n_23975, n32553);
  not g53526 (n_23976, n32557);
  and g53527 (n32558, n_23975, n_23976);
  not g53528 (n_23977, n32558);
  and g53529 (n32559, pi0789, n_23977);
  not g53530 (n_23978, n32549);
  not g53531 (n_23979, n32559);
  and g53532 (n32560, n_23978, n_23979);
  and g53533 (n32561, n_12524, n32560);
  and g53534 (n32562, n17969, n32444);
  not g53535 (n_23980, n32561);
  not g53536 (n_23981, n32562);
  and g53537 (n32563, n_23980, n_23981);
  not g53538 (n_23982, n32563);
  and g53539 (n32564, n_12368, n_23982);
  and g53540 (n32565, n17779, n32444);
  not g53541 (n_23983, n32564);
  not g53542 (n_23984, n32565);
  and g53543 (n32566, n_23983, n_23984);
  not g53544 (n_23985, n32566);
  and g53545 (n32567, n_12392, n_23985);
  and g53546 (n32568, n17804, n32444);
  not g53547 (n_23986, n32567);
  not g53548 (n_23987, n32568);
  and g53549 (n32569, n_23986, n_23987);
  not g53550 (n_23988, n32569);
  and g53551 (n32570, pi0644, n_23988);
  and g53552 (n32571, n_11819, n32444);
  not g53553 (n_23989, n32571);
  and g53554 (n32572, n_12395, n_23989);
  not g53555 (n_23990, n32570);
  and g53556 (n32573, n_23990, n32572);
  not g53557 (n_23991, n32573);
  and g53558 (n32574, pi1160, n_23991);
  not g53559 (n_23992, n32506);
  and g53560 (n32575, n_23992, n32574);
  and g53561 (n32576, pi0644, n_23932);
  not g53562 (n_23993, n32576);
  and g53563 (n32577, n_12395, n_23993);
  and g53564 (n32578, n_11819, n_23988);
  and g53565 (n32579, pi0644, n32444);
  not g53566 (n_23994, n32579);
  and g53567 (n32580, pi0715, n_23994);
  not g53568 (n_23995, n32578);
  and g53569 (n32581, n_23995, n32580);
  not g53570 (n_23996, n32581);
  and g53571 (n32582, n_12405, n_23996);
  not g53572 (n_23997, n32577);
  and g53573 (n32583, n_23997, n32582);
  not g53574 (n_23998, n32575);
  not g53575 (n_23999, n32583);
  and g53576 (n32584, n_23998, n_23999);
  not g53577 (n_24000, n32584);
  and g53578 (n32585, pi0790, n_24000);
  and g53579 (n32586, n_12354, n32485);
  and g53580 (n32587, n_14557, n32563);
  and g53581 (n32588, pi0629, n32489);
  not g53582 (n_24001, n32586);
  not g53583 (n_24002, n32588);
  and g53584 (n32589, n_24001, n_24002);
  not g53585 (n_24003, n32587);
  and g53586 (n32590, n_24003, n32589);
  not g53587 (n_24004, n32590);
  and g53588 (n32591, pi0792, n_24004);
  and g53589 (n32592, pi0609, n32469);
  not g53590 (n_24005, n32519);
  and g53591 (n32593, n_16236, n_24005);
  and g53592 (n32594, n_5790, n17629);
  and g53593 (n32595, pi0193, n17631);
  not g53594 (n_24006, n32595);
  and g53595 (n32596, pi0739, n_24006);
  not g53596 (n_24007, n32594);
  and g53597 (n32597, n_24007, n32596);
  and g53598 (n32598, pi0193, n_12240);
  and g53599 (n32599, n_5790, n_12230);
  not g53600 (n_24008, n32598);
  and g53601 (n32600, n_16204, n_24008);
  not g53602 (n_24009, n32599);
  and g53603 (n32601, n_24009, n32600);
  not g53604 (n_24010, n32597);
  not g53605 (n_24011, n32601);
  and g53606 (n32602, n_24010, n_24011);
  not g53607 (n_24012, n32602);
  and g53608 (n32603, n_162, n_24012);
  and g53609 (n32604, pi0193, n17605);
  and g53610 (n32605, n_5790, n_12180);
  not g53611 (n_24013, n32605);
  and g53612 (n32606, pi0739, n_24013);
  not g53613 (n_24014, n32604);
  and g53614 (n32607, n_24014, n32606);
  and g53615 (n32608, n_5790, n17404);
  and g53616 (n32609, pi0193, n17485);
  not g53617 (n_24015, n32609);
  and g53618 (n32610, n_16204, n_24015);
  not g53619 (n_24016, n32608);
  and g53620 (n32611, n_24016, n32610);
  not g53621 (n_24017, n32607);
  and g53622 (n32612, pi0039, n_24017);
  not g53623 (n_24018, n32611);
  and g53624 (n32613, n_24018, n32612);
  not g53625 (n_24019, n32603);
  and g53626 (n32614, n_161, n_24019);
  not g53627 (n_24020, n32613);
  and g53628 (n32615, n_24020, n32614);
  and g53629 (n32616, n_16204, n24055);
  not g53630 (n_24021, n32616);
  and g53631 (n32617, n_12250, n_24021);
  not g53632 (n_24022, n32617);
  and g53633 (n32618, n_162, n_24022);
  not g53634 (n_24023, n32618);
  and g53635 (n32619, n_5790, n_24023);
  and g53636 (n32620, n_12120, n_23746);
  not g53637 (n_24024, n32620);
  and g53638 (n32621, pi0193, n_24024);
  and g53639 (n32622, n6284, n32621);
  not g53640 (n_24025, n32622);
  and g53641 (n32623, pi0038, n_24025);
  not g53642 (n_24026, n32619);
  and g53643 (n32624, n_24026, n32623);
  not g53644 (n_24027, n32624);
  and g53645 (n32625, pi0690, n_24027);
  not g53646 (n_24028, n32615);
  and g53647 (n32626, n_24028, n32625);
  not g53648 (n_24029, n32626);
  and g53649 (n32627, n2571, n_24029);
  not g53650 (n_24030, n32593);
  and g53651 (n32628, n_24030, n32627);
  not g53652 (n_24031, n32628);
  and g53653 (n32629, n_23943, n_24031);
  and g53654 (n32630, n_11753, n32629);
  and g53655 (n32631, pi0625, n32521);
  not g53656 (n_24032, n32631);
  and g53657 (n32632, n_11757, n_24032);
  not g53658 (n_24033, n32630);
  and g53659 (n32633, n_24033, n32632);
  and g53660 (n32634, n_11823, n_23898);
  not g53661 (n_24034, n32633);
  and g53662 (n32635, n_24034, n32634);
  and g53663 (n32636, n_11753, n32521);
  and g53664 (n32637, pi0625, n32629);
  not g53665 (n_24035, n32636);
  and g53666 (n32638, pi1153, n_24035);
  not g53667 (n_24036, n32637);
  and g53668 (n32639, n_24036, n32638);
  and g53669 (n32640, pi0608, n_23899);
  not g53670 (n_24037, n32639);
  and g53671 (n32641, n_24037, n32640);
  not g53672 (n_24038, n32635);
  not g53673 (n_24039, n32641);
  and g53674 (n32642, n_24038, n_24039);
  not g53675 (n_24040, n32642);
  and g53676 (n32643, pi0778, n_24040);
  and g53677 (n32644, n_11749, n32629);
  not g53678 (n_24041, n32643);
  not g53679 (n_24042, n32644);
  and g53680 (n32645, n_24041, n_24042);
  not g53681 (n_24043, n32645);
  and g53682 (n32646, n_11971, n_24043);
  not g53683 (n_24044, n32592);
  and g53684 (n32647, n_11768, n_24044);
  not g53685 (n_24045, n32646);
  and g53686 (n32648, n_24045, n32647);
  and g53687 (n32649, n_11767, n_23955);
  not g53688 (n_24046, n32648);
  and g53689 (n32650, n_24046, n32649);
  and g53690 (n32651, n_11971, n32469);
  and g53691 (n32652, pi0609, n_24043);
  not g53692 (n_24047, n32651);
  and g53693 (n32653, pi1155, n_24047);
  not g53694 (n_24048, n32652);
  and g53695 (n32654, n_24048, n32653);
  and g53696 (n32655, pi0660, n_23956);
  not g53697 (n_24049, n32654);
  and g53698 (n32656, n_24049, n32655);
  not g53699 (n_24050, n32650);
  not g53700 (n_24051, n32656);
  and g53701 (n32657, n_24050, n_24051);
  not g53702 (n_24052, n32657);
  and g53703 (n32658, pi0785, n_24052);
  and g53704 (n32659, n_11964, n_24043);
  not g53705 (n_24053, n32658);
  not g53706 (n_24054, n32659);
  and g53707 (n32660, n_24053, n_24054);
  not g53708 (n_24055, n32660);
  and g53709 (n32661, n_11984, n_24055);
  and g53710 (n32662, pi0618, n32472);
  not g53711 (n_24056, n32662);
  and g53712 (n32663, n_11413, n_24056);
  not g53713 (n_24057, n32661);
  and g53714 (n32664, n_24057, n32663);
  and g53715 (n32665, n_11412, n_23965);
  not g53716 (n_24058, n32664);
  and g53717 (n32666, n_24058, n32665);
  and g53718 (n32667, n_11984, n32472);
  and g53719 (n32668, pi0618, n_24055);
  not g53720 (n_24059, n32667);
  and g53721 (n32669, pi1154, n_24059);
  not g53722 (n_24060, n32668);
  and g53723 (n32670, n_24060, n32669);
  and g53724 (n32671, pi0627, n_23966);
  not g53725 (n_24061, n32670);
  and g53726 (n32672, n_24061, n32671);
  not g53727 (n_24062, n32666);
  not g53728 (n_24063, n32672);
  and g53729 (n32673, n_24062, n_24063);
  not g53730 (n_24064, n32673);
  and g53731 (n32674, pi0781, n_24064);
  and g53732 (n32675, n_11981, n_24055);
  not g53733 (n_24065, n32674);
  not g53734 (n_24066, n32675);
  and g53735 (n32676, n_24065, n_24066);
  and g53736 (n32677, n_12315, n32676);
  not g53737 (n_24067, n32475);
  and g53738 (n32678, pi0619, n_24067);
  not g53739 (n_24068, n32676);
  and g53740 (n32679, n_11821, n_24068);
  not g53741 (n_24069, n32678);
  and g53742 (n32680, n_11405, n_24069);
  not g53743 (n_24070, n32679);
  and g53744 (n32681, n_24070, n32680);
  and g53745 (n32682, n_11403, n_23975);
  not g53746 (n_24071, n32681);
  and g53747 (n32683, n_24071, n32682);
  and g53748 (n32684, n_11821, n_24067);
  and g53749 (n32685, pi0619, n_24068);
  not g53750 (n_24072, n32684);
  and g53751 (n32686, pi1159, n_24072);
  not g53752 (n_24073, n32685);
  and g53753 (n32687, n_24073, n32686);
  and g53754 (n32688, pi0648, n_23976);
  not g53755 (n_24074, n32687);
  and g53756 (n32689, n_24074, n32688);
  not g53757 (n_24075, n32683);
  and g53758 (n32690, pi0789, n_24075);
  not g53759 (n_24076, n32689);
  and g53760 (n32691, n_24076, n32690);
  not g53761 (n_24077, n32677);
  and g53762 (n32692, n17970, n_24077);
  not g53763 (n_24078, n32691);
  and g53764 (n32693, n_24078, n32692);
  and g53765 (n32694, n17871, n32477);
  not g53766 (n_24079, n32560);
  and g53767 (n32695, n_12320, n_24079);
  and g53768 (n32696, pi0626, n_23882);
  not g53769 (n_24080, n32696);
  and g53770 (n32697, n16629, n_24080);
  not g53771 (n_24081, n32695);
  and g53772 (n32698, n_24081, n32697);
  and g53773 (n32699, pi0626, n_24079);
  and g53774 (n32700, n_12320, n_23882);
  not g53775 (n_24082, n32700);
  and g53776 (n32701, n16628, n_24082);
  not g53777 (n_24083, n32699);
  and g53778 (n32702, n_24083, n32701);
  not g53779 (n_24084, n32694);
  not g53780 (n_24085, n32698);
  and g53781 (n32703, n_24084, n_24085);
  not g53782 (n_24086, n32702);
  and g53783 (n32704, n_24086, n32703);
  not g53784 (n_24087, n32704);
  and g53785 (n32705, pi0788, n_24087);
  not g53786 (n_24088, n32705);
  and g53787 (n32706, n_14638, n_24088);
  not g53788 (n_24089, n32693);
  and g53789 (n32707, n_24089, n32706);
  not g53790 (n_24090, n32591);
  not g53791 (n_24091, n32707);
  and g53792 (n32708, n_24090, n_24091);
  not g53793 (n_24092, n32708);
  and g53794 (n32709, n_14387, n_24092);
  not g53795 (n_24093, n32495);
  and g53796 (n32710, n17802, n_24093);
  and g53797 (n32711, n_14548, n32566);
  not g53798 (n_24094, n32499);
  and g53799 (n32712, n17801, n_24094);
  not g53800 (n_24095, n32710);
  not g53801 (n_24096, n32712);
  and g53802 (n32713, n_24095, n_24096);
  not g53803 (n_24097, n32711);
  and g53804 (n32714, n_24097, n32713);
  not g53805 (n_24098, n32714);
  and g53806 (n32715, pi0787, n_24098);
  and g53807 (n32716, n_11819, n32582);
  and g53808 (n32717, pi0644, n32574);
  not g53809 (n_24099, n32716);
  and g53810 (n32718, pi0790, n_24099);
  not g53811 (n_24100, n32717);
  and g53812 (n32719, n_24100, n32718);
  not g53813 (n_24101, n32709);
  not g53814 (n_24102, n32715);
  and g53815 (n32720, n_24101, n_24102);
  not g53816 (n_24103, n32719);
  and g53817 (n32721, n_24103, n32720);
  not g53818 (n_24104, n32585);
  not g53819 (n_24105, n32721);
  and g53820 (n32722, n_24104, n_24105);
  not g53821 (n_24106, n32722);
  and g53822 (n32723, n_4226, n_24106);
  not g53823 (n_24107, n32443);
  and g53824 (n32724, n_12415, n_24107);
  not g53825 (n_24108, n32723);
  and g53826 (n32725, n_24108, n32724);
  not g53827 (n_24109, n32442);
  not g53828 (n_24110, n32725);
  and g53829 (po0350, n_24109, n_24110);
  and g53830 (n32727, n_11115, n_11751);
  not g53831 (n_24111, n32727);
  and g53832 (n32728, n16635, n_24111);
  and g53833 (n32729, pi0194, n_17520);
  and g53834 (n32730, n_11115, n24388);
  not g53835 (n_24112, n32730);
  and g53836 (n32731, pi0730, n_24112);
  and g53837 (n32732, n_11115, n_11743);
  and g53838 (n32733, n_16117, n32732);
  not g53839 (n_24113, n32733);
  and g53840 (n32734, n2571, n_24113);
  not g53841 (n_24114, n32731);
  and g53842 (n32735, n_24114, n32734);
  not g53843 (n_24115, n32729);
  not g53844 (n_24116, n32735);
  and g53845 (n32736, n_24115, n_24116);
  not g53846 (n_24117, n32736);
  and g53847 (n32737, n_11749, n_24117);
  and g53848 (n32738, n_11753, n32727);
  and g53849 (n32739, pi0625, n32736);
  not g53850 (n_24118, n32738);
  and g53851 (n32740, pi1153, n_24118);
  not g53852 (n_24119, n32739);
  and g53853 (n32741, n_24119, n32740);
  and g53854 (n32742, n_11753, n32736);
  and g53855 (n32743, pi0625, n32727);
  not g53856 (n_24120, n32743);
  and g53857 (n32744, n_11757, n_24120);
  not g53858 (n_24121, n32742);
  and g53859 (n32745, n_24121, n32744);
  not g53860 (n_24122, n32741);
  not g53861 (n_24123, n32745);
  and g53862 (n32746, n_24122, n_24123);
  not g53863 (n_24124, n32746);
  and g53864 (n32747, pi0778, n_24124);
  not g53865 (n_24125, n32737);
  not g53866 (n_24126, n32747);
  and g53867 (n32748, n_24125, n_24126);
  not g53868 (n_24127, n32748);
  and g53869 (n32749, n_11773, n_24127);
  and g53870 (n32750, n17075, n_24111);
  not g53871 (n_24128, n32749);
  not g53872 (n_24129, n32750);
  and g53873 (n32751, n_24128, n_24129);
  and g53874 (n32752, n_11777, n32751);
  and g53875 (n32753, n16639, n32727);
  not g53876 (n_24130, n32752);
  not g53877 (n_24131, n32753);
  and g53878 (n32754, n_24130, n_24131);
  and g53879 (n32755, n_11780, n32754);
  not g53880 (n_24132, n32728);
  not g53881 (n_24133, n32755);
  and g53882 (n32756, n_24132, n_24133);
  and g53883 (n32757, n_11783, n32756);
  and g53884 (n32758, n16631, n32727);
  not g53885 (n_24134, n32757);
  not g53886 (n_24135, n32758);
  and g53887 (n32759, n_24134, n_24135);
  and g53888 (n32760, n_11787, n32759);
  and g53889 (n32761, n_11789, n32727);
  not g53890 (n_24136, n32759);
  and g53891 (n32762, pi0628, n_24136);
  not g53892 (n_24137, n32761);
  and g53893 (n32763, pi1156, n_24137);
  not g53894 (n_24138, n32762);
  and g53895 (n32764, n_24138, n32763);
  and g53896 (n32765, pi0628, n32727);
  and g53897 (n32766, n_11789, n_24136);
  not g53898 (n_24139, n32765);
  and g53899 (n32767, n_11794, n_24139);
  not g53900 (n_24140, n32766);
  and g53901 (n32768, n_24140, n32767);
  not g53902 (n_24141, n32764);
  not g53903 (n_24142, n32768);
  and g53904 (n32769, n_24141, n_24142);
  not g53905 (n_24143, n32769);
  and g53906 (n32770, pi0792, n_24143);
  not g53907 (n_24144, n32760);
  not g53908 (n_24145, n32770);
  and g53909 (n32771, n_24144, n_24145);
  not g53910 (n_24146, n32771);
  and g53911 (n32772, n_11803, n_24146);
  and g53912 (n32773, n_11806, n32727);
  and g53913 (n32774, pi0647, n32771);
  not g53914 (n_24147, n32773);
  and g53915 (n32775, pi1157, n_24147);
  not g53916 (n_24148, n32774);
  and g53917 (n32776, n_24148, n32775);
  and g53918 (n32777, n_11806, n32771);
  and g53919 (n32778, pi0647, n32727);
  not g53920 (n_24149, n32778);
  and g53921 (n32779, n_11810, n_24149);
  not g53922 (n_24150, n32777);
  and g53923 (n32780, n_24150, n32779);
  not g53924 (n_24151, n32776);
  not g53925 (n_24152, n32780);
  and g53926 (n32781, n_24151, n_24152);
  not g53927 (n_24153, n32781);
  and g53928 (n32782, pi0787, n_24153);
  not g53929 (n_24154, n32772);
  not g53930 (n_24155, n32782);
  and g53931 (n32783, n_24154, n_24155);
  and g53932 (n32784, n_11819, n32783);
  and g53933 (n32785, n_11984, n32727);
  and g53934 (n32786, pi0194, n_11417);
  and g53935 (n32787, n_11115, n19439);
  and g53936 (n32788, pi0194, n24447);
  not g53937 (n_24156, n32787);
  not g53938 (n_24157, n32788);
  and g53939 (n32789, n_24156, n_24157);
  not g53940 (n_24158, n32789);
  and g53941 (n32790, pi0748, n_24158);
  not g53942 (n_24159, n32732);
  and g53943 (n32791, n_16089, n_24159);
  not g53944 (n_24160, n32790);
  not g53945 (n_24161, n32791);
  and g53946 (n32792, n_24160, n_24161);
  not g53947 (n_24162, n32792);
  and g53948 (n32793, n2571, n_24162);
  not g53949 (n_24163, n32786);
  not g53950 (n_24164, n32793);
  and g53951 (n32794, n_24163, n_24164);
  not g53952 (n_24165, n32794);
  and g53953 (n32795, n_11960, n_24165);
  and g53954 (n32796, n17117, n_24111);
  not g53955 (n_24166, n32795);
  not g53956 (n_24167, n32796);
  and g53957 (n32797, n_24166, n_24167);
  not g53958 (n_24168, n32797);
  and g53959 (n32798, n_11964, n_24168);
  and g53960 (n32799, n_11967, n_24111);
  and g53961 (n32800, pi0609, n32795);
  not g53962 (n_24169, n32799);
  not g53963 (n_24170, n32800);
  and g53964 (n32801, n_24169, n_24170);
  not g53965 (n_24171, n32801);
  and g53966 (n32802, pi1155, n_24171);
  and g53967 (n32803, n_11972, n_24111);
  and g53968 (n32804, n_11971, n32795);
  not g53969 (n_24172, n32803);
  not g53970 (n_24173, n32804);
  and g53971 (n32805, n_24172, n_24173);
  not g53972 (n_24174, n32805);
  and g53973 (n32806, n_11768, n_24174);
  not g53974 (n_24175, n32802);
  not g53975 (n_24176, n32806);
  and g53976 (n32807, n_24175, n_24176);
  not g53977 (n_24177, n32807);
  and g53978 (n32808, pi0785, n_24177);
  not g53979 (n_24178, n32798);
  not g53980 (n_24179, n32808);
  and g53981 (n32809, n_24178, n_24179);
  and g53982 (n32810, pi0618, n32809);
  not g53983 (n_24180, n32785);
  and g53984 (n32811, pi1154, n_24180);
  not g53985 (n_24181, n32810);
  and g53986 (n32812, n_24181, n32811);
  and g53987 (n32813, n_16117, n32792);
  and g53988 (n32814, pi0194, n19496);
  and g53989 (n32815, n_11115, n_13718);
  not g53990 (n_24182, n32815);
  and g53991 (n32816, pi0748, n_24182);
  not g53992 (n_24183, n32814);
  and g53993 (n32817, n_24183, n32816);
  and g53994 (n32818, pi0194, n_17658);
  and g53995 (n32819, n_11115, n19477);
  not g53996 (n_24184, n32818);
  and g53997 (n32820, n_16089, n_24184);
  not g53998 (n_24185, n32819);
  and g53999 (n32821, n_24185, n32820);
  not g54000 (n_24186, n32817);
  and g54001 (n32822, pi0730, n_24186);
  not g54002 (n_24187, n32821);
  and g54003 (n32823, n_24187, n32822);
  not g54004 (n_24188, n32813);
  and g54005 (n32824, n2571, n_24188);
  not g54006 (n_24189, n32823);
  and g54007 (n32825, n_24189, n32824);
  not g54008 (n_24190, n32825);
  and g54009 (n32826, n_24163, n_24190);
  and g54010 (n32827, n_11753, n32826);
  and g54011 (n32828, pi0625, n32794);
  not g54012 (n_24191, n32828);
  and g54013 (n32829, n_11757, n_24191);
  not g54014 (n_24192, n32827);
  and g54015 (n32830, n_24192, n32829);
  and g54016 (n32831, n_11823, n_24122);
  not g54017 (n_24193, n32830);
  and g54018 (n32832, n_24193, n32831);
  and g54019 (n32833, n_11753, n32794);
  and g54020 (n32834, pi0625, n32826);
  not g54021 (n_24194, n32833);
  and g54022 (n32835, pi1153, n_24194);
  not g54023 (n_24195, n32834);
  and g54024 (n32836, n_24195, n32835);
  and g54025 (n32837, pi0608, n_24123);
  not g54026 (n_24196, n32836);
  and g54027 (n32838, n_24196, n32837);
  not g54028 (n_24197, n32832);
  not g54029 (n_24198, n32838);
  and g54030 (n32839, n_24197, n_24198);
  not g54031 (n_24199, n32839);
  and g54032 (n32840, pi0778, n_24199);
  and g54033 (n32841, n_11749, n32826);
  not g54034 (n_24200, n32840);
  not g54035 (n_24201, n32841);
  and g54036 (n32842, n_24200, n_24201);
  not g54037 (n_24202, n32842);
  and g54038 (n32843, n_11971, n_24202);
  and g54039 (n32844, pi0609, n32748);
  not g54040 (n_24203, n32844);
  and g54041 (n32845, n_11768, n_24203);
  not g54042 (n_24204, n32843);
  and g54043 (n32846, n_24204, n32845);
  and g54044 (n32847, n_11767, n_24175);
  not g54045 (n_24205, n32846);
  and g54046 (n32848, n_24205, n32847);
  and g54047 (n32849, n_11971, n32748);
  and g54048 (n32850, pi0609, n_24202);
  not g54049 (n_24206, n32849);
  and g54050 (n32851, pi1155, n_24206);
  not g54051 (n_24207, n32850);
  and g54052 (n32852, n_24207, n32851);
  and g54053 (n32853, pi0660, n_24176);
  not g54054 (n_24208, n32852);
  and g54055 (n32854, n_24208, n32853);
  not g54056 (n_24209, n32848);
  not g54057 (n_24210, n32854);
  and g54058 (n32855, n_24209, n_24210);
  not g54059 (n_24211, n32855);
  and g54060 (n32856, pi0785, n_24211);
  and g54061 (n32857, n_11964, n_24202);
  not g54062 (n_24212, n32856);
  not g54063 (n_24213, n32857);
  and g54064 (n32858, n_24212, n_24213);
  not g54065 (n_24214, n32858);
  and g54066 (n32859, n_11984, n_24214);
  and g54067 (n32860, pi0618, n32751);
  not g54068 (n_24215, n32860);
  and g54069 (n32861, n_11413, n_24215);
  not g54070 (n_24216, n32859);
  and g54071 (n32862, n_24216, n32861);
  not g54072 (n_24217, n32812);
  and g54073 (n32863, n_11412, n_24217);
  not g54074 (n_24218, n32862);
  and g54075 (n32864, n_24218, n32863);
  and g54076 (n32865, n_11984, n32809);
  and g54077 (n32866, pi0618, n32727);
  not g54078 (n_24219, n32866);
  and g54079 (n32867, n_11413, n_24219);
  not g54080 (n_24220, n32865);
  and g54081 (n32868, n_24220, n32867);
  and g54082 (n32869, n_11984, n32751);
  and g54083 (n32870, pi0618, n_24214);
  not g54084 (n_24221, n32869);
  and g54085 (n32871, pi1154, n_24221);
  not g54086 (n_24222, n32870);
  and g54087 (n32872, n_24222, n32871);
  not g54088 (n_24223, n32868);
  and g54089 (n32873, pi0627, n_24223);
  not g54090 (n_24224, n32872);
  and g54091 (n32874, n_24224, n32873);
  not g54092 (n_24225, n32864);
  not g54093 (n_24226, n32874);
  and g54094 (n32875, n_24225, n_24226);
  not g54095 (n_24227, n32875);
  and g54096 (n32876, pi0781, n_24227);
  and g54097 (n32877, n_11981, n_24214);
  not g54098 (n_24228, n32876);
  not g54099 (n_24229, n32877);
  and g54100 (n32878, n_24228, n_24229);
  not g54101 (n_24230, n32878);
  and g54102 (n32879, n_11821, n_24230);
  not g54103 (n_24231, n32754);
  and g54104 (n32880, pi0619, n_24231);
  not g54105 (n_24232, n32880);
  and g54106 (n32881, n_11405, n_24232);
  not g54107 (n_24233, n32879);
  and g54108 (n32882, n_24233, n32881);
  and g54109 (n32883, n_11821, n32727);
  not g54110 (n_24234, n32809);
  and g54111 (n32884, n_11981, n_24234);
  and g54112 (n32885, n_24217, n_24223);
  not g54113 (n_24235, n32885);
  and g54114 (n32886, pi0781, n_24235);
  not g54115 (n_24236, n32884);
  not g54116 (n_24237, n32886);
  and g54117 (n32887, n_24236, n_24237);
  and g54118 (n32888, pi0619, n32887);
  not g54119 (n_24238, n32883);
  and g54120 (n32889, pi1159, n_24238);
  not g54121 (n_24239, n32888);
  and g54122 (n32890, n_24239, n32889);
  not g54123 (n_24240, n32890);
  and g54124 (n32891, n_11403, n_24240);
  not g54125 (n_24241, n32882);
  and g54126 (n32892, n_24241, n32891);
  and g54127 (n32893, pi0619, n_24230);
  and g54128 (n32894, n_11821, n_24231);
  not g54129 (n_24242, n32894);
  and g54130 (n32895, pi1159, n_24242);
  not g54131 (n_24243, n32893);
  and g54132 (n32896, n_24243, n32895);
  and g54133 (n32897, n_11821, n32887);
  and g54134 (n32898, pi0619, n32727);
  not g54135 (n_24244, n32898);
  and g54136 (n32899, n_11405, n_24244);
  not g54137 (n_24245, n32897);
  and g54138 (n32900, n_24245, n32899);
  not g54139 (n_24246, n32900);
  and g54140 (n32901, pi0648, n_24246);
  not g54141 (n_24247, n32896);
  and g54142 (n32902, n_24247, n32901);
  not g54143 (n_24248, n32892);
  not g54144 (n_24249, n32902);
  and g54145 (n32903, n_24248, n_24249);
  not g54146 (n_24250, n32903);
  and g54147 (n32904, pi0789, n_24250);
  and g54148 (n32905, n_12315, n_24230);
  not g54149 (n_24251, n32904);
  not g54150 (n_24252, n32905);
  and g54151 (n32906, n_24251, n_24252);
  and g54152 (n32907, n_12318, n32906);
  and g54153 (n32908, n_12320, n32906);
  not g54154 (n_24253, n32756);
  and g54155 (n32909, pi0626, n_24253);
  not g54156 (n_24254, n32909);
  and g54157 (n32910, n_11395, n_24254);
  not g54158 (n_24255, n32908);
  and g54159 (n32911, n_24255, n32910);
  not g54160 (n_24256, n32887);
  and g54161 (n32912, n_12315, n_24256);
  and g54162 (n32913, n_24240, n_24246);
  not g54163 (n_24257, n32913);
  and g54164 (n32914, pi0789, n_24257);
  not g54165 (n_24258, n32912);
  not g54166 (n_24259, n32914);
  and g54167 (n32915, n_24258, n_24259);
  not g54168 (n_24260, n32915);
  and g54169 (n32916, n_12320, n_24260);
  and g54170 (n32917, pi0626, n_24111);
  not g54171 (n_24261, n32917);
  and g54172 (n32918, pi0641, n_24261);
  not g54173 (n_24262, n32916);
  and g54174 (n32919, n_24262, n32918);
  not g54175 (n_24263, n32919);
  and g54176 (n32920, n_11397, n_24263);
  not g54177 (n_24264, n32911);
  and g54178 (n32921, n_24264, n32920);
  and g54179 (n32922, pi0626, n32906);
  and g54180 (n32923, n_12320, n_24253);
  not g54181 (n_24265, n32923);
  and g54182 (n32924, pi0641, n_24265);
  not g54183 (n_24266, n32922);
  and g54184 (n32925, n_24266, n32924);
  and g54185 (n32926, pi0626, n_24260);
  and g54186 (n32927, n_12320, n_24111);
  not g54187 (n_24267, n32927);
  and g54188 (n32928, n_11395, n_24267);
  not g54189 (n_24268, n32926);
  and g54190 (n32929, n_24268, n32928);
  not g54191 (n_24269, n32929);
  and g54192 (n32930, pi1158, n_24269);
  not g54193 (n_24270, n32925);
  and g54194 (n32931, n_24270, n32930);
  not g54195 (n_24271, n32921);
  not g54196 (n_24272, n32931);
  and g54197 (n32932, n_24271, n_24272);
  not g54198 (n_24273, n32932);
  and g54199 (n32933, pi0788, n_24273);
  not g54200 (n_24274, n32907);
  not g54201 (n_24275, n32933);
  and g54202 (n32934, n_24274, n_24275);
  and g54203 (n32935, n_11789, n32934);
  and g54204 (n32936, n_12524, n32915);
  and g54205 (n32937, n17969, n32727);
  not g54206 (n_24276, n32936);
  not g54207 (n_24277, n32937);
  and g54208 (n32938, n_24276, n_24277);
  not g54209 (n_24278, n32938);
  and g54210 (n32939, pi0628, n_24278);
  not g54211 (n_24279, n32939);
  and g54212 (n32940, n_11794, n_24279);
  not g54213 (n_24280, n32935);
  and g54214 (n32941, n_24280, n32940);
  and g54215 (n32942, n_12354, n_24141);
  not g54216 (n_24281, n32941);
  and g54217 (n32943, n_24281, n32942);
  and g54218 (n32944, pi0628, n32934);
  and g54219 (n32945, n_11789, n_24278);
  not g54220 (n_24282, n32945);
  and g54221 (n32946, pi1156, n_24282);
  not g54222 (n_24283, n32944);
  and g54223 (n32947, n_24283, n32946);
  and g54224 (n32948, pi0629, n_24142);
  not g54225 (n_24284, n32947);
  and g54226 (n32949, n_24284, n32948);
  not g54227 (n_24285, n32943);
  not g54228 (n_24286, n32949);
  and g54229 (n32950, n_24285, n_24286);
  not g54230 (n_24287, n32950);
  and g54231 (n32951, pi0792, n_24287);
  and g54232 (n32952, n_11787, n32934);
  not g54233 (n_24288, n32951);
  not g54234 (n_24289, n32952);
  and g54235 (n32953, n_24288, n_24289);
  not g54236 (n_24290, n32953);
  and g54237 (n32954, n_11806, n_24290);
  and g54238 (n32955, n_12368, n_24278);
  and g54239 (n32956, n17779, n32727);
  not g54240 (n_24291, n32955);
  not g54241 (n_24292, n32956);
  and g54242 (n32957, n_24291, n_24292);
  not g54243 (n_24293, n32957);
  and g54244 (n32958, pi0647, n_24293);
  not g54245 (n_24294, n32958);
  and g54246 (n32959, n_11810, n_24294);
  not g54247 (n_24295, n32954);
  and g54248 (n32960, n_24295, n32959);
  and g54249 (n32961, n_12375, n_24151);
  not g54250 (n_24296, n32960);
  and g54251 (n32962, n_24296, n32961);
  and g54252 (n32963, pi0647, n_24290);
  and g54253 (n32964, n_11806, n_24293);
  not g54254 (n_24297, n32964);
  and g54255 (n32965, pi1157, n_24297);
  not g54256 (n_24298, n32963);
  and g54257 (n32966, n_24298, n32965);
  and g54258 (n32967, pi0630, n_24152);
  not g54259 (n_24299, n32966);
  and g54260 (n32968, n_24299, n32967);
  not g54261 (n_24300, n32962);
  not g54262 (n_24301, n32968);
  and g54263 (n32969, n_24300, n_24301);
  not g54264 (n_24302, n32969);
  and g54265 (n32970, pi0787, n_24302);
  and g54266 (n32971, n_11803, n_24290);
  not g54267 (n_24303, n32970);
  not g54268 (n_24304, n32971);
  and g54269 (n32972, n_24303, n_24304);
  not g54270 (n_24305, n32972);
  and g54271 (n32973, pi0644, n_24305);
  not g54272 (n_24306, n32784);
  and g54273 (n32974, pi0715, n_24306);
  not g54274 (n_24307, n32973);
  and g54275 (n32975, n_24307, n32974);
  and g54276 (n32976, n17804, n_24111);
  and g54277 (n32977, n_12392, n32957);
  not g54278 (n_24308, n32976);
  not g54279 (n_24309, n32977);
  and g54280 (n32978, n_24308, n_24309);
  and g54281 (n32979, pi0644, n32978);
  and g54282 (n32980, n_11819, n32727);
  not g54283 (n_24310, n32980);
  and g54284 (n32981, n_12395, n_24310);
  not g54285 (n_24311, n32979);
  and g54286 (n32982, n_24311, n32981);
  not g54287 (n_24312, n32982);
  and g54288 (n32983, pi1160, n_24312);
  not g54289 (n_24313, n32975);
  and g54290 (n32984, n_24313, n32983);
  and g54291 (n32985, n_11819, n_24305);
  and g54292 (n32986, pi0644, n32783);
  not g54293 (n_24314, n32986);
  and g54294 (n32987, n_12395, n_24314);
  not g54295 (n_24315, n32985);
  and g54296 (n32988, n_24315, n32987);
  and g54297 (n32989, n_11819, n32978);
  and g54298 (n32990, pi0644, n32727);
  not g54299 (n_24316, n32990);
  and g54300 (n32991, pi0715, n_24316);
  not g54301 (n_24317, n32989);
  and g54302 (n32992, n_24317, n32991);
  not g54303 (n_24318, n32992);
  and g54304 (n32993, n_12405, n_24318);
  not g54305 (n_24319, n32988);
  and g54306 (n32994, n_24319, n32993);
  not g54307 (n_24320, n32984);
  and g54308 (n32995, pi0790, n_24320);
  not g54309 (n_24321, n32994);
  and g54310 (n32996, n_24321, n32995);
  and g54311 (n32997, n_12411, n32972);
  not g54312 (n_24322, n32997);
  and g54313 (n32998, n_4226, n_24322);
  not g54314 (n_24323, n32996);
  and g54315 (n32999, n_24323, n32998);
  and g54316 (n33000, n_11115, po1038);
  not g54317 (n_24324, n33000);
  and g54318 (n33001, n_12415, n_24324);
  not g54319 (n_24325, n32999);
  and g54320 (n33002, n_24325, n33001);
  and g54321 (n33003, n_11115, n_12418);
  and g54322 (n33004, pi0730, n16645);
  not g54323 (n_24326, n33003);
  not g54324 (n_24327, n33004);
  and g54325 (n33005, n_24326, n_24327);
  and g54326 (n33006, n_11749, n33005);
  and g54327 (n33007, n_11753, n33004);
  not g54328 (n_24328, n33005);
  not g54329 (n_24329, n33007);
  and g54330 (n33008, n_24328, n_24329);
  not g54331 (n_24330, n33008);
  and g54332 (n33009, pi1153, n_24330);
  and g54333 (n33010, n_11757, n_24326);
  and g54334 (n33011, n_24329, n33010);
  not g54335 (n_24331, n33009);
  not g54336 (n_24332, n33011);
  and g54337 (n33012, n_24331, n_24332);
  not g54338 (n_24333, n33012);
  and g54339 (n33013, pi0778, n_24333);
  not g54340 (n_24334, n33006);
  not g54341 (n_24335, n33013);
  and g54342 (n33014, n_24334, n_24335);
  and g54343 (n33015, n_12429, n33014);
  and g54344 (n33016, n_12430, n33015);
  and g54345 (n33017, n_12431, n33016);
  and g54346 (n33018, n_12432, n33017);
  and g54347 (n33019, n_12436, n33018);
  and g54348 (n33020, n_11806, n33019);
  and g54349 (n33021, pi0647, n33003);
  not g54350 (n_24336, n33021);
  and g54351 (n33022, n_11810, n_24336);
  not g54352 (n_24337, n33020);
  and g54353 (n33023, n_24337, n33022);
  and g54354 (n33024, pi0630, n33023);
  and g54355 (n33025, pi0748, n17244);
  not g54356 (n_24338, n33025);
  and g54357 (n33026, n_24326, n_24338);
  not g54358 (n_24339, n33026);
  and g54359 (n33027, n_12448, n_24339);
  not g54360 (n_24340, n33027);
  and g54361 (n33028, n_11964, n_24340);
  and g54362 (n33029, n_12451, n_24339);
  not g54363 (n_24341, n33029);
  and g54364 (n33030, pi1155, n_24341);
  and g54365 (n33031, n_12453, n33027);
  not g54366 (n_24342, n33031);
  and g54367 (n33032, n_11768, n_24342);
  not g54368 (n_24343, n33030);
  not g54369 (n_24344, n33032);
  and g54370 (n33033, n_24343, n_24344);
  not g54371 (n_24345, n33033);
  and g54372 (n33034, pi0785, n_24345);
  not g54373 (n_24346, n33028);
  not g54374 (n_24347, n33034);
  and g54375 (n33035, n_24346, n_24347);
  not g54376 (n_24348, n33035);
  and g54377 (n33036, n_11981, n_24348);
  and g54378 (n33037, n_12461, n33035);
  not g54379 (n_24349, n33037);
  and g54380 (n33038, pi1154, n_24349);
  and g54381 (n33039, n_12463, n33035);
  not g54382 (n_24350, n33039);
  and g54383 (n33040, n_11413, n_24350);
  not g54384 (n_24351, n33038);
  not g54385 (n_24352, n33040);
  and g54386 (n33041, n_24351, n_24352);
  not g54387 (n_24353, n33041);
  and g54388 (n33042, pi0781, n_24353);
  not g54389 (n_24354, n33036);
  not g54390 (n_24355, n33042);
  and g54391 (n33043, n_24354, n_24355);
  not g54392 (n_24356, n33043);
  and g54393 (n33044, n_12315, n_24356);
  and g54394 (n33045, n_11821, n33003);
  and g54395 (n33046, pi0619, n33043);
  not g54396 (n_24357, n33045);
  and g54397 (n33047, pi1159, n_24357);
  not g54398 (n_24358, n33046);
  and g54399 (n33048, n_24358, n33047);
  and g54400 (n33049, n_11821, n33043);
  and g54401 (n33050, pi0619, n33003);
  not g54402 (n_24359, n33050);
  and g54403 (n33051, n_11405, n_24359);
  not g54404 (n_24360, n33049);
  and g54405 (n33052, n_24360, n33051);
  not g54406 (n_24361, n33048);
  not g54407 (n_24362, n33052);
  and g54408 (n33053, n_24361, n_24362);
  not g54409 (n_24363, n33053);
  and g54410 (n33054, pi0789, n_24363);
  not g54411 (n_24364, n33044);
  not g54412 (n_24365, n33054);
  and g54413 (n33055, n_24364, n_24365);
  and g54414 (n33056, n_12524, n33055);
  and g54415 (n33057, n17969, n33003);
  not g54416 (n_24366, n33056);
  not g54417 (n_24367, n33057);
  and g54418 (n33058, n_24366, n_24367);
  not g54419 (n_24368, n33058);
  and g54420 (n33059, n_12368, n_24368);
  and g54421 (n33060, n17779, n33003);
  not g54422 (n_24369, n33059);
  not g54423 (n_24370, n33060);
  and g54424 (n33061, n_24369, n_24370);
  and g54425 (n33062, n_14548, n33061);
  not g54426 (n_24371, n33019);
  and g54427 (n33063, pi0647, n_24371);
  and g54428 (n33064, n_11806, n_24326);
  not g54429 (n_24372, n33063);
  not g54430 (n_24373, n33064);
  and g54431 (n33065, n_24372, n_24373);
  not g54432 (n_24374, n33065);
  and g54433 (n33066, n17801, n_24374);
  not g54434 (n_24375, n33024);
  not g54435 (n_24376, n33066);
  and g54436 (n33067, n_24375, n_24376);
  not g54437 (n_24377, n33062);
  and g54438 (n33068, n_24377, n33067);
  not g54439 (n_24378, n33068);
  and g54440 (n33069, pi0787, n_24378);
  and g54441 (n33070, n17871, n33017);
  not g54442 (n_24379, n33055);
  and g54443 (n33071, n_12320, n_24379);
  and g54444 (n33072, pi0626, n_24326);
  not g54445 (n_24380, n33072);
  and g54446 (n33073, n16629, n_24380);
  not g54447 (n_24381, n33071);
  and g54448 (n33074, n_24381, n33073);
  and g54449 (n33075, pi0626, n_24379);
  and g54450 (n33076, n_12320, n_24326);
  not g54451 (n_24382, n33076);
  and g54452 (n33077, n16628, n_24382);
  not g54453 (n_24383, n33075);
  and g54454 (n33078, n_24383, n33077);
  not g54455 (n_24384, n33070);
  not g54456 (n_24385, n33074);
  and g54457 (n33079, n_24384, n_24385);
  not g54458 (n_24386, n33078);
  and g54459 (n33080, n_24386, n33079);
  not g54460 (n_24387, n33080);
  and g54461 (n33081, pi0788, n_24387);
  and g54462 (n33082, pi0618, n33015);
  and g54463 (n33083, pi0609, n33014);
  and g54464 (n33084, n_11866, n_24328);
  and g54465 (n33085, pi0625, n33084);
  not g54466 (n_24388, n33084);
  and g54467 (n33086, n33026, n_24388);
  not g54468 (n_24389, n33085);
  not g54469 (n_24390, n33086);
  and g54470 (n33087, n_24389, n_24390);
  not g54471 (n_24391, n33087);
  and g54472 (n33088, n33010, n_24391);
  and g54473 (n33089, n_11823, n_24331);
  not g54474 (n_24392, n33088);
  and g54475 (n33090, n_24392, n33089);
  and g54476 (n33091, pi1153, n33026);
  and g54477 (n33092, n_24389, n33091);
  and g54478 (n33093, pi0608, n_24332);
  not g54479 (n_24393, n33092);
  and g54480 (n33094, n_24393, n33093);
  not g54481 (n_24394, n33090);
  not g54482 (n_24395, n33094);
  and g54483 (n33095, n_24394, n_24395);
  not g54484 (n_24396, n33095);
  and g54485 (n33096, pi0778, n_24396);
  and g54486 (n33097, n_11749, n_24390);
  not g54487 (n_24397, n33096);
  not g54488 (n_24398, n33097);
  and g54489 (n33098, n_24397, n_24398);
  not g54490 (n_24399, n33098);
  and g54491 (n33099, n_11971, n_24399);
  not g54492 (n_24400, n33083);
  and g54493 (n33100, n_11768, n_24400);
  not g54494 (n_24401, n33099);
  and g54495 (n33101, n_24401, n33100);
  and g54496 (n33102, n_11767, n_24343);
  not g54497 (n_24402, n33101);
  and g54498 (n33103, n_24402, n33102);
  and g54499 (n33104, n_11971, n33014);
  and g54500 (n33105, pi0609, n_24399);
  not g54501 (n_24403, n33104);
  and g54502 (n33106, pi1155, n_24403);
  not g54503 (n_24404, n33105);
  and g54504 (n33107, n_24404, n33106);
  and g54505 (n33108, pi0660, n_24344);
  not g54506 (n_24405, n33107);
  and g54507 (n33109, n_24405, n33108);
  not g54508 (n_24406, n33103);
  not g54509 (n_24407, n33109);
  and g54510 (n33110, n_24406, n_24407);
  not g54511 (n_24408, n33110);
  and g54512 (n33111, pi0785, n_24408);
  and g54513 (n33112, n_11964, n_24399);
  not g54514 (n_24409, n33111);
  not g54515 (n_24410, n33112);
  and g54516 (n33113, n_24409, n_24410);
  not g54517 (n_24411, n33113);
  and g54518 (n33114, n_11984, n_24411);
  not g54519 (n_24412, n33082);
  and g54520 (n33115, n_11413, n_24412);
  not g54521 (n_24413, n33114);
  and g54522 (n33116, n_24413, n33115);
  and g54523 (n33117, n_11412, n_24351);
  not g54524 (n_24414, n33116);
  and g54525 (n33118, n_24414, n33117);
  and g54526 (n33119, n_11984, n33015);
  and g54527 (n33120, pi0618, n_24411);
  not g54528 (n_24415, n33119);
  and g54529 (n33121, pi1154, n_24415);
  not g54530 (n_24416, n33120);
  and g54531 (n33122, n_24416, n33121);
  and g54532 (n33123, pi0627, n_24352);
  not g54533 (n_24417, n33122);
  and g54534 (n33124, n_24417, n33123);
  not g54535 (n_24418, n33118);
  not g54536 (n_24419, n33124);
  and g54537 (n33125, n_24418, n_24419);
  not g54538 (n_24420, n33125);
  and g54539 (n33126, pi0781, n_24420);
  and g54540 (n33127, n_11981, n_24411);
  not g54541 (n_24421, n33126);
  not g54542 (n_24422, n33127);
  and g54543 (n33128, n_24421, n_24422);
  and g54544 (n33129, n_12315, n33128);
  not g54545 (n_24423, n33128);
  and g54546 (n33130, n_11821, n_24423);
  and g54547 (n33131, pi0619, n33016);
  not g54548 (n_24424, n33131);
  and g54549 (n33132, n_11405, n_24424);
  not g54550 (n_24425, n33130);
  and g54551 (n33133, n_24425, n33132);
  and g54552 (n33134, n_11403, n_24361);
  not g54553 (n_24426, n33133);
  and g54554 (n33135, n_24426, n33134);
  and g54555 (n33136, pi0619, n_24423);
  and g54556 (n33137, n_11821, n33016);
  not g54557 (n_24427, n33137);
  and g54558 (n33138, pi1159, n_24427);
  not g54559 (n_24428, n33136);
  and g54560 (n33139, n_24428, n33138);
  and g54561 (n33140, pi0648, n_24362);
  not g54562 (n_24429, n33139);
  and g54563 (n33141, n_24429, n33140);
  not g54564 (n_24430, n33135);
  and g54565 (n33142, pi0789, n_24430);
  not g54566 (n_24431, n33141);
  and g54567 (n33143, n_24431, n33142);
  not g54568 (n_24432, n33129);
  and g54569 (n33144, n17970, n_24432);
  not g54570 (n_24433, n33143);
  and g54571 (n33145, n_24433, n33144);
  not g54572 (n_24434, n33081);
  not g54573 (n_24435, n33145);
  and g54574 (n33146, n_24434, n_24435);
  not g54575 (n_24436, n33146);
  and g54576 (n33147, n_14638, n_24436);
  and g54577 (n33148, n17854, n_24368);
  and g54578 (n33149, n20851, n33018);
  not g54579 (n_24437, n33148);
  not g54580 (n_24438, n33149);
  and g54581 (n33150, n_24437, n_24438);
  not g54582 (n_24439, n33150);
  and g54583 (n33151, n_12354, n_24439);
  and g54584 (n33152, n20855, n33018);
  and g54585 (n33153, n17853, n_24368);
  not g54586 (n_24440, n33152);
  not g54587 (n_24441, n33153);
  and g54588 (n33154, n_24440, n_24441);
  not g54589 (n_24442, n33154);
  and g54590 (n33155, pi0629, n_24442);
  not g54591 (n_24443, n33151);
  not g54592 (n_24444, n33155);
  and g54593 (n33156, n_24443, n_24444);
  not g54594 (n_24445, n33156);
  and g54595 (n33157, pi0792, n_24445);
  not g54596 (n_24446, n33157);
  and g54597 (n33158, n_14387, n_24446);
  not g54598 (n_24447, n33147);
  and g54599 (n33159, n_24447, n33158);
  not g54600 (n_24448, n33069);
  not g54601 (n_24449, n33159);
  and g54602 (n33160, n_24448, n_24449);
  and g54603 (n33161, n_12411, n33160);
  and g54604 (n33162, n_11803, n_24371);
  and g54605 (n33163, pi1157, n_24374);
  not g54606 (n_24450, n33023);
  not g54607 (n_24451, n33163);
  and g54608 (n33164, n_24450, n_24451);
  not g54609 (n_24452, n33164);
  and g54610 (n33165, pi0787, n_24452);
  not g54611 (n_24453, n33162);
  not g54612 (n_24454, n33165);
  and g54613 (n33166, n_24453, n_24454);
  and g54614 (n33167, n_11819, n33166);
  and g54615 (n33168, pi0644, n33160);
  not g54616 (n_24455, n33167);
  and g54617 (n33169, pi0715, n_24455);
  not g54618 (n_24456, n33168);
  and g54619 (n33170, n_24456, n33169);
  not g54620 (n_24457, n33061);
  and g54621 (n33171, n_12392, n_24457);
  and g54622 (n33172, n17804, n33003);
  not g54623 (n_24458, n33171);
  not g54624 (n_24459, n33172);
  and g54625 (n33173, n_24458, n_24459);
  not g54626 (n_24460, n33173);
  and g54627 (n33174, pi0644, n_24460);
  and g54628 (n33175, n_11819, n33003);
  not g54629 (n_24461, n33175);
  and g54630 (n33176, n_12395, n_24461);
  not g54631 (n_24462, n33174);
  and g54632 (n33177, n_24462, n33176);
  not g54633 (n_24463, n33177);
  and g54634 (n33178, pi1160, n_24463);
  not g54635 (n_24464, n33170);
  and g54636 (n33179, n_24464, n33178);
  and g54637 (n33180, n_11819, n_24460);
  and g54638 (n33181, pi0644, n33003);
  not g54639 (n_24465, n33181);
  and g54640 (n33182, pi0715, n_24465);
  not g54641 (n_24466, n33180);
  and g54642 (n33183, n_24466, n33182);
  and g54643 (n33184, pi0644, n33166);
  and g54644 (n33185, n_11819, n33160);
  not g54645 (n_24467, n33184);
  and g54646 (n33186, n_12395, n_24467);
  not g54647 (n_24468, n33185);
  and g54648 (n33187, n_24468, n33186);
  not g54649 (n_24469, n33183);
  and g54650 (n33188, n_12405, n_24469);
  not g54651 (n_24470, n33187);
  and g54652 (n33189, n_24470, n33188);
  not g54653 (n_24471, n33179);
  not g54654 (n_24472, n33189);
  and g54655 (n33190, n_24471, n_24472);
  not g54656 (n_24473, n33190);
  and g54657 (n33191, pi0790, n_24473);
  not g54658 (n_24474, n33161);
  and g54659 (n33192, pi0832, n_24474);
  not g54660 (n_24475, n33191);
  and g54661 (n33193, n_24475, n33192);
  not g54662 (n_24476, n33002);
  not g54663 (n_24477, n33193);
  and g54664 (po0351, n_24476, n_24477);
  and g54665 (n33195, n_5671, n16565);
  and g54666 (n33196, n_5669, n33195);
  not g54667 (n_24478, n33196);
  and g54668 (n33197, pi0195, n_24478);
  and g54669 (n33198, n_7426, n16193);
  and g54670 (n33199, n_3120, n16168);
  and g54671 (n33200, n16167, n_11279);
  not g54678 (n_24482, n33203);
  and g54679 (n33204, pi0232, n_24482);
  not g54680 (n_24483, n33204);
  and g54681 (n33205, n_11284, n_24483);
  not g54682 (n_24484, n33205);
  and g54683 (n33206, pi0039, n_24484);
  and g54684 (n33207, n13910, n_11023);
  not g54685 (n_24485, n33207);
  and g54686 (n33208, n_162, n_24485);
  and g54693 (n33212, n_1493, n9326);
  not g54694 (n_24489, n33212);
  and g54695 (n33213, n_11303, n_24489);
  not g54696 (n_24490, n33213);
  and g54697 (n33214, n9036, n_24490);
  not g54698 (n_24491, n33214);
  and g54699 (n33215, n9291, n_24491);
  and g54700 (n33216, n_11043, n16511);
  and g54701 (n33217, pi0192, n16520);
  not g54702 (n_24492, n33215);
  not g54703 (n_24493, n33216);
  and g54704 (n33218, n_24492, n_24493);
  not g54705 (n_24494, n33217);
  and g54706 (n33219, n_24494, n33218);
  not g54707 (n_24495, n33219);
  and g54708 (n33220, pi0232, n_24495);
  not g54709 (n_24496, n33220);
  and g54710 (n33221, n_11311, n_24496);
  not g54711 (n_24497, n33221);
  and g54712 (n33222, pi0039, n_24497);
  and g54713 (n33223, pi0192, n16539);
  and g54714 (n33224, n_11314, n_11031);
  and g54715 (n33225, pi0171, n13737);
  not g54716 (n_24498, n33224);
  not g54717 (n_24499, n33225);
  and g54718 (n33226, n_24498, n_24499);
  not g54719 (n_24500, n33226);
  and g54720 (n33227, pi0299, n_24500);
  and g54721 (n33228, n_11043, n16533);
  not g54728 (n_24504, n33231);
  and g54729 (n33232, n16536, n_24504);
  not g54730 (n_24505, n33222);
  and g54731 (n33233, n2608, n_24505);
  not g54732 (n_24506, n33232);
  and g54733 (n33234, n_24506, n33233);
  not g54734 (n_24507, n33234);
  and g54735 (n33235, n_172, n_24507);
  not g54736 (n_24508, n33235);
  and g54737 (n33236, n16508, n_24508);
  not g54738 (n_24509, n33236);
  and g54739 (n33237, n_174, n_24509);
  not g54740 (n_24510, n33237);
  and g54741 (n33238, n16507, n_24510);
  not g54742 (n_24511, n33238);
  and g54743 (n33239, n_176, n_24511);
  not g54744 (n_24512, n33239);
  and g54745 (n33240, n_11338, n_24512);
  not g54746 (n_24513, n33240);
  and g54747 (n33241, n2529, n_24513);
  and g54748 (n33242, n9883, n33197);
  not g54749 (n_24514, n33241);
  and g54750 (n33243, n_24514, n33242);
  or g54751 (po0352, n33211, n33243);
  and g54752 (n33245, n13132, n16492);
  and g54753 (n33246, n_1673, n9039);
  not g54754 (n_24515, n16492);
  not g54755 (n_24516, n33246);
  and g54756 (n33247, n_24515, n_24516);
  not g54757 (n_24517, n33247);
  and g54758 (n33248, n13130, n_24517);
  not g54759 (n_24518, n33245);
  and g54760 (n33249, pi0232, n_24518);
  not g54761 (n_24519, n33248);
  and g54762 (n33250, n_24519, n33249);
  not g54763 (n_24520, n33250);
  and g54764 (n33251, n_11284, n_24520);
  not g54765 (n_24521, n33251);
  and g54766 (n33252, pi0039, n_24521);
  and g54767 (n33253, n13910, n16287);
  not g54768 (n_24522, n33253);
  and g54769 (n33254, n_162, n_24522);
  not g54770 (n_24523, n33254);
  and g54771 (n33255, n_161, n_24523);
  not g54772 (n_24524, n33252);
  and g54773 (n33256, n_24524, n33255);
  not g54774 (n_24525, n33256);
  and g54775 (n33257, pi0194, n_24525);
  and g54776 (n33258, pi0299, n_24521);
  not g54777 (n_24526, n33258);
  and g54778 (n33259, n_7428, n_24526);
  not g54779 (n_24527, n33259);
  and g54780 (n33260, pi0039, n_24527);
  and g54781 (n33261, n13910, n_11111);
  not g54782 (n_24528, n33261);
  and g54783 (n33262, n_162, n_24528);
  not g54784 (n_24529, n33262);
  and g54785 (n33263, n_161, n_24529);
  not g54786 (n_24530, n33260);
  and g54787 (n33264, n_24530, n33263);
  not g54788 (n_24531, n33264);
  and g54789 (n33265, n_11115, n_24531);
  not g54790 (n_24532, n33257);
  and g54791 (n33266, n10197, n_24532);
  not g54792 (n_24533, n33265);
  and g54793 (n33267, n_24533, n33266);
  not g54794 (n_24534, n33267);
  and g54795 (n33268, n_5669, n_24534);
  and g54796 (n33269, n_1673, n9326);
  not g54797 (n_24535, n33269);
  and g54798 (n33270, n_11303, n_24535);
  not g54799 (n_24536, n33270);
  and g54800 (n33271, n9036, n_24536);
  not g54801 (n_24537, n33271);
  and g54802 (n33272, n9291, n_24537);
  not g54803 (n_24538, n33272);
  and g54804 (n33273, n_11299, n_24538);
  not g54805 (n_24539, n33273);
  and g54806 (n33274, pi0232, n_24539);
  not g54807 (n_24540, n33274);
  and g54808 (n33275, n_11311, n_24540);
  and g54809 (n33276, pi0232, n16520);
  not g54810 (n_24541, n33276);
  and g54811 (n33277, n33275, n_24541);
  not g54812 (n_24542, n33277);
  and g54813 (n33278, pi0039, n_24542);
  and g54814 (n33279, n_161, pi0194);
  not g54815 (n_24543, n33278);
  and g54816 (n33280, n_24543, n33279);
  not g54817 (n_24544, n33275);
  and g54818 (n33281, pi0039, n_24544);
  and g54819 (n33282, n_161, n_11115);
  not g54820 (n_24545, n33281);
  and g54821 (n33283, n_24545, n33282);
  not g54822 (n_24546, n33280);
  not g54823 (n_24547, n33283);
  and g54824 (n33284, n_24546, n_24547);
  not g54825 (n_24548, n16536);
  not g54826 (n_24549, n33284);
  and g54827 (n33285, n_24548, n_24549);
  and g54828 (n33286, n_11314, n_11125);
  and g54829 (n33287, pi0170, n13737);
  not g54830 (n_24550, n33286);
  not g54831 (n_24551, n33287);
  and g54832 (n33288, n_24550, n_24551);
  not g54833 (n_24552, n33288);
  and g54834 (n33289, pi0299, n_24552);
  not g54835 (n_24553, n16539);
  and g54836 (n33290, n_24553, n33280);
  and g54837 (n33291, n_11316, n33283);
  not g54838 (n_24554, n33290);
  not g54839 (n_24555, n33291);
  and g54840 (n33292, n_24554, n_24555);
  not g54841 (n_24556, n33289);
  and g54842 (n33293, pi0232, n_24556);
  not g54843 (n_24557, n33292);
  and g54844 (n33294, n_24557, n33293);
  not g54845 (n_24558, n33285);
  not g54846 (n_24559, n33294);
  and g54847 (n33295, n_24558, n_24559);
  not g54848 (n_24560, n33295);
  and g54849 (n33296, n_164, n_24560);
  not g54850 (n_24561, n33296);
  and g54851 (n33297, n_172, n_24561);
  not g54852 (n_24562, n33297);
  and g54853 (n33298, n16508, n_24562);
  not g54854 (n_24563, n33298);
  and g54855 (n33299, n_174, n_24563);
  not g54856 (n_24564, n33299);
  and g54857 (n33300, n16507, n_24564);
  not g54858 (n_24565, n33300);
  and g54859 (n33301, n_176, n_24565);
  not g54860 (n_24566, n33301);
  and g54861 (n33302, n_11338, n_24566);
  not g54862 (n_24567, n33302);
  and g54863 (n33303, n2529, n_24567);
  not g54864 (n_24568, n33303);
  and g54865 (n33304, n9883, n_24568);
  not g54866 (n_24569, n33304);
  and g54867 (n33305, pi0196, n_24569);
  not g54868 (n_24570, n33195);
  not g54869 (n_24571, n33268);
  and g54870 (n33306, n_24570, n_24571);
  not g54871 (n_24572, n33305);
  and g54872 (n33307, n_24572, n33306);
  and g54873 (n33308, pi0195, n_5669);
  not g54874 (n_24573, n33308);
  and g54875 (n33309, n_24534, n_24573);
  and g54876 (n33310, n_24569, n33308);
  not g54877 (n_24574, n33309);
  and g54878 (n33311, n33195, n_24574);
  not g54879 (n_24575, n33310);
  and g54880 (n33312, n_24575, n33311);
  or g54881 (po0353, n33307, n33312);
  and g54882 (n33314, n_6219, n_12418);
  and g54883 (n33315, n_14479, pi0947);
  and g54884 (n33316, n_14424, n20902);
  not g54885 (n_24576, n33315);
  not g54886 (n_24577, n33316);
  and g54887 (n33317, n_24576, n_24577);
  not g54888 (n_24578, n33317);
  and g54889 (n33318, n2926, n_24578);
  not g54890 (n_24579, n33314);
  and g54891 (n33319, pi0832, n_24579);
  not g54892 (n_24580, n33318);
  and g54893 (n33320, n_24580, n33319);
  and g54894 (n33321, n_6219, n_14814);
  and g54895 (n33322, n16641, n_24576);
  and g54896 (n33323, pi0197, n_11740);
  not g54897 (n_24581, n33322);
  and g54898 (n33324, pi0038, n_24581);
  not g54899 (n_24582, n33323);
  and g54900 (n33325, n_24582, n33324);
  and g54901 (n33326, n_6219, n_11674);
  and g54902 (n33327, n16958, n33315);
  not g54903 (n_24583, n33326);
  and g54904 (n33328, n_162, n_24583);
  not g54905 (n_24584, n33327);
  and g54906 (n33329, n_24584, n33328);
  and g54907 (n33330, n_6219, n_14891);
  and g54908 (n33331, pi0197, n_15009);
  not g54909 (n_24585, n33331);
  and g54910 (n33332, pi0299, n_24585);
  not g54911 (n_24586, n33330);
  and g54912 (n33333, n_24586, n33332);
  and g54913 (n33334, n_6219, n_11719);
  not g54914 (n_24587, n33334);
  and g54915 (n33335, n21019, n_24587);
  not g54916 (n_24588, n33335);
  and g54917 (n33336, n_14479, n_24588);
  not g54918 (n_24589, n33333);
  and g54919 (n33337, n_24589, n33336);
  and g54920 (n33338, n_6219, pi0767);
  and g54921 (n33339, n_11736, n33338);
  not g54922 (n_24590, n33339);
  and g54923 (n33340, pi0039, n_24590);
  not g54924 (n_24591, n33337);
  and g54925 (n33341, n_24591, n33340);
  not g54926 (n_24592, n33329);
  and g54927 (n33342, n_161, n_24592);
  not g54928 (n_24593, n33341);
  and g54929 (n33343, n_24593, n33342);
  not g54930 (n_24594, n33325);
  not g54931 (n_24595, n33343);
  and g54932 (n33344, n_24594, n_24595);
  not g54933 (n_24596, n33344);
  and g54934 (n33345, pi0698, n_24596);
  and g54935 (n33346, n_14975, n33329);
  and g54936 (n33347, n21111, n_24587);
  and g54937 (n33348, pi0197, n21108);
  and g54938 (n33349, n_6219, n21092);
  not g54939 (n_24597, n33348);
  and g54940 (n33350, pi0299, n_24597);
  not g54941 (n_24598, n33349);
  and g54942 (n33351, n_24598, n33350);
  not g54943 (n_24599, n33347);
  and g54944 (n33352, pi0767, n_24599);
  not g54945 (n_24600, n33351);
  and g54946 (n33353, n_24600, n33352);
  and g54947 (n33354, n_6219, n21064);
  and g54948 (n33355, pi0197, n21080);
  not g54949 (n_24601, n33355);
  and g54950 (n33356, n_14479, n_24601);
  not g54951 (n_24602, n33354);
  and g54952 (n33357, n_24602, n33356);
  not g54953 (n_24603, n33353);
  and g54954 (n33358, pi0039, n_24603);
  not g54955 (n_24604, n33357);
  and g54956 (n33359, n_24604, n33358);
  not g54957 (n_24605, n33346);
  not g54958 (n_24606, n33359);
  and g54959 (n33360, n_24605, n_24606);
  not g54960 (n_24607, n33360);
  and g54961 (n33361, n_161, n_24607);
  and g54962 (n33362, n_6219, n_11418);
  and g54963 (n33363, pi0767, pi0947);
  not g54964 (n_24608, n33363);
  and g54965 (n33364, n_162, n_24608);
  and g54966 (n33365, n21239, n33364);
  not g54967 (n_24609, n33362);
  and g54968 (n33366, pi0038, n_24609);
  not g54969 (n_24610, n33365);
  and g54970 (n33367, n_24610, n33366);
  not g54971 (n_24611, n33367);
  and g54972 (n33368, n_14424, n_24611);
  not g54973 (n_24612, n33361);
  and g54974 (n33369, n_24612, n33368);
  not g54975 (n_24613, n33345);
  not g54976 (n_24614, n33369);
  and g54977 (n33370, n_24613, n_24614);
  not g54978 (n_24615, n33370);
  and g54979 (n33371, n10197, n_24615);
  not g54980 (n_24616, n33321);
  and g54981 (n33372, n_12415, n_24616);
  not g54982 (n_24617, n33371);
  and g54983 (n33373, n_24617, n33372);
  not g54984 (n_24618, n33320);
  not g54985 (n_24619, n33373);
  and g54986 (po0354, n_24618, n_24619);
  and g54987 (n33375, n2530, n_11674);
  not g54988 (n_24620, n33375);
  and g54989 (n33376, n18591, n_24620);
  not g54990 (n_24621, n33376);
  and g54991 (n33377, pi0198, n_24621);
  and g54992 (n33378, pi0198, n_11543);
  and g54993 (n33379, pi0198, n_11445);
  not g54994 (n_24622, po1101);
  not g54995 (n_24623, n33379);
  and g54996 (n33380, n_24622, n_24623);
  not g54997 (n_24624, n33380);
  and g54998 (n33381, n33378, n_24624);
  and g54999 (n33382, n6192, n_11479);
  and g55000 (n33383, n_3138, n_11556);
  not g55001 (n_24625, n33382);
  and g55002 (n33384, pi0198, n_24625);
  not g55003 (n_24626, n33383);
  and g55004 (n33385, n_24626, n33384);
  and g55005 (n33386, n_3162, n33385);
  not g55006 (n_24627, n33381);
  not g55007 (n_24628, n33386);
  and g55008 (n33387, n_24627, n_24628);
  not g55009 (n_24629, n33387);
  and g55010 (n33388, pi0215, n_24629);
  and g55011 (n33389, n3448, n_24623);
  and g55012 (n33390, pi0198, n_11513);
  not g55013 (n_24630, n33390);
  and g55014 (n33391, po1101, n_24630);
  not g55015 (n_24631, n33391);
  and g55016 (n33392, n_24624, n_24631);
  and g55017 (n33393, n6242, n33392);
  not g55018 (n_24632, n17143);
  and g55019 (n33394, pi0198, n_24632);
  and g55020 (n33395, n_3162, n33394);
  not g55021 (n_24633, n33393);
  and g55022 (n33396, n_9350, n_24633);
  not g55023 (n_24634, n33395);
  and g55024 (n33397, n_24634, n33396);
  not g55025 (n_24635, n33389);
  and g55026 (n33398, n_36, n_24635);
  not g55027 (n_24636, n33397);
  and g55028 (n33399, n_24636, n33398);
  not g55029 (n_24637, n33388);
  and g55030 (n33400, pi0299, n_24637);
  not g55031 (n_24638, n33399);
  and g55032 (n33401, n_24638, n33400);
  and g55033 (n33402, n_3119, n33385);
  not g55034 (n_24639, n33402);
  and g55035 (n33403, n_24627, n_24639);
  not g55036 (n_24640, n33403);
  and g55037 (n33404, pi0223, n_24640);
  and g55038 (n33405, n2603, n_24623);
  and g55039 (n33406, n_3119, n33394);
  and g55040 (n33407, n6205, n33392);
  not g55041 (n_24641, n33407);
  and g55042 (n33408, n_9349, n_24641);
  not g55043 (n_24642, n33406);
  and g55044 (n33409, n_24642, n33408);
  not g55045 (n_24643, n33405);
  and g55046 (n33410, n_223, n_24643);
  not g55047 (n_24644, n33409);
  and g55048 (n33411, n_24644, n33410);
  not g55049 (n_24645, n33404);
  and g55050 (n33412, n_234, n_24645);
  not g55051 (n_24646, n33411);
  and g55052 (n33413, n_24646, n33412);
  not g55058 (n_24649, n33377);
  not g55059 (n_24650, n33416);
  and g55060 (n33417, n_24649, n_24650);
  not g55061 (n_24651, n19149);
  and g55062 (n33418, n_24651, n33417);
  not g55063 (n_24652, n33417);
  and g55064 (n33419, n16639, n_24652);
  and g55065 (n33420, pi0198, n_11417);
  and g55066 (n33421, pi0039, pi0198);
  not g55067 (n_24653, n33421);
  and g55068 (n33422, pi0038, n_24653);
  and g55069 (n33423, pi0198, n_11432);
  and g55070 (n33424, pi0634, n16644);
  and g55071 (n33425, n16667, n33424);
  not g55072 (n_24655, n33423);
  not g55073 (n_24656, n33425);
  and g55074 (n33426, n_24655, n_24656);
  not g55075 (n_24657, n33426);
  and g55076 (n33427, n_162, n_24657);
  not g55077 (n_24658, n33427);
  and g55078 (n33428, n33422, n_24658);
  and g55079 (n33429, pi0198, n16721);
  and g55080 (n33430, pi0634, n_11479);
  and g55081 (n33431, n16658, n33430);
  not g55082 (n_24659, n33429);
  not g55083 (n_24660, n33431);
  and g55084 (n33432, n_24659, n_24660);
  not g55085 (n_24661, n33432);
  and g55086 (n33433, n6195, n_24661);
  and g55087 (n33434, n_11502, n33385);
  and g55088 (n33435, n6192, n33432);
  and g55089 (n33436, n_11450, n_24623);
  not g55090 (n_24662, n33436);
  and g55091 (n33437, pi0634, n_24662);
  not g55092 (n_24663, n33437);
  and g55093 (n33438, n_24623, n_24663);
  and g55094 (n33439, n_3102, n33438);
  and g55095 (n33440, n6197, n33432);
  not g55096 (n_24664, n33439);
  not g55097 (n_24665, n33440);
  and g55098 (n33441, n_24664, n_24665);
  not g55099 (n_24666, n33441);
  and g55100 (n33442, n_3138, n_24666);
  not g55101 (n_24667, n33435);
  and g55102 (n33443, n17323, n_24667);
  not g55103 (n_24668, n33442);
  and g55104 (n33444, n_24668, n33443);
  not g55105 (n_24669, n33433);
  not g55106 (n_24670, n33434);
  and g55107 (n33445, n_24669, n_24670);
  not g55108 (n_24671, n33444);
  and g55109 (n33446, n_24671, n33445);
  and g55110 (n33447, n_3119, n33446);
  and g55111 (n33448, n33378, n33434);
  not g55112 (n_24672, n33438);
  and g55113 (n33449, n6197, n_24672);
  and g55114 (n33450, n_3102, n_24661);
  not g55115 (n_24673, n33449);
  not g55116 (n_24674, n33450);
  and g55117 (n33451, n_24673, n_24674);
  and g55118 (n33452, n6192, n33451);
  and g55119 (n33453, n_3138, n33438);
  not g55120 (n_24675, n33453);
  and g55121 (n33454, n17323, n_24675);
  not g55122 (n_24676, n33452);
  and g55123 (n33455, n_24676, n33454);
  not g55124 (n_24677, n33451);
  and g55125 (n33456, n6195, n_24677);
  not g55126 (n_24678, n33448);
  not g55127 (n_24679, n33456);
  and g55128 (n33457, n_24678, n_24679);
  not g55129 (n_24680, n33455);
  and g55130 (n33458, n_24680, n33457);
  and g55131 (n33459, n6205, n33458);
  not g55132 (n_24681, n33447);
  and g55133 (n33460, pi0223, n_24681);
  not g55134 (n_24682, n33459);
  and g55135 (n33461, n_24682, n33460);
  and g55136 (n33462, pi0680, n33437);
  not g55137 (n_24683, n33462);
  and g55138 (n33463, n_24623, n_24683);
  and g55139 (n33464, n2603, n33463);
  and g55140 (n33465, pi0198, n16681);
  and g55141 (n33466, pi0634, n16686);
  not g55142 (n_24684, n33465);
  not g55143 (n_24685, n33466);
  and g55144 (n33467, n_24684, n_24685);
  not g55145 (n_24686, n33467);
  and g55146 (n33468, n_3102, n_24686);
  not g55147 (n_24687, n33468);
  and g55148 (n33469, n_24673, n_24687);
  not g55149 (n_24688, n33469);
  and g55150 (n33470, n6195, n_24688);
  and g55151 (n33471, n6192, n33469);
  not g55152 (n_24689, n33471);
  and g55153 (n33472, n33454, n_24689);
  and g55154 (n33473, n_3138, n_24623);
  and g55155 (n33474, n6192, n_24630);
  not g55156 (n_24690, n33473);
  and g55157 (n33475, n_11502, n_24690);
  not g55158 (n_24691, n33474);
  and g55159 (n33476, n_24691, n33475);
  not g55160 (n_24692, n33470);
  not g55161 (n_24693, n33476);
  and g55162 (n33477, n_24692, n_24693);
  not g55163 (n_24694, n33472);
  and g55164 (n33478, n_24694, n33477);
  not g55165 (n_24695, n33478);
  and g55166 (n33479, n6205, n_24695);
  and g55167 (n33480, pi0198, n16753);
  and g55168 (n33481, n6195, n_24686);
  and g55169 (n33482, n6192, n33467);
  and g55170 (n33483, n6197, n33467);
  not g55171 (n_24696, n33483);
  and g55172 (n33484, n_24664, n_24696);
  not g55173 (n_24697, n33484);
  and g55174 (n33485, n_3138, n_24697);
  not g55175 (n_24698, n33482);
  and g55176 (n33486, n17323, n_24698);
  not g55177 (n_24699, n33485);
  and g55178 (n33487, n_24699, n33486);
  not g55179 (n_24700, n33480);
  not g55180 (n_24701, n33481);
  and g55181 (n33488, n_24700, n_24701);
  not g55182 (n_24702, n33487);
  and g55183 (n33489, n_24702, n33488);
  not g55184 (n_24703, n33489);
  and g55185 (n33490, n_3119, n_24703);
  not g55186 (n_24704, n33479);
  and g55187 (n33491, n_9349, n_24704);
  not g55188 (n_24705, n33490);
  and g55189 (n33492, n_24705, n33491);
  not g55190 (n_24706, n33464);
  and g55191 (n33493, n_223, n_24706);
  not g55192 (n_24707, n33492);
  and g55193 (n33494, n_24707, n33493);
  not g55194 (n_24708, n33461);
  and g55195 (n33495, n_234, n_24708);
  not g55196 (n_24709, n33494);
  and g55197 (n33496, n_24709, n33495);
  and g55198 (n33497, n_3162, n33446);
  and g55199 (n33498, n6242, n33458);
  not g55200 (n_24710, n33497);
  and g55201 (n33499, pi0215, n_24710);
  not g55202 (n_24711, n33498);
  and g55203 (n33500, n_24711, n33499);
  and g55204 (n33501, n3448, n33463);
  and g55205 (n33502, n_3162, n_24703);
  and g55206 (n33503, n6242, n_24695);
  not g55207 (n_24712, n33502);
  and g55208 (n33504, n_9350, n_24712);
  not g55209 (n_24713, n33503);
  and g55210 (n33505, n_24713, n33504);
  not g55211 (n_24714, n33501);
  and g55212 (n33506, n_36, n_24714);
  not g55213 (n_24715, n33505);
  and g55214 (n33507, n_24715, n33506);
  not g55215 (n_24716, n33500);
  and g55216 (n33508, pi0299, n_24716);
  not g55217 (n_24717, n33507);
  and g55218 (n33509, n_24717, n33508);
  not g55219 (n_24718, n33496);
  not g55220 (n_24719, n33509);
  and g55221 (n33510, n_24718, n_24719);
  not g55222 (n_24720, n33510);
  and g55223 (n33511, pi0039, n_24720);
  and g55224 (n33512, pi0634, pi0680);
  and g55225 (n33513, pi0198, n16931);
  and g55226 (n33514, n_11634, n33512);
  not g55227 (n_24721, n33513);
  and g55228 (n33515, n_24721, n33514);
  not g55229 (n_24722, n33515);
  and g55230 (n33516, n_11643, n_24722);
  not g55231 (n_24723, n33516);
  and g55232 (n33517, n_234, n_24723);
  and g55233 (n33518, n_305, n16923);
  and g55234 (n33519, pi0198, n_11655);
  not g55235 (n_24724, n33518);
  not g55236 (n_24725, n33519);
  and g55237 (n33520, n_24724, n_24725);
  not g55238 (n_24726, n33520);
  and g55239 (n33521, n33512, n_24726);
  and g55240 (n33522, pi0198, n_11670);
  not g55241 (n_24727, n33512);
  and g55242 (n33523, n_24727, n33522);
  not g55243 (n_24728, n33521);
  not g55244 (n_24729, n33523);
  and g55245 (n33524, n_24728, n_24729);
  not g55246 (n_24730, n33524);
  and g55247 (n33525, pi0299, n_24730);
  not g55248 (n_24731, n33517);
  and g55249 (n33526, n_162, n_24731);
  not g55250 (n_24732, n33525);
  and g55251 (n33527, n_24732, n33526);
  not g55252 (n_24733, n33511);
  not g55253 (n_24734, n33527);
  and g55254 (n33528, n_24733, n_24734);
  not g55255 (n_24735, n33528);
  and g55256 (n33529, n_161, n_24735);
  not g55257 (n_24736, n33428);
  and g55258 (n33530, n2571, n_24736);
  not g55259 (n_24737, n33529);
  and g55260 (n33531, n_24737, n33530);
  not g55261 (n_24738, n33420);
  not g55262 (n_24739, n33531);
  and g55263 (n33532, n_24738, n_24739);
  not g55264 (n_24740, n33532);
  and g55265 (n33533, n_11749, n_24740);
  and g55266 (n33534, n_11753, n33417);
  and g55267 (n33535, pi0625, n33532);
  not g55268 (n_24741, n33534);
  and g55269 (n33536, pi1153, n_24741);
  not g55270 (n_24742, n33535);
  and g55271 (n33537, n_24742, n33536);
  and g55272 (n33538, n_11753, n33532);
  and g55273 (n33539, pi0625, n33417);
  not g55274 (n_24743, n33539);
  and g55275 (n33540, n_11757, n_24743);
  not g55276 (n_24744, n33538);
  and g55277 (n33541, n_24744, n33540);
  not g55278 (n_24745, n33537);
  not g55279 (n_24746, n33541);
  and g55280 (n33542, n_24745, n_24746);
  not g55281 (n_24747, n33542);
  and g55282 (n33543, pi0778, n_24747);
  not g55283 (n_24748, n33533);
  not g55284 (n_24749, n33543);
  and g55285 (n33544, n_24748, n_24749);
  and g55286 (n33545, n_11773, n33544);
  and g55287 (n33546, n17075, n33417);
  not g55288 (n_24750, n33545);
  not g55289 (n_24751, n33546);
  and g55290 (n33547, n_24750, n_24751);
  and g55291 (n33548, n_11777, n33547);
  not g55292 (n_24752, n33419);
  not g55293 (n_24753, n33548);
  and g55294 (n33549, n_24752, n_24753);
  and g55295 (n33550, n_11780, n33549);
  and g55296 (n33551, n_11783, n33550);
  not g55297 (n_24754, n33418);
  not g55298 (n_24755, n33551);
  and g55299 (n33552, n_24754, n_24755);
  and g55300 (n33553, n_11787, n33552);
  not g55301 (n_24756, n33552);
  and g55302 (n33554, pi0628, n_24756);
  and g55303 (n33555, n_11789, n33417);
  not g55304 (n_24757, n33554);
  not g55305 (n_24758, n33555);
  and g55306 (n33556, n_24757, n_24758);
  and g55307 (n33557, pi1156, n33556);
  and g55308 (n33558, pi0628, n33417);
  and g55309 (n33559, n_11789, n_24756);
  not g55310 (n_24759, n33558);
  and g55311 (n33560, n_11794, n_24759);
  not g55312 (n_24760, n33559);
  and g55313 (n33561, n_24760, n33560);
  not g55314 (n_24761, n33557);
  not g55315 (n_24762, n33561);
  and g55316 (n33562, n_24761, n_24762);
  not g55317 (n_24763, n33562);
  and g55318 (n33563, pi0792, n_24763);
  not g55319 (n_24764, n33553);
  not g55320 (n_24765, n33563);
  and g55321 (n33564, n_24764, n_24765);
  and g55322 (n33565, n_11806, n33564);
  and g55323 (n33566, pi0647, n33417);
  not g55324 (n_24766, n33566);
  and g55325 (n33567, n_11810, n_24766);
  not g55326 (n_24767, n33565);
  and g55327 (n33568, n_24767, n33567);
  and g55328 (n33569, pi0630, n33568);
  and g55329 (n33570, n17779, n_24652);
  and g55330 (n33571, n_11836, n_11839);
  not g55331 (n_24769, n33571);
  and g55332 (n33572, pi0633, n_24769);
  not g55333 (n_24770, n33572);
  and g55334 (n33573, n_11643, n_24770);
  not g55335 (n_24771, n33573);
  and g55336 (n33574, n_11843, n_24771);
  and g55337 (n33575, n_234, n33574);
  and g55338 (n33576, pi0603, pi0633);
  not g55339 (n_24772, n33522);
  not g55340 (n_24773, n33576);
  and g55341 (n33577, n_24772, n_24773);
  and g55342 (n33578, pi0198, n_11832);
  and g55343 (n33579, n_305, n17230);
  not g55344 (n_24774, n33578);
  not g55345 (n_24775, n33579);
  and g55346 (n33580, n_24774, n_24775);
  and g55347 (n33581, n33576, n33580);
  not g55348 (n_24776, n33577);
  not g55349 (n_24777, n33581);
  and g55350 (n33582, n_24776, n_24777);
  and g55351 (n33583, pi0299, n33582);
  not g55352 (n_24778, n33575);
  and g55353 (n33584, n_162, n_24778);
  not g55354 (n_24779, n33583);
  and g55355 (n33585, n_24779, n33584);
  and g55356 (n33586, pi0633, n17239);
  not g55357 (n_24780, n33385);
  not g55358 (n_24781, n33586);
  and g55359 (n33587, n_24780, n_24781);
  not g55360 (n_24782, n33587);
  and g55361 (n33588, n_3139, n_24782);
  and g55362 (n33589, pi0633, n16653);
  and g55363 (n33590, n_11865, n33589);
  and g55364 (n33591, n_11479, n33590);
  not g55365 (n_24783, n33591);
  and g55366 (n33592, n_24659, n_24783);
  not g55367 (n_24784, n33592);
  and g55368 (n33593, n17188, n_24784);
  not g55369 (n_24785, n33588);
  not g55370 (n_24786, n33593);
  and g55371 (n33594, n_24785, n_24786);
  and g55372 (n33595, n_3119, n33594);
  not g55373 (n_24787, n33590);
  and g55374 (n33596, n_24623, n_24787);
  not g55375 (n_24788, n33596);
  and g55376 (n33597, pi0603, n_24788);
  and g55377 (n33598, n_11512, n33379);
  not g55378 (n_24789, n33597);
  not g55379 (n_24790, n33598);
  and g55380 (n33599, n_24789, n_24790);
  and g55381 (n33600, n_11867, n33599);
  and g55382 (n33601, n6197, n_24788);
  not g55383 (n_24791, n33378);
  and g55384 (n33602, n_24791, n_24783);
  not g55385 (n_24792, n33601);
  and g55386 (n33603, n_24792, n33602);
  not g55387 (n_24793, n33603);
  and g55388 (n33604, pi0603, n_24793);
  and g55389 (n33605, n17167, n_24790);
  not g55390 (n_24794, n33604);
  and g55391 (n33606, n_24794, n33605);
  not g55392 (n_24795, n33600);
  not g55393 (n_24796, n33606);
  and g55394 (n33607, n_24795, n_24796);
  and g55395 (n33608, n_3139, n33607);
  and g55396 (n33609, n_24791, n_24794);
  not g55397 (n_24797, n33609);
  and g55398 (n33610, n6195, n_24797);
  not g55399 (n_24798, n33608);
  not g55400 (n_24799, n33610);
  and g55401 (n33611, n_24798, n_24799);
  and g55402 (n33612, n6205, n33611);
  not g55403 (n_24800, n33595);
  and g55404 (n33613, pi0223, n_24800);
  not g55405 (n_24801, n33612);
  and g55406 (n33614, n_24801, n33613);
  and g55407 (n33615, n2603, n33599);
  and g55408 (n33616, pi0642, n_24789);
  and g55409 (n33617, pi0633, n17147);
  not g55410 (n_24802, n33617);
  and g55411 (n33618, n_24684, n_24802);
  not g55412 (n_24803, n33618);
  and g55413 (n33619, n_3102, n_24803);
  not g55414 (n_24804, n33619);
  and g55415 (n33620, n_24792, n_24804);
  not g55416 (n_24805, n33620);
  and g55417 (n33621, pi0603, n_24805);
  not g55418 (n_24806, n33621);
  and g55419 (n33622, n_3087, n_24806);
  not g55420 (n_24807, n33616);
  and g55421 (n33623, n6191, n_24807);
  not g55422 (n_24808, n33622);
  and g55423 (n33624, n_24808, n33623);
  not g55424 (n_24809, n6191);
  and g55425 (n33625, n_24809, n33597);
  not g55426 (n_24810, n33625);
  and g55427 (n33626, n_24790, n_24810);
  not g55428 (n_24811, n33624);
  and g55429 (n33627, n_24811, n33626);
  and g55430 (n33628, n_3139, n33627);
  and g55431 (n33629, n_11512, n33390);
  not g55432 (n_24812, n33629);
  and g55433 (n33630, n6195, n_24812);
  and g55434 (n33631, n_24806, n33630);
  not g55435 (n_24813, n33628);
  not g55436 (n_24814, n33631);
  and g55437 (n33632, n_24813, n_24814);
  and g55438 (n33633, n6205, n33632);
  and g55439 (n33634, pi0603, n_24803);
  and g55440 (n33635, n17167, n33634);
  and g55441 (n33636, pi0198, n17149);
  and g55442 (n33637, n6197, n33618);
  and g55443 (n33638, n_3102, n33596);
  and g55444 (n33639, pi0603, n_11867);
  not g55445 (n_24815, n33638);
  and g55446 (n33640, n_24815, n33639);
  not g55447 (n_24816, n33637);
  and g55448 (n33641, n_24816, n33640);
  not g55449 (n_24817, n33635);
  not g55450 (n_24818, n33636);
  and g55451 (n33642, n_24817, n_24818);
  not g55452 (n_24819, n33641);
  and g55453 (n33643, n_24819, n33642);
  and g55454 (n33644, n_3139, n33643);
  and g55455 (n33645, n6195, n_24684);
  not g55456 (n_24820, n33634);
  and g55457 (n33646, n_24820, n33645);
  not g55458 (n_24821, n33644);
  not g55459 (n_24822, n33646);
  and g55460 (n33647, n_24821, n_24822);
  and g55461 (n33648, n_3119, n33647);
  not g55462 (n_24823, n33648);
  and g55463 (n33649, n_9349, n_24823);
  not g55464 (n_24824, n33633);
  and g55465 (n33650, n_24824, n33649);
  not g55466 (n_24825, n33615);
  and g55467 (n33651, n_223, n_24825);
  not g55468 (n_24826, n33650);
  and g55469 (n33652, n_24826, n33651);
  not g55470 (n_24827, n33614);
  not g55471 (n_24828, n33652);
  and g55472 (n33653, n_24827, n_24828);
  not g55473 (n_24829, n33653);
  and g55474 (n33654, n_234, n_24829);
  and g55475 (n33655, n_3162, n33594);
  and g55476 (n33656, n6242, n33611);
  not g55477 (n_24830, n33655);
  and g55478 (n33657, pi0215, n_24830);
  not g55479 (n_24831, n33656);
  and g55480 (n33658, n_24831, n33657);
  and g55481 (n33659, n3448, n33599);
  and g55482 (n33660, n_3162, n33647);
  and g55483 (n33661, n6242, n33632);
  not g55484 (n_24832, n33660);
  and g55485 (n33662, n_9350, n_24832);
  not g55486 (n_24833, n33661);
  and g55487 (n33663, n_24833, n33662);
  not g55488 (n_24834, n33659);
  and g55489 (n33664, n_36, n_24834);
  not g55490 (n_24835, n33663);
  and g55491 (n33665, n_24835, n33664);
  not g55492 (n_24836, n33658);
  not g55493 (n_24837, n33665);
  and g55494 (n33666, n_24836, n_24837);
  not g55495 (n_24838, n33666);
  and g55496 (n33667, pi0299, n_24838);
  not g55497 (n_24839, n33654);
  and g55498 (n33668, pi0039, n_24839);
  not g55499 (n_24840, n33667);
  and g55500 (n33669, n_24840, n33668);
  not g55501 (n_24841, n33585);
  not g55502 (n_24842, n33669);
  and g55503 (n33670, n_24841, n_24842);
  not g55504 (n_24843, n33670);
  and g55505 (n33671, n_161, n_24843);
  and g55506 (n33672, pi0633, n17168);
  and g55507 (n33673, n16667, n33672);
  not g55508 (n_24844, n33673);
  and g55509 (n33674, n_24655, n_24844);
  not g55510 (n_24845, n33674);
  and g55511 (n33675, n_162, n_24845);
  not g55512 (n_24846, n33675);
  and g55513 (n33676, n33422, n_24846);
  not g55514 (n_24847, n33676);
  and g55515 (n33677, n2571, n_24847);
  not g55516 (n_24848, n33671);
  and g55517 (n33678, n_24848, n33677);
  not g55518 (n_24849, n33678);
  and g55519 (n33679, n_24738, n_24849);
  not g55520 (n_24850, n33679);
  and g55521 (n33680, n_11960, n_24850);
  and g55522 (n33681, n17117, n_24652);
  not g55523 (n_24851, n33680);
  not g55524 (n_24852, n33681);
  and g55525 (n33682, n_24851, n_24852);
  not g55526 (n_24853, n33682);
  and g55527 (n33683, n_11964, n_24853);
  and g55528 (n33684, n_11967, n_24652);
  and g55529 (n33685, pi0609, n33680);
  not g55530 (n_24854, n33684);
  not g55531 (n_24855, n33685);
  and g55532 (n33686, n_24854, n_24855);
  not g55533 (n_24856, n33686);
  and g55534 (n33687, pi1155, n_24856);
  and g55535 (n33688, n_11972, n_24652);
  and g55536 (n33689, n_11971, n33680);
  not g55537 (n_24857, n33688);
  not g55538 (n_24858, n33689);
  and g55539 (n33690, n_24857, n_24858);
  not g55540 (n_24859, n33690);
  and g55541 (n33691, n_11768, n_24859);
  not g55542 (n_24860, n33687);
  not g55543 (n_24861, n33691);
  and g55544 (n33692, n_24860, n_24861);
  not g55545 (n_24862, n33692);
  and g55546 (n33693, pi0785, n_24862);
  not g55547 (n_24863, n33683);
  not g55548 (n_24864, n33693);
  and g55549 (n33694, n_24863, n_24864);
  not g55550 (n_24865, n33694);
  and g55551 (n33695, n_11981, n_24865);
  and g55552 (n33696, n_11984, n33417);
  and g55553 (n33697, pi0618, n33694);
  not g55554 (n_24866, n33696);
  and g55555 (n33698, pi1154, n_24866);
  not g55556 (n_24867, n33697);
  and g55557 (n33699, n_24867, n33698);
  and g55558 (n33700, n_11984, n33694);
  and g55559 (n33701, pi0618, n33417);
  not g55560 (n_24868, n33701);
  and g55561 (n33702, n_11413, n_24868);
  not g55562 (n_24869, n33700);
  and g55563 (n33703, n_24869, n33702);
  not g55564 (n_24870, n33699);
  not g55565 (n_24871, n33703);
  and g55566 (n33704, n_24870, n_24871);
  not g55567 (n_24872, n33704);
  and g55568 (n33705, pi0781, n_24872);
  not g55569 (n_24873, n33695);
  not g55570 (n_24874, n33705);
  and g55571 (n33706, n_24873, n_24874);
  not g55572 (n_24875, n33706);
  and g55573 (n33707, n_12315, n_24875);
  and g55574 (n33708, n_11821, n33417);
  and g55575 (n33709, pi0619, n33706);
  not g55576 (n_24876, n33708);
  and g55577 (n33710, pi1159, n_24876);
  not g55578 (n_24877, n33709);
  and g55579 (n33711, n_24877, n33710);
  and g55580 (n33712, n_11821, n33706);
  and g55581 (n33713, pi0619, n33417);
  not g55582 (n_24878, n33713);
  and g55583 (n33714, n_11405, n_24878);
  not g55584 (n_24879, n33712);
  and g55585 (n33715, n_24879, n33714);
  not g55586 (n_24880, n33711);
  not g55587 (n_24881, n33715);
  and g55588 (n33716, n_24880, n_24881);
  not g55589 (n_24882, n33716);
  and g55590 (n33717, pi0789, n_24882);
  not g55591 (n_24883, n33707);
  not g55592 (n_24884, n33717);
  and g55593 (n33718, n_24883, n_24884);
  and g55594 (n33719, n_12524, n33718);
  and g55595 (n33720, n17969, n33417);
  not g55596 (n_24885, n33719);
  not g55597 (n_24886, n33720);
  and g55598 (n33721, n_24885, n_24886);
  and g55599 (n33722, n_12368, n33721);
  not g55600 (n_24887, n33570);
  not g55601 (n_24888, n33722);
  and g55602 (n33723, n_24887, n_24888);
  not g55603 (n_24889, n33723);
  and g55604 (n33724, n_14548, n_24889);
  not g55605 (n_24890, n33564);
  and g55606 (n33725, pi0647, n_24890);
  and g55607 (n33726, n_11806, n_24652);
  not g55608 (n_24891, n33725);
  not g55609 (n_24892, n33726);
  and g55610 (n33727, n_24891, n_24892);
  not g55611 (n_24893, n33727);
  and g55612 (n33728, n17801, n_24893);
  not g55613 (n_24894, n33569);
  not g55614 (n_24895, n33728);
  and g55615 (n33729, n_24894, n_24895);
  not g55616 (n_24896, n33724);
  and g55617 (n33730, n_24896, n33729);
  not g55618 (n_24897, n33730);
  and g55619 (n33731, pi0787, n_24897);
  and g55620 (n33732, pi0629, n33561);
  and g55621 (n33733, n_14557, n33721);
  and g55622 (n33734, n17776, n33556);
  not g55623 (n_24898, n33732);
  not g55624 (n_24899, n33734);
  and g55625 (n33735, n_24898, n_24899);
  not g55626 (n_24900, n33733);
  and g55627 (n33736, n_24900, n33735);
  not g55628 (n_24901, n33736);
  and g55629 (n33737, pi0792, n_24901);
  and g55630 (n33738, n16635, n33417);
  not g55631 (n_24902, n33550);
  not g55632 (n_24903, n33738);
  and g55633 (n33739, n_24902, n_24903);
  not g55634 (n_24904, n33739);
  and g55635 (n33740, n17871, n_24904);
  not g55636 (n_24905, n33718);
  and g55637 (n33741, n_12320, n_24905);
  and g55638 (n33742, pi0626, n_24652);
  not g55639 (n_24906, n33742);
  and g55640 (n33743, n16629, n_24906);
  not g55641 (n_24907, n33741);
  and g55642 (n33744, n_24907, n33743);
  and g55643 (n33745, pi0626, n_24905);
  and g55644 (n33746, n_12320, n_24652);
  not g55645 (n_24908, n33746);
  and g55646 (n33747, n16628, n_24908);
  not g55647 (n_24909, n33745);
  and g55648 (n33748, n_24909, n33747);
  not g55649 (n_24910, n33740);
  not g55650 (n_24911, n33744);
  and g55651 (n33749, n_24910, n_24911);
  not g55652 (n_24912, n33748);
  and g55653 (n33750, n_24912, n33749);
  not g55654 (n_24913, n33750);
  and g55655 (n33751, pi0788, n_24913);
  and g55656 (n33752, pi0609, n33544);
  and g55657 (n33753, pi0634, n17645);
  not g55658 (n_24914, n33753);
  and g55659 (n33754, n33674, n_24914);
  not g55660 (n_24915, n33754);
  and g55661 (n33755, n_162, n_24915);
  not g55662 (n_24916, n33755);
  and g55663 (n33756, n33422, n_24916);
  and g55664 (n33757, n_24727, n33582);
  and g55665 (n33758, n_11512, n_24726);
  and g55666 (n33759, n_305, n_12032);
  and g55667 (n33760, n17122, n33759);
  not g55668 (n_24917, n17230);
  and g55669 (n33761, n_24917, n33519);
  not g55670 (n_24918, pi0633);
  not g55671 (n_24919, n33760);
  and g55672 (n33762, n_24918, n_24919);
  not g55673 (n_24920, n33761);
  and g55674 (n33763, n_24920, n33762);
  and g55675 (n33764, pi0198, n_12032);
  not g55680 (n_24922, n33763);
  and g55681 (n33768, pi0603, n_24922);
  not g55682 (n_24923, n33767);
  and g55683 (n33769, n_24923, n33768);
  not g55684 (n_24924, n33758);
  not g55685 (n_24925, n33769);
  and g55686 (n33770, n_24924, n_24925);
  not g55687 (n_24926, n33770);
  and g55688 (n33771, n33512, n_24926);
  not g55689 (n_24927, n33757);
  and g55690 (n33772, pi0299, n_24927);
  not g55691 (n_24928, n33771);
  and g55692 (n33773, n_24928, n33772);
  and g55693 (n33774, n_11502, n33574);
  and g55694 (n33775, n_11512, n33516);
  and g55695 (n33776, pi0198, n_24918);
  and g55696 (n33777, pi0634, n_12032);
  not g55697 (n_24929, n33776);
  and g55698 (n33778, n_24929, n33777);
  and g55699 (n33779, n_11835, n33778);
  not g55700 (n_24930, pi0634);
  and g55701 (n33780, n_24930, n16929);
  and g55702 (n33781, pi0634, n16932);
  and g55703 (n33782, n_11917, n33781);
  not g55704 (n_24931, n33780);
  not g55705 (n_24932, n33782);
  and g55706 (n33783, n_24931, n_24932);
  not g55707 (n_24933, n33783);
  and g55708 (n33784, n_24918, n_24933);
  not g55714 (n_24936, n33775);
  and g55715 (n33788, pi0680, n_24936);
  not g55716 (n_24937, n33787);
  and g55717 (n33789, n_24937, n33788);
  not g55718 (n_24938, n33774);
  and g55719 (n33790, n_234, n_24938);
  not g55720 (n_24939, n33789);
  and g55721 (n33791, n_24939, n33790);
  not g55722 (n_24940, n33773);
  not g55723 (n_24941, n33791);
  and g55724 (n33792, n_24940, n_24941);
  not g55725 (n_24942, n33792);
  and g55726 (n33793, n_162, n_24942);
  and g55727 (n33794, n17355, n33437);
  not g55728 (n_24943, n33794);
  and g55729 (n33795, n33599, n_24943);
  and g55730 (n33796, n2603, n33795);
  and g55731 (n33797, n_11502, n33627);
  and g55732 (n33798, n_11512, n_24672);
  and g55733 (n33799, n17159, n33777);
  not g55734 (n_24944, n33799);
  and g55735 (n33800, n33596, n_24944);
  not g55736 (n_24945, n33800);
  and g55737 (n33801, pi0603, n_24945);
  not g55738 (n_24946, n33798);
  not g55739 (n_24947, n33801);
  and g55740 (n33802, n_24946, n_24947);
  not g55741 (n_24948, n33802);
  and g55742 (n33803, n_24809, n_24948);
  and g55743 (n33804, n6197, n_24945);
  and g55744 (n33805, pi0634, n17424);
  not g55745 (n_24949, n33805);
  and g55746 (n33806, n33618, n_24949);
  not g55747 (n_24950, n33806);
  and g55748 (n33807, n_3102, n_24950);
  not g55749 (n_24951, n33804);
  not g55750 (n_24952, n33807);
  and g55751 (n33808, n_24951, n_24952);
  not g55752 (n_24953, n33808);
  and g55753 (n33809, pi0603, n_24953);
  and g55754 (n33810, n_3087, n33809);
  and g55755 (n33811, pi0642, n33801);
  not g55756 (n_24954, n33811);
  and g55757 (n33812, n_24946, n_24954);
  not g55758 (n_24955, n33810);
  and g55759 (n33813, n_24955, n33812);
  not g55760 (n_24956, n33813);
  and g55761 (n33814, n6191, n_24956);
  not g55762 (n_24957, n33803);
  and g55763 (n33815, n_11455, n_24957);
  not g55764 (n_24958, n33814);
  and g55765 (n33816, n_24958, n33815);
  and g55766 (n33817, n_11512, n_24688);
  not g55767 (n_24959, n33817);
  and g55768 (n33818, n16657, n_24959);
  not g55769 (n_24960, n33809);
  and g55770 (n33819, n_24960, n33818);
  not g55771 (n_24961, n33816);
  not g55772 (n_24962, n33819);
  and g55773 (n33820, n_24961, n_24962);
  not g55774 (n_24963, n33820);
  and g55775 (n33821, pi0680, n_24963);
  not g55776 (n_24964, n33797);
  not g55777 (n_24965, n33821);
  and g55778 (n33822, n_24964, n_24965);
  and g55779 (n33823, n6205, n33822);
  not g55780 (n_24966, n33643);
  and g55781 (n33824, n_11502, n_24966);
  and g55782 (n33825, n_11512, n33484);
  and g55783 (n33826, n_11867, n33801);
  not g55784 (n_24967, n33640);
  not g55785 (n_24968, n33826);
  and g55786 (n33827, n_24967, n_24968);
  and g55787 (n33828, n_3138, n33827);
  not g55788 (n_24969, n33827);
  and g55789 (n33829, n_3102, n_24969);
  not g55790 (n_24970, n33829);
  and g55791 (n33830, n33806, n_24970);
  not g55792 (n_24971, n33828);
  not g55793 (n_24972, n33830);
  and g55794 (n33831, n_24971, n_24972);
  not g55795 (n_24973, n33825);
  not g55796 (n_24974, n33831);
  and g55797 (n33832, n_24973, n_24974);
  not g55798 (n_24975, n33832);
  and g55799 (n33833, n17323, n_24975);
  and g55800 (n33834, n_11866, n_24686);
  not g55801 (n_24976, n33834);
  and g55802 (n33835, n_24820, n_24976);
  not g55803 (n_24977, n33835);
  and g55804 (n33836, n6195, n_24977);
  not g55805 (n_24978, n33824);
  not g55806 (n_24979, n33836);
  and g55807 (n33837, n_24978, n_24979);
  not g55808 (n_24980, n33833);
  and g55809 (n33838, n_24980, n33837);
  not g55810 (n_24981, n33838);
  and g55811 (n33839, n_3119, n_24981);
  not g55812 (n_24982, n33839);
  and g55813 (n33840, n_9349, n_24982);
  not g55814 (n_24983, n33823);
  and g55815 (n33841, n_24983, n33840);
  not g55816 (n_24984, n33796);
  and g55817 (n33842, n_223, n_24984);
  not g55818 (n_24985, n33841);
  and g55819 (n33843, n_24985, n33842);
  and g55820 (n33844, n_11502, n_24782);
  and g55821 (n33845, n17191, n33759);
  and g55822 (n33846, n17144, n33764);
  not g55823 (n_24986, n33846);
  and g55824 (n33847, n_24659, n_24986);
  not g55825 (n_24987, n33845);
  and g55826 (n33848, n_24987, n33847);
  not g55827 (n_24988, n33848);
  and g55828 (n33849, pi0634, n_24988);
  and g55829 (n33850, n_24930, n33429);
  not g55830 (n_24989, n33850);
  and g55831 (n33851, n_24783, n_24989);
  not g55832 (n_24990, n33849);
  and g55833 (n33852, n_24990, n33851);
  not g55834 (n_24991, n33852);
  and g55835 (n33853, pi0603, n_24991);
  and g55836 (n33854, n_11512, n_24661);
  not g55837 (n_24992, n33853);
  not g55838 (n_24993, n33854);
  and g55839 (n33855, n_24992, n_24993);
  not g55840 (n_24994, n33855);
  and g55841 (n33856, n6195, n_24994);
  and g55842 (n33857, n17167, n33853);
  and g55843 (n33858, n_11512, n33441);
  and g55844 (n33859, n_24969, n_24991);
  not g55851 (n_24998, n33862);
  and g55852 (n33863, n17323, n_24998);
  not g55853 (n_24999, n33844);
  not g55854 (n_25000, n33856);
  and g55855 (n33864, n_24999, n_25000);
  not g55856 (n_25001, n33863);
  and g55857 (n33865, n_25001, n33864);
  and g55858 (n33866, n_3119, n33865);
  and g55859 (n33867, n_11502, n33607);
  and g55860 (n33868, n_3102, n_24991);
  not g55861 (n_25002, n33868);
  and g55862 (n33869, n_24951, n_25002);
  not g55863 (n_25003, n33869);
  and g55864 (n33870, pi0603, n_25003);
  and g55865 (n33871, n_11512, n_24677);
  not g55866 (n_25004, n33870);
  not g55867 (n_25005, n33871);
  and g55868 (n33872, n_25004, n_25005);
  not g55869 (n_25006, n33872);
  and g55870 (n33873, n6195, n_25006);
  and g55871 (n33874, n_11867, n33802);
  and g55872 (n33875, n17167, n_24946);
  and g55873 (n33876, n_25004, n33875);
  not g55874 (n_25007, n33874);
  and g55875 (n33877, n17323, n_25007);
  not g55876 (n_25008, n33876);
  and g55877 (n33878, n_25008, n33877);
  not g55878 (n_25009, n33867);
  not g55879 (n_25010, n33873);
  and g55880 (n33879, n_25009, n_25010);
  not g55881 (n_25011, n33878);
  and g55882 (n33880, n_25011, n33879);
  and g55883 (n33881, n6205, n33880);
  not g55884 (n_25012, n33866);
  and g55885 (n33882, pi0223, n_25012);
  not g55886 (n_25013, n33881);
  and g55887 (n33883, n_25013, n33882);
  not g55888 (n_25014, n33843);
  not g55889 (n_25015, n33883);
  and g55890 (n33884, n_25014, n_25015);
  not g55891 (n_25016, n33884);
  and g55892 (n33885, n_234, n_25016);
  and g55893 (n33886, n3448, n33795);
  and g55894 (n33887, n6242, n33822);
  and g55895 (n33888, n_3162, n_24981);
  not g55896 (n_25017, n33888);
  and g55897 (n33889, n_9350, n_25017);
  not g55898 (n_25018, n33887);
  and g55899 (n33890, n_25018, n33889);
  not g55900 (n_25019, n33886);
  and g55901 (n33891, n_36, n_25019);
  not g55902 (n_25020, n33890);
  and g55903 (n33892, n_25020, n33891);
  and g55904 (n33893, n_3162, n33865);
  and g55905 (n33894, n6242, n33880);
  not g55906 (n_25021, n33893);
  and g55907 (n33895, pi0215, n_25021);
  not g55908 (n_25022, n33894);
  and g55909 (n33896, n_25022, n33895);
  not g55910 (n_25023, n33892);
  not g55911 (n_25024, n33896);
  and g55912 (n33897, n_25023, n_25024);
  not g55913 (n_25025, n33897);
  and g55914 (n33898, pi0299, n_25025);
  not g55915 (n_25026, n33885);
  and g55916 (n33899, pi0039, n_25026);
  not g55917 (n_25027, n33898);
  and g55918 (n33900, n_25027, n33899);
  not g55919 (n_25028, n33793);
  not g55920 (n_25029, n33900);
  and g55921 (n33901, n_25028, n_25029);
  not g55922 (n_25030, n33901);
  and g55923 (n33902, n_161, n_25030);
  not g55924 (n_25031, n33756);
  and g55925 (n33903, n2571, n_25031);
  not g55926 (n_25032, n33902);
  and g55927 (n33904, n_25032, n33903);
  not g55928 (n_25033, n33904);
  and g55929 (n33905, n_24738, n_25033);
  and g55930 (n33906, n_11753, n33905);
  and g55931 (n33907, pi0625, n33679);
  not g55932 (n_25034, n33907);
  and g55933 (n33908, n_11757, n_25034);
  not g55934 (n_25035, n33906);
  and g55935 (n33909, n_25035, n33908);
  and g55936 (n33910, n_11823, n_24745);
  not g55937 (n_25036, n33909);
  and g55938 (n33911, n_25036, n33910);
  and g55939 (n33912, n_11753, n33679);
  and g55940 (n33913, pi0625, n33905);
  not g55941 (n_25037, n33912);
  and g55942 (n33914, pi1153, n_25037);
  not g55943 (n_25038, n33913);
  and g55944 (n33915, n_25038, n33914);
  and g55945 (n33916, pi0608, n_24746);
  not g55946 (n_25039, n33915);
  and g55947 (n33917, n_25039, n33916);
  not g55948 (n_25040, n33911);
  not g55949 (n_25041, n33917);
  and g55950 (n33918, n_25040, n_25041);
  not g55951 (n_25042, n33918);
  and g55952 (n33919, pi0778, n_25042);
  and g55953 (n33920, n_11749, n33905);
  not g55954 (n_25043, n33919);
  not g55955 (n_25044, n33920);
  and g55956 (n33921, n_25043, n_25044);
  not g55957 (n_25045, n33921);
  and g55958 (n33922, n_11971, n_25045);
  not g55959 (n_25046, n33752);
  and g55960 (n33923, n_11768, n_25046);
  not g55961 (n_25047, n33922);
  and g55962 (n33924, n_25047, n33923);
  and g55963 (n33925, n_11767, n_24860);
  not g55964 (n_25048, n33924);
  and g55965 (n33926, n_25048, n33925);
  and g55966 (n33927, n_11971, n33544);
  and g55967 (n33928, pi0609, n_25045);
  not g55968 (n_25049, n33927);
  and g55969 (n33929, pi1155, n_25049);
  not g55970 (n_25050, n33928);
  and g55971 (n33930, n_25050, n33929);
  and g55972 (n33931, pi0660, n_24861);
  not g55973 (n_25051, n33930);
  and g55974 (n33932, n_25051, n33931);
  not g55975 (n_25052, n33926);
  not g55976 (n_25053, n33932);
  and g55977 (n33933, n_25052, n_25053);
  not g55978 (n_25054, n33933);
  and g55979 (n33934, pi0785, n_25054);
  and g55980 (n33935, n_11964, n_25045);
  not g55981 (n_25055, n33934);
  not g55982 (n_25056, n33935);
  and g55983 (n33936, n_25055, n_25056);
  not g55984 (n_25057, n33936);
  and g55985 (n33937, n_11984, n_25057);
  not g55986 (n_25058, n33547);
  and g55987 (n33938, pi0618, n_25058);
  not g55988 (n_25059, n33938);
  and g55989 (n33939, n_11413, n_25059);
  not g55990 (n_25060, n33937);
  and g55991 (n33940, n_25060, n33939);
  and g55992 (n33941, n_11412, n_24870);
  not g55993 (n_25061, n33940);
  and g55994 (n33942, n_25061, n33941);
  and g55995 (n33943, pi0618, n_25057);
  and g55996 (n33944, n_11984, n_25058);
  not g55997 (n_25062, n33944);
  and g55998 (n33945, pi1154, n_25062);
  not g55999 (n_25063, n33943);
  and g56000 (n33946, n_25063, n33945);
  and g56001 (n33947, pi0627, n_24871);
  not g56002 (n_25064, n33946);
  and g56003 (n33948, n_25064, n33947);
  not g56004 (n_25065, n33942);
  not g56005 (n_25066, n33948);
  and g56006 (n33949, n_25065, n_25066);
  not g56007 (n_25067, n33949);
  and g56008 (n33950, pi0781, n_25067);
  and g56009 (n33951, n_11981, n_25057);
  not g56010 (n_25068, n33950);
  not g56011 (n_25069, n33951);
  and g56012 (n33952, n_25068, n_25069);
  and g56013 (n33953, n_12315, n33952);
  not g56014 (n_25070, n33952);
  and g56015 (n33954, n_11821, n_25070);
  and g56016 (n33955, pi0619, n33549);
  not g56017 (n_25071, n33955);
  and g56018 (n33956, n_11405, n_25071);
  not g56019 (n_25072, n33954);
  and g56020 (n33957, n_25072, n33956);
  and g56021 (n33958, n_11403, n_24880);
  not g56022 (n_25073, n33957);
  and g56023 (n33959, n_25073, n33958);
  and g56024 (n33960, n_11821, n33549);
  and g56025 (n33961, pi0619, n_25070);
  not g56026 (n_25074, n33960);
  and g56027 (n33962, pi1159, n_25074);
  not g56028 (n_25075, n33961);
  and g56029 (n33963, n_25075, n33962);
  and g56030 (n33964, pi0648, n_24881);
  not g56031 (n_25076, n33963);
  and g56032 (n33965, n_25076, n33964);
  not g56033 (n_25077, n33959);
  and g56034 (n33966, pi0789, n_25077);
  not g56035 (n_25078, n33965);
  and g56036 (n33967, n_25078, n33966);
  not g56037 (n_25079, n33953);
  and g56038 (n33968, n17970, n_25079);
  not g56039 (n_25080, n33967);
  and g56040 (n33969, n_25080, n33968);
  not g56041 (n_25081, n33751);
  not g56042 (n_25082, n33969);
  and g56043 (n33970, n_25081, n_25082);
  not g56044 (n_25083, n33737);
  not g56045 (n_25084, n33970);
  and g56046 (n33971, n_25083, n_25084);
  and g56047 (n33972, n20364, n33736);
  not g56048 (n_25085, n33972);
  and g56049 (n33973, n_14387, n_25085);
  not g56050 (n_25086, n33971);
  and g56051 (n33974, n_25086, n33973);
  not g56052 (n_25087, n33731);
  not g56053 (n_25088, n33974);
  and g56054 (n33975, n_25087, n_25088);
  not g56055 (n_25089, n33975);
  and g56056 (n33976, n_12411, n_25089);
  and g56057 (n33977, n_11803, n_24890);
  and g56058 (n33978, pi1157, n_24893);
  not g56059 (n_25090, n33568);
  not g56060 (n_25091, n33978);
  and g56061 (n33979, n_25090, n_25091);
  not g56062 (n_25092, n33979);
  and g56063 (n33980, pi0787, n_25092);
  not g56064 (n_25093, n33977);
  not g56065 (n_25094, n33980);
  and g56066 (n33981, n_25093, n_25094);
  and g56067 (n33982, n_11819, n33981);
  and g56068 (n33983, pi0644, n33975);
  not g56069 (n_25095, n33982);
  and g56070 (n33984, pi0715, n_25095);
  not g56071 (n_25096, n33983);
  and g56072 (n33985, n_25096, n33984);
  and g56073 (n33986, n_12392, n33723);
  and g56074 (n33987, n17804, n33417);
  not g56075 (n_25097, n33986);
  not g56076 (n_25098, n33987);
  and g56077 (n33988, n_25097, n_25098);
  not g56078 (n_25099, n33988);
  and g56079 (n33989, pi0644, n_25099);
  and g56080 (n33990, n_11819, n33417);
  not g56081 (n_25100, n33990);
  and g56082 (n33991, n_12395, n_25100);
  not g56083 (n_25101, n33989);
  and g56084 (n33992, n_25101, n33991);
  not g56085 (n_25102, n33992);
  and g56086 (n33993, pi1160, n_25102);
  not g56087 (n_25103, n33985);
  and g56088 (n33994, n_25103, n33993);
  and g56089 (n33995, n_11819, n_25099);
  and g56090 (n33996, pi0644, n33417);
  not g56091 (n_25104, n33996);
  and g56092 (n33997, pi0715, n_25104);
  not g56093 (n_25105, n33995);
  and g56094 (n33998, n_25105, n33997);
  and g56095 (n33999, pi0644, n33981);
  and g56096 (n34000, n_11819, n33975);
  not g56097 (n_25106, n33999);
  and g56098 (n34001, n_12395, n_25106);
  not g56099 (n_25107, n34000);
  and g56100 (n34002, n_25107, n34001);
  not g56101 (n_25108, n33998);
  and g56102 (n34003, n_12405, n_25108);
  not g56103 (n_25109, n34002);
  and g56104 (n34004, n_25109, n34003);
  not g56105 (n_25110, n33994);
  and g56106 (n34005, pi0790, n_25110);
  not g56107 (n_25111, n34004);
  and g56108 (n34006, n_25111, n34005);
  not g56109 (n_25112, n33976);
  not g56110 (n_25113, n34006);
  and g56111 (n34007, n_25112, n_25113);
  not g56112 (n_25114, n34007);
  and g56113 (n34008, n_4226, n_25114);
  and g56114 (n34009, pi0198, po1038);
  or g56115 (po0355, n34008, n34009);
  and g56116 (n34011, pi0199, n_11751);
  not g56117 (n_25115, n34011);
  and g56118 (n34012, n_11821, n_25115);
  not g56119 (n_25117, pi0617);
  and g56120 (n34013, n_25117, n_25115);
  not g56121 (n_25118, n19432);
  and g56122 (n34014, n_7044, n_25118);
  not g56123 (n_25119, n34014);
  and g56124 (n34015, n19438, n_25119);
  and g56125 (n34016, n_7044, n_14476);
  and g56126 (n34017, pi0199, n17221);
  not g56127 (n_25120, n34016);
  and g56128 (n34018, n_161, n_25120);
  not g56129 (n_25121, n34017);
  and g56130 (n34019, n_25121, n34018);
  not g56131 (n_25122, n34015);
  not g56132 (n_25123, n34019);
  and g56133 (n34020, n_25122, n_25123);
  not g56134 (n_25124, n34020);
  and g56135 (n34021, n2571, n_25124);
  and g56136 (n34022, pi0199, n_11417);
  not g56137 (n_25125, n34022);
  and g56138 (n34023, pi0617, n_25125);
  not g56139 (n_25126, n34021);
  and g56140 (n34024, n_25126, n34023);
  not g56141 (n_25127, n34013);
  not g56142 (n_25128, n34024);
  and g56143 (n34025, n_25127, n_25128);
  not g56144 (n_25129, n34025);
  and g56145 (n34026, n_11960, n_25129);
  and g56146 (n34027, n17117, n_25115);
  not g56147 (n_25130, n34026);
  not g56148 (n_25131, n34027);
  and g56149 (n34028, n_25130, n_25131);
  and g56150 (n34029, n_11964, n34028);
  and g56151 (n34030, n_11971, n_25115);
  not g56152 (n_25132, n34028);
  and g56153 (n34031, pi0609, n_25132);
  not g56154 (n_25133, n34030);
  and g56155 (n34032, pi1155, n_25133);
  not g56156 (n_25134, n34031);
  and g56157 (n34033, n_25134, n34032);
  and g56158 (n34034, n_11971, n_25132);
  and g56159 (n34035, pi0609, n_25115);
  not g56160 (n_25135, n34035);
  and g56161 (n34036, n_11768, n_25135);
  not g56162 (n_25136, n34034);
  and g56163 (n34037, n_25136, n34036);
  not g56164 (n_25137, n34033);
  not g56165 (n_25138, n34037);
  and g56166 (n34038, n_25137, n_25138);
  not g56167 (n_25139, n34038);
  and g56168 (n34039, pi0785, n_25139);
  not g56169 (n_25140, n34029);
  not g56170 (n_25141, n34039);
  and g56171 (n34040, n_25140, n_25141);
  not g56172 (n_25142, n34040);
  and g56173 (n34041, n_11981, n_25142);
  and g56174 (n34042, n_11984, n_25115);
  and g56175 (n34043, pi0618, n34040);
  not g56176 (n_25143, n34042);
  and g56177 (n34044, pi1154, n_25143);
  not g56178 (n_25144, n34043);
  and g56179 (n34045, n_25144, n34044);
  and g56180 (n34046, pi0618, n_25115);
  and g56181 (n34047, n_11984, n34040);
  not g56182 (n_25145, n34046);
  and g56183 (n34048, n_11413, n_25145);
  not g56184 (n_25146, n34047);
  and g56185 (n34049, n_25146, n34048);
  not g56186 (n_25147, n34045);
  not g56187 (n_25148, n34049);
  and g56188 (n34050, n_25147, n_25148);
  not g56189 (n_25149, n34050);
  and g56190 (n34051, pi0781, n_25149);
  not g56191 (n_25150, n34041);
  not g56192 (n_25151, n34051);
  and g56193 (n34052, n_25150, n_25151);
  and g56194 (n34053, pi0619, n34052);
  not g56195 (n_25152, n34012);
  and g56196 (n34054, pi1159, n_25152);
  not g56197 (n_25153, n34053);
  and g56198 (n34055, n_25153, n34054);
  and g56199 (n34056, n_11753, n_25115);
  not g56200 (n_25155, pi0637);
  and g56201 (n34057, n_25155, n_25115);
  and g56202 (n34058, n_7044, n_11418);
  not g56203 (n_25156, n34058);
  and g56204 (n34059, n19899, n_25156);
  not g56205 (n_25157, n16840);
  and g56206 (n34060, pi0199, n_25157);
  and g56207 (n34061, n_7044, n_11500);
  not g56208 (n_25158, n34061);
  and g56209 (n34062, pi0039, n_25158);
  not g56210 (n_25159, n34060);
  and g56211 (n34063, n_25159, n34062);
  and g56212 (n34064, pi0199, n_11660);
  and g56213 (n34065, n_7044, n16926);
  not g56214 (n_25160, n34064);
  and g56215 (n34066, n_162, n_25160);
  not g56216 (n_25161, n34065);
  and g56217 (n34067, n_25161, n34066);
  not g56218 (n_25162, n34067);
  and g56219 (n34068, n_161, n_25162);
  not g56220 (n_25163, n34063);
  and g56221 (n34069, n_25163, n34068);
  not g56222 (n_25164, n34059);
  not g56223 (n_25165, n34069);
  and g56224 (n34070, n_25164, n_25165);
  not g56225 (n_25166, n34070);
  and g56226 (n34071, n2571, n_25166);
  and g56227 (n34072, pi0637, n_25125);
  not g56228 (n_25167, n34071);
  and g56229 (n34073, n_25167, n34072);
  not g56230 (n_25168, n34057);
  not g56231 (n_25169, n34073);
  and g56232 (n34074, n_25168, n_25169);
  not g56233 (n_25170, n34074);
  and g56234 (n34075, pi0625, n_25170);
  not g56235 (n_25171, n34056);
  and g56236 (n34076, pi1153, n_25171);
  not g56237 (n_25172, n34075);
  and g56238 (n34077, n_25172, n34076);
  and g56239 (n34078, n_25155, n34025);
  and g56240 (n34079, pi0199, n19476);
  and g56241 (n34080, n2571, n_17658);
  not g56242 (n_25173, n34080);
  and g56243 (n34081, n_7044, n_25173);
  and g56249 (n34085, n2571, n19496);
  not g56250 (n_25176, n34085);
  and g56251 (n34086, n_7044, n_25176);
  and g56252 (n34087, pi0199, n19488);
  not g56253 (n_25177, n34087);
  and g56254 (n34088, pi0617, n_25177);
  not g56255 (n_25178, n34086);
  and g56256 (n34089, n_25178, n34088);
  not g56257 (n_25179, n34089);
  and g56258 (n34090, n_25125, n_25179);
  not g56259 (n_25180, n34084);
  and g56260 (n34091, n_25180, n34090);
  not g56261 (n_25181, n34091);
  and g56262 (n34092, pi0637, n_25181);
  not g56263 (n_25182, n34078);
  not g56264 (n_25183, n34092);
  and g56265 (n34093, n_25182, n_25183);
  and g56266 (n34094, n_11753, n34093);
  and g56267 (n34095, pi0625, n_25129);
  not g56268 (n_25184, n34095);
  and g56269 (n34096, n_11757, n_25184);
  not g56270 (n_25185, n34094);
  and g56271 (n34097, n_25185, n34096);
  not g56272 (n_25186, n34077);
  and g56273 (n34098, n_11823, n_25186);
  not g56274 (n_25187, n34097);
  and g56275 (n34099, n_25187, n34098);
  and g56276 (n34100, n_11753, n_25170);
  and g56277 (n34101, pi0625, n_25115);
  not g56278 (n_25188, n34101);
  and g56279 (n34102, n_11757, n_25188);
  not g56280 (n_25189, n34100);
  and g56281 (n34103, n_25189, n34102);
  and g56282 (n34104, pi0625, n34093);
  and g56283 (n34105, n_11753, n_25129);
  not g56284 (n_25190, n34105);
  and g56285 (n34106, pi1153, n_25190);
  not g56286 (n_25191, n34104);
  and g56287 (n34107, n_25191, n34106);
  not g56288 (n_25192, n34103);
  and g56289 (n34108, pi0608, n_25192);
  not g56290 (n_25193, n34107);
  and g56291 (n34109, n_25193, n34108);
  not g56292 (n_25194, n34099);
  not g56293 (n_25195, n34109);
  and g56294 (n34110, n_25194, n_25195);
  not g56295 (n_25196, n34110);
  and g56296 (n34111, pi0778, n_25196);
  and g56297 (n34112, n_11749, n34093);
  not g56298 (n_25197, n34111);
  not g56299 (n_25198, n34112);
  and g56300 (n34113, n_25197, n_25198);
  not g56301 (n_25199, n34113);
  and g56302 (n34114, n_11971, n_25199);
  and g56303 (n34115, n_11749, n34074);
  and g56304 (n34116, n_25186, n_25192);
  not g56305 (n_25200, n34116);
  and g56306 (n34117, pi0778, n_25200);
  not g56307 (n_25201, n34115);
  not g56308 (n_25202, n34117);
  and g56309 (n34118, n_25201, n_25202);
  and g56310 (n34119, pi0609, n34118);
  not g56311 (n_25203, n34119);
  and g56312 (n34120, n_11768, n_25203);
  not g56313 (n_25204, n34114);
  and g56314 (n34121, n_25204, n34120);
  and g56315 (n34122, n_11767, n_25137);
  not g56316 (n_25205, n34121);
  and g56317 (n34123, n_25205, n34122);
  and g56318 (n34124, n_11971, n34118);
  and g56319 (n34125, pi0609, n_25199);
  not g56320 (n_25206, n34124);
  and g56321 (n34126, pi1155, n_25206);
  not g56322 (n_25207, n34125);
  and g56323 (n34127, n_25207, n34126);
  and g56324 (n34128, pi0660, n_25138);
  not g56325 (n_25208, n34127);
  and g56326 (n34129, n_25208, n34128);
  not g56327 (n_25209, n34123);
  not g56328 (n_25210, n34129);
  and g56329 (n34130, n_25209, n_25210);
  not g56330 (n_25211, n34130);
  and g56331 (n34131, pi0785, n_25211);
  and g56332 (n34132, n_11964, n_25199);
  not g56333 (n_25212, n34131);
  not g56334 (n_25213, n34132);
  and g56335 (n34133, n_25212, n_25213);
  not g56336 (n_25214, n34133);
  and g56337 (n34134, n_11984, n_25214);
  and g56338 (n34135, n17075, n_25115);
  and g56339 (n34136, n_11773, n34118);
  not g56340 (n_25215, n34135);
  not g56341 (n_25216, n34136);
  and g56342 (n34137, n_25215, n_25216);
  not g56343 (n_25217, n34137);
  and g56344 (n34138, pi0618, n_25217);
  not g56345 (n_25218, n34138);
  and g56346 (n34139, n_11413, n_25218);
  not g56347 (n_25219, n34134);
  and g56348 (n34140, n_25219, n34139);
  and g56349 (n34141, n_11412, n_25147);
  not g56350 (n_25220, n34140);
  and g56351 (n34142, n_25220, n34141);
  and g56352 (n34143, pi0618, n_25214);
  and g56353 (n34144, n_11984, n_25217);
  not g56354 (n_25221, n34144);
  and g56355 (n34145, pi1154, n_25221);
  not g56356 (n_25222, n34143);
  and g56357 (n34146, n_25222, n34145);
  and g56358 (n34147, pi0627, n_25148);
  not g56359 (n_25223, n34146);
  and g56360 (n34148, n_25223, n34147);
  not g56361 (n_25224, n34142);
  not g56362 (n_25225, n34148);
  and g56363 (n34149, n_25224, n_25225);
  not g56364 (n_25226, n34149);
  and g56365 (n34150, pi0781, n_25226);
  and g56366 (n34151, n_11981, n_25214);
  not g56367 (n_25227, n34150);
  not g56368 (n_25228, n34151);
  and g56369 (n34152, n_25227, n_25228);
  not g56370 (n_25229, n34152);
  and g56371 (n34153, n_11821, n_25229);
  and g56372 (n34154, n_11777, n34137);
  and g56373 (n34155, n16639, n34011);
  not g56374 (n_25230, n34154);
  not g56375 (n_25231, n34155);
  and g56376 (n34156, n_25230, n_25231);
  and g56377 (n34157, pi0619, n34156);
  not g56378 (n_25232, n34157);
  and g56379 (n34158, n_11405, n_25232);
  not g56380 (n_25233, n34153);
  and g56381 (n34159, n_25233, n34158);
  not g56382 (n_25234, n34055);
  and g56383 (n34160, n_11403, n_25234);
  not g56384 (n_25235, n34159);
  and g56385 (n34161, n_25235, n34160);
  and g56386 (n34162, pi0619, n_25115);
  and g56387 (n34163, n_11821, n34052);
  not g56388 (n_25236, n34162);
  and g56389 (n34164, n_11405, n_25236);
  not g56390 (n_25237, n34163);
  and g56391 (n34165, n_25237, n34164);
  and g56392 (n34166, n_11821, n34156);
  and g56393 (n34167, pi0619, n_25229);
  not g56394 (n_25238, n34166);
  and g56395 (n34168, pi1159, n_25238);
  not g56396 (n_25239, n34167);
  and g56397 (n34169, n_25239, n34168);
  not g56398 (n_25240, n34165);
  and g56399 (n34170, pi0648, n_25240);
  not g56400 (n_25241, n34169);
  and g56401 (n34171, n_25241, n34170);
  not g56402 (n_25242, n34161);
  not g56403 (n_25243, n34171);
  and g56404 (n34172, n_25242, n_25243);
  not g56405 (n_25244, n34172);
  and g56406 (n34173, pi0789, n_25244);
  and g56407 (n34174, n_12315, n_25229);
  not g56408 (n_25245, n34173);
  not g56409 (n_25246, n34174);
  and g56410 (n34175, n_25245, n_25246);
  and g56411 (n34176, n_12318, n34175);
  and g56412 (n34177, n_12320, n34175);
  and g56413 (n34178, n16635, n_25115);
  and g56414 (n34179, n_11780, n34156);
  not g56415 (n_25247, n34178);
  not g56416 (n_25248, n34179);
  and g56417 (n34180, n_25247, n_25248);
  and g56418 (n34181, pi0626, n34180);
  not g56419 (n_25249, n34181);
  and g56420 (n34182, n_11395, n_25249);
  not g56421 (n_25250, n34177);
  and g56422 (n34183, n_25250, n34182);
  not g56423 (n_25251, n34052);
  and g56424 (n34184, n_12315, n_25251);
  and g56425 (n34185, n_25234, n_25240);
  not g56426 (n_25252, n34185);
  and g56427 (n34186, pi0789, n_25252);
  not g56428 (n_25253, n34184);
  not g56429 (n_25254, n34186);
  and g56430 (n34187, n_25253, n_25254);
  not g56431 (n_25255, n34187);
  and g56432 (n34188, n_12320, n_25255);
  and g56433 (n34189, pi0626, n34011);
  not g56434 (n_25256, n34189);
  and g56435 (n34190, pi0641, n_25256);
  not g56436 (n_25257, n34188);
  and g56437 (n34191, n_25257, n34190);
  not g56438 (n_25258, n34191);
  and g56439 (n34192, n_11397, n_25258);
  not g56440 (n_25259, n34183);
  and g56441 (n34193, n_25259, n34192);
  and g56442 (n34194, n_12320, n34180);
  and g56443 (n34195, pi0626, n34175);
  not g56444 (n_25260, n34194);
  and g56445 (n34196, pi0641, n_25260);
  not g56446 (n_25261, n34195);
  and g56447 (n34197, n_25261, n34196);
  and g56448 (n34198, pi0626, n_25255);
  and g56449 (n34199, n_12320, n34011);
  not g56450 (n_25262, n34199);
  and g56451 (n34200, n_11395, n_25262);
  not g56452 (n_25263, n34198);
  and g56453 (n34201, n_25263, n34200);
  not g56454 (n_25264, n34201);
  and g56455 (n34202, pi1158, n_25264);
  not g56456 (n_25265, n34197);
  and g56457 (n34203, n_25265, n34202);
  not g56458 (n_25266, n34193);
  not g56459 (n_25267, n34203);
  and g56460 (n34204, n_25266, n_25267);
  not g56461 (n_25268, n34204);
  and g56462 (n34205, pi0788, n_25268);
  not g56463 (n_25269, n34176);
  not g56464 (n_25270, n34205);
  and g56465 (n34206, n_25269, n_25270);
  and g56466 (n34207, n_11789, n34206);
  and g56467 (n34208, n_12524, n_25255);
  and g56468 (n34209, n17969, n34011);
  not g56469 (n_25271, n34208);
  not g56470 (n_25272, n34209);
  and g56471 (n34210, n_25271, n_25272);
  and g56472 (n34211, pi0628, n34210);
  not g56473 (n_25273, n34211);
  and g56474 (n34212, n_11794, n_25273);
  not g56475 (n_25274, n34207);
  and g56476 (n34213, n_25274, n34212);
  and g56477 (n34214, n_11789, n_25115);
  and g56478 (n34215, n_11783, n34180);
  and g56479 (n34216, n16631, n34011);
  not g56480 (n_25275, n34215);
  not g56481 (n_25276, n34216);
  and g56482 (n34217, n_25275, n_25276);
  and g56483 (n34218, pi0628, n34217);
  not g56484 (n_25277, n34214);
  and g56485 (n34219, pi1156, n_25277);
  not g56486 (n_25278, n34218);
  and g56487 (n34220, n_25278, n34219);
  not g56488 (n_25279, n34220);
  and g56489 (n34221, n_12354, n_25279);
  not g56490 (n_25280, n34213);
  and g56491 (n34222, n_25280, n34221);
  and g56492 (n34223, pi0628, n34206);
  and g56493 (n34224, n_11789, n34210);
  not g56494 (n_25281, n34224);
  and g56495 (n34225, pi1156, n_25281);
  not g56496 (n_25282, n34223);
  and g56497 (n34226, n_25282, n34225);
  and g56498 (n34227, pi0628, n_25115);
  and g56499 (n34228, n_11789, n34217);
  not g56500 (n_25283, n34227);
  and g56501 (n34229, n_11794, n_25283);
  not g56502 (n_25284, n34228);
  and g56503 (n34230, n_25284, n34229);
  not g56504 (n_25285, n34230);
  and g56505 (n34231, pi0629, n_25285);
  not g56506 (n_25286, n34226);
  and g56507 (n34232, n_25286, n34231);
  not g56508 (n_25287, n34222);
  not g56509 (n_25288, n34232);
  and g56510 (n34233, n_25287, n_25288);
  not g56511 (n_25289, n34233);
  and g56512 (n34234, pi0792, n_25289);
  and g56513 (n34235, n_11787, n34206);
  not g56514 (n_25290, n34234);
  not g56515 (n_25291, n34235);
  and g56516 (n34236, n_25290, n_25291);
  not g56517 (n_25292, n34236);
  and g56518 (n34237, n_11806, n_25292);
  not g56519 (n_25293, n34210);
  and g56520 (n34238, n_12368, n_25293);
  and g56521 (n34239, n17779, n34011);
  not g56522 (n_25294, n34238);
  not g56523 (n_25295, n34239);
  and g56524 (n34240, n_25294, n_25295);
  and g56525 (n34241, pi0647, n34240);
  not g56526 (n_25296, n34241);
  and g56527 (n34242, n_11810, n_25296);
  not g56528 (n_25297, n34237);
  and g56529 (n34243, n_25297, n34242);
  and g56530 (n34244, n_11806, n_25115);
  not g56531 (n_25298, n34217);
  and g56532 (n34245, n_11787, n_25298);
  and g56533 (n34246, n_25279, n_25285);
  not g56534 (n_25299, n34246);
  and g56535 (n34247, pi0792, n_25299);
  not g56536 (n_25300, n34245);
  not g56537 (n_25301, n34247);
  and g56538 (n34248, n_25300, n_25301);
  and g56539 (n34249, pi0647, n34248);
  not g56540 (n_25302, n34244);
  and g56541 (n34250, pi1157, n_25302);
  not g56542 (n_25303, n34249);
  and g56543 (n34251, n_25303, n34250);
  not g56544 (n_25304, n34251);
  and g56545 (n34252, n_12375, n_25304);
  not g56546 (n_25305, n34243);
  and g56547 (n34253, n_25305, n34252);
  and g56548 (n34254, pi0647, n_25292);
  and g56549 (n34255, n_11806, n34240);
  not g56550 (n_25306, n34255);
  and g56551 (n34256, pi1157, n_25306);
  not g56552 (n_25307, n34254);
  and g56553 (n34257, n_25307, n34256);
  and g56554 (n34258, pi0647, n_25115);
  and g56555 (n34259, n_11806, n34248);
  not g56556 (n_25308, n34258);
  and g56557 (n34260, n_11810, n_25308);
  not g56558 (n_25309, n34259);
  and g56559 (n34261, n_25309, n34260);
  not g56560 (n_25310, n34261);
  and g56561 (n34262, pi0630, n_25310);
  not g56562 (n_25311, n34257);
  and g56563 (n34263, n_25311, n34262);
  not g56564 (n_25312, n34253);
  not g56565 (n_25313, n34263);
  and g56566 (n34264, n_25312, n_25313);
  not g56567 (n_25314, n34264);
  and g56568 (n34265, pi0787, n_25314);
  and g56569 (n34266, n_11803, n_25292);
  not g56570 (n_25315, n34265);
  not g56571 (n_25316, n34266);
  and g56572 (n34267, n_25315, n_25316);
  and g56573 (n34268, n_12411, n34267);
  not g56574 (n_25317, n34248);
  and g56575 (n34269, n_11803, n_25317);
  and g56576 (n34270, n_25304, n_25310);
  not g56577 (n_25318, n34270);
  and g56578 (n34271, pi0787, n_25318);
  not g56579 (n_25319, n34269);
  not g56580 (n_25320, n34271);
  and g56581 (n34272, n_25319, n_25320);
  and g56582 (n34273, n_11819, n34272);
  not g56583 (n_25321, n34267);
  and g56584 (n34274, pi0644, n_25321);
  not g56585 (n_25322, n34273);
  and g56586 (n34275, pi0715, n_25322);
  not g56587 (n_25323, n34274);
  and g56588 (n34276, n_25323, n34275);
  and g56589 (n34277, n17804, n_25115);
  and g56590 (n34278, n_12392, n34240);
  not g56591 (n_25324, n34277);
  not g56592 (n_25325, n34278);
  and g56593 (n34279, n_25324, n_25325);
  not g56594 (n_25326, n34279);
  and g56595 (n34280, pi0644, n_25326);
  and g56596 (n34281, n_11819, n_25115);
  not g56597 (n_25327, n34281);
  and g56598 (n34282, n_12395, n_25327);
  not g56599 (n_25328, n34280);
  and g56600 (n34283, n_25328, n34282);
  not g56601 (n_25329, n34283);
  and g56602 (n34284, pi1160, n_25329);
  not g56603 (n_25330, n34276);
  and g56604 (n34285, n_25330, n34284);
  and g56605 (n34286, n_11819, n_25321);
  and g56606 (n34287, pi0644, n34272);
  not g56607 (n_25331, n34287);
  and g56608 (n34288, n_12395, n_25331);
  not g56609 (n_25332, n34286);
  and g56610 (n34289, n_25332, n34288);
  and g56611 (n34290, n_11819, n_25326);
  and g56612 (n34291, pi0644, n_25115);
  not g56613 (n_25333, n34291);
  and g56614 (n34292, pi0715, n_25333);
  not g56615 (n_25334, n34290);
  and g56616 (n34293, n_25334, n34292);
  not g56617 (n_25335, n34293);
  and g56618 (n34294, n_12405, n_25335);
  not g56619 (n_25336, n34289);
  and g56620 (n34295, n_25336, n34294);
  not g56621 (n_25337, n34285);
  and g56622 (n34296, pi0790, n_25337);
  not g56623 (n_25338, n34295);
  and g56624 (n34297, n_25338, n34296);
  not g56625 (n_25339, n34268);
  not g56626 (n_25340, n34297);
  and g56627 (n34298, n_25339, n_25340);
  not g56628 (n_25341, n34298);
  and g56629 (n34299, n_4226, n_25341);
  and g56630 (n34300, pi0199, po1038);
  or g56631 (po0356, n34299, n34300);
  and g56632 (n34302, pi0200, n_11751);
  not g56633 (n_25343, pi0606);
  not g56634 (n_25344, n34302);
  and g56635 (n34303, n_25343, n_25344);
  and g56636 (n34304, pi0200, n_11417);
  and g56637 (n34305, n_7045, n_25118);
  not g56638 (n_25345, n34305);
  and g56639 (n34306, n19438, n_25345);
  and g56640 (n34307, n_7045, n_14476);
  and g56641 (n34308, pi0200, n17221);
  not g56642 (n_25346, n34307);
  and g56643 (n34309, n_161, n_25346);
  not g56644 (n_25347, n34308);
  and g56645 (n34310, n_25347, n34309);
  not g56646 (n_25348, n34306);
  not g56647 (n_25349, n34310);
  and g56648 (n34311, n_25348, n_25349);
  not g56649 (n_25350, n34311);
  and g56650 (n34312, n2571, n_25350);
  not g56651 (n_25351, n34304);
  and g56652 (n34313, pi0606, n_25351);
  not g56653 (n_25352, n34312);
  and g56654 (n34314, n_25352, n34313);
  not g56655 (n_25353, n34303);
  not g56656 (n_25354, n34314);
  and g56657 (n34315, n_25353, n_25354);
  not g56658 (n_25355, n34315);
  and g56659 (n34316, n_11960, n_25355);
  and g56660 (n34317, n17117, n_25344);
  not g56661 (n_25356, n34316);
  not g56662 (n_25357, n34317);
  and g56663 (n34318, n_25356, n_25357);
  and g56664 (n34319, n_11964, n34318);
  and g56665 (n34320, n_11971, n_25344);
  not g56666 (n_25358, n34318);
  and g56667 (n34321, pi0609, n_25358);
  not g56668 (n_25359, n34320);
  and g56669 (n34322, pi1155, n_25359);
  not g56670 (n_25360, n34321);
  and g56671 (n34323, n_25360, n34322);
  and g56672 (n34324, n_11971, n_25358);
  and g56673 (n34325, pi0609, n_25344);
  not g56674 (n_25361, n34325);
  and g56675 (n34326, n_11768, n_25361);
  not g56676 (n_25362, n34324);
  and g56677 (n34327, n_25362, n34326);
  not g56678 (n_25363, n34323);
  not g56679 (n_25364, n34327);
  and g56680 (n34328, n_25363, n_25364);
  not g56681 (n_25365, n34328);
  and g56682 (n34329, pi0785, n_25365);
  not g56683 (n_25366, n34319);
  not g56684 (n_25367, n34329);
  and g56685 (n34330, n_25366, n_25367);
  not g56686 (n_25368, n34330);
  and g56687 (n34331, n_11981, n_25368);
  and g56688 (n34332, n_11984, n_25344);
  and g56689 (n34333, pi0618, n34330);
  not g56690 (n_25369, n34332);
  and g56691 (n34334, pi1154, n_25369);
  not g56692 (n_25370, n34333);
  and g56693 (n34335, n_25370, n34334);
  and g56694 (n34336, pi0618, n_25344);
  and g56695 (n34337, n_11984, n34330);
  not g56696 (n_25371, n34336);
  and g56697 (n34338, n_11413, n_25371);
  not g56698 (n_25372, n34337);
  and g56699 (n34339, n_25372, n34338);
  not g56700 (n_25373, n34335);
  not g56701 (n_25374, n34339);
  and g56702 (n34340, n_25373, n_25374);
  not g56703 (n_25375, n34340);
  and g56704 (n34341, pi0781, n_25375);
  not g56705 (n_25376, n34331);
  not g56706 (n_25377, n34341);
  and g56707 (n34342, n_25376, n_25377);
  not g56708 (n_25378, n34342);
  and g56709 (n34343, n_12315, n_25378);
  and g56710 (n34344, n_11821, n_25344);
  and g56711 (n34345, pi0619, n34342);
  not g56712 (n_25379, n34344);
  and g56713 (n34346, pi1159, n_25379);
  not g56714 (n_25380, n34345);
  and g56715 (n34347, n_25380, n34346);
  and g56716 (n34348, pi0619, n_25344);
  and g56717 (n34349, n_11821, n34342);
  not g56718 (n_25381, n34348);
  and g56719 (n34350, n_11405, n_25381);
  not g56720 (n_25382, n34349);
  and g56721 (n34351, n_25382, n34350);
  not g56722 (n_25383, n34347);
  not g56723 (n_25384, n34351);
  and g56724 (n34352, n_25383, n_25384);
  not g56725 (n_25385, n34352);
  and g56726 (n34353, pi0789, n_25385);
  not g56727 (n_25386, n34343);
  not g56728 (n_25387, n34353);
  and g56729 (n34354, n_25386, n_25387);
  not g56730 (n_25388, n34354);
  and g56731 (n34355, n_12524, n_25388);
  and g56732 (n34356, n17969, n34302);
  not g56733 (n_25389, n34355);
  not g56734 (n_25390, n34356);
  and g56735 (n34357, n_25389, n_25390);
  not g56736 (n_25391, n34357);
  and g56737 (n34358, n_12368, n_25391);
  and g56738 (n34359, n17779, n34302);
  not g56739 (n_25392, n34358);
  not g56740 (n_25393, n34359);
  and g56741 (n34360, n_25392, n_25393);
  not g56742 (n_25394, n34360);
  and g56743 (n34361, n_12392, n_25394);
  and g56744 (n34362, n17804, n34302);
  not g56745 (n_25395, n34361);
  not g56746 (n_25396, n34362);
  and g56747 (n34363, n_25395, n_25396);
  and g56748 (n34364, n_11819, n34363);
  and g56749 (n34365, pi0644, n_25344);
  not g56750 (n_25397, n34365);
  and g56751 (n34366, pi0715, n_25397);
  not g56752 (n_25398, n34364);
  and g56753 (n34367, n_25398, n34366);
  and g56754 (n34368, n16635, n_25344);
  and g56755 (n34369, n17075, n_25344);
  not g56756 (n_25400, pi0643);
  and g56757 (n34370, n_25400, n_25344);
  and g56758 (n34371, n_7045, n_11418);
  not g56759 (n_25401, n34371);
  and g56760 (n34372, n19899, n_25401);
  and g56761 (n34373, n_7045, n16733);
  and g56762 (n34374, pi0200, n16823);
  not g56763 (n_25402, n34373);
  and g56764 (n34375, n_234, n_25402);
  not g56765 (n_25403, n34374);
  and g56766 (n34376, n_25403, n34375);
  and g56767 (n34377, n_7045, n16747);
  and g56768 (n34378, pi0200, n16838);
  not g56769 (n_25404, n34377);
  and g56770 (n34379, pi0299, n_25404);
  not g56771 (n_25405, n34378);
  and g56772 (n34380, n_25405, n34379);
  not g56773 (n_25406, n34376);
  not g56774 (n_25407, n34380);
  and g56775 (n34381, n_25406, n_25407);
  not g56776 (n_25408, n34381);
  and g56777 (n34382, pi0039, n_25408);
  and g56778 (n34383, n_7045, n_12243);
  and g56779 (n34384, pi0200, n16948);
  not g56780 (n_25409, n34383);
  and g56781 (n34385, n_162, n_25409);
  not g56782 (n_25410, n34384);
  and g56783 (n34386, n_25410, n34385);
  not g56784 (n_25411, n34382);
  not g56785 (n_25412, n34386);
  and g56786 (n34387, n_25411, n_25412);
  not g56787 (n_25413, n34387);
  and g56788 (n34388, n_161, n_25413);
  not g56789 (n_25414, n34372);
  not g56790 (n_25415, n34388);
  and g56791 (n34389, n_25414, n_25415);
  not g56792 (n_25416, n34389);
  and g56793 (n34390, n2571, n_25416);
  and g56794 (n34391, pi0643, n_25351);
  not g56795 (n_25417, n34390);
  and g56796 (n34392, n_25417, n34391);
  not g56797 (n_25418, n34370);
  not g56798 (n_25419, n34392);
  and g56799 (n34393, n_25418, n_25419);
  and g56800 (n34394, n_11749, n34393);
  and g56801 (n34395, n_11753, n_25344);
  not g56802 (n_25420, n34393);
  and g56803 (n34396, pi0625, n_25420);
  not g56804 (n_25421, n34395);
  and g56805 (n34397, pi1153, n_25421);
  not g56806 (n_25422, n34396);
  and g56807 (n34398, n_25422, n34397);
  and g56808 (n34399, n_11753, n_25420);
  and g56809 (n34400, pi0625, n_25344);
  not g56810 (n_25423, n34400);
  and g56811 (n34401, n_11757, n_25423);
  not g56812 (n_25424, n34399);
  and g56813 (n34402, n_25424, n34401);
  not g56814 (n_25425, n34398);
  not g56815 (n_25426, n34402);
  and g56816 (n34403, n_25425, n_25426);
  not g56817 (n_25427, n34403);
  and g56818 (n34404, pi0778, n_25427);
  not g56819 (n_25428, n34394);
  not g56820 (n_25429, n34404);
  and g56821 (n34405, n_25428, n_25429);
  and g56822 (n34406, n_11773, n34405);
  not g56823 (n_25430, n34369);
  not g56824 (n_25431, n34406);
  and g56825 (n34407, n_25430, n_25431);
  and g56826 (n34408, n_11777, n34407);
  and g56827 (n34409, n16639, n34302);
  not g56828 (n_25432, n34408);
  not g56829 (n_25433, n34409);
  and g56830 (n34410, n_25432, n_25433);
  and g56831 (n34411, n_11780, n34410);
  not g56832 (n_25434, n34368);
  not g56833 (n_25435, n34411);
  and g56834 (n34412, n_25434, n_25435);
  and g56835 (n34413, n_11783, n34412);
  and g56836 (n34414, n16631, n34302);
  not g56837 (n_25436, n34413);
  not g56838 (n_25437, n34414);
  and g56839 (n34415, n_25436, n_25437);
  not g56840 (n_25438, n34415);
  and g56841 (n34416, n_11787, n_25438);
  and g56842 (n34417, pi0628, n_25344);
  and g56843 (n34418, n_11789, n34415);
  not g56844 (n_25439, n34417);
  and g56845 (n34419, n_11794, n_25439);
  not g56846 (n_25440, n34418);
  and g56847 (n34420, n_25440, n34419);
  and g56848 (n34421, n_11789, n_25344);
  and g56849 (n34422, pi0628, n34415);
  not g56850 (n_25441, n34421);
  and g56851 (n34423, pi1156, n_25441);
  not g56852 (n_25442, n34422);
  and g56853 (n34424, n_25442, n34423);
  not g56854 (n_25443, n34420);
  not g56855 (n_25444, n34424);
  and g56856 (n34425, n_25443, n_25444);
  not g56857 (n_25445, n34425);
  and g56858 (n34426, pi0792, n_25445);
  not g56859 (n_25446, n34416);
  not g56860 (n_25447, n34426);
  and g56861 (n34427, n_25446, n_25447);
  not g56862 (n_25448, n34427);
  and g56863 (n34428, n_11803, n_25448);
  and g56864 (n34429, pi0647, n_25448);
  and g56865 (n34430, n_11806, n34302);
  not g56866 (n_25449, n34429);
  not g56867 (n_25450, n34430);
  and g56868 (n34431, n_25449, n_25450);
  not g56869 (n_25451, n34431);
  and g56870 (n34432, pi1157, n_25451);
  and g56871 (n34433, pi0647, n_25344);
  and g56872 (n34434, n_11806, n34427);
  not g56873 (n_25452, n34433);
  and g56874 (n34435, n_11810, n_25452);
  not g56875 (n_25453, n34434);
  and g56876 (n34436, n_25453, n34435);
  not g56877 (n_25454, n34432);
  not g56878 (n_25455, n34436);
  and g56879 (n34437, n_25454, n_25455);
  not g56880 (n_25456, n34437);
  and g56881 (n34438, pi0787, n_25456);
  not g56882 (n_25457, n34428);
  not g56883 (n_25458, n34438);
  and g56884 (n34439, n_25457, n_25458);
  and g56885 (n34440, pi0644, n34439);
  and g56886 (n34441, n_12354, n34424);
  and g56887 (n34442, n_14557, n_25391);
  and g56888 (n34443, pi0629, n34420);
  not g56889 (n_25459, n34441);
  not g56890 (n_25460, n34443);
  and g56891 (n34444, n_25459, n_25460);
  not g56892 (n_25461, n34442);
  and g56893 (n34445, n_25461, n34444);
  not g56894 (n_25462, n34445);
  and g56895 (n34446, pi0792, n_25462);
  and g56896 (n34447, pi0609, n34405);
  and g56897 (n34448, n_25400, n34315);
  and g56898 (n34449, n_13724, n_13721);
  not g56899 (n_25463, n34449);
  and g56900 (n34450, n_7045, n_25463);
  and g56901 (n34451, pi0038, pi0200);
  and g56902 (n34452, n19485, n34451);
  and g56903 (n34453, n_7045, n_13722);
  and g56904 (n34454, pi0200, n_17822);
  not g56905 (n_25464, n34453);
  and g56906 (n34455, n_161, n_25464);
  not g56907 (n_25465, n34454);
  and g56908 (n34456, n_25465, n34455);
  and g56916 (n34461, n_17518, n_12023);
  not g56917 (n_25469, n34461);
  and g56918 (n34462, n34372, n_25469);
  not g56919 (n_25470, n19467);
  and g56920 (n34463, n_7045, n_25470);
  and g56921 (n34464, pi0200, n_13708);
  not g56922 (n_25471, n34463);
  and g56923 (n34465, n_161, n_25471);
  not g56924 (n_25472, n34464);
  and g56925 (n34466, n_25472, n34465);
  not g56926 (n_25473, n34462);
  not g56927 (n_25474, n34466);
  and g56928 (n34467, n_25473, n_25474);
  and g56929 (n34468, n_25343, n2571);
  not g56930 (n_25475, n34467);
  and g56931 (n34469, n_25475, n34468);
  not g56932 (n_25476, n34460);
  and g56933 (n34470, n_25351, n_25476);
  not g56934 (n_25477, n34469);
  and g56935 (n34471, n_25477, n34470);
  not g56936 (n_25478, n34471);
  and g56937 (n34472, pi0643, n_25478);
  not g56938 (n_25479, n34448);
  not g56939 (n_25480, n34472);
  and g56940 (n34473, n_25479, n_25480);
  and g56941 (n34474, n_11753, n34473);
  and g56942 (n34475, pi0625, n_25355);
  not g56943 (n_25481, n34475);
  and g56944 (n34476, n_11757, n_25481);
  not g56945 (n_25482, n34474);
  and g56946 (n34477, n_25482, n34476);
  and g56947 (n34478, n_11823, n_25425);
  not g56948 (n_25483, n34477);
  and g56949 (n34479, n_25483, n34478);
  and g56950 (n34480, pi0625, n34473);
  and g56951 (n34481, n_11753, n_25355);
  not g56952 (n_25484, n34481);
  and g56953 (n34482, pi1153, n_25484);
  not g56954 (n_25485, n34480);
  and g56955 (n34483, n_25485, n34482);
  and g56956 (n34484, pi0608, n_25426);
  not g56957 (n_25486, n34483);
  and g56958 (n34485, n_25486, n34484);
  not g56959 (n_25487, n34479);
  not g56960 (n_25488, n34485);
  and g56961 (n34486, n_25487, n_25488);
  not g56962 (n_25489, n34486);
  and g56963 (n34487, pi0778, n_25489);
  and g56964 (n34488, n_11749, n34473);
  not g56965 (n_25490, n34487);
  not g56966 (n_25491, n34488);
  and g56967 (n34489, n_25490, n_25491);
  not g56968 (n_25492, n34489);
  and g56969 (n34490, n_11971, n_25492);
  not g56970 (n_25493, n34447);
  and g56971 (n34491, n_11768, n_25493);
  not g56972 (n_25494, n34490);
  and g56973 (n34492, n_25494, n34491);
  and g56974 (n34493, n_11767, n_25363);
  not g56975 (n_25495, n34492);
  and g56976 (n34494, n_25495, n34493);
  and g56977 (n34495, n_11971, n34405);
  and g56978 (n34496, pi0609, n_25492);
  not g56979 (n_25496, n34495);
  and g56980 (n34497, pi1155, n_25496);
  not g56981 (n_25497, n34496);
  and g56982 (n34498, n_25497, n34497);
  and g56983 (n34499, pi0660, n_25364);
  not g56984 (n_25498, n34498);
  and g56985 (n34500, n_25498, n34499);
  not g56986 (n_25499, n34494);
  not g56987 (n_25500, n34500);
  and g56988 (n34501, n_25499, n_25500);
  not g56989 (n_25501, n34501);
  and g56990 (n34502, pi0785, n_25501);
  and g56991 (n34503, n_11964, n_25492);
  not g56992 (n_25502, n34502);
  not g56993 (n_25503, n34503);
  and g56994 (n34504, n_25502, n_25503);
  not g56995 (n_25504, n34504);
  and g56996 (n34505, n_11984, n_25504);
  not g56997 (n_25505, n34407);
  and g56998 (n34506, pi0618, n_25505);
  not g56999 (n_25506, n34506);
  and g57000 (n34507, n_11413, n_25506);
  not g57001 (n_25507, n34505);
  and g57002 (n34508, n_25507, n34507);
  and g57003 (n34509, n_11412, n_25373);
  not g57004 (n_25508, n34508);
  and g57005 (n34510, n_25508, n34509);
  and g57006 (n34511, pi0618, n_25504);
  and g57007 (n34512, n_11984, n_25505);
  not g57008 (n_25509, n34512);
  and g57009 (n34513, pi1154, n_25509);
  not g57010 (n_25510, n34511);
  and g57011 (n34514, n_25510, n34513);
  and g57012 (n34515, pi0627, n_25374);
  not g57013 (n_25511, n34514);
  and g57014 (n34516, n_25511, n34515);
  not g57015 (n_25512, n34510);
  not g57016 (n_25513, n34516);
  and g57017 (n34517, n_25512, n_25513);
  not g57018 (n_25514, n34517);
  and g57019 (n34518, pi0781, n_25514);
  and g57020 (n34519, n_11981, n_25504);
  not g57021 (n_25515, n34518);
  not g57022 (n_25516, n34519);
  and g57023 (n34520, n_25515, n_25516);
  and g57024 (n34521, n_12315, n34520);
  not g57025 (n_25517, n34520);
  and g57026 (n34522, n_11821, n_25517);
  and g57027 (n34523, pi0619, n34410);
  not g57028 (n_25518, n34523);
  and g57029 (n34524, n_11405, n_25518);
  not g57030 (n_25519, n34522);
  and g57031 (n34525, n_25519, n34524);
  and g57032 (n34526, n_11403, n_25383);
  not g57033 (n_25520, n34525);
  and g57034 (n34527, n_25520, n34526);
  and g57035 (n34528, pi0619, n_25517);
  and g57036 (n34529, n_11821, n34410);
  not g57037 (n_25521, n34529);
  and g57038 (n34530, pi1159, n_25521);
  not g57039 (n_25522, n34528);
  and g57040 (n34531, n_25522, n34530);
  and g57041 (n34532, pi0648, n_25384);
  not g57042 (n_25523, n34531);
  and g57043 (n34533, n_25523, n34532);
  not g57044 (n_25524, n34527);
  and g57045 (n34534, pi0789, n_25524);
  not g57046 (n_25525, n34533);
  and g57047 (n34535, n_25525, n34534);
  not g57048 (n_25526, n34521);
  and g57049 (n34536, n17970, n_25526);
  not g57050 (n_25527, n34535);
  and g57051 (n34537, n_25527, n34536);
  not g57052 (n_25528, n34412);
  and g57053 (n34538, n17871, n_25528);
  and g57054 (n34539, pi0626, n34302);
  and g57055 (n34540, n_12320, n_25388);
  not g57056 (n_25529, n34539);
  and g57057 (n34541, n16629, n_25529);
  not g57058 (n_25530, n34540);
  and g57059 (n34542, n_25530, n34541);
  and g57060 (n34543, n_12320, n34302);
  and g57061 (n34544, pi0626, n_25388);
  not g57062 (n_25531, n34543);
  and g57063 (n34545, n16628, n_25531);
  not g57064 (n_25532, n34544);
  and g57065 (n34546, n_25532, n34545);
  not g57066 (n_25533, n34538);
  not g57067 (n_25534, n34542);
  and g57068 (n34547, n_25533, n_25534);
  not g57069 (n_25535, n34546);
  and g57070 (n34548, n_25535, n34547);
  not g57071 (n_25536, n34548);
  and g57072 (n34549, pi0788, n_25536);
  not g57073 (n_25537, n34549);
  and g57074 (n34550, n_14638, n_25537);
  not g57075 (n_25538, n34537);
  and g57076 (n34551, n_25538, n34550);
  not g57077 (n_25539, n34446);
  not g57078 (n_25540, n34551);
  and g57079 (n34552, n_25539, n_25540);
  not g57080 (n_25541, n34552);
  and g57081 (n34553, n_14387, n_25541);
  and g57082 (n34554, pi0630, n34436);
  and g57083 (n34555, n_14548, n_25394);
  and g57084 (n34556, n17801, n_25451);
  not g57085 (n_25542, n34554);
  not g57086 (n_25543, n34555);
  and g57087 (n34557, n_25542, n_25543);
  not g57088 (n_25544, n34556);
  and g57089 (n34558, n_25544, n34557);
  not g57090 (n_25545, n34558);
  and g57091 (n34559, pi0787, n_25545);
  not g57092 (n_25546, n34553);
  not g57093 (n_25547, n34559);
  and g57094 (n34560, n_25546, n_25547);
  and g57095 (n34561, n_11819, n34560);
  not g57096 (n_25548, n34440);
  and g57097 (n34562, n_12395, n_25548);
  not g57098 (n_25549, n34561);
  and g57099 (n34563, n_25549, n34562);
  not g57100 (n_25550, n34367);
  and g57101 (n34564, n_12405, n_25550);
  not g57102 (n_25551, n34563);
  and g57103 (n34565, n_25551, n34564);
  and g57104 (n34566, n_11819, n34439);
  and g57105 (n34567, pi0644, n34560);
  not g57106 (n_25552, n34566);
  and g57107 (n34568, pi0715, n_25552);
  not g57108 (n_25553, n34567);
  and g57109 (n34569, n_25553, n34568);
  and g57110 (n34570, pi0644, n34363);
  and g57111 (n34571, n_11819, n_25344);
  not g57112 (n_25554, n34571);
  and g57113 (n34572, n_12395, n_25554);
  not g57114 (n_25555, n34570);
  and g57115 (n34573, n_25555, n34572);
  not g57116 (n_25556, n34573);
  and g57117 (n34574, pi1160, n_25556);
  not g57118 (n_25557, n34569);
  and g57119 (n34575, n_25557, n34574);
  not g57120 (n_25558, n34565);
  not g57121 (n_25559, n34575);
  and g57122 (n34576, n_25558, n_25559);
  not g57123 (n_25560, n34576);
  and g57124 (n34577, pi0790, n_25560);
  and g57125 (n34578, n_12411, n34560);
  not g57126 (n_25561, n34577);
  not g57127 (n_25562, n34578);
  and g57128 (n34579, n_25561, n_25562);
  not g57129 (n_25563, n34579);
  and g57130 (n34580, n_4226, n_25563);
  and g57131 (n34581, n_7045, po1038);
  not g57132 (n_25564, n34580);
  not g57133 (n_25565, n34581);
  and g57134 (po0357, n_25564, n_25565);
  and g57135 (n34583, pi0233, pi0237);
  and g57136 (n34584, pi0057, pi0332);
  and g57137 (n34585, n2572, n6573);
  and g57138 (n34586, n2521, n34585);
  not g57139 (n_25568, n34586);
  and g57140 (n34587, n_4, n_25568);
  not g57141 (n_25569, n34587);
  and g57142 (n34588, n6304, n_25569);
  and g57143 (n34589, pi0332, n_3240);
  not g57144 (n_25570, n34589);
  and g57145 (n34590, pi0059, n_25570);
  not g57146 (n_25571, n34588);
  and g57147 (n34591, n_25571, n34590);
  and g57148 (n34592, pi0332, n_3243);
  not g57149 (n_25572, n34592);
  and g57150 (n34593, n_792, n_25572);
  and g57151 (n34594, pi0055, n34587);
  and g57152 (n34595, pi0074, pi0332);
  not g57153 (n_25573, n34595);
  and g57154 (n34596, n_176, n_25573);
  and g57155 (n34597, n2726, n11086);
  and g57156 (n34598, pi0468, n6192);
  and g57157 (n34599, n_234, pi0587);
  not g57158 (n_25574, n34599);
  and g57159 (n34600, n_14939, n_25574);
  not g57160 (n_25575, n34600);
  and g57161 (n34601, n_3100, n_25575);
  not g57162 (n_25576, n34598);
  not g57163 (n_25577, n34601);
  and g57164 (n34602, n_25576, n_25577);
  not g57165 (n_25578, n34602);
  and g57166 (n34603, n34597, n_25578);
  not g57167 (n_25579, n34603);
  and g57168 (n34604, n_4, n_25579);
  not g57169 (n_25580, n34604);
  and g57170 (n34605, n7363, n_25580);
  and g57171 (n34606, n2521, n6585);
  not g57172 (n_25581, n34606);
  and g57173 (n34607, n_4, n_25581);
  not g57174 (n_25582, n34607);
  and g57175 (n34608, n15625, n_25582);
  and g57176 (n34609, pi0332, n_240);
  not g57177 (n_25583, n34608);
  not g57178 (n_25584, n34609);
  and g57179 (n34610, n_25583, n_25584);
  not g57180 (n_25585, n34605);
  and g57181 (n34611, n_25585, n34610);
  not g57182 (n_25586, n34611);
  and g57183 (n34612, n_168, n_25586);
  not g57184 (n_25587, n34612);
  and g57185 (n34613, n34596, n_25587);
  not g57186 (n_25588, n34594);
  and g57187 (n34614, n2529, n_25588);
  not g57188 (n_25589, n34613);
  and g57189 (n34615, n_25589, n34614);
  not g57190 (n_25590, n34615);
  and g57191 (n34616, n34593, n_25590);
  not g57192 (n_25591, n34591);
  and g57193 (n34617, n_796, n_25591);
  not g57194 (n_25592, n34616);
  and g57195 (n34618, n_25592, n34617);
  not g57196 (n_25593, n34584);
  not g57197 (n_25594, n34618);
  and g57198 (n34619, n_25593, n_25594);
  not g57199 (n_25595, n34583);
  not g57200 (n_25596, n34619);
  and g57201 (n34620, n_25595, n_25596);
  and g57202 (n34621, n_4, n_3138);
  not g57203 (n_25597, n34621);
  and g57204 (n34622, n_3149, n_25597);
  and g57205 (n34623, pi0096, pi0210);
  and g57206 (n34624, pi0332, n34623);
  and g57207 (n34625, n_142, pi0070);
  and g57208 (n34626, n_139, n_3052);
  and g57209 (n34627, pi0032, n34626);
  not g57210 (n_25598, n34625);
  not g57211 (n_25599, n34627);
  and g57212 (n34628, n_25598, n_25599);
  not g57213 (n_25600, n34628);
  and g57214 (n34629, n_271, n_25600);
  and g57215 (n34630, n_142, n_135);
  and g57216 (n34631, pi0070, n34630);
  not g57217 (n_25601, n34631);
  and g57218 (n34632, n_4, n_25601);
  not g57219 (n_25602, n34629);
  and g57220 (n34633, n_25602, n34632);
  not g57221 (n_25603, n34624);
  not g57222 (n_25604, n34633);
  and g57223 (n34634, n_25603, n_25604);
  and g57224 (n34635, n_3102, n34634);
  not g57225 (n_25605, n34635);
  and g57226 (n34636, n6192, n_25605);
  not g57227 (n_25606, n34636);
  and g57228 (n34637, n34622, n_25606);
  not g57229 (n_25607, n34634);
  and g57230 (n34638, n6192, n_25607);
  and g57231 (n34639, pi0332, pi0468);
  and g57232 (n34640, n_3100, n_25604);
  not g57233 (n_25608, n34639);
  not g57234 (n_25609, n34640);
  and g57235 (n34641, n_25608, n_25609);
  and g57236 (n34642, n_3138, n34641);
  not g57237 (n_25610, n34638);
  and g57238 (n34643, pi0947, n_25610);
  not g57239 (n_25611, n34642);
  and g57240 (n34644, n_25611, n34643);
  not g57241 (n_25612, n34637);
  not g57242 (n_25613, n34644);
  and g57243 (n34645, n_25612, n_25613);
  not g57244 (n_25614, n34645);
  and g57245 (n34646, pi0057, n_25614);
  and g57246 (n34647, n_3240, n34645);
  and g57247 (n34648, n_204, n34645);
  not g57248 (n_25615, n34626);
  and g57249 (n34649, pi0032, n_25615);
  and g57250 (n34650, n_144, n2736);
  not g57251 (n_25616, n34649);
  and g57252 (n34651, n_25616, n34650);
  and g57253 (n34652, n2706, n34651);
  and g57254 (n34653, n2728, n34652);
  not g57255 (n_25617, n34653);
  and g57256 (n34654, n34628, n_25617);
  not g57257 (n_25618, n34654);
  and g57258 (n34655, n_271, n_25618);
  and g57259 (n34656, n_144, n2975);
  not g57260 (n_25619, n34656);
  and g57261 (n34657, n_139, n_25619);
  not g57262 (n_25620, n34657);
  and g57263 (n34658, n34630, n_25620);
  and g57264 (n34659, pi0210, n34658);
  not g57265 (n_25621, n34655);
  and g57266 (n34660, n_4, n_25621);
  not g57267 (n_25622, n34659);
  and g57268 (n34661, n_25622, n34660);
  not g57269 (n_25623, n34661);
  and g57270 (n34662, n_25603, n_25623);
  and g57271 (n34663, n_3102, n34662);
  not g57272 (n_25624, n34663);
  and g57273 (n34664, n6192, n_25624);
  not g57274 (n_25625, n34664);
  and g57275 (n34665, n34622, n_25625);
  not g57276 (n_25626, n34662);
  and g57277 (n34666, n6192, n_25626);
  and g57278 (n34667, n_3100, n_25623);
  not g57279 (n_25627, n34667);
  and g57280 (n34668, n_25608, n_25627);
  and g57281 (n34669, n_3138, n34668);
  not g57282 (n_25628, n34666);
  and g57283 (n34670, pi0947, n_25628);
  not g57284 (n_25629, n34669);
  and g57285 (n34671, n_25629, n34670);
  not g57286 (n_25630, n34665);
  not g57287 (n_25631, n34671);
  and g57288 (n34672, n_25630, n_25631);
  and g57289 (n34673, n2572, n34672);
  not g57290 (n_25632, n34648);
  not g57291 (n_25633, n34673);
  and g57292 (n34674, n_25632, n_25633);
  not g57293 (n_25634, n34674);
  and g57294 (n34675, n6304, n_25634);
  not g57295 (n_25635, n34647);
  and g57296 (n34676, pi0059, n_25635);
  not g57297 (n_25636, n34675);
  and g57298 (n34677, n_25636, n34676);
  and g57299 (n34678, n_3243, n34645);
  and g57300 (n34679, pi0055, n34674);
  and g57301 (n34680, n_168, n2611);
  and g57302 (n34681, pi0299, n_25614);
  and g57303 (n34682, pi0096, pi0198);
  and g57304 (n34683, pi0332, n34682);
  and g57305 (n34684, n_305, n_25600);
  not g57306 (n_25637, n34684);
  and g57307 (n34685, n34632, n_25637);
  not g57308 (n_25638, n34683);
  not g57309 (n_25639, n34685);
  and g57310 (n34686, n_25638, n_25639);
  not g57311 (n_25640, n34686);
  and g57312 (n34687, n6192, n_25640);
  and g57313 (n34688, n6583, n_25639);
  not g57314 (n_25641, n34688);
  and g57315 (n34689, n34621, n_25641);
  not g57321 (n_25644, n34680);
  not g57322 (n_25645, n34692);
  and g57323 (n34693, n_25644, n_25645);
  not g57324 (n_25646, n34681);
  and g57325 (n34694, n_25646, n34693);
  and g57326 (n34695, n2726, n2962);
  and g57327 (n34696, n34651, n34695);
  not g57328 (n_25647, n34696);
  and g57329 (n34697, n34628, n_25647);
  not g57330 (n_25648, n34697);
  and g57331 (n34698, n_271, n_25648);
  and g57332 (n34699, n_144, n2517);
  and g57333 (n34700, n34695, n34699);
  not g57334 (n_25649, n34700);
  and g57335 (n34701, n_139, n_25649);
  not g57336 (n_25650, n34701);
  and g57337 (n34702, n34630, n_25650);
  and g57338 (n34703, pi0210, n34702);
  not g57339 (n_25651, n34698);
  and g57340 (n34704, n_4, n_25651);
  not g57341 (n_25652, n34703);
  and g57342 (n34705, n_25652, n34704);
  not g57343 (n_25653, n34705);
  and g57344 (n34706, n_25603, n_25653);
  and g57345 (n34707, n_3102, n34706);
  not g57346 (n_25654, n34707);
  and g57347 (n34708, n6192, n_25654);
  not g57348 (n_25655, n34708);
  and g57349 (n34709, n34622, n_25655);
  not g57350 (n_25656, n34706);
  and g57351 (n34710, n6192, n_25656);
  and g57352 (n34711, n_3100, n_25653);
  not g57353 (n_25657, n34711);
  and g57354 (n34712, n_25608, n_25657);
  and g57355 (n34713, n_3138, n34712);
  not g57356 (n_25658, n34710);
  and g57357 (n34714, pi0947, n_25658);
  not g57358 (n_25659, n34713);
  and g57359 (n34715, n_25659, n34714);
  not g57360 (n_25660, n34709);
  and g57361 (n34716, pi0299, n_25660);
  not g57362 (n_25661, n34715);
  and g57363 (n34717, n_25661, n34716);
  and g57364 (n34718, n_3105, n_25597);
  and g57365 (n34719, n_305, n_25648);
  and g57366 (n34720, pi0198, n34702);
  not g57367 (n_25662, n34719);
  and g57368 (n34721, n_4, n_25662);
  not g57369 (n_25663, n34720);
  and g57370 (n34722, n_25663, n34721);
  not g57371 (n_25664, n34722);
  and g57372 (n34723, n_25638, n_25664);
  and g57373 (n34724, n_3102, n34723);
  not g57374 (n_25665, n34724);
  and g57375 (n34725, n6192, n_25665);
  not g57376 (n_25666, n34725);
  and g57377 (n34726, n34718, n_25666);
  not g57378 (n_25667, n34723);
  and g57379 (n34727, n6192, n_25667);
  and g57380 (n34728, n_3100, n_25664);
  and g57381 (n34729, n_3138, n_25608);
  not g57382 (n_25668, n34728);
  and g57383 (n34730, n_25668, n34729);
  not g57384 (n_25669, n34727);
  and g57385 (n34731, pi0587, n_25669);
  not g57386 (n_25670, n34730);
  and g57387 (n34732, n_25670, n34731);
  not g57388 (n_25671, n34726);
  and g57389 (n34733, n_234, n_25671);
  not g57390 (n_25672, n34732);
  and g57391 (n34734, n_25672, n34733);
  not g57392 (n_25673, n34717);
  not g57393 (n_25674, n34734);
  and g57394 (n34735, n_25673, n_25674);
  not g57395 (n_25675, n34735);
  and g57396 (n34736, n7363, n_25675);
  not g57397 (n_25676, n34672);
  and g57398 (n34737, pi0299, n_25676);
  and g57399 (n34738, n_305, n_25618);
  and g57400 (n34739, pi0198, n34658);
  not g57401 (n_25677, n34738);
  and g57402 (n34740, n_4, n_25677);
  not g57403 (n_25678, n34739);
  and g57404 (n34741, n_25678, n34740);
  not g57405 (n_25679, n34741);
  and g57406 (n34742, n_25638, n_25679);
  and g57407 (n34743, n_3102, n34742);
  not g57408 (n_25680, n34743);
  and g57409 (n34744, n6192, n_25680);
  not g57410 (n_25681, n34744);
  and g57411 (n34745, n34718, n_25681);
  not g57412 (n_25682, n34742);
  and g57413 (n34746, n6192, n_25682);
  and g57414 (n34747, n_3100, n_25679);
  not g57415 (n_25683, n34747);
  and g57416 (n34748, n34729, n_25683);
  not g57417 (n_25684, n34746);
  and g57418 (n34749, pi0587, n_25684);
  not g57419 (n_25685, n34748);
  and g57420 (n34750, n_25685, n34749);
  not g57421 (n_25686, n34745);
  not g57422 (n_25687, n34750);
  and g57423 (n34751, n_25686, n_25687);
  not g57424 (n_25688, n34751);
  and g57425 (n34752, n_234, n_25688);
  not g57426 (n_25689, n34737);
  and g57427 (n34753, n15625, n_25689);
  not g57428 (n_25690, n34752);
  and g57429 (n34754, n_25690, n34753);
  not g57430 (n_25691, n34736);
  not g57431 (n_25692, n34754);
  and g57432 (n34755, n_25691, n_25692);
  not g57433 (n_25693, n34755);
  and g57434 (n34756, n_168, n_25693);
  not g57435 (n_25694, n34694);
  and g57436 (n34757, n_176, n_25694);
  not g57437 (n_25695, n34756);
  and g57438 (n34758, n_25695, n34757);
  not g57439 (n_25696, n34679);
  and g57440 (n34759, n2529, n_25696);
  not g57441 (n_25697, n34758);
  and g57442 (n34760, n_25697, n34759);
  not g57443 (n_25698, n34678);
  and g57444 (n34761, n_792, n_25698);
  not g57445 (n_25699, n34760);
  and g57446 (n34762, n_25699, n34761);
  not g57447 (n_25700, n34677);
  not g57448 (n_25701, n34762);
  and g57449 (n34763, n_25700, n_25701);
  not g57450 (n_25702, n34763);
  and g57451 (n34764, n_796, n_25702);
  not g57452 (n_25703, n34646);
  not g57453 (n_25704, n34764);
  and g57454 (n34765, n_25703, n_25704);
  not g57455 (n_25705, n34765);
  and g57456 (n34766, n34583, n_25705);
  not g57457 (n_25706, n34620);
  not g57458 (n_25707, n34766);
  and g57459 (n34767, n_25706, n_25707);
  not g57460 (n_25709, pi0201);
  not g57461 (n_25710, n34767);
  and g57462 (n34768, n_25709, n_25710);
  not g57463 (n_25711, n16479);
  and g57464 (n34769, n_3445, n_25711);
  and g57465 (n34770, n6583, n34682);
  not g57466 (n_25712, n34770);
  and g57467 (n34771, n16479, n_25712);
  not g57468 (n_25713, n34623);
  and g57469 (n34772, n_25711, n_25713);
  not g57470 (n_25714, n34769);
  not g57471 (n_25715, n34771);
  and g57472 (n34773, n_25714, n_25715);
  not g57473 (n_25716, n34772);
  and g57474 (n34774, n_25716, n34773);
  and g57475 (n34775, n34583, n34774);
  not g57476 (n_25717, n34775);
  and g57477 (n34776, pi0201, n_25717);
  not g57478 (n_25718, n34768);
  not g57479 (n_25719, n34776);
  and g57480 (po0358, n_25718, n_25719);
  not g57481 (n_25720, pi0233);
  and g57482 (n34778, n_25720, pi0237);
  not g57483 (n_25721, n34778);
  and g57484 (n34779, n_25596, n_25721);
  and g57485 (n34780, n_25705, n34778);
  not g57486 (n_25722, n34779);
  not g57487 (n_25723, n34780);
  and g57488 (n34781, n_25722, n_25723);
  not g57489 (n_25725, pi0202);
  not g57490 (n_25726, n34781);
  and g57491 (n34782, n_25725, n_25726);
  and g57492 (n34783, n34774, n34778);
  not g57493 (n_25727, n34783);
  and g57494 (n34784, pi0202, n_25727);
  not g57495 (n_25728, n34782);
  not g57496 (n_25729, n34784);
  and g57497 (po0359, n_25728, n_25729);
  not g57498 (n_25730, pi0237);
  and g57499 (n34786, n_25720, n_25730);
  not g57500 (n_25731, n34786);
  and g57501 (n34787, n_25596, n_25731);
  and g57502 (n34788, n_25705, n34786);
  not g57503 (n_25732, n34787);
  not g57504 (n_25733, n34788);
  and g57505 (n34789, n_25732, n_25733);
  not g57506 (n_25735, pi0203);
  not g57507 (n_25736, n34789);
  and g57508 (n34790, n_25735, n_25736);
  and g57509 (n34791, n34774, n34786);
  not g57510 (n_25737, n34791);
  and g57511 (n34792, pi0203, n_25737);
  not g57512 (n_25738, n34790);
  not g57513 (n_25739, n34792);
  and g57514 (po0360, n_25738, n_25739);
  and g57515 (n34794, n2572, n6310);
  and g57516 (n34795, n2521, n34794);
  not g57517 (n_25740, n34795);
  and g57518 (n34796, n_4, n_25740);
  not g57519 (n_25741, n34796);
  and g57520 (n34797, n6304, n_25741);
  not g57521 (n_25742, n34797);
  and g57522 (n34798, n34590, n_25742);
  and g57523 (n34799, pi0055, n34796);
  and g57524 (n34800, n_3100, pi0602);
  and g57525 (n34801, pi0468, n6195);
  not g57526 (n_25743, n34800);
  not g57527 (n_25744, n34801);
  and g57528 (n34802, n_25743, n_25744);
  not g57529 (n_25745, n34802);
  and g57530 (n34803, n_234, n_25745);
  not g57531 (n_25746, n34803);
  and g57532 (n34804, n_3246, n_25746);
  not g57533 (n_25747, n34804);
  and g57534 (n34805, n2521, n_25747);
  not g57535 (n_25748, n34805);
  and g57536 (n34806, n_4, n_25748);
  not g57537 (n_25749, n34806);
  and g57538 (n34807, n15625, n_25749);
  and g57539 (n34808, n_234, n_3106);
  and g57540 (n34809, pi0299, n_3148);
  not g57541 (n_25750, n34808);
  and g57542 (n34810, n_3100, n_25750);
  not g57543 (n_25751, n34809);
  and g57544 (n34811, n_25751, n34810);
  not g57545 (n_25752, n34811);
  and g57546 (n34812, n_25744, n_25752);
  not g57547 (n_25753, n34812);
  and g57548 (n34813, n34597, n_25753);
  not g57549 (n_25754, n34813);
  and g57550 (n34814, n_4, n_25754);
  not g57551 (n_25755, n34814);
  and g57552 (n34815, n7363, n_25755);
  not g57553 (n_25756, n34807);
  not g57554 (n_25757, n34815);
  and g57555 (n34816, n_25756, n_25757);
  not g57556 (n_25758, n34816);
  and g57557 (n34817, n_168, n_25758);
  and g57558 (n34818, n34596, n_25584);
  not g57559 (n_25759, n34817);
  and g57560 (n34819, n_25759, n34818);
  not g57561 (n_25760, n34799);
  and g57562 (n34820, n2529, n_25760);
  not g57563 (n_25761, n34819);
  and g57564 (n34821, n_25761, n34820);
  not g57565 (n_25762, n34821);
  and g57566 (n34822, n34593, n_25762);
  not g57567 (n_25763, n34798);
  and g57568 (n34823, n_796, n_25763);
  not g57569 (n_25764, n34822);
  and g57570 (n34824, n_25764, n34823);
  not g57571 (n_25765, n34824);
  and g57572 (n34825, n_25593, n_25765);
  not g57573 (n_25766, n34825);
  and g57574 (n34826, n_25595, n_25766);
  and g57575 (n34827, n_4, n_3139);
  not g57576 (n_25767, n34827);
  and g57577 (n34828, n_3148, n_25767);
  and g57578 (n34829, n6195, n_25605);
  not g57579 (n_25768, n34829);
  and g57580 (n34830, n34828, n_25768);
  and g57581 (n34831, n6195, n_25607);
  and g57582 (n34832, n_3139, n34641);
  not g57583 (n_25769, n34831);
  and g57584 (n34833, pi0907, n_25769);
  not g57585 (n_25770, n34832);
  and g57586 (n34834, n_25770, n34833);
  not g57587 (n_25771, n34830);
  not g57588 (n_25772, n34834);
  and g57589 (n34835, n_25771, n_25772);
  not g57590 (n_25773, n34835);
  and g57591 (n34836, pi0057, n_25773);
  and g57592 (n34837, n_3240, n34835);
  and g57593 (n34838, n_204, n34835);
  and g57594 (n34839, n6195, n_25626);
  and g57595 (n34840, n_3139, n34668);
  not g57596 (n_25774, n34839);
  and g57597 (n34841, pi0907, n_25774);
  not g57598 (n_25775, n34840);
  and g57599 (n34842, n_25775, n34841);
  and g57600 (n34843, pi0332, n_11455);
  not g57601 (n_25776, n34843);
  and g57602 (n34844, pi0680, n_25776);
  and g57603 (n34845, n_25624, n34844);
  not g57604 (n_25777, n34845);
  and g57605 (n34846, n34828, n_25777);
  not g57606 (n_25778, n34842);
  not g57607 (n_25779, n34846);
  and g57608 (n34847, n_25778, n_25779);
  and g57609 (n34848, n2572, n34847);
  not g57610 (n_25780, n34838);
  not g57611 (n_25781, n34848);
  and g57612 (n34849, n_25780, n_25781);
  not g57613 (n_25782, n34849);
  and g57614 (n34850, n6304, n_25782);
  not g57615 (n_25783, n34837);
  and g57616 (n34851, pi0059, n_25783);
  not g57617 (n_25784, n34850);
  and g57618 (n34852, n_25784, n34851);
  and g57619 (n34853, n_3243, n34835);
  and g57620 (n34854, pi0055, n34849);
  and g57621 (n34855, pi0299, n34847);
  and g57622 (n34856, n6195, n34682);
  not g57623 (n_25785, n34856);
  and g57624 (n34857, pi0332, n_25785);
  not g57625 (n_25786, n34857);
  and g57626 (n34858, n_234, n_25786);
  and g57627 (n34859, n6326, n34742);
  not g57628 (n_25787, n34859);
  and g57629 (n34860, n34858, n_25787);
  not g57630 (n_25788, n34855);
  not g57631 (n_25789, n34860);
  and g57632 (n34861, n_25788, n_25789);
  not g57633 (n_25790, n34861);
  and g57634 (n34862, n15625, n_25790);
  and g57635 (n34863, n6326, n34723);
  not g57636 (n_25791, n34863);
  and g57637 (n34864, n34858, n_25791);
  and g57638 (n34865, n6195, n_25654);
  not g57639 (n_25792, n34865);
  and g57640 (n34866, n34828, n_25792);
  and g57641 (n34867, n6195, n_25656);
  and g57642 (n34868, n_3139, n34712);
  not g57643 (n_25793, n34867);
  and g57644 (n34869, pi0907, n_25793);
  not g57645 (n_25794, n34868);
  and g57646 (n34870, n_25794, n34869);
  not g57647 (n_25795, n34866);
  and g57648 (n34871, pi0299, n_25795);
  not g57649 (n_25796, n34870);
  and g57650 (n34872, n_25796, n34871);
  not g57651 (n_25797, n34864);
  not g57652 (n_25798, n34872);
  and g57653 (n34873, n_25797, n_25798);
  not g57654 (n_25799, n34873);
  and g57655 (n34874, n7363, n_25799);
  not g57656 (n_25800, n34862);
  not g57657 (n_25801, n34874);
  and g57658 (n34875, n_25800, n_25801);
  not g57659 (n_25802, n34875);
  and g57660 (n34876, n_168, n_25802);
  and g57661 (n34877, pi0299, n_25773);
  and g57662 (n34878, n34686, n_25745);
  not g57663 (n_25803, n34878);
  and g57664 (n34879, n_25786, n_25803);
  not g57665 (n_25804, n34879);
  and g57666 (n34880, n_234, n_25804);
  not g57667 (n_25805, n34880);
  and g57668 (n34881, n_25644, n_25805);
  not g57669 (n_25806, n34877);
  and g57670 (n34882, n_25806, n34881);
  not g57671 (n_25807, n34882);
  and g57672 (n34883, n_176, n_25807);
  not g57673 (n_25808, n34876);
  and g57674 (n34884, n_25808, n34883);
  not g57675 (n_25809, n34854);
  and g57676 (n34885, n2529, n_25809);
  not g57677 (n_25810, n34884);
  and g57678 (n34886, n_25810, n34885);
  not g57679 (n_25811, n34853);
  and g57680 (n34887, n_792, n_25811);
  not g57681 (n_25812, n34886);
  and g57682 (n34888, n_25812, n34887);
  not g57683 (n_25813, n34852);
  not g57684 (n_25814, n34888);
  and g57685 (n34889, n_25813, n_25814);
  not g57686 (n_25815, n34889);
  and g57687 (n34890, n_796, n_25815);
  not g57688 (n_25816, n34836);
  not g57689 (n_25817, n34890);
  and g57690 (n34891, n_25816, n_25817);
  not g57691 (n_25818, n34891);
  and g57692 (n34892, n34583, n_25818);
  not g57693 (n_25819, n34826);
  not g57694 (n_25820, n34892);
  and g57695 (n34893, n_25819, n_25820);
  not g57696 (n_25822, pi0204);
  not g57697 (n_25823, n34893);
  and g57698 (n34894, n_25822, n_25823);
  not g57699 (n_25824, n6310);
  and g57700 (n34895, n_25824, n_25711);
  and g57701 (n34896, n6326, n34682);
  not g57702 (n_25825, n34896);
  and g57703 (n34897, n16479, n_25825);
  not g57704 (n_25826, n34895);
  and g57705 (n34898, n_25716, n_25826);
  not g57706 (n_25827, n34897);
  and g57707 (n34899, n_25827, n34898);
  and g57708 (n34900, n34583, n34899);
  not g57709 (n_25828, n34900);
  and g57710 (n34901, pi0204, n_25828);
  not g57711 (n_25829, n34894);
  not g57712 (n_25830, n34901);
  and g57713 (po0361, n_25829, n_25830);
  and g57714 (n34903, n_25721, n_25766);
  and g57715 (n34904, n34778, n_25818);
  not g57716 (n_25831, n34903);
  not g57717 (n_25832, n34904);
  and g57718 (n34905, n_25831, n_25832);
  not g57719 (n_25834, pi0205);
  not g57720 (n_25835, n34905);
  and g57721 (n34906, n_25834, n_25835);
  and g57722 (n34907, n34778, n34899);
  not g57723 (n_25836, n34907);
  and g57724 (n34908, pi0205, n_25836);
  not g57725 (n_25837, n34906);
  not g57726 (n_25838, n34908);
  and g57727 (po0362, n_25837, n_25838);
  and g57728 (n34910, pi0233, n_25730);
  not g57729 (n_25839, n34910);
  and g57730 (n34911, n_25766, n_25839);
  and g57731 (n34912, n_25818, n34910);
  not g57732 (n_25840, n34911);
  not g57733 (n_25841, n34912);
  and g57734 (n34913, n_25840, n_25841);
  not g57735 (n_25843, pi0206);
  not g57736 (n_25844, n34913);
  and g57737 (n34914, n_25843, n_25844);
  and g57738 (n34915, n34899, n34910);
  not g57739 (n_25845, n34915);
  and g57740 (n34916, pi0206, n_25845);
  not g57741 (n_25846, n34914);
  not g57742 (n_25847, n34916);
  and g57743 (po0363, n_25846, n_25847);
  and g57744 (n34918, n_13449, n24385);
  and g57745 (n34919, n19151, n34918);
  and g57746 (n34920, n_13453, n34919);
  not g57747 (n_25848, n34920);
  and g57748 (n34921, pi0207, n_25848);
  and g57749 (n34922, n16635, n_11751);
  and g57750 (n34923, n2571, n24388);
  not g57751 (n_25849, n34923);
  and g57752 (n34924, n_11749, n_25849);
  and g57753 (n34925, n_11753, n_11751);
  and g57754 (n34926, pi0625, n_25849);
  not g57755 (n_25850, n34925);
  not g57756 (n_25851, n34926);
  and g57757 (n34927, n_25850, n_25851);
  not g57758 (n_25852, n34927);
  and g57759 (n34928, pi1153, n_25852);
  and g57760 (n34929, pi0625, n_11751);
  and g57761 (n34930, n_11753, n_25849);
  not g57762 (n_25853, n34929);
  not g57763 (n_25854, n34930);
  and g57764 (n34931, n_25853, n_25854);
  not g57765 (n_25855, n34931);
  and g57766 (n34932, n_11757, n_25855);
  not g57767 (n_25856, n34928);
  not g57768 (n_25857, n34932);
  and g57769 (n34933, n_25856, n_25857);
  not g57770 (n_25858, n34933);
  and g57771 (n34934, pi0778, n_25858);
  not g57772 (n_25859, n34924);
  not g57773 (n_25860, n34934);
  and g57774 (n34935, n_25859, n_25860);
  not g57775 (n_25861, n34935);
  and g57776 (n34936, n_11773, n_25861);
  and g57777 (n34937, n_11751, n17075);
  not g57778 (n_25862, n34936);
  not g57779 (n_25863, n34937);
  and g57780 (n34938, n_25862, n_25863);
  and g57781 (n34939, n_11777, n34938);
  and g57782 (n34940, n16639, n17059);
  not g57783 (n_25864, n34939);
  not g57784 (n_25865, n34940);
  and g57785 (n34941, n_25864, n_25865);
  and g57786 (n34942, n_11780, n34941);
  not g57787 (n_25866, n34922);
  not g57788 (n_25867, n34942);
  and g57789 (n34943, n_25866, n_25867);
  and g57790 (n34944, n_11783, n34943);
  and g57791 (n34945, n16631, n17059);
  not g57792 (n_25868, n34944);
  not g57793 (n_25869, n34945);
  and g57794 (n34946, n_25868, n_25869);
  not g57795 (n_25870, n34946);
  and g57796 (n34947, n_13453, n_25870);
  and g57797 (n34948, n17059, n17856);
  not g57798 (n_25871, n34947);
  not g57799 (n_25872, n34948);
  and g57800 (n34949, n_25871, n_25872);
  not g57801 (n_25873, pi0207);
  not g57802 (n_25874, n34949);
  and g57803 (n34950, n_25873, n_25874);
  not g57804 (n_25875, n34921);
  not g57805 (n_25876, n34950);
  and g57806 (n34951, n_25875, n_25876);
  not g57807 (n_25878, n34951);
  and g57808 (n34952, pi0710, n_25878);
  and g57809 (n34953, n_25873, n_11751);
  not g57810 (n_25879, pi0710);
  not g57811 (n_25880, n34953);
  and g57812 (n34954, n_25879, n_25880);
  not g57813 (n_25881, n34952);
  not g57814 (n_25882, n34954);
  and g57815 (n34955, n_25881, n_25882);
  not g57816 (n_25883, n34955);
  and g57817 (n34956, n_11803, n_25883);
  and g57818 (n34957, n_11806, n34955);
  and g57819 (n34958, pi0647, n34953);
  not g57820 (n_25884, n34958);
  and g57821 (n34959, n_11810, n_25884);
  not g57822 (n_25885, n34957);
  and g57823 (n34960, n_25885, n34959);
  and g57824 (n34961, n_11806, n34953);
  and g57825 (n34962, pi0647, n34955);
  not g57826 (n_25886, n34961);
  and g57827 (n34963, pi1157, n_25886);
  not g57828 (n_25887, n34962);
  and g57829 (n34964, n_25887, n34963);
  not g57830 (n_25888, n34960);
  not g57831 (n_25889, n34964);
  and g57832 (n34965, n_25888, n_25889);
  not g57833 (n_25890, n34965);
  and g57834 (n34966, pi0787, n_25890);
  not g57835 (n_25891, n34956);
  not g57836 (n_25892, n34966);
  and g57837 (n34967, n_25891, n_25892);
  and g57838 (n34968, n_11819, n34967);
  and g57839 (n34969, n_12375, n34964);
  and g57840 (n34970, n_11751, n17117);
  and g57841 (n34971, n2571, n19439);
  not g57842 (n_25893, n34971);
  and g57843 (n34972, n_11960, n_25893);
  not g57844 (n_25894, n34970);
  not g57845 (n_25895, n34972);
  and g57846 (n34973, n_25894, n_25895);
  not g57847 (n_25896, n34973);
  and g57848 (n34974, n_11964, n_25896);
  and g57849 (n34975, n_11751, n_11972);
  and g57850 (n34976, n_11971, n34972);
  not g57851 (n_25897, n34975);
  not g57852 (n_25898, n34976);
  and g57853 (n34977, n_25897, n_25898);
  not g57854 (n_25899, n34977);
  and g57855 (n34978, n_11768, n_25899);
  and g57856 (n34979, n_11751, n_11967);
  and g57857 (n34980, pi0609, n34972);
  not g57858 (n_25900, n34979);
  not g57859 (n_25901, n34980);
  and g57860 (n34981, n_25900, n_25901);
  not g57861 (n_25902, n34981);
  and g57862 (n34982, pi1155, n_25902);
  not g57863 (n_25903, n34978);
  not g57864 (n_25904, n34982);
  and g57865 (n34983, n_25903, n_25904);
  not g57866 (n_25905, n34983);
  and g57867 (n34984, pi0785, n_25905);
  not g57868 (n_25906, n34974);
  not g57869 (n_25907, n34984);
  and g57870 (n34985, n_25906, n_25907);
  not g57871 (n_25908, n34985);
  and g57872 (n34986, n_11981, n_25908);
  and g57873 (n34987, n_11984, n34985);
  and g57874 (n34988, pi0618, n17059);
  not g57875 (n_25909, n34988);
  and g57876 (n34989, n_11413, n_25909);
  not g57877 (n_25910, n34987);
  and g57878 (n34990, n_25910, n34989);
  and g57879 (n34991, n_11984, n17059);
  and g57880 (n34992, pi0618, n34985);
  not g57881 (n_25911, n34991);
  and g57882 (n34993, pi1154, n_25911);
  not g57883 (n_25912, n34992);
  and g57884 (n34994, n_25912, n34993);
  not g57885 (n_25913, n34990);
  not g57886 (n_25914, n34994);
  and g57887 (n34995, n_25913, n_25914);
  not g57888 (n_25915, n34995);
  and g57889 (n34996, pi0781, n_25915);
  not g57890 (n_25916, n34986);
  not g57891 (n_25917, n34996);
  and g57892 (n34997, n_25916, n_25917);
  not g57893 (n_25918, n34997);
  and g57894 (n34998, n_12315, n_25918);
  and g57895 (n34999, n_11821, n34997);
  and g57896 (n35000, pi0619, n17059);
  not g57897 (n_25919, n35000);
  and g57898 (n35001, n_11405, n_25919);
  not g57899 (n_25920, n34999);
  and g57900 (n35002, n_25920, n35001);
  and g57901 (n35003, n_11821, n17059);
  and g57902 (n35004, pi0619, n34997);
  not g57903 (n_25921, n35003);
  and g57904 (n35005, pi1159, n_25921);
  not g57905 (n_25922, n35004);
  and g57906 (n35006, n_25922, n35005);
  not g57907 (n_25923, n35002);
  not g57908 (n_25924, n35006);
  and g57909 (n35007, n_25923, n_25924);
  not g57910 (n_25925, n35007);
  and g57911 (n35008, pi0789, n_25925);
  not g57912 (n_25926, n34998);
  not g57913 (n_25927, n35008);
  and g57914 (n35009, n_25926, n_25927);
  and g57915 (n35010, n_12524, n35009);
  and g57916 (n35011, n17059, n17969);
  not g57917 (n_25928, n35010);
  not g57918 (n_25929, n35011);
  and g57919 (n35012, n_25928, n_25929);
  not g57920 (n_25930, n35012);
  and g57921 (n35013, n_12368, n_25930);
  and g57922 (n35014, n17059, n17779);
  not g57923 (n_25931, n35013);
  not g57924 (n_25932, n35014);
  and g57925 (n35015, n_25931, n_25932);
  not g57926 (n_25933, n35015);
  and g57927 (n35016, n_25873, n_25933);
  and g57928 (n35017, n2571, n_17784);
  and g57929 (n35018, n_11960, n35017);
  and g57930 (n35019, n_14288, n35018);
  and g57931 (n35020, n_14295, n35019);
  and g57932 (n35021, n_14294, n35020);
  and g57933 (n35022, n_12524, n35021);
  and g57934 (n35023, n_12368, n35022);
  not g57935 (n_25934, n35023);
  and g57936 (n35024, pi0207, n_25934);
  not g57937 (n_25936, n35024);
  and g57938 (n35025, pi0623, n_25936);
  not g57939 (n_25937, n35016);
  and g57940 (n35026, n_25937, n35025);
  not g57941 (n_25938, pi0623);
  and g57942 (n35027, n_25938, n34953);
  not g57943 (n_25939, n35026);
  not g57944 (n_25940, n35027);
  and g57945 (n35028, n_25939, n_25940);
  and g57946 (n35029, n_14548, n35028);
  and g57947 (n35030, pi0630, n34960);
  not g57948 (n_25941, n34969);
  not g57949 (n_25942, n35029);
  and g57950 (n35031, n_25941, n_25942);
  not g57951 (n_25943, n35030);
  and g57952 (n35032, n_25943, n35031);
  not g57953 (n_25944, n35032);
  and g57954 (n35033, pi0787, n_25944);
  not g57955 (n_25945, n35028);
  and g57956 (n35034, n_25879, n_25945);
  and g57957 (n35035, n_11789, n_11751);
  and g57958 (n35036, pi0628, n34946);
  not g57959 (n_25946, n35035);
  not g57960 (n_25947, n35036);
  and g57961 (n35037, n_25946, n_25947);
  not g57962 (n_25948, n35037);
  and g57963 (n35038, n_12354, n_25948);
  not g57964 (n_25949, n35038);
  and g57965 (n35039, n_25946, n_25949);
  not g57966 (n_25950, n35039);
  and g57967 (n35040, pi1156, n_25950);
  and g57968 (n35041, pi0628, n_11751);
  and g57969 (n35042, n_11794, n35041);
  and g57970 (n35043, n_11789, n34946);
  not g57971 (n_25951, n35041);
  not g57972 (n_25952, n35043);
  and g57973 (n35044, n_25951, n_25952);
  not g57974 (n_25953, n35044);
  and g57975 (n35045, n17777, n_25953);
  not g57976 (n_25954, n35042);
  not g57977 (n_25955, n35045);
  and g57978 (n35046, n_25954, n_25955);
  not g57979 (n_25956, n35040);
  and g57980 (n35047, n_25956, n35046);
  not g57981 (n_25957, n35047);
  and g57982 (n35048, pi0792, n_25957);
  and g57983 (n35049, pi1159, n_11751);
  and g57984 (n35050, pi0619, n34941);
  and g57985 (n35051, pi1154, n_11751);
  not g57986 (n_25958, n34938);
  and g57987 (n35052, pi0618, n_25958);
  and g57988 (n35053, pi1155, n_11751);
  and g57989 (n35054, pi0609, n_25861);
  not g57990 (n_25959, n19477);
  and g57991 (n35055, n2571, n_25959);
  not g57992 (n_25960, n35055);
  and g57993 (n35056, n_11749, n_25960);
  and g57994 (n35057, n_11753, n_25960);
  not g57995 (n_25961, n35057);
  and g57996 (n35058, n_25853, n_25961);
  not g57997 (n_25962, n35058);
  and g57998 (n35059, n_11757, n_25962);
  and g57999 (n35060, n_11823, n_25856);
  not g58000 (n_25963, n35059);
  and g58001 (n35061, n_25963, n35060);
  and g58002 (n35062, pi0625, n_25960);
  not g58003 (n_25964, n35062);
  and g58004 (n35063, n_25850, n_25964);
  not g58005 (n_25965, n35063);
  and g58006 (n35064, pi1153, n_25965);
  and g58007 (n35065, pi0608, n_25857);
  not g58008 (n_25966, n35064);
  and g58009 (n35066, n_25966, n35065);
  not g58010 (n_25967, n35061);
  and g58011 (n35067, pi0778, n_25967);
  not g58012 (n_25968, n35066);
  and g58013 (n35068, n_25968, n35067);
  not g58014 (n_25969, n35056);
  not g58015 (n_25970, n35068);
  and g58016 (n35069, n_25969, n_25970);
  not g58017 (n_25971, n35069);
  and g58018 (n35070, n_11971, n_25971);
  not g58019 (n_25972, n35054);
  not g58020 (n_25973, n35070);
  and g58021 (n35071, n_25972, n_25973);
  not g58022 (n_25974, n35071);
  and g58023 (n35072, n_11768, n_25974);
  not g58024 (n_25975, n35053);
  and g58025 (n35073, n_11767, n_25975);
  not g58026 (n_25976, n35072);
  and g58027 (n35074, n_25976, n35073);
  and g58028 (n35075, n_11768, n_11751);
  and g58029 (n35076, n_11971, n_25861);
  and g58030 (n35077, pi0609, n_25971);
  not g58031 (n_25977, n35076);
  not g58032 (n_25978, n35077);
  and g58033 (n35078, n_25977, n_25978);
  not g58034 (n_25979, n35078);
  and g58035 (n35079, pi1155, n_25979);
  not g58036 (n_25980, n35075);
  and g58037 (n35080, pi0660, n_25980);
  not g58038 (n_25981, n35079);
  and g58039 (n35081, n_25981, n35080);
  not g58040 (n_25982, n35074);
  not g58041 (n_25983, n35081);
  and g58042 (n35082, n_25982, n_25983);
  not g58043 (n_25984, n35082);
  and g58044 (n35083, pi0785, n_25984);
  and g58045 (n35084, n_11964, n35069);
  not g58046 (n_25985, n35083);
  not g58047 (n_25986, n35084);
  and g58048 (n35085, n_25985, n_25986);
  and g58049 (n35086, n_11984, n35085);
  not g58050 (n_25987, n35052);
  not g58051 (n_25988, n35086);
  and g58052 (n35087, n_25987, n_25988);
  not g58053 (n_25989, n35087);
  and g58054 (n35088, n_11413, n_25989);
  not g58055 (n_25990, n35051);
  and g58056 (n35089, n_11412, n_25990);
  not g58057 (n_25991, n35088);
  and g58058 (n35090, n_25991, n35089);
  and g58059 (n35091, n_11413, n_11751);
  and g58060 (n35092, n_11984, n_25958);
  and g58061 (n35093, pi0618, n35085);
  not g58062 (n_25992, n35092);
  not g58063 (n_25993, n35093);
  and g58064 (n35094, n_25992, n_25993);
  not g58065 (n_25994, n35094);
  and g58066 (n35095, pi1154, n_25994);
  not g58067 (n_25995, n35091);
  and g58068 (n35096, pi0627, n_25995);
  not g58069 (n_25996, n35095);
  and g58070 (n35097, n_25996, n35096);
  not g58071 (n_25997, n35090);
  not g58072 (n_25998, n35097);
  and g58073 (n35098, n_25997, n_25998);
  not g58074 (n_25999, n35098);
  and g58075 (n35099, pi0781, n_25999);
  not g58076 (n_26000, n35085);
  and g58077 (n35100, n_11981, n_26000);
  not g58078 (n_26001, n35099);
  not g58079 (n_26002, n35100);
  and g58080 (n35101, n_26001, n_26002);
  and g58081 (n35102, n_11821, n35101);
  not g58082 (n_26003, n35050);
  not g58083 (n_26004, n35102);
  and g58084 (n35103, n_26003, n_26004);
  not g58085 (n_26005, n35103);
  and g58086 (n35104, n_11405, n_26005);
  not g58087 (n_26006, n35049);
  and g58088 (n35105, n_11403, n_26006);
  not g58089 (n_26007, n35104);
  and g58090 (n35106, n_26007, n35105);
  and g58091 (n35107, n_11405, n_11751);
  and g58092 (n35108, n_11821, n34941);
  and g58093 (n35109, pi0619, n35101);
  not g58094 (n_26008, n35108);
  not g58095 (n_26009, n35109);
  and g58096 (n35110, n_26008, n_26009);
  not g58097 (n_26010, n35110);
  and g58098 (n35111, pi1159, n_26010);
  not g58099 (n_26011, n35107);
  and g58100 (n35112, pi0648, n_26011);
  not g58101 (n_26012, n35111);
  and g58102 (n35113, n_26012, n35112);
  not g58103 (n_26013, n35106);
  not g58104 (n_26014, n35113);
  and g58105 (n35114, n_26013, n_26014);
  not g58106 (n_26015, n35114);
  and g58107 (n35115, pi0789, n_26015);
  not g58108 (n_26016, n35101);
  and g58109 (n35116, n_12315, n_26016);
  not g58110 (n_26017, n35115);
  not g58111 (n_26018, n35116);
  and g58112 (n35117, n_26017, n_26018);
  not g58113 (n_26019, n35117);
  and g58114 (n35118, n_12318, n_26019);
  and g58115 (n35119, pi0641, n_11751);
  and g58116 (n35120, pi0626, n34943);
  and g58117 (n35121, n_12320, n_26019);
  not g58118 (n_26020, n35120);
  and g58119 (n35122, n_11395, n_26020);
  not g58120 (n_26021, n35121);
  and g58121 (n35123, n_26021, n35122);
  not g58122 (n_26022, n35119);
  and g58123 (n35124, n_11397, n_26022);
  not g58124 (n_26023, n35123);
  and g58125 (n35125, n_26023, n35124);
  and g58126 (n35126, n_11395, n_11751);
  and g58127 (n35127, n_12320, n34943);
  and g58128 (n35128, pi0626, n_26019);
  not g58129 (n_26024, n35127);
  and g58130 (n35129, pi0641, n_26024);
  not g58131 (n_26025, n35128);
  and g58132 (n35130, n_26025, n35129);
  not g58133 (n_26026, n35126);
  and g58134 (n35131, pi1158, n_26026);
  not g58135 (n_26027, n35130);
  and g58136 (n35132, n_26027, n35131);
  not g58137 (n_26028, n35125);
  not g58138 (n_26029, n35132);
  and g58139 (n35133, n_26028, n_26029);
  not g58140 (n_26030, n35133);
  and g58141 (n35134, pi0788, n_26030);
  not g58142 (n_26031, n35118);
  and g58143 (n35135, n_14638, n_26031);
  not g58144 (n_26032, n35134);
  and g58145 (n35136, n_26032, n35135);
  not g58146 (n_26033, n35048);
  not g58147 (n_26034, n35136);
  and g58148 (n35137, n_26033, n_26034);
  not g58149 (n_26035, n35137);
  and g58150 (n35138, n_25873, n_26035);
  not g58151 (n_26036, n34918);
  and g58152 (n35139, pi0609, n_26036);
  and g58153 (n35140, n_11749, n_25173);
  and g58154 (n35141, n_11753, n34080);
  not g58155 (n_26037, n35141);
  and g58156 (n35142, n_11757, n_26037);
  and g58157 (n35143, pi0625, n24385);
  not g58158 (n_26038, n35143);
  and g58159 (n35144, pi1153, n_26038);
  not g58160 (n_26039, n35144);
  and g58161 (n35145, n_11823, n_26039);
  not g58162 (n_26040, n35142);
  and g58163 (n35146, n_26040, n35145);
  and g58164 (n35147, pi0625, n34080);
  not g58165 (n_26041, n35147);
  and g58166 (n35148, pi1153, n_26041);
  and g58167 (n35149, n_11753, n24385);
  not g58168 (n_26042, n35149);
  and g58169 (n35150, n_11757, n_26042);
  not g58170 (n_26043, n35150);
  and g58171 (n35151, pi0608, n_26043);
  not g58172 (n_26044, n35148);
  and g58173 (n35152, n_26044, n35151);
  not g58174 (n_26045, n35146);
  and g58175 (n35153, pi0778, n_26045);
  not g58176 (n_26046, n35152);
  and g58177 (n35154, n_26046, n35153);
  not g58178 (n_26047, n35140);
  not g58179 (n_26048, n35154);
  and g58180 (n35155, n_26047, n_26048);
  not g58181 (n_26049, n35155);
  and g58182 (n35156, n_11971, n_26049);
  not g58183 (n_26050, n35139);
  and g58184 (n35157, n17073, n_26050);
  not g58185 (n_26051, n35156);
  and g58186 (n35158, n_26051, n35157);
  and g58187 (n35159, pi0609, n_26049);
  and g58188 (n35160, n_11971, n_26036);
  not g58189 (n_26052, n35160);
  and g58190 (n35161, n17072, n_26052);
  not g58191 (n_26053, n35159);
  and g58192 (n35162, n_26053, n35161);
  not g58193 (n_26054, n35158);
  not g58194 (n_26055, n35162);
  and g58195 (n35163, n_26054, n_26055);
  not g58196 (n_26056, n35163);
  and g58197 (n35164, pi0785, n_26056);
  and g58198 (n35165, n_11964, n35155);
  not g58199 (n_26057, n35164);
  not g58200 (n_26058, n35165);
  and g58201 (n35166, n_26057, n_26058);
  and g58202 (n35167, n_11981, n35166);
  and g58203 (n35168, n_11984, n35166);
  and g58204 (n35169, n_11773, n34918);
  not g58205 (n_26059, n35169);
  and g58206 (n35170, pi0618, n_26059);
  not g58207 (n_26060, n35170);
  and g58208 (n35171, n16637, n_26060);
  not g58209 (n_26061, n35168);
  and g58210 (n35172, n_26061, n35171);
  and g58211 (n35173, n_11984, n_26059);
  and g58212 (n35174, pi0618, n35166);
  not g58213 (n_26062, n35173);
  and g58214 (n35175, n16636, n_26062);
  not g58215 (n_26063, n35174);
  and g58216 (n35176, n_26063, n35175);
  not g58217 (n_26064, n35172);
  and g58218 (n35177, pi0781, n_26064);
  not g58219 (n_26065, n35176);
  and g58220 (n35178, n_26065, n35177);
  not g58221 (n_26066, n35167);
  and g58222 (n35179, n_16916, n_26066);
  not g58223 (n_26067, n35178);
  and g58224 (n35180, n_26067, n35179);
  and g58225 (n35181, n19150, n34918);
  and g58226 (n35182, n16634, n20231);
  and g58227 (n35183, n35181, n35182);
  not g58228 (n_26068, n35180);
  not g58229 (n_26069, n35183);
  and g58230 (n35184, n_26068, n_26069);
  and g58231 (n35185, n_12318, n35184);
  and g58232 (n35186, n_11780, n35181);
  not g58233 (n_26070, n35186);
  and g58234 (n35187, pi0626, n_26070);
  not g58235 (n_26071, n35187);
  and g58236 (n35188, n_11395, n_26071);
  and g58237 (n35189, n_12320, n35184);
  and g58238 (n35190, n_11397, n35188);
  not g58239 (n_26072, n35189);
  and g58240 (n35191, n_26072, n35190);
  and g58241 (n35192, pi0626, n35184);
  and g58242 (n35193, n_12320, n_26070);
  not g58243 (n_26073, n35193);
  and g58244 (n35194, pi0641, n_26073);
  and g58245 (n35195, pi1158, n35194);
  not g58246 (n_26074, n35192);
  and g58247 (n35196, n_26074, n35195);
  not g58248 (n_26075, n35191);
  and g58249 (n35197, pi0788, n_26075);
  not g58250 (n_26076, n35196);
  and g58251 (n35198, n_26076, n35197);
  not g58252 (n_26077, n35185);
  and g58253 (n35199, n_14638, n_26077);
  not g58254 (n_26078, n35198);
  and g58255 (n35200, n_26078, n35199);
  and g58256 (n35201, n17779, n17855);
  and g58257 (n35202, n34919, n35201);
  not g58258 (n_26079, n35200);
  not g58259 (n_26080, n35202);
  and g58260 (n35203, n_26079, n_26080);
  not g58261 (n_26081, n35203);
  and g58262 (n35204, pi0207, n_26081);
  not g58263 (n_26082, n35204);
  and g58264 (n35205, n_25938, n_26082);
  not g58265 (n_26083, n35138);
  and g58266 (n35206, n_26083, n35205);
  not g58267 (n_26084, n34919);
  and g58268 (n35207, n_11794, n_26084);
  not g58269 (n_26085, n35022);
  and g58270 (n35208, pi1156, n_26085);
  not g58271 (n_26086, n35207);
  and g58272 (n35209, n20566, n_26086);
  not g58273 (n_26087, n35208);
  and g58274 (n35210, n_26087, n35209);
  and g58275 (n35211, pi1156, n_26084);
  and g58276 (n35212, n_11794, n_26085);
  not g58277 (n_26088, n35211);
  and g58278 (n35213, n20568, n_26088);
  not g58279 (n_26089, n35212);
  and g58280 (n35214, n_26089, n35213);
  not g58281 (n_26090, n35210);
  not g58282 (n_26091, n35214);
  and g58283 (n35215, n_26090, n_26091);
  not g58284 (n_26092, n35215);
  and g58285 (n35216, pi0792, n_26092);
  and g58286 (n35217, n17868, n35021);
  not g58287 (n_26093, n35020);
  and g58288 (n35218, n_11405, n_26093);
  not g58289 (n_26094, n35181);
  and g58290 (n35219, pi1159, n_26094);
  and g58296 (n35223, pi1159, n_26093);
  and g58297 (n35224, n_11405, n_26094);
  not g58303 (n_26099, n35222);
  and g58304 (n35228, pi0789, n_26099);
  not g58305 (n_26100, n35227);
  and g58306 (n35229, n_26100, n35228);
  not g58307 (n_26101, n35229);
  and g58308 (n35230, pi0789, n_26101);
  and g58309 (n35231, n_11413, n_26060);
  and g58310 (n35232, n20233, n35019);
  not g58311 (n_26102, n35232);
  and g58312 (n35233, n_11412, n_26102);
  not g58313 (n_26103, n35231);
  and g58314 (n35234, n_26103, n35233);
  and g58315 (n35235, n20232, n35019);
  and g58316 (n35236, n_11749, n_25176);
  and g58317 (n35237, n_11753, n34085);
  and g58318 (n35238, pi0625, n35017);
  not g58319 (n_26104, n35238);
  and g58320 (n35239, n_11757, n_26104);
  not g58321 (n_26105, n35237);
  and g58322 (n35240, n_26105, n35239);
  not g58323 (n_26106, n35240);
  and g58324 (n35241, n35145, n_26106);
  and g58325 (n35242, n_11753, n35017);
  and g58326 (n35243, pi0625, n34085);
  not g58327 (n_26107, n35242);
  and g58328 (n35244, pi1153, n_26107);
  not g58329 (n_26108, n35243);
  and g58330 (n35245, n_26108, n35244);
  not g58331 (n_26109, n35245);
  and g58332 (n35246, n35151, n_26109);
  not g58333 (n_26110, n35241);
  and g58334 (n35247, pi0778, n_26110);
  not g58335 (n_26111, n35246);
  and g58336 (n35248, n_26111, n35247);
  not g58337 (n_26112, n35236);
  not g58338 (n_26113, n35248);
  and g58339 (n35249, n_26112, n_26113);
  not g58340 (n_26114, n35249);
  and g58341 (n35250, n_11964, n_26114);
  and g58342 (n35251, n20223, n35018);
  and g58343 (n35252, n_11971, n_26114);
  and g58344 (n35253, n_11768, n_26050);
  not g58345 (n_26115, n35252);
  and g58346 (n35254, n_26115, n35253);
  not g58347 (n_26116, n35251);
  and g58348 (n35255, n_11767, n_26116);
  not g58349 (n_26117, n35254);
  and g58350 (n35256, n_26117, n35255);
  and g58351 (n35257, n20222, n35018);
  and g58352 (n35258, pi0609, n_26114);
  and g58353 (n35259, pi1155, n_26052);
  not g58354 (n_26118, n35258);
  and g58355 (n35260, n_26118, n35259);
  not g58356 (n_26119, n35257);
  and g58357 (n35261, pi0660, n_26119);
  not g58358 (n_26120, n35260);
  and g58359 (n35262, n_26120, n35261);
  not g58360 (n_26121, n35256);
  not g58361 (n_26122, n35262);
  and g58362 (n35263, n_26121, n_26122);
  not g58363 (n_26123, n35263);
  and g58364 (n35264, pi0785, n_26123);
  not g58365 (n_26124, n35250);
  not g58366 (n_26125, n35264);
  and g58367 (n35265, n_26124, n_26125);
  not g58368 (n_26126, n35265);
  and g58369 (n35266, pi0618, n_26126);
  and g58370 (n35267, pi1154, n_26062);
  not g58371 (n_26127, n35266);
  and g58372 (n35268, n_26127, n35267);
  not g58373 (n_26128, n35235);
  and g58374 (n35269, pi0627, n_26128);
  not g58375 (n_26129, n35268);
  and g58376 (n35270, n_26129, n35269);
  not g58377 (n_26130, n35234);
  not g58378 (n_26131, n35270);
  and g58379 (n35271, n_26130, n_26131);
  not g58380 (n_26132, n35271);
  and g58381 (n35272, pi0781, n_26132);
  and g58382 (n35273, n_11984, n_11412);
  not g58383 (n_26133, n35273);
  and g58384 (n35274, pi0781, n_26133);
  not g58385 (n_26134, n35274);
  and g58386 (n35275, n_26126, n_26134);
  and g58387 (n35276, n_16914, n35229);
  not g58388 (n_26135, n35275);
  not g58389 (n_26136, n35276);
  and g58390 (n35277, n_26135, n_26136);
  not g58391 (n_26137, n35272);
  and g58392 (n35278, n_26137, n35277);
  not g58393 (n_26138, n35230);
  not g58394 (n_26139, n35278);
  and g58395 (n35279, n_26138, n_26139);
  and g58396 (n35280, n_12320, n35279);
  not g58397 (n_26140, n35280);
  and g58398 (n35281, n35188, n_26140);
  not g58399 (n_26141, n35217);
  and g58400 (n35282, n_11397, n_26141);
  not g58401 (n_26142, n35281);
  and g58402 (n35283, n_26142, n35282);
  and g58403 (n35284, n17869, n35021);
  and g58404 (n35285, pi0626, n35279);
  not g58405 (n_26143, n35285);
  and g58406 (n35286, n35194, n_26143);
  not g58407 (n_26144, n35284);
  and g58408 (n35287, pi1158, n_26144);
  not g58409 (n_26145, n35286);
  and g58410 (n35288, n_26145, n35287);
  not g58411 (n_26146, n35283);
  not g58412 (n_26147, n35288);
  and g58413 (n35289, n_26146, n_26147);
  not g58414 (n_26148, n35289);
  and g58415 (n35290, pi0788, n_26148);
  and g58416 (n35291, n_12318, n35279);
  not g58417 (n_26149, n35291);
  and g58418 (n35292, n_14638, n_26149);
  not g58419 (n_26150, n35290);
  and g58420 (n35293, n_26150, n35292);
  not g58421 (n_26151, n35216);
  not g58422 (n_26152, n35293);
  and g58423 (n35294, n_26151, n_26152);
  not g58424 (n_26153, n35294);
  and g58425 (n35295, pi0207, n_26153);
  and g58426 (n35296, n2571, n19488);
  not g58427 (n_26154, n35296);
  and g58428 (n35297, n_11749, n_26154);
  and g58429 (n35298, n_11753, n34971);
  and g58430 (n35299, pi0625, n35296);
  not g58431 (n_26155, n35299);
  and g58432 (n35300, pi1153, n_26155);
  not g58433 (n_26156, n35298);
  and g58434 (n35301, n_26156, n35300);
  not g58435 (n_26157, n35301);
  and g58436 (n35302, n35065, n_26157);
  and g58437 (n35303, n_11753, n35296);
  and g58438 (n35304, pi0625, n34971);
  not g58439 (n_26158, n35303);
  and g58440 (n35305, n_11757, n_26158);
  not g58441 (n_26159, n35304);
  and g58442 (n35306, n_26159, n35305);
  not g58443 (n_26160, n35306);
  and g58444 (n35307, n35060, n_26160);
  not g58445 (n_26161, n35302);
  and g58446 (n35308, pi0778, n_26161);
  not g58447 (n_26162, n35307);
  and g58448 (n35309, n_26162, n35308);
  not g58449 (n_26163, n35297);
  not g58450 (n_26164, n35309);
  and g58451 (n35310, n_26163, n_26164);
  not g58452 (n_26165, n35310);
  and g58453 (n35311, n_11971, n_26165);
  not g58454 (n_26166, n35311);
  and g58455 (n35312, n_25972, n_26166);
  not g58456 (n_26167, n35312);
  and g58457 (n35313, n_11768, n_26167);
  and g58458 (n35314, n_11767, n_25904);
  not g58459 (n_26168, n35313);
  and g58460 (n35315, n_26168, n35314);
  and g58461 (n35316, pi0609, n_26165);
  not g58462 (n_26169, n35316);
  and g58463 (n35317, n_25977, n_26169);
  not g58464 (n_26170, n35317);
  and g58465 (n35318, pi1155, n_26170);
  and g58466 (n35319, pi0660, n_25903);
  not g58467 (n_26171, n35318);
  and g58468 (n35320, n_26171, n35319);
  not g58469 (n_26172, n35315);
  not g58470 (n_26173, n35320);
  and g58471 (n35321, n_26172, n_26173);
  not g58472 (n_26174, n35321);
  and g58473 (n35322, pi0785, n_26174);
  and g58474 (n35323, n_11964, n35310);
  not g58475 (n_26175, n35322);
  not g58476 (n_26176, n35323);
  and g58477 (n35324, n_26175, n_26176);
  and g58478 (n35325, n_11984, n35324);
  not g58479 (n_26177, n35325);
  and g58480 (n35326, n_25987, n_26177);
  not g58481 (n_26178, n35326);
  and g58482 (n35327, n_11413, n_26178);
  and g58483 (n35328, n_11412, n_25914);
  not g58484 (n_26179, n35327);
  and g58485 (n35329, n_26179, n35328);
  and g58486 (n35330, pi0618, n35324);
  not g58487 (n_26180, n35330);
  and g58488 (n35331, n_25992, n_26180);
  not g58489 (n_26181, n35331);
  and g58490 (n35332, pi1154, n_26181);
  and g58491 (n35333, pi0627, n_25913);
  not g58492 (n_26182, n35332);
  and g58493 (n35334, n_26182, n35333);
  not g58494 (n_26183, n35329);
  not g58495 (n_26184, n35334);
  and g58496 (n35335, n_26183, n_26184);
  not g58497 (n_26185, n35335);
  and g58498 (n35336, pi0781, n_26185);
  not g58499 (n_26186, n35324);
  and g58500 (n35337, n_11981, n_26186);
  not g58501 (n_26187, n35336);
  not g58502 (n_26188, n35337);
  and g58503 (n35338, n_26187, n_26188);
  and g58504 (n35339, n_12315, n35338);
  and g58505 (n35340, n_11821, n35338);
  not g58506 (n_26189, n35340);
  and g58507 (n35341, n_26003, n_26189);
  not g58508 (n_26190, n35341);
  and g58509 (n35342, n_11405, n_26190);
  and g58510 (n35343, n_11403, n_25924);
  not g58511 (n_26191, n35342);
  and g58512 (n35344, n_26191, n35343);
  and g58513 (n35345, pi0619, n35338);
  not g58514 (n_26192, n35345);
  and g58515 (n35346, n_26008, n_26192);
  not g58516 (n_26193, n35346);
  and g58517 (n35347, pi1159, n_26193);
  and g58518 (n35348, pi0648, n_25923);
  not g58519 (n_26194, n35347);
  and g58520 (n35349, n_26194, n35348);
  not g58521 (n_26195, n35344);
  and g58522 (n35350, pi0789, n_26195);
  not g58523 (n_26196, n35349);
  and g58524 (n35351, n_26196, n35350);
  not g58525 (n_26197, n35339);
  and g58526 (n35352, n17970, n_26197);
  not g58527 (n_26198, n35351);
  and g58528 (n35353, n_26198, n35352);
  not g58529 (n_26199, n34943);
  and g58530 (n35354, pi0641, n_26199);
  and g58531 (n35355, n17865, n_26026);
  not g58532 (n_26200, n35354);
  and g58533 (n35356, n_26200, n35355);
  and g58534 (n35357, n_11401, n_12446);
  and g58535 (n35358, n35009, n35357);
  and g58536 (n35359, n_11395, n_26199);
  and g58537 (n35360, n17866, n_26022);
  not g58538 (n_26201, n35359);
  and g58539 (n35361, n_26201, n35360);
  not g58540 (n_26202, n35356);
  not g58541 (n_26203, n35361);
  and g58542 (n35362, n_26202, n_26203);
  not g58543 (n_26204, n35358);
  and g58544 (n35363, n_26204, n35362);
  not g58545 (n_26205, n35363);
  and g58546 (n35364, pi0788, n_26205);
  not g58547 (n_26206, n35364);
  and g58548 (n35365, n_14638, n_26206);
  not g58549 (n_26207, n35353);
  and g58550 (n35366, n_26207, n35365);
  and g58551 (n35367, n_14557, n35012);
  and g58552 (n35368, pi1156, n35038);
  not g58553 (n_26208, n35367);
  and g58554 (n35369, n_25955, n_26208);
  not g58555 (n_26209, n35368);
  and g58556 (n35370, n_26209, n35369);
  not g58557 (n_26210, n35370);
  and g58558 (n35371, pi0792, n_26210);
  not g58559 (n_26211, n35366);
  not g58560 (n_26212, n35371);
  and g58561 (n35372, n_26211, n_26212);
  not g58562 (n_26213, n35372);
  and g58563 (n35373, n_25873, n_26213);
  not g58564 (n_26214, n35295);
  and g58565 (n35374, pi0623, n_26214);
  not g58566 (n_26215, n35373);
  and g58567 (n35375, n_26215, n35374);
  not g58568 (n_26216, n35375);
  and g58569 (n35376, pi0710, n_26216);
  not g58570 (n_26217, n35206);
  and g58571 (n35377, n_26217, n35376);
  not g58572 (n_26218, n35034);
  and g58573 (n35378, n_14387, n_26218);
  not g58574 (n_26219, n35377);
  and g58575 (n35379, n_26219, n35378);
  not g58576 (n_26220, n35033);
  not g58577 (n_26221, n35379);
  and g58578 (n35380, n_26220, n_26221);
  and g58579 (n35381, pi0644, n35380);
  not g58580 (n_26222, n34968);
  and g58581 (n35382, pi0715, n_26222);
  not g58582 (n_26223, n35381);
  and g58583 (n35383, n_26223, n35382);
  and g58584 (n35384, n17804, n_25880);
  and g58585 (n35385, n_12392, n35028);
  not g58586 (n_26224, n35384);
  not g58587 (n_26225, n35385);
  and g58588 (n35386, n_26224, n_26225);
  and g58589 (n35387, pi0644, n35386);
  and g58590 (n35388, n_11819, n34953);
  not g58591 (n_26226, n35388);
  and g58592 (n35389, n_12395, n_26226);
  not g58593 (n_26227, n35387);
  and g58594 (n35390, n_26227, n35389);
  not g58595 (n_26228, n35390);
  and g58596 (n35391, pi1160, n_26228);
  not g58597 (n_26229, n35383);
  and g58598 (n35392, n_26229, n35391);
  and g58599 (n35393, pi0644, n34967);
  and g58600 (n35394, n_11819, n35380);
  not g58601 (n_26230, n35393);
  and g58602 (n35395, n_12395, n_26230);
  not g58603 (n_26231, n35394);
  and g58604 (n35396, n_26231, n35395);
  and g58605 (n35397, n_11819, n35386);
  and g58606 (n35398, pi0644, n34953);
  not g58607 (n_26232, n35398);
  and g58608 (n35399, pi0715, n_26232);
  not g58609 (n_26233, n35397);
  and g58610 (n35400, n_26233, n35399);
  not g58611 (n_26234, n35400);
  and g58612 (n35401, n_12405, n_26234);
  not g58613 (n_26235, n35396);
  and g58614 (n35402, n_26235, n35401);
  not g58615 (n_26236, n35392);
  not g58616 (n_26237, n35402);
  and g58617 (n35403, n_26236, n_26237);
  not g58618 (n_26238, n35403);
  and g58619 (n35404, pi0790, n_26238);
  and g58620 (n35405, n_12411, n35380);
  not g58621 (n_26239, n35404);
  not g58622 (n_26240, n35405);
  and g58623 (n35406, n_26239, n_26240);
  not g58624 (n_26241, n35406);
  and g58625 (n35407, n_4226, n_26241);
  and g58626 (n35408, n_25873, po1038);
  or g58627 (po0364, n35407, n35408);
  and g58628 (n35410, pi0208, n_25848);
  not g58629 (n_26242, pi0208);
  and g58630 (n35411, n_26242, n_25874);
  not g58631 (n_26243, n35410);
  not g58632 (n_26244, n35411);
  and g58633 (n35412, n_26243, n_26244);
  not g58634 (n_26246, n35412);
  and g58635 (n35413, pi0638, n_26246);
  and g58636 (n35414, n_26242, n_11751);
  not g58637 (n_26247, pi0638);
  not g58638 (n_26248, n35414);
  and g58639 (n35415, n_26247, n_26248);
  not g58640 (n_26249, n35413);
  not g58641 (n_26250, n35415);
  and g58642 (n35416, n_26249, n_26250);
  not g58643 (n_26251, n35416);
  and g58644 (n35417, n_11803, n_26251);
  and g58645 (n35418, n_11806, n35416);
  and g58646 (n35419, pi0647, n35414);
  not g58647 (n_26252, n35419);
  and g58648 (n35420, n_11810, n_26252);
  not g58649 (n_26253, n35418);
  and g58650 (n35421, n_26253, n35420);
  and g58651 (n35422, n_11806, n35414);
  and g58652 (n35423, pi0647, n35416);
  not g58653 (n_26254, n35422);
  and g58654 (n35424, pi1157, n_26254);
  not g58655 (n_26255, n35423);
  and g58656 (n35425, n_26255, n35424);
  not g58657 (n_26256, n35421);
  not g58658 (n_26257, n35425);
  and g58659 (n35426, n_26256, n_26257);
  not g58660 (n_26258, n35426);
  and g58661 (n35427, pi0787, n_26258);
  not g58662 (n_26259, n35417);
  not g58663 (n_26260, n35427);
  and g58664 (n35428, n_26259, n_26260);
  and g58665 (n35429, n_11819, n35428);
  and g58666 (n35430, n_12375, n35425);
  and g58667 (n35431, n_26242, n_25933);
  and g58668 (n35432, pi0208, n_25934);
  not g58669 (n_26262, n35432);
  and g58670 (n35433, pi0607, n_26262);
  not g58671 (n_26263, n35431);
  and g58672 (n35434, n_26263, n35433);
  not g58673 (n_26264, pi0607);
  and g58674 (n35435, n_26264, n35414);
  not g58675 (n_26265, n35434);
  not g58676 (n_26266, n35435);
  and g58677 (n35436, n_26265, n_26266);
  and g58678 (n35437, n_14548, n35436);
  and g58679 (n35438, pi0630, n35421);
  not g58680 (n_26267, n35430);
  not g58681 (n_26268, n35437);
  and g58682 (n35439, n_26267, n_26268);
  not g58683 (n_26269, n35438);
  and g58684 (n35440, n_26269, n35439);
  not g58685 (n_26270, n35440);
  and g58686 (n35441, pi0787, n_26270);
  not g58687 (n_26271, n35436);
  and g58688 (n35442, n_26247, n_26271);
  and g58689 (n35443, n_26242, n_26035);
  and g58690 (n35444, pi0208, n_26081);
  not g58691 (n_26272, n35444);
  and g58692 (n35445, n_26264, n_26272);
  not g58693 (n_26273, n35443);
  and g58694 (n35446, n_26273, n35445);
  and g58695 (n35447, pi0208, n_26153);
  and g58696 (n35448, n_26242, n_26213);
  not g58697 (n_26274, n35447);
  and g58698 (n35449, pi0607, n_26274);
  not g58699 (n_26275, n35448);
  and g58700 (n35450, n_26275, n35449);
  not g58701 (n_26276, n35450);
  and g58702 (n35451, pi0638, n_26276);
  not g58703 (n_26277, n35446);
  and g58704 (n35452, n_26277, n35451);
  not g58705 (n_26278, n35442);
  and g58706 (n35453, n_14387, n_26278);
  not g58707 (n_26279, n35452);
  and g58708 (n35454, n_26279, n35453);
  not g58709 (n_26280, n35441);
  not g58710 (n_26281, n35454);
  and g58711 (n35455, n_26280, n_26281);
  and g58712 (n35456, pi0644, n35455);
  not g58713 (n_26282, n35429);
  and g58714 (n35457, pi0715, n_26282);
  not g58715 (n_26283, n35456);
  and g58716 (n35458, n_26283, n35457);
  and g58717 (n35459, n17804, n_26248);
  and g58718 (n35460, n_12392, n35436);
  not g58719 (n_26284, n35459);
  not g58720 (n_26285, n35460);
  and g58721 (n35461, n_26284, n_26285);
  and g58722 (n35462, pi0644, n35461);
  and g58723 (n35463, n_11819, n35414);
  not g58724 (n_26286, n35463);
  and g58725 (n35464, n_12395, n_26286);
  not g58726 (n_26287, n35462);
  and g58727 (n35465, n_26287, n35464);
  not g58728 (n_26288, n35465);
  and g58729 (n35466, pi1160, n_26288);
  not g58730 (n_26289, n35458);
  and g58731 (n35467, n_26289, n35466);
  and g58732 (n35468, pi0644, n35428);
  and g58733 (n35469, n_11819, n35455);
  not g58734 (n_26290, n35468);
  and g58735 (n35470, n_12395, n_26290);
  not g58736 (n_26291, n35469);
  and g58737 (n35471, n_26291, n35470);
  and g58738 (n35472, n_11819, n35461);
  and g58739 (n35473, pi0644, n35414);
  not g58740 (n_26292, n35473);
  and g58741 (n35474, pi0715, n_26292);
  not g58742 (n_26293, n35472);
  and g58743 (n35475, n_26293, n35474);
  not g58744 (n_26294, n35475);
  and g58745 (n35476, n_12405, n_26294);
  not g58746 (n_26295, n35471);
  and g58747 (n35477, n_26295, n35476);
  not g58748 (n_26296, n35467);
  not g58749 (n_26297, n35477);
  and g58750 (n35478, n_26296, n_26297);
  not g58751 (n_26298, n35478);
  and g58752 (n35479, pi0790, n_26298);
  and g58753 (n35480, n_12411, n35455);
  not g58754 (n_26299, n35479);
  not g58755 (n_26300, n35480);
  and g58756 (n35481, n_26299, n_26300);
  not g58757 (n_26301, n35481);
  and g58758 (n35482, n_4226, n_26301);
  and g58759 (n35483, n_26242, po1038);
  or g58760 (po0365, n35482, n35483);
  and g58761 (n35485, n10197, n17052);
  not g58762 (n_26303, pi0639);
  and g58763 (n35486, n_26303, n35485);
  and g58764 (n35487, pi0715, n17059);
  and g58765 (n35488, n_14387, n_26035);
  and g58766 (n35489, n_11806, n_11751);
  and g58767 (n35490, pi0647, n34949);
  not g58768 (n_26304, n35489);
  not g58769 (n_26305, n35490);
  and g58770 (n35491, n_26304, n_26305);
  not g58771 (n_26306, n35491);
  and g58772 (n35492, n_12375, n_26306);
  not g58773 (n_26307, n35492);
  and g58774 (n35493, n_26304, n_26307);
  not g58775 (n_26308, n35493);
  and g58776 (n35494, pi1157, n_26308);
  and g58777 (n35495, pi0647, n_11751);
  and g58778 (n35496, n_11810, n35495);
  and g58779 (n35497, n_11806, n34949);
  not g58780 (n_26309, n35495);
  not g58781 (n_26310, n35497);
  and g58782 (n35498, n_26309, n_26310);
  not g58783 (n_26311, n35498);
  and g58784 (n35499, n17802, n_26311);
  not g58785 (n_26312, n35496);
  not g58786 (n_26313, n35499);
  and g58787 (n35500, n_26312, n_26313);
  not g58788 (n_26314, n35494);
  and g58789 (n35501, n_26314, n35500);
  not g58790 (n_26315, n35501);
  and g58791 (n35502, pi0787, n_26315);
  not g58792 (n_26316, n35488);
  not g58793 (n_26317, n35502);
  and g58794 (n35503, n_26316, n_26317);
  not g58795 (n_26318, n35503);
  and g58796 (n35504, n_11819, n_26318);
  and g58797 (n35505, n_13598, n34949);
  and g58798 (n35506, n_11751, n19342);
  not g58799 (n_26319, n35505);
  not g58800 (n_26320, n35506);
  and g58801 (n35507, n_26319, n_26320);
  not g58802 (n_26321, n35507);
  and g58803 (n35508, pi0644, n_26321);
  not g58804 (n_26322, n35508);
  and g58805 (n35509, n_12395, n_26322);
  not g58806 (n_26323, n35504);
  and g58807 (n35510, n_26323, n35509);
  not g58808 (n_26324, n35487);
  and g58809 (n35511, n_12405, n_26324);
  not g58810 (n_26325, n35510);
  and g58811 (n35512, n_26325, n35511);
  and g58812 (n35513, n_12395, n17059);
  and g58813 (n35514, pi0644, n_26318);
  and g58814 (n35515, n_11819, n_26321);
  not g58815 (n_26326, n35515);
  and g58816 (n35516, pi0715, n_26326);
  not g58817 (n_26327, n35514);
  and g58818 (n35517, n_26327, n35516);
  not g58819 (n_26328, n35513);
  and g58820 (n35518, pi1160, n_26328);
  not g58821 (n_26329, n35517);
  and g58822 (n35519, n_26329, n35518);
  not g58823 (n_26330, n35512);
  not g58824 (n_26331, n35519);
  and g58825 (n35520, n_26330, n_26331);
  not g58826 (n_26332, n35520);
  and g58827 (n35521, pi0790, n_26332);
  and g58828 (n35522, n_12411, n_26318);
  not g58829 (n_26333, n35522);
  and g58830 (n35523, n_4226, n_26333);
  not g58831 (n_26334, n35521);
  and g58832 (n35524, n_26334, n35523);
  and g58833 (n35525, pi0639, n35524);
  not g58834 (n_26336, pi0622);
  not g58835 (n_26337, n35486);
  and g58836 (n35526, n_26336, n_26337);
  not g58837 (n_26338, n35525);
  and g58838 (n35527, n_26338, n35526);
  and g58839 (n35528, n_11751, n17804);
  and g58840 (n35529, n_12392, n35015);
  not g58841 (n_26339, n35528);
  not g58842 (n_26340, n35529);
  and g58843 (n35530, n_26339, n_26340);
  not g58844 (n_26341, n35530);
  and g58845 (n35531, n_12411, n_26341);
  and g58846 (n35532, pi0644, n_26341);
  and g58847 (n35533, n_11819, n_11751);
  not g58848 (n_26342, n35532);
  not g58849 (n_26343, n35533);
  and g58850 (n35534, n_26342, n_26343);
  and g58851 (n35535, pi1160, n35534);
  and g58852 (n35536, n_11819, n_26341);
  and g58853 (n35537, pi0644, n_11751);
  not g58854 (n_26344, n35536);
  not g58855 (n_26345, n35537);
  and g58856 (n35538, n_26344, n_26345);
  and g58857 (n35539, n_12405, n35538);
  not g58858 (n_26346, n35535);
  and g58859 (n35540, pi0790, n_26346);
  not g58860 (n_26347, n35539);
  and g58861 (n35541, n_26347, n35540);
  not g58862 (n_26348, n35531);
  and g58863 (n35542, n_4226, n_26348);
  not g58864 (n_26349, n35541);
  and g58865 (n35543, n_26349, n35542);
  and g58866 (n35544, n_26303, n35543);
  and g58867 (n35545, pi0715, n35538);
  and g58868 (n35546, n_14387, n_26213);
  and g58869 (n35547, n_14548, n35015);
  and g58870 (n35548, pi1157, n35492);
  not g58871 (n_26350, n35547);
  and g58872 (n35549, n_26313, n_26350);
  not g58873 (n_26351, n35548);
  and g58874 (n35550, n_26351, n35549);
  not g58875 (n_26352, n35550);
  and g58876 (n35551, pi0787, n_26352);
  not g58877 (n_26353, n35546);
  not g58878 (n_26354, n35551);
  and g58879 (n35552, n_26353, n_26354);
  not g58880 (n_26355, n35552);
  and g58881 (n35553, n_11819, n_26355);
  not g58882 (n_26356, n35553);
  and g58883 (n35554, n35509, n_26356);
  not g58884 (n_26357, n35545);
  and g58885 (n35555, n_12405, n_26357);
  not g58886 (n_26358, n35554);
  and g58887 (n35556, n_26358, n35555);
  and g58888 (n35557, n_12395, n35534);
  and g58889 (n35558, pi0644, n_26355);
  not g58890 (n_26359, n35558);
  and g58891 (n35559, n35516, n_26359);
  not g58892 (n_26360, n35557);
  and g58893 (n35560, pi1160, n_26360);
  not g58894 (n_26361, n35559);
  and g58895 (n35561, n_26361, n35560);
  not g58896 (n_26362, n35556);
  not g58897 (n_26363, n35561);
  and g58898 (n35562, n_26362, n_26363);
  not g58899 (n_26364, n35562);
  and g58900 (n35563, pi0790, n_26364);
  and g58901 (n35564, n_12411, n_26355);
  not g58902 (n_26365, n35564);
  and g58903 (n35565, n_4226, n_26365);
  not g58904 (n_26366, n35563);
  and g58905 (n35566, n_26366, n35565);
  and g58906 (n35567, pi0639, n35566);
  not g58907 (n_26367, n35544);
  and g58908 (n35568, pi0622, n_26367);
  not g58909 (n_26368, n35567);
  and g58910 (n35569, n_26368, n35568);
  not g58911 (n_26369, n35527);
  not g58912 (n_26370, n35569);
  and g58913 (n35570, n_26369, n_26370);
  not g58914 (n_26372, pi0209);
  not g58915 (n_26373, n35570);
  and g58916 (n35571, n_26372, n_26373);
  and g58917 (n35572, n_11819, pi1160);
  and g58918 (n35573, pi0644, n_12405);
  not g58919 (n_26374, n35572);
  not g58920 (n_26375, n35573);
  and g58921 (n35574, n_26374, n_26375);
  not g58922 (n_26376, n35574);
  and g58923 (n35575, pi0790, n_26376);
  and g58924 (n35576, n23684, n35022);
  not g58925 (n_26377, n35575);
  and g58926 (n35577, n_4226, n_26377);
  and g58927 (n35578, n35576, n35577);
  and g58928 (n35579, pi0622, n35578);
  not g58929 (n_26378, n35579);
  and g58930 (n35580, n_26303, n_26378);
  and g58931 (n35581, n_14387, n_26081);
  and g58932 (n35582, n17804, n19341);
  and g58933 (n35583, n34920, n35582);
  not g58934 (n_26379, n35581);
  not g58935 (n_26380, n35583);
  and g58936 (n35584, n_26379, n_26380);
  and g58937 (n35585, n_12411, n35584);
  and g58938 (n35586, n_13598, n34920);
  not g58939 (n_26381, n35586);
  and g58940 (n35587, n_11819, n_26381);
  not g58941 (n_26382, n35587);
  and g58942 (n35588, pi0715, n_26382);
  and g58943 (n35589, pi0644, n35584);
  and g58944 (n35590, pi1160, n35588);
  not g58945 (n_26383, n35589);
  and g58946 (n35591, n_26383, n35590);
  and g58947 (n35592, pi0644, n_26381);
  not g58948 (n_26384, n35592);
  and g58949 (n35593, n_12395, n_26384);
  and g58950 (n35594, n_11819, n35584);
  and g58951 (n35595, n_12405, n35593);
  not g58952 (n_26385, n35594);
  and g58953 (n35596, n_26385, n35595);
  not g58954 (n_26386, n35591);
  and g58955 (n35597, pi0790, n_26386);
  not g58956 (n_26387, n35596);
  and g58957 (n35598, n_26387, n35597);
  not g58958 (n_26388, n35585);
  and g58959 (n35599, n_4226, n_26388);
  not g58960 (n_26389, n35598);
  and g58961 (n35600, n_26389, n35599);
  not g58962 (n_26390, n35600);
  and g58963 (n35601, n_26336, n_26390);
  and g58964 (n35602, n_11819, pi0715);
  and g58965 (n35603, n35576, n35602);
  and g58966 (n35604, pi0647, n34920);
  not g58967 (n_26391, n35604);
  and g58968 (n35605, pi1157, n_26391);
  and g58969 (n35606, pi0647, n35023);
  and g58970 (n35607, n_11806, n_26153);
  not g58971 (n_26392, n35606);
  and g58972 (n35608, n_11810, n_26392);
  not g58973 (n_26393, n35607);
  and g58974 (n35609, n_26393, n35608);
  not g58975 (n_26394, n35605);
  and g58976 (n35610, n_12375, n_26394);
  not g58977 (n_26395, n35609);
  and g58978 (n35611, n_26395, n35610);
  and g58979 (n35612, n_11806, n34920);
  not g58980 (n_26396, n35612);
  and g58981 (n35613, n_11810, n_26396);
  and g58982 (n35614, n_11806, n35023);
  and g58983 (n35615, pi0647, n_26153);
  not g58984 (n_26397, n35614);
  and g58985 (n35616, pi1157, n_26397);
  not g58986 (n_26398, n35615);
  and g58987 (n35617, n_26398, n35616);
  not g58988 (n_26399, n35613);
  and g58989 (n35618, pi0630, n_26399);
  not g58990 (n_26400, n35617);
  and g58991 (n35619, n_26400, n35618);
  not g58992 (n_26401, n35611);
  not g58993 (n_26402, n35619);
  and g58994 (n35620, n_26401, n_26402);
  not g58995 (n_26403, n35620);
  and g58996 (n35621, pi0787, n_26403);
  and g58997 (n35622, n_11803, n_26153);
  not g58998 (n_26404, n35621);
  not g58999 (n_26405, n35622);
  and g59000 (n35623, n_26404, n_26405);
  and g59001 (n35624, n_11819, n35623);
  not g59002 (n_26406, n35624);
  and g59003 (n35625, n35593, n_26406);
  not g59004 (n_26407, n35603);
  and g59005 (n35626, n_12405, n_26407);
  not g59006 (n_26408, n35625);
  and g59007 (n35627, n_26408, n35626);
  and g59008 (n35628, pi0644, n_12395);
  and g59009 (n35629, n35576, n35628);
  and g59010 (n35630, pi0644, n35623);
  not g59011 (n_26409, n35630);
  and g59012 (n35631, n35588, n_26409);
  not g59013 (n_26410, n35629);
  and g59014 (n35632, pi1160, n_26410);
  not g59015 (n_26411, n35631);
  and g59016 (n35633, n_26411, n35632);
  not g59017 (n_26412, n35627);
  not g59018 (n_26413, n35633);
  and g59019 (n35634, n_26412, n_26413);
  not g59020 (n_26414, n35634);
  and g59021 (n35635, pi0790, n_26414);
  and g59022 (n35636, n_12411, n35623);
  not g59023 (n_26415, n35636);
  and g59024 (n35637, n_4226, n_26415);
  not g59025 (n_26416, n35635);
  and g59026 (n35638, n_26416, n35637);
  and g59027 (n35639, pi0622, pi0639);
  not g59028 (n_26417, n35638);
  and g59029 (n35640, n_26417, n35639);
  or g59036 (po0366, n35571, n35643);
  and g59037 (n35645, pi0210, n_11418);
  and g59038 (n35646, pi0634, n20902);
  and g59039 (n35647, pi0633, pi0947);
  not g59040 (n_26421, n35646);
  not g59041 (n_26422, n35647);
  and g59042 (n35648, n_26421, n_26422);
  not g59043 (n_26423, n35648);
  and g59044 (n35649, n16641, n_26423);
  not g59045 (n_26424, n35645);
  and g59046 (n35650, pi0038, n_26424);
  not g59047 (n_26425, n35649);
  and g59048 (n35651, n_26425, n35650);
  and g59049 (n35652, n_11651, n_26423);
  not g59050 (n_26426, n35652);
  and g59051 (n35653, pi0299, n_26426);
  and g59052 (n35654, n_11652, n35653);
  and g59053 (n35655, pi0210, n_11671);
  and g59054 (n35656, n16930, n_26423);
  not g59055 (n_26427, n35655);
  and g59056 (n35657, n_234, n_26427);
  not g59057 (n_26428, n35656);
  and g59058 (n35658, n_26428, n35657);
  not g59059 (n_26429, n35654);
  and g59060 (n35659, n_162, n_26429);
  not g59061 (n_26430, n35658);
  and g59062 (n35660, n_26430, n35659);
  and g59063 (n35661, pi0210, n_11445);
  not g59064 (n_26431, n33589);
  not g59065 (n_26432, n35661);
  and g59066 (n35662, n_26431, n_26432);
  and g59067 (n35663, n6227, n35662);
  not g59068 (n_26433, n35663);
  and g59069 (n35664, pi0947, n_26433);
  and g59070 (n35665, pi0210, n16721);
  and g59071 (n35666, pi0633, n_11479);
  not g59072 (n_26434, n35665);
  not g59073 (n_26435, n35666);
  and g59074 (n35667, n_26434, n_26435);
  and g59075 (n35668, n_3140, n35667);
  not g59076 (n_26436, n35668);
  and g59077 (n35669, n35664, n_26436);
  and g59078 (n35670, pi0634, n16653);
  not g59079 (n_26437, n35670);
  and g59080 (n35671, n_26432, n_26437);
  and g59081 (n35672, n6227, n35671);
  not g59082 (n_26438, n35672);
  and g59083 (n35673, pi0907, n_26438);
  not g59084 (n_26439, n33430);
  and g59085 (n35674, n_26439, n_26434);
  and g59086 (n35675, n_3140, n35674);
  not g59087 (n_26440, n35675);
  and g59088 (n35676, n35673, n_26440);
  and g59089 (n35677, n6227, n16652);
  and g59090 (n35678, n2926, n35677);
  not g59091 (n_26441, n35678);
  and g59092 (n35679, n35665, n_26441);
  not g59093 (n_26442, n35676);
  not g59094 (n_26443, n35679);
  and g59095 (n35680, n_26442, n_26443);
  not g59096 (n_26444, n35680);
  and g59097 (n35681, n_3149, n_26444);
  not g59098 (n_26445, n35669);
  and g59099 (n35682, n_3119, n_26445);
  not g59100 (n_26446, n35681);
  and g59101 (n35683, n_26446, n35682);
  and g59102 (n35684, n_24622, n35662);
  not g59103 (n_26447, n35684);
  and g59104 (n35685, pi0947, n_26447);
  not g59105 (n_26448, n35667);
  and g59106 (n35686, n_3102, n_26448);
  and g59107 (n35687, po1101, n35662);
  not g59108 (n_26449, n35687);
  and g59109 (n35688, n_3120, n_26449);
  not g59110 (n_26450, n35686);
  not g59111 (n_26451, n35688);
  and g59112 (n35689, n_26450, n_26451);
  not g59113 (n_26452, n35689);
  and g59114 (n35690, n35685, n_26452);
  not g59115 (n_26453, n35671);
  and g59116 (n35691, n_3120, n_26453);
  not g59117 (n_26454, n35691);
  and g59118 (n35692, pi0907, n_26454);
  not g59119 (n_26455, n35674);
  and g59120 (n35693, n6198, n_26455);
  not g59121 (n_26456, n35693);
  and g59122 (n35694, n35692, n_26456);
  and g59123 (n35695, n_24622, n35661);
  and g59124 (n35696, pi0210, po1101);
  and g59125 (n35697, n_11543, n35696);
  not g59126 (n_26457, n35695);
  not g59127 (n_26458, n35697);
  and g59128 (n35698, n_26457, n_26458);
  and g59129 (n35699, n_3148, n35698);
  not g59130 (n_26459, n35694);
  and g59131 (n35700, n_3149, n_26459);
  not g59132 (n_26460, n35699);
  and g59133 (n35701, n_26460, n35700);
  not g59134 (n_26461, n35690);
  and g59135 (n35702, n6205, n_26461);
  not g59136 (n_26462, n35701);
  and g59137 (n35703, n_26462, n35702);
  not g59138 (n_26463, n35683);
  and g59139 (n35704, pi0223, n_26463);
  not g59140 (n_26464, n35703);
  and g59141 (n35705, n_26464, n35704);
  and g59142 (n35706, n16653, n_26423);
  not g59143 (n_26465, n35706);
  and g59144 (n35707, n_26432, n_26465);
  and g59145 (n35708, n2603, n35707);
  and g59146 (n35709, pi0210, n16681);
  and g59147 (n35710, pi0633, n_11448);
  not g59148 (n_26466, n35709);
  not g59149 (n_26467, n35710);
  and g59150 (n35711, n_26466, n_26467);
  not g59151 (n_26468, n35711);
  and g59152 (n35712, n_3102, n_26468);
  not g59153 (n_26469, n35712);
  and g59154 (n35713, n_26451, n_26469);
  not g59155 (n_26470, n35713);
  and g59156 (n35714, n35685, n_26470);
  and g59157 (n35715, pi0634, n_11448);
  not g59158 (n_26471, n35715);
  and g59159 (n35716, n_26466, n_26471);
  not g59160 (n_26472, n35716);
  and g59161 (n35717, n6198, n_26472);
  not g59162 (n_26473, n35717);
  and g59163 (n35718, n35692, n_26473);
  and g59164 (n35719, n_11513, n35696);
  not g59165 (n_26474, n35719);
  and g59166 (n35720, n_26457, n_26474);
  and g59167 (n35721, n_3148, n35720);
  not g59168 (n_26475, n35718);
  and g59169 (n35722, n_3149, n_26475);
  not g59170 (n_26476, n35721);
  and g59171 (n35723, n_26476, n35722);
  not g59172 (n_26477, n35714);
  and g59173 (n35724, n6205, n_26477);
  not g59174 (n_26478, n35723);
  and g59175 (n35725, n_26478, n35724);
  and g59176 (n35726, n_3140, n35716);
  not g59177 (n_26479, n35726);
  and g59178 (n35727, n35673, n_26479);
  and g59179 (n35728, pi0210, n_24632);
  and g59180 (n35729, n_3148, n35728);
  not g59181 (n_26480, n35727);
  not g59182 (n_26481, n35729);
  and g59183 (n35730, n_26480, n_26481);
  not g59184 (n_26482, n35730);
  and g59185 (n35731, n_3149, n_26482);
  and g59186 (n35732, n_3140, n35711);
  not g59187 (n_26483, n35732);
  and g59188 (n35733, n35664, n_26483);
  not g59189 (n_26484, n35733);
  and g59190 (n35734, n_3119, n_26484);
  not g59191 (n_26485, n35731);
  and g59192 (n35735, n_26485, n35734);
  not g59193 (n_26486, n35725);
  not g59194 (n_26487, n35735);
  and g59195 (n35736, n_26486, n_26487);
  not g59196 (n_26488, n35736);
  and g59197 (n35737, n_9349, n_26488);
  not g59198 (n_26489, n35708);
  and g59199 (n35738, n_223, n_26489);
  not g59200 (n_26490, n35737);
  and g59201 (n35739, n_26490, n35738);
  not g59202 (n_26491, n35705);
  and g59203 (n35740, n_234, n_26491);
  not g59204 (n_26492, n35739);
  and g59205 (n35741, n_26492, n35740);
  and g59206 (n35742, n_11720, n_26443);
  and g59207 (n35743, n6241, n35698);
  not g59208 (n_26493, n35742);
  and g59209 (n35744, n_3148, n_26493);
  not g59210 (n_26494, n35743);
  and g59211 (n35745, n_26494, n35744);
  not g59212 (n_26495, n35745);
  and g59213 (n35746, n_26442, n_26495);
  not g59214 (n_26496, n35746);
  and g59215 (n35747, n_3149, n_26496);
  not g59216 (n_26497, n35747);
  and g59217 (n35748, n_26445, n_26497);
  not g59218 (n_26498, n35748);
  and g59219 (n35749, pi0215, n_26498);
  and g59220 (n35750, n3448, n35707);
  not g59221 (n_26499, n35728);
  and g59222 (n35751, n_11720, n_26499);
  and g59223 (n35752, n6241, n35720);
  not g59224 (n_26500, n35752);
  and g59225 (n35753, n_3148, n_26500);
  not g59226 (n_26501, n35751);
  and g59227 (n35754, n_26501, n35753);
  not g59228 (n_26502, n35754);
  and g59229 (n35755, n_26480, n_26502);
  not g59230 (n_26503, n35755);
  and g59231 (n35756, n_3149, n_26503);
  and g59232 (n35757, n_9350, n_26484);
  not g59233 (n_26504, n35756);
  and g59234 (n35758, n_26504, n35757);
  not g59235 (n_26505, n35750);
  and g59236 (n35759, n_36, n_26505);
  not g59237 (n_26506, n35758);
  and g59238 (n35760, n_26506, n35759);
  not g59239 (n_26507, n35749);
  and g59240 (n35761, pi0299, n_26507);
  not g59241 (n_26508, n35760);
  and g59242 (n35762, n_26508, n35761);
  not g59243 (n_26509, n35762);
  and g59244 (n35763, pi0039, n_26509);
  not g59245 (n_26510, n35741);
  and g59246 (n35764, n_26510, n35763);
  not g59247 (n_26511, n35660);
  and g59248 (n35765, n_161, n_26511);
  not g59249 (n_26512, n35764);
  and g59250 (n35766, n_26512, n35765);
  not g59251 (n_26513, n35651);
  not g59252 (n_26514, n35766);
  and g59253 (n35767, n_26513, n_26514);
  not g59254 (n_26515, n35767);
  and g59255 (n35768, n10197, n_26515);
  and g59256 (n35769, n_271, n_14814);
  not g59257 (n_26516, n35768);
  not g59258 (n_26517, n35769);
  and g59259 (po0367, n_26516, n_26517);
  and g59260 (n35771, n2571, n_15421);
  and g59261 (n35772, n_25343, n35771);
  and g59262 (n35773, n2571, n_15420);
  and g59263 (n35774, pi0606, n35773);
  not g59264 (n_26518, n35772);
  and g59265 (n35775, pi0643, n_26518);
  not g59266 (n_26519, n35774);
  and g59267 (n35776, n_26519, n35775);
  and g59268 (n35777, n_25343, n17059);
  and g59269 (n35778, n2571, n_15424);
  and g59270 (n35779, pi0606, n35778);
  not g59271 (n_26520, n35777);
  and g59272 (n35780, n_25400, n_26520);
  not g59273 (n_26521, n35779);
  and g59274 (n35781, n_26521, n35780);
  not g59275 (n_26522, n35781);
  and g59276 (n35782, n_4226, n_26522);
  not g59277 (n_26523, n35776);
  and g59278 (n35783, n_26523, n35782);
  not g59279 (n_26524, n35783);
  and g59280 (n35784, pi0211, n_26524);
  and g59281 (n35785, n2571, n21628);
  not g59282 (n_26525, n35785);
  and g59283 (n35786, n_25343, n_26525);
  and g59284 (n35787, n2571, n21625);
  not g59285 (n_26526, n35787);
  and g59286 (n35788, pi0606, n_26526);
  not g59287 (n_26527, n35786);
  and g59288 (n35789, pi0643, n_26527);
  not g59289 (n_26528, n35788);
  and g59290 (n35790, n_26528, n35789);
  and g59291 (n35791, n2571, n21034);
  and g59292 (n35792, pi0606, n_25400);
  and g59293 (n35793, n35791, n35792);
  not g59294 (n_26529, n35790);
  not g59295 (n_26530, n35793);
  and g59296 (n35794, n_26529, n_26530);
  and g59297 (n35795, n_7075, n_4226);
  not g59298 (n_26531, n35794);
  and g59299 (n35796, n_26531, n35795);
  or g59300 (po0368, n35784, n35796);
  and g59301 (n35798, n_26264, n35771);
  and g59302 (n35799, pi0607, n35773);
  not g59303 (n_26532, n35798);
  and g59304 (n35800, pi0638, n_26532);
  not g59305 (n_26533, n35799);
  and g59306 (n35801, n_26533, n35800);
  and g59307 (n35802, n_26264, n17059);
  and g59308 (n35803, pi0607, n35778);
  not g59309 (n_26534, n35802);
  and g59310 (n35804, n_26247, n_26534);
  not g59311 (n_26535, n35803);
  and g59312 (n35805, n_26535, n35804);
  not g59313 (n_26536, n35805);
  and g59314 (n35806, n_4226, n_26536);
  not g59315 (n_26537, n35801);
  and g59316 (n35807, n_26537, n35806);
  not g59317 (n_26538, pi0212);
  not g59318 (n_26539, n35807);
  and g59319 (n35808, n_26538, n_26539);
  and g59320 (n35809, pi0607, n_26526);
  and g59321 (n35810, n_26264, n_26525);
  not g59322 (n_26540, n35809);
  and g59323 (n35811, pi0638, n_26540);
  not g59324 (n_26541, n35810);
  and g59325 (n35812, n_26541, n35811);
  and g59326 (n35813, pi0607, n_26247);
  and g59327 (n35814, n35791, n35813);
  not g59328 (n_26542, n35812);
  not g59329 (n_26543, n35814);
  and g59330 (n35815, n_26542, n_26543);
  and g59331 (n35816, pi0212, n_4226);
  not g59332 (n_26544, n35815);
  and g59333 (n35817, n_26544, n35816);
  or g59334 (po0369, n35808, n35817);
  and g59335 (n35819, pi0213, n_4226);
  and g59336 (n35820, pi0622, n_26526);
  and g59337 (n35821, n_26336, n_26525);
  not g59338 (n_26546, n35820);
  and g59339 (n35822, pi0639, n_26546);
  not g59340 (n_26547, n35821);
  and g59341 (n35823, n_26547, n35822);
  and g59342 (n35824, pi0622, n_26303);
  and g59343 (n35825, n35791, n35824);
  not g59344 (n_26548, n35823);
  not g59345 (n_26549, n35825);
  and g59346 (n35826, n_26548, n_26549);
  not g59347 (n_26550, n35826);
  and g59348 (n35827, n35819, n_26550);
  and g59349 (n35828, n_26303, n35778);
  and g59350 (n35829, pi0639, n35773);
  not g59351 (n_26551, n35828);
  and g59352 (n35830, pi0622, n_26551);
  not g59353 (n_26552, n35829);
  and g59354 (n35831, n_26552, n35830);
  and g59355 (n35832, n_26303, n17059);
  and g59356 (n35833, pi0639, n35771);
  not g59357 (n_26553, n35832);
  and g59358 (n35834, n_26336, n_26553);
  not g59359 (n_26554, n35833);
  and g59360 (n35835, n_26554, n35834);
  not g59361 (n_26555, n35835);
  and g59362 (n35836, n_4226, n_26555);
  not g59363 (n_26556, n35831);
  and g59364 (n35837, n_26556, n35836);
  not g59365 (n_26557, pi0213);
  not g59366 (n_26558, n35837);
  and g59367 (n35838, n_26557, n_26558);
  or g59368 (po0370, n35827, n35838);
  and g59369 (n35840, n_25938, n35771);
  and g59370 (n35841, pi0623, n35773);
  not g59371 (n_26559, n35840);
  and g59372 (n35842, pi0710, n_26559);
  not g59373 (n_26560, n35841);
  and g59374 (n35843, n_26560, n35842);
  and g59375 (n35844, n_25938, n17059);
  and g59376 (n35845, pi0623, n35778);
  not g59377 (n_26561, n35844);
  and g59378 (n35846, n_25879, n_26561);
  not g59379 (n_26562, n35845);
  and g59380 (n35847, n_26562, n35846);
  not g59381 (n_26563, n35847);
  and g59382 (n35848, n_4226, n_26563);
  not g59383 (n_26564, n35843);
  and g59384 (n35849, n_26564, n35848);
  not g59385 (n_26565, pi0214);
  not g59386 (n_26566, n35849);
  and g59387 (n35850, n_26565, n_26566);
  and g59388 (n35851, pi0623, n_26526);
  and g59389 (n35852, n_25938, n_26525);
  not g59390 (n_26567, n35851);
  and g59391 (n35853, pi0710, n_26567);
  not g59392 (n_26568, n35852);
  and g59393 (n35854, n_26568, n35853);
  and g59394 (n35855, pi0623, n_25879);
  and g59395 (n35856, n35791, n35855);
  not g59396 (n_26569, n35854);
  not g59397 (n_26570, n35856);
  and g59398 (n35857, n_26569, n_26570);
  and g59399 (n35858, pi0214, n_4226);
  not g59400 (n_26571, n35857);
  and g59401 (n35859, n_26571, n35858);
  or g59402 (po0371, n35850, n35859);
  and g59403 (n35861, pi0215, n_14814);
  and g59404 (n35862, pi0681, pi0907);
  and g59405 (n35863, n_3149, n35862);
  and g59406 (n35864, pi0642, pi0947);
  not g59407 (n_26572, n35863);
  not g59408 (n_26573, n35864);
  and g59409 (n35865, n_26572, n_26573);
  not g59410 (n_26574, n35865);
  and g59411 (n35866, n16641, n_26574);
  and g59412 (n35867, pi0215, n_11418);
  not g59413 (n_26575, n35866);
  and g59414 (n35868, pi0038, n_26575);
  not g59415 (n_26576, n35867);
  and g59416 (n35869, n_26576, n35868);
  and g59417 (n35870, pi0215, n_11670);
  and g59418 (n35871, n16941, n_26574);
  not g59419 (n_26577, n35870);
  and g59420 (n35872, pi0299, n_26577);
  not g59421 (n_26578, n35871);
  and g59422 (n35873, n_26578, n35872);
  and g59423 (n35874, n16930, n_26574);
  and g59424 (n35875, pi0215, n_11671);
  not g59425 (n_26579, n35874);
  and g59426 (n35876, n_234, n_26579);
  not g59427 (n_26580, n35875);
  and g59428 (n35877, n_26580, n35876);
  not g59429 (n_26581, n35873);
  and g59430 (n35878, n_162, n_26581);
  not g59431 (n_26582, n35877);
  and g59432 (n35879, n_26582, n35878);
  and g59433 (n35880, n_3149, n21326);
  and g59434 (n35881, n16656, n16963);
  and g59435 (n35882, n_3139, n_11558);
  not g59436 (n_26583, n35881);
  and g59437 (n35883, n_3087, n_26583);
  not g59438 (n_26584, n35882);
  and g59439 (n35884, n_26584, n35883);
  not g59440 (n_26585, n35884);
  and g59441 (n35885, pi0947, n_26585);
  not g59442 (n_26586, n35885);
  and g59443 (n35886, n_26572, n_26586);
  not g59444 (n_26587, n35880);
  and g59445 (n35887, n_26587, n35886);
  not g59446 (n_26588, n35887);
  and g59447 (n35888, pi0299, n_26588);
  and g59448 (n35889, n2603, n_26574);
  and g59449 (n35890, n2603, n_11445);
  not g59450 (n_26589, n35862);
  and g59451 (n35891, n21431, n_26589);
  and g59452 (n35892, n_3087, n17143);
  not g59453 (n_26590, n35892);
  and g59454 (n35893, n_3119, n_26590);
  and g59455 (n35894, n_3087, n16684);
  not g59456 (n_26591, n35894);
  and g59457 (n35895, n6195, n_26591);
  and g59458 (n35896, n16769, n17167);
  and g59459 (n35897, n_24809, n16653);
  and g59460 (n35898, n_3087, n35897);
  not g59461 (n_26592, n35898);
  and g59462 (n35899, n_3139, n_26592);
  not g59463 (n_26593, n35896);
  and g59464 (n35900, n_26593, n35899);
  not g59465 (n_26594, n35895);
  not g59466 (n_26595, n35900);
  and g59467 (n35901, n_26594, n_26595);
  not g59468 (n_26596, n35901);
  and g59469 (n35902, n6205, n_26596);
  not g59470 (n_26597, n35893);
  and g59471 (n35903, pi0947, n_26597);
  not g59472 (n_26598, n35902);
  and g59473 (n35904, n_26598, n35903);
  not g59474 (n_26599, n35904);
  and g59475 (n35905, n_9349, n_26599);
  not g59476 (n_26600, n35891);
  and g59477 (n35906, n_26600, n35905);
  not g59480 (n_26602, n35890);
  and g59484 (n35910, n_3119, n_26585);
  and g59485 (n35911, n6195, n_11543);
  and g59486 (n35912, n_3139, n_11549);
  not g59487 (n_26604, n35911);
  and g59488 (n35913, n_3087, n_26604);
  not g59489 (n_26605, n35912);
  and g59490 (n35914, n_26605, n35913);
  not g59491 (n_26606, n35914);
  and g59492 (n35915, n6205, n_26606);
  not g59493 (n_26607, n35910);
  and g59494 (n35916, pi0947, n_26607);
  not g59495 (n_26608, n35915);
  and g59496 (n35917, n_26608, n35916);
  not g59497 (n_26609, n35917);
  and g59498 (n35918, n_14930, n_26609);
  and g59499 (n35919, pi0223, n_26572);
  not g59500 (n_26610, n35918);
  and g59501 (n35920, n_26610, n35919);
  not g59502 (n_26611, n35920);
  and g59503 (n35921, n_234, n_26611);
  not g59504 (n_26612, n35909);
  and g59505 (n35922, n_26612, n35921);
  not g59506 (n_26613, n35888);
  not g59507 (n_26614, n35922);
  and g59508 (n35923, n_26613, n_26614);
  not g59509 (n_26615, n35923);
  and g59510 (n35924, pi0215, n_26615);
  and g59511 (n35925, n16653, n35889);
  and g59512 (n35926, n16702, n35862);
  not g59513 (n_26616, n35926);
  and g59514 (n35927, n_3149, n_26616);
  and g59515 (n35928, pi0642, n16657);
  and g59516 (n35929, n_3139, n16699);
  not g59517 (n_26617, n35929);
  and g59518 (n35930, n_11848, n_26617);
  and g59519 (n35931, n35928, n35930);
  and g59520 (n35932, pi0642, n_11455);
  and g59521 (n35933, n_12078, n35932);
  not g59522 (n_26618, n35933);
  and g59523 (n35934, pi0947, n_26618);
  not g59524 (n_26619, n35931);
  and g59525 (n35935, n_26619, n35934);
  not g59526 (n_26620, n35927);
  not g59527 (n_26621, n35935);
  and g59528 (n35936, n_26620, n_26621);
  not g59529 (n_26622, n35936);
  and g59530 (n35937, n_3119, n_26622);
  and g59531 (n35938, n16653, n35932);
  and g59532 (n35939, n_11685, n35928);
  and g59533 (n35940, n_11698, n35939);
  not g59534 (n_26623, n35938);
  not g59535 (n_26624, n35940);
  and g59536 (n35941, n_26623, n_26624);
  not g59537 (n_26625, n35941);
  and g59538 (n35942, pi0947, n_26625);
  and g59539 (n35943, n16776, n35863);
  not g59540 (n_26626, n35942);
  and g59541 (n35944, n6205, n_26626);
  not g59542 (n_26627, n35943);
  and g59543 (n35945, n_26627, n35944);
  not g59544 (n_26628, n35937);
  and g59545 (n35946, n_9349, n_26628);
  not g59546 (n_26629, n35945);
  and g59547 (n35947, n_26629, n35946);
  not g59548 (n_26630, n35925);
  and g59549 (n35948, n_223, n_26630);
  not g59550 (n_26631, n35947);
  and g59551 (n35949, n_26631, n35948);
  and g59552 (n35950, n6205, n_11549);
  not g59553 (n_26632, n35950);
  and g59554 (n35951, n35862, n_26632);
  not g59555 (n_26633, n35951);
  and g59556 (n35952, n_3149, n_26633);
  and g59557 (n35953, pi0947, n_11556);
  not g59558 (n_26634, n35953);
  and g59559 (n35954, n_11558, n_26634);
  and g59560 (n35955, n_3119, n35954);
  and g59561 (n35956, n_11686, n35939);
  and g59562 (n35957, pi0947, n_26623);
  not g59563 (n_26635, n35956);
  and g59564 (n35958, n_26635, n35957);
  not g59565 (n_26636, n35955);
  not g59566 (n_26637, n35958);
  and g59567 (n35959, n_26636, n_26637);
  not g59568 (n_26638, n35952);
  and g59569 (n35960, n_26638, n35959);
  not g59570 (n_26639, n35960);
  and g59571 (n35961, pi0223, n_26639);
  not g59572 (n_26640, n35949);
  not g59573 (n_26641, n35961);
  and g59574 (n35962, n_26640, n_26641);
  not g59575 (n_26642, n35962);
  and g59576 (n35963, n_234, n_26642);
  and g59577 (n35964, n17026, n_26574);
  and g59578 (n35965, n_9350, n35936);
  not g59579 (n_26643, n35964);
  and g59580 (n35966, pi0299, n_26643);
  not g59581 (n_26644, n35965);
  and g59582 (n35967, n_26644, n35966);
  not g59583 (n_26645, n35967);
  and g59584 (n35968, n_36, n_26645);
  not g59585 (n_26646, n35963);
  and g59586 (n35969, n_26646, n35968);
  not g59587 (n_26647, n35924);
  not g59588 (n_26648, n35969);
  and g59589 (n35970, n_26647, n_26648);
  not g59590 (n_26649, n35970);
  and g59591 (n35971, pi0039, n_26649);
  not g59592 (n_26650, n35879);
  and g59593 (n35972, n_161, n_26650);
  not g59594 (n_26651, n35971);
  and g59595 (n35973, n_26651, n35972);
  not g59596 (n_26652, n35869);
  and g59597 (n35974, n10197, n_26652);
  not g59598 (n_26653, n35973);
  and g59599 (n35975, n_26653, n35974);
  or g59600 (po0372, n35861, n35975);
  and g59601 (n35977, pi0662, pi0907);
  and g59602 (n35978, n_3149, n35977);
  and g59603 (n35979, pi0614, pi0947);
  not g59604 (n_26654, n35978);
  not g59605 (n_26655, n35979);
  and g59606 (n35980, n_26654, n_26655);
  not g59607 (n_26656, n35980);
  and g59608 (n35981, n16641, n_26656);
  and g59609 (n35982, pi0216, n_11418);
  not g59610 (n_26657, n35981);
  and g59611 (n35983, pi0038, n_26657);
  not g59612 (n_26658, n35982);
  and g59613 (n35984, n_26658, n35983);
  and g59614 (n35985, pi0216, n_11670);
  and g59615 (n35986, n16941, n_26656);
  not g59616 (n_26659, n35985);
  and g59617 (n35987, pi0299, n_26659);
  not g59618 (n_26660, n35986);
  and g59619 (n35988, n_26660, n35987);
  and g59620 (n35989, n16930, n_26656);
  and g59621 (n35990, pi0216, n_11671);
  not g59622 (n_26661, n35989);
  and g59623 (n35991, n_234, n_26661);
  not g59624 (n_26662, n35990);
  and g59625 (n35992, n_26662, n35991);
  not g59626 (n_26663, n35988);
  and g59627 (n35993, n_162, n_26663);
  not g59628 (n_26664, n35992);
  and g59629 (n35994, n_26664, n35993);
  and g59630 (n35995, n_26632, n35977);
  not g59631 (n_26665, n35995);
  and g59632 (n35996, n_3149, n_26665);
  and g59633 (n35997, n_11686, n16997);
  and g59634 (n35998, pi0947, n_11700);
  not g59635 (n_26666, n35997);
  and g59636 (n35999, n_26666, n35998);
  not g59637 (n_26667, n35999);
  and g59638 (n36000, n_26636, n_26667);
  not g59639 (n_26668, n35996);
  and g59640 (n36001, n_26668, n36000);
  not g59641 (n_26669, n36001);
  and g59642 (n36002, pi0223, n_26669);
  and g59643 (n36003, n2603, n_26656);
  and g59644 (n36004, n16653, n36003);
  and g59645 (n36005, n35930, n35979);
  and g59646 (n36006, n16702, n35978);
  not g59647 (n_26670, n36005);
  not g59648 (n_26671, n36006);
  and g59649 (n36007, n_26670, n_26671);
  and g59650 (n36008, n_3119, n36007);
  and g59651 (n36009, n16776, n35978);
  not g59652 (n_26672, n17001);
  and g59653 (n36010, pi0947, n_26672);
  not g59654 (n_26673, n36010);
  and g59655 (n36011, n6205, n_26673);
  not g59656 (n_26674, n36009);
  and g59657 (n36012, n_26674, n36011);
  not g59658 (n_26675, n36008);
  and g59659 (n36013, n_9349, n_26675);
  not g59660 (n_26676, n36012);
  and g59661 (n36014, n_26676, n36013);
  not g59662 (n_26677, n36004);
  and g59663 (n36015, n_223, n_26677);
  not g59664 (n_26678, n36014);
  and g59665 (n36016, n_26678, n36015);
  not g59666 (n_26679, n36002);
  and g59667 (n36017, n_20, n_26679);
  not g59668 (n_26680, n36016);
  and g59669 (n36018, n_26680, n36017);
  and g59670 (n36019, n_3091, n16799);
  not g59671 (n_26681, n16978);
  and g59672 (n36020, n_3139, n_26681);
  not g59673 (n_26682, n36019);
  and g59674 (n36021, n_26682, n36020);
  and g59675 (n36022, n_3090, n_26604);
  not g59676 (n_26683, n36021);
  and g59677 (n36023, n_26683, n36022);
  not g59678 (n_26684, n36023);
  and g59679 (n36024, n6205, n_26684);
  not g59680 (n_26685, n17452);
  and g59681 (n36025, n_26685, n_24625);
  and g59682 (n36026, n_24626, n36025);
  not g59683 (n_26686, n36026);
  and g59684 (n36027, n17002, n_26686);
  and g59685 (n36028, n_3090, n_11479);
  and g59686 (n36029, n6195, n36028);
  not g59687 (n_26687, n36027);
  not g59688 (n_26688, n36029);
  and g59689 (n36030, n_26687, n_26688);
  and g59690 (n36031, n_3119, n36030);
  not g59691 (n_26689, n36031);
  and g59692 (n36032, pi0947, n_26689);
  not g59693 (n_26690, n36024);
  and g59694 (n36033, n_26690, n36032);
  not g59695 (n_26691, n36033);
  and g59696 (n36034, n_14930, n_26691);
  and g59697 (n36035, pi0223, n_26654);
  not g59698 (n_26692, n36034);
  and g59699 (n36036, n_26692, n36035);
  and g59700 (n36037, n_3090, n17143);
  not g59701 (n_26693, n36037);
  and g59702 (n36038, pi0947, n_26693);
  and g59703 (n36039, n_3149, n_11712);
  not g59705 (n_26694, n36038);
  not g59707 (n_26695, n36039);
  not g59709 (n_26696, n17008);
  and g59710 (n36043, pi0947, n_26696);
  and g59711 (n36044, n_3149, n17011);
  not g59712 (n_26697, n35977);
  and g59713 (n36045, n_26697, n36044);
  not g59714 (n_26698, n36043);
  not g59715 (n_26699, n36045);
  and g59716 (n36046, n_26698, n_26699);
  not g59717 (n_26700, n36046);
  and g59718 (n36047, n6205, n_26700);
  not g59719 (n_26701, n36042);
  and g59720 (n36048, n_9349, n_26701);
  not g59721 (n_26702, n36047);
  and g59722 (n36049, n_26702, n36048);
  not g59728 (n_26705, n36036);
  and g59729 (n36053, pi0216, n_26705);
  not g59730 (n_26706, n36052);
  and g59731 (n36054, n_26706, n36053);
  not g59732 (n_26707, n36018);
  and g59733 (n36055, n_234, n_26707);
  not g59734 (n_26708, n36054);
  and g59735 (n36056, n_26708, n36055);
  not g59736 (n_26709, n36007);
  and g59737 (n36057, n5777, n_26709);
  and g59738 (n36058, n17026, n_26656);
  and g59739 (n36059, n_3149, n20994);
  and g59740 (n36060, n_26654, n_26694);
  not g59741 (n_26710, n36059);
  and g59742 (n36061, n_26710, n36060);
  not g59743 (n_26711, n36061);
  and g59744 (n36062, pi0216, n_26711);
  not g59745 (n_26712, n36057);
  not g59746 (n_26713, n36058);
  and g59747 (n36063, n_26712, n_26713);
  not g59748 (n_26714, n36062);
  and g59749 (n36064, n_26714, n36063);
  not g59750 (n_26715, n36064);
  and g59751 (n36065, n_36, n_26715);
  and g59752 (n36066, n16814, n35977);
  not g59753 (n_26716, n36066);
  and g59754 (n36067, n_3149, n_26716);
  and g59755 (n36068, pi0947, n16723);
  not g59756 (n_26717, n36068);
  and g59757 (n36069, n_26667, n_26717);
  not g59758 (n_26718, n36067);
  and g59759 (n36070, n_26718, n36069);
  not g59760 (n_26719, n36070);
  and g59761 (n36071, n_20, n_26719);
  and g59762 (n36072, pi0947, n36030);
  not g59767 (n_26721, n36071);
  and g59768 (n36076, pi0215, n_26721);
  not g59769 (n_26722, n36075);
  and g59770 (n36077, n_26722, n36076);
  not g59771 (n_26723, n36077);
  and g59772 (n36078, pi0299, n_26723);
  not g59773 (n_26724, n36065);
  and g59774 (n36079, n_26724, n36078);
  not g59775 (n_26725, n36056);
  and g59776 (n36080, pi0039, n_26725);
  not g59777 (n_26726, n36079);
  and g59778 (n36081, n_26726, n36080);
  not g59779 (n_26727, n35994);
  and g59780 (n36082, n_161, n_26727);
  not g59781 (n_26728, n36081);
  and g59782 (n36083, n_26728, n36082);
  not g59783 (n_26729, n35984);
  not g59784 (n_26730, n36083);
  and g59785 (n36084, n_26729, n_26730);
  not g59786 (n_26731, n36084);
  and g59787 (n36085, n10197, n_26731);
  and g59788 (n36086, n_20, n_14814);
  not g59789 (n_26732, n36085);
  not g59790 (n_26733, n36086);
  and g59791 (po0373, n_26732, n_26733);
  not g59792 (n_26735, pi0695);
  and g59793 (n36088, n_26735, n35600);
  not g59794 (n_26736, n36088);
  and g59795 (n36089, pi0217, n_26736);
  not g59796 (n_26737, n35485);
  and g59797 (n36090, pi0695, n_26737);
  not g59798 (n_26738, n35524);
  and g59799 (n36091, n_26735, n_26738);
  not g59800 (n_26739, n36090);
  and g59801 (n36092, n_5623, n_26739);
  not g59802 (n_26740, n36091);
  and g59803 (n36093, n_26740, n36092);
  not g59804 (n_26742, pi0612);
  not g59805 (n_26743, n36089);
  and g59806 (n36094, n_26742, n_26743);
  not g59807 (n_26744, n36093);
  and g59808 (n36095, n_26744, n36094);
  and g59809 (n36096, n_26735, n35638);
  and g59810 (n36097, pi0695, n35578);
  not g59811 (n_26745, n36097);
  and g59812 (n36098, pi0217, n_26745);
  not g59813 (n_26746, n36096);
  and g59814 (n36099, n_26746, n36098);
  not g59815 (n_26747, n35543);
  and g59816 (n36100, pi0695, n_26747);
  not g59817 (n_26748, n35566);
  and g59818 (n36101, n_26735, n_26748);
  not g59819 (n_26749, n36100);
  and g59820 (n36102, n_5623, n_26749);
  not g59821 (n_26750, n36101);
  and g59822 (n36103, n_26750, n36102);
  not g59823 (n_26751, n36099);
  and g59824 (n36104, pi0612, n_26751);
  not g59825 (n_26752, n36103);
  and g59826 (n36105, n_26752, n36104);
  or g59827 (po0374, n36095, n36105);
  and g59828 (n36107, n_25731, n_25766);
  and g59829 (n36108, n34786, n_25818);
  not g59830 (n_26753, n36107);
  not g59831 (n_26754, n36108);
  and g59832 (n36109, n_26753, n_26754);
  not g59833 (n_26756, pi0218);
  not g59834 (n_26757, n36109);
  and g59835 (n36110, n_26756, n_26757);
  and g59836 (n36111, n34786, n34899);
  not g59837 (n_26758, n36111);
  and g59838 (n36112, pi0218, n_26758);
  not g59839 (n_26759, n36110);
  not g59840 (n_26760, n36112);
  and g59841 (po0375, n_26759, n_26760);
  and g59842 (n36114, n_6791, n_4226);
  and g59843 (n36115, pi0617, n_26526);
  and g59844 (n36116, n_25117, n_26525);
  not g59845 (n_26761, n36115);
  and g59846 (n36117, pi0637, n_26761);
  not g59847 (n_26762, n36116);
  and g59848 (n36118, n_26762, n36117);
  and g59849 (n36119, pi0617, n_25155);
  and g59850 (n36120, n35791, n36119);
  not g59851 (n_26763, n36118);
  not g59852 (n_26764, n36120);
  and g59853 (n36121, n_26763, n_26764);
  not g59854 (n_26765, n36121);
  and g59855 (n36122, n36114, n_26765);
  and g59856 (n36123, n_25117, n35771);
  and g59857 (n36124, pi0617, n35773);
  not g59858 (n_26766, n36123);
  and g59859 (n36125, pi0637, n_26766);
  not g59860 (n_26767, n36124);
  and g59861 (n36126, n_26767, n36125);
  and g59862 (n36127, n_25117, n17059);
  and g59863 (n36128, pi0617, n35778);
  not g59864 (n_26768, n36127);
  and g59865 (n36129, n_25155, n_26768);
  not g59866 (n_26769, n36128);
  and g59867 (n36130, n_26769, n36129);
  not g59868 (n_26770, n36130);
  and g59869 (n36131, n_4226, n_26770);
  not g59870 (n_26771, n36126);
  and g59871 (n36132, n_26771, n36131);
  not g59872 (n_26772, n36132);
  and g59873 (n36133, pi0219, n_26772);
  or g59874 (po0376, n36122, n36133);
  and g59875 (n36135, n_25596, n_25839);
  and g59876 (n36136, n_25705, n34910);
  not g59877 (n_26773, n36135);
  not g59878 (n_26774, n36136);
  and g59879 (n36137, n_26773, n_26774);
  not g59880 (n_26776, pi0220);
  not g59881 (n_26777, n36137);
  and g59882 (n36138, n_26776, n_26777);
  and g59883 (n36139, n34774, n34910);
  not g59884 (n_26778, n36139);
  and g59885 (n36140, pi0220, n_26778);
  not g59886 (n_26779, n36138);
  not g59887 (n_26780, n36140);
  and g59888 (po0377, n_26779, n_26780);
  and g59889 (n36142, pi0661, pi0907);
  and g59890 (n36143, n_3149, n36142);
  and g59891 (n36144, pi0616, pi0947);
  not g59892 (n_26781, n36143);
  not g59893 (n_26782, n36144);
  and g59894 (n36145, n_26781, n_26782);
  not g59895 (n_26783, n36145);
  and g59896 (n36146, n16641, n_26783);
  and g59897 (n36147, pi0221, n_11418);
  not g59898 (n_26784, n36146);
  and g59899 (n36148, pi0038, n_26784);
  not g59900 (n_26785, n36147);
  and g59901 (n36149, n_26785, n36148);
  and g59902 (n36150, pi0221, n_11670);
  and g59903 (n36151, n16941, n_26783);
  not g59904 (n_26786, n36150);
  and g59905 (n36152, pi0299, n_26786);
  not g59906 (n_26787, n36151);
  and g59907 (n36153, n_26787, n36152);
  and g59908 (n36154, n16930, n_26783);
  and g59909 (n36155, pi0221, n_11671);
  not g59910 (n_26788, n36154);
  and g59911 (n36156, n_234, n_26788);
  not g59912 (n_26789, n36155);
  and g59913 (n36157, n_26789, n36156);
  not g59914 (n_26790, n36153);
  and g59915 (n36158, n_162, n_26790);
  not g59916 (n_26791, n36157);
  and g59917 (n36159, n_26791, n36158);
  not g59918 (n_26792, n16980);
  and g59919 (n36160, pi0947, n_26792);
  not g59920 (n_26793, n36160);
  and g59921 (n36161, n_26781, n_26793);
  and g59922 (n36162, n35950, n_26793);
  not g59923 (n_26794, n36161);
  and g59924 (n36163, n_26636, n_26794);
  not g59925 (n_26795, n36162);
  and g59926 (n36164, n_26795, n36163);
  not g59927 (n_26796, n36164);
  and g59928 (n36165, pi0223, n_26796);
  and g59929 (n36166, n16653, n_26783);
  and g59930 (n36167, n2603, n36166);
  not g59931 (n_26797, n36167);
  and g59932 (n36168, n_223, n_26797);
  and g59933 (n36169, n16976, n_11698);
  not g59934 (n_26798, n36169);
  and g59935 (n36170, n_11688, n_26798);
  not g59936 (n_26799, n36170);
  and g59937 (n36171, pi0947, n_26799);
  and g59938 (n36172, n16776, n36143);
  not g59939 (n_26800, n36171);
  and g59940 (n36173, n6205, n_26800);
  not g59941 (n_26801, n36172);
  and g59942 (n36174, n_26801, n36173);
  and g59943 (n36175, n35930, n36144);
  and g59944 (n36176, n16702, n36143);
  not g59945 (n_26802, n36175);
  not g59946 (n_26803, n36176);
  and g59947 (n36177, n_26802, n_26803);
  and g59948 (n36178, n_3119, n36177);
  not g59949 (n_26804, n36178);
  and g59950 (n36179, n_9349, n_26804);
  not g59951 (n_26805, n36174);
  and g59952 (n36180, n_26805, n36179);
  not g59953 (n_26806, n36180);
  and g59954 (n36181, n36168, n_26806);
  not g59955 (n_26807, n36165);
  and g59956 (n36182, n_26, n_26807);
  not g59957 (n_26808, n36181);
  and g59958 (n36183, n_26808, n36182);
  and g59959 (n36184, n_26590, n_26619);
  not g59960 (n_26809, n36184);
  and g59961 (n36185, n16984, n_26809);
  and g59962 (n36186, n_3102, n16774);
  not g59963 (n_26810, n36186);
  and g59964 (n36187, n_11460, n_26810);
  not g59965 (n_26811, n36187);
  and g59966 (n36188, n16981, n_26811);
  not g59967 (n_26812, n36185);
  and g59968 (n36189, pi0947, n_26812);
  not g59969 (n_26813, n36188);
  and g59970 (n36190, n_26813, n36189);
  not g59971 (n_26814, n36190);
  and g59972 (n36191, n_26695, n_26814);
  not g59973 (n_26815, n36191);
  and g59974 (n36192, n_3119, n_26815);
  and g59975 (n36193, n16774, n16981);
  and g59976 (n36194, n_11699, n17008);
  not g59977 (n_26816, n36194);
  and g59978 (n36195, n16984, n_26816);
  not g59979 (n_26817, n36193);
  not g59980 (n_26818, n36195);
  and g59981 (n36196, n_26817, n_26818);
  not g59982 (n_26819, n36196);
  and g59983 (n36197, pi0947, n_26819);
  not g59984 (n_26820, n36044);
  and g59985 (n36198, n6205, n_26820);
  not g59986 (n_26821, n36197);
  and g59987 (n36199, n_26821, n36198);
  not g59988 (n_26822, n36192);
  and g59989 (n36200, n_26781, n_26822);
  not g59990 (n_26823, n36199);
  and g59991 (n36201, n_26823, n36200);
  not g59992 (n_26824, n36201);
  and g59993 (n36202, n_9349, n_26824);
  and g59994 (n36203, n_26602, n36168);
  not g59995 (n_26825, n36202);
  and g59996 (n36204, n_26825, n36203);
  and g59997 (n36205, n_3149, n16990);
  not g59998 (n_26826, n16987);
  and g59999 (n36206, pi0947, n_26826);
  not g60000 (n_26827, n36206);
  and g60001 (n36207, n6205, n_26827);
  not g60002 (n_26828, n36205);
  and g60003 (n36208, n_26828, n36207);
  and g60004 (n36209, n_3149, n_11684);
  and g60005 (n36210, n_11556, n_11546);
  not g60006 (n_26829, n36210);
  and g60007 (n36211, n_3139, n_26829);
  and g60008 (n36212, n_3091, n_26583);
  not g60009 (n_26830, n36211);
  and g60010 (n36213, n_26830, n36212);
  not g60011 (n_26831, n36213);
  and g60012 (n36214, pi0947, n_26831);
  not g60013 (n_26832, n36209);
  not g60014 (n_26833, n36214);
  and g60015 (n36215, n_26832, n_26833);
  not g60016 (n_26834, n36215);
  and g60017 (n36216, n_3119, n_26834);
  not g60023 (n_26837, n36219);
  and g60024 (n36220, pi0221, n_26837);
  not g60025 (n_26838, n36204);
  and g60026 (n36221, n_26838, n36220);
  not g60027 (n_26839, n36183);
  and g60028 (n36222, n_234, n_26839);
  not g60029 (n_26840, n36221);
  and g60030 (n36223, n_26840, n36222);
  not g60031 (n_26841, n36142);
  and g60032 (n36224, n_14885, n_26841);
  not g60033 (n_26842, n36224);
  and g60034 (n36225, n_3149, n_26842);
  and g60035 (n36226, pi0221, n_26814);
  not g60036 (n_26843, n36225);
  and g60037 (n36227, n_26843, n36226);
  not g60038 (n_26844, n36177);
  and g60039 (n36228, pi0216, n_26844);
  and g60040 (n36229, n_20, n36166);
  not g60041 (n_26845, n36229);
  and g60042 (n36230, n_26, n_26845);
  not g60043 (n_26846, n36228);
  and g60044 (n36231, n_26846, n36230);
  not g60045 (n_26847, n36231);
  and g60046 (n36232, n_36, n_26847);
  not g60047 (n_26848, n36227);
  and g60048 (n36233, n_26848, n36232);
  not g60052 (n_26849, n35954);
  and g60053 (n36237, n_26849, n_26794);
  not g60054 (n_26850, n36237);
  and g60055 (n36238, n_26, n_26850);
  not g60056 (n_26851, n36238);
  and g60057 (n36239, pi0215, n_26851);
  not g60058 (n_26852, n36236);
  and g60059 (n36240, n_26852, n36239);
  not g60060 (n_26853, n36240);
  and g60061 (n36241, pi0299, n_26853);
  not g60062 (n_26854, n36233);
  and g60063 (n36242, n_26854, n36241);
  not g60064 (n_26855, n36223);
  and g60065 (n36243, pi0039, n_26855);
  not g60066 (n_26856, n36242);
  and g60067 (n36244, n_26856, n36243);
  not g60068 (n_26857, n36159);
  and g60069 (n36245, n_161, n_26857);
  not g60070 (n_26858, n36244);
  and g60071 (n36246, n_26858, n36245);
  not g60072 (n_26859, n36149);
  not g60073 (n_26860, n36246);
  and g60074 (n36247, n_26859, n_26860);
  not g60075 (n_26861, n36247);
  and g60076 (n36248, n10197, n_26861);
  and g60077 (n36249, n_26, n_14814);
  not g60078 (n_26862, n36248);
  not g60079 (n_26863, n36249);
  and g60080 (po0378, n_26862, n_26863);
  and g60081 (n36251, n_223, n_15206);
  not g60082 (n_26864, n36251);
  and g60083 (n36252, n_11717, n_26864);
  not g60084 (n_26865, n36252);
  and g60085 (n36253, n_234, n_26865);
  not g60086 (n_26866, n36253);
  and g60087 (n36254, pi0039, n_26866);
  and g60088 (n36255, n_11735, n36254);
  and g60089 (n36256, n_161, n_12667);
  not g60090 (n_26867, n36255);
  and g60091 (n36257, n_26867, n36256);
  not g60092 (n_26868, n36257);
  and g60093 (n36258, n18591, n_26868);
  not g60094 (n_26869, n36258);
  and g60095 (n36259, pi0222, n_26869);
  not g60096 (n_26870, n36259);
  and g60097 (n36260, n_24651, n_26870);
  and g60098 (n36261, pi0222, n_11417);
  and g60099 (n36262, pi0222, n_11418);
  not g60100 (n_26871, n36262);
  and g60101 (n36263, pi0038, n_26871);
  and g60102 (n36264, pi0661, n16646);
  not g60103 (n_26872, n36264);
  and g60104 (n36265, n36263, n_26872);
  and g60105 (n36266, pi0661, pi0680);
  not g60106 (n_26873, n36266);
  and g60107 (n36267, n16918, n_26873);
  and g60108 (n36268, n_226, n_12231);
  and g60109 (n36269, pi0222, n16935);
  and g60116 (n36273, pi0222, n16944);
  and g60117 (n36274, n16923, n_26873);
  and g60118 (n36275, n_226, n_12235);
  not g60125 (n_26880, n36272);
  and g60126 (n36279, n_162, n_26880);
  not g60127 (n_26881, n36278);
  and g60128 (n36280, n_26881, n36279);
  and g60129 (n36281, n_3096, n_11712);
  and g60130 (n36282, pi0680, n16758);
  not g60131 (n_26882, n36282);
  and g60132 (n36283, n_11509, n_26882);
  not g60133 (n_26883, n36283);
  and g60134 (n36284, pi0661, n_26883);
  not g60135 (n_26884, n36281);
  not g60136 (n_26885, n36284);
  and g60137 (n36285, n_26884, n_26885);
  and g60138 (n36286, n_3119, n36285);
  and g60139 (n36287, n_3096, n16994);
  and g60140 (n36288, n_11675, n_11526);
  and g60141 (n36289, n_3093, n16995);
  not g60142 (n_26886, n36288);
  not g60143 (n_26887, n36289);
  and g60144 (n36290, n_26886, n_26887);
  not g60145 (n_26888, n36290);
  and g60146 (n36291, n16656, n_26888);
  not g60147 (n_26889, n16786);
  and g60148 (n36292, pi0661, n_26889);
  not g60149 (n_26890, n36287);
  not g60150 (n_26891, n36291);
  and g60151 (n36293, n_26890, n_26891);
  not g60152 (n_26892, n36292);
  and g60153 (n36294, n_26892, n36293);
  and g60154 (n36295, n6205, n36294);
  not g60155 (n_26893, n36286);
  and g60156 (n36296, pi0222, n_26893);
  not g60157 (n_26894, n36295);
  and g60158 (n36297, n_26894, n36296);
  not g60159 (n_26895, n16690);
  and g60160 (n36298, n_26895, n36266);
  and g60161 (n36299, n6205, n36298);
  and g60162 (n36300, pi0661, n16703);
  and g60163 (n36301, n_3119, n36300);
  not g60164 (n_26896, n36299);
  and g60165 (n36302, pi0224, n_26896);
  not g60166 (n_26897, n36301);
  and g60167 (n36303, n_26897, n36302);
  and g60168 (n36304, pi0661, n16739);
  not g60169 (n_26898, n36304);
  and g60170 (n36305, n_219, n_26898);
  not g60171 (n_26899, n36305);
  and g60172 (n36306, n_226, n_26899);
  not g60173 (n_26900, n36303);
  and g60174 (n36307, n_26900, n36306);
  not g60175 (n_26901, n36307);
  and g60176 (n36308, n_223, n_26901);
  not g60177 (n_26902, n36297);
  and g60178 (n36309, n_26902, n36308);
  and g60179 (n36310, n_226, pi0661);
  and g60180 (n36311, n16729, n36310);
  and g60181 (n36312, n_3096, n16960);
  and g60182 (n36313, n16656, n16966);
  not g60183 (n_26903, n16818);
  and g60184 (n36314, pi0661, n_26903);
  not g60185 (n_26904, n36312);
  not g60186 (n_26905, n36314);
  and g60187 (n36315, n_26904, n_26905);
  not g60188 (n_26906, n36313);
  and g60189 (n36316, n_26906, n36315);
  and g60190 (n36317, n_3119, n36316);
  and g60191 (n36318, n_3096, n_11694);
  and g60192 (n36319, n_11555, n_11554);
  not g60193 (n_26907, n36319);
  and g60194 (n36320, pi0661, n_26907);
  not g60195 (n_26908, n36318);
  not g60196 (n_26909, n36320);
  and g60197 (n36321, n_26908, n_26909);
  and g60198 (n36322, n6205, n36321);
  not g60199 (n_26910, n36317);
  and g60200 (n36323, pi0222, n_26910);
  not g60201 (n_26911, n36322);
  and g60202 (n36324, n_26911, n36323);
  not g60203 (n_26912, n36311);
  and g60204 (n36325, pi0223, n_26912);
  not g60205 (n_26913, n36324);
  and g60206 (n36326, n_26913, n36325);
  not g60207 (n_26914, n36309);
  not g60208 (n_26915, n36326);
  and g60209 (n36327, n_26914, n_26915);
  not g60210 (n_26916, n36327);
  and g60211 (n36328, n_234, n_26916);
  and g60212 (n36329, n16744, n36310);
  and g60213 (n36330, n_3162, n36316);
  and g60214 (n36331, n6242, n36321);
  not g60215 (n_26917, n36330);
  and g60216 (n36332, pi0222, n_26917);
  not g60217 (n_26918, n36331);
  and g60218 (n36333, n_26918, n36332);
  not g60219 (n_26919, n36329);
  not g60220 (n_26920, n36333);
  and g60221 (n36334, n_26919, n_26920);
  not g60222 (n_26921, n36334);
  and g60223 (n36335, pi0215, n_26921);
  and g60224 (n36336, pi0222, n_11445);
  not g60225 (n_26922, n36336);
  and g60226 (n36337, n3448, n_26922);
  and g60227 (n36338, n_26898, n36337);
  and g60228 (n36339, n_3162, n36285);
  and g60229 (n36340, n6242, n36294);
  not g60230 (n_26923, n36339);
  and g60231 (n36341, pi0222, n_26923);
  not g60232 (n_26924, n36340);
  and g60233 (n36342, n_26924, n36341);
  not g60234 (n_26925, n36300);
  and g60235 (n36343, n_3162, n_26925);
  not g60236 (n_26926, n36298);
  and g60237 (n36344, n6242, n_26926);
  not g60238 (n_26927, n36343);
  and g60239 (n36345, n_226, n_26927);
  not g60240 (n_26928, n36344);
  and g60241 (n36346, n_26928, n36345);
  not g60242 (n_26929, n36346);
  and g60243 (n36347, n_9350, n_26929);
  not g60244 (n_26930, n36342);
  and g60245 (n36348, n_26930, n36347);
  not g60246 (n_26931, n36338);
  and g60247 (n36349, n_36, n_26931);
  not g60248 (n_26932, n36348);
  and g60249 (n36350, n_26932, n36349);
  not g60250 (n_26933, n36335);
  and g60251 (n36351, pi0299, n_26933);
  not g60252 (n_26934, n36350);
  and g60253 (n36352, n_26934, n36351);
  not g60254 (n_26935, n36328);
  not g60255 (n_26936, n36352);
  and g60256 (n36353, n_26935, n_26936);
  not g60257 (n_26937, n36353);
  and g60258 (n36354, pi0039, n_26937);
  not g60259 (n_26938, n36280);
  not g60260 (n_26939, n36354);
  and g60261 (n36355, n_26938, n_26939);
  not g60262 (n_26940, n36355);
  and g60263 (n36356, n_161, n_26940);
  not g60264 (n_26941, n36265);
  and g60265 (n36357, n2571, n_26941);
  not g60266 (n_26942, n36356);
  and g60267 (n36358, n_26942, n36357);
  not g60268 (n_26943, n36261);
  not g60269 (n_26944, n36358);
  and g60270 (n36359, n_26943, n_26944);
  not g60271 (n_26945, n36359);
  and g60272 (n36360, n_11749, n_26945);
  and g60273 (n36361, pi0625, n36359);
  and g60274 (n36362, n_11753, n_26870);
  not g60275 (n_26946, n36362);
  and g60276 (n36363, pi1153, n_26946);
  not g60277 (n_26947, n36361);
  and g60278 (n36364, n_26947, n36363);
  and g60279 (n36365, n_11753, n36359);
  and g60280 (n36366, pi0625, n_26870);
  not g60281 (n_26948, n36366);
  and g60282 (n36367, n_11757, n_26948);
  not g60283 (n_26949, n36365);
  and g60284 (n36368, n_26949, n36367);
  not g60285 (n_26950, n36364);
  not g60286 (n_26951, n36368);
  and g60287 (n36369, n_26950, n_26951);
  not g60288 (n_26952, n36369);
  and g60289 (n36370, pi0778, n_26952);
  not g60290 (n_26953, n36360);
  not g60291 (n_26954, n36370);
  and g60292 (n36371, n_26953, n_26954);
  not g60293 (n_26955, n36371);
  and g60294 (n36372, n_11773, n_26955);
  and g60295 (n36373, n17075, n36259);
  not g60296 (n_26956, n36372);
  not g60297 (n_26957, n36373);
  and g60298 (n36374, n_26956, n_26957);
  not g60299 (n_26958, n36374);
  and g60300 (n36375, n_11777, n_26958);
  and g60301 (n36376, n16639, n36259);
  not g60302 (n_26959, n36375);
  not g60303 (n_26960, n36376);
  and g60304 (n36377, n_26959, n_26960);
  and g60305 (n36378, n_11780, n36377);
  and g60306 (n36379, n_11783, n36378);
  not g60307 (n_26961, n36260);
  not g60308 (n_26962, n36379);
  and g60309 (n36380, n_26961, n_26962);
  not g60310 (n_26963, n36380);
  and g60311 (n36381, n_13453, n_26963);
  and g60312 (n36382, n17856, n_26870);
  not g60313 (n_26964, n36381);
  not g60314 (n_26965, n36382);
  and g60315 (n36383, n_26964, n_26965);
  and g60316 (n36384, n_11803, n36383);
  not g60317 (n_26966, n36383);
  and g60318 (n36385, n_11806, n_26966);
  and g60319 (n36386, pi0647, n_26870);
  not g60320 (n_26967, n36386);
  and g60321 (n36387, n_11810, n_26967);
  not g60322 (n_26968, n36385);
  and g60323 (n36388, n_26968, n36387);
  and g60324 (n36389, pi0647, n_26966);
  and g60325 (n36390, n_11806, n_26870);
  not g60326 (n_26969, n36390);
  and g60327 (n36391, pi1157, n_26969);
  not g60328 (n_26970, n36389);
  and g60329 (n36392, n_26970, n36391);
  not g60330 (n_26971, n36388);
  not g60331 (n_26972, n36392);
  and g60332 (n36393, n_26971, n_26972);
  not g60333 (n_26973, n36393);
  and g60334 (n36394, pi0787, n_26973);
  not g60335 (n_26974, n36384);
  not g60336 (n_26975, n36394);
  and g60337 (n36395, n_26974, n_26975);
  and g60338 (n36396, n_11819, n36395);
  and g60339 (n36397, pi0628, n_26870);
  and g60340 (n36398, n_11789, n_26963);
  not g60341 (n_26976, n36397);
  and g60342 (n36399, n17777, n_26976);
  not g60343 (n_26977, n36398);
  and g60344 (n36400, n_26977, n36399);
  and g60345 (n36401, n17969, n_26870);
  and g60346 (n36402, pi0616, n17280);
  not g60347 (n_26978, n36402);
  and g60348 (n36403, n36263, n_26978);
  and g60349 (n36404, n_3091, n17233);
  and g60350 (n36405, n_226, n_11923);
  and g60351 (n36406, pi0222, n17139);
  and g60358 (n36410, n_3139, n17235);
  not g60359 (n_26982, n36410);
  and g60360 (n36411, n_11925, n_26982);
  not g60361 (n_26983, n36411);
  and g60362 (n36412, pi0616, n_26983);
  and g60363 (n36413, n_226, n36412);
  and g60364 (n36414, n_11494, n36413);
  not g60365 (n_26984, n17182);
  and g60366 (n36415, pi0616, n_26984);
  not g60367 (n_26985, n36415);
  and g60368 (n36416, n16814, n_26985);
  not g60369 (n_26986, n16656);
  not g60370 (n_26987, n36416);
  and g60371 (n36417, n_26986, n_26987);
  and g60372 (n36418, n_11675, n_11558);
  and g60373 (n36419, n_11676, n_26985);
  not g60374 (n_26988, n36418);
  and g60375 (n36420, n_26988, n36419);
  not g60376 (n_26989, n36420);
  and g60377 (n36421, n16656, n_26989);
  not g60378 (n_26990, n36417);
  not g60379 (n_26991, n36421);
  and g60380 (n36422, n_26990, n_26991);
  and g60381 (n36423, n_3162, n36422);
  not g60382 (n_26992, n17169);
  and g60383 (n36424, pi0616, n_26992);
  not g60384 (n_26993, n36424);
  and g60385 (n36425, n_11548, n_26993);
  not g60386 (n_26994, n36425);
  and g60387 (n36426, n_26986, n_26994);
  and g60388 (n36427, pi0616, n17168);
  not g60389 (n_26995, n36427);
  and g60390 (n36428, n6193, n_26995);
  and g60391 (n36429, n16797, n36428);
  and g60392 (n36430, n_11675, n36425);
  not g60393 (n_26996, n36429);
  and g60394 (n36431, n16656, n_26996);
  not g60395 (n_26997, n36430);
  and g60396 (n36432, n_26997, n36431);
  not g60397 (n_26998, n36426);
  not g60398 (n_26999, n36432);
  and g60399 (n36433, n_26998, n_26999);
  and g60400 (n36434, n6242, n36433);
  not g60401 (n_27000, n36423);
  and g60402 (n36435, pi0222, n_27000);
  not g60403 (n_27001, n36434);
  and g60404 (n36436, n_27001, n36435);
  not g60405 (n_27002, n36414);
  not g60406 (n_27003, n36436);
  and g60407 (n36437, n_27002, n_27003);
  not g60408 (n_27004, n36437);
  and g60409 (n36438, pi0215, n_27004);
  and g60410 (n36439, n16978, n17168);
  not g60411 (n_27005, n36439);
  and g60412 (n36440, n36337, n_27005);
  and g60413 (n36441, n_11525, n_26993);
  not g60414 (n_27006, n36441);
  and g60415 (n36442, n_26986, n_27006);
  and g60416 (n36443, n16684, n36428);
  and g60417 (n36444, n_11675, n36441);
  not g60418 (n_27007, n36443);
  and g60419 (n36445, n16656, n_27007);
  not g60420 (n_27008, n36444);
  and g60421 (n36446, n_27008, n36445);
  not g60422 (n_27009, n36442);
  not g60423 (n_27010, n36446);
  and g60424 (n36447, n_27009, n_27010);
  and g60425 (n36448, n6242, n36447);
  and g60426 (n36449, pi0616, n_11856);
  and g60427 (n36450, n_3091, n36187);
  not g60428 (n_27011, n36449);
  not g60429 (n_27012, n36450);
  and g60430 (n36451, n_27011, n_27012);
  not g60431 (n_27013, n36451);
  and g60432 (n36452, n_26986, n_27013);
  and g60433 (n36453, n17147, n_26995);
  not g60434 (n_27014, n36453);
  and g60435 (n36454, n_11854, n_27014);
  not g60436 (n_27015, n36454);
  and g60437 (n36455, n6193, n_27015);
  and g60438 (n36456, n_11675, n36451);
  not g60439 (n_27016, n36455);
  and g60440 (n36457, n16656, n_27016);
  not g60441 (n_27017, n36456);
  and g60442 (n36458, n_27017, n36457);
  not g60443 (n_27018, n36452);
  not g60444 (n_27019, n36458);
  and g60445 (n36459, n_27018, n_27019);
  and g60446 (n36460, n_3162, n36459);
  not g60447 (n_27020, n36448);
  and g60448 (n36461, pi0222, n_27020);
  not g60449 (n_27021, n36460);
  and g60450 (n36462, n_27021, n36461);
  and g60451 (n36463, n_11932, n_26982);
  not g60452 (n_27022, n36463);
  and g60453 (n36464, pi0616, n_27022);
  not g60454 (n_27023, n36464);
  and g60455 (n36465, n6242, n_27023);
  and g60456 (n36466, n_12078, n36427);
  not g60457 (n_27024, n36466);
  and g60458 (n36467, n_26986, n_27024);
  and g60459 (n36468, pi0616, n6193);
  and g60460 (n36469, n17375, n36468);
  and g60461 (n36470, n_11675, n36466);
  not g60462 (n_27025, n36469);
  and g60463 (n36471, n16656, n_27025);
  not g60464 (n_27026, n36470);
  and g60465 (n36472, n_27026, n36471);
  not g60466 (n_27027, n36467);
  not g60467 (n_27028, n36472);
  and g60468 (n36473, n_27027, n_27028);
  not g60469 (n_27029, n36473);
  and g60470 (n36474, n_3162, n_27029);
  not g60471 (n_27030, n36465);
  and g60472 (n36475, n_226, n_27030);
  not g60473 (n_27031, n36474);
  and g60474 (n36476, n_27031, n36475);
  not g60475 (n_27032, n36476);
  and g60476 (n36477, n_9350, n_27032);
  not g60477 (n_27033, n36462);
  and g60478 (n36478, n_27033, n36477);
  not g60479 (n_27034, n36440);
  and g60480 (n36479, n_36, n_27034);
  not g60481 (n_27035, n36478);
  and g60482 (n36480, n_27035, n36479);
  not g60483 (n_27036, n36438);
  and g60484 (n36481, pi0299, n_27036);
  not g60485 (n_27037, n36480);
  and g60486 (n36482, n_27037, n36481);
  and g60487 (n36483, n6205, n36464);
  and g60488 (n36484, n_3119, n36473);
  not g60489 (n_27038, n36483);
  and g60490 (n36485, pi0224, n_27038);
  not g60491 (n_27039, n36484);
  and g60492 (n36486, n_27039, n36485);
  and g60493 (n36487, n_219, n_27005);
  not g60494 (n_27040, n36487);
  and g60495 (n36488, n_226, n_27040);
  not g60496 (n_27041, n36486);
  and g60497 (n36489, n_27041, n36488);
  and g60498 (n36490, n6205, n36447);
  and g60499 (n36491, n_3119, n36459);
  not g60500 (n_27042, n36490);
  and g60501 (n36492, pi0222, n_27042);
  not g60502 (n_27043, n36491);
  and g60503 (n36493, n_27043, n36492);
  not g60504 (n_27044, n36489);
  and g60505 (n36494, n_223, n_27044);
  not g60506 (n_27045, n36493);
  and g60507 (n36495, n_27045, n36494);
  and g60508 (n36496, n_11484, n36413);
  and g60509 (n36497, n_3119, n36422);
  and g60510 (n36498, n6205, n36433);
  not g60511 (n_27046, n36497);
  and g60512 (n36499, pi0222, n_27046);
  not g60513 (n_27047, n36498);
  and g60514 (n36500, n_27047, n36499);
  not g60515 (n_27048, n36496);
  and g60516 (n36501, pi0223, n_27048);
  not g60517 (n_27049, n36500);
  and g60518 (n36502, n_27049, n36501);
  not g60519 (n_27050, n36495);
  not g60520 (n_27051, n36502);
  and g60521 (n36503, n_27050, n_27051);
  not g60522 (n_27052, n36503);
  and g60523 (n36504, n_234, n_27052);
  not g60524 (n_27053, n36482);
  and g60525 (n36505, pi0039, n_27053);
  not g60526 (n_27054, n36504);
  and g60527 (n36506, n_27054, n36505);
  not g60528 (n_27055, n36409);
  and g60529 (n36507, n_161, n_27055);
  not g60530 (n_27056, n36506);
  and g60531 (n36508, n_27056, n36507);
  not g60532 (n_27057, n36403);
  and g60533 (n36509, n2571, n_27057);
  not g60534 (n_27058, n36508);
  and g60535 (n36510, n_27058, n36509);
  not g60536 (n_27059, n36510);
  and g60537 (n36511, n_26943, n_27059);
  not g60538 (n_27060, n36511);
  and g60539 (n36512, n_11960, n_27060);
  and g60540 (n36513, n17117, n36259);
  not g60541 (n_27061, n36512);
  not g60542 (n_27062, n36513);
  and g60543 (n36514, n_27061, n_27062);
  not g60544 (n_27063, n36514);
  and g60545 (n36515, n_11964, n_27063);
  and g60546 (n36516, pi0609, n36514);
  and g60547 (n36517, n_11971, n_26870);
  not g60548 (n_27064, n36517);
  and g60549 (n36518, pi1155, n_27064);
  not g60550 (n_27065, n36516);
  and g60551 (n36519, n_27065, n36518);
  and g60552 (n36520, n_11971, n36514);
  and g60553 (n36521, pi0609, n_26870);
  not g60554 (n_27066, n36521);
  and g60555 (n36522, n_11768, n_27066);
  not g60556 (n_27067, n36520);
  and g60557 (n36523, n_27067, n36522);
  not g60558 (n_27068, n36519);
  not g60559 (n_27069, n36523);
  and g60560 (n36524, n_27068, n_27069);
  not g60561 (n_27070, n36524);
  and g60562 (n36525, pi0785, n_27070);
  not g60563 (n_27071, n36515);
  not g60564 (n_27072, n36525);
  and g60565 (n36526, n_27071, n_27072);
  not g60566 (n_27073, n36526);
  and g60567 (n36527, n_11981, n_27073);
  and g60568 (n36528, pi0618, n36526);
  and g60569 (n36529, n_11984, n_26870);
  not g60570 (n_27074, n36529);
  and g60571 (n36530, pi1154, n_27074);
  not g60572 (n_27075, n36528);
  and g60573 (n36531, n_27075, n36530);
  and g60574 (n36532, n_11984, n36526);
  and g60575 (n36533, pi0618, n_26870);
  not g60576 (n_27076, n36533);
  and g60577 (n36534, n_11413, n_27076);
  not g60578 (n_27077, n36532);
  and g60579 (n36535, n_27077, n36534);
  not g60580 (n_27078, n36531);
  not g60581 (n_27079, n36535);
  and g60582 (n36536, n_27078, n_27079);
  not g60583 (n_27080, n36536);
  and g60584 (n36537, pi0781, n_27080);
  not g60585 (n_27081, n36527);
  not g60586 (n_27082, n36537);
  and g60587 (n36538, n_27081, n_27082);
  not g60588 (n_27083, n36538);
  and g60589 (n36539, n_12315, n_27083);
  and g60590 (n36540, pi0619, n36538);
  and g60591 (n36541, n_11821, n_26870);
  not g60592 (n_27084, n36541);
  and g60593 (n36542, pi1159, n_27084);
  not g60594 (n_27085, n36540);
  and g60595 (n36543, n_27085, n36542);
  and g60596 (n36544, n_11821, n36538);
  and g60597 (n36545, pi0619, n_26870);
  not g60598 (n_27086, n36545);
  and g60599 (n36546, n_11405, n_27086);
  not g60600 (n_27087, n36544);
  and g60601 (n36547, n_27087, n36546);
  not g60602 (n_27088, n36543);
  not g60603 (n_27089, n36547);
  and g60604 (n36548, n_27088, n_27089);
  not g60605 (n_27090, n36548);
  and g60606 (n36549, pi0789, n_27090);
  not g60607 (n_27091, n36539);
  not g60608 (n_27092, n36549);
  and g60609 (n36550, n_27091, n_27092);
  and g60610 (n36551, n_12524, n36550);
  not g60611 (n_27093, n36401);
  not g60612 (n_27094, n36551);
  and g60613 (n36552, n_27093, n_27094);
  and g60614 (n36553, n_14557, n36552);
  and g60615 (n36554, n_11789, n_26870);
  and g60616 (n36555, pi0628, n_26963);
  not g60617 (n_27095, n36554);
  and g60618 (n36556, n17776, n_27095);
  not g60619 (n_27096, n36555);
  and g60620 (n36557, n_27096, n36556);
  not g60621 (n_27097, n36400);
  not g60622 (n_27098, n36557);
  and g60623 (n36558, n_27097, n_27098);
  not g60624 (n_27099, n36553);
  and g60625 (n36559, n_27099, n36558);
  not g60626 (n_27100, n36559);
  and g60627 (n36560, pi0792, n_27100);
  and g60628 (n36561, pi0609, n36371);
  and g60629 (n36562, n16667, n17493);
  and g60630 (n36563, n_226, n_3091);
  and g60631 (n36564, n_162, pi0616);
  and g60632 (n36565, n36266, n36564);
  not g60633 (n_27101, n36563);
  not g60634 (n_27102, n36565);
  and g60635 (n36566, n_27101, n_27102);
  not g60636 (n_27103, n36566);
  and g60637 (n36567, n36562, n_27103);
  and g60638 (n36568, n_26873, n_26995);
  and g60639 (n36569, n_3091, n_12023);
  not g60640 (n_27104, n36568);
  not g60641 (n_27105, n36569);
  and g60642 (n36570, n_27104, n_27105);
  and g60643 (n36571, n16641, n36570);
  not g60644 (n_27106, n36571);
  and g60645 (n36572, n_26871, n_27106);
  not g60646 (n_27107, n36567);
  not g60647 (n_27108, n36572);
  and g60648 (n36573, n_27107, n_27108);
  not g60649 (n_27109, n36573);
  and g60650 (n36574, pi0038, n_27109);
  and g60651 (n36575, n_3096, pi0681);
  and g60652 (n36576, n_26994, n36575);
  and g60653 (n36577, n_11502, n36425);
  not g60654 (n_27110, n17504);
  and g60655 (n36578, pi0616, n_27110);
  not g60656 (n_27111, n36578);
  and g60657 (n36579, pi0680, n_27111);
  and g60658 (n36580, n_12016, n36579);
  not g60659 (n_27112, n36577);
  and g60660 (n36581, pi0661, n_27112);
  not g60661 (n_27113, n36580);
  and g60662 (n36582, n_27113, n36581);
  not g60663 (n_27114, n36576);
  and g60664 (n36583, n_26999, n_27114);
  not g60665 (n_27115, n36582);
  and g60666 (n36584, n_27115, n36583);
  not g60667 (n_27116, n36584);
  and g60668 (n36585, n6242, n_27116);
  and g60669 (n36586, n_26987, n36575);
  and g60670 (n36587, n_11502, n36416);
  and g60671 (n36588, n_12158, n17493);
  not g60672 (n_27117, n36588);
  and g60673 (n36589, pi0616, n_27117);
  not g60674 (n_27118, n36589);
  and g60675 (n36590, pi0680, n_27118);
  and g60676 (n36591, n17330, n36590);
  not g60677 (n_27119, n36591);
  and g60678 (n36592, pi0661, n_27119);
  not g60679 (n_27120, n36587);
  and g60680 (n36593, n_27120, n36592);
  not g60681 (n_27121, n36586);
  and g60682 (n36594, n_26991, n_27121);
  not g60683 (n_27122, n36593);
  and g60684 (n36595, n_27122, n36594);
  not g60685 (n_27123, n36595);
  and g60686 (n36596, n_3162, n_27123);
  not g60687 (n_27124, n36585);
  and g60688 (n36597, pi0222, n_27124);
  not g60689 (n_27125, n36596);
  and g60690 (n36598, n_27125, n36597);
  and g60691 (n36599, n17444, n36266);
  not g60692 (n_27126, n36412);
  not g60693 (n_27127, n36599);
  and g60694 (n36600, n_27126, n_27127);
  not g60695 (n_27128, n36600);
  and g60696 (n36601, n6242, n_27128);
  and g60697 (n36602, pi0616, n17237);
  not g60698 (n_27129, n36602);
  and g60699 (n36603, n_3096, n_27129);
  and g60700 (n36604, n_11479, n36439);
  not g60701 (n_27130, n36604);
  and g60702 (n36605, n6195, n_27130);
  and g60703 (n36606, n_11502, n36602);
  not g60704 (n_27131, n17559);
  and g60705 (n36607, n_11999, n_27131);
  and g60706 (n36608, pi0616, n36607);
  not g60707 (n_27132, n36608);
  and g60708 (n36609, pi0680, n_27132);
  and g60709 (n36610, n17458, n36609);
  not g60710 (n_27133, n36606);
  and g60711 (n36611, pi0661, n_27133);
  not g60712 (n_27134, n36610);
  and g60713 (n36612, n_27134, n36611);
  not g60714 (n_27135, n36603);
  not g60715 (n_27136, n36605);
  and g60716 (n36613, n_27135, n_27136);
  not g60717 (n_27137, n36612);
  and g60718 (n36614, n_27137, n36613);
  and g60719 (n36615, n_3162, n36614);
  not g60720 (n_27138, n36601);
  and g60721 (n36616, n_226, n_27138);
  not g60722 (n_27139, n36615);
  and g60723 (n36617, n_27139, n36616);
  not g60724 (n_27140, n36617);
  and g60725 (n36618, pi0215, n_27140);
  not g60726 (n_27141, n36598);
  and g60727 (n36619, n_27141, n36618);
  not g60728 (n_27142, n17548);
  and g60729 (n36620, pi0616, n_27142);
  and g60730 (n36621, n_3091, n_12066);
  not g60731 (n_27143, n36620);
  not g60732 (n_27144, n36621);
  and g60733 (n36622, n_27143, n_27144);
  and g60734 (n36623, n_27104, n36622);
  not g60735 (n_27145, n36623);
  and g60736 (n36624, n36337, n_27145);
  and g60737 (n36625, n_27013, n36575);
  and g60738 (n36626, pi0603, n16681);
  and g60739 (n36627, n6197, n16754);
  not g60740 (n_27146, n36627);
  and g60741 (n36628, n_11998, n_27146);
  and g60742 (n36629, n_11512, n36628);
  not g60743 (n_27147, n36626);
  and g60744 (n36630, n_12033, n_27147);
  not g60745 (n_27148, n36629);
  and g60746 (n36631, n_27148, n36630);
  and g60747 (n36632, n_3087, n36631);
  and g60748 (n36633, n_12200, n36628);
  not g60749 (n_27149, n36633);
  and g60750 (n36634, pi0642, n_27149);
  not g60751 (n_27150, n36632);
  and g60752 (n36635, n6191, n_27150);
  not g60753 (n_27151, n36634);
  and g60754 (n36636, n_27151, n36635);
  and g60755 (n36637, n17452, n36633);
  not g60756 (n_27152, n36628);
  and g60757 (n36638, n17493, n_27152);
  not g60758 (n_27153, n36638);
  and g60759 (n36639, pi0616, n_27153);
  not g60764 (n_27156, n36636);
  and g60766 (n36643, n_11502, n36451);
  not g60767 (n_27157, n36642);
  and g60768 (n36644, pi0661, n_27157);
  not g60769 (n_27158, n36643);
  and g60770 (n36645, n_27158, n36644);
  not g60771 (n_27159, n36625);
  and g60772 (n36646, n_27019, n_27159);
  not g60773 (n_27160, n36645);
  and g60774 (n36647, n_27160, n36646);
  not g60775 (n_27161, n36647);
  and g60776 (n36648, n_3162, n_27161);
  and g60777 (n36649, n_27006, n36575);
  and g60778 (n36650, n_11502, n36441);
  and g60779 (n36651, n_12030, n36579);
  not g60780 (n_27162, n36650);
  and g60781 (n36652, pi0661, n_27162);
  not g60782 (n_27163, n36651);
  and g60783 (n36653, n_27163, n36652);
  not g60784 (n_27164, n36649);
  and g60785 (n36654, n_27010, n_27164);
  not g60786 (n_27165, n36653);
  and g60787 (n36655, n_27165, n36654);
  not g60788 (n_27166, n36655);
  and g60789 (n36656, n6242, n_27166);
  not g60790 (n_27167, n36656);
  and g60791 (n36657, pi0222, n_27167);
  not g60792 (n_27168, n36648);
  and g60793 (n36658, n_27168, n36657);
  and g60794 (n36659, n_27024, n36575);
  and g60795 (n36660, n_11502, n36466);
  and g60796 (n36661, pi0616, n17578);
  not g60797 (n_27169, n36661);
  and g60798 (n36662, pi0680, n_27169);
  and g60799 (n36663, n_12087, n36662);
  not g60800 (n_27170, n36660);
  and g60801 (n36664, pi0661, n_27170);
  not g60802 (n_27171, n36663);
  and g60803 (n36665, n_27171, n36664);
  not g60804 (n_27172, n36659);
  and g60805 (n36666, n_27028, n_27172);
  not g60806 (n_27173, n36665);
  and g60807 (n36667, n_27173, n36666);
  and g60808 (n36668, n_3162, n36667);
  and g60809 (n36669, n_11675, n36439);
  and g60810 (n36670, n17246, n36468);
  not g60811 (n_27174, n36669);
  and g60812 (n36671, n16656, n_27174);
  not g60813 (n_27175, n36670);
  and g60814 (n36672, n_27175, n36671);
  and g60815 (n36673, n_27005, n36575);
  and g60816 (n36674, n_11502, n36439);
  and g60817 (n36675, pi0680, n_12073);
  and g60818 (n36676, n_27143, n36675);
  not g60819 (n_27176, n36674);
  and g60820 (n36677, pi0661, n_27176);
  not g60821 (n_27177, n36676);
  and g60822 (n36678, n_27177, n36677);
  not g60823 (n_27178, n36672);
  not g60824 (n_27179, n36673);
  and g60825 (n36679, n_27178, n_27179);
  not g60826 (n_27180, n36678);
  and g60827 (n36680, n_27180, n36679);
  and g60828 (n36681, n6242, n36680);
  not g60829 (n_27181, n36681);
  and g60830 (n36682, n_226, n_27181);
  not g60831 (n_27182, n36668);
  and g60832 (n36683, n_27182, n36682);
  not g60833 (n_27183, n36658);
  not g60834 (n_27184, n36683);
  and g60835 (n36684, n_27183, n_27184);
  not g60836 (n_27185, n36684);
  and g60837 (n36685, n_9350, n_27185);
  not g60838 (n_27186, n36624);
  and g60839 (n36686, n_36, n_27186);
  not g60840 (n_27187, n36685);
  and g60841 (n36687, n_27187, n36686);
  not g60842 (n_27188, n36619);
  and g60843 (n36688, pi0299, n_27188);
  not g60844 (n_27189, n36687);
  and g60845 (n36689, n_27189, n36688);
  not g60846 (n_27190, n36622);
  and g60847 (n36690, n36266, n_27190);
  and g60848 (n36691, n_26873, n_27005);
  not g60849 (n_27191, n36691);
  and g60850 (n36692, n_226, n_27191);
  not g60851 (n_27192, n36690);
  and g60852 (n36693, n_27192, n36692);
  not g60853 (n_27193, n3351);
  not g60854 (n_27194, n36693);
  and g60855 (n36694, n_27193, n_27194);
  and g60856 (n36695, n_3119, n36667);
  and g60857 (n36696, n6205, n36680);
  not g60858 (n_27195, n36696);
  and g60859 (n36697, pi0224, n_27195);
  not g60860 (n_27196, n36695);
  and g60861 (n36698, n_27196, n36697);
  not g60862 (n_27197, n36694);
  not g60863 (n_27198, n36698);
  and g60864 (n36699, n_27197, n_27198);
  and g60865 (n36700, n6205, n36655);
  and g60866 (n36701, n_3119, n36647);
  not g60867 (n_27199, n36700);
  and g60868 (n36702, pi0222, n_27199);
  not g60869 (n_27200, n36701);
  and g60870 (n36703, n_27200, n36702);
  not g60871 (n_27201, n36699);
  not g60872 (n_27202, n36703);
  and g60873 (n36704, n_27201, n_27202);
  not g60874 (n_27203, n36704);
  and g60875 (n36705, n_223, n_27203);
  and g60876 (n36706, n6205, n_27116);
  and g60877 (n36707, n_3119, n_27123);
  not g60878 (n_27204, n36706);
  and g60879 (n36708, pi0222, n_27204);
  not g60880 (n_27205, n36707);
  and g60881 (n36709, n_27205, n36708);
  and g60882 (n36710, n6205, n_27128);
  and g60883 (n36711, n_3119, n36614);
  not g60884 (n_27206, n36710);
  and g60885 (n36712, n_226, n_27206);
  not g60886 (n_27207, n36711);
  and g60887 (n36713, n_27207, n36712);
  not g60888 (n_27208, n36713);
  and g60889 (n36714, pi0223, n_27208);
  not g60890 (n_27209, n36709);
  and g60891 (n36715, n_27209, n36714);
  not g60892 (n_27210, n36715);
  and g60893 (n36716, n_234, n_27210);
  not g60894 (n_27211, n36705);
  and g60895 (n36717, n_27211, n36716);
  not g60896 (n_27212, n36717);
  and g60897 (n36718, pi0039, n_27212);
  not g60898 (n_27213, n36689);
  and g60899 (n36719, n_27213, n36718);
  and g60900 (n36720, pi0661, n17618);
  and g60901 (n36721, pi0616, n17226);
  not g60902 (n_27214, n36721);
  and g60903 (n36722, n_226, n_27214);
  not g60904 (n_27215, n36720);
  and g60905 (n36723, n_27215, n36722);
  and g60906 (n36724, n_3091, n17226);
  and g60907 (n36725, n17617, n_26873);
  and g60908 (n36726, n_11512, n_11648);
  not g60909 (n_27216, n17367);
  and g60910 (n36727, n_27216, n_12232);
  not g60911 (n_27217, n36726);
  and g60912 (n36728, n_27217, n36727);
  not g60913 (n_27218, n36724);
  not g60914 (n_27219, n36728);
  and g60915 (n36729, n_27218, n_27219);
  not g60916 (n_27220, n36725);
  and g60917 (n36730, n_27220, n36729);
  not g60918 (n_27221, n36730);
  and g60919 (n36731, pi0222, n_27221);
  not g60920 (n_27222, n36723);
  not g60921 (n_27223, n36731);
  and g60922 (n36732, n_27222, n_27223);
  not g60923 (n_27224, n36732);
  and g60924 (n36733, n_234, n_27224);
  and g60925 (n36734, n_3091, n17231);
  and g60926 (n36735, n17622, n_26873);
  and g60927 (n36736, n_11512, n_11655);
  and g60928 (n36737, n_11833, n_27216);
  not g60929 (n_27225, n36736);
  and g60930 (n36738, n_27225, n36737);
  not g60931 (n_27226, n36734);
  not g60932 (n_27227, n36738);
  and g60933 (n36739, n_27226, n_27227);
  not g60934 (n_27228, n36735);
  and g60935 (n36740, n_27228, n36739);
  not g60936 (n_27229, n36740);
  and g60937 (n36741, pi0222, n_27229);
  and g60938 (n36742, pi0661, n17623);
  and g60939 (n36743, pi0616, n17231);
  not g60940 (n_27230, n36743);
  and g60941 (n36744, n_226, n_27230);
  not g60942 (n_27231, n36742);
  and g60943 (n36745, n_27231, n36744);
  not g60944 (n_27232, n36741);
  not g60945 (n_27233, n36745);
  and g60946 (n36746, n_27232, n_27233);
  not g60947 (n_27234, n36746);
  and g60948 (n36747, pi0299, n_27234);
  not g60949 (n_27235, n36733);
  and g60950 (n36748, n_162, n_27235);
  not g60951 (n_27236, n36747);
  and g60952 (n36749, n_27236, n36748);
  not g60953 (n_27237, n36749);
  and g60954 (n36750, n_161, n_27237);
  not g60955 (n_27238, n36719);
  and g60956 (n36751, n_27238, n36750);
  not g60957 (n_27239, n36574);
  and g60958 (n36752, n2571, n_27239);
  not g60959 (n_27240, n36751);
  and g60960 (n36753, n_27240, n36752);
  not g60961 (n_27241, n36753);
  and g60962 (n36754, n_26943, n_27241);
  and g60963 (n36755, n_11753, n36754);
  and g60964 (n36756, pi0625, n36511);
  not g60965 (n_27242, n36756);
  and g60966 (n36757, n_11757, n_27242);
  not g60967 (n_27243, n36755);
  and g60968 (n36758, n_27243, n36757);
  and g60969 (n36759, n_11823, n_26950);
  not g60970 (n_27244, n36758);
  and g60971 (n36760, n_27244, n36759);
  and g60972 (n36761, n_11753, n36511);
  and g60973 (n36762, pi0625, n36754);
  not g60974 (n_27245, n36761);
  and g60975 (n36763, pi1153, n_27245);
  not g60976 (n_27246, n36762);
  and g60977 (n36764, n_27246, n36763);
  and g60978 (n36765, pi0608, n_26951);
  not g60979 (n_27247, n36764);
  and g60980 (n36766, n_27247, n36765);
  not g60981 (n_27248, n36760);
  not g60982 (n_27249, n36766);
  and g60983 (n36767, n_27248, n_27249);
  not g60984 (n_27250, n36767);
  and g60985 (n36768, pi0778, n_27250);
  and g60986 (n36769, n_11749, n36754);
  not g60987 (n_27251, n36768);
  not g60988 (n_27252, n36769);
  and g60989 (n36770, n_27251, n_27252);
  not g60990 (n_27253, n36770);
  and g60991 (n36771, n_11971, n_27253);
  not g60992 (n_27254, n36561);
  and g60993 (n36772, n_11768, n_27254);
  not g60994 (n_27255, n36771);
  and g60995 (n36773, n_27255, n36772);
  and g60996 (n36774, n_11767, n_27068);
  not g60997 (n_27256, n36773);
  and g60998 (n36775, n_27256, n36774);
  and g60999 (n36776, n_11971, n36371);
  and g61000 (n36777, pi0609, n_27253);
  not g61001 (n_27257, n36776);
  and g61002 (n36778, pi1155, n_27257);
  not g61003 (n_27258, n36777);
  and g61004 (n36779, n_27258, n36778);
  and g61005 (n36780, pi0660, n_27069);
  not g61006 (n_27259, n36779);
  and g61007 (n36781, n_27259, n36780);
  not g61008 (n_27260, n36775);
  not g61009 (n_27261, n36781);
  and g61010 (n36782, n_27260, n_27261);
  not g61011 (n_27262, n36782);
  and g61012 (n36783, pi0785, n_27262);
  and g61013 (n36784, n_11964, n_27253);
  not g61014 (n_27263, n36783);
  not g61015 (n_27264, n36784);
  and g61016 (n36785, n_27263, n_27264);
  not g61017 (n_27265, n36785);
  and g61018 (n36786, n_11984, n_27265);
  and g61019 (n36787, pi0618, n36374);
  not g61020 (n_27266, n36787);
  and g61021 (n36788, n_11413, n_27266);
  not g61022 (n_27267, n36786);
  and g61023 (n36789, n_27267, n36788);
  and g61024 (n36790, n_11412, n_27078);
  not g61025 (n_27268, n36789);
  and g61026 (n36791, n_27268, n36790);
  and g61027 (n36792, n_11984, n36374);
  and g61028 (n36793, pi0618, n_27265);
  not g61029 (n_27269, n36792);
  and g61030 (n36794, pi1154, n_27269);
  not g61031 (n_27270, n36793);
  and g61032 (n36795, n_27270, n36794);
  and g61033 (n36796, pi0627, n_27079);
  not g61034 (n_27271, n36795);
  and g61035 (n36797, n_27271, n36796);
  not g61036 (n_27272, n36791);
  not g61037 (n_27273, n36797);
  and g61038 (n36798, n_27272, n_27273);
  not g61039 (n_27274, n36798);
  and g61040 (n36799, pi0781, n_27274);
  and g61041 (n36800, n_11981, n_27265);
  not g61042 (n_27275, n36799);
  not g61043 (n_27276, n36800);
  and g61044 (n36801, n_27275, n_27276);
  and g61045 (n36802, n_12315, n36801);
  and g61046 (n36803, n_12320, n36550);
  and g61047 (n36804, pi0626, n_26870);
  not g61048 (n_27277, n36804);
  and g61049 (n36805, n16629, n_27277);
  not g61050 (n_27278, n36803);
  and g61051 (n36806, n_27278, n36805);
  and g61052 (n36807, n16635, n_26870);
  not g61053 (n_27279, n36807);
  and g61054 (n36808, n17871, n_27279);
  not g61055 (n_27280, n36378);
  and g61056 (n36809, n_27280, n36808);
  and g61057 (n36810, pi0626, n36550);
  and g61058 (n36811, n_12320, n_26870);
  not g61059 (n_27281, n36811);
  and g61060 (n36812, n16628, n_27281);
  not g61061 (n_27282, n36810);
  and g61062 (n36813, n_27282, n36812);
  not g61063 (n_27283, n36806);
  not g61064 (n_27284, n36809);
  and g61065 (n36814, n_27283, n_27284);
  not g61066 (n_27285, n36813);
  and g61067 (n36815, n_27285, n36814);
  not g61068 (n_27286, n36815);
  and g61069 (n36816, pi0788, n_27286);
  not g61070 (n_27287, n36801);
  and g61071 (n36817, n_11821, n_27287);
  and g61072 (n36818, pi0619, n36377);
  not g61073 (n_27288, n36818);
  and g61074 (n36819, n_11405, n_27288);
  not g61075 (n_27289, n36817);
  and g61076 (n36820, n_27289, n36819);
  and g61077 (n36821, n_11403, n_27088);
  not g61078 (n_27290, n36820);
  and g61079 (n36822, n_27290, n36821);
  and g61080 (n36823, pi0619, n_27287);
  and g61081 (n36824, n_11821, n36377);
  not g61082 (n_27291, n36824);
  and g61083 (n36825, pi1159, n_27291);
  not g61084 (n_27292, n36823);
  and g61085 (n36826, n_27292, n36825);
  and g61086 (n36827, pi0648, n_27089);
  not g61087 (n_27293, n36826);
  and g61088 (n36828, n_27293, n36827);
  not g61089 (n_27294, n36822);
  and g61090 (n36829, pi0789, n_27294);
  not g61091 (n_27295, n36828);
  and g61092 (n36830, n_27295, n36829);
  not g61093 (n_27296, n36802);
  not g61094 (n_27297, n36816);
  and g61095 (n36831, n_27296, n_27297);
  not g61096 (n_27298, n36830);
  and g61097 (n36832, n_27298, n36831);
  not g61098 (n_27299, n17970);
  and g61099 (n36833, n_27299, n36815);
  not g61100 (n_27300, n36833);
  and g61101 (n36834, n_14638, n_27300);
  not g61102 (n_27301, n36832);
  and g61103 (n36835, n_27301, n36834);
  not g61104 (n_27302, n36560);
  not g61105 (n_27303, n36835);
  and g61106 (n36836, n_27302, n_27303);
  not g61107 (n_27304, n36836);
  and g61108 (n36837, n_14387, n_27304);
  and g61109 (n36838, n_12375, n36392);
  and g61110 (n36839, n_12368, n36552);
  and g61111 (n36840, n17779, n36259);
  not g61112 (n_27305, n36839);
  not g61113 (n_27306, n36840);
  and g61114 (n36841, n_27305, n_27306);
  not g61115 (n_27307, n36841);
  and g61116 (n36842, n_14548, n_27307);
  and g61117 (n36843, pi0630, n36388);
  not g61118 (n_27308, n36838);
  not g61119 (n_27309, n36843);
  and g61120 (n36844, n_27308, n_27309);
  not g61121 (n_27310, n36842);
  and g61122 (n36845, n_27310, n36844);
  not g61123 (n_27311, n36845);
  and g61124 (n36846, pi0787, n_27311);
  not g61125 (n_27312, n36837);
  not g61126 (n_27313, n36846);
  and g61127 (n36847, n_27312, n_27313);
  and g61128 (n36848, pi0644, n36847);
  not g61129 (n_27314, n36396);
  and g61130 (n36849, pi0715, n_27314);
  not g61131 (n_27315, n36848);
  and g61132 (n36850, n_27315, n36849);
  and g61133 (n36851, n17804, n_26870);
  and g61134 (n36852, n_12392, n36841);
  not g61135 (n_27316, n36851);
  not g61136 (n_27317, n36852);
  and g61137 (n36853, n_27316, n_27317);
  not g61138 (n_27318, n36853);
  and g61139 (n36854, pi0644, n_27318);
  and g61140 (n36855, n_11819, n_26870);
  not g61141 (n_27319, n36855);
  and g61142 (n36856, n_12395, n_27319);
  not g61143 (n_27320, n36854);
  and g61144 (n36857, n_27320, n36856);
  not g61145 (n_27321, n36857);
  and g61146 (n36858, pi1160, n_27321);
  not g61147 (n_27322, n36850);
  and g61148 (n36859, n_27322, n36858);
  and g61149 (n36860, pi0644, n36395);
  and g61150 (n36861, n_11819, n36847);
  not g61151 (n_27323, n36860);
  and g61152 (n36862, n_12395, n_27323);
  not g61153 (n_27324, n36861);
  and g61154 (n36863, n_27324, n36862);
  and g61155 (n36864, n_11819, n_27318);
  and g61156 (n36865, pi0644, n_26870);
  not g61157 (n_27325, n36865);
  and g61158 (n36866, pi0715, n_27325);
  not g61159 (n_27326, n36864);
  and g61160 (n36867, n_27326, n36866);
  not g61161 (n_27327, n36867);
  and g61162 (n36868, n_12405, n_27327);
  not g61163 (n_27328, n36863);
  and g61164 (n36869, n_27328, n36868);
  not g61165 (n_27329, n36859);
  not g61166 (n_27330, n36869);
  and g61167 (n36870, n_27329, n_27330);
  not g61168 (n_27331, n36870);
  and g61169 (n36871, pi0790, n_27331);
  and g61170 (n36872, n_12411, n36847);
  not g61171 (n_27332, n36871);
  not g61172 (n_27333, n36872);
  and g61173 (n36873, n_27332, n_27333);
  not g61174 (n_27334, n36873);
  and g61175 (n36874, n_4226, n_27334);
  and g61176 (n36875, n_226, po1038);
  not g61177 (n_27335, n36874);
  not g61178 (n_27336, n36875);
  and g61179 (po0379, n_27335, n_27336);
  and g61180 (n36877, n_234, n_11697);
  not g61181 (n_27337, n36877);
  and g61182 (n36878, pi0039, n_27337);
  and g61183 (n36879, n_11735, n36878);
  and g61184 (n36880, n14873, n_12667);
  not g61185 (n_27338, n36879);
  and g61186 (n36881, n_27338, n36880);
  not g61187 (n_27339, n36881);
  and g61188 (n36882, n18591, n_27339);
  not g61189 (n_27340, n36882);
  and g61190 (n36883, pi0223, n_27340);
  not g61191 (n_27341, n36883);
  and g61192 (n36884, n_24651, n_27341);
  and g61193 (n36885, n17075, n_27341);
  and g61194 (n36886, pi0223, n_11417);
  and g61195 (n36887, pi0680, pi0681);
  not g61196 (n_27342, n36887);
  and g61197 (n36888, n16918, n_27342);
  and g61198 (n36889, n_223, n_12231);
  and g61199 (n36890, pi0223, n16935);
  and g61206 (n36894, pi0223, n16944);
  and g61207 (n36895, n16923, n_27342);
  and g61208 (n36896, n_223, n_12235);
  not g61215 (n_27349, n36893);
  and g61216 (n36900, n_162, n_27349);
  not g61217 (n_27350, n36899);
  and g61218 (n36901, n_27350, n36900);
  and g61219 (n36902, pi0681, n16739);
  not g61220 (n_27351, n36902);
  and g61221 (n36903, n2603, n_27351);
  and g61222 (n36904, n_26895, n36887);
  and g61223 (n36905, n6205, n36904);
  and g61224 (n36906, pi0681, n16703);
  and g61225 (n36907, n_3119, n36906);
  not g61226 (n_27352, n36905);
  and g61227 (n36908, n_9349, n_27352);
  not g61228 (n_27353, n36907);
  and g61229 (n36909, n_27353, n36908);
  not g61230 (n_27354, n36903);
  not g61231 (n_27355, n36909);
  and g61232 (n36910, n_27354, n_27355);
  not g61233 (n_27356, n36910);
  and g61234 (n36911, n_223, n_27356);
  and g61235 (n36912, pi0681, n_26907);
  not g61236 (n_27357, n36912);
  and g61237 (n36913, n_11693, n_27357);
  not g61238 (n_27358, n36913);
  and g61239 (n36914, n6205, n_27358);
  and g61240 (n36915, pi0681, n_26903);
  not g61241 (n_27359, n36915);
  and g61242 (n36916, n_11683, n_27359);
  not g61243 (n_27360, n36916);
  and g61244 (n36917, n_3119, n_27360);
  not g61245 (n_27361, n36914);
  and g61246 (n36918, pi0223, n_27361);
  not g61247 (n_27362, n36917);
  and g61248 (n36919, n_27362, n36918);
  not g61249 (n_27363, n36919);
  and g61250 (n36920, n_234, n_27363);
  not g61251 (n_27364, n36911);
  and g61252 (n36921, n_27364, n36920);
  and g61253 (n36922, n_223, pi0681);
  and g61254 (n36923, n16744, n36922);
  and g61255 (n36924, n6242, n36913);
  and g61256 (n36925, n_3162, n36916);
  not g61257 (n_27365, n36924);
  and g61258 (n36926, pi0223, n_27365);
  not g61259 (n_27366, n36925);
  and g61260 (n36927, n_27366, n36926);
  not g61261 (n_27367, n36923);
  and g61262 (n36928, pi0215, n_27367);
  not g61263 (n_27368, n36927);
  and g61264 (n36929, n_27368, n36928);
  and g61265 (n36930, pi0223, n_11445);
  not g61266 (n_27369, n36930);
  and g61267 (n36931, n3448, n_27369);
  and g61268 (n36932, n_27351, n36931);
  and g61269 (n36933, pi0681, n_26883);
  and g61270 (n36934, n_3162, n_11711);
  not g61271 (n_27370, n36933);
  and g61272 (n36935, n_27370, n36934);
  and g61273 (n36936, pi0681, n_26889);
  and g61274 (n36937, n6242, n_11705);
  not g61275 (n_27371, n36936);
  and g61276 (n36938, n_27371, n36937);
  not g61277 (n_27372, n36935);
  and g61278 (n36939, pi0223, n_27372);
  not g61279 (n_27373, n36938);
  and g61280 (n36940, n_27373, n36939);
  not g61281 (n_27374, n36906);
  and g61282 (n36941, n_3162, n_27374);
  not g61283 (n_27375, n36904);
  and g61284 (n36942, n6242, n_27375);
  not g61285 (n_27376, n36941);
  and g61286 (n36943, n_223, n_27376);
  not g61287 (n_27377, n36942);
  and g61288 (n36944, n_27377, n36943);
  not g61289 (n_27378, n36944);
  and g61290 (n36945, n_9350, n_27378);
  not g61291 (n_27379, n36940);
  and g61292 (n36946, n_27379, n36945);
  not g61293 (n_27380, n36932);
  not g61294 (n_27381, n36946);
  and g61295 (n36947, n_27380, n_27381);
  not g61296 (n_27382, n36947);
  and g61297 (n36948, n_36, n_27382);
  not g61298 (n_27383, n36929);
  and g61299 (n36949, pi0299, n_27383);
  not g61300 (n_27384, n36948);
  and g61301 (n36950, n_27384, n36949);
  not g61302 (n_27385, n36921);
  and g61303 (n36951, pi0039, n_27385);
  not g61304 (n_27386, n36950);
  and g61305 (n36952, n_27386, n36951);
  not g61306 (n_27387, n36901);
  not g61307 (n_27388, n36952);
  and g61308 (n36953, n_27387, n_27388);
  not g61309 (n_27389, n36953);
  and g61310 (n36954, n_161, n_27389);
  and g61311 (n36955, pi0681, n16646);
  and g61312 (n36956, pi0223, n_11418);
  not g61313 (n_27390, n36955);
  and g61314 (n36957, pi0038, n_27390);
  not g61315 (n_27391, n36956);
  and g61316 (n36958, n_27391, n36957);
  not g61317 (n_27392, n36958);
  and g61318 (n36959, n2571, n_27392);
  not g61319 (n_27393, n36954);
  and g61320 (n36960, n_27393, n36959);
  not g61321 (n_27394, n36886);
  not g61322 (n_27395, n36960);
  and g61323 (n36961, n_27394, n_27395);
  not g61324 (n_27396, n36961);
  and g61325 (n36962, n_11749, n_27396);
  and g61326 (n36963, pi0625, n36961);
  and g61327 (n36964, n_11753, n_27341);
  not g61328 (n_27397, n36964);
  and g61329 (n36965, pi1153, n_27397);
  not g61330 (n_27398, n36963);
  and g61331 (n36966, n_27398, n36965);
  and g61332 (n36967, n_11753, n36961);
  and g61333 (n36968, pi0625, n_27341);
  not g61334 (n_27399, n36968);
  and g61335 (n36969, n_11757, n_27399);
  not g61336 (n_27400, n36967);
  and g61337 (n36970, n_27400, n36969);
  not g61338 (n_27401, n36966);
  not g61339 (n_27402, n36970);
  and g61340 (n36971, n_27401, n_27402);
  not g61341 (n_27403, n36971);
  and g61342 (n36972, pi0778, n_27403);
  not g61343 (n_27404, n36962);
  not g61344 (n_27405, n36972);
  and g61345 (n36973, n_27404, n_27405);
  and g61346 (n36974, n_11773, n36973);
  not g61347 (n_27406, n36885);
  not g61348 (n_27407, n36974);
  and g61349 (n36975, n_27406, n_27407);
  and g61350 (n36976, n_11777, n36975);
  and g61351 (n36977, n16639, n36883);
  not g61352 (n_27408, n36976);
  not g61353 (n_27409, n36977);
  and g61354 (n36978, n_27408, n_27409);
  and g61355 (n36979, n_11780, n36978);
  and g61356 (n36980, n_11783, n36979);
  not g61357 (n_27410, n36884);
  not g61358 (n_27411, n36980);
  and g61359 (n36981, n_27410, n_27411);
  not g61360 (n_27412, n36981);
  and g61361 (n36982, n_13453, n_27412);
  and g61362 (n36983, n17856, n_27341);
  not g61363 (n_27413, n36982);
  not g61364 (n_27414, n36983);
  and g61365 (n36984, n_27413, n_27414);
  and g61366 (n36985, n_11803, n36984);
  not g61367 (n_27415, n36984);
  and g61368 (n36986, n_11806, n_27415);
  and g61369 (n36987, pi0647, n_27341);
  not g61370 (n_27416, n36987);
  and g61371 (n36988, n_11810, n_27416);
  not g61372 (n_27417, n36986);
  and g61373 (n36989, n_27417, n36988);
  and g61374 (n36990, pi0647, n_27415);
  and g61375 (n36991, n_11806, n_27341);
  not g61376 (n_27418, n36991);
  and g61377 (n36992, pi1157, n_27418);
  not g61378 (n_27419, n36990);
  and g61379 (n36993, n_27419, n36992);
  not g61380 (n_27420, n36989);
  not g61381 (n_27421, n36993);
  and g61382 (n36994, n_27420, n_27421);
  not g61383 (n_27422, n36994);
  and g61384 (n36995, pi0787, n_27422);
  not g61385 (n_27423, n36985);
  not g61386 (n_27424, n36995);
  and g61387 (n36996, n_27423, n_27424);
  and g61388 (n36997, n_11819, n36996);
  and g61389 (n36998, n_12375, n36993);
  and g61390 (n36999, n17969, n_27341);
  and g61391 (n37000, n17117, n_27341);
  and g61392 (n37001, pi0039, pi0223);
  not g61393 (n_27425, n37001);
  and g61394 (n37002, pi0038, n_27425);
  and g61395 (n37003, pi0642, n17168);
  not g61396 (n_27426, n37003);
  and g61397 (n37004, n16667, n_27426);
  and g61398 (n37005, n_223, n_11432);
  not g61399 (n_27427, n37005);
  and g61400 (n37006, n_162, n_27427);
  not g61401 (n_27428, n37004);
  and g61402 (n37007, n_27428, n37006);
  not g61403 (n_27429, n37007);
  and g61404 (n37008, n37002, n_27429);
  and g61405 (n37009, n_223, pi0642);
  and g61406 (n37010, n17226, n37009);
  not g61407 (n_27430, n37010);
  and g61408 (n37011, n_234, n_27430);
  and g61409 (n37012, n_3087, n17226);
  not g61410 (n_27431, n37012);
  and g61411 (n37013, pi0223, n_27431);
  and g61412 (n37014, n17137, n37013);
  not g61413 (n_27432, n37014);
  and g61414 (n37015, n37011, n_27432);
  and g61415 (n37016, n17231, n37009);
  not g61416 (n_27433, n37016);
  and g61417 (n37017, pi0299, n_27433);
  and g61418 (n37018, n6190, n17230);
  and g61419 (n37019, pi0223, n_11834);
  not g61420 (n_27434, n37018);
  and g61421 (n37020, n_27434, n37019);
  not g61422 (n_27435, n37020);
  and g61423 (n37021, n37017, n_27435);
  not g61424 (n_27436, n37021);
  and g61425 (n37022, n_162, n_27436);
  not g61426 (n_27437, n37015);
  and g61427 (n37023, n_27437, n37022);
  and g61428 (n37024, n35897, n_27426);
  and g61429 (n37025, pi0642, n_26992);
  not g61430 (n_27438, n37025);
  and g61431 (n37026, n36425, n_27438);
  not g61432 (n_27439, n37024);
  not g61433 (n_27440, n37026);
  and g61434 (n37027, n_27439, n_27440);
  and g61435 (n37028, pi0681, n37027);
  and g61436 (n37029, n6194, n37004);
  and g61437 (n37030, n16797, n37029);
  not g61438 (n_27441, n37027);
  and g61439 (n37031, n_11707, n_27441);
  not g61440 (n_27442, n37030);
  and g61441 (n37032, n_3098, n_27442);
  not g61442 (n_27443, n37031);
  and g61443 (n37033, n_27443, n37032);
  not g61444 (n_27444, n37028);
  not g61445 (n_27445, n37033);
  and g61446 (n37034, n_27444, n_27445);
  and g61447 (n37035, n6205, n37034);
  and g61448 (n37036, n_3087, n_11558);
  not g61449 (n_27446, n17183);
  and g61450 (n37037, pi0642, n_27446);
  not g61451 (n_27447, n37036);
  not g61452 (n_27448, n37037);
  and g61453 (n37038, n_27447, n_27448);
  and g61454 (n37039, n_11707, n37038);
  and g61455 (n37040, pi0642, n_26984);
  not g61456 (n_27449, n37040);
  and g61457 (n37041, n6194, n_27449);
  and g61458 (n37042, n_11479, n37041);
  not g61459 (n_27450, n37042);
  and g61460 (n37043, n_3098, n_27450);
  not g61461 (n_27451, n37039);
  and g61462 (n37044, n_27451, n37043);
  not g61463 (n_27452, n37038);
  and g61464 (n37045, pi0681, n_27452);
  not g61465 (n_27453, n37044);
  not g61466 (n_27454, n37045);
  and g61467 (n37046, n_27453, n_27454);
  and g61468 (n37047, n_3119, n37046);
  not g61469 (n_27455, n37047);
  and g61470 (n37048, pi0223, n_27455);
  not g61471 (n_27456, n37035);
  and g61472 (n37049, n_27456, n37048);
  and g61473 (n37050, pi0642, n17235);
  not g61474 (n_27457, n37050);
  and g61475 (n37051, n2603, n_27457);
  and g61476 (n37052, n_11707, n37050);
  not g61477 (n_27458, n37052);
  and g61478 (n37053, n_3098, n_27458);
  and g61479 (n37054, pi0642, n6194);
  and g61480 (n37055, n17246, n37054);
  not g61481 (n_27459, n37055);
  and g61482 (n37056, n37053, n_27459);
  and g61483 (n37057, pi0681, n_27457);
  not g61484 (n_27460, n37056);
  not g61485 (n_27461, n37057);
  and g61486 (n37058, n_27460, n_27461);
  and g61487 (n37059, n6205, n37058);
  and g61488 (n37060, n_12078, n37003);
  not g61489 (n_27462, n37060);
  and g61490 (n37061, pi0681, n_27462);
  and g61491 (n37062, n17375, n37054);
  and g61492 (n37063, n_11707, n37060);
  not g61493 (n_27463, n37062);
  and g61494 (n37064, n_3098, n_27463);
  not g61495 (n_27464, n37063);
  and g61496 (n37065, n_27464, n37064);
  not g61497 (n_27465, n37061);
  not g61498 (n_27466, n37065);
  and g61499 (n37066, n_27465, n_27466);
  and g61500 (n37067, n_3119, n37066);
  not g61501 (n_27467, n37059);
  and g61502 (n37068, n_9349, n_27467);
  not g61503 (n_27468, n37067);
  and g61504 (n37069, n_27468, n37068);
  not g61505 (n_27469, n37051);
  and g61506 (n37070, n_223, n_27469);
  not g61507 (n_27470, n37069);
  and g61508 (n37071, n_27470, n37070);
  not g61509 (n_27471, n37049);
  and g61510 (n37072, n_234, n_27471);
  not g61511 (n_27472, n37071);
  and g61512 (n37073, n_27472, n37072);
  and g61513 (n37074, n17236, n37054);
  not g61514 (n_27473, n37074);
  and g61515 (n37075, n37053, n_27473);
  and g61516 (n37076, n16723, n37043);
  not g61517 (n_27474, n37075);
  not g61518 (n_27475, n37076);
  and g61519 (n37077, n_27474, n_27475);
  and g61520 (n37078, pi0642, n17237);
  not g61521 (n_27476, n37078);
  and g61522 (n37079, pi0681, n_27476);
  not g61523 (n_27477, n37079);
  and g61524 (n37080, n37077, n_27477);
  not g61525 (n_27478, n37080);
  and g61526 (n37081, pi0947, n_27478);
  and g61527 (n37082, n6242, n_27474);
  and g61528 (n37083, n37050, n37082);
  and g61529 (n37084, n_14829, n37080);
  not g61530 (n_27479, n37083);
  and g61531 (n37085, n_3149, n_27479);
  not g61532 (n_27480, n37084);
  and g61533 (n37086, n_27480, n37085);
  not g61534 (n_27481, n37081);
  and g61535 (n37087, n_223, n_27481);
  not g61536 (n_27482, n37086);
  and g61537 (n37088, n_27482, n37087);
  and g61538 (n37089, n_3162, n37046);
  and g61539 (n37090, n6242, n37034);
  not g61540 (n_27483, n37089);
  and g61541 (n37091, pi0223, n_27483);
  not g61542 (n_27484, n37090);
  and g61543 (n37092, n_27484, n37091);
  not g61544 (n_27485, n37088);
  not g61545 (n_27486, n37092);
  and g61546 (n37093, n_27485, n_27486);
  not g61547 (n_27487, n37093);
  and g61548 (n37094, pi0215, n_27487);
  and g61549 (n37095, n36931, n_27457);
  not g61550 (n_27488, n37066);
  and g61551 (n37096, pi0947, n_27488);
  and g61552 (n37097, n20923, n37058);
  and g61553 (n37098, n_14829, n37066);
  not g61554 (n_27489, n37097);
  and g61555 (n37099, n_3149, n_27489);
  not g61556 (n_27490, n37098);
  and g61557 (n37100, n_27490, n37099);
  not g61558 (n_27491, n37096);
  and g61559 (n37101, n_223, n_27491);
  not g61560 (n_27492, n37100);
  and g61561 (n37102, n_27492, n37101);
  and g61562 (n37103, pi0642, n_11856);
  and g61563 (n37104, n_3087, n_11503);
  not g61564 (n_27493, n37103);
  not g61565 (n_27494, n37104);
  and g61566 (n37105, n_27493, n_27494);
  not g61567 (n_27495, n37105);
  and g61568 (n37106, pi0681, n_27495);
  and g61569 (n37107, n_11707, n37105);
  and g61570 (n37108, n17014, n_27426);
  not g61571 (n_27496, n37108);
  and g61572 (n37109, n_3098, n_27496);
  not g61573 (n_27497, n37107);
  and g61574 (n37110, n_27497, n37109);
  not g61575 (n_27498, n37110);
  and g61576 (n37111, n_3162, n_27498);
  not g61577 (n_27499, n37106);
  and g61578 (n37112, n_27499, n37111);
  and g61579 (n37113, n6191, n_27438);
  and g61580 (n37114, n_11518, n37113);
  not g61581 (n_27500, n37114);
  and g61582 (n37115, n_27439, n_27500);
  and g61583 (n37116, pi0681, n37115);
  not g61584 (n_27501, n37115);
  and g61585 (n37117, n_11707, n_27501);
  and g61586 (n37118, n_11864, n_26591);
  not g61587 (n_27502, n37118);
  and g61588 (n37119, n6194, n_27502);
  not g61589 (n_27503, n37119);
  and g61590 (n37120, n_3098, n_27503);
  not g61591 (n_27504, n37117);
  and g61592 (n37121, n_27504, n37120);
  not g61593 (n_27505, n37121);
  and g61594 (n37122, n6242, n_27505);
  not g61595 (n_27506, n37116);
  and g61596 (n37123, n_27506, n37122);
  not g61597 (n_27507, n37112);
  and g61598 (n37124, pi0223, n_27507);
  not g61599 (n_27508, n37123);
  and g61600 (n37125, n_27508, n37124);
  not g61601 (n_27509, n37102);
  and g61602 (n37126, n_9350, n_27509);
  not g61603 (n_27510, n37125);
  and g61604 (n37127, n_27510, n37126);
  not g61605 (n_27511, n37095);
  and g61606 (n37128, n_36, n_27511);
  not g61607 (n_27512, n37127);
  and g61608 (n37129, n_27512, n37128);
  not g61609 (n_27513, n37094);
  and g61610 (n37130, pi0299, n_27513);
  not g61611 (n_27514, n37129);
  and g61612 (n37131, n_27514, n37130);
  not g61613 (n_27515, n37073);
  and g61614 (n37132, pi0039, n_27515);
  not g61615 (n_27516, n37131);
  and g61616 (n37133, n_27516, n37132);
  not g61617 (n_27517, n37023);
  and g61618 (n37134, n_161, n_27517);
  not g61619 (n_27518, n37133);
  and g61620 (n37135, n_27518, n37134);
  not g61621 (n_27519, n37008);
  and g61622 (n37136, n2571, n_27519);
  not g61623 (n_27520, n37135);
  and g61624 (n37137, n_27520, n37136);
  not g61625 (n_27521, n37137);
  and g61626 (n37138, n_27394, n_27521);
  and g61627 (n37139, n_11960, n37138);
  not g61628 (n_27522, n37000);
  not g61629 (n_27523, n37139);
  and g61630 (n37140, n_27522, n_27523);
  and g61631 (n37141, n_11964, n37140);
  not g61632 (n_27524, n37140);
  and g61633 (n37142, pi0609, n_27524);
  and g61634 (n37143, n_11971, n_27341);
  not g61635 (n_27525, n37143);
  and g61636 (n37144, pi1155, n_27525);
  not g61637 (n_27526, n37142);
  and g61638 (n37145, n_27526, n37144);
  and g61639 (n37146, n_11971, n_27524);
  and g61640 (n37147, pi0609, n_27341);
  not g61641 (n_27527, n37147);
  and g61642 (n37148, n_11768, n_27527);
  not g61643 (n_27528, n37146);
  and g61644 (n37149, n_27528, n37148);
  not g61645 (n_27529, n37145);
  not g61646 (n_27530, n37149);
  and g61647 (n37150, n_27529, n_27530);
  not g61648 (n_27531, n37150);
  and g61649 (n37151, pi0785, n_27531);
  not g61650 (n_27532, n37141);
  not g61651 (n_27533, n37151);
  and g61652 (n37152, n_27532, n_27533);
  not g61653 (n_27534, n37152);
  and g61654 (n37153, n_11981, n_27534);
  and g61655 (n37154, pi0618, n37152);
  and g61656 (n37155, n_11984, n_27341);
  not g61657 (n_27535, n37155);
  and g61658 (n37156, pi1154, n_27535);
  not g61659 (n_27536, n37154);
  and g61660 (n37157, n_27536, n37156);
  and g61661 (n37158, n_11984, n37152);
  and g61662 (n37159, pi0618, n_27341);
  not g61663 (n_27537, n37159);
  and g61664 (n37160, n_11413, n_27537);
  not g61665 (n_27538, n37158);
  and g61666 (n37161, n_27538, n37160);
  not g61667 (n_27539, n37157);
  not g61668 (n_27540, n37161);
  and g61669 (n37162, n_27539, n_27540);
  not g61670 (n_27541, n37162);
  and g61671 (n37163, pi0781, n_27541);
  not g61672 (n_27542, n37153);
  not g61673 (n_27543, n37163);
  and g61674 (n37164, n_27542, n_27543);
  not g61675 (n_27544, n37164);
  and g61676 (n37165, n_12315, n_27544);
  and g61677 (n37166, pi0619, n37164);
  and g61678 (n37167, n_11821, n_27341);
  not g61679 (n_27545, n37167);
  and g61680 (n37168, pi1159, n_27545);
  not g61681 (n_27546, n37166);
  and g61682 (n37169, n_27546, n37168);
  and g61683 (n37170, n_11821, n37164);
  and g61684 (n37171, pi0619, n_27341);
  not g61685 (n_27547, n37171);
  and g61686 (n37172, n_11405, n_27547);
  not g61687 (n_27548, n37170);
  and g61688 (n37173, n_27548, n37172);
  not g61689 (n_27549, n37169);
  not g61690 (n_27550, n37173);
  and g61691 (n37174, n_27549, n_27550);
  not g61692 (n_27551, n37174);
  and g61693 (n37175, pi0789, n_27551);
  not g61694 (n_27552, n37165);
  not g61695 (n_27553, n37175);
  and g61696 (n37176, n_27552, n_27553);
  and g61697 (n37177, n_12524, n37176);
  not g61698 (n_27554, n36999);
  not g61699 (n_27555, n37177);
  and g61700 (n37178, n_27554, n_27555);
  and g61701 (n37179, n_12368, n37178);
  and g61702 (n37180, n17779, n36883);
  not g61703 (n_27556, n37179);
  not g61704 (n_27557, n37180);
  and g61705 (n37181, n_27556, n_27557);
  not g61706 (n_27558, n37181);
  and g61707 (n37182, n_14548, n_27558);
  and g61708 (n37183, pi0630, n36989);
  not g61709 (n_27559, n36998);
  not g61710 (n_27560, n37183);
  and g61711 (n37184, n_27559, n_27560);
  not g61712 (n_27561, n37182);
  and g61713 (n37185, n_27561, n37184);
  not g61714 (n_27562, n37185);
  and g61715 (n37186, pi0787, n_27562);
  and g61716 (n37187, pi0628, n_27341);
  and g61717 (n37188, n_11789, n_27412);
  not g61718 (n_27563, n37187);
  and g61719 (n37189, n17777, n_27563);
  not g61720 (n_27564, n37188);
  and g61721 (n37190, n_27564, n37189);
  and g61722 (n37191, n_14557, n37178);
  and g61723 (n37192, n_11789, n_27341);
  and g61724 (n37193, pi0628, n_27412);
  not g61725 (n_27565, n37192);
  and g61726 (n37194, n17776, n_27565);
  not g61727 (n_27566, n37193);
  and g61728 (n37195, n_27566, n37194);
  not g61729 (n_27567, n37190);
  not g61730 (n_27568, n37195);
  and g61731 (n37196, n_27567, n_27568);
  not g61732 (n_27569, n37191);
  and g61733 (n37197, n_27569, n37196);
  not g61734 (n_27570, n37197);
  and g61735 (n37198, pi0792, n_27570);
  and g61736 (n37199, n16635, n_27341);
  not g61737 (n_27571, n36979);
  not g61738 (n_27572, n37199);
  and g61739 (n37200, n_27571, n_27572);
  not g61740 (n_27573, n37200);
  and g61741 (n37201, n17871, n_27573);
  and g61742 (n37202, n_12320, n36883);
  not g61743 (n_27574, n37176);
  and g61744 (n37203, pi0626, n_27574);
  not g61745 (n_27575, n37202);
  and g61746 (n37204, n16628, n_27575);
  not g61747 (n_27576, n37203);
  and g61748 (n37205, n_27576, n37204);
  and g61749 (n37206, pi0626, n36883);
  and g61750 (n37207, n_12320, n_27574);
  not g61751 (n_27577, n37206);
  and g61752 (n37208, n16629, n_27577);
  not g61753 (n_27578, n37207);
  and g61754 (n37209, n_27578, n37208);
  not g61755 (n_27579, n37201);
  not g61756 (n_27580, n37205);
  and g61757 (n37210, n_27579, n_27580);
  not g61758 (n_27581, n37209);
  and g61759 (n37211, n_27581, n37210);
  not g61760 (n_27582, n37211);
  and g61761 (n37212, pi0788, n_27582);
  and g61762 (n37213, pi0609, n36973);
  and g61763 (n37214, n_27342, n37003);
  and g61764 (n37215, n_3087, n_12007);
  not g61765 (n_27583, n37215);
  and g61766 (n37216, n36887, n_27583);
  not g61767 (n_27584, n36562);
  and g61768 (n37217, n_27584, n37216);
  not g61769 (n_27585, n37214);
  not g61770 (n_27586, n37217);
  and g61771 (n37218, n_27585, n_27586);
  and g61772 (n37219, n_27342, n37004);
  and g61773 (n37220, pi0642, n17493);
  not g61774 (n_27587, n37220);
  and g61775 (n37221, n_27583, n_27587);
  not g61776 (n_27588, n37221);
  and g61777 (n37222, n16667, n_27588);
  and g61778 (n37223, n36887, n37222);
  not g61779 (n_27589, n37219);
  and g61780 (n37224, pi0223, n_27589);
  not g61781 (n_27590, n37223);
  and g61782 (n37225, n_27590, n37224);
  not g61783 (n_27591, n37225);
  and g61784 (n37226, n37218, n_27591);
  not g61785 (n_27592, n37226);
  and g61786 (n37227, n37006, n_27592);
  not g61787 (n_27593, n37227);
  and g61788 (n37228, n37002, n_27593);
  and g61789 (n37229, n17618, n36922);
  and g61790 (n37230, n17617, n_27342);
  and g61791 (n37231, n_27219, n37013);
  not g61792 (n_27594, n37230);
  and g61793 (n37232, n_27594, n37231);
  not g61794 (n_27595, n37229);
  and g61795 (n37233, n37011, n_27595);
  not g61796 (n_27596, n37232);
  and g61797 (n37234, n_27596, n37233);
  and g61798 (n37235, n17623, n36922);
  and g61799 (n37236, n17622, n_27342);
  not g61804 (n_27598, n37235);
  and g61805 (n37240, n37017, n_27598);
  not g61806 (n_27599, n37239);
  and g61807 (n37241, n_27599, n37240);
  not g61808 (n_27600, n37234);
  and g61809 (n37242, n_162, n_27600);
  not g61810 (n_27601, n37241);
  and g61811 (n37243, n_27601, n37242);
  and g61812 (n37244, n_27342, n_27444);
  and g61813 (n37245, n_11425, n37222);
  not g61814 (n_27602, n37245);
  and g61815 (n37246, n_24809, n_27602);
  not g61816 (n_27603, n37246);
  and g61817 (n37247, pi0680, n_27603);
  and g61818 (n37248, pi0642, n_27110);
  and g61819 (n37249, n_3090, n17343);
  not g61820 (n_27604, n37248);
  not g61821 (n_27605, n37249);
  and g61822 (n37250, n_27604, n_27605);
  not g61823 (n_27606, n37250);
  and g61824 (n37251, n_3091, n_27606);
  not g61825 (n_27607, n37251);
  and g61826 (n37252, n37247, n_27607);
  not g61827 (n_27608, n37244);
  not g61828 (n_27609, n37252);
  and g61829 (n37253, n_27608, n_27609);
  not g61830 (n_27610, n37253);
  and g61831 (n37254, n_27445, n_27610);
  not g61832 (n_27611, n37254);
  and g61833 (n37255, n6242, n_27611);
  and g61834 (n37256, n_11502, n37038);
  and g61835 (n37257, pi0642, n_27117);
  and g61836 (n37258, n_24809, n17325);
  not g61842 (n_27614, n37261);
  and g61843 (n37262, pi0681, n_27614);
  not g61844 (n_27615, n37256);
  and g61845 (n37263, n_27615, n37262);
  not g61846 (n_27616, n37263);
  and g61847 (n37264, n_27453, n_27616);
  not g61848 (n_27617, n37264);
  and g61849 (n37265, n_3162, n_27617);
  not g61850 (n_27618, n37265);
  and g61851 (n37266, pi0223, n_27618);
  not g61852 (n_27619, n37255);
  and g61853 (n37267, n_27619, n37266);
  and g61854 (n37268, n_11502, n_27457);
  and g61855 (n37269, n_12007, n_27604);
  not g61856 (n_27620, n37269);
  and g61857 (n37270, n35897, n_27620);
  not g61858 (n_27621, n37270);
  and g61859 (n37271, pi0680, n_27621);
  and g61860 (n37272, pi0642, n_27142);
  not g61861 (n_27622, n37272);
  and g61862 (n37273, n6191, n_27622);
  and g61863 (n37274, n_12105, n37273);
  not g61864 (n_27623, n37274);
  and g61865 (n37275, n37271, n_27623);
  not g61866 (n_27624, n37268);
  not g61867 (n_27625, n37275);
  and g61868 (n37276, n_27624, n_27625);
  not g61869 (n_27626, n37276);
  and g61870 (n37277, pi0681, n_27626);
  not g61871 (n_27627, n37277);
  and g61872 (n37278, n37082, n_27627);
  and g61873 (n37279, n_27342, n_27477);
  and g61874 (n37280, n_3087, n_24809);
  and g61875 (n37281, n_12103, n37280);
  and g61876 (n37282, n17454, n17559);
  not g61877 (n_27628, n37282);
  and g61878 (n37283, n17167, n_27628);
  and g61879 (n37284, pi0642, n36607);
  not g61886 (n_27632, n37279);
  not g61887 (n_27633, n37287);
  and g61888 (n37288, n_27632, n_27633);
  and g61889 (n37289, n_3162, n37077);
  not g61890 (n_27634, n37288);
  and g61891 (n37290, n_27634, n37289);
  not g61892 (n_27635, n37278);
  and g61893 (n37291, n_223, n_27635);
  not g61894 (n_27636, n37290);
  and g61895 (n37292, n_27636, n37291);
  not g61896 (n_27637, n37292);
  and g61897 (n37293, pi0215, n_27637);
  not g61898 (n_27638, n37267);
  and g61899 (n37294, n_27638, n37293);
  and g61900 (n37295, n_27342, n_27506);
  and g61901 (n37296, n_12026, n_27604);
  not g61902 (n_27639, n37296);
  and g61903 (n37297, n6191, n_27639);
  not g61904 (n_27640, n37297);
  and g61905 (n37298, n37247, n_27640);
  not g61906 (n_27641, n37295);
  not g61907 (n_27642, n37298);
  and g61908 (n37299, n_27641, n_27642);
  not g61909 (n_27643, n37299);
  and g61910 (n37300, n37122, n_27643);
  and g61911 (n37301, n_27342, n_27499);
  and g61912 (n37302, pi0642, n_27153);
  not g61913 (n_27644, n36631);
  and g61914 (n37303, n17167, n_27644);
  and g61915 (n37304, n36633, n37280);
  not g61922 (n_27648, n37301);
  not g61923 (n_27649, n37307);
  and g61924 (n37308, n_27648, n_27649);
  not g61925 (n_27650, n37308);
  and g61926 (n37309, n37111, n_27650);
  not g61927 (n_27651, n37309);
  and g61928 (n37310, pi0223, n_27651);
  not g61929 (n_27652, n37300);
  and g61930 (n37311, n_27652, n37310);
  and g61931 (n37312, n_3087, n_12193);
  not g61932 (n_27653, n37312);
  and g61933 (n37313, n37273, n_27653);
  not g61934 (n_27654, n37313);
  and g61935 (n37314, n37271, n_27654);
  not g61936 (n_27655, n37314);
  and g61937 (n37315, n_27624, n_27655);
  not g61938 (n_27656, n37315);
  and g61939 (n37316, pi0681, n_27656);
  not g61940 (n_27657, n37316);
  and g61941 (n37317, n_27460, n_27657);
  not g61942 (n_27658, n37317);
  and g61943 (n37318, n6242, n_27658);
  and g61944 (n37319, n_27342, n_27465);
  and g61945 (n37320, pi0642, n17578);
  and g61946 (n37321, n_12076, n37280);
  not g61952 (n_27661, n37319);
  not g61953 (n_27662, n37324);
  and g61954 (n37325, n_27661, n_27662);
  not g61955 (n_27663, n37325);
  and g61956 (n37326, n_27466, n_27663);
  not g61957 (n_27664, n37326);
  and g61958 (n37327, n_3162, n_27664);
  not g61959 (n_27665, n37318);
  and g61960 (n37328, n_223, n_27665);
  not g61961 (n_27666, n37327);
  and g61962 (n37329, n_27666, n37328);
  not g61963 (n_27667, n37311);
  and g61964 (n37330, n_9350, n_27667);
  not g61965 (n_27668, n37329);
  and g61966 (n37331, n_27668, n37330);
  not g61967 (n_27669, n37218);
  and g61968 (n37332, n16653, n_27669);
  and g61969 (n37333, n_223, n37332);
  and g61970 (n37334, n36931, n_27591);
  not g61971 (n_27670, n37333);
  and g61972 (n37335, n_27670, n37334);
  not g61973 (n_27671, n37335);
  and g61974 (n37336, n_36, n_27671);
  not g61975 (n_27672, n37331);
  and g61976 (n37337, n_27672, n37336);
  not g61977 (n_27673, n37294);
  and g61978 (n37338, pi0299, n_27673);
  not g61979 (n_27674, n37337);
  and g61980 (n37339, n_27674, n37338);
  and g61981 (n37340, n6205, n37254);
  and g61982 (n37341, n_3119, n37264);
  not g61983 (n_27675, n37341);
  and g61984 (n37342, pi0223, n_27675);
  not g61985 (n_27676, n37340);
  and g61986 (n37343, n_27676, n37342);
  not g61987 (n_27677, n37332);
  and g61988 (n37344, n2603, n_27677);
  and g61989 (n37345, n_3119, n37326);
  and g61990 (n37346, n6205, n37317);
  not g61991 (n_27678, n37345);
  and g61992 (n37347, n_9349, n_27678);
  not g61993 (n_27679, n37346);
  and g61994 (n37348, n_27679, n37347);
  not g61995 (n_27680, n37344);
  and g61996 (n37349, n_223, n_27680);
  not g61997 (n_27681, n37348);
  and g61998 (n37350, n_27681, n37349);
  not g61999 (n_27682, n37343);
  and g62000 (n37351, n_234, n_27682);
  not g62001 (n_27683, n37350);
  and g62002 (n37352, n_27683, n37351);
  not g62003 (n_27684, n37352);
  and g62004 (n37353, pi0039, n_27684);
  not g62005 (n_27685, n37339);
  and g62006 (n37354, n_27685, n37353);
  not g62007 (n_27686, n37243);
  and g62008 (n37355, n_161, n_27686);
  not g62009 (n_27687, n37354);
  and g62010 (n37356, n_27687, n37355);
  not g62011 (n_27688, n37228);
  and g62012 (n37357, n2571, n_27688);
  not g62013 (n_27689, n37356);
  and g62014 (n37358, n_27689, n37357);
  not g62015 (n_27690, n37358);
  and g62016 (n37359, n_27394, n_27690);
  and g62017 (n37360, n_11753, n37359);
  and g62018 (n37361, pi0625, n37138);
  not g62019 (n_27691, n37361);
  and g62020 (n37362, n_11757, n_27691);
  not g62021 (n_27692, n37360);
  and g62022 (n37363, n_27692, n37362);
  not g62023 (n_27693, n37363);
  and g62024 (n37364, n_11823, n_27693);
  and g62025 (n37365, n_27401, n37364);
  and g62026 (n37366, n_11753, n37138);
  and g62027 (n37367, pi0625, n37359);
  not g62028 (n_27694, n37366);
  and g62029 (n37368, pi1153, n_27694);
  not g62030 (n_27695, n37367);
  and g62031 (n37369, n_27695, n37368);
  not g62032 (n_27696, n37369);
  and g62033 (n37370, pi0608, n_27696);
  and g62034 (n37371, n_27402, n37370);
  not g62035 (n_27697, n37365);
  not g62036 (n_27698, n37371);
  and g62037 (n37372, n_27697, n_27698);
  not g62038 (n_27699, n37372);
  and g62039 (n37373, pi0778, n_27699);
  and g62040 (n37374, n_11749, n37359);
  not g62041 (n_27700, n37373);
  not g62042 (n_27701, n37374);
  and g62043 (n37375, n_27700, n_27701);
  not g62044 (n_27702, n37375);
  and g62045 (n37376, n_11971, n_27702);
  not g62046 (n_27703, n37213);
  and g62047 (n37377, n_11768, n_27703);
  not g62048 (n_27704, n37376);
  and g62049 (n37378, n_27704, n37377);
  and g62050 (n37379, n_11767, n_27529);
  not g62051 (n_27705, n37378);
  and g62052 (n37380, n_27705, n37379);
  and g62053 (n37381, n_11971, n36973);
  and g62054 (n37382, pi0609, n_27702);
  not g62055 (n_27706, n37381);
  and g62056 (n37383, pi1155, n_27706);
  not g62057 (n_27707, n37382);
  and g62058 (n37384, n_27707, n37383);
  and g62059 (n37385, pi0660, n_27530);
  not g62060 (n_27708, n37384);
  and g62061 (n37386, n_27708, n37385);
  not g62062 (n_27709, n37380);
  not g62063 (n_27710, n37386);
  and g62064 (n37387, n_27709, n_27710);
  not g62065 (n_27711, n37387);
  and g62066 (n37388, pi0785, n_27711);
  and g62067 (n37389, n_11964, n_27702);
  not g62068 (n_27712, n37388);
  not g62069 (n_27713, n37389);
  and g62070 (n37390, n_27712, n_27713);
  not g62071 (n_27714, n37390);
  and g62072 (n37391, n_11984, n_27714);
  not g62073 (n_27715, n36975);
  and g62074 (n37392, pi0618, n_27715);
  not g62075 (n_27716, n37392);
  and g62076 (n37393, n_11413, n_27716);
  not g62077 (n_27717, n37391);
  and g62078 (n37394, n_27717, n37393);
  and g62079 (n37395, n_11412, n_27539);
  not g62080 (n_27718, n37394);
  and g62081 (n37396, n_27718, n37395);
  and g62082 (n37397, pi0618, n_27714);
  and g62083 (n37398, n_11984, n_27715);
  not g62084 (n_27719, n37398);
  and g62085 (n37399, pi1154, n_27719);
  not g62086 (n_27720, n37397);
  and g62087 (n37400, n_27720, n37399);
  and g62088 (n37401, pi0627, n_27540);
  not g62089 (n_27721, n37400);
  and g62090 (n37402, n_27721, n37401);
  not g62091 (n_27722, n37396);
  not g62092 (n_27723, n37402);
  and g62093 (n37403, n_27722, n_27723);
  not g62094 (n_27724, n37403);
  and g62095 (n37404, pi0781, n_27724);
  and g62096 (n37405, n_11981, n_27714);
  not g62097 (n_27725, n37404);
  not g62098 (n_27726, n37405);
  and g62099 (n37406, n_27725, n_27726);
  and g62100 (n37407, n_12315, n37406);
  not g62101 (n_27727, n37406);
  and g62102 (n37408, n_11821, n_27727);
  and g62103 (n37409, pi0619, n36978);
  not g62104 (n_27728, n37409);
  and g62105 (n37410, n_11405, n_27728);
  not g62106 (n_27729, n37408);
  and g62107 (n37411, n_27729, n37410);
  and g62108 (n37412, n_11403, n_27549);
  not g62109 (n_27730, n37411);
  and g62110 (n37413, n_27730, n37412);
  and g62111 (n37414, n_11821, n36978);
  and g62112 (n37415, pi0619, n_27727);
  not g62113 (n_27731, n37414);
  and g62114 (n37416, pi1159, n_27731);
  not g62115 (n_27732, n37415);
  and g62116 (n37417, n_27732, n37416);
  and g62117 (n37418, pi0648, n_27550);
  not g62118 (n_27733, n37417);
  and g62119 (n37419, n_27733, n37418);
  not g62120 (n_27734, n37413);
  and g62121 (n37420, pi0789, n_27734);
  not g62122 (n_27735, n37419);
  and g62123 (n37421, n_27735, n37420);
  not g62124 (n_27736, n37407);
  and g62125 (n37422, n17970, n_27736);
  not g62126 (n_27737, n37421);
  and g62127 (n37423, n_27737, n37422);
  not g62128 (n_27738, n37212);
  not g62129 (n_27739, n37423);
  and g62130 (n37424, n_27738, n_27739);
  not g62131 (n_27740, n37198);
  not g62132 (n_27741, n37424);
  and g62133 (n37425, n_27740, n_27741);
  and g62134 (n37426, n20364, n37197);
  not g62135 (n_27742, n37426);
  and g62136 (n37427, n_14387, n_27742);
  not g62137 (n_27743, n37425);
  and g62138 (n37428, n_27743, n37427);
  not g62139 (n_27744, n37186);
  not g62140 (n_27745, n37428);
  and g62141 (n37429, n_27744, n_27745);
  and g62142 (n37430, pi0644, n37429);
  not g62143 (n_27746, n36997);
  and g62144 (n37431, pi0715, n_27746);
  not g62145 (n_27747, n37430);
  and g62146 (n37432, n_27747, n37431);
  and g62147 (n37433, n17804, n_27341);
  and g62148 (n37434, n_12392, n37181);
  not g62149 (n_27748, n37433);
  not g62150 (n_27749, n37434);
  and g62151 (n37435, n_27748, n_27749);
  not g62152 (n_27750, n37435);
  and g62153 (n37436, pi0644, n_27750);
  and g62154 (n37437, n_11819, n_27341);
  not g62155 (n_27751, n37437);
  and g62156 (n37438, n_12395, n_27751);
  not g62157 (n_27752, n37436);
  and g62158 (n37439, n_27752, n37438);
  not g62159 (n_27753, n37439);
  and g62160 (n37440, pi1160, n_27753);
  not g62161 (n_27754, n37432);
  and g62162 (n37441, n_27754, n37440);
  and g62163 (n37442, pi0644, n36996);
  and g62164 (n37443, n_11819, n37429);
  not g62165 (n_27755, n37442);
  and g62166 (n37444, n_12395, n_27755);
  not g62167 (n_27756, n37443);
  and g62168 (n37445, n_27756, n37444);
  and g62169 (n37446, n_11819, n_27750);
  and g62170 (n37447, pi0644, n_27341);
  not g62171 (n_27757, n37447);
  and g62172 (n37448, pi0715, n_27757);
  not g62173 (n_27758, n37446);
  and g62174 (n37449, n_27758, n37448);
  not g62175 (n_27759, n37449);
  and g62176 (n37450, n_12405, n_27759);
  not g62177 (n_27760, n37445);
  and g62178 (n37451, n_27760, n37450);
  not g62179 (n_27761, n37441);
  not g62180 (n_27762, n37451);
  and g62181 (n37452, n_27761, n_27762);
  not g62182 (n_27763, n37452);
  and g62183 (n37453, pi0790, n_27763);
  and g62184 (n37454, n_12411, n37429);
  not g62185 (n_27764, n37453);
  not g62186 (n_27765, n37454);
  and g62187 (n37455, n_27764, n_27765);
  not g62188 (n_27766, n37455);
  and g62189 (n37456, n_4226, n_27766);
  and g62190 (n37457, n_223, po1038);
  not g62191 (n_27767, n37456);
  not g62192 (n_27768, n37457);
  and g62193 (po0380, n_27767, n_27768);
  and g62194 (n37459, pi0224, n_26869);
  not g62195 (n_27769, n37459);
  and g62196 (n37460, n_24651, n_27769);
  and g62197 (n37461, pi0224, n_11417);
  and g62198 (n37462, pi0224, n_11418);
  not g62199 (n_27770, n37462);
  and g62200 (n37463, pi0038, n_27770);
  and g62201 (n37464, pi0662, n16646);
  not g62202 (n_27771, n37464);
  and g62203 (n37465, n37463, n_27771);
  and g62204 (n37466, pi0662, pi0680);
  not g62205 (n_27772, n37466);
  and g62206 (n37467, n16918, n_27772);
  and g62207 (n37468, n_219, n_12231);
  and g62208 (n37469, pi0224, n16935);
  and g62215 (n37473, pi0224, n16944);
  and g62216 (n37474, n16923, n_27772);
  and g62217 (n37475, n_219, n_12235);
  not g62224 (n_27779, n37472);
  and g62225 (n37479, n_162, n_27779);
  not g62226 (n_27780, n37478);
  and g62227 (n37480, n_27780, n37479);
  and g62228 (n37481, pi0662, n16655);
  and g62229 (n37482, n_11675, n_26883);
  not g62230 (n_27781, n37482);
  and g62231 (n37483, n17018, n_27781);
  and g62232 (n37484, n_3119, n37483);
  and g62233 (n37485, pi0662, n_26889);
  and g62234 (n37486, n_3093, n_11706);
  not g62235 (n_27782, n37485);
  not g62236 (n_27783, n37486);
  and g62237 (n37487, n_27782, n_27783);
  and g62238 (n37488, n6205, n37487);
  not g62239 (n_27784, n37484);
  and g62240 (n37489, pi0224, n_27784);
  not g62241 (n_27785, n37488);
  and g62242 (n37490, n_27785, n37489);
  and g62243 (n37491, pi0662, n16703);
  not g62244 (n_27786, n37491);
  and g62245 (n37492, n_3119, n_27786);
  and g62246 (n37493, n_26895, n37466);
  not g62247 (n_27787, n37493);
  and g62248 (n37494, n6205, n_27787);
  not g62249 (n_27788, n37492);
  and g62250 (n37495, n5810, n_27788);
  not g62251 (n_27789, n37494);
  and g62252 (n37496, n_27789, n37495);
  and g62259 (n37500, n_219, pi0662);
  and g62260 (n37501, n16729, n37500);
  and g62261 (n37502, n_3093, n_11694);
  and g62262 (n37503, pi0662, n_26907);
  not g62263 (n_27793, n37502);
  not g62264 (n_27794, n37503);
  and g62265 (n37504, n_27793, n_27794);
  and g62266 (n37505, n6205, n37504);
  and g62267 (n37506, n_3093, n_11684);
  and g62268 (n37507, pi0662, n_26903);
  not g62269 (n_27795, n37506);
  not g62270 (n_27796, n37507);
  and g62271 (n37508, n_27795, n_27796);
  and g62272 (n37509, n_3119, n37508);
  not g62273 (n_27797, n37505);
  and g62274 (n37510, pi0224, n_27797);
  not g62275 (n_27798, n37509);
  and g62276 (n37511, n_27798, n37510);
  not g62277 (n_27799, n37501);
  and g62278 (n37512, pi0223, n_27799);
  not g62279 (n_27800, n37511);
  and g62280 (n37513, n_27800, n37512);
  not g62281 (n_27801, n37513);
  and g62282 (n37514, n_234, n_27801);
  not g62283 (n_27802, n37499);
  and g62284 (n37515, n_27802, n37514);
  and g62285 (n37516, pi0224, n_11445);
  not g62286 (n_27803, n37516);
  and g62287 (n37517, n3448, n_27803);
  and g62288 (n37518, n16658, n37466);
  not g62289 (n_27804, n37518);
  and g62290 (n37519, n37517, n_27804);
  and g62291 (n37520, n_3162, n37483);
  and g62292 (n37521, n6242, n37487);
  not g62293 (n_27805, n37520);
  and g62294 (n37522, pi0224, n_27805);
  not g62295 (n_27806, n37521);
  and g62296 (n37523, n_27806, n37522);
  and g62297 (n37524, n_3162, n_27786);
  and g62298 (n37525, n6242, n_27787);
  not g62299 (n_27807, n37524);
  and g62300 (n37526, n_219, n_27807);
  not g62301 (n_27808, n37525);
  and g62302 (n37527, n_27808, n37526);
  not g62303 (n_27809, n37527);
  and g62304 (n37528, n_9350, n_27809);
  not g62305 (n_27810, n37523);
  and g62306 (n37529, n_27810, n37528);
  not g62307 (n_27811, n37519);
  not g62308 (n_27812, n37529);
  and g62309 (n37530, n_27811, n_27812);
  not g62310 (n_27813, n37530);
  and g62311 (n37531, n_36, n_27813);
  and g62312 (n37532, n16744, n37500);
  and g62313 (n37533, n6242, n37504);
  and g62314 (n37534, n_3162, n37508);
  not g62315 (n_27814, n37533);
  and g62316 (n37535, pi0224, n_27814);
  not g62317 (n_27815, n37534);
  and g62318 (n37536, n_27815, n37535);
  not g62319 (n_27816, n37532);
  and g62320 (n37537, pi0215, n_27816);
  not g62321 (n_27817, n37536);
  and g62322 (n37538, n_27817, n37537);
  not g62323 (n_27818, n37538);
  and g62324 (n37539, pi0299, n_27818);
  not g62325 (n_27819, n37531);
  and g62326 (n37540, n_27819, n37539);
  not g62327 (n_27820, n37515);
  and g62328 (n37541, pi0039, n_27820);
  not g62329 (n_27821, n37540);
  and g62330 (n37542, n_27821, n37541);
  not g62331 (n_27822, n37480);
  not g62332 (n_27823, n37542);
  and g62333 (n37543, n_27822, n_27823);
  not g62334 (n_27824, n37543);
  and g62335 (n37544, n_161, n_27824);
  not g62336 (n_27825, n37465);
  and g62337 (n37545, n2571, n_27825);
  not g62338 (n_27826, n37544);
  and g62339 (n37546, n_27826, n37545);
  not g62340 (n_27827, n37461);
  not g62341 (n_27828, n37546);
  and g62342 (n37547, n_27827, n_27828);
  not g62343 (n_27829, n37547);
  and g62344 (n37548, n_11749, n_27829);
  and g62345 (n37549, pi0625, n37547);
  and g62346 (n37550, n_11753, n_27769);
  not g62347 (n_27830, n37550);
  and g62348 (n37551, pi1153, n_27830);
  not g62349 (n_27831, n37549);
  and g62350 (n37552, n_27831, n37551);
  and g62351 (n37553, n_11753, n37547);
  and g62352 (n37554, pi0625, n_27769);
  not g62353 (n_27832, n37554);
  and g62354 (n37555, n_11757, n_27832);
  not g62355 (n_27833, n37553);
  and g62356 (n37556, n_27833, n37555);
  not g62357 (n_27834, n37552);
  not g62358 (n_27835, n37556);
  and g62359 (n37557, n_27834, n_27835);
  not g62360 (n_27836, n37557);
  and g62361 (n37558, pi0778, n_27836);
  not g62362 (n_27837, n37548);
  not g62363 (n_27838, n37558);
  and g62364 (n37559, n_27837, n_27838);
  not g62365 (n_27839, n37559);
  and g62366 (n37560, n_11773, n_27839);
  and g62367 (n37561, n17075, n37459);
  not g62368 (n_27840, n37560);
  not g62369 (n_27841, n37561);
  and g62370 (n37562, n_27840, n_27841);
  not g62371 (n_27842, n37562);
  and g62372 (n37563, n_11777, n_27842);
  and g62373 (n37564, n16639, n37459);
  not g62374 (n_27843, n37563);
  not g62375 (n_27844, n37564);
  and g62376 (n37565, n_27843, n_27844);
  and g62377 (n37566, n_11780, n37565);
  and g62378 (n37567, n_11783, n37566);
  not g62379 (n_27845, n37460);
  not g62380 (n_27846, n37567);
  and g62381 (n37568, n_27845, n_27846);
  not g62382 (n_27847, n37568);
  and g62383 (n37569, n_13453, n_27847);
  and g62384 (n37570, n17856, n_27769);
  not g62385 (n_27848, n37569);
  not g62386 (n_27849, n37570);
  and g62387 (n37571, n_27848, n_27849);
  and g62388 (n37572, n_11803, n37571);
  not g62389 (n_27850, n37571);
  and g62390 (n37573, n_11806, n_27850);
  and g62391 (n37574, pi0647, n_27769);
  not g62392 (n_27851, n37574);
  and g62393 (n37575, n_11810, n_27851);
  not g62394 (n_27852, n37573);
  and g62395 (n37576, n_27852, n37575);
  and g62396 (n37577, pi0647, n_27850);
  and g62397 (n37578, n_11806, n_27769);
  not g62398 (n_27853, n37578);
  and g62399 (n37579, pi1157, n_27853);
  not g62400 (n_27854, n37577);
  and g62401 (n37580, n_27854, n37579);
  not g62402 (n_27855, n37576);
  not g62403 (n_27856, n37580);
  and g62404 (n37581, n_27855, n_27856);
  not g62405 (n_27857, n37581);
  and g62406 (n37582, pi0787, n_27857);
  not g62407 (n_27858, n37572);
  not g62408 (n_27859, n37582);
  and g62409 (n37583, n_27858, n_27859);
  and g62410 (n37584, n_11819, n37583);
  and g62411 (n37585, pi0628, n_27769);
  and g62412 (n37586, n_11789, n_27847);
  not g62413 (n_27860, n37585);
  and g62414 (n37587, n17777, n_27860);
  not g62415 (n_27861, n37586);
  and g62416 (n37588, n_27861, n37587);
  and g62417 (n37589, n17969, n_27769);
  and g62418 (n37590, pi0614, n17280);
  not g62419 (n_27862, n37590);
  and g62420 (n37591, n37463, n_27862);
  and g62421 (n37592, pi0614, n17226);
  and g62422 (n37593, n_219, n37592);
  and g62423 (n37594, n_3090, n17226);
  not g62424 (n_27863, n37594);
  and g62425 (n37595, pi0224, n_27863);
  and g62426 (n37596, n17137, n37595);
  not g62427 (n_27864, n37593);
  and g62428 (n37597, n_234, n_27864);
  not g62429 (n_27865, n37596);
  and g62430 (n37598, n_27865, n37597);
  and g62431 (n37599, pi0614, n17231);
  and g62432 (n37600, pi0224, n17122);
  not g62433 (n_27866, n37600);
  and g62434 (n37601, n37599, n_27866);
  and g62435 (n37602, pi0224, n_11670);
  not g62436 (n_27867, n37601);
  not g62437 (n_27868, n37602);
  and g62438 (n37603, n_27867, n_27868);
  and g62439 (n37604, pi0299, n37603);
  not g62440 (n_27869, n37598);
  and g62441 (n37605, n_162, n_27869);
  not g62442 (n_27870, n37604);
  and g62443 (n37606, n_27870, n37605);
  and g62444 (n37607, pi0614, n_26983);
  and g62445 (n37608, n_219, n37607);
  and g62446 (n37609, n_11494, n37608);
  and g62447 (n37610, pi0614, n_27446);
  not g62448 (n_27871, n37610);
  and g62449 (n37611, n_26686, n_27871);
  not g62450 (n_27872, n37611);
  and g62451 (n37612, n_11502, n_27872);
  and g62452 (n37613, pi0680, n_11880);
  not g62453 (n_27873, n36028);
  and g62454 (n37614, n_27873, n37613);
  not g62455 (n_27874, n37612);
  not g62456 (n_27875, n37614);
  and g62457 (n37615, n_27874, n_27875);
  not g62458 (n_27876, n37615);
  and g62459 (n37616, n16657, n_27876);
  and g62460 (n37617, n_11455, n_27872);
  not g62461 (n_27877, n37616);
  not g62462 (n_27878, n37617);
  and g62463 (n37618, n_27877, n_27878);
  and g62464 (n37619, n_3162, n37618);
  and g62465 (n37620, pi0614, n17168);
  not g62466 (n_27879, n37620);
  and g62467 (n37621, n16653, n_27879);
  not g62468 (n_27880, n37621);
  and g62469 (n37622, n_3138, n_27880);
  not g62470 (n_27881, n37622);
  and g62471 (n37623, n_11548, n_27881);
  not g62472 (n_27882, n37623);
  and g62473 (n37624, n_11455, n_27882);
  and g62474 (n37625, n_11502, n_27882);
  and g62475 (n37626, pi0680, n37620);
  not g62476 (n_27883, n37626);
  and g62477 (n37627, n_11686, n_27883);
  not g62478 (n_27884, n37625);
  and g62479 (n37628, n_27884, n37627);
  not g62480 (n_27885, n37628);
  and g62481 (n37629, n16657, n_27885);
  not g62482 (n_27886, n37624);
  not g62483 (n_27887, n37629);
  and g62484 (n37630, n_27886, n_27887);
  and g62485 (n37631, n6242, n37630);
  not g62486 (n_27888, n37619);
  and g62487 (n37632, pi0224, n_27888);
  not g62488 (n_27889, n37631);
  and g62489 (n37633, n_27889, n37632);
  not g62490 (n_27890, n37609);
  not g62491 (n_27891, n37633);
  and g62492 (n37634, n_27890, n_27891);
  not g62493 (n_27892, n37634);
  and g62494 (n37635, pi0215, n_27892);
  and g62495 (n37636, n16999, n17168);
  not g62496 (n_27893, n37636);
  and g62497 (n37637, n37517, n_27893);
  and g62498 (n37638, pi0614, n_11856);
  and g62499 (n37639, n_3090, pi0616);
  and g62500 (n37640, n16699, n37639);
  and g62501 (n37641, n_3102, n16772);
  and g62502 (n37642, n6191, n_11460);
  not g62503 (n_27894, n37641);
  and g62504 (n37643, n_27894, n37642);
  not g62505 (n_27895, n37638);
  not g62506 (n_27896, n37640);
  and g62507 (n37644, n_27895, n_27896);
  not g62508 (n_27897, n37643);
  and g62509 (n37645, n_27897, n37644);
  not g62510 (n_27898, n37645);
  and g62511 (n37646, n_11455, n_27898);
  and g62512 (n37647, n_11502, n_27898);
  and g62513 (n37648, pi0614, n17375);
  not g62514 (n_27899, n37648);
  and g62515 (n37649, pi0680, n_27899);
  and g62516 (n37650, n16681, n37649);
  not g62517 (n_27900, n37650);
  and g62518 (n37651, n_27883, n_27900);
  not g62519 (n_27901, n37647);
  and g62520 (n37652, n_27901, n37651);
  not g62521 (n_27902, n37652);
  and g62522 (n37653, n16657, n_27902);
  not g62523 (n_27903, n37646);
  not g62524 (n_27904, n37653);
  and g62525 (n37654, n_27903, n_27904);
  and g62526 (n37655, n_3162, n37654);
  and g62527 (n37656, n_11525, n_27881);
  not g62528 (n_27905, n37656);
  and g62529 (n37657, n_11455, n_27905);
  and g62530 (n37658, n_11502, n_27905);
  and g62531 (n37659, n_11698, n_27883);
  not g62532 (n_27906, n37658);
  and g62533 (n37660, n_27906, n37659);
  not g62534 (n_27907, n37660);
  and g62535 (n37661, n16657, n_27907);
  not g62536 (n_27908, n37657);
  not g62537 (n_27909, n37661);
  and g62538 (n37662, n_27908, n_27909);
  and g62539 (n37663, n6242, n37662);
  not g62540 (n_27910, n37655);
  and g62541 (n37664, pi0224, n_27910);
  not g62542 (n_27911, n37663);
  and g62543 (n37665, n_27911, n37664);
  and g62544 (n37666, n_12078, n37620);
  not g62545 (n_27912, n37666);
  and g62546 (n37667, n_11502, n_27912);
  not g62547 (n_27913, n37649);
  not g62548 (n_27914, n37667);
  and g62549 (n37668, n_27913, n_27914);
  not g62550 (n_27915, n37668);
  and g62551 (n37669, n16657, n_27915);
  and g62552 (n37670, n_11455, n_27912);
  not g62553 (n_27916, n37669);
  not g62554 (n_27917, n37670);
  and g62555 (n37671, n_27916, n_27917);
  not g62556 (n_27918, n37671);
  and g62557 (n37672, n_3162, n_27918);
  and g62558 (n37673, pi0614, n_27022);
  not g62559 (n_27919, n37673);
  and g62560 (n37674, n6242, n_27919);
  not g62561 (n_27920, n37674);
  and g62562 (n37675, n_219, n_27920);
  not g62563 (n_27921, n37672);
  and g62564 (n37676, n_27921, n37675);
  not g62565 (n_27922, n37676);
  and g62566 (n37677, n_9350, n_27922);
  not g62567 (n_27923, n37665);
  and g62568 (n37678, n_27923, n37677);
  not g62569 (n_27924, n37637);
  and g62570 (n37679, n_36, n_27924);
  not g62571 (n_27925, n37678);
  and g62572 (n37680, n_27925, n37679);
  not g62573 (n_27926, n37635);
  and g62574 (n37681, pi0299, n_27926);
  not g62575 (n_27927, n37680);
  and g62576 (n37682, n_27927, n37681);
  and g62577 (n37683, n_11484, n37608);
  and g62578 (n37684, n_3119, n37618);
  and g62579 (n37685, n6205, n37630);
  not g62580 (n_27928, n37684);
  and g62581 (n37686, pi0224, n_27928);
  not g62582 (n_27929, n37685);
  and g62583 (n37687, n_27929, n37686);
  not g62584 (n_27930, n37683);
  and g62585 (n37688, pi0223, n_27930);
  not g62586 (n_27931, n37687);
  and g62587 (n37689, n_27931, n37688);
  and g62588 (n37690, pi0614, n17268);
  and g62589 (n37691, n6205, n_27919);
  and g62590 (n37692, n_3119, n_27918);
  not g62591 (n_27932, n37691);
  and g62592 (n37693, n5810, n_27932);
  not g62593 (n_27933, n37692);
  and g62594 (n37694, n_27933, n37693);
  and g62595 (n37695, n_3119, n37654);
  and g62596 (n37696, n6205, n37662);
  not g62597 (n_27934, n37695);
  and g62598 (n37697, pi0224, n_27934);
  not g62599 (n_27935, n37696);
  and g62600 (n37698, n_27935, n37697);
  not g62607 (n_27939, n37689);
  not g62608 (n_27940, n37701);
  and g62609 (n37702, n_27939, n_27940);
  not g62610 (n_27941, n37702);
  and g62611 (n37703, n_234, n_27941);
  not g62612 (n_27942, n37682);
  and g62613 (n37704, pi0039, n_27942);
  not g62614 (n_27943, n37703);
  and g62615 (n37705, n_27943, n37704);
  not g62616 (n_27944, n37606);
  and g62617 (n37706, n_161, n_27944);
  not g62618 (n_27945, n37705);
  and g62619 (n37707, n_27945, n37706);
  not g62620 (n_27946, n37591);
  and g62621 (n37708, n2571, n_27946);
  not g62622 (n_27947, n37707);
  and g62623 (n37709, n_27947, n37708);
  not g62624 (n_27948, n37709);
  and g62625 (n37710, n_27827, n_27948);
  not g62626 (n_27949, n37710);
  and g62627 (n37711, n_11960, n_27949);
  and g62628 (n37712, n17117, n37459);
  not g62629 (n_27950, n37711);
  not g62630 (n_27951, n37712);
  and g62631 (n37713, n_27950, n_27951);
  not g62632 (n_27952, n37713);
  and g62633 (n37714, n_11964, n_27952);
  and g62634 (n37715, pi0609, n37713);
  and g62635 (n37716, n_11971, n_27769);
  not g62636 (n_27953, n37716);
  and g62637 (n37717, pi1155, n_27953);
  not g62638 (n_27954, n37715);
  and g62639 (n37718, n_27954, n37717);
  and g62640 (n37719, n_11971, n37713);
  and g62641 (n37720, pi0609, n_27769);
  not g62642 (n_27955, n37720);
  and g62643 (n37721, n_11768, n_27955);
  not g62644 (n_27956, n37719);
  and g62645 (n37722, n_27956, n37721);
  not g62646 (n_27957, n37718);
  not g62647 (n_27958, n37722);
  and g62648 (n37723, n_27957, n_27958);
  not g62649 (n_27959, n37723);
  and g62650 (n37724, pi0785, n_27959);
  not g62651 (n_27960, n37714);
  not g62652 (n_27961, n37724);
  and g62653 (n37725, n_27960, n_27961);
  not g62654 (n_27962, n37725);
  and g62655 (n37726, n_11981, n_27962);
  and g62656 (n37727, pi0618, n37725);
  and g62657 (n37728, n_11984, n_27769);
  not g62658 (n_27963, n37728);
  and g62659 (n37729, pi1154, n_27963);
  not g62660 (n_27964, n37727);
  and g62661 (n37730, n_27964, n37729);
  and g62662 (n37731, n_11984, n37725);
  and g62663 (n37732, pi0618, n_27769);
  not g62664 (n_27965, n37732);
  and g62665 (n37733, n_11413, n_27965);
  not g62666 (n_27966, n37731);
  and g62667 (n37734, n_27966, n37733);
  not g62668 (n_27967, n37730);
  not g62669 (n_27968, n37734);
  and g62670 (n37735, n_27967, n_27968);
  not g62671 (n_27969, n37735);
  and g62672 (n37736, pi0781, n_27969);
  not g62673 (n_27970, n37726);
  not g62674 (n_27971, n37736);
  and g62675 (n37737, n_27970, n_27971);
  not g62676 (n_27972, n37737);
  and g62677 (n37738, n_12315, n_27972);
  and g62678 (n37739, pi0619, n37737);
  and g62679 (n37740, n_11821, n_27769);
  not g62680 (n_27973, n37740);
  and g62681 (n37741, pi1159, n_27973);
  not g62682 (n_27974, n37739);
  and g62683 (n37742, n_27974, n37741);
  and g62684 (n37743, n_11821, n37737);
  and g62685 (n37744, pi0619, n_27769);
  not g62686 (n_27975, n37744);
  and g62687 (n37745, n_11405, n_27975);
  not g62688 (n_27976, n37743);
  and g62689 (n37746, n_27976, n37745);
  not g62690 (n_27977, n37742);
  not g62691 (n_27978, n37746);
  and g62692 (n37747, n_27977, n_27978);
  not g62693 (n_27979, n37747);
  and g62694 (n37748, pi0789, n_27979);
  not g62695 (n_27980, n37738);
  not g62696 (n_27981, n37748);
  and g62697 (n37749, n_27980, n_27981);
  and g62698 (n37750, n_12524, n37749);
  not g62699 (n_27982, n37589);
  not g62700 (n_27983, n37750);
  and g62701 (n37751, n_27982, n_27983);
  and g62702 (n37752, n_14557, n37751);
  and g62703 (n37753, n_11789, n_27769);
  and g62704 (n37754, pi0628, n_27847);
  not g62705 (n_27984, n37753);
  and g62706 (n37755, n17776, n_27984);
  not g62707 (n_27985, n37754);
  and g62708 (n37756, n_27985, n37755);
  not g62709 (n_27986, n37588);
  not g62710 (n_27987, n37756);
  and g62711 (n37757, n_27986, n_27987);
  not g62712 (n_27988, n37752);
  and g62713 (n37758, n_27988, n37757);
  not g62714 (n_27989, n37758);
  and g62715 (n37759, pi0792, n_27989);
  and g62716 (n37760, pi0609, n37559);
  and g62717 (n37761, pi0662, n17355);
  and g62718 (n37762, n16641, n37761);
  not g62719 (n_27990, n37762);
  and g62720 (n37763, n37591, n_27990);
  and g62721 (n37764, n17617, n37466);
  not g62722 (n_27991, n37592);
  not g62723 (n_27992, n37764);
  and g62724 (n37765, n_27991, n_27992);
  not g62725 (n_27993, n37765);
  and g62726 (n37766, n_219, n_27993);
  and g62727 (n37767, n17617, n_27772);
  and g62728 (n37768, n_27219, n37595);
  not g62729 (n_27994, n37767);
  and g62730 (n37769, n_27994, n37768);
  not g62731 (n_27995, n37766);
  not g62732 (n_27996, n37769);
  and g62733 (n37770, n_27995, n_27996);
  not g62734 (n_27997, n37770);
  and g62735 (n37771, n_234, n_27997);
  and g62736 (n37772, n_27772, n37603);
  and g62737 (n37773, n_3090, n17231);
  not g62738 (n_27998, n37773);
  and g62739 (n37774, n_27227, n_27998);
  not g62740 (n_27999, n37774);
  and g62741 (n37775, pi0224, n_27999);
  not g62742 (n_28000, n17622);
  and g62743 (n37776, n_219, n_28000);
  not g62744 (n_28001, n37599);
  and g62745 (n37777, n_28001, n37776);
  not g62746 (n_28002, n37775);
  not g62747 (n_28003, n37777);
  and g62748 (n37778, n_28002, n_28003);
  not g62749 (n_28004, n37778);
  and g62750 (n37779, n37466, n_28004);
  not g62751 (n_28005, n37772);
  and g62752 (n37780, pi0299, n_28005);
  not g62753 (n_28006, n37779);
  and g62754 (n37781, n_28006, n37780);
  not g62755 (n_28007, n37771);
  not g62756 (n_28008, n37781);
  and g62757 (n37782, n_28007, n_28008);
  not g62758 (n_28009, n37782);
  and g62759 (n37783, n_162, n_28009);
  and g62760 (n37784, n17407, n37466);
  not g62761 (n_28010, n37784);
  and g62762 (n37785, n_27893, n_28010);
  not g62763 (n_28011, n37785);
  and g62764 (n37786, n_219, n_28011);
  and g62765 (n37787, n_226, n37786);
  and g62766 (n37788, n_12066, n37639);
  not g62767 (n_28012, n37788);
  and g62768 (n37789, n_27143, n_28012);
  not g62769 (n_28013, n37789);
  and g62770 (n37790, pi0680, n_28013);
  not g62771 (n_28014, n36675);
  and g62772 (n37791, n_28014, n_27893);
  not g62773 (n_28015, n37790);
  not g62774 (n_28016, n37791);
  and g62775 (n37792, n_28015, n_28016);
  not g62776 (n_28017, n37792);
  and g62777 (n37793, pi0662, n_28017);
  and g62778 (n37794, n_3093, n_27919);
  not g62779 (n_28018, n37793);
  not g62780 (n_28019, n37794);
  and g62781 (n37795, n_28018, n_28019);
  not g62782 (n_28020, n37795);
  and g62783 (n37796, n6205, n_28020);
  and g62784 (n37797, n_3093, n_26986);
  and g62785 (n37798, n_27912, n37797);
  and g62786 (n37799, n_3090, n17434);
  and g62787 (n37800, pi0614, n_12201);
  not g62788 (n_28021, n37800);
  and g62789 (n37801, pi0680, n_28021);
  not g62790 (n_28022, n37799);
  and g62791 (n37802, n_28022, n37801);
  not g62792 (n_28023, n37802);
  and g62793 (n37803, n_27914, n_28023);
  not g62794 (n_28024, n37803);
  and g62795 (n37804, pi0662, n_28024);
  not g62796 (n_28025, n37798);
  and g62797 (n37805, n_27916, n_28025);
  not g62798 (n_28026, n37804);
  and g62799 (n37806, n_28026, n37805);
  not g62800 (n_28027, n37806);
  and g62801 (n37807, n_3119, n_28027);
  not g62802 (n_28028, n37796);
  and g62803 (n37808, n5810, n_28028);
  not g62804 (n_28029, n37807);
  and g62805 (n37809, n_28029, n37808);
  and g62806 (n37810, n_27905, n37797);
  not g62807 (n_28030, n24055);
  and g62808 (n37811, n_3090, n_28030);
  and g62809 (n37812, pi0614, n_27584);
  not g62810 (n_28031, n37811);
  not g62811 (n_28032, n37812);
  and g62812 (n37813, n_28031, n_28032);
  and g62813 (n37814, n_11425, n37813);
  not g62814 (n_28033, n37814);
  and g62815 (n37815, pi0616, n_28033);
  and g62816 (n37816, pi0614, n_27110);
  not g62817 (n_28034, n37816);
  and g62818 (n37817, n_12028, n_28034);
  not g62819 (n_28035, n37817);
  and g62820 (n37818, n_3091, n_28035);
  not g62821 (n_28036, n37815);
  not g62822 (n_28037, n37818);
  and g62823 (n37819, n_28036, n_28037);
  not g62824 (n_28038, n37819);
  and g62825 (n37820, pi0680, n_28038);
  not g62826 (n_28039, n37820);
  and g62827 (n37821, n_27906, n_28039);
  not g62828 (n_28040, n37821);
  and g62829 (n37822, pi0662, n_28040);
  not g62830 (n_28041, n37810);
  and g62831 (n37823, n_27909, n_28041);
  not g62832 (n_28042, n37822);
  and g62833 (n37824, n_28042, n37823);
  and g62834 (n37825, n6205, n37824);
  and g62835 (n37826, n_27898, n37797);
  and g62836 (n37827, pi0614, n_27153);
  and g62837 (n37828, n36633, n37639);
  not g62838 (n_28043, n37827);
  not g62839 (n_28044, n37828);
  and g62840 (n37829, n_28043, n_28044);
  and g62841 (n37830, n_27156, n37829);
  not g62842 (n_28045, n37830);
  and g62843 (n37831, pi0680, n_28045);
  not g62844 (n_28046, n37831);
  and g62845 (n37832, n_27901, n_28046);
  not g62846 (n_28047, n37832);
  and g62847 (n37833, pi0662, n_28047);
  not g62848 (n_28048, n37826);
  and g62849 (n37834, n_27904, n_28048);
  not g62850 (n_28049, n37833);
  and g62851 (n37835, n_28049, n37834);
  and g62852 (n37836, n_3119, n37835);
  not g62853 (n_28050, n37836);
  and g62854 (n37837, pi0224, n_28050);
  not g62855 (n_28051, n37825);
  and g62856 (n37838, n_28051, n37837);
  and g62863 (n37842, pi0680, n_12099);
  not g62864 (n_28055, n37842);
  and g62865 (n37843, n_27893, n_28055);
  not g62866 (n_28056, n37843);
  and g62867 (n37844, n_28015, n_28056);
  not g62868 (n_28057, n37844);
  and g62869 (n37845, pi0662, n_28057);
  not g62870 (n_28058, n37607);
  and g62871 (n37846, n_3093, n_28058);
  not g62872 (n_28059, n37845);
  not g62873 (n_28060, n37846);
  and g62874 (n37847, n_28059, n_28060);
  not g62875 (n_28061, n37847);
  and g62876 (n37848, n_219, n_28061);
  and g62877 (n37849, n_27882, n37797);
  and g62878 (n37850, n_12013, n_28034);
  not g62879 (n_28062, n37850);
  and g62880 (n37851, n_3091, n_28062);
  not g62881 (n_28063, n37851);
  and g62882 (n37852, n_28036, n_28063);
  not g62883 (n_28064, n37852);
  and g62884 (n37853, pi0680, n_28064);
  not g62885 (n_28065, n37853);
  and g62886 (n37854, n_27884, n_28065);
  not g62887 (n_28066, n37854);
  and g62888 (n37855, pi0662, n_28066);
  not g62889 (n_28067, n37849);
  and g62890 (n37856, n_27887, n_28067);
  not g62891 (n_28068, n37855);
  and g62892 (n37857, n_28068, n37856);
  and g62893 (n37858, pi0224, n37857);
  not g62894 (n_28069, n37848);
  and g62895 (n37859, n6205, n_28069);
  not g62896 (n_28070, n37858);
  and g62897 (n37860, n_28070, n37859);
  and g62898 (n37861, n_27872, n37797);
  and g62899 (n37862, pi0614, n_27117);
  not g62900 (n_28071, n37862);
  and g62901 (n37863, n17330, n_28071);
  not g62902 (n_28072, n37863);
  and g62903 (n37864, pi0680, n_28072);
  not g62904 (n_28073, n37864);
  and g62905 (n37865, n_27874, n_28073);
  not g62906 (n_28074, n37865);
  and g62907 (n37866, pi0662, n_28074);
  not g62908 (n_28075, n37861);
  and g62909 (n37867, n_27877, n_28075);
  not g62910 (n_28076, n37866);
  and g62911 (n37868, n_28076, n37867);
  and g62912 (n37869, pi0224, n37868);
  and g62913 (n37870, n_11556, n37607);
  not g62914 (n_28077, n37870);
  and g62915 (n37871, n_3093, n_28077);
  and g62916 (n37872, pi0614, n_11502);
  and g62917 (n37873, n17237, n37872);
  and g62918 (n37874, pi0614, n36607);
  and g62919 (n37875, n_3090, n17451);
  not g62925 (n_28080, n37873);
  and g62926 (n37879, pi0662, n_28080);
  not g62927 (n_28081, n37878);
  and g62928 (n37880, n_28081, n37879);
  not g62929 (n_28082, n37871);
  not g62930 (n_28083, n37880);
  and g62931 (n37881, n_28082, n_28083);
  not g62932 (n_28084, n37881);
  and g62933 (n37882, n_219, n_28084);
  not g62934 (n_28085, n37882);
  and g62935 (n37883, n_3119, n_28085);
  not g62936 (n_28086, n37869);
  and g62937 (n37884, n_28086, n37883);
  not g62938 (n_28087, n37884);
  and g62939 (n37885, pi0223, n_28087);
  not g62940 (n_28088, n37860);
  and g62941 (n37886, n_28088, n37885);
  not g62942 (n_28089, n37841);
  not g62943 (n_28090, n37886);
  and g62944 (n37887, n_28089, n_28090);
  not g62945 (n_28091, n37887);
  and g62946 (n37888, n_234, n_28091);
  not g62947 (n_28092, n37868);
  and g62948 (n37889, n_3162, n_28092);
  not g62949 (n_28093, n37857);
  and g62950 (n37890, n6242, n_28093);
  not g62951 (n_28094, n37889);
  and g62952 (n37891, pi0224, n_28094);
  not g62953 (n_28095, n37890);
  and g62954 (n37892, n_28095, n37891);
  and g62955 (n37893, n6242, n37847);
  and g62956 (n37894, n_3162, n37881);
  not g62957 (n_28096, n37894);
  and g62958 (n37895, n_219, n_28096);
  not g62959 (n_28097, n37893);
  and g62960 (n37896, n_28097, n37895);
  not g62961 (n_28098, n37896);
  and g62962 (n37897, pi0215, n_28098);
  not g62963 (n_28099, n37892);
  and g62964 (n37898, n_28099, n37897);
  and g62965 (n37899, n37466, n37813);
  and g62966 (n37900, n_27772, n_27879);
  and g62967 (n37901, n16667, n37900);
  not g62968 (n_28100, n37901);
  and g62969 (n37902, pi0224, n_28100);
  not g62970 (n_28101, n37899);
  and g62971 (n37903, n_28101, n37902);
  not g62972 (n_28102, n37903);
  and g62973 (n37904, n37517, n_28102);
  not g62974 (n_28103, n37786);
  and g62975 (n37905, n_28103, n37904);
  and g62976 (n37906, n_219, n_28020);
  and g62977 (n37907, pi0224, n37824);
  not g62978 (n_28104, n37906);
  and g62979 (n37908, n6242, n_28104);
  not g62980 (n_28105, n37907);
  and g62981 (n37909, n_28105, n37908);
  and g62982 (n37910, n_219, n_28027);
  and g62983 (n37911, pi0224, n37835);
  not g62984 (n_28106, n37910);
  and g62985 (n37912, n_3162, n_28106);
  not g62986 (n_28107, n37911);
  and g62987 (n37913, n_28107, n37912);
  not g62988 (n_28108, n37909);
  and g62989 (n37914, n_9350, n_28108);
  not g62990 (n_28109, n37913);
  and g62991 (n37915, n_28109, n37914);
  not g62992 (n_28110, n37905);
  and g62993 (n37916, n_36, n_28110);
  not g62994 (n_28111, n37915);
  and g62995 (n37917, n_28111, n37916);
  not g62996 (n_28112, n37898);
  and g62997 (n37918, pi0299, n_28112);
  not g62998 (n_28113, n37917);
  and g62999 (n37919, n_28113, n37918);
  not g63000 (n_28114, n37888);
  and g63001 (n37920, pi0039, n_28114);
  not g63002 (n_28115, n37919);
  and g63003 (n37921, n_28115, n37920);
  not g63004 (n_28116, n37783);
  and g63005 (n37922, n_161, n_28116);
  not g63006 (n_28117, n37921);
  and g63007 (n37923, n_28117, n37922);
  not g63008 (n_28118, n37763);
  and g63009 (n37924, n2571, n_28118);
  not g63010 (n_28119, n37923);
  and g63011 (n37925, n_28119, n37924);
  not g63012 (n_28120, n37925);
  and g63013 (n37926, n_27827, n_28120);
  and g63014 (n37927, n_11753, n37926);
  and g63015 (n37928, pi0625, n37710);
  not g63016 (n_28121, n37928);
  and g63017 (n37929, n_11757, n_28121);
  not g63018 (n_28122, n37927);
  and g63019 (n37930, n_28122, n37929);
  and g63020 (n37931, n_11823, n_27834);
  not g63021 (n_28123, n37930);
  and g63022 (n37932, n_28123, n37931);
  and g63023 (n37933, n_11753, n37710);
  and g63024 (n37934, pi0625, n37926);
  not g63025 (n_28124, n37933);
  and g63026 (n37935, pi1153, n_28124);
  not g63027 (n_28125, n37934);
  and g63028 (n37936, n_28125, n37935);
  and g63029 (n37937, pi0608, n_27835);
  not g63030 (n_28126, n37936);
  and g63031 (n37938, n_28126, n37937);
  not g63032 (n_28127, n37932);
  not g63033 (n_28128, n37938);
  and g63034 (n37939, n_28127, n_28128);
  not g63035 (n_28129, n37939);
  and g63036 (n37940, pi0778, n_28129);
  and g63037 (n37941, n_11749, n37926);
  not g63038 (n_28130, n37940);
  not g63039 (n_28131, n37941);
  and g63040 (n37942, n_28130, n_28131);
  not g63041 (n_28132, n37942);
  and g63042 (n37943, n_11971, n_28132);
  not g63043 (n_28133, n37760);
  and g63044 (n37944, n_11768, n_28133);
  not g63045 (n_28134, n37943);
  and g63046 (n37945, n_28134, n37944);
  and g63047 (n37946, n_11767, n_27957);
  not g63048 (n_28135, n37945);
  and g63049 (n37947, n_28135, n37946);
  and g63050 (n37948, n_11971, n37559);
  and g63051 (n37949, pi0609, n_28132);
  not g63052 (n_28136, n37948);
  and g63053 (n37950, pi1155, n_28136);
  not g63054 (n_28137, n37949);
  and g63055 (n37951, n_28137, n37950);
  and g63056 (n37952, pi0660, n_27958);
  not g63057 (n_28138, n37951);
  and g63058 (n37953, n_28138, n37952);
  not g63059 (n_28139, n37947);
  not g63060 (n_28140, n37953);
  and g63061 (n37954, n_28139, n_28140);
  not g63062 (n_28141, n37954);
  and g63063 (n37955, pi0785, n_28141);
  and g63064 (n37956, n_11964, n_28132);
  not g63065 (n_28142, n37955);
  not g63066 (n_28143, n37956);
  and g63067 (n37957, n_28142, n_28143);
  not g63068 (n_28144, n37957);
  and g63069 (n37958, n_11984, n_28144);
  and g63070 (n37959, pi0618, n37562);
  not g63071 (n_28145, n37959);
  and g63072 (n37960, n_11413, n_28145);
  not g63073 (n_28146, n37958);
  and g63074 (n37961, n_28146, n37960);
  and g63075 (n37962, n_11412, n_27967);
  not g63076 (n_28147, n37961);
  and g63077 (n37963, n_28147, n37962);
  and g63078 (n37964, n_11984, n37562);
  and g63079 (n37965, pi0618, n_28144);
  not g63080 (n_28148, n37964);
  and g63081 (n37966, pi1154, n_28148);
  not g63082 (n_28149, n37965);
  and g63083 (n37967, n_28149, n37966);
  and g63084 (n37968, pi0627, n_27968);
  not g63085 (n_28150, n37967);
  and g63086 (n37969, n_28150, n37968);
  not g63087 (n_28151, n37963);
  not g63088 (n_28152, n37969);
  and g63089 (n37970, n_28151, n_28152);
  not g63090 (n_28153, n37970);
  and g63091 (n37971, pi0781, n_28153);
  and g63092 (n37972, n_11981, n_28144);
  not g63093 (n_28154, n37971);
  not g63094 (n_28155, n37972);
  and g63095 (n37973, n_28154, n_28155);
  and g63096 (n37974, n_12315, n37973);
  not g63097 (n_28156, n37973);
  and g63098 (n37975, n_11821, n_28156);
  and g63099 (n37976, pi0619, n37565);
  not g63100 (n_28157, n37976);
  and g63101 (n37977, n_11405, n_28157);
  not g63102 (n_28158, n37975);
  and g63103 (n37978, n_28158, n37977);
  and g63104 (n37979, n_11403, n_27977);
  not g63105 (n_28159, n37978);
  and g63106 (n37980, n_28159, n37979);
  and g63107 (n37981, pi0619, n_28156);
  and g63108 (n37982, n_11821, n37565);
  not g63109 (n_28160, n37982);
  and g63110 (n37983, pi1159, n_28160);
  not g63111 (n_28161, n37981);
  and g63112 (n37984, n_28161, n37983);
  and g63113 (n37985, pi0648, n_27978);
  not g63114 (n_28162, n37984);
  and g63115 (n37986, n_28162, n37985);
  not g63116 (n_28163, n37980);
  and g63117 (n37987, pi0789, n_28163);
  not g63118 (n_28164, n37986);
  and g63119 (n37988, n_28164, n37987);
  not g63120 (n_28165, n37974);
  and g63121 (n37989, n17970, n_28165);
  not g63122 (n_28166, n37988);
  and g63123 (n37990, n_28166, n37989);
  and g63124 (n37991, n16635, n_27769);
  not g63125 (n_28167, n37566);
  not g63126 (n_28168, n37991);
  and g63127 (n37992, n_28167, n_28168);
  not g63128 (n_28169, n37992);
  and g63129 (n37993, n17871, n_28169);
  and g63130 (n37994, n_12320, n37459);
  not g63131 (n_28170, n37749);
  and g63132 (n37995, pi0626, n_28170);
  not g63133 (n_28171, n37994);
  and g63134 (n37996, n16628, n_28171);
  not g63135 (n_28172, n37995);
  and g63136 (n37997, n_28172, n37996);
  and g63137 (n37998, pi0626, n37459);
  and g63138 (n37999, n_12320, n_28170);
  not g63139 (n_28173, n37998);
  and g63140 (n38000, n16629, n_28173);
  not g63141 (n_28174, n37999);
  and g63142 (n38001, n_28174, n38000);
  not g63143 (n_28175, n37993);
  not g63144 (n_28176, n37997);
  and g63145 (n38002, n_28175, n_28176);
  not g63146 (n_28177, n38001);
  and g63147 (n38003, n_28177, n38002);
  not g63148 (n_28178, n38003);
  and g63149 (n38004, pi0788, n_28178);
  not g63150 (n_28179, n38004);
  and g63151 (n38005, n_14638, n_28179);
  not g63152 (n_28180, n37990);
  and g63153 (n38006, n_28180, n38005);
  not g63154 (n_28181, n37759);
  not g63155 (n_28182, n38006);
  and g63156 (n38007, n_28181, n_28182);
  not g63157 (n_28183, n38007);
  and g63158 (n38008, n_14387, n_28183);
  and g63159 (n38009, n_12375, n37580);
  and g63160 (n38010, n_12368, n37751);
  and g63161 (n38011, n17779, n37459);
  not g63162 (n_28184, n38010);
  not g63163 (n_28185, n38011);
  and g63164 (n38012, n_28184, n_28185);
  not g63165 (n_28186, n38012);
  and g63166 (n38013, n_14548, n_28186);
  and g63167 (n38014, pi0630, n37576);
  not g63168 (n_28187, n38009);
  not g63169 (n_28188, n38014);
  and g63170 (n38015, n_28187, n_28188);
  not g63171 (n_28189, n38013);
  and g63172 (n38016, n_28189, n38015);
  not g63173 (n_28190, n38016);
  and g63174 (n38017, pi0787, n_28190);
  not g63175 (n_28191, n38008);
  not g63176 (n_28192, n38017);
  and g63177 (n38018, n_28191, n_28192);
  and g63178 (n38019, pi0644, n38018);
  not g63179 (n_28193, n37584);
  and g63180 (n38020, pi0715, n_28193);
  not g63181 (n_28194, n38019);
  and g63182 (n38021, n_28194, n38020);
  and g63183 (n38022, n17804, n_27769);
  and g63184 (n38023, n_12392, n38012);
  not g63185 (n_28195, n38022);
  not g63186 (n_28196, n38023);
  and g63187 (n38024, n_28195, n_28196);
  not g63188 (n_28197, n38024);
  and g63189 (n38025, pi0644, n_28197);
  and g63190 (n38026, n_11819, n_27769);
  not g63191 (n_28198, n38026);
  and g63192 (n38027, n_12395, n_28198);
  not g63193 (n_28199, n38025);
  and g63194 (n38028, n_28199, n38027);
  not g63195 (n_28200, n38028);
  and g63196 (n38029, pi1160, n_28200);
  not g63197 (n_28201, n38021);
  and g63198 (n38030, n_28201, n38029);
  and g63199 (n38031, pi0644, n37583);
  and g63200 (n38032, n_11819, n38018);
  not g63201 (n_28202, n38031);
  and g63202 (n38033, n_12395, n_28202);
  not g63203 (n_28203, n38032);
  and g63204 (n38034, n_28203, n38033);
  and g63205 (n38035, n_11819, n_28197);
  and g63206 (n38036, pi0644, n_27769);
  not g63207 (n_28204, n38036);
  and g63208 (n38037, pi0715, n_28204);
  not g63209 (n_28205, n38035);
  and g63210 (n38038, n_28205, n38037);
  not g63211 (n_28206, n38038);
  and g63212 (n38039, n_12405, n_28206);
  not g63213 (n_28207, n38034);
  and g63214 (n38040, n_28207, n38039);
  not g63215 (n_28208, n38030);
  not g63216 (n_28209, n38040);
  and g63217 (n38041, n_28208, n_28209);
  not g63218 (n_28210, n38041);
  and g63219 (n38042, pi0790, n_28210);
  and g63220 (n38043, n_12411, n38018);
  not g63221 (n_28211, n38042);
  not g63222 (n_28212, n38043);
  and g63223 (n38044, n_28211, n_28212);
  not g63224 (n_28213, n38044);
  and g63225 (n38045, n_4226, n_28213);
  and g63226 (n38046, n_219, po1038);
  not g63227 (n_28214, n38045);
  not g63228 (n_28215, n38046);
  and g63229 (po0381, n_28214, n_28215);
  and g63230 (n38048, n2547, n2625);
  and g63231 (n38049, n3330, n38048);
  and g63232 (n38050, n_158, n38049);
  not g63233 (n_28216, n38050);
  and g63234 (n38051, n_824, n_28216);
  and g63235 (n38052, pi0062, n38049);
  and g63236 (n38053, n2534, n38048);
  not g63237 (n_28217, n38053);
  and g63238 (n38054, pi0054, n_28217);
  and g63239 (n38055, pi0092, n2533);
  and g63240 (n38056, n38048, n38055);
  and g63241 (n38057, n_3066, n6263);
  not g63242 (n_28218, n38057);
  and g63243 (n38058, n_186, n_28218);
  not g63244 (n_28219, n38058);
  and g63245 (n38059, n7301, n_28219);
  not g63246 (n_28220, n38059);
  and g63247 (n38060, pi0075, n_28220);
  and g63248 (n38061, pi0087, n38048);
  and g63249 (n38062, n6286, n_28219);
  and g63250 (n38063, pi0038, n_186);
  and g63251 (n38064, pi0039, n2547);
  and g63252 (n38065, n_345, n_523);
  not g63253 (n_28221, n38065);
  and g63254 (n38066, pi0137, n_28221);
  not g63255 (n_28222, n38066);
  and g63256 (n38067, n_480, n_28222);
  not g63257 (n_28223, n38067);
  and g63258 (n38068, n_4, n_28223);
  and g63259 (n38069, n2517, n11417);
  not g63260 (n_28224, n38069);
  and g63261 (n38070, n2738, n_28224);
  and g63262 (n38071, n_186, n2713);
  not g63263 (n_28225, n38070);
  and g63264 (n38072, n_28225, n38071);
  not g63265 (n_28226, n11417);
  and g63266 (n38073, n3168, n_28226);
  and g63267 (n38074, n_473, n38073);
  not g63268 (n_28227, n38074);
  and g63269 (n38075, n2746, n_28227);
  not g63270 (n_28228, n38075);
  and g63271 (n38076, n2744, n_28228);
  not g63272 (n_28229, n38076);
  and g63273 (n38077, n_330, n_28229);
  not g63274 (n_28230, n38077);
  and g63275 (n38078, n_144, n_28230);
  not g63276 (n_28231, n38078);
  and g63277 (n38079, n3088, n_28231);
  not g63278 (n_28232, n38072);
  and g63279 (n38080, pi0332, n_28232);
  not g63280 (n_28233, n38079);
  and g63281 (n38081, n_28233, n38080);
  not g63282 (n_28234, n38068);
  not g63283 (n_28235, n38081);
  and g63284 (n38082, n_28234, n_28235);
  not g63285 (n_28236, n38082);
  and g63286 (n38083, pi0210, n_28236);
  and g63287 (n38084, n2922, n_28225);
  not g63288 (n_28237, n38084);
  and g63289 (n38085, pi1093, n_28237);
  and g63290 (n38086, n2922, n2933);
  and g63291 (n38087, n2517, n_4103);
  and g63292 (n38088, n_516, n38087);
  not g63293 (n_28238, n38088);
  and g63294 (n38089, n_142, n_28238);
  not g63295 (n_28239, n38089);
  and g63296 (n38090, n38086, n_28239);
  not g63297 (n_28240, n38090);
  and g63298 (n38091, n_3206, n_28240);
  and g63299 (n38092, n_7455, n38084);
  and g63300 (n38093, n11416, n38087);
  and g63301 (n38094, n38086, n38093);
  not g63302 (n_28241, n38092);
  not g63303 (n_28242, n38094);
  and g63304 (n38095, n_28241, n_28242);
  and g63305 (n38096, n38091, n38095);
  not g63306 (n_28243, n38085);
  not g63307 (n_28244, n38096);
  and g63308 (n38097, n_28243, n_28244);
  not g63309 (n_28245, n38097);
  and g63310 (n38098, n11549, n_28245);
  and g63311 (n38099, n_485, n_28229);
  not g63312 (n_28246, n38099);
  and g63313 (n38100, n_144, n_28246);
  not g63314 (n_28247, n38100);
  and g63315 (n38101, n_345, n_28247);
  not g63316 (n_28248, n38101);
  and g63317 (n38102, pi0137, n_28248);
  and g63318 (n38103, n_7455, n3023);
  not g63319 (n_28249, n38103);
  and g63320 (n38104, n38091, n_28249);
  and g63321 (n38105, n_540, n38087);
  not g63322 (n_28250, n38105);
  and g63323 (n38106, n_142, n_28250);
  not g63324 (n_28251, n38106);
  and g63325 (n38107, n38086, n_28251);
  and g63326 (n38108, pi1093, n_28249);
  not g63327 (n_28252, n38107);
  and g63328 (n38109, n_28252, n38108);
  not g63329 (n_28253, n38104);
  not g63330 (n_28254, n38109);
  and g63331 (n38110, n_28253, n_28254);
  not g63332 (n_28255, n38110);
  and g63333 (n38111, n11517, n_28255);
  and g63334 (n38112, n38095, n38111);
  not g63335 (n_28256, n38098);
  not g63336 (n_28257, n38112);
  and g63337 (n38113, n_28256, n_28257);
  not g63338 (n_28258, n38102);
  and g63339 (n38114, n_28258, n38113);
  not g63340 (n_28259, n38114);
  and g63341 (n38115, pi0332, n_28259);
  and g63342 (n38116, n_345, n_530);
  not g63343 (n_28260, n38116);
  and g63344 (n38117, pi0137, n_28260);
  and g63345 (n38118, pi1093, n_560);
  not g63346 (n_28261, n38118);
  and g63347 (n38119, n_28253, n_28261);
  not g63348 (n_28262, n38119);
  and g63349 (n38120, n11549, n_28262);
  not g63350 (n_28263, n38111);
  not g63351 (n_28264, n38120);
  and g63352 (n38121, n_28263, n_28264);
  not g63353 (n_28265, n38117);
  and g63354 (n38122, n_28265, n38121);
  not g63355 (n_28266, n38122);
  and g63356 (n38123, n_4, n_28266);
  not g63357 (n_28267, n38115);
  not g63358 (n_28268, n38123);
  and g63359 (n38124, n_28267, n_28268);
  and g63360 (n38125, n_272, n38124);
  and g63361 (n38126, n_186, n_28237);
  not g63362 (n_28269, n38126);
  and g63363 (n38127, n_28258, n_28269);
  not g63364 (n_28270, n38127);
  and g63365 (n38128, pi0332, n_28270);
  and g63366 (n38129, n_561, n_28265);
  not g63367 (n_28271, n38129);
  and g63368 (n38130, n_4, n_28271);
  not g63369 (n_28272, n38128);
  not g63370 (n_28273, n38130);
  and g63371 (n38131, n_28272, n_28273);
  and g63372 (n38132, n2640, n38131);
  not g63373 (n_28274, n38125);
  and g63374 (n38133, n_271, n_28274);
  not g63375 (n_28275, n38132);
  and g63376 (n38134, n_28275, n38133);
  not g63377 (n_28276, n38083);
  and g63378 (n38135, pi0299, n_28276);
  not g63379 (n_28277, n38134);
  and g63380 (n38136, n_28277, n38135);
  and g63381 (n38137, pi0198, n_28236);
  and g63382 (n38138, n6260, n38131);
  and g63383 (n38139, n_3261, n38124);
  not g63384 (n_28278, n38138);
  and g63385 (n38140, n_305, n_28278);
  not g63386 (n_28279, n38139);
  and g63387 (n38141, n_28279, n38140);
  not g63388 (n_28280, n38137);
  and g63389 (n38142, n_234, n_28280);
  not g63390 (n_28281, n38141);
  and g63391 (n38143, n_28281, n38142);
  not g63392 (n_28282, n38136);
  not g63393 (n_28283, n38143);
  and g63394 (n38144, n_28282, n_28283);
  not g63395 (n_28284, n38144);
  and g63396 (n38145, n_162, n_28284);
  not g63397 (n_28285, n38064);
  and g63398 (n38146, n_161, n_28285);
  not g63399 (n_28286, n38145);
  and g63400 (n38147, n_28286, n38146);
  not g63401 (n_28287, n38063);
  and g63402 (n38148, n6137, n_28287);
  not g63403 (n_28288, n38147);
  and g63404 (n38149, n_28288, n38148);
  not g63405 (n_28289, n38062);
  not g63406 (n_28290, n38149);
  and g63407 (n38150, n_28289, n_28290);
  not g63408 (n_28291, n38150);
  and g63409 (n38151, n_172, n_28291);
  not g63410 (n_28292, n38061);
  and g63411 (n38152, n_171, n_28292);
  not g63412 (n_28293, n38151);
  and g63413 (n38153, n_28293, n38152);
  not g63414 (n_28294, n38060);
  and g63415 (n38154, n_174, n_28294);
  not g63416 (n_28295, n38153);
  and g63417 (n38155, n_28295, n38154);
  not g63418 (n_28296, n38056);
  and g63419 (n38156, n_167, n_28296);
  not g63420 (n_28297, n38155);
  and g63421 (n38157, n_28297, n38156);
  not g63422 (n_28298, n38054);
  and g63423 (n38158, n_168, n_28298);
  not g63424 (n_28299, n38157);
  and g63425 (n38159, n_28299, n38158);
  and g63426 (n38160, pi0074, n6128);
  and g63427 (n38161, n38048, n38160);
  not g63428 (n_28300, n38161);
  and g63429 (n38162, n_176, n_28300);
  not g63430 (n_28301, n38159);
  and g63431 (n38163, n_28301, n38162);
  not g63432 (n_28302, n38163);
  and g63433 (n38164, n7348, n_28302);
  and g63434 (n38165, pi0056, n2536);
  and g63435 (n38166, n38048, n38165);
  not g63436 (n_28303, n38164);
  not g63437 (n_28304, n38166);
  and g63438 (n38167, n_28303, n_28304);
  not g63439 (n_28305, n38167);
  and g63440 (n38168, n_158, n_28305);
  not g63441 (n_28306, n38052);
  and g63442 (n38169, n3328, n_28306);
  not g63443 (n_28307, n38168);
  and g63444 (n38170, n_28307, n38169);
  not g63445 (n_28308, n38051);
  and g63446 (n38171, n_3030, n_28308);
  not g63447 (n_28309, n38170);
  and g63448 (po0382, n_28309, n38171);
  and g63449 (n38173, pi0228, pi0231);
  not g63450 (n_28311, n38173);
  and g63451 (n38174, n_4038, n_28311);
  not g63452 (n_28312, n38174);
  and g63453 (n38175, pi0056, n_28312);
  and g63454 (n38176, pi0055, n_28311);
  not g63455 (n_28313, n7364);
  and g63456 (n38177, n_28313, n_28311);
  not g63457 (n_28314, n38177);
  and g63458 (n38178, pi0074, n_28314);
  and g63459 (n38179, pi0054, n_28311);
  and g63460 (n38180, n_9345, n_28311);
  not g63461 (n_28315, n38180);
  and g63462 (n38181, pi0075, n_28315);
  and g63463 (n38182, pi0087, n_28311);
  and g63464 (n38183, n_4043, n38182);
  and g63465 (n38184, n_9347, n_28311);
  not g63466 (n_28316, n38184);
  and g63467 (n38185, pi0100, n_28316);
  not g63468 (n_28317, n2730);
  and g63469 (n38186, n_28317, n_643);
  not g63470 (n_28318, n38186);
  and g63471 (n38187, n_139, n_28318);
  not g63472 (n_28319, n38187);
  and g63473 (n38188, n_138, n_28319);
  not g63474 (n_28320, n38188);
  and g63475 (n38189, n2748, n_28320);
  not g63476 (n_28321, n38189);
  and g63477 (n38190, n3168, n_28321);
  not g63478 (n_28322, n38190);
  and g63479 (n38191, n2746, n_28322);
  not g63480 (n_28323, n38191);
  and g63481 (n38192, n2744, n_28323);
  not g63482 (n_28324, n38192);
  and g63483 (n38193, n_3071, n_28324);
  not g63484 (n_28325, n38193);
  and g63485 (n38194, n_144, n_28325);
  not g63486 (n_28326, n38194);
  and g63487 (n38195, n2742, n_28326);
  not g63488 (n_28327, n38195);
  and g63489 (n38196, n_162, n_28327);
  and g63490 (n38197, n_161, n_880);
  not g63491 (n_28328, n38196);
  and g63492 (n38198, n_28328, n38197);
  and g63493 (n38199, n_188, n38198);
  not g63494 (n_28329, n38199);
  and g63495 (n38200, n_28311, n_28329);
  not g63496 (n_28330, n38200);
  and g63497 (n38201, n_164, n_28330);
  not g63498 (n_28331, n38185);
  and g63499 (n38202, n_172, n_28331);
  not g63500 (n_28332, n38201);
  and g63501 (n38203, n_28332, n38202);
  not g63502 (n_28333, n38183);
  and g63503 (n38204, n_171, n_28333);
  not g63504 (n_28334, n38203);
  and g63505 (n38205, n_28334, n38204);
  not g63506 (n_28335, n38181);
  and g63507 (n38206, n_174, n_28335);
  not g63508 (n_28336, n38205);
  and g63509 (n38207, n_28336, n38206);
  and g63510 (n38208, pi0092, n_28311);
  and g63511 (n38209, n_4041, n38208);
  not g63512 (n_28337, n38207);
  not g63513 (n_28338, n38209);
  and g63514 (n38210, n_28337, n_28338);
  not g63515 (n_28339, n38210);
  and g63516 (n38211, n_167, n_28339);
  not g63517 (n_28340, n38179);
  and g63518 (n38212, n_168, n_28340);
  not g63519 (n_28341, n38211);
  and g63520 (n38213, n_28341, n38212);
  not g63521 (n_28342, n38178);
  and g63522 (n38214, n_176, n_28342);
  not g63523 (n_28343, n38213);
  and g63524 (n38215, n_28343, n38214);
  not g63525 (n_28344, n38176);
  and g63526 (n38216, n_157, n_28344);
  not g63527 (n_28345, n38215);
  and g63528 (n38217, n_28345, n38216);
  not g63529 (n_28346, n38175);
  and g63530 (n38218, n_158, n_28346);
  not g63531 (n_28347, n38217);
  and g63532 (n38219, n_28347, n38218);
  and g63533 (n38220, pi0062, n_28311);
  and g63534 (n38221, n_4036, n38220);
  not g63535 (n_28348, n38219);
  not g63536 (n_28349, n38221);
  and g63537 (n38222, n_28348, n_28349);
  not g63538 (n_28350, n38222);
  and g63539 (n38223, n3328, n_28350);
  and g63540 (n38224, n_824, n_28311);
  not g63541 (n_28351, n38223);
  not g63542 (n_28352, n38224);
  and g63543 (po0383, n_28351, n_28352);
  and g63544 (n38226, n13080, n_8712);
  and g63545 (n38227, n6480, n38226);
  not g63546 (n_28353, n38227);
  and g63547 (n38228, n_3286, n_28353);
  not g63548 (n_28354, n38228);
  and g63549 (n38229, pi1093, n_28354);
  and g63550 (n38230, n2708, n6420);
  and g63551 (n38231, n_109, n_355);
  not g63552 (n_28355, n38231);
  and g63553 (n38232, n38230, n_28355);
  not g63554 (n_28356, n38232);
  and g63555 (n38233, n_134, n_28356);
  and g63556 (n38234, n11022, n38230);
  and g63557 (n38235, n_7196, n38234);
  not g63558 (n_28357, n8903);
  and g63559 (n38236, n_28357, n38233);
  not g63560 (n_28358, n38235);
  and g63561 (n38237, n_28358, n38236);
  not g63562 (n_28359, n38237);
  and g63563 (n38238, n6480, n_28359);
  not g63564 (n_28360, n38229);
  not g63565 (n_28361, n38238);
  and g63566 (n38239, n_28360, n_28361);
  not g63567 (n_28362, n38234);
  and g63568 (n38240, n38233, n_28362);
  not g63569 (n_28363, n38240);
  and g63570 (n38241, n6480, n_28363);
  not g63571 (n_28364, n38241);
  and g63572 (n38242, n10074, n_28364);
  and g63573 (n38243, n_6605, n11022);
  and g63574 (n38244, n2754, n11031);
  and g63575 (n38245, n11029, n38244);
  not g63576 (n_28365, n38243);
  and g63577 (n38246, n38231, n_28365);
  not g63578 (n_28366, n38245);
  and g63579 (n38247, n_28366, n38246);
  not g63580 (n_28367, n38247);
  and g63581 (n38248, n38230, n_28367);
  not g63582 (n_28368, n38248);
  and g63583 (n38249, n_134, n_28368);
  not g63584 (n_28369, n38249);
  and g63585 (n38250, n6480, n_28369);
  not g63586 (n_28370, n6215);
  and g63587 (n38251, pi0829, n_28370);
  not g63588 (n_28371, n38250);
  and g63589 (n38252, n_28371, n38251);
  not g63590 (n_28372, n38239);
  not g63591 (n_28373, n38242);
  and g63592 (n38253, n_28372, n_28373);
  not g63593 (n_28374, n38252);
  and g63594 (n38254, n_28374, n38253);
  not g63595 (n_28375, n38254);
  and g63596 (n38255, n_162, n_28375);
  not g63597 (n_28376, n11471);
  or g63598 (po0384, n_28376, n38255);
  and g63599 (n38257, n_162, pi0228);
  not g63600 (n_28377, n11420);
  not g63601 (n_28378, n11425);
  and g63602 (n38258, n_28377, n_28378);
  not g63603 (n_28379, n38258);
  and g63604 (n38259, pi0039, n_28379);
  and g63605 (n38260, n6391, n38259);
  not g63606 (n_28380, n2930);
  not g63607 (n_28381, n8904);
  and g63608 (n38261, n_28380, n_28381);
  not g63614 (n_28383, n38260);
  not g63615 (n_28384, n38265);
  and g63616 (n38266, n_28383, n_28384);
  not g63617 (n_28385, n38266);
  and g63618 (n38267, n10200, n_28385);
  or g63619 (po0385, n38257, n38267);
  and g63620 (n38269, n_3039, n10197);
  and g63621 (n38270, pi0120, n6218);
  not g63622 (n_28386, n38270);
  and g63623 (n38271, n16652, n_28386);
  not g63624 (n_28387, n35677);
  not g63625 (n_28388, n38271);
  and g63626 (n38272, n_28387, n_28388);
  not g63627 (n_28389, n38272);
  and g63628 (n38273, n_3119, n_28389);
  and g63629 (n38274, n_3120, n16652);
  not g63630 (n_28390, n38274);
  and g63631 (n38275, n_28388, n_28390);
  not g63632 (n_28391, n38275);
  and g63633 (n38276, n6205, n_28391);
  not g63634 (n_28392, n38273);
  and g63635 (n38277, pi0223, n_28392);
  not g63636 (n_28393, n38276);
  and g63637 (n38278, n_28393, n38277);
  and g63638 (n38279, n2603, n16652);
  and g63639 (n38280, n_3130, n7517);
  and g63640 (n38281, n16661, n38280);
  not g63641 (n_28394, n38280);
  and g63642 (n38282, n16649, n_28394);
  not g63643 (n_28395, n38281);
  and g63644 (n38283, pi1091, n_28395);
  not g63645 (n_28396, n38282);
  and g63646 (n38284, n_28396, n38283);
  and g63647 (n38285, n6383, n16661);
  not g63648 (n_28397, n6383);
  and g63649 (n38286, n_28397, n16649);
  not g63650 (n_28398, n38285);
  and g63651 (n38287, n_3128, n_28398);
  not g63652 (n_28399, n38286);
  and g63653 (n38288, n_28399, n38287);
  not g63654 (n_28400, n38284);
  not g63655 (n_28401, n38288);
  and g63656 (n38289, n_28400, n_28401);
  not g63657 (n_28402, n38289);
  and g63658 (n38290, n_9389, n_28402);
  not g63659 (n_28403, n38290);
  and g63660 (n38291, n_11426, n_28403);
  and g63661 (n38292, n_3140, n38291);
  not g63662 (n_28404, n38292);
  and g63663 (n38293, n_28387, n_28404);
  and g63664 (n38294, n_3119, n38293);
  and g63665 (n38295, n6198, n38291);
  not g63666 (n_28405, n38295);
  and g63667 (n38296, n_28390, n_28405);
  and g63668 (n38297, n6205, n38296);
  not g63669 (n_28406, n38294);
  and g63670 (n38298, n_9349, n_28406);
  not g63671 (n_28407, n38297);
  and g63672 (n38299, n_28407, n38298);
  not g63673 (n_28408, n38279);
  and g63674 (n38300, n_223, n_28408);
  not g63675 (n_28409, n38299);
  and g63676 (n38301, n_28409, n38300);
  not g63677 (n_28410, n38278);
  and g63678 (n38302, n_234, n_28410);
  not g63679 (n_28411, n38301);
  and g63680 (n38303, n_28411, n38302);
  and g63681 (n38304, n_3162, n_28389);
  and g63682 (n38305, n6242, n_28391);
  not g63683 (n_28412, n38304);
  and g63684 (n38306, pi0215, n_28412);
  not g63685 (n_28413, n38305);
  and g63686 (n38307, n_28413, n38306);
  and g63687 (n38308, n_3162, n38293);
  and g63688 (n38309, n6242, n38296);
  not g63689 (n_28414, n38308);
  and g63690 (n38310, n_9350, n_28414);
  not g63691 (n_28415, n38309);
  and g63692 (n38311, n_28415, n38310);
  not g63693 (n_28416, n16825);
  and g63694 (n38312, n_36, n_28416);
  not g63695 (n_28417, n38311);
  and g63696 (n38313, n_28417, n38312);
  not g63697 (n_28418, n38307);
  and g63698 (n38314, pi0299, n_28418);
  not g63699 (n_28419, n38313);
  and g63700 (n38315, n_28419, n38314);
  not g63701 (n_28420, n38303);
  not g63702 (n_28421, n38315);
  and g63703 (n38316, n_28420, n_28421);
  not g63704 (n_28422, n38316);
  and g63705 (n38317, pi0039, n_28422);
  and g63706 (n38318, n6170, n16854);
  not g63707 (n_28423, n16856);
  and g63708 (n38319, n_28423, n38318);
  not g63709 (n_28424, n38319);
  and g63710 (n38320, n_143, n_28424);
  not g63711 (n_28425, n38320);
  and g63712 (n38321, n10289, n_28425);
  not g63713 (n_28426, n38321);
  and g63714 (n38322, pi0252, n_28426);
  and g63715 (n38323, n6277, n_11592);
  not g63716 (n_28427, n38322);
  and g63717 (n38324, n_28427, n38323);
  and g63718 (n38325, n_7462, n16866);
  not g63719 (n_28428, n38324);
  and g63720 (n38326, n_3206, n_28428);
  not g63721 (n_28429, n38325);
  and g63722 (n38327, n_28429, n38326);
  and g63723 (n38328, n_3066, n_3279);
  and g63724 (n38329, n_7196, n16866);
  not g63725 (n_28430, n38329);
  and g63726 (n38330, n_11605, n_28430);
  not g63727 (n_28431, n38330);
  and g63728 (n38331, n38328, n_28431);
  and g63729 (n38332, pi0829, pi1091);
  and g63730 (n38333, n16907, n38332);
  not g63731 (n_28432, n38333);
  and g63732 (n38334, n_3126, n_28432);
  not g63733 (n_28433, n16902);
  and g63734 (n38335, pi0824, n_28433);
  not g63735 (n_28434, n38334);
  and g63736 (n38336, n_3279, n_28434);
  not g63737 (n_28435, n38335);
  and g63738 (n38337, n_28435, n38336);
  not g63739 (n_28436, n16866);
  not g63740 (n_28437, n38337);
  and g63741 (n38338, n_28436, n_28437);
  and g63742 (n38339, n38332, n38334);
  not g63743 (n_28438, n38339);
  and g63744 (n38340, n_28435, n_28438);
  and g63745 (n38341, n2932, n_3279);
  not g63746 (n_28439, n38340);
  and g63747 (n38342, n_28439, n38341);
  not g63748 (n_28440, n38328);
  not g63749 (n_28441, n38338);
  and g63750 (n38343, n_28440, n_28441);
  not g63751 (n_28442, n38342);
  and g63752 (n38344, n_28442, n38343);
  not g63753 (n_28443, n38331);
  and g63754 (n38345, pi1093, n_28443);
  not g63755 (n_28444, n38344);
  and g63756 (n38346, n_28444, n38345);
  not g63757 (n_28445, n38327);
  and g63758 (n38347, n_162, n_28445);
  not g63759 (n_28446, n38346);
  and g63760 (n38348, n_28446, n38347);
  not g63761 (n_28447, n38317);
  and g63762 (n38349, n_161, n_28447);
  not g63763 (n_28448, n38348);
  and g63764 (n38350, n_28448, n38349);
  not g63765 (n_28449, n38350);
  and g63766 (po0387, n38269, n_28449);
  and g63767 (n38352, n_105, n_436);
  not g63768 (n_28450, n38352);
  and g63769 (n38353, n6443, n_28450);
  not g63770 (n_28451, n38353);
  and g63771 (n38354, n2462, n_28451);
  not g63772 (n_28452, n38354);
  and g63773 (n38355, n2873, n_28452);
  not g63774 (n_28453, n38355);
  and g63775 (n38356, n2785, n_28453);
  not g63776 (n_28454, n38356);
  and g63777 (n38357, n2877, n_28454);
  not g63778 (n_28455, n38357);
  and g63779 (n38358, n2719, n_28455);
  not g63780 (n_28456, n38358);
  and g63781 (n38359, n_333, n_28456);
  not g63782 (n_28457, n38359);
  and g63783 (n38360, n_119, n_28457);
  not g63784 (n_28458, n38360);
  and g63785 (n38361, n2783, n_28458);
  not g63786 (n_28459, n38361);
  and g63787 (n38362, n2781, n_28459);
  not g63788 (n_28460, n38362);
  and g63789 (n38363, n_453, n_28460);
  not g63790 (n_28461, n38363);
  and g63791 (n38364, n_123, n_28461);
  not g63792 (n_28462, n38364);
  and g63793 (n38365, n2775, n_28462);
  not g63794 (n_28463, n38365);
  and g63795 (n38366, n2889, n_28463);
  not g63796 (n_28464, n38366);
  and g63797 (n38367, n_459, n_28464);
  not g63798 (n_28465, n38367);
  and g63799 (n38368, n2765, n_28465);
  not g63800 (n_28466, n38368);
  and g63801 (n38369, n2764, n_28466);
  not g63802 (n_28467, n38369);
  and g63803 (n38370, n2757, n_28467);
  not g63804 (n_28468, n38370);
  and g63805 (n38371, n3108, n_28468);
  not g63806 (n_28469, n38371);
  and g63807 (n38372, n2504, n_28469);
  not g63808 (n_28470, n38372);
  and g63809 (n38373, n15635, n_28470);
  not g63810 (n_28471, n38373);
  and g63811 (n38374, n_139, n_28471);
  not g63812 (n_28472, n38374);
  and g63813 (n38375, n_622, n_28472);
  not g63814 (n_28473, n38375);
  and g63815 (n38376, n_138, n_28473);
  not g63816 (n_28474, n38376);
  and g63817 (n38377, n2748, n_28474);
  not g63818 (n_28475, n38377);
  and g63819 (n38378, n3168, n_28475);
  not g63820 (n_28476, n38378);
  and g63821 (n38379, n2746, n_28476);
  and g63822 (n38380, n_6603, n2743);
  not g63823 (n_28477, n38380);
  and g63824 (n38381, n_142, n_28477);
  not g63825 (n_28478, n38379);
  and g63826 (n38382, n_28478, n38381);
  not g63827 (n_28479, n38382);
  and g63828 (n38383, n_875, n_28479);
  not g63829 (n_28480, n38383);
  and g63830 (n38384, n_144, n_28480);
  not g63831 (n_28481, n38384);
  and g63832 (n38385, n_345, n_28481);
  not g63833 (n_28482, n38385);
  and g63834 (n38386, n_162, n_28482);
  not g63835 (n_28483, n7307);
  not g63836 (n_28484, n7309);
  and g63837 (n38387, n_28483, n_28484);
  not g63838 (n_28485, n6217);
  or g63839 (po0950, n_6605, n_28485);
  not g63840 (n_28487, po0950);
  and g63841 (n38389, n6381, n_28487);
  not g63842 (n_28488, n38387);
  and g63843 (n38390, n_28488, n38389);
  and g63844 (n38391, n6185, n11369);
  not g63845 (n_28489, n38390);
  and g63846 (n38392, n_28489, n38391);
  not g63847 (n_28490, n38392);
  and g63848 (n38393, n_880, n_28490);
  not g63849 (n_28491, n38386);
  and g63850 (n38394, n_28491, n38393);
  not g63851 (n_28492, n38394);
  and g63852 (n38395, n_161, n_28492);
  not g63853 (n_28493, n38395);
  and g63854 (n38396, n6137, n_28493);
  not g63855 (n_28494, n6286);
  and g63856 (n38397, n_172, n_28494);
  not g63857 (n_28495, n38396);
  and g63858 (n38398, n_28495, n38397);
  not g63859 (n_28496, n38398);
  and g63860 (n38399, n_3037, n_28496);
  not g63861 (n_28497, n38399);
  and g63862 (n38400, n2569, n_28497);
  not g63863 (n_28498, n38400);
  and g63864 (n38401, n7306, n_28498);
  not g63865 (n_28499, n38401);
  and g63866 (n38402, n_167, n_28499);
  not g63867 (n_28500, n38402);
  and g63868 (n38403, n_4020, n_28500);
  not g63869 (n_28501, n38403);
  and g63870 (n38404, n8879, n_28501);
  not g63871 (n_28502, n38404);
  and g63872 (n38405, n15712, n_28502);
  not g63873 (n_28503, n38405);
  and g63874 (n38406, n_157, n_28503);
  not g63875 (n_28504, n38406);
  and g63876 (n38407, n_3223, n_28504);
  not g63877 (n_28505, n38407);
  and g63878 (n38408, n_158, n_28505);
  not g63879 (n_28506, n38408);
  and g63880 (n38409, n_3227, n_28506);
  not g63881 (n_28507, n38409);
  and g63882 (n38410, n3328, n_28507);
  not g63883 (n_28508, n38410);
  and g63884 (po0389, n6123, n_28508);
  not g63885 (n_28510, pi0230);
  and g63886 (n38412, n_28510, n_25720);
  and g63887 (n38413, n_26538, n_26565);
  not g63888 (n_28511, n38413);
  and g63889 (n38414, n_7075, n_28511);
  not g63890 (n_28512, n38414);
  and g63891 (n38415, pi0219, n_28512);
  not g63892 (n_28513, n38415);
  and g63893 (n38416, po1038, n_28513);
  and g63894 (n38417, pi1142, n_6933);
  and g63895 (n38418, pi0211, pi1143);
  and g63896 (n38419, n_7075, pi1144);
  not g63897 (n_28514, n38418);
  not g63898 (n_28515, n38419);
  and g63899 (n38420, n_28514, n_28515);
  and g63900 (n38421, n_26538, pi0214);
  and g63901 (n38422, pi0212, n_26565);
  not g63902 (n_28516, n38421);
  not g63903 (n_28517, n38422);
  and g63904 (n38423, n_28516, n_28517);
  not g63905 (n_28518, n38420);
  not g63906 (n_28519, n38423);
  and g63907 (n38424, n_28518, n_28519);
  and g63908 (n38425, n_7075, pi1143);
  and g63909 (n38426, n10843, n38425);
  not g63910 (n_28520, n38424);
  not g63911 (n_28521, n38426);
  and g63912 (n38427, n_28520, n_28521);
  not g63913 (n_28522, n38427);
  and g63914 (n38428, n_6791, n_28522);
  not g63915 (n_28523, n38417);
  not g63916 (n_28524, n38428);
  and g63917 (n38429, n_28523, n_28524);
  not g63918 (n_28525, n38429);
  and g63919 (n38430, n38416, n_28525);
  and g63920 (n38431, pi0299, n_28518);
  and g63921 (n38432, pi0199, pi1142);
  not g63922 (n_28526, n38432);
  and g63923 (n38433, n_7045, n_28526);
  and g63924 (n38434, n_7044, pi1144);
  not g63925 (n_28527, n38434);
  and g63926 (n38435, n38433, n_28527);
  and g63927 (n38436, n_7044, pi1143);
  not g63928 (n_28528, n38436);
  and g63929 (n38437, pi0200, n_28528);
  not g63930 (n_28529, n38435);
  not g63931 (n_28530, n38437);
  and g63932 (n38438, n_28529, n_28530);
  not g63933 (n_28531, n38438);
  and g63934 (n38439, n_234, n_28531);
  not g63935 (n_28532, n38439);
  and g63936 (n38440, n_25873, n_28532);
  and g63937 (n38441, pi0207, n_234);
  and g63938 (n38442, n38433, n_28528);
  and g63939 (n38443, n_7044, pi1142);
  not g63940 (n_28533, n38443);
  and g63941 (n38444, pi0200, n_28533);
  not g63942 (n_28534, n38444);
  and g63943 (n38445, n38441, n_28534);
  not g63944 (n_28535, n38442);
  and g63945 (n38446, n_28535, n38445);
  not g63946 (n_28536, n38440);
  not g63947 (n_28537, n38446);
  and g63948 (n38447, n_28536, n_28537);
  not g63949 (n_28538, n38447);
  and g63950 (n38448, pi0208, n_28538);
  and g63951 (n38449, pi0207, n_26242);
  and g63952 (n38450, n38438, n38449);
  not g63953 (n_28539, n38448);
  not g63954 (n_28540, n38450);
  and g63955 (n38451, n_28539, n_28540);
  not g63956 (n_28541, n38451);
  and g63957 (n38452, n_234, n_28541);
  not g63958 (n_28542, n38452);
  and g63959 (n38453, n_26565, n_28542);
  not g63960 (n_28543, n38431);
  and g63961 (n38454, n_28543, n38453);
  and g63962 (n38455, pi0211, pi1142);
  not g63963 (n_28544, n38425);
  not g63964 (n_28545, n38455);
  and g63965 (n38456, n_28544, n_28545);
  not g63966 (n_28546, n38456);
  and g63967 (n38457, pi0299, n_28546);
  not g63968 (n_28547, n38457);
  and g63969 (n38458, pi0214, n_28547);
  and g63970 (n38459, n_28542, n38458);
  not g63971 (n_28548, n38459);
  and g63972 (n38460, pi0212, n_28548);
  not g63973 (n_28549, n38454);
  and g63974 (n38461, n_28549, n38460);
  and g63975 (n38462, n_28543, n_28542);
  not g63976 (n_28550, n38453);
  and g63977 (n38463, n_26538, n_28550);
  not g63978 (n_28551, n38462);
  and g63979 (n38464, n_28551, n38463);
  not g63980 (n_28552, n38461);
  and g63981 (n38465, n_6791, n_28552);
  not g63982 (n_28553, n38464);
  and g63983 (n38466, n_28553, n38465);
  and g63984 (n38467, n_28512, n38452);
  and g63985 (n38468, n_234, n38451);
  and g63986 (n38469, pi0299, n_1311);
  not g63987 (n_28554, n38469);
  and g63988 (n38470, n38414, n_28554);
  not g63989 (n_28555, n38468);
  and g63990 (n38471, n_28555, n38470);
  not g63991 (n_28556, n38467);
  and g63992 (n38472, pi0219, n_28556);
  not g63993 (n_28557, n38471);
  and g63994 (n38473, n_28557, n38472);
  not g63995 (n_28558, n38473);
  and g63996 (n38474, n_4226, n_28558);
  not g63997 (n_28559, n38466);
  and g63998 (n38475, n_28559, n38474);
  not g63999 (n_28560, n38430);
  not g64000 (n_28561, n38475);
  and g64001 (n38476, n_28560, n_28561);
  and g64002 (n38477, pi0213, n38476);
  and g64003 (n38478, n_7075, pi1157);
  and g64004 (n38479, pi0211, pi1156);
  not g64005 (n_28562, n38478);
  not g64006 (n_28563, n38479);
  and g64007 (n38480, n_28562, n_28563);
  not g64008 (n_28564, n38480);
  and g64009 (n38481, pi0214, n_28564);
  not g64010 (n_28565, n38481);
  and g64011 (n38482, n_26538, n_28565);
  and g64012 (n38483, n_7075, pi1156);
  and g64013 (n38484, pi0211, pi1155);
  not g64014 (n_28566, n38483);
  not g64015 (n_28567, n38484);
  and g64016 (n38485, n_28566, n_28567);
  not g64017 (n_28568, n38485);
  and g64018 (n38486, n_26565, n_28568);
  and g64019 (n38487, n_7075, pi1155);
  and g64020 (n38488, pi0211, pi1154);
  not g64021 (n_28569, n38487);
  not g64022 (n_28570, n38488);
  and g64023 (n38489, n_28569, n_28570);
  not g64024 (n_28571, n38489);
  and g64025 (n38490, pi0214, n_28571);
  not g64026 (n_28572, n38486);
  not g64027 (n_28573, n38490);
  and g64028 (n38491, n_28572, n_28573);
  and g64029 (n38492, pi0212, n38491);
  not g64030 (n_28574, n38482);
  not g64031 (n_28575, n38492);
  and g64032 (n38493, n_28574, n_28575);
  not g64033 (n_28576, n38493);
  and g64034 (n38494, n_6791, n_28576);
  and g64035 (n38495, n_7075, pi1154);
  not g64036 (n_28577, n38495);
  and g64037 (n38496, n_26565, n_28577);
  and g64038 (n38497, n_7075, pi1153);
  not g64039 (n_28578, n38497);
  and g64040 (n38498, n10843, n_28578);
  and g64041 (n38499, n_7075, pi0214);
  and g64042 (n38500, pi1155, n38499);
  not g64043 (n_28579, n38500);
  and g64044 (n38501, n_26538, n_28579);
  not g64045 (n_28580, n38496);
  not g64046 (n_28581, n38498);
  and g64047 (n38502, n_28580, n_28581);
  not g64048 (n_28582, n38501);
  and g64049 (n38503, n_28582, n38502);
  not g64050 (n_28583, n38503);
  and g64051 (n38504, pi0219, n_28583);
  not g64052 (n_28584, n38504);
  and g64053 (n38505, po1038, n_28584);
  not g64054 (n_28585, n38494);
  and g64055 (n38506, n_28585, n38505);
  not g64056 (n_28586, n38506);
  and g64057 (n38507, n_26557, n_28586);
  and g64058 (n38508, n_6791, pi0299);
  and g64059 (n38509, n38493, n38508);
  and g64060 (n38510, pi0299, pi1155);
  and g64061 (n38511, n38421, n38510);
  and g64062 (n38512, pi0299, pi1153);
  not g64063 (n_28587, n38512);
  and g64064 (n38513, pi0214, n_28587);
  and g64065 (n38514, pi0299, pi1154);
  not g64066 (n_28588, n38514);
  and g64067 (n38515, n_26565, n_28588);
  not g64068 (n_28589, n38513);
  and g64069 (n38516, pi0212, n_28589);
  not g64070 (n_28590, n38515);
  and g64071 (n38517, n_28590, n38516);
  not g64072 (n_28591, n38511);
  not g64073 (n_28592, n38517);
  and g64074 (n38518, n_28591, n_28592);
  and g64075 (n38519, n_7075, pi0219);
  not g64076 (n_28593, n38518);
  and g64077 (n38520, n_28593, n38519);
  not g64078 (n_28594, n38509);
  not g64079 (n_28595, n38520);
  and g64080 (n38521, n_28594, n_28595);
  and g64081 (n38522, n_28542, n38521);
  not g64082 (n_28596, n38522);
  and g64083 (n38523, n_4226, n_28596);
  not g64084 (n_28597, n38523);
  and g64085 (n38524, n38507, n_28597);
  not g64086 (n_28598, n38524);
  and g64087 (n38525, pi0209, n_28598);
  not g64088 (n_28599, n38477);
  and g64089 (n38526, n_28599, n38525);
  and g64090 (n38527, n_7075, n10843);
  and g64091 (n38528, pi0299, n_1124);
  and g64092 (n38529, n_7045, pi1155);
  and g64093 (n38530, pi0199, n38529);
  and g64094 (n38531, n_234, n38530);
  not g64095 (n_28600, n38531);
  and g64096 (n38532, n_11794, n_28600);
  not g64097 (n_28601, n11444);
  and g64098 (n38533, n_234, n_28601);
  not g64099 (n_28602, n38530);
  and g64100 (n38534, pi1156, n_28602);
  and g64101 (n38535, n38533, n38534);
  not g64102 (n_28603, n38532);
  not g64103 (n_28604, n38535);
  and g64104 (n38536, n_28603, n_28604);
  and g64105 (n38537, pi0207, n38536);
  not g64106 (n_28605, n38537);
  and g64107 (n38538, n_234, n_28605);
  not g64108 (n_28606, n38538);
  and g64109 (n38539, n_26242, n_28606);
  and g64110 (n38540, n_11810, n38539);
  not g64111 (n_28607, n38528);
  and g64112 (n38541, n_28607, n38540);
  and g64113 (n38542, n_26242, pi1157);
  and g64114 (n38543, pi0299, pi1143);
  and g64115 (n38544, n_11768, n_7047);
  and g64116 (n38545, pi0200, n_234);
  not g64117 (n_28608, n38545);
  and g64118 (n38546, pi1155, n_28608);
  not g64119 (n_28609, n38544);
  not g64120 (n_28610, n38546);
  and g64121 (n38547, n_28609, n_28610);
  and g64122 (n38548, pi0199, n_11768);
  and g64123 (n38549, pi0199, pi0200);
  not g64124 (n_28611, n38549);
  and g64125 (n38550, n_234, n_28611);
  not g64126 (n_28612, n38548);
  and g64127 (n38551, pi1156, n_28612);
  and g64128 (n38552, n38550, n38551);
  not g64129 (n_28613, n38552);
  and g64130 (n38553, n38547, n_28613);
  and g64131 (n38554, pi0207, n_28607);
  not g64132 (n_28614, n38553);
  and g64133 (n38555, n_28614, n38554);
  not g64134 (n_28615, n38543);
  not g64135 (n_28616, n38555);
  and g64136 (n38556, n_28615, n_28616);
  not g64137 (n_28617, n38556);
  and g64138 (n38557, n38542, n_28617);
  not g64139 (n_28618, n38550);
  and g64140 (n38558, pi1153, n_28618);
  not g64141 (n_28619, n38558);
  and g64142 (n38559, pi1154, n_28619);
  and g64143 (n38560, n11384, n38529);
  and g64144 (n38561, n_7046, n_28611);
  and g64145 (n38562, n_11757, n_7385);
  and g64146 (n38563, pi1154, n38561);
  not g64147 (n_28620, n38562);
  and g64148 (n38564, n_28620, n38563);
  not g64149 (n_28621, n38560);
  not g64150 (n_28622, n38564);
  and g64151 (n38565, n_28621, n_28622);
  not g64152 (n_28623, n38565);
  and g64153 (n38566, n38559, n_28623);
  and g64154 (n38567, n_7044, n_11768);
  and g64155 (n38568, n_7045, n_234);
  and g64156 (n38569, pi0199, n_11757);
  not g64157 (n_28624, n38569);
  and g64158 (n38570, n38568, n_28624);
  not g64159 (n_28625, n38567);
  and g64160 (n38571, n_11413, n_28625);
  and g64161 (n38572, n38570, n38571);
  not g64162 (n_28626, n38566);
  not g64163 (n_28627, n38572);
  and g64164 (n38573, n_28626, n_28627);
  and g64165 (n38574, pi0207, n38573);
  and g64166 (n38575, n_28615, n38574);
  and g64167 (n38576, n_7044, pi1155);
  and g64168 (n38577, n38545, n38576);
  not g64169 (n_28628, n38577);
  and g64170 (n38578, n_11413, n_28628);
  and g64171 (n38579, n_28615, n38578);
  and g64172 (n38580, n_11768, n38543);
  not g64173 (n_28629, n38561);
  and g64174 (n38581, n_234, n_28629);
  not g64175 (n_28630, n38581);
  and g64176 (n38582, pi1155, n_28630);
  and g64177 (n38583, n_28607, n38582);
  and g64178 (n38584, n_7045, n_11768);
  and g64179 (n38585, n11373, n38584);
  not g64180 (n_28631, n38585);
  and g64181 (n38586, pi1154, n_28631);
  not g64182 (n_28632, n38580);
  and g64183 (n38587, n_28632, n38586);
  not g64184 (n_28633, n38583);
  and g64185 (n38588, n_28633, n38587);
  not g64186 (n_28634, n38579);
  and g64187 (n38589, n_11794, n_28634);
  not g64188 (n_28635, n38588);
  and g64189 (n38590, n_28635, n38589);
  not g64190 (n_28636, n38576);
  and g64191 (n38591, pi0200, n_28636);
  not g64192 (n_28637, n38591);
  and g64193 (n38592, n_234, n_28637);
  not g64194 (n_28638, n38592);
  and g64195 (n38593, pi1154, n_28638);
  and g64196 (n38594, n_28615, n38593);
  not g64197 (n_28639, n11373);
  and g64198 (n38595, pi1155, n_28639);
  not g64199 (n_28640, n38595);
  and g64200 (n38596, n_28609, n_28640);
  not g64201 (n_28641, n38596);
  and g64202 (n38597, n_28607, n_28641);
  not g64203 (n_28642, n38597);
  and g64204 (n38598, n_11413, n_28642);
  not g64205 (n_28643, n38594);
  and g64206 (n38599, pi1156, n_28643);
  not g64207 (n_28644, n38598);
  and g64208 (n38600, n_28644, n38599);
  not g64209 (n_28645, n38590);
  not g64210 (n_28646, n38600);
  and g64211 (n38601, n_28645, n_28646);
  and g64212 (n38602, n_25873, n38601);
  not g64213 (n_28647, n38575);
  and g64214 (n38603, pi0208, n_28647);
  not g64215 (n_28648, n38602);
  and g64216 (n38604, n_28648, n38603);
  not g64217 (n_28649, n38541);
  not g64218 (n_28650, n38557);
  and g64219 (n38605, n_28649, n_28650);
  not g64220 (n_28651, n38604);
  and g64221 (n38606, n_28651, n38605);
  and g64222 (n38607, n38527, n38606);
  and g64223 (n38608, n_7077, n_28511);
  not g64224 (n_28652, n38606);
  and g64225 (n38609, pi0211, n_28652);
  and g64226 (n38610, pi0299, n_5);
  not g64227 (n_28653, n38610);
  and g64228 (n38611, n38540, n_28653);
  and g64229 (n38612, pi0299, pi1144);
  and g64230 (n38613, pi0207, n_28653);
  and g64231 (n38614, n_28614, n38613);
  not g64232 (n_28654, n38612);
  not g64233 (n_28655, n38614);
  and g64234 (n38615, n_28654, n_28655);
  not g64235 (n_28656, n38615);
  and g64236 (n38616, n38542, n_28656);
  and g64237 (n38617, n38574, n_28654);
  and g64238 (n38618, n38578, n_28654);
  and g64239 (n38619, n_11768, n38612);
  and g64240 (n38620, n38582, n_28653);
  not g64241 (n_28657, n38619);
  and g64242 (n38621, n38586, n_28657);
  not g64243 (n_28658, n38620);
  and g64244 (n38622, n_28658, n38621);
  not g64245 (n_28659, n38618);
  and g64246 (n38623, n_11794, n_28659);
  not g64247 (n_28660, n38622);
  and g64248 (n38624, n_28660, n38623);
  and g64249 (n38625, n38593, n_28654);
  and g64250 (n38626, n_28641, n_28653);
  not g64251 (n_28661, n38626);
  and g64252 (n38627, n_11413, n_28661);
  not g64253 (n_28662, n38625);
  and g64254 (n38628, pi1156, n_28662);
  not g64255 (n_28663, n38627);
  and g64256 (n38629, n_28663, n38628);
  not g64257 (n_28664, n38624);
  not g64258 (n_28665, n38629);
  and g64259 (n38630, n_28664, n_28665);
  and g64260 (n38631, n_25873, n38630);
  not g64261 (n_28666, n38617);
  and g64262 (n38632, pi0208, n_28666);
  not g64263 (n_28667, n38631);
  and g64264 (n38633, n_28667, n38632);
  not g64265 (n_28668, n38611);
  not g64266 (n_28669, n38616);
  and g64267 (n38634, n_28668, n_28669);
  not g64268 (n_28670, n38633);
  and g64269 (n38635, n_28670, n38634);
  not g64270 (n_28671, n38635);
  and g64271 (n38636, n_7075, n_28671);
  not g64272 (n_28672, n38609);
  and g64273 (n38637, n38608, n_28672);
  not g64274 (n_28673, n38636);
  and g64275 (n38638, n_28673, n38637);
  not g64276 (n_28674, n38607);
  not g64277 (n_28675, n38638);
  and g64278 (n38639, n_28674, n_28675);
  not g64279 (n_28676, n38639);
  and g64280 (n38640, n_6791, n_28676);
  and g64281 (n38641, n_234, n38561);
  not g64282 (n_28677, n38584);
  and g64283 (n38642, n_28677, n38641);
  and g64284 (n38643, n_28603, n38642);
  and g64285 (n38644, pi0207, n38643);
  not g64286 (n_28678, n38644);
  and g64287 (n38645, n_26242, n_28678);
  and g64288 (n38646, n10810, n_28637);
  not g64289 (n_28679, n38578);
  and g64290 (n38647, n_28679, n38646);
  and g64291 (n38648, pi0200, n_11768);
  not g64292 (n_28680, n38648);
  and g64293 (n38649, n11384, n_28680);
  and g64294 (n38650, pi1156, n38649);
  not g64295 (n_28681, n38647);
  not g64296 (n_28682, n38650);
  and g64297 (n38651, n_28681, n_28682);
  and g64298 (n38652, n_25873, n38651);
  not g64299 (n_28683, n38574);
  not g64300 (n_28684, n38652);
  and g64301 (n38653, n_28683, n_28684);
  not g64302 (n_28685, n38653);
  and g64303 (n38654, pi0208, n_28685);
  not g64304 (n_28686, n38645);
  not g64305 (n_28687, n38654);
  and g64306 (n38655, n_28686, n_28687);
  not g64307 (n_28688, n38655);
  and g64308 (n38656, n_11810, n_28688);
  and g64309 (n38657, n_11794, n_28612);
  and g64310 (n38658, n38568, n38657);
  not g64311 (n_28689, n38658);
  and g64312 (n38659, n_28613, n_28689);
  not g64313 (n_28690, n38659);
  and g64314 (n38660, pi0207, n_28690);
  not g64315 (n_28691, n38660);
  and g64316 (n38661, n_26242, n_28691);
  not g64317 (n_28692, n38661);
  and g64318 (n38662, n_28687, n_28692);
  not g64319 (n_28693, n38662);
  and g64320 (n38663, pi1157, n_28693);
  not g64321 (n_28694, n38656);
  not g64322 (n_28695, n38663);
  and g64323 (n38664, n_28694, n_28695);
  and g64324 (n38665, n_6791, n_28511);
  not g64325 (n_28696, n38665);
  and g64326 (n38666, n_28512, n_28696);
  not g64327 (n_28697, n38664);
  and g64328 (n38667, n_28697, n38666);
  not g64329 (n_28698, n38539);
  and g64330 (n38668, n_11810, n_28698);
  not g64331 (n_28699, n38547);
  and g64332 (n38669, n_11794, n_28699);
  not g64333 (n_28700, n38529);
  and g64334 (n38670, n11373, n_28700);
  not g64335 (n_28701, n38670);
  and g64336 (n38671, pi1156, n_28701);
  not g64337 (n_28702, n38669);
  not g64338 (n_28703, n38671);
  and g64339 (n38672, n_28702, n_28703);
  and g64340 (n38673, pi0207, n38672);
  and g64341 (n38674, n_25873, n_234);
  not g64342 (n_28704, n38674);
  and g64343 (n38675, n_26242, n_28704);
  not g64344 (n_28705, n38673);
  and g64345 (n38676, n_28705, n38675);
  not g64346 (n_28706, n38676);
  and g64347 (n38677, pi1157, n_28706);
  not g64348 (n_28707, n38668);
  and g64349 (n38678, n_28554, n_28707);
  not g64350 (n_28708, n38677);
  and g64351 (n38679, n_28708, n38678);
  and g64352 (n38680, pi0299, pi1142);
  and g64353 (n38681, pi1153, n38585);
  and g64354 (n38682, pi1153, n_28608);
  and g64355 (n38683, n_11757, n_7047);
  not g64356 (n_28709, n38682);
  not g64357 (n_28710, n38683);
  and g64358 (n38684, n_28709, n_28710);
  not g64359 (n_28711, n38684);
  and g64360 (n38685, pi1155, n_28711);
  not g64361 (n_28712, n38681);
  not g64362 (n_28713, n38685);
  and g64363 (n38686, n_28712, n_28713);
  not g64364 (n_28714, n38686);
  and g64365 (n38687, n_11413, n_28714);
  and g64366 (n38688, n_28624, n38641);
  not g64367 (n_28715, n38688);
  and g64368 (n38689, n_28640, n_28715);
  not g64369 (n_28716, n38689);
  and g64370 (n38690, pi1154, n_28716);
  not g64371 (n_28717, n38687);
  not g64372 (n_28718, n38690);
  and g64373 (n38691, n_28717, n_28718);
  not g64374 (n_28719, n38691);
  and g64375 (n38692, n_234, n_28719);
  not g64376 (n_28720, n38680);
  and g64377 (n38693, pi0207, n_28720);
  not g64378 (n_28721, n38692);
  and g64379 (n38694, n_28721, n38693);
  and g64380 (n38695, n_28628, n_28720);
  and g64381 (n38696, n_11413, n_11794);
  not g64382 (n_28722, n38695);
  and g64383 (n38697, n_28722, n38696);
  and g64384 (n38698, pi1156, n_28641);
  and g64385 (n38699, pi0199, n_7045);
  not g64386 (n_28723, n38699);
  and g64387 (n38700, n_234, n_28723);
  not g64388 (n_28724, n38700);
  and g64389 (n38701, n_11768, n_28724);
  not g64390 (n_28725, n38582);
  not g64391 (n_28726, n38701);
  and g64392 (n38702, n_28725, n_28726);
  not g64393 (n_28727, n38702);
  and g64394 (n38703, pi1154, n_28727);
  not g64395 (n_28728, n38698);
  not g64396 (n_28729, n38703);
  and g64397 (n38704, n_28728, n_28729);
  not g64398 (n_28730, n38704);
  and g64399 (n38705, n_28554, n_28730);
  not g64400 (n_28731, n38697);
  and g64401 (n38706, n_25873, n_28731);
  not g64402 (n_28732, n38705);
  and g64403 (n38707, n_28732, n38706);
  not g64404 (n_28733, n38707);
  and g64405 (n38708, pi0208, n_28733);
  not g64406 (n_28734, n38694);
  and g64407 (n38709, n_28734, n38708);
  not g64408 (n_28735, n38666);
  and g64420 (n38716, pi0213, n_28560);
  not g64421 (n_28741, n38715);
  and g64422 (n38717, n_28741, n38716);
  and g64423 (n38718, pi0211, n_28697);
  and g64424 (n38719, n_26565, n_28697);
  not g64425 (n_28742, n38719);
  and g64426 (n38720, n_26538, n_28742);
  not g64427 (n_28743, n38510);
  and g64428 (n38721, n_25873, n_28743);
  not g64429 (n_28744, n38721);
  and g64430 (n38722, n_26242, n_28744);
  and g64431 (n38723, n_7385, n_28610);
  not g64432 (n_28745, n38723);
  and g64433 (n38724, pi1156, n_28745);
  and g64434 (n38725, n_11794, n_28608);
  and g64435 (n38726, n_28726, n38725);
  not g64436 (n_28746, n38724);
  not g64437 (n_28747, n38726);
  and g64438 (n38727, n_28746, n_28747);
  and g64439 (n38728, pi0207, n38727);
  and g64440 (n38729, pi1157, n38722);
  not g64441 (n_28748, n38728);
  and g64442 (n38730, n_28748, n38729);
  and g64443 (n38731, n_11768, n_7385);
  and g64444 (n38732, n_234, n38532);
  not g64445 (n_28749, n38731);
  and g64446 (n38733, n_28630, n_28749);
  not g64447 (n_28750, n38732);
  and g64448 (n38734, n_28750, n38733);
  and g64449 (n38735, n38722, n38734);
  and g64450 (n38736, pi0207, n38691);
  and g64451 (n38737, n38651, n38721);
  not g64452 (n_28751, n38737);
  and g64453 (n38738, pi0208, n_28751);
  not g64454 (n_28752, n38736);
  and g64455 (n38739, n_28752, n38738);
  not g64456 (n_28753, n38730);
  not g64457 (n_28754, n38735);
  and g64458 (n38740, n_28753, n_28754);
  not g64459 (n_28755, n38739);
  and g64460 (n38741, n_28755, n38740);
  and g64461 (n38742, n38499, n38741);
  not g64462 (n_28756, n38742);
  and g64463 (n38743, n38720, n_28756);
  and g64464 (n38744, n_7075, n_26565);
  and g64465 (n38745, pi0299, n_11413);
  not g64466 (n_28757, n38745);
  and g64467 (n38746, pi1157, n_28757);
  and g64468 (n38747, n38676, n38746);
  and g64469 (n38748, n38651, n_28729);
  not g64470 (n_28758, n38748);
  and g64471 (n38749, n_25873, n_28758);
  and g64472 (n38750, n_234, n38689);
  not g64473 (n_28759, n38750);
  and g64474 (n38751, pi1154, n_28759);
  not g64475 (n_28760, n38751);
  and g64476 (n38752, n_28627, n_28760);
  not g64477 (n_28761, n38752);
  and g64478 (n38753, pi0207, n_28761);
  not g64479 (n_28762, n38749);
  not g64480 (n_28763, n38753);
  and g64481 (n38754, n_28762, n_28763);
  not g64482 (n_28764, n38754);
  and g64483 (n38755, pi0208, n_28764);
  and g64484 (n38756, n_28588, n_28678);
  not g64485 (n_28765, n38756);
  and g64486 (n38757, n_26242, n_28765);
  and g64487 (n38758, n_11810, n38757);
  not g64488 (n_28766, n38747);
  not g64489 (n_28767, n38758);
  and g64490 (n38759, n_28766, n_28767);
  not g64491 (n_28768, n38755);
  and g64492 (n38760, n_28768, n38759);
  and g64493 (n38761, n38744, n38760);
  and g64494 (n38762, pi1153, n_28724);
  not g64495 (n_28769, n38762);
  and g64496 (n38763, n38565, n_28769);
  not g64497 (n_28770, n38763);
  and g64498 (n38764, pi0207, n_28770);
  and g64499 (n38765, pi0299, n_11768);
  not g64500 (n_28771, n38533);
  and g64501 (n38766, pi1155, n_28771);
  not g64502 (n_28772, n38765);
  not g64503 (n_28773, n38766);
  and g64504 (n38767, n_28772, n_28773);
  and g64505 (n38768, n38704, n38767);
  and g64506 (n38769, pi0299, n_11757);
  not g64507 (n_28774, n38769);
  and g64508 (n38770, n_25873, n_28774);
  not g64509 (n_28775, n38768);
  and g64510 (n38771, n_28775, n38770);
  not g64511 (n_28776, n38764);
  not g64512 (n_28777, n38771);
  and g64513 (n38772, n_28776, n_28777);
  not g64514 (n_28778, n38772);
  and g64515 (n38773, pi0208, n_28778);
  and g64516 (n38774, n_28707, n_28774);
  and g64517 (n38775, n_28708, n38774);
  not g64518 (n_28779, n38773);
  and g64519 (n38776, n38499, n_28779);
  not g64520 (n_28780, n38775);
  and g64521 (n38777, n_28780, n38776);
  not g64522 (n_28781, n38761);
  and g64523 (n38778, pi0212, n_28781);
  not g64524 (n_28782, n38777);
  and g64525 (n38779, n_28782, n38778);
  not g64526 (n_28783, n38743);
  not g64527 (n_28784, n38779);
  and g64528 (n38780, n_28783, n_28784);
  not g64529 (n_28785, n38718);
  not g64530 (n_28786, n38780);
  and g64531 (n38781, n_28785, n_28786);
  not g64532 (n_28787, n38781);
  and g64533 (n38782, pi0219, n_28787);
  not g64534 (n_28788, n10484);
  not g64535 (n_28789, n38744);
  and g64536 (n38783, n_28788, n_28789);
  not g64537 (n_28790, n38741);
  and g64538 (n38784, n_28790, n38783);
  not g64539 (n_28791, n38760);
  and g64540 (n38785, n10484, n_28791);
  and g64541 (n38786, n_28603, n38539);
  and g64542 (n38787, pi0299, pi1156);
  not g64543 (n_28792, n38787);
  and g64544 (n38788, n_28691, n_28792);
  not g64545 (n_28793, n38788);
  and g64546 (n38789, n38542, n_28793);
  not g64547 (n_28794, n38573);
  and g64548 (n38790, pi0207, n_28794);
  and g64549 (n38791, n_28681, n_28728);
  not g64550 (n_28795, n38791);
  and g64551 (n38792, n_25873, n_28795);
  and g64552 (n38793, pi0207, n38787);
  not g64553 (n_28796, n38792);
  not g64554 (n_28797, n38793);
  and g64555 (n38794, n_28796, n_28797);
  not g64556 (n_28798, n38790);
  and g64557 (n38795, n_28798, n38794);
  not g64558 (n_28799, n38795);
  and g64559 (n38796, pi0208, n_28799);
  not g64560 (n_28800, n38786);
  not g64561 (n_28801, n38789);
  and g64562 (n38797, n_28800, n_28801);
  not g64563 (n_28802, n38796);
  and g64564 (n38798, n_28802, n38797);
  not g64565 (n_28803, n38798);
  and g64566 (n38799, n38744, n_28803);
  not g64567 (n_28804, n38784);
  not g64568 (n_28805, n38799);
  and g64569 (n38800, n_28804, n_28805);
  not g64570 (n_28806, n38785);
  and g64571 (n38801, n_28806, n38800);
  not g64572 (n_28807, n38801);
  and g64573 (n38802, pi0212, n_28807);
  and g64574 (n38803, pi0211, n_28803);
  and g64575 (n38804, n_25873, n38768);
  and g64576 (n38805, n38441, n38763);
  not g64577 (n_28808, n38805);
  and g64578 (n38806, pi0208, n_28808);
  not g64579 (n_28809, n38804);
  and g64580 (n38807, n_28809, n38806);
  not g64581 (n_28810, n38807);
  and g64582 (n38808, n38677, n_28810);
  not g64583 (n_28811, n38808);
  and g64584 (n38809, n_7075, n_28811);
  and g64585 (n38810, n_28694, n38809);
  not g64586 (n_28812, n38803);
  and g64587 (n38811, pi0214, n_28812);
  not g64588 (n_28813, n38810);
  and g64589 (n38812, n_28813, n38811);
  not g64590 (n_28814, n38812);
  and g64591 (n38813, n38720, n_28814);
  not g64592 (n_28815, n38802);
  and g64593 (n38814, n_6791, n_28815);
  not g64594 (n_28816, n38813);
  and g64595 (n38815, n_28816, n38814);
  not g64596 (n_28817, n38815);
  and g64597 (n38816, n_4226, n_28817);
  not g64598 (n_28818, n38782);
  and g64599 (n38817, n_28818, n38816);
  not g64600 (n_28819, n38817);
  and g64601 (n38818, n38507, n_28819);
  not g64602 (n_28820, n38717);
  and g64603 (n38819, n_26372, n_28820);
  not g64604 (n_28821, n38818);
  and g64605 (n38820, n_28821, n38819);
  not g64606 (n_28822, n38526);
  not g64607 (n_28823, n38820);
  and g64608 (n38821, n_28822, n_28823);
  not g64609 (n_28824, n38821);
  and g64610 (n38822, pi0230, n_28824);
  or g64611 (po0390, n38412, n38822);
  and g64612 (n38824, n_6900, n38651);
  and g64613 (n38825, n_25873, n_26242);
  not g64614 (n_28825, n38825);
  and g64615 (n38826, n_6900, n_28825);
  and g64616 (n38827, n_7044, n38584);
  and g64617 (n38828, n_11413, n_28621);
  not g64618 (n_28826, n38827);
  and g64619 (n38829, n38550, n_28826);
  not g64620 (n_28827, n38828);
  and g64621 (n38830, n_28827, n38829);
  and g64622 (n38831, pi0207, n38830);
  not g64623 (n_28828, n38826);
  not g64624 (n_28829, n38831);
  and g64625 (n38832, n_28828, n_28829);
  not g64626 (n_28830, n38824);
  not g64627 (n_28831, n38832);
  and g64628 (n38833, n_28830, n_28831);
  and g64629 (n38834, n_28512, n38833);
  not g64630 (n_28832, n38834);
  and g64631 (n38835, pi0219, n_28832);
  and g64632 (n38836, n_25873, n38514);
  and g64633 (n38837, pi0207, n_28758);
  not g64634 (n_28833, n38836);
  not g64635 (n_28834, n38837);
  and g64636 (n38838, n_28833, n_28834);
  not g64637 (n_28835, n38838);
  and g64638 (n38839, n_26242, n_28835);
  and g64639 (n38840, n_11768, n10809);
  not g64640 (n_28836, n38840);
  and g64641 (n38841, n_28611, n_28836);
  not g64642 (n_28837, n38841);
  and g64643 (n38842, n_234, n_28837);
  not g64644 (n_28838, n38842);
  and g64645 (n38843, n_28827, n_28838);
  and g64646 (n38844, pi0207, n38843);
  not g64647 (n_28839, n38844);
  and g64648 (n38845, n_28762, n_28839);
  not g64649 (n_28840, n38845);
  and g64650 (n38846, pi0208, n_28840);
  not g64651 (n_28841, n38839);
  not g64652 (n_28842, n38846);
  and g64653 (n38847, n_28841, n_28842);
  not g64654 (n_28843, n38847);
  and g64655 (n38848, n_7075, n_28843);
  and g64656 (n38849, n_28511, n38848);
  not g64657 (n_28844, n38849);
  and g64658 (n38850, n38835, n_28844);
  not g64659 (n_28845, n38833);
  and g64660 (n38851, n_26565, n_28845);
  not g64661 (n_28846, n38851);
  and g64662 (n38852, n_26538, n_28846);
  and g64663 (n38853, pi0207, n_28795);
  not g64664 (n_28847, n38853);
  and g64665 (n38854, n_28792, n_28847);
  not g64666 (n_28848, n38854);
  and g64667 (n38855, n_26242, n_28848);
  and g64668 (n38856, n38794, n_28829);
  not g64669 (n_28849, n38856);
  and g64670 (n38857, pi0208, n_28849);
  not g64671 (n_28850, n38855);
  not g64672 (n_28851, n38857);
  and g64673 (n38858, n_28850, n_28851);
  not g64674 (n_28852, n38858);
  and g64675 (n38859, n_7075, n_28852);
  and g64676 (n38860, n_28743, n38651);
  not g64677 (n_28853, n38860);
  and g64678 (n38861, n38722, n_28853);
  and g64679 (n38862, pi0207, n_28743);
  not g64680 (n_28854, n38830);
  and g64681 (n38863, n_28854, n38862);
  not g64682 (n_28855, n38863);
  and g64683 (n38864, pi0208, n_28855);
  and g64684 (n38865, n_28751, n38864);
  not g64685 (n_28856, n38861);
  not g64686 (n_28857, n38865);
  and g64687 (n38866, n_28856, n_28857);
  not g64688 (n_28858, n38866);
  and g64689 (n38867, pi0211, n_28858);
  not g64690 (n_28859, n38859);
  not g64691 (n_28860, n38867);
  and g64692 (n38868, n_28859, n_28860);
  and g64693 (n38869, pi0214, n38868);
  not g64694 (n_28861, n38869);
  and g64695 (n38870, n38852, n_28861);
  and g64696 (n38871, pi0211, n_28843);
  and g64697 (n38872, n_7075, n_28858);
  not g64698 (n_28862, n38872);
  and g64699 (n38873, pi0214, n_28862);
  not g64700 (n_28863, n38871);
  and g64701 (n38874, n_28863, n38873);
  and g64702 (n38875, n_26565, n38868);
  not g64703 (n_28864, n38874);
  and g64704 (n38876, pi0212, n_28864);
  not g64705 (n_28865, n38875);
  and g64706 (n38877, n_28865, n38876);
  not g64707 (n_28866, n38870);
  and g64708 (n38878, n_6791, n_28866);
  not g64709 (n_28867, n38877);
  and g64710 (n38879, n_28867, n38878);
  not g64711 (n_28868, n38850);
  and g64712 (n38880, n35819, n_28868);
  not g64713 (n_28869, n38879);
  and g64714 (n38881, n_28869, n38880);
  and g64715 (n38882, pi0211, pi1153);
  not g64716 (n_28870, n38882);
  and g64717 (n38883, n_28577, n_28870);
  and g64718 (n38884, n_7077, n38883);
  not g64719 (n_28871, n38884);
  and g64720 (n38885, n38665, n_28871);
  and g64721 (n38886, n_28581, n38885);
  and g64722 (n38887, po1038, n38886);
  not g64723 (n_28873, pi1152);
  not g64724 (n_28874, n38887);
  and g64725 (n38888, n_28873, n_28874);
  and g64726 (n38889, pi0207, n38767);
  and g64727 (n38890, n38704, n38889);
  not g64728 (n_28875, n38890);
  and g64729 (n38891, n38675, n_28875);
  not g64730 (n_28876, n38843);
  and g64731 (n38892, n38441, n_28876);
  not g64732 (n_28877, n38892);
  and g64733 (n38893, pi0208, n_28877);
  and g64734 (n38894, n_28809, n38893);
  not g64735 (n_28878, n38891);
  not g64736 (n_28879, n38894);
  and g64737 (n38895, n_28878, n_28879);
  not g64738 (n_28880, n38895);
  and g64739 (n38896, n_28774, n_28880);
  and g64740 (n38897, pi0211, n38896);
  not g64741 (n_28881, n38848);
  not g64742 (n_28882, n38897);
  and g64743 (n38898, n_28881, n_28882);
  and g64744 (n38899, pi0214, n38898);
  not g64745 (n_28883, n38899);
  and g64746 (n38900, n38852, n_28883);
  not g64747 (n_28884, n38900);
  and g64748 (n38901, n_6791, n_28884);
  not g64749 (n_28885, n38898);
  and g64750 (n38902, n_26565, n_28885);
  not g64751 (n_28886, n38896);
  and g64752 (n38903, n_7075, n_28886);
  not g64753 (n_28887, n38903);
  and g64754 (n38904, pi0214, n_28887);
  and g64755 (n38905, pi0211, n_28845);
  not g64756 (n_28888, n38905);
  and g64757 (n38906, n38904, n_28888);
  not g64758 (n_28889, n38902);
  not g64759 (n_28890, n38906);
  and g64760 (n38907, n_28889, n_28890);
  not g64761 (n_28891, n38907);
  and g64762 (n38908, pi0212, n_28891);
  not g64763 (n_28892, n38908);
  and g64764 (n38909, n38901, n_28892);
  and g64765 (n38910, pi0219, n_28845);
  not g64766 (n_28893, n38910);
  and g64767 (n38911, n_4226, n_28893);
  not g64768 (n_28894, n38909);
  and g64769 (n38912, n_28894, n38911);
  not g64770 (n_28895, n38912);
  and g64771 (n38913, n38888, n_28895);
  and g64772 (n38914, pi1153, n_28789);
  not g64773 (n_28896, n38499);
  and g64774 (n38915, n_28580, n_28896);
  not g64775 (n_28897, n38914);
  not g64776 (n_28898, n38915);
  and g64777 (n38916, n_28897, n_28898);
  not g64778 (n_28899, n38916);
  and g64779 (n38917, pi0212, n_28899);
  not g64780 (n_28900, n38883);
  and g64781 (n38918, n38421, n_28900);
  not g64782 (n_28901, n38918);
  and g64783 (n38919, n_6791, n_28901);
  not g64784 (n_28902, n38917);
  and g64785 (n38920, n_28902, n38919);
  not g64786 (n_28903, n38920);
  and g64787 (n38921, n38416, n_28903);
  not g64788 (n_28904, n38921);
  and g64789 (n38922, pi1152, n_28904);
  and g64790 (n38923, n_28880, n38904);
  not g64791 (n_28905, n38923);
  and g64792 (n38924, n_28889, n_28905);
  not g64793 (n_28906, n38924);
  and g64794 (n38925, pi0212, n_28906);
  not g64795 (n_28907, n38925);
  and g64796 (n38926, n38901, n_28907);
  and g64797 (n38927, n38414, n_28880);
  not g64798 (n_28908, n38927);
  and g64799 (n38928, n38835, n_28908);
  not g64800 (n_28909, n38928);
  and g64801 (n38929, n_4226, n_28909);
  not g64802 (n_28910, n38926);
  and g64803 (n38930, n_28910, n38929);
  not g64804 (n_28911, n38930);
  and g64805 (n38931, n38922, n_28911);
  not g64806 (n_28912, n38913);
  and g64807 (n38932, n_26557, n_28912);
  not g64808 (n_28913, n38931);
  and g64809 (n38933, n_28913, n38932);
  not g64810 (n_28914, n38881);
  and g64811 (n38934, pi0209, n_28914);
  not g64812 (n_28915, n38933);
  and g64813 (n38935, n_28915, n38934);
  and g64814 (n38936, n_7044, pi1153);
  and g64815 (n38937, pi0200, n38936);
  and g64816 (n38938, n_234, n38937);
  not g64817 (n_28916, n38938);
  and g64818 (n38939, n_11413, n_28916);
  and g64819 (n38940, pi1154, n38545);
  not g64820 (n_28917, n38936);
  and g64821 (n38941, n_28917, n38940);
  not g64822 (n_28918, n38939);
  not g64823 (n_28919, n38941);
  and g64824 (n38942, n_28918, n_28919);
  not g64825 (n_28920, n38942);
  and g64826 (n38943, n38700, n_28920);
  not g64827 (n_28921, n38943);
  and g64828 (n38944, n38675, n_28921);
  and g64829 (n38945, n_7045, n_11757);
  not g64830 (n_28922, n38945);
  and g64831 (n38946, n_7044, n_28922);
  not g64832 (n_28923, n38946);
  and g64833 (n38947, n_234, n_28923);
  and g64834 (n38948, n_28723, n38947);
  and g64835 (n38949, pi0207, n38948);
  and g64836 (n38950, n_25873, n38943);
  not g64837 (n_28924, n38949);
  and g64838 (n38951, pi0208, n_28924);
  not g64839 (n_28925, n38950);
  and g64840 (n38952, n_28925, n38951);
  not g64841 (n_28926, n38944);
  not g64842 (n_28927, n38952);
  and g64843 (n38953, n_28926, n_28927);
  and g64844 (n38954, n_7075, n38953);
  and g64845 (n38955, n_234, n10809);
  not g64846 (n_28928, n38955);
  and g64847 (n38956, n_11757, n_28928);
  not g64848 (n_28929, n38956);
  and g64849 (n38957, n38559, n_28929);
  and g64850 (n38958, n_7044, n_11757);
  not g64851 (n_28930, n38958);
  and g64852 (n38959, n38641, n_28930);
  not g64853 (n_28931, n38957);
  not g64854 (n_28932, n38959);
  and g64855 (n38960, n_28931, n_28932);
  and g64856 (n38961, n_6900, n38960);
  and g64857 (n38962, n_11757, n10809);
  not g64858 (n_28933, n38962);
  and g64859 (n38963, n38550, n_28933);
  not g64860 (n_28934, n38963);
  and g64861 (n38964, n10487, n_28934);
  not g64862 (n_28935, n38964);
  and g64863 (n38965, n_28825, n_28935);
  not g64864 (n_28936, n38961);
  and g64865 (n38966, n_28936, n38965);
  not g64866 (n_28937, n38966);
  and g64867 (n38967, pi0211, n_28937);
  not g64868 (n_28938, n38954);
  not g64869 (n_28939, n38967);
  and g64870 (n38968, n_28938, n_28939);
  and g64871 (n38969, n_28511, n38968);
  and g64872 (n38970, pi0219, n_28511);
  and g64873 (n38971, pi0219, n_28937);
  not g64874 (n_28940, n38970);
  not g64875 (n_28941, n38971);
  and g64876 (n38972, n_28940, n_28941);
  not g64877 (n_28942, n38969);
  not g64878 (n_28943, n38972);
  and g64879 (n38973, n_28942, n_28943);
  not g64880 (n_28944, n38973);
  and g64881 (n38974, n_4226, n_28944);
  and g64882 (n38975, n_25873, n38512);
  not g64883 (n_28945, n38568);
  and g64884 (n38976, n_11757, n_28945);
  not g64885 (n_28946, n38976);
  and g64886 (n38977, n_28630, n_28946);
  and g64887 (n38978, pi1154, n_28639);
  and g64888 (n38979, n_28946, n38978);
  not g64889 (n_28947, n38977);
  not g64890 (n_28948, n38979);
  and g64891 (n38980, n_28947, n_28948);
  not g64892 (n_28949, n38980);
  and g64893 (n38981, pi0207, n_28949);
  not g64894 (n_28950, n38975);
  not g64895 (n_28951, n38981);
  and g64896 (n38982, n_28950, n_28951);
  not g64897 (n_28952, n38982);
  and g64898 (n38983, n_26242, n_28952);
  and g64899 (n38984, n_25873, n_28949);
  and g64900 (n38985, n_234, n38549);
  not g64901 (n_28953, n38985);
  and g64902 (n38986, pi0207, n_28953);
  and g64903 (n38987, n_28710, n38986);
  not g64904 (n_28954, n38984);
  not g64905 (n_28955, n38987);
  and g64906 (n38988, n_28954, n_28955);
  not g64907 (n_28956, n38988);
  and g64908 (n38989, pi0208, n_28956);
  not g64909 (n_28957, n38983);
  not g64910 (n_28958, n38989);
  and g64911 (n38990, n_28957, n_28958);
  not g64912 (n_28959, n38990);
  and g64913 (n38991, n_7075, n_28959);
  not g64914 (n_28960, n38953);
  and g64915 (n38992, pi0211, n_28960);
  not g64916 (n_28961, n38991);
  and g64917 (n38993, pi0214, n_28961);
  not g64918 (n_28962, n38992);
  and g64919 (n38994, n_28962, n38993);
  not g64920 (n_28963, n38960);
  and g64921 (n38995, pi0207, n_28963);
  not g64922 (n_28964, n38995);
  and g64923 (n38996, n_28588, n_28964);
  not g64924 (n_28965, n38996);
  and g64925 (n38997, n_26242, n_28965);
  not g64926 (n_28966, n38948);
  and g64927 (n38998, pi0207, n_28966);
  and g64928 (n38999, n_28757, n38998);
  and g64929 (n39000, pi1154, n_7047);
  not g64930 (n_28967, n39000);
  and g64931 (n39001, n_28931, n_28967);
  and g64932 (n39002, n_28932, n39001);
  not g64933 (n_28968, n39002);
  and g64934 (n39003, n_25873, n_28968);
  not g64935 (n_28969, n38999);
  not g64936 (n_28970, n39003);
  and g64937 (n39004, n_28969, n_28970);
  not g64938 (n_28971, n39004);
  and g64939 (n39005, pi0208, n_28971);
  not g64940 (n_28972, n38997);
  not g64941 (n_28973, n39005);
  and g64942 (n39006, n_28972, n_28973);
  not g64943 (n_28974, n39006);
  and g64944 (n39007, n_7075, n_28974);
  and g64945 (n39008, pi0211, n_28959);
  not g64946 (n_28975, n39007);
  not g64947 (n_28976, n39008);
  and g64948 (n39009, n_28975, n_28976);
  and g64949 (n39010, n_26565, n39009);
  not g64950 (n_28977, n38994);
  and g64951 (n39011, pi0212, n_28977);
  not g64952 (n_28978, n39010);
  and g64953 (n39012, n_28978, n39011);
  and g64954 (n39013, n_26565, n_28937);
  not g64955 (n_28979, n39013);
  and g64956 (n39014, n_26538, n_28979);
  and g64957 (n39015, pi0214, n39009);
  not g64958 (n_28980, n39015);
  and g64959 (n39016, n39014, n_28980);
  not g64960 (n_28981, n39012);
  and g64961 (n39017, n_6791, n_28981);
  not g64962 (n_28982, n39016);
  and g64963 (n39018, n_28982, n39017);
  not g64964 (n_28983, n39018);
  and g64965 (n39019, n38974, n_28983);
  not g64966 (n_28984, n39019);
  and g64967 (n39020, n38922, n_28984);
  and g64968 (n39021, pi0200, n_11757);
  not g64969 (n_28985, n39021);
  and g64970 (n39022, n11384, n_28985);
  not g64971 (n_28986, n39022);
  and g64972 (n39023, pi1154, n_28986);
  not g64973 (n_28987, n39023);
  and g64974 (n39024, n_28918, n_28987);
  and g64975 (n39025, n38826, n39024);
  and g64976 (n39026, pi0208, n38441);
  and g64977 (n39027, pi1153, n_7047);
  and g64978 (n39028, n39026, n39027);
  not g64979 (n_28988, n39025);
  not g64980 (n_28989, n39028);
  and g64981 (n39029, n_28988, n_28989);
  and g64982 (n39030, pi0219, n39029);
  not g64983 (n_28990, n39030);
  and g64984 (n39031, n_4226, n_28990);
  and g64985 (n39032, pi1153, n_11413);
  and g64986 (n39033, n_28771, n39032);
  not g64987 (n_28991, n39033);
  and g64988 (n39034, n_28948, n_28991);
  not g64989 (n_28992, n39034);
  and g64990 (n39035, pi0207, n_28992);
  not g64991 (n_28993, n39035);
  and g64992 (n39036, n_28950, n_28993);
  not g64993 (n_28994, n39036);
  and g64994 (n39037, n_26242, n_28994);
  and g64995 (n39038, n_25873, n_28992);
  and g64996 (n39039, pi0207, n_7047);
  and g64997 (n39040, pi1153, n39039);
  not g64998 (n_28995, n39038);
  not g64999 (n_28996, n39040);
  and g65000 (n39041, n_28995, n_28996);
  not g65001 (n_28997, n39041);
  and g65002 (n39042, pi0208, n_28997);
  not g65003 (n_28998, n39037);
  not g65004 (n_28999, n39042);
  and g65005 (n39043, n_28998, n_28999);
  and g65006 (n39044, n38527, n39043);
  and g65007 (n39045, pi1153, n_28639);
  not g65008 (n_29000, n39045);
  and g65009 (n39046, n_28710, n_29000);
  not g65010 (n_29001, n39046);
  and g65011 (n39047, pi1154, n_29001);
  not g65012 (n_29002, n39047);
  and g65013 (n39048, n_28916, n_29002);
  not g65014 (n_29003, n39048);
  and g65015 (n39049, pi0207, n_29003);
  not g65016 (n_29004, n39049);
  and g65017 (n39050, n_28833, n_29004);
  not g65018 (n_29005, n39050);
  and g65019 (n39051, n_26242, n_29005);
  and g65020 (n39052, n_234, n_11757);
  not g65021 (n_29006, n39052);
  and g65022 (n39053, n_7047, n_29006);
  and g65023 (n39054, n_28757, n39053);
  not g65024 (n_29007, n39054);
  and g65025 (n39055, pi0207, n_29007);
  and g65026 (n39056, n_25873, n39048);
  not g65027 (n_29008, n39055);
  and g65028 (n39057, pi0208, n_29008);
  not g65029 (n_29009, n39056);
  and g65030 (n39058, n_29009, n39057);
  not g65031 (n_29010, n39051);
  not g65032 (n_29011, n39058);
  and g65033 (n39059, n_29010, n_29011);
  and g65034 (n39060, n_7075, n39059);
  and g65035 (n39061, pi0211, n39043);
  not g65036 (n_29012, n39060);
  not g65037 (n_29013, n39061);
  and g65038 (n39062, n_29012, n_29013);
  not g65039 (n_29014, n39062);
  and g65040 (n39063, n38608, n_29014);
  not g65041 (n_29015, n39044);
  not g65042 (n_29016, n39063);
  and g65043 (n39064, n_29015, n_29016);
  not g65044 (n_29017, n39064);
  and g65045 (n39065, n_6791, n_29017);
  not g65046 (n_29018, n38608);
  and g65047 (n39066, n_28896, n_29018);
  and g65048 (n39067, n39029, n39066);
  not g65049 (n_29019, n39067);
  and g65050 (n39068, n39031, n_29019);
  not g65051 (n_29020, n39065);
  and g65052 (n39069, n_29020, n39068);
  not g65053 (n_29021, n39069);
  and g65054 (n39070, n38888, n_29021);
  not g65055 (n_29022, n39020);
  not g65056 (n_29023, n39070);
  and g65057 (n39071, n_29022, n_29023);
  and g65058 (n39072, n_26557, n39071);
  and g65059 (n39073, n_28873, n_4226);
  not g65060 (n_29024, n39029);
  and g65061 (n39074, n38413, n_29024);
  not g65062 (n_29025, n38937);
  and g65063 (n39075, n_234, n_29025);
  not g65064 (n_29026, n39075);
  and g65065 (n39076, n_11413, n_29026);
  and g65066 (n39077, n_28772, n39076);
  and g65067 (n39078, n_28749, n39047);
  not g65068 (n_29027, n39077);
  not g65069 (n_29028, n39078);
  and g65070 (n39079, n_29027, n_29028);
  and g65071 (n39080, pi0207, n39079);
  not g65072 (n_29029, n39080);
  and g65073 (n39081, n38722, n_29029);
  and g65074 (n39082, n_25873, n39079);
  and g65075 (n39083, n_28772, n39053);
  not g65076 (n_29030, n39083);
  and g65077 (n39084, pi0207, n_29030);
  not g65078 (n_29031, n39084);
  and g65079 (n39085, pi0208, n_29031);
  not g65080 (n_29032, n39082);
  and g65081 (n39086, n_29032, n39085);
  not g65082 (n_29033, n39081);
  not g65083 (n_29034, n39086);
  and g65084 (n39087, n_29033, n_29034);
  and g65085 (n39088, n_7075, n39087);
  and g65086 (n39089, pi0211, n39059);
  not g65087 (n_29035, n39088);
  and g65088 (n39090, n10843, n_29035);
  not g65089 (n_29036, n39089);
  and g65090 (n39091, n_29036, n39090);
  and g65091 (n39092, n_7075, n_28792);
  and g65092 (n39093, n39029, n39092);
  and g65093 (n39094, pi0211, n39087);
  not g65094 (n_29037, n39093);
  and g65095 (n39095, n_28519, n_29037);
  not g65096 (n_29038, n39094);
  and g65097 (n39096, n_29038, n39095);
  not g65098 (n_29039, n39091);
  not g65099 (n_29040, n39096);
  and g65100 (n39097, n_29039, n_29040);
  not g65101 (n_29041, n39097);
  and g65102 (n39098, n_6791, n_29041);
  and g65103 (n39099, pi0211, n39029);
  not g65104 (n_29042, n39099);
  and g65105 (n39100, n38970, n_29042);
  and g65106 (n39101, n_29012, n39100);
  not g65107 (n_29043, n39074);
  not g65108 (n_29044, n39101);
  and g65109 (n39102, n_29043, n_29044);
  not g65110 (n_29045, n39098);
  and g65111 (n39103, n_29045, n39102);
  not g65112 (n_29046, n39103);
  and g65113 (n39104, n39073, n_29046);
  and g65114 (n39105, n_28512, n38966);
  and g65115 (n39106, n_28511, n39007);
  not g65116 (n_29047, n39105);
  not g65117 (n_29048, n39106);
  and g65118 (n39107, n_29047, n_29048);
  not g65119 (n_29049, n39107);
  and g65120 (n39108, pi0219, n_29049);
  and g65121 (n39109, n_26538, n39013);
  and g65122 (n39110, pi0211, n_28974);
  and g65123 (n39111, n_7044, n_11413);
  and g65124 (n39112, n_7045, n39111);
  and g65125 (n39113, n38674, n39112);
  and g65126 (n39114, n38722, n_28921);
  not g65127 (n_29050, n39114);
  and g65128 (n39115, n_28927, n_29050);
  not g65129 (n_29051, n39113);
  and g65130 (n39116, n_28772, n_29051);
  not g65131 (n_29052, n39115);
  and g65132 (n39117, n_29052, n39116);
  and g65133 (n39118, n_7075, n39117);
  not g65134 (n_29053, n39118);
  and g65135 (n39119, n10843, n_29053);
  not g65136 (n_29054, n39110);
  and g65137 (n39120, n_29054, n39119);
  and g65138 (n39121, n_26242, n_28792);
  and g65139 (n39122, n_28964, n39121);
  and g65140 (n39123, pi0299, n_11794);
  not g65141 (n_29055, n39123);
  and g65142 (n39124, n38998, n_29055);
  and g65143 (n39125, n_28792, n38960);
  not g65144 (n_29056, n39125);
  and g65145 (n39126, n_25873, n_29056);
  not g65146 (n_29057, n39124);
  and g65147 (n39127, pi0208, n_29057);
  not g65148 (n_29058, n39126);
  and g65149 (n39128, n_29058, n39127);
  not g65150 (n_29059, n39122);
  and g65151 (n39129, n_7075, n_29059);
  not g65152 (n_29060, n39128);
  and g65153 (n39130, n_29060, n39129);
  and g65154 (n39131, pi0211, n39117);
  not g65155 (n_29061, n39130);
  and g65156 (n39132, n_28519, n_29061);
  not g65157 (n_29062, n39131);
  and g65158 (n39133, n_29062, n39132);
  not g65165 (n_29066, n39108);
  not g65166 (n_29067, n39136);
  and g65167 (n39137, n_29066, n_29067);
  and g65168 (n39138, pi1152, n_4226);
  not g65169 (n_29068, n39137);
  and g65170 (n39139, n_29068, n39138);
  not g65171 (n_29069, n39104);
  not g65172 (n_29070, n39139);
  and g65173 (n39140, n_29069, n_29070);
  not g65174 (n_29071, n39140);
  and g65175 (n39141, pi0213, n_29071);
  not g65176 (n_29072, n39141);
  and g65177 (n39142, n_26372, n_29072);
  not g65178 (n_29073, n39072);
  and g65179 (n39143, n_29073, n39142);
  not g65180 (n_29074, n38935);
  not g65181 (n_29075, n39143);
  and g65182 (n39144, n_29074, n_29075);
  and g65183 (n39145, pi0219, n_28577);
  not g65184 (n_29076, n38491);
  and g65185 (n39146, pi0212, n_29076);
  and g65186 (n39147, pi0214, n_28568);
  and g65187 (n39148, n_26538, n39147);
  not g65188 (n_29077, n39148);
  and g65189 (n39149, n_6791, n_29077);
  not g65190 (n_29078, n39146);
  and g65191 (n39150, n_29078, n39149);
  not g65192 (n_29079, n39145);
  not g65197 (n_29081, n39144);
  not g65198 (n_29082, n39153);
  and g65199 (n39154, n_29081, n_29082);
  not g65200 (n_29083, n39154);
  and g65201 (n39155, pi0230, n_29083);
  and g65202 (n39156, n_28510, pi0234);
  or g65203 (po0391, n39155, n39156);
  and g65204 (n39158, pi0219, n_28569);
  and g65205 (n39159, pi0219, n_29018);
  and g65206 (n39160, n_26538, n38481);
  and g65207 (n39161, n_26565, n_28564);
  not g65208 (n_29084, n39147);
  not g65209 (n_29085, n39161);
  and g65210 (n39162, n_29084, n_29085);
  not g65211 (n_29086, n39162);
  and g65212 (n39163, pi0212, n_29086);
  not g65213 (n_29087, n39163);
  and g65214 (n39164, n_6791, n_29087);
  not g65215 (n_29088, n39160);
  and g65216 (n39165, n_29088, n39164);
  not g65217 (n_29089, n39158);
  not g65218 (n_29090, n39159);
  and g65223 (n39169, pi0208, pi1157);
  and g65224 (n39170, n_28682, n_28773);
  not g65225 (n_29092, n39170);
  and g65226 (n39171, pi0207, n_29092);
  not g65227 (n_29093, n38727);
  and g65228 (n39172, n_25873, n_29093);
  not g65229 (n_29094, n39171);
  not g65230 (n_29095, n39172);
  and g65231 (n39173, n_29094, n_29095);
  not g65232 (n_29096, n39173);
  and g65233 (n39174, n39169, n_29096);
  and g65234 (n39175, n_25873, n38734);
  not g65235 (n_29097, n39175);
  and g65236 (n39176, n_29094, n_29097);
  not g65237 (n_29098, n39176);
  and g65238 (n39177, pi0208, n_29098);
  not g65239 (n_29099, n39177);
  and g65240 (n39178, n_28754, n_29099);
  not g65241 (n_29100, n39178);
  and g65242 (n39179, n_11810, n_29100);
  not g65243 (n_29101, n39174);
  and g65244 (n39180, n_28753, n_29101);
  not g65245 (n_29102, n39179);
  and g65246 (n39181, n_29102, n39180);
  not g65247 (n_29103, n39181);
  and g65248 (n39182, pi0211, n_29103);
  and g65249 (n39183, n_11794, n38577);
  not g65250 (n_29104, n39183);
  and g65251 (n39184, n_28728, n_29104);
  not g65252 (n_29105, n39184);
  and g65253 (n39185, pi0207, n_29105);
  and g65254 (n39186, n_28689, n_28703);
  not g65255 (n_29106, n39186);
  and g65256 (n39187, n_25873, n_29106);
  not g65257 (n_29107, n39185);
  not g65258 (n_29108, n39187);
  and g65259 (n39188, n_29107, n_29108);
  not g65260 (n_29109, n39188);
  and g65261 (n39189, n39169, n_29109);
  and g65262 (n39190, n_25873, n38536);
  not g65263 (n_29110, n39190);
  and g65264 (n39191, n_29107, n_29110);
  not g65265 (n_29111, n39191);
  and g65266 (n39192, pi0208, n_29111);
  not g65267 (n_29112, n39192);
  and g65268 (n39193, n_28800, n_29112);
  not g65269 (n_29113, n39193);
  and g65270 (n39194, n_11810, n_29113);
  not g65271 (n_29114, n39189);
  and g65272 (n39195, n_28801, n_29114);
  not g65273 (n_29115, n39194);
  and g65274 (n39196, n_29115, n39195);
  not g65275 (n_29116, n39196);
  and g65276 (n39197, n_7075, n_29116);
  not g65277 (n_29117, n39182);
  and g65278 (n39198, n10843, n_29117);
  not g65279 (n_29118, n39197);
  and g65280 (n39199, n_29118, n39198);
  and g65281 (n39200, n10487, n_28682);
  and g65282 (n39201, n_29104, n39200);
  not g65283 (n_29119, n38643);
  and g65284 (n39202, n_25873, n_29119);
  not g65285 (n_29120, n39201);
  not g65286 (n_29121, n39202);
  and g65287 (n39203, n_29120, n_29121);
  and g65288 (n39204, n_28686, n39203);
  not g65289 (n_29122, n39204);
  and g65290 (n39205, n_11810, n_29122);
  and g65291 (n39206, n_25873, n38659);
  not g65292 (n_29123, n39206);
  and g65293 (n39207, n_29120, n_29123);
  and g65294 (n39208, n_28692, n39207);
  not g65295 (n_29124, n39208);
  and g65296 (n39209, pi1157, n_29124);
  not g65297 (n_29125, n39205);
  not g65298 (n_29126, n39209);
  and g65299 (n39210, n_29125, n_29126);
  not g65300 (n_29127, n39210);
  and g65301 (n39211, n38413, n_29127);
  and g65302 (n39212, pi0211, n_29116);
  and g65303 (n39213, n_25873, n38672);
  not g65304 (n_29128, n39213);
  and g65305 (n39214, pi0208, n_29128);
  and g65306 (n39215, n_28728, n38889);
  not g65307 (n_29129, n39215);
  and g65308 (n39216, n39214, n_29129);
  not g65309 (n_29130, n39216);
  and g65310 (n39217, n_28706, n_29130);
  and g65311 (n39218, pi1157, n39217);
  and g65312 (n39219, n_7075, n_29125);
  not g65313 (n_29131, n39218);
  and g65314 (n39220, n_29131, n39219);
  not g65315 (n_29132, n39220);
  and g65316 (n39221, n38608, n_29132);
  not g65317 (n_29133, n39212);
  and g65318 (n39222, n_29133, n39221);
  not g65319 (n_29134, n39211);
  not g65320 (n_29135, n39222);
  and g65321 (n39223, n_29134, n_29135);
  not g65322 (n_29136, n39199);
  and g65323 (n39224, n_29136, n39223);
  not g65324 (n_29137, n39224);
  and g65325 (n39225, n_6791, n_29137);
  and g65326 (n39226, n_7075, n39181);
  and g65327 (n39227, pi0211, n_29127);
  not g65328 (n_29138, n39227);
  and g65329 (n39228, n_28519, n_29138);
  not g65330 (n_29139, n39226);
  and g65331 (n39229, n_29139, n39228);
  and g65332 (n39230, n38423, n39210);
  not g65333 (n_29140, n39230);
  and g65334 (n39231, pi0219, n_29140);
  not g65335 (n_29141, n39229);
  and g65336 (n39232, n_29141, n39231);
  not g65337 (n_29142, n39232);
  and g65338 (n39233, pi0209, n_29142);
  not g65339 (n_29143, n39225);
  and g65340 (n39234, n_29143, n39233);
  and g65341 (n39235, n_28719, n38722);
  and g65342 (n39236, n_25873, n38691);
  and g65343 (n39237, pi0208, n_29029);
  not g65344 (n_29144, n39236);
  and g65345 (n39238, n_29144, n39237);
  not g65346 (n_29145, n39235);
  not g65347 (n_29146, n39238);
  and g65348 (n39239, n_29145, n_29146);
  not g65349 (n_29147, n39239);
  and g65350 (n39240, pi0211, n_29147);
  not g65351 (n_29148, n39024);
  and g65352 (n39241, n10487, n_29148);
  and g65353 (n39242, n_28794, n_28825);
  not g65354 (n_29149, n39242);
  and g65355 (n39243, n_6900, n_29149);
  not g65356 (n_29150, n39241);
  not g65357 (n_29151, n39243);
  and g65358 (n39244, n_29150, n_29151);
  not g65359 (n_29152, n39244);
  and g65360 (n39245, n_28792, n_29152);
  not g65361 (n_29153, n39245);
  and g65362 (n39246, n_7075, n_29153);
  not g65363 (n_29154, n39240);
  and g65364 (n39247, n10843, n_29154);
  not g65365 (n_29155, n39246);
  and g65366 (n39248, n_29155, n39247);
  and g65367 (n39249, n38413, n_29152);
  and g65368 (n39250, n38675, n_28808);
  and g65369 (n39251, n38674, n38763);
  not g65370 (n_29156, n39076);
  and g65371 (n39252, n_29002, n_29156);
  and g65372 (n39253, pi0207, n39252);
  not g65373 (n_29157, n39251);
  and g65374 (n39254, pi0208, n_29157);
  not g65375 (n_29158, n39253);
  and g65376 (n39255, n_29158, n39254);
  not g65377 (n_29159, n39250);
  not g65378 (n_29160, n39255);
  and g65379 (n39256, n_29159, n_29160);
  not g65380 (n_29161, n39256);
  and g65381 (n39257, pi1157, n_29161);
  and g65382 (n39258, n_11810, n39244);
  not g65383 (n_29162, n39257);
  and g65384 (n39259, n_7075, n_29162);
  not g65385 (n_29163, n39258);
  and g65386 (n39260, n_29163, n39259);
  and g65387 (n39261, pi0211, n39245);
  not g65388 (n_29164, n39260);
  not g65389 (n_29165, n39261);
  and g65390 (n39262, n_29164, n_29165);
  not g65391 (n_29166, n39262);
  and g65392 (n39263, n38608, n_29166);
  not g65393 (n_29167, n39248);
  not g65394 (n_29168, n39249);
  and g65395 (n39264, n_29167, n_29168);
  not g65396 (n_29169, n39263);
  and g65397 (n39265, n_29169, n39264);
  not g65398 (n_29170, n39265);
  and g65399 (n39266, n_6791, n_29170);
  and g65400 (n39267, n_7075, n39239);
  and g65401 (n39268, pi0211, n_29152);
  not g65402 (n_29171, n39268);
  and g65403 (n39269, n_28519, n_29171);
  not g65404 (n_29172, n39267);
  and g65405 (n39270, n_29172, n39269);
  and g65406 (n39271, n38423, n39244);
  not g65407 (n_29173, n39271);
  and g65408 (n39272, pi0219, n_29173);
  not g65409 (n_29174, n39270);
  and g65410 (n39273, n_29174, n39272);
  not g65411 (n_29175, n39273);
  and g65412 (n39274, n_26372, n_29175);
  not g65413 (n_29176, n39266);
  and g65414 (n39275, n_29176, n39274);
  not g65415 (n_29177, n39234);
  not g65416 (n_29178, n39275);
  and g65417 (n39276, n_29177, n_29178);
  not g65418 (n_29179, n39276);
  and g65419 (n39277, n_4226, n_29179);
  not g65420 (n_29180, n39168);
  and g65421 (n39278, pi0213, n_29180);
  not g65422 (n_29181, n39277);
  and g65423 (n39279, n_29181, n39278);
  and g65424 (n39280, pi0219, n_28578);
  not g65425 (n_29182, n39280);
  and g65426 (n39281, po1038, n_29182);
  and g65427 (n39282, n_28571, n38608);
  and g65428 (n39283, n10843, n_28900);
  not g65429 (n_29183, n39282);
  and g65430 (n39284, n_6791, n_29183);
  not g65431 (n_29184, n39283);
  and g65432 (n39285, n_29184, n39284);
  and g65433 (n39286, n_29090, n39281);
  not g65434 (n_29185, n39285);
  and g65435 (n39287, n_29185, n39286);
  not g65436 (n_29186, n39217);
  and g65437 (n39288, pi1157, n_29186);
  and g65438 (n39289, pi0299, n_11810);
  not g65439 (n_29187, n39289);
  and g65440 (n39290, n_29115, n_29187);
  not g65441 (n_29188, n39288);
  and g65442 (n39291, n_29188, n39290);
  not g65443 (n_29189, n39291);
  and g65444 (n39292, n_28774, n_29189);
  not g65445 (n_29190, n39292);
  and g65446 (n39293, n_7075, n_29190);
  not g65447 (n_29191, n39293);
  and g65448 (n39294, n39228, n_29191);
  not g65449 (n_29192, n39294);
  and g65450 (n39295, n39231, n_29192);
  not g65451 (n_29193, n38767);
  and g65452 (n39296, n_28679, n_29193);
  not g65453 (n_29194, n39296);
  and g65454 (n39297, n_28682, n_29194);
  not g65455 (n_29195, n39297);
  and g65456 (n39298, pi0207, n_29195);
  and g65457 (n39299, pi1154, n_28604);
  not g65458 (n_29196, n38642);
  not g65459 (n_29197, n39299);
  and g65460 (n39300, n_29196, n_29197);
  and g65461 (n39301, n_25873, n_28750);
  not g65462 (n_29198, n39300);
  and g65463 (n39302, n_29198, n39301);
  not g65464 (n_29199, n39298);
  not g65465 (n_29200, n39302);
  and g65466 (n39303, n_29199, n_29200);
  not g65467 (n_29201, n39303);
  and g65468 (n39304, pi0208, n_29201);
  not g65469 (n_29202, n38757);
  not g65470 (n_29203, n39304);
  and g65471 (n39305, n_29202, n_29203);
  not g65472 (n_29204, n39305);
  and g65473 (n39306, n_11810, n_29204);
  and g65474 (n39307, n38746, n_29186);
  not g65475 (n_29205, n39306);
  not g65476 (n_29206, n39307);
  and g65477 (n39308, n_29205, n_29206);
  not g65478 (n_29207, n39308);
  and g65479 (n39309, n_7075, n_29207);
  and g65480 (n39310, pi0211, n39292);
  not g65481 (n_29208, n39309);
  and g65482 (n39311, n10843, n_29208);
  not g65483 (n_29209, n39310);
  and g65484 (n39312, n_29209, n39311);
  and g65485 (n39313, pi0211, n39308);
  not g65486 (n_29210, n39313);
  and g65487 (n39314, n_29139, n_29210);
  not g65488 (n_29211, n39314);
  and g65489 (n39315, n38608, n_29211);
  not g65490 (n_29212, n39315);
  and g65491 (n39316, n_29134, n_29212);
  not g65492 (n_29213, n39312);
  and g65493 (n39317, n_29213, n39316);
  not g65494 (n_29214, n39317);
  and g65495 (n39318, n_6791, n_29214);
  not g65496 (n_29215, n39295);
  not g65497 (n_29216, n39318);
  and g65498 (n39319, n_29215, n_29216);
  not g65499 (n_29217, n39319);
  and g65500 (n39320, pi0209, n_29217);
  and g65501 (n39321, n_28776, n_28950);
  not g65502 (n_29218, n39321);
  and g65503 (n39322, n_26242, n_29218);
  and g65504 (n39323, n_25873, n_28770);
  not g65505 (n_29219, n39323);
  and g65506 (n39324, n_28993, n_29219);
  not g65507 (n_29220, n39324);
  and g65508 (n39325, pi0208, n_29220);
  not g65509 (n_29221, n39322);
  not g65510 (n_29222, n39325);
  and g65511 (n39326, n_29221, n_29222);
  and g65512 (n39327, n_7075, n39326);
  not g65513 (n_29223, n39327);
  and g65514 (n39328, n39269, n_29223);
  not g65515 (n_29224, n39328);
  and g65516 (n39329, n39272, n_29224);
  and g65517 (n39330, n_28763, n_28833);
  not g65518 (n_29225, n39330);
  and g65519 (n39331, n_26242, n_29225);
  and g65520 (n39332, n_25873, n_28761);
  not g65521 (n_29226, n39332);
  and g65522 (n39333, n_29004, n_29226);
  not g65523 (n_29227, n39333);
  and g65524 (n39334, pi0208, n_29227);
  not g65525 (n_29228, n39331);
  not g65526 (n_29229, n39334);
  and g65527 (n39335, n_29228, n_29229);
  and g65528 (n39336, pi0211, n39335);
  not g65529 (n_29230, n39336);
  and g65530 (n39337, n_29172, n_29230);
  not g65531 (n_29231, n39337);
  and g65532 (n39338, n_28519, n_29231);
  not g65533 (n_29232, n39335);
  and g65534 (n39339, n_7075, n_29232);
  not g65535 (n_29233, n39326);
  and g65536 (n39340, pi0211, n_29233);
  not g65537 (n_29234, n39340);
  and g65538 (n39341, n10843, n_29234);
  not g65539 (n_29235, n39339);
  and g65540 (n39342, n_29235, n39341);
  not g65541 (n_29236, n39342);
  and g65542 (n39343, n_29168, n_29236);
  not g65543 (n_29237, n39338);
  and g65544 (n39344, n_29237, n39343);
  not g65545 (n_29238, n39344);
  and g65546 (n39345, n_6791, n_29238);
  not g65547 (n_29239, n39329);
  not g65548 (n_29240, n39345);
  and g65549 (n39346, n_29239, n_29240);
  not g65550 (n_29241, n39346);
  and g65551 (n39347, n_26372, n_29241);
  not g65552 (n_29242, n39347);
  and g65553 (n39348, n_4226, n_29242);
  not g65554 (n_29243, n39320);
  and g65555 (n39349, n_29243, n39348);
  not g65556 (n_29244, n39287);
  and g65557 (n39350, n_26557, n_29244);
  not g65558 (n_29245, n39349);
  and g65559 (n39351, n_29245, n39350);
  not g65560 (n_29246, n39279);
  not g65561 (n_29247, n39351);
  and g65562 (n39352, n_29246, n_29247);
  not g65563 (n_29248, n39352);
  and g65564 (n39353, pi0230, n_29248);
  and g65565 (n39354, n_28510, n_1106);
  not g65566 (n_29249, n39353);
  not g65567 (n_29250, n39354);
  and g65568 (po0392, n_29249, n_29250);
  and g65569 (n39356, n_164, n38198);
  not g65570 (n_29251, n39356);
  and g65571 (n39357, n38397, n_29251);
  not g65572 (n_29252, n39357);
  and g65573 (n39358, n_3037, n_29252);
  not g65574 (n_29253, n39358);
  and g65575 (n39359, n_171, n_29253);
  not g65576 (n_29254, n39359);
  and g65577 (n39360, n_3993, n_29254);
  not g65578 (n_29255, n39360);
  and g65579 (n39361, n_174, n_29255);
  not g65580 (n_29256, n39361);
  and g65581 (n39362, n13654, n_29256);
  not g65582 (n_29257, n39362);
  and g65583 (n39363, n_168, n_29257);
  not g65584 (n_29258, n39363);
  and g65585 (n39364, n6131, n_29258);
  not g65586 (n_29259, n39364);
  and g65587 (n39365, n_157, n_29259);
  not g65588 (n_29260, n39365);
  and g65589 (n39366, n_3223, n_29260);
  not g65590 (n_29261, n39366);
  and g65591 (n39367, n_158, n_29261);
  not g65592 (n_29262, n39367);
  and g65593 (po0393, n13662, n_29262);
  and g65594 (n39369, pi0211, pi1157);
  and g65595 (n39370, n_7075, pi1158);
  not g65596 (n_29263, n39369);
  not g65597 (n_29264, n39370);
  and g65598 (n39371, n_29263, n_29264);
  not g65599 (n_29265, n39371);
  and g65600 (n39372, n38421, n_29265);
  not g65601 (n_29266, n39372);
  and g65602 (n39373, n39164, n_29266);
  and g65603 (n39374, n_6791, po1038);
  and g65604 (n39375, n38421, n38483);
  and g65605 (n39376, po1038, n39375);
  not g65606 (n_29267, n39374);
  not g65607 (n_29268, n39376);
  and g65608 (n39377, n_29267, n_29268);
  and g65609 (n39378, pi0214, n38495);
  and g65610 (n39379, pi1155, n38744);
  not g65611 (n_29269, n39378);
  not g65612 (n_29270, n39379);
  and g65613 (n39380, n_29269, n_29270);
  not g65614 (n_29271, n39380);
  and g65615 (n39381, pi0212, n_29271);
  and g65616 (n39382, po1038, n39381);
  not g65617 (n_29272, n39382);
  and g65618 (n39383, n39377, n_29272);
  not g65619 (n_29273, n39373);
  not g65620 (n_29274, n39383);
  and g65621 (n39384, n_29273, n_29274);
  not g65622 (n_29275, n39384);
  and g65623 (n39385, n_26557, n_29275);
  and g65624 (n39386, n38508, n_29273);
  and g65625 (n39387, pi0199, pi1143);
  not g65626 (n_29276, n39387);
  and g65627 (n39388, n_7045, n_29276);
  and g65628 (n39389, n_28527, n39388);
  and g65629 (n39390, n_28530, n39026);
  not g65630 (n_29277, n39389);
  and g65631 (n39391, n_29277, n39390);
  and g65632 (n39392, pi0200, n_28527);
  and g65633 (n39393, n_7044, pi1145);
  not g65634 (n_29278, n39393);
  and g65635 (n39394, n39388, n_29278);
  not g65636 (n_29279, n39392);
  and g65637 (n39395, n38826, n_29279);
  not g65638 (n_29280, n39394);
  and g65639 (n39396, n_29280, n39395);
  not g65640 (n_29281, n39391);
  not g65641 (n_29282, n39396);
  and g65642 (n39397, n_29281, n_29282);
  not g65643 (n_29283, n39397);
  and g65644 (n39398, n_234, n_29283);
  and g65645 (n39399, n38421, n38787);
  and g65646 (n39400, pi0214, n_28588);
  and g65647 (n39401, n_26565, n_28743);
  not g65648 (n_29284, n39400);
  and g65649 (n39402, pi0212, n_29284);
  not g65650 (n_29285, n39401);
  and g65651 (n39403, n_29285, n39402);
  not g65652 (n_29286, n39399);
  not g65653 (n_29287, n39403);
  and g65654 (n39404, n_29286, n_29287);
  not g65655 (n_29288, n39404);
  and g65656 (n39405, n38519, n_29288);
  not g65657 (n_29289, n39398);
  not g65658 (n_29290, n39405);
  and g65659 (n39406, n_29289, n_29290);
  not g65660 (n_29291, n39386);
  and g65661 (n39407, n_29291, n39406);
  not g65662 (n_29292, n39407);
  and g65663 (n39408, n_4226, n_29292);
  not g65664 (n_29293, n39408);
  and g65665 (n39409, n39385, n_29293);
  and g65666 (n39410, pi0219, n_28544);
  and g65667 (n39411, n10843, n38420);
  and g65668 (n39412, n_7075, pi1145);
  and g65669 (n39413, pi0211, pi1144);
  not g65670 (n_29294, n39412);
  not g65671 (n_29295, n39413);
  and g65672 (n39414, n_29294, n_29295);
  and g65673 (n39415, n_7077, n39414);
  not g65674 (n_29296, n39411);
  and g65675 (n39416, n_28511, n_29296);
  not g65676 (n_29297, n39415);
  and g65677 (n39417, n_29297, n39416);
  not g65678 (n_29298, n39417);
  and g65679 (n39418, n_6791, n_29298);
  not g65680 (n_29299, n39410);
  and g65681 (n39419, n38416, n_29299);
  not g65682 (n_29300, n39418);
  and g65683 (n39420, n_29300, n39419);
  and g65684 (n39421, n38508, n39417);
  and g65685 (n39422, pi0299, n38970);
  and g65686 (n39423, n38425, n39422);
  not g65687 (n_29301, n39423);
  and g65688 (n39424, n_29289, n_29301);
  not g65689 (n_29302, n39421);
  and g65690 (n39425, n_29302, n39424);
  not g65691 (n_29303, n39425);
  and g65692 (n39426, n_4226, n_29303);
  not g65693 (n_29304, n39420);
  not g65694 (n_29305, n39426);
  and g65695 (n39427, n_29304, n_29305);
  and g65696 (n39428, pi0213, n39427);
  not g65697 (n_29306, n39409);
  and g65698 (n39429, pi0209, n_29306);
  not g65699 (n_29307, n39428);
  and g65700 (n39430, n_29307, n39429);
  and g65701 (n39431, n38449, n38568);
  and g65702 (n39432, pi1158, n38955);
  and g65703 (n39433, n_7044, n_11397);
  not g65704 (n_29308, n39433);
  and g65705 (n39434, pi1156, n_29308);
  not g65706 (n_29309, n39432);
  not g65707 (n_29310, n39434);
  and g65708 (n39435, n_29309, n_29310);
  not g65709 (n_29311, n39435);
  and g65710 (n39436, n39431, n_29311);
  and g65711 (n39437, pi0207, n38651);
  and g65712 (n39438, pi0208, n_29121);
  not g65713 (n_29312, n39437);
  and g65714 (n39439, n_29312, n39438);
  not g65715 (n_29313, n39436);
  not g65716 (n_29314, n39439);
  and g65717 (n39440, n_29313, n_29314);
  not g65718 (n_29315, n39440);
  and g65719 (n39441, n_11810, n_29315);
  and g65720 (n39442, pi1156, n38699);
  and g65721 (n39443, n_7045, n_11397);
  not g65722 (n_29316, n39443);
  and g65723 (n39444, n_7044, n_29316);
  not g65724 (n_29317, n39442);
  not g65725 (n_29318, n39444);
  and g65726 (n39445, n_29317, n_29318);
  not g65727 (n_29319, n39445);
  and g65728 (n39446, n38441, n_29319);
  and g65729 (n39447, n_26242, n39446);
  and g65730 (n39448, pi0208, n_29123);
  and g65731 (n39449, n_29312, n39448);
  not g65732 (n_29320, n39447);
  not g65733 (n_29321, n39449);
  and g65734 (n39450, n_29320, n_29321);
  not g65735 (n_29322, n39450);
  and g65736 (n39451, pi1157, n_29322);
  not g65737 (n_29323, n39441);
  not g65738 (n_29324, n39451);
  and g65739 (n39452, n_29323, n_29324);
  and g65740 (n39453, n_28512, n39452);
  and g65741 (n39454, n_7045, pi0207);
  and g65742 (n39455, n_29311, n39454);
  not g65743 (n_29325, n39455);
  and g65744 (n39456, n_11810, n_29325);
  and g65745 (n39457, pi1156, n_28953);
  not g65746 (n_29326, n38641);
  and g65747 (n39458, n_11397, n_29326);
  not g65748 (n_29327, n39458);
  and g65749 (n39459, n39457, n_29327);
  not g65750 (n_29328, n39459);
  and g65751 (n39460, n_29318, n_29328);
  not g65752 (n_29329, n39460);
  and g65753 (n39461, n38441, n_29329);
  not g65754 (n_29330, n39456);
  and g65755 (n39462, n_26242, n_29330);
  and g65756 (n39463, n39461, n39462);
  not g65757 (n_29331, n39463);
  and g65758 (n39464, n_26242, n_29331);
  and g65759 (n39465, n_28615, n39464);
  not g65760 (n_29332, n38536);
  and g65761 (n39466, n_234, n_29332);
  and g65762 (n39467, n_7045, pi1157);
  and g65763 (n39468, n_7044, n39467);
  not g65764 (n_29333, n39468);
  and g65765 (n39469, n39466, n_29333);
  and g65766 (n39470, n_25873, n_28607);
  not g65767 (n_29334, n39469);
  and g65768 (n39471, n_29334, n39470);
  not g65769 (n_29335, n38601);
  and g65770 (n39472, pi0207, n_29335);
  not g65771 (n_29336, n39471);
  and g65772 (n39473, pi0208, n_29336);
  not g65773 (n_29337, n39472);
  and g65774 (n39474, n_29337, n39473);
  not g65775 (n_29338, n39465);
  not g65776 (n_29339, n39474);
  and g65777 (n39475, n_29338, n_29339);
  not g65778 (n_29340, n39475);
  and g65779 (n39476, n38414, n_29340);
  not g65780 (n_29341, n39453);
  not g65781 (n_29342, n39476);
  and g65782 (n39477, n_29341, n_29342);
  not g65783 (n_29343, n39477);
  and g65784 (n39478, pi0219, n_29343);
  and g65785 (n39479, n_26565, n39452);
  not g65786 (n_29344, n39479);
  and g65787 (n39480, n_26538, n_29344);
  and g65788 (n39481, pi0299, n_986);
  not g65789 (n_29345, n39481);
  and g65790 (n39482, n_25873, n_29345);
  and g65791 (n39483, n_29334, n39482);
  and g65792 (n39484, pi0299, pi1145);
  not g65793 (n_29346, n39484);
  and g65794 (n39485, n38578, n_29346);
  and g65795 (n39486, n_28727, n_29345);
  not g65796 (n_29347, n39486);
  and g65797 (n39487, pi1154, n_29347);
  not g65798 (n_29348, n39485);
  and g65799 (n39488, n_11794, n_29348);
  not g65800 (n_29349, n39487);
  and g65801 (n39489, n_29349, n39488);
  and g65802 (n39490, n38593, n_29346);
  and g65803 (n39491, n_28641, n_29345);
  not g65804 (n_29350, n39491);
  and g65805 (n39492, n_11413, n_29350);
  not g65806 (n_29351, n39490);
  and g65807 (n39493, pi1156, n_29351);
  not g65808 (n_29352, n39492);
  and g65809 (n39494, n_29352, n39493);
  not g65810 (n_29353, n39489);
  not g65811 (n_29354, n39494);
  and g65812 (n39495, n_29353, n_29354);
  not g65813 (n_29355, n39495);
  and g65814 (n39496, pi0207, n_29355);
  not g65815 (n_29356, n39483);
  and g65816 (n39497, pi0208, n_29356);
  not g65817 (n_29357, n39496);
  and g65818 (n39498, n_29357, n39497);
  not g65819 (n_29358, n38725);
  and g65820 (n39499, n38641, n_29358);
  and g65821 (n39500, pi1157, n_29309);
  not g65822 (n_29359, n39499);
  and g65823 (n39501, n_29359, n39500);
  not g65824 (n_29360, n39501);
  and g65825 (n39502, pi0207, n_29360);
  and g65826 (n39503, n_234, n39442);
  and g65827 (n39504, n_11810, n_29309);
  not g65828 (n_29361, n39503);
  and g65829 (n39505, n_29361, n39504);
  not g65830 (n_29362, n39505);
  and g65831 (n39506, n39502, n_29362);
  and g65832 (n39507, n_26242, n_29346);
  not g65833 (n_29363, n39506);
  and g65834 (n39508, n_29363, n39507);
  not g65835 (n_29364, n39498);
  not g65836 (n_29365, n39508);
  and g65837 (n39509, n_29364, n_29365);
  not g65838 (n_29366, n39509);
  and g65839 (n39510, n_7075, n_29366);
  and g65840 (n39511, n_28654, n39464);
  and g65841 (n39512, n_25873, n_28653);
  and g65842 (n39513, n_29334, n39512);
  not g65843 (n_29367, n38630);
  and g65844 (n39514, pi0207, n_29367);
  not g65845 (n_29368, n39513);
  and g65846 (n39515, pi0208, n_29368);
  not g65847 (n_29369, n39514);
  and g65848 (n39516, n_29369, n39515);
  not g65849 (n_29370, n39511);
  not g65850 (n_29371, n39516);
  and g65851 (n39517, n_29370, n_29371);
  not g65852 (n_29372, n39517);
  and g65853 (n39518, pi0211, n_29372);
  not g65854 (n_29373, n39510);
  not g65855 (n_29374, n39518);
  and g65856 (n39519, n_29373, n_29374);
  not g65857 (n_29375, n39519);
  and g65858 (n39520, pi0214, n_29375);
  not g65859 (n_29376, n39520);
  and g65860 (n39521, n39480, n_29376);
  and g65861 (n39522, n_7075, n39517);
  and g65862 (n39523, pi0211, n39475);
  not g65863 (n_29377, n39522);
  and g65864 (n39524, pi0214, n_29377);
  not g65865 (n_29378, n39523);
  and g65866 (n39525, n_29378, n39524);
  and g65867 (n39526, n_26565, n_29375);
  not g65868 (n_29379, n39525);
  and g65869 (n39527, pi0212, n_29379);
  not g65870 (n_29380, n39526);
  and g65871 (n39528, n_29380, n39527);
  not g65872 (n_29381, n39521);
  and g65873 (n39529, n_6791, n_29381);
  not g65874 (n_29382, n39528);
  and g65875 (n39530, n_29382, n39529);
  not g65876 (n_29383, n39478);
  and g65877 (n39531, n_4226, n_29383);
  not g65878 (n_29384, n39530);
  and g65879 (n39532, n_29384, n39531);
  and g65880 (n39533, pi0213, n_29304);
  not g65881 (n_29385, n39532);
  and g65882 (n39534, n_29385, n39533);
  and g65883 (n39535, n_28847, n_29108);
  not g65884 (n_29386, n39535);
  and g65885 (n39536, n39169, n_29386);
  not g65886 (n_29387, n39446);
  and g65887 (n39537, n_28792, n_29387);
  not g65888 (n_29388, n39537);
  and g65889 (n39538, n38542, n_29388);
  and g65890 (n39539, n39121, n_29325);
  and g65891 (n39540, pi0208, n_29110);
  and g65892 (n39541, n_28847, n39540);
  not g65893 (n_29389, n39539);
  and g65894 (n39542, n_11810, n_29389);
  not g65895 (n_29390, n39541);
  and g65896 (n39543, n_29390, n39542);
  not g65897 (n_29391, n39536);
  not g65898 (n_29392, n39538);
  and g65899 (n39544, n_29391, n_29392);
  not g65900 (n_29393, n39543);
  and g65901 (n39545, n_29393, n39544);
  and g65902 (n39546, n38421, n39545);
  and g65903 (n39547, pi0207, n_28853);
  not g65904 (n_29394, n39547);
  and g65905 (n39548, n_29095, n_29394);
  not g65906 (n_29395, n39548);
  and g65907 (n39549, n39169, n_29395);
  not g65908 (n_29396, n39461);
  and g65909 (n39550, n_28743, n_29396);
  not g65910 (n_29397, n39550);
  and g65911 (n39551, n38542, n_29397);
  and g65912 (n39552, n_29097, n_29394);
  not g65913 (n_29398, n39552);
  and g65914 (n39553, pi0208, n_29398);
  and g65915 (n39554, n_26242, n38510);
  not g65916 (n_29399, n39554);
  and g65917 (n39555, n_29313, n_29399);
  not g65918 (n_29400, n39553);
  and g65919 (n39556, n_29400, n39555);
  not g65920 (n_29401, n39556);
  and g65921 (n39557, n_11810, n_29401);
  not g65922 (n_29402, n39549);
  not g65923 (n_29403, n39551);
  and g65924 (n39558, n_29402, n_29403);
  not g65925 (n_29404, n39557);
  and g65926 (n39559, n_29404, n39558);
  not g65927 (n_29405, n39559);
  and g65928 (n39560, n_26565, n_29405);
  not g65929 (n_29406, n38672);
  and g65930 (n39561, n_25873, n_29406);
  and g65931 (n39562, n_28757, n39561);
  not g65932 (n_29407, n39562);
  and g65933 (n39563, pi1157, n_29407);
  and g65934 (n39564, n_11810, n_29313);
  and g65935 (n39565, n_29200, n39564);
  not g65936 (n_29408, n39563);
  not g65937 (n_29409, n39565);
  and g65938 (n39566, n_29408, n_29409);
  and g65939 (n39567, pi0208, n_28834);
  not g65940 (n_29410, n39566);
  and g65941 (n39568, n_29410, n39567);
  not g65942 (n_29411, n39564);
  and g65943 (n39569, n39461, n_29411);
  and g65944 (n39570, n_26242, n_28588);
  not g65945 (n_29412, n39569);
  and g65946 (n39571, n_29412, n39570);
  not g65947 (n_29413, n39571);
  and g65948 (n39572, pi0214, n_29413);
  not g65949 (n_29414, n39568);
  and g65950 (n39573, n_29414, n39572);
  not g65951 (n_29415, n39573);
  and g65952 (n39574, pi0212, n_29415);
  not g65953 (n_29416, n39560);
  and g65954 (n39575, n_29416, n39574);
  not g65955 (n_29417, n39546);
  not g65956 (n_29418, n39575);
  and g65957 (n39576, n_29417, n_29418);
  not g65958 (n_29419, n39576);
  and g65959 (n39577, n_7075, n_29419);
  not g65960 (n_29420, n39577);
  and g65961 (n39578, n_29341, n_29420);
  not g65962 (n_29421, n39578);
  and g65963 (n39579, pi0219, n_29421);
  and g65964 (n39580, n_234, n39445);
  not g65965 (n_29422, n39580);
  and g65966 (n39581, n38675, n_29422);
  and g65967 (n39582, n_28875, n39214);
  not g65968 (n_29423, n39581);
  not g65969 (n_29424, n39582);
  and g65970 (n39583, n_29423, n_29424);
  not g65971 (n_29425, n39583);
  and g65972 (n39584, pi1157, n_29425);
  not g65973 (n_29426, n39584);
  and g65974 (n39585, n_29323, n_29426);
  and g65975 (n39586, pi0211, n39585);
  and g65976 (n39587, n38441, n39442);
  not g65977 (n_29427, n39039);
  and g65978 (n39588, n_234, n_29427);
  not g65979 (n_29428, n39588);
  and g65980 (n39589, pi1158, n_29428);
  not g65981 (n_29429, n39587);
  and g65982 (n39590, n_26242, n_29429);
  not g65983 (n_29430, n39589);
  and g65984 (n39591, n_29430, n39590);
  and g65985 (n39592, n_11397, n38651);
  and g65986 (n39593, pi1158, n38768);
  not g65987 (n_29431, n39592);
  and g65988 (n39594, pi0207, n_29431);
  not g65989 (n_29432, n39593);
  and g65990 (n39595, n_29432, n39594);
  and g65991 (n39596, pi0299, n_11397);
  not g65992 (n_29433, n39596);
  and g65993 (n39597, n_25873, n_29433);
  not g65994 (n_29434, n39466);
  and g65995 (n39598, n_29434, n39597);
  not g65996 (n_29435, n39598);
  and g65997 (n39599, pi0208, n_29435);
  not g65998 (n_29436, n39595);
  and g65999 (n39600, n_29436, n39599);
  not g66000 (n_29437, n39591);
  and g66001 (n39601, n_11810, n_29437);
  not g66002 (n_29438, n39600);
  and g66003 (n39602, n_29438, n39601);
  and g66004 (n39603, n39561, n_29433);
  not g66005 (n_29439, n39603);
  and g66006 (n39604, n_29436, n_29439);
  not g66007 (n_29440, n39604);
  and g66008 (n39605, n39169, n_29440);
  not g66009 (n_29441, n39502);
  and g66010 (n39606, n_29441, n_29430);
  not g66011 (n_29442, n39606);
  and g66012 (n39607, n38542, n_29442);
  not g66013 (n_29443, n39607);
  and g66014 (n39608, n_7075, n_29443);
  not g66015 (n_29444, n39602);
  and g66016 (n39609, n_29444, n39608);
  not g66017 (n_29445, n39605);
  and g66018 (n39610, n_29445, n39609);
  not g66019 (n_29446, n39586);
  not g66020 (n_29447, n39610);
  and g66021 (n39611, n_29446, n_29447);
  not g66022 (n_29448, n39611);
  and g66023 (n39612, pi0214, n_29448);
  not g66024 (n_29449, n39612);
  and g66025 (n39613, n39480, n_29449);
  not g66026 (n_29450, n39545);
  and g66027 (n39614, n38783, n_29450);
  and g66028 (n39615, n10484, n_29405);
  not g66029 (n_29451, n39585);
  and g66030 (n39616, n38744, n_29451);
  not g66031 (n_29452, n39614);
  not g66032 (n_29453, n39615);
  and g66033 (n39617, n_29452, n_29453);
  not g66034 (n_29454, n39616);
  and g66035 (n39618, n_29454, n39617);
  not g66036 (n_29455, n39618);
  and g66037 (n39619, pi0212, n_29455);
  not g66038 (n_29456, n39619);
  and g66039 (n39620, n_6791, n_29456);
  not g66040 (n_29457, n39613);
  and g66041 (n39621, n_29457, n39620);
  not g66042 (n_29458, n39579);
  and g66043 (n39622, n_4226, n_29458);
  not g66044 (n_29459, n39621);
  and g66045 (n39623, n_29459, n39622);
  not g66046 (n_29460, n39623);
  and g66047 (n39624, n39385, n_29460);
  not g66048 (n_29461, n39534);
  and g66049 (n39625, n_26372, n_29461);
  not g66050 (n_29462, n39624);
  and g66051 (n39626, n_29462, n39625);
  not g66052 (n_29463, n39430);
  not g66053 (n_29464, n39626);
  and g66054 (n39627, n_29463, n_29464);
  not g66055 (n_29465, n39627);
  and g66056 (n39628, pi0230, n_29465);
  and g66057 (n39629, n_28510, n_25730);
  or g66058 (po0394, n39628, n39629);
  and g66059 (n39631, n_7075, n_11757);
  and g66060 (n39632, pi0219, n39631);
  not g66061 (n_29466, n39632);
  and g66062 (n39633, n38416, n_29466);
  and g66063 (n39634, n_29185, n39633);
  not g66064 (n_29468, pi1151);
  and g66065 (n39635, n_29468, n_4226);
  and g66066 (n39636, n10809, n38826);
  not g66067 (n_29469, n39636);
  and g66068 (n39637, n_234, n_29469);
  not g66069 (n_29470, n39637);
  and g66070 (n39638, n_8688, n_29470);
  and g66071 (n39639, n38826, n38955);
  not g66072 (n_29471, n39639);
  and g66073 (n39640, n_26565, n_29471);
  and g66074 (n39641, n_26538, n39640);
  not g66075 (n_29472, n39641);
  and g66076 (n39642, n39638, n_29472);
  and g66077 (n39643, pi1153, n39642);
  not g66078 (n_29473, n39643);
  and g66079 (n39644, n_28696, n_29473);
  and g66080 (n39645, n38882, n_29470);
  and g66081 (n39646, pi1153, n39639);
  not g66082 (n_29474, n39646);
  and g66083 (n39647, n_28588, n_29474);
  not g66084 (n_29475, n39647);
  and g66085 (n39648, n_7075, n_29475);
  not g66086 (n_29476, n39645);
  and g66087 (n39649, n10843, n_29476);
  not g66088 (n_29477, n39648);
  and g66089 (n39650, n_29477, n39649);
  and g66090 (n39651, pi0299, n_28571);
  not g66091 (n_29478, n39651);
  and g66092 (n39652, n_28519, n_29478);
  and g66093 (n39653, n_29474, n39652);
  not g66094 (n_29479, n39650);
  not g66095 (n_29480, n39653);
  and g66096 (n39654, n_29479, n_29480);
  not g66097 (n_29481, n39654);
  and g66098 (n39655, n_6791, n_29481);
  not g66099 (n_29482, n39644);
  and g66100 (n39656, n39635, n_29482);
  not g66101 (n_29483, n39655);
  and g66102 (n39657, n_29483, n39656);
  and g66103 (n39658, n_6900, n38568);
  and g66104 (n39659, n_28825, n39658);
  and g66105 (n39660, n38561, n39026);
  not g66106 (n_29484, n39659);
  not g66107 (n_29485, n39660);
  and g66108 (n39661, n_29484, n_29485);
  not g66109 (n_29486, n39661);
  and g66110 (n39662, n_28933, n_29486);
  not g66111 (n_29487, n39662);
  and g66112 (n39663, n_26565, n_29487);
  not g66113 (n_29488, n39663);
  and g66114 (n39664, n_26538, n_29488);
  and g66115 (n39665, n38568, n_28930);
  and g66116 (n39666, n_11757, n_28724);
  not g66117 (n_29489, n39666);
  and g66118 (n39667, n_28709, n_29489);
  not g66119 (n_29490, n39667);
  and g66120 (n39668, pi1155, n_29490);
  not g66121 (n_29491, n39665);
  not g66122 (n_29492, n39668);
  and g66123 (n39669, n_29491, n_29492);
  and g66124 (n39670, n38441, n_28629);
  not g66125 (n_29493, n39670);
  and g66126 (n39671, pi0208, n_29493);
  not g66127 (n_29494, n38722);
  not g66128 (n_29495, n39671);
  and g66129 (n39672, n_29494, n_29495);
  not g66130 (n_29496, n39669);
  not g66131 (n_29497, n39672);
  and g66132 (n39673, n_29496, n_29497);
  not g66133 (n_29498, n39673);
  and g66134 (n39674, n_29485, n_29498);
  not g66135 (n_29499, n39674);
  and g66136 (n39675, n_234, n_29499);
  and g66137 (n39676, pi0214, n_29478);
  not g66138 (n_29500, n39675);
  and g66139 (n39677, n_29500, n39676);
  not g66140 (n_29501, n39677);
  and g66141 (n39678, n39664, n_29501);
  and g66142 (n39679, n_28588, n38783);
  and g66143 (n39680, n_29487, n39679);
  and g66144 (n39681, n38744, n39674);
  not g66145 (n_29502, n39454);
  and g66146 (n39682, n_234, n_29502);
  not g66147 (n_29503, n39682);
  and g66148 (n39683, n_26242, n_29503);
  and g66149 (n39684, pi0200, n38674);
  not g66150 (n_29504, n39684);
  and g66151 (n39685, n39671, n_29504);
  not g66152 (n_29505, n39683);
  not g66153 (n_29506, n39685);
  and g66154 (n39686, n_29505, n_29506);
  not g66155 (n_29507, n39686);
  and g66156 (n39687, n_28710, n_29507);
  not g66157 (n_29508, n39687);
  and g66158 (n39688, n10484, n_29508);
  not g66165 (n_29512, n39691);
  and g66166 (n39692, n_6791, n_29512);
  not g66167 (n_29513, n39678);
  and g66168 (n39693, n_29513, n39692);
  and g66169 (n39694, pi1151, n_4226);
  and g66170 (n39695, n_7075, n_29507);
  and g66171 (n39696, pi0211, n_29486);
  not g66172 (n_29514, n39695);
  not g66173 (n_29515, n39696);
  and g66174 (n39697, n_29514, n_29515);
  not g66175 (n_29516, n39697);
  and g66176 (n39698, n_28710, n_29516);
  and g66177 (n39699, n38413, n_29487);
  not g66178 (n_29517, n39699);
  and g66179 (n39700, n39698, n_29517);
  not g66180 (n_29518, n39700);
  and g66181 (n39701, pi0219, n_29518);
  not g66182 (n_29519, n39701);
  and g66183 (n39702, n39694, n_29519);
  not g66184 (n_29520, n39693);
  and g66185 (n39703, n_29520, n39702);
  not g66186 (n_29521, n39657);
  and g66187 (n39704, n_28873, n_29521);
  not g66188 (n_29522, n39703);
  and g66189 (n39705, n_29522, n39704);
  and g66190 (n39706, n_7409, n_29000);
  not g66191 (n_29523, n39706);
  and g66192 (n39707, pi0207, n_29523);
  not g66193 (n_29524, n39707);
  and g66194 (n39708, n_28950, n_29524);
  not g66195 (n_29525, n39708);
  and g66196 (n39709, n_26242, n_29525);
  and g66197 (n39710, pi0200, pi0207);
  not g66198 (n_29526, n39710);
  and g66199 (n39711, n_7044, n_29526);
  not g66200 (n_29527, n39711);
  and g66201 (n39712, n_234, n_29527);
  not g66202 (n_29528, n39712);
  and g66203 (n39713, pi0208, n_29528);
  and g66204 (n39714, n_25873, n10809);
  not g66205 (n_29529, n39714);
  and g66206 (n39715, n_234, n_29529);
  not g66207 (n_29530, n39715);
  and g66208 (n39716, n_11757, n_29530);
  not g66209 (n_29531, n39716);
  and g66210 (n39717, n39713, n_29531);
  not g66211 (n_29532, n39709);
  not g66212 (n_29533, n39717);
  and g66213 (n39718, n_29532, n_29533);
  not g66214 (n_29534, n39718);
  and g66215 (n39719, pi0211, n_29534);
  not g66216 (n_29535, n38947);
  and g66217 (n39720, n_25873, n_29535);
  not g66218 (n_29536, n39720);
  and g66219 (n39721, n_29427, n_29536);
  not g66220 (n_29537, n39721);
  and g66221 (n39722, pi0208, n_29537);
  and g66222 (n39723, n38675, n_29535);
  not g66223 (n_29538, n39722);
  not g66224 (n_29539, n39723);
  and g66225 (n39724, n_29538, n_29539);
  and g66226 (n39725, n_7075, n_28757);
  not g66227 (n_29540, n39724);
  and g66228 (n39726, n_29540, n39725);
  not g66229 (n_29541, n39719);
  not g66230 (n_29542, n39726);
  and g66231 (n39727, n_29541, n_29542);
  not g66232 (n_29543, n39727);
  and g66233 (n39728, n10843, n_29543);
  and g66234 (n39729, pi0299, n38489);
  and g66235 (n39730, n_28519, n_29540);
  not g66236 (n_29544, n39729);
  and g66237 (n39731, n_29544, n39730);
  not g66238 (n_29545, n39728);
  not g66239 (n_29546, n39731);
  and g66240 (n39732, n_29545, n_29546);
  not g66241 (n_29547, n39732);
  and g66242 (n39733, n_6791, n_29547);
  and g66243 (n39734, n_6900, n38945);
  and g66244 (n39735, n_28828, n_29502);
  not g66245 (n_29548, n39735);
  and g66246 (n39736, n11384, n_29548);
  not g66247 (n_29549, n39734);
  and g66248 (n39737, n_29549, n39736);
  and g66249 (n39738, n_7075, n38512);
  and g66250 (n39739, n_28511, n39738);
  not g66251 (n_29550, n39737);
  not g66252 (n_29551, n39739);
  and g66253 (n39740, n_29550, n_29551);
  not g66254 (n_29552, n39740);
  and g66255 (n39741, n_28696, n_29552);
  not g66256 (n_29553, n39733);
  not g66257 (n_29554, n39741);
  and g66258 (n39742, n_29553, n_29554);
  not g66259 (n_29555, n39742);
  and g66260 (n39743, n39635, n_29555);
  and g66261 (n39744, n38441, n38561);
  and g66262 (n39745, pi0208, n38550);
  and g66263 (n39746, n_29529, n39745);
  not g66264 (n_29556, n39744);
  not g66265 (n_29557, n39746);
  and g66266 (n39747, n_29556, n_29557);
  and g66267 (n39748, n_26565, n39747);
  and g66268 (n39749, n_29474, n39748);
  not g66269 (n_29558, n39749);
  and g66270 (n39750, n_26538, n_29558);
  and g66271 (n39751, n_26565, n39750);
  not g66272 (n_29559, n38986);
  and g66273 (n39752, n38948, n_29559);
  not g66274 (n_29560, n39752);
  and g66275 (n39753, pi0208, n_29560);
  and g66276 (n39754, n38675, n_28924);
  not g66277 (n_29561, n39753);
  not g66278 (n_29562, n39754);
  and g66279 (n39755, n_29561, n_29562);
  not g66280 (n_29563, n39755);
  and g66281 (n39756, n_7075, n_29563);
  and g66282 (n39757, n_28772, n39756);
  and g66283 (n39758, pi0211, n_29563);
  and g66284 (n39759, n_28757, n39758);
  not g66285 (n_29564, n39757);
  not g66286 (n_29565, n39759);
  and g66287 (n39760, n_29564, n_29565);
  not g66288 (n_29566, n39760);
  and g66289 (n39761, n_28519, n_29566);
  and g66290 (n39762, n_29476, n39747);
  and g66291 (n39763, n_29542, n39762);
  not g66292 (n_29567, n39763);
  and g66293 (n39764, n10843, n_29567);
  and g66300 (n39768, pi0219, n39747);
  and g66301 (n39769, n_29473, n39768);
  not g66302 (n_29571, n39769);
  and g66303 (n39770, n39694, n_29571);
  not g66304 (n_29572, n39767);
  and g66305 (n39771, n_29572, n39770);
  not g66306 (n_29573, n39771);
  and g66307 (n39772, pi1152, n_29573);
  not g66308 (n_29574, n39743);
  and g66309 (n39773, n_29574, n39772);
  not g66310 (n_29575, n39705);
  not g66311 (n_29576, n39773);
  and g66312 (n39774, n_29575, n_29576);
  not g66313 (n_29577, n39774);
  and g66314 (n39775, n_26372, n_29577);
  and g66315 (n39776, n38641, n39032);
  not g66316 (n_29578, n39776);
  and g66317 (n39777, n10487, n_29578);
  and g66318 (n39778, n_28931, n39777);
  not g66319 (n_29579, n39778);
  and g66320 (n39779, n_29151, n_29579);
  not g66321 (n_29580, n39779);
  and g66322 (n39780, n_26565, n_29580);
  and g66323 (n39781, n_26538, n39780);
  and g66324 (n39782, pi0211, n39779);
  and g66325 (n39783, pi1153, n_28630);
  not g66326 (n_29581, n39783);
  and g66327 (n39784, n_28931, n_29581);
  not g66328 (n_29582, n39784);
  and g66329 (n39785, pi0207, n_29582);
  not g66330 (n_29583, n39785);
  and g66331 (n39786, n_29219, n_29583);
  not g66332 (n_29584, n39786);
  and g66333 (n39787, pi0208, n_29584);
  not g66334 (n_29585, n39787);
  and g66335 (n39788, n_29221, n_29585);
  not g66336 (n_29586, n39788);
  and g66337 (n39789, n_7075, n_29586);
  not g66338 (n_29587, n39782);
  not g66339 (n_29588, n39789);
  and g66340 (n39790, n_29587, n_29588);
  and g66341 (n39791, n38970, n39790);
  and g66342 (n39792, n_28618, n39084);
  and g66343 (n39793, n_11413, n_29006);
  and g66344 (n39794, n_28630, n39793);
  not g66345 (n_29589, n39794);
  and g66346 (n39795, pi0207, n_29589);
  and g66347 (n39796, n39001, n39795);
  not g66348 (n_29590, n39796);
  and g66349 (n39797, pi0208, n_29590);
  not g66350 (n_29591, n39792);
  and g66351 (n39798, n_29591, n39797);
  and g66352 (n39799, n_29144, n39798);
  not g66353 (n_29592, n39799);
  and g66354 (n39800, n_29145, n_29592);
  not g66355 (n_29593, n39800);
  and g66356 (n39801, n_7075, n_29593);
  and g66357 (n39802, n39001, n_29578);
  not g66358 (n_29594, n39802);
  and g66359 (n39803, pi0207, n_29594);
  not g66360 (n_29595, n39803);
  and g66361 (n39804, n_29226, n_29595);
  not g66362 (n_29596, n39804);
  and g66363 (n39805, pi0208, n_29596);
  not g66364 (n_29597, n39805);
  and g66365 (n39806, n_29228, n_29597);
  not g66366 (n_29598, n39806);
  and g66367 (n39807, pi0211, n_29598);
  not g66368 (n_29599, n39801);
  and g66369 (n39808, n38421, n_29599);
  not g66370 (n_29600, n39807);
  and g66371 (n39809, n_29600, n39808);
  and g66372 (n39810, n10484, n_29586);
  and g66373 (n39811, n38744, n_29593);
  and g66374 (n39812, n38783, n_29598);
  not g66381 (n_29604, n39809);
  not g66382 (n_29605, n39815);
  and g66383 (n39816, n_29604, n_29605);
  not g66384 (n_29606, n39816);
  and g66385 (n39817, n_6791, n_29606);
  not g66386 (n_29607, n39781);
  not g66392 (n_29610, n39820);
  and g66393 (n39821, pi0209, n_29610);
  not g66394 (n_29611, n39775);
  not g66395 (n_29612, n39821);
  and g66396 (n39822, n_29611, n_29612);
  not g66397 (n_29613, n39634);
  not g66398 (n_29614, n39822);
  and g66399 (n39823, n_29613, n_29614);
  not g66400 (n_29615, n39823);
  and g66401 (n39824, pi0213, n_29615);
  and g66402 (n39825, n_7075, n38608);
  and g66403 (n39826, pi1153, n39825);
  and g66404 (n39827, n39374, n39826);
  not g66405 (n_29616, n39827);
  and g66406 (n39828, n_29468, n_29616);
  and g66407 (n39829, pi0219, n_29471);
  not g66408 (n_29617, n39829);
  and g66409 (n39830, n_4226, n_29617);
  and g66410 (n39831, n_8688, n_29474);
  not g66411 (n_29618, n39640);
  and g66412 (n39832, pi0212, n_29618);
  not g66413 (n_29619, n39831);
  and g66414 (n39833, n_29619, n39832);
  not g66415 (n_29620, n39833);
  and g66416 (n39834, n_6791, n_29620);
  and g66417 (n39835, n39640, n39643);
  and g66418 (n39836, n38421, n39738);
  and g66424 (n39840, n39643, n39830);
  not g66425 (n_29623, n39839);
  and g66426 (n39841, n_29623, n39840);
  not g66427 (n_29624, n39841);
  and g66428 (n39842, n39828, n_29624);
  not g66429 (n_29625, n39826);
  and g66430 (n39843, n10486, n_29625);
  not g66431 (n_29626, n39843);
  and g66432 (n39844, n38416, n_29626);
  not g66433 (n_29627, n39844);
  and g66434 (n39845, pi1151, n_29627);
  and g66435 (n39846, n_26565, n39698);
  and g66436 (n39847, n_29487, n39831);
  not g66437 (n_29628, n39847);
  and g66438 (n39848, pi0214, n_29628);
  not g66439 (n_29629, n39848);
  and g66440 (n39849, pi0212, n_29629);
  not g66441 (n_29630, n39846);
  and g66442 (n39850, n_29630, n39849);
  and g66443 (n39851, n_26538, n_29518);
  not g66444 (n_29631, n39850);
  not g66445 (n_29632, n39851);
  and g66446 (n39852, n_29631, n_29632);
  not g66447 (n_29633, n39852);
  and g66448 (n39853, n_6791, n_29633);
  and g66449 (n39854, n_7075, pi0299);
  not g66450 (n_29634, n39854);
  and g66451 (n39855, n_29474, n_29634);
  and g66452 (n39856, n_29487, n39855);
  not g66453 (n_29635, n39856);
  and g66454 (n39857, n_29517, n_29635);
  not g66455 (n_29636, n39857);
  and g66456 (n39858, pi0219, n_29636);
  not g66457 (n_29637, n39858);
  and g66458 (n39859, n_4226, n_29637);
  not g66459 (n_29638, n39853);
  and g66460 (n39860, n_29638, n39859);
  not g66461 (n_29639, n39860);
  and g66462 (n39861, n39845, n_29639);
  not g66463 (n_29640, n39842);
  and g66464 (n39862, n_28873, n_29640);
  not g66465 (n_29641, n39861);
  and g66466 (n39863, n_29641, n39862);
  and g66467 (n39864, n_6792, n38665);
  and g66468 (n39865, po1038, n39864);
  not g66469 (n_29642, n39631);
  and g66470 (n39866, n_7077, n_29642);
  not g66471 (n_29643, n38527);
  not g66472 (n_29644, n39866);
  and g66473 (n39867, n_29643, n_29644);
  not g66474 (n_29645, n39867);
  and g66475 (n39868, n39865, n_29645);
  and g66476 (n39869, n_6933, n38416);
  not g66477 (n_29646, n39869);
  and g66478 (n39870, pi1151, n_29646);
  not g66479 (n_29647, n39868);
  and g66480 (n39871, n_29647, n39870);
  and g66481 (n39872, n_29474, n39747);
  not g66482 (n_29648, n39756);
  and g66483 (n39873, n_29648, n39872);
  and g66484 (n39874, pi0214, n39873);
  not g66485 (n_29649, n39874);
  and g66486 (n39875, n_29558, n_29649);
  not g66487 (n_29650, n39875);
  and g66488 (n39876, n_26538, n_29650);
  not g66489 (n_29651, n39873);
  not g66490 (n_29652, n39876);
  and g66491 (n39877, n_29651, n_29652);
  not g66492 (n_29653, n39877);
  and g66493 (n39878, pi0219, n_29653);
  not g66494 (n_29654, n39878);
  and g66495 (n39879, n_4226, n_29654);
  and g66496 (n39880, pi1153, n_29470);
  not g66497 (n_29655, n39758);
  not g66498 (n_29656, n39880);
  and g66499 (n39881, n_29655, n_29656);
  and g66500 (n39882, pi0214, n39747);
  and g66501 (n39883, n39881, n39882);
  not g66502 (n_29657, n39883);
  and g66503 (n39884, n39750, n_29657);
  and g66504 (n39885, pi0214, n39755);
  and g66505 (n39886, n39748, n39881);
  not g66506 (n_29658, n39885);
  and g66507 (n39887, pi0212, n_29658);
  not g66508 (n_29659, n39886);
  and g66509 (n39888, n_29659, n39887);
  not g66510 (n_29660, n39884);
  and g66511 (n39889, n_6791, n_29660);
  not g66512 (n_29661, n39888);
  and g66513 (n39890, n_29661, n39889);
  not g66514 (n_29662, n39890);
  and g66515 (n39891, n39879, n_29662);
  not g66516 (n_29663, n39891);
  and g66517 (n39892, n39871, n_29663);
  and g66518 (n39893, n_29468, n_29647);
  and g66519 (n39894, pi0219, n_29550);
  not g66520 (n_29664, n39894);
  and g66521 (n39895, n_4226, n_29664);
  and g66522 (n39896, n_7075, n39718);
  not g66523 (n_29665, n39896);
  and g66524 (n39897, n39730, n_29665);
  and g66525 (n39898, n_29018, n39737);
  and g66526 (n39899, pi0299, n38527);
  not g66533 (n_29669, n39902);
  and g66534 (n39903, n39895, n_29669);
  not g66535 (n_29670, n39903);
  and g66536 (n39904, n39893, n_29670);
  not g66537 (n_29671, n39904);
  and g66538 (n39905, pi1152, n_29671);
  not g66539 (n_29672, n39892);
  and g66540 (n39906, n_29672, n39905);
  not g66541 (n_29673, n39863);
  not g66542 (n_29674, n39906);
  and g66543 (n39907, n_29673, n_29674);
  and g66544 (n39908, n_26372, n39907);
  and g66545 (n39909, n_6791, n38608);
  not g66546 (n_29675, n39909);
  and g66547 (n39910, n_29580, n_29675);
  and g66548 (n39911, n39790, n39909);
  not g66549 (n_29676, n39910);
  and g66550 (n39912, n_4226, n_29676);
  not g66551 (n_29677, n39911);
  and g66552 (n39913, n_29677, n39912);
  not g66553 (n_29678, n39913);
  and g66554 (n39914, n39828, n_29678);
  and g66555 (n39915, n_29157, n39797);
  not g66556 (n_29679, n39915);
  and g66557 (n39916, n_29159, n_29679);
  not g66558 (n_29680, n39916);
  and g66559 (n39917, n_7075, n_29680);
  not g66560 (n_29681, n39917);
  and g66561 (n39918, n_29587, n_29681);
  and g66562 (n39919, n_28511, n39918);
  not g66563 (n_29682, n39919);
  and g66564 (n39920, n_29607, n_29682);
  not g66565 (n_29683, n39920);
  and g66566 (n39921, pi0219, n_29683);
  not g66567 (n_29684, n39921);
  and g66568 (n39922, n_4226, n_29684);
  and g66569 (n39923, pi0214, n39790);
  not g66570 (n_29685, n39780);
  not g66571 (n_29686, n39923);
  and g66572 (n39924, n_29685, n_29686);
  not g66573 (n_29687, n39924);
  and g66574 (n39925, n_26538, n_29687);
  not g66575 (n_29688, n39790);
  and g66576 (n39926, n_26565, n_29688);
  and g66577 (n39927, pi0211, n_29680);
  and g66578 (n39928, n_7075, n39779);
  not g66579 (n_29689, n39927);
  not g66580 (n_29690, n39928);
  and g66581 (n39929, n_29689, n_29690);
  not g66582 (n_29691, n39929);
  and g66583 (n39930, pi0214, n_29691);
  not g66584 (n_29692, n39926);
  and g66585 (n39931, pi0212, n_29692);
  not g66586 (n_29693, n39930);
  and g66587 (n39932, n_29693, n39931);
  not g66588 (n_29694, n39925);
  not g66589 (n_29695, n39932);
  and g66590 (n39933, n_29694, n_29695);
  not g66591 (n_29696, n39933);
  and g66592 (n39934, n_6791, n_29696);
  not g66593 (n_29697, n39934);
  and g66594 (n39935, n39922, n_29697);
  not g66595 (n_29698, n39935);
  and g66596 (n39936, n39845, n_29698);
  not g66597 (n_29699, n39914);
  and g66598 (n39937, n_28873, n_29699);
  not g66599 (n_29700, n39936);
  and g66600 (n39938, n_29700, n39937);
  and g66601 (n39939, n_29588, n_29689);
  not g66602 (n_29701, n39939);
  and g66603 (n39940, n_26565, n_29701);
  not g66604 (n_29702, n39918);
  and g66605 (n39941, pi0214, n_29702);
  not g66606 (n_29703, n39940);
  not g66607 (n_29704, n39941);
  and g66608 (n39942, n_29703, n_29704);
  not g66609 (n_29705, n39942);
  and g66610 (n39943, pi0212, n_29705);
  and g66611 (n39944, pi0214, n39939);
  and g66612 (n39945, n_26538, n_29685);
  not g66613 (n_29706, n39944);
  and g66614 (n39946, n_29706, n39945);
  not g66615 (n_29707, n39946);
  and g66616 (n39947, n_6791, n_29707);
  not g66617 (n_29708, n39943);
  and g66618 (n39948, n_29708, n39947);
  and g66619 (n39949, pi0219, n_29580);
  not g66620 (n_29709, n39949);
  and g66621 (n39950, n_4226, n_29709);
  not g66622 (n_29710, n39948);
  and g66623 (n39951, n_29710, n39950);
  not g66624 (n_29711, n39951);
  and g66625 (n39952, n39893, n_29711);
  and g66626 (n39953, pi0214, n_29680);
  not g66627 (n_29712, n39953);
  and g66628 (n39954, n_29703, n_29712);
  not g66629 (n_29713, n39954);
  and g66630 (n39955, pi0212, n_29713);
  not g66631 (n_29714, n39955);
  and g66632 (n39956, n39947, n_29714);
  not g66633 (n_29715, n39956);
  and g66634 (n39957, n39922, n_29715);
  not g66635 (n_29716, n39957);
  and g66636 (n39958, n39871, n_29716);
  not g66637 (n_29717, n39952);
  and g66638 (n39959, pi1152, n_29717);
  not g66639 (n_29718, n39958);
  and g66640 (n39960, n_29718, n39959);
  not g66641 (n_29719, n39938);
  and g66642 (n39961, pi0209, n_29719);
  not g66643 (n_29720, n39960);
  and g66644 (n39962, n_29720, n39961);
  not g66645 (n_29721, n39908);
  and g66646 (n39963, n_26557, n_29721);
  not g66647 (n_29722, n39962);
  and g66648 (n39964, n_29722, n39963);
  not g66649 (n_29723, n39824);
  not g66650 (n_29724, n39964);
  and g66651 (n39965, n_29723, n_29724);
  not g66652 (n_29725, n39965);
  and g66653 (n39966, pi0230, n_29725);
  and g66654 (n39967, n_28510, pi0238);
  or g66655 (po0395, n39966, n39967);
  not g66656 (n_29726, n38651);
  and g66657 (n39969, n38449, n_29726);
  not g66658 (n_29727, n39969);
  and g66659 (n39970, pi0212, n_29727);
  not g66660 (n_29728, n39970);
  and g66661 (n39971, n_4226, n_29728);
  and g66662 (n39972, n_26565, n39969);
  not g66663 (n_29729, n39972);
  and g66664 (n39973, n_26538, n_29729);
  and g66665 (n39974, n_6791, n39973);
  and g66666 (n39975, pi0299, pi1158);
  not g66667 (n_29730, n38449);
  and g66668 (n39976, n_29730, n39975);
  and g66669 (n39977, n_26242, n39595);
  not g66670 (n_29731, n39976);
  not g66671 (n_29732, n39977);
  and g66672 (n39978, n_29731, n_29732);
  not g66673 (n_29733, n39978);
  and g66674 (n39979, n_7075, n_29733);
  and g66675 (n39980, n_11810, n_29727);
  and g66676 (n39981, pi0208, pi0299);
  not g66677 (n_29734, n39981);
  and g66678 (n39982, pi1157, n_29734);
  and g66679 (n39983, n_28878, n39982);
  not g66680 (n_29735, n39980);
  and g66681 (n39984, pi0211, n_29735);
  not g66682 (n_29736, n39983);
  and g66683 (n39985, n_29736, n39984);
  not g66684 (n_29737, n39979);
  not g66685 (n_29738, n39985);
  and g66686 (n39986, n_29737, n_29738);
  not g66687 (n_29739, n39986);
  and g66688 (n39987, pi0214, n_29739);
  not g66689 (n_29740, n39987);
  and g66690 (n39988, n39974, n_29740);
  and g66691 (n39989, pi0219, n39973);
  and g66692 (n39990, pi0211, n_29727);
  not g66693 (n_29741, n39990);
  and g66694 (n39991, pi0214, n_29741);
  and g66695 (n39992, n_28850, n39092);
  not g66696 (n_29742, n39992);
  and g66697 (n39993, n39991, n_29742);
  not g66698 (n_29743, n39993);
  and g66699 (n39994, n39989, n_29743);
  and g66705 (n39998, n_6791, n_29266);
  not g66706 (n_29746, n39377);
  not g66707 (n_29747, n39998);
  and g66708 (n39999, n_29746, n_29747);
  and g66709 (n40000, n39447, n_29411);
  and g66710 (n40001, n_26565, n40000);
  not g66711 (n_29748, n40001);
  and g66712 (n40002, n_26538, n_29748);
  and g66713 (n40003, n_6791, n40002);
  and g66714 (n40004, n_29423, n39982);
  not g66715 (n_29749, n40004);
  and g66716 (n40005, n_29411, n_29749);
  not g66717 (n_29750, n40005);
  and g66718 (n40006, pi0211, n_29750);
  not g66719 (n_29751, n39975);
  and g66720 (n40007, pi0208, n_29751);
  not g66721 (n_29752, n38542);
  not g66722 (n_29753, n40007);
  and g66723 (n40008, n_29752, n_29753);
  and g66724 (n40009, n_29437, n40008);
  not g66725 (n_29754, n40009);
  and g66726 (n40010, n39608, n_29754);
  not g66727 (n_29755, n40006);
  and g66728 (n40011, pi0214, n_29755);
  not g66729 (n_29756, n40010);
  and g66730 (n40012, n_29756, n40011);
  not g66731 (n_29757, n40012);
  and g66732 (n40013, n40003, n_29757);
  not g66733 (n_29758, n40000);
  and g66734 (n40014, pi0212, n_29758);
  not g66735 (n_29759, n40014);
  and g66736 (n40015, n_4226, n_29759);
  and g66737 (n40016, pi0219, n40002);
  and g66738 (n40017, pi0211, n_29758);
  and g66739 (n40018, n39092, n_29758);
  not g66740 (n_29760, n40018);
  and g66741 (n40019, pi0214, n_29760);
  not g66742 (n_29761, n40017);
  and g66743 (n40020, n_29761, n40019);
  not g66744 (n_29762, n40020);
  and g66745 (n40021, n40016, n_29762);
  and g66757 (n40028, po1038, n_29079);
  not g66758 (n_29768, n39149);
  and g66759 (n40029, n38421, n_29768);
  and g66760 (n40030, n40028, n40029);
  and g66761 (n40031, pi0211, n_28743);
  and g66762 (n40032, n_29331, n40031);
  not g66763 (n_29769, n40032);
  and g66764 (n40033, n40019, n_29769);
  not g66765 (n_29770, n40033);
  and g66766 (n40034, n40003, n_29770);
  and g66767 (n40035, n_7075, n_28588);
  and g66768 (n40036, n_29331, n40035);
  and g66769 (n40037, pi0214, n_29761);
  not g66770 (n_29771, n40036);
  and g66771 (n40038, n_29771, n40037);
  not g66772 (n_29772, n40038);
  and g66773 (n40039, n40016, n_29772);
  not g66774 (n_29773, n40034);
  and g66775 (n40040, n40015, n_29773);
  not g66776 (n_29774, n40039);
  and g66777 (n40041, n_29774, n40040);
  not g66778 (n_29775, n40041);
  and g66779 (n40042, pi0209, n_29775);
  and g66780 (n40043, n_28588, n_28841);
  not g66781 (n_29776, n40043);
  and g66782 (n40044, n39991, n_29776);
  not g66783 (n_29777, n40044);
  and g66784 (n40045, n39989, n_29777);
  and g66785 (n40046, n_28856, n40031);
  not g66786 (n_29778, n40046);
  and g66787 (n40047, pi0214, n_29778);
  and g66788 (n40048, n_29742, n40047);
  not g66789 (n_29779, n40048);
  and g66790 (n40049, n39974, n_29779);
  not g66791 (n_29780, n40049);
  and g66792 (n40050, n39971, n_29780);
  not g66793 (n_29781, n40045);
  and g66794 (n40051, n_29781, n40050);
  not g66795 (n_29782, n40051);
  and g66796 (n40052, n_26372, n_29782);
  not g66797 (n_29783, n40042);
  not g66798 (n_29784, n40052);
  and g66799 (n40053, n_29783, n_29784);
  not g66800 (n_29785, n40030);
  and g66801 (n40054, n_26557, n_29785);
  not g66802 (n_29786, n40053);
  and g66803 (n40055, n_29786, n40054);
  not g66804 (n_29787, n40027);
  not g66805 (n_29788, n40055);
  and g66806 (n40056, n_29787, n_29788);
  not g66807 (n_29789, n40056);
  and g66808 (n40057, pi0230, n_29789);
  and g66809 (n40058, n_28510, n_906);
  not g66810 (n_29790, n40057);
  not g66811 (n_29791, n40058);
  and g66812 (po0396, n_29790, n_29791);
  and g66813 (n40060, n_4226, n39736);
  not g66814 (n_29792, n39830);
  not g66815 (n_29793, n40060);
  and g66816 (n40061, n_29792, n_29793);
  not g66817 (n_29794, n39736);
  and g66818 (n40062, n_26565, n_29794);
  not g66819 (n_29795, n40062);
  and g66820 (n40063, n_26538, n_29795);
  and g66821 (n40064, n11384, n38449);
  not g66822 (n_29796, n40064);
  and g66823 (n40065, n_234, n_29796);
  not g66824 (n_29797, n39713);
  and g66825 (n40066, n_29797, n40065);
  and g66826 (n40067, pi0214, n40066);
  not g66827 (n_29798, n40067);
  and g66828 (n40068, n40063, n_29798);
  not g66829 (n_29799, n40068);
  and g66830 (n40069, n_6791, n_29799);
  and g66831 (n40070, pi0211, n39736);
  not g66832 (n_29800, n40066);
  and g66833 (n40071, n_7075, n_29800);
  not g66834 (n_29801, n40070);
  and g66835 (n40072, pi0214, n_29801);
  not g66836 (n_29802, n40071);
  and g66837 (n40073, n_29802, n40072);
  not g66838 (n_29803, n40073);
  and g66839 (n40074, pi0212, n_29803);
  and g66840 (n40075, n_29800, n40074);
  not g66841 (n_29804, n40075);
  and g66842 (n40076, n40069, n_29804);
  not g66843 (n_29805, n40061);
  not g66844 (n_29806, n40076);
  and g66845 (n40077, n_29805, n_29806);
  not g66846 (n_29807, n39865);
  not g66847 (n_29808, n40077);
  and g66848 (n40078, n_29807, n_29808);
  not g66849 (n_29810, pi1147);
  and g66850 (n40079, n_29810, n40078);
  and g66851 (n40080, n_7075, po1038);
  not g66852 (n_29811, n40080);
  and g66853 (n40081, n_29267, n_29811);
  not g66854 (n_29812, n40081);
  and g66855 (n40082, n_28511, n_29812);
  and g66856 (n40083, pi0299, n_28511);
  and g66857 (n40084, n_4226, n_28513);
  and g66858 (n40085, n40083, n40084);
  and g66859 (n40086, n38550, n_28825);
  and g66860 (n40087, n_4226, n40086);
  not g66861 (n_29813, n40085);
  not g66862 (n_29814, n40087);
  and g66863 (n40088, n_29813, n_29814);
  not g66864 (n_29815, n40082);
  and g66865 (n40089, n_29815, n40088);
  and g66866 (n40090, pi1147, n40089);
  not g66867 (n_29817, n40090);
  and g66868 (n40091, pi1149, n_29817);
  not g66869 (n_29818, n40079);
  and g66870 (n40092, n_29818, n40091);
  and g66871 (n40093, pi0211, n38421);
  and g66872 (n40094, pi0212, n38783);
  not g66873 (n_29819, n40093);
  not g66874 (n_29820, n40094);
  and g66875 (n40095, n_29819, n_29820);
  not g66876 (n_29821, n40095);
  and g66877 (n40096, n39374, n_29821);
  and g66878 (n40097, n_28828, n_29427);
  and g66879 (n40098, n_6900, n38533);
  not g66880 (n_29822, n40097);
  not g66881 (n_29823, n40098);
  and g66882 (n40099, n_29822, n_29823);
  and g66883 (n40100, n39715, n40099);
  and g66884 (n40101, pi0299, n10484);
  not g66885 (n_29824, n40100);
  not g66886 (n_29825, n40101);
  and g66887 (n40102, n_29824, n_29825);
  not g66888 (n_29826, n40102);
  and g66889 (n40103, n_26538, n_29826);
  not g66890 (n_29827, n40103);
  and g66891 (n40104, n_6791, n_29827);
  not g66892 (n_29828, n40099);
  and g66893 (n40105, n_234, n_29828);
  not g66894 (n_29829, n40105);
  and g66895 (n40106, pi0214, n_29829);
  and g66896 (n40107, n_26565, n40100);
  not g66897 (n_29830, n40107);
  and g66898 (n40108, n_26538, n_29830);
  not g66899 (n_29831, n40106);
  and g66900 (n40109, n_29831, n40108);
  and g66901 (n40110, n_7075, n_29829);
  not g66902 (n_29832, n40110);
  and g66903 (n40111, n_29824, n_29832);
  not g66904 (n_29833, n40111);
  and g66905 (n40112, pi0214, n_29833);
  not g66906 (n_29834, n40112);
  and g66907 (n40113, pi0212, n_29834);
  and g66908 (n40114, n_26565, n_29829);
  not g66909 (n_29835, n40114);
  and g66910 (n40115, n40113, n_29835);
  not g66911 (n_29836, n40109);
  not g66912 (n_29837, n40115);
  and g66913 (n40116, n_29836, n_29837);
  and g66914 (n40117, n_8688, n_29824);
  and g66915 (n40118, n_29831, n40117);
  not g66916 (n_29838, n40118);
  and g66917 (n40119, pi0212, n_29838);
  and g66918 (n40120, n40116, n40119);
  not g66919 (n_29839, n40120);
  and g66920 (n40121, n40104, n_29839);
  and g66921 (n40122, pi0219, n_29824);
  not g66922 (n_29840, n40122);
  and g66923 (n40123, n_4226, n_29840);
  not g66924 (n_29841, n40121);
  and g66925 (n40124, n_29841, n40123);
  not g66926 (n_29842, n40096);
  not g66927 (n_29843, n40124);
  and g66928 (n40125, n_29842, n_29843);
  and g66929 (n40126, n_29810, n40125);
  not g66930 (n_29844, n39747);
  and g66931 (n40127, n_4226, n_29844);
  and g66932 (n40128, pi0212, n_28789);
  and g66933 (n40129, n_6791, n_29819);
  not g66934 (n_29845, n40128);
  and g66935 (n40130, n_29845, n40129);
  not g66936 (n_29846, n40130);
  and g66937 (n40131, n38416, n_29846);
  and g66938 (n40132, n40085, n_29846);
  not g66939 (n_29847, n40127);
  not g66940 (n_29848, n40131);
  and g66941 (n40133, n_29847, n_29848);
  not g66942 (n_29849, n40132);
  and g66943 (n40134, n_29849, n40133);
  and g66944 (n40135, pi1147, n40134);
  not g66945 (n_29850, pi1149);
  not g66946 (n_29851, n40135);
  and g66947 (n40136, n_29850, n_29851);
  not g66948 (n_29852, n40126);
  and g66949 (n40137, n_29852, n40136);
  not g66950 (n_29853, n40092);
  not g66951 (n_29854, n40137);
  and g66952 (n40138, n_29853, n_29854);
  not g66953 (n_29856, n40138);
  and g66954 (n40139, pi1148, n_29856);
  and g66955 (n40140, n16479, n39636);
  and g66956 (n40141, n_6791, n_25711);
  and g66957 (n40142, n39825, n40141);
  not g66958 (n_29857, n40140);
  not g66959 (n_29858, n40142);
  and g66960 (n40143, n_29857, n_29858);
  and g66961 (n40144, n_29810, n40143);
  not g66962 (n_29859, n39825);
  and g66963 (n40145, n10486, n_29859);
  not g66964 (n_29860, n40145);
  and g66965 (n40146, n38416, n_29860);
  and g66966 (n40147, n_7075, n_29486);
  and g66967 (n40148, pi0211, n_29507);
  not g66968 (n_29861, n40148);
  and g66969 (n40149, pi0214, n_29861);
  not g66970 (n_29862, n40147);
  and g66971 (n40150, n_29862, n40149);
  not g66972 (n_29863, n40150);
  and g66973 (n40151, n10843, n_29863);
  and g66974 (n40152, n_26565, n39661);
  not g66975 (n_29864, n40152);
  and g66976 (n40153, n_26538, n_29864);
  and g66977 (n40154, pi0214, n39697);
  not g66978 (n_29865, n40154);
  and g66979 (n40155, n40153, n_29865);
  not g66980 (n_29866, n40155);
  and g66981 (n40156, n_6791, n_29866);
  and g66982 (n40157, pi0212, n_29863);
  and g66983 (n40158, n_29516, n40157);
  not g66984 (n_29867, n40158);
  and g66985 (n40159, n40156, n_29867);
  not g66986 (n_29868, n40151);
  and g66987 (n40160, n_29868, n40159);
  and g66988 (n40161, pi0212, n_29516);
  not g66989 (n_29869, n40161);
  and g66990 (n40162, pi0219, n_29869);
  and g66991 (n40163, n_29866, n40162);
  not g66992 (n_29870, n40163);
  and g66993 (n40164, n_4226, n_29870);
  not g66994 (n_29871, n40160);
  and g66995 (n40165, n_29871, n40164);
  not g66996 (n_29872, n40146);
  not g66997 (n_29873, n40165);
  and g66998 (n40166, n_29872, n_29873);
  and g66999 (n40167, pi1147, n40166);
  not g67000 (n_29874, n40144);
  and g67001 (n40168, pi1149, n_29874);
  not g67002 (n_29875, n40167);
  and g67003 (n40169, n_29875, n40168);
  and g67004 (n40170, n_26538, n_29825);
  and g67005 (n40171, n39747, n40170);
  and g67006 (n40172, n39747, n_29634);
  not g67007 (n_29876, n39748);
  not g67008 (n_29877, n40172);
  and g67009 (n40173, n_29876, n_29877);
  and g67010 (n40174, n_26565, n13061);
  not g67011 (n_29878, n40174);
  and g67012 (n40175, pi0212, n_29878);
  not g67013 (n_29879, n40173);
  and g67014 (n40176, n_29879, n40175);
  not g67015 (n_29880, n40171);
  not g67016 (n_29881, n40176);
  and g67017 (n40177, n_29880, n_29881);
  not g67018 (n_29882, n40177);
  and g67019 (n40178, n_6791, n_29882);
  and g67020 (n40179, n38700, n_29526);
  not g67021 (n_29883, n40179);
  and g67022 (n40180, pi0208, n_29883);
  not g67023 (n_29884, n40180);
  and g67024 (n40181, n_7044, n_29884);
  not g67025 (n_29885, n40181);
  and g67026 (n40182, n_29844, n_29885);
  not g67027 (n_29886, n40182);
  and g67028 (n40183, n_234, n_29886);
  and g67029 (n40184, n_6791, n40183);
  not g67030 (n_29887, n40178);
  not g67031 (n_29888, n40184);
  and g67032 (n40185, n_29887, n_29888);
  not g67033 (n_29889, n40185);
  and g67034 (n40186, n_7075, n_29889);
  and g67035 (n40187, n_8688, n39882);
  and g67036 (n40188, n_26565, n40172);
  not g67037 (n_29890, n40188);
  and g67038 (n40189, pi0212, n_29890);
  not g67039 (n_29891, n40187);
  and g67040 (n40190, n_29891, n40189);
  and g67041 (n40191, n_26538, n40173);
  not g67042 (n_29892, n40191);
  and g67043 (n40192, n_6791, n_29892);
  not g67044 (n_29893, n40190);
  and g67045 (n40193, n_29893, n40192);
  and g67046 (n40194, pi0219, n_29634);
  not g67047 (n_29894, n40194);
  and g67048 (n40195, n40084, n_29894);
  not g67049 (n_29895, n40195);
  and g67050 (n40196, n_29847, n_29895);
  not g67051 (n_29896, n40193);
  not g67052 (n_29897, n40196);
  and g67053 (n40197, n_29896, n_29897);
  not g67054 (n_29898, n40183);
  and g67055 (n40198, n_29898, n40197);
  not g67056 (n_29899, n40186);
  and g67057 (n40199, n_29899, n40198);
  not g67058 (n_29900, n40199);
  and g67059 (n40200, n_29646, n_29900);
  and g67060 (n40201, pi1147, n_29850);
  not g67061 (n_29901, n40200);
  and g67062 (n40202, n_29901, n40201);
  not g67063 (n_29902, n40169);
  not g67064 (n_29903, n40202);
  and g67065 (n40203, n_29902, n_29903);
  not g67066 (n_29904, pi1148);
  not g67067 (n_29905, n40203);
  and g67068 (n40204, n_29904, n_29905);
  not g67069 (n_29906, n40139);
  not g67070 (n_29907, n40204);
  and g67071 (n40205, n_29906, n_29907);
  not g67072 (n_29908, n40205);
  and g67073 (n40206, pi0213, n_29908);
  and g67074 (n40207, n10846, n38665);
  and g67075 (n40208, po1038, n40207);
  and g67076 (n40209, n_7075, pi1146);
  and g67077 (n40210, pi0211, pi1145);
  not g67078 (n_29909, n40209);
  not g67079 (n_29910, n40210);
  and g67080 (n40211, n_29909, n_29910);
  not g67081 (n_29911, n40211);
  and g67082 (n40212, pi0214, n_29911);
  and g67083 (n40213, pi0211, pi1146);
  and g67084 (n40214, n_26565, n40213);
  not g67085 (n_29912, n40212);
  not g67086 (n_29913, n40214);
  and g67087 (n40215, n_29912, n_29913);
  not g67088 (n_29914, n40215);
  and g67089 (n40216, pi0212, n_29914);
  and g67090 (n40217, n38421, n40213);
  not g67091 (n_29915, n40216);
  not g67092 (n_29916, n40217);
  and g67093 (n40218, n_29915, n_29916);
  and g67094 (n40219, n_28940, n40218);
  and g67095 (n40220, po1038, n39412);
  not g67096 (n_29917, n40220);
  and g67097 (n40221, n_29267, n_29917);
  not g67098 (n_29918, n40219);
  not g67099 (n_29919, n40221);
  and g67100 (n40222, n_29918, n_29919);
  not g67101 (n_29920, n40208);
  and g67102 (n40223, pi1147, n_29920);
  not g67103 (n_29921, n40222);
  and g67104 (n40224, n_29921, n40223);
  and g67105 (n40225, n_7075, n39484);
  not g67106 (n_29922, n40225);
  and g67107 (n40226, pi0219, n_29922);
  not g67108 (n_29923, n40226);
  and g67109 (n40227, n40084, n_29923);
  not g67110 (n_29924, n40227);
  and g67111 (n40228, n_29847, n_29924);
  and g67112 (n40229, n38413, n_29844);
  not g67113 (n_29925, n40229);
  and g67114 (n40230, n_6791, n_29925);
  and g67115 (n40231, pi0299, n_29911);
  not g67116 (n_29926, n40231);
  and g67117 (n40232, n39747, n_29926);
  not g67118 (n_29927, n40232);
  and g67119 (n40233, n10843, n_29927);
  and g67120 (n40234, pi0299, pi1146);
  and g67121 (n40235, pi0211, n40234);
  not g67122 (n_29928, n40235);
  and g67123 (n40236, n_29634, n_29928);
  and g67124 (n40237, n39747, n40236);
  not g67125 (n_29929, n40237);
  and g67126 (n40238, n38608, n_29929);
  not g67127 (n_29930, n40233);
  and g67128 (n40239, n40230, n_29930);
  not g67129 (n_29931, n40238);
  and g67130 (n40240, n_29931, n40239);
  not g67131 (n_29932, n40228);
  not g67132 (n_29933, n40240);
  and g67133 (n40241, n_29932, n_29933);
  not g67134 (n_29934, n40241);
  and g67135 (n40242, n40224, n_29934);
  and g67136 (n40243, n_4226, n40100);
  and g67137 (n40244, n_29810, n_29921);
  and g67138 (n40245, pi0219, n40227);
  not g67139 (n_29935, n40218);
  and g67140 (n40246, pi0299, n_29935);
  and g67141 (n40247, n36114, n40246);
  not g67142 (n_29936, n40245);
  not g67143 (n_29937, n40247);
  and g67144 (n40248, n_29936, n_29937);
  and g67145 (n40249, n40244, n40248);
  not g67146 (n_29938, n40243);
  and g67147 (n40250, n_29938, n40249);
  not g67148 (n_29939, n40242);
  and g67149 (n40251, pi1148, n_29939);
  not g67150 (n_29940, n40250);
  and g67151 (n40252, n_29940, n40251);
  and g67152 (n40253, n39412, n39422);
  and g67153 (n40254, n_28696, n40182);
  and g67154 (n40255, n_803, n13061);
  not g67155 (n_29941, n40255);
  and g67156 (n40256, n38608, n_29941);
  not g67157 (n_29942, n40256);
  and g67158 (n40257, n_29930, n_29942);
  and g67159 (n40258, n_6791, n_29898);
  not g67160 (n_29943, n40257);
  and g67161 (n40259, n_29943, n40258);
  not g67162 (n_29944, n40253);
  not g67163 (n_29945, n40254);
  and g67164 (n40260, n_29944, n_29945);
  not g67165 (n_29946, n40259);
  and g67166 (n40261, n_29946, n40260);
  not g67167 (n_29947, n40261);
  and g67168 (n40262, n_4226, n_29947);
  not g67169 (n_29948, n40262);
  and g67170 (n40263, n40224, n_29948);
  not g67171 (n_29949, n40249);
  and g67172 (n40264, n_29904, n_29949);
  not g67173 (n_29950, n40263);
  and g67174 (n40265, n_29950, n40264);
  not g67175 (n_29951, n40252);
  not g67176 (n_29952, n40265);
  and g67177 (n40266, n_29951, n_29952);
  not g67178 (n_29953, n40266);
  and g67179 (n40267, n_29850, n_29953);
  and g67180 (n40268, pi0219, n39661);
  not g67181 (n_29954, n40268);
  and g67182 (n40269, n_4226, n_29954);
  not g67183 (n_29955, n40269);
  and g67184 (n40270, n_29924, n_29955);
  and g67185 (n40271, n_234, n39685);
  not g67186 (n_29956, n39431);
  not g67187 (n_29957, n40271);
  and g67188 (n40272, n_29956, n_29957);
  not g67189 (n_29958, n40234);
  and g67190 (n40273, n_29958, n40272);
  not g67191 (n_29959, n40273);
  and g67192 (n40274, pi0211, n_29959);
  not g67193 (n_29960, n40274);
  and g67194 (n40275, n_29514, n_29960);
  and g67195 (n40276, pi0214, n40275);
  not g67196 (n_29961, n40276);
  and g67197 (n40277, n40153, n_29961);
  and g67198 (n40278, pi0214, n_29926);
  and g67199 (n40279, n40272, n40278);
  and g67200 (n40280, n_26565, n40275);
  not g67201 (n_29962, n40279);
  and g67202 (n40281, pi0212, n_29962);
  not g67203 (n_29963, n40280);
  and g67204 (n40282, n_29963, n40281);
  not g67205 (n_29964, n40277);
  and g67206 (n40283, n_6791, n_29964);
  not g67207 (n_29965, n40282);
  and g67208 (n40284, n_29965, n40283);
  not g67209 (n_29966, n40270);
  not g67210 (n_29967, n40284);
  and g67211 (n40285, n_29966, n_29967);
  not g67212 (n_29968, n40285);
  and g67213 (n40286, n40224, n_29968);
  and g67214 (n40287, n_29857, n40249);
  not g67215 (n_29969, n40287);
  and g67216 (n40288, n_29904, n_29969);
  not g67217 (n_29970, n40286);
  and g67218 (n40289, n_29970, n40288);
  not g67219 (n_29971, n40086);
  and g67220 (n40290, pi0219, n_29971);
  not g67221 (n_29972, n40290);
  and g67222 (n40291, n_4226, n_29972);
  and g67223 (n40292, pi0211, n_29971);
  and g67224 (n40293, pi0214, pi0299);
  not g67225 (n_29973, n40293);
  and g67226 (n40294, n_29971, n_29973);
  not g67227 (n_29974, n40294);
  and g67228 (n40295, n_26538, n_29974);
  not g67229 (n_29975, n40292);
  and g67230 (n40296, n_29975, n40295);
  and g67231 (n40297, n_234, n_29971);
  not g67232 (n_29976, n40297);
  and g67233 (n40298, pi0212, n_29976);
  and g67234 (n40299, pi0299, n40128);
  not g67235 (n_29977, n40299);
  and g67236 (n40300, n40298, n_29977);
  not g67237 (n_29978, n40296);
  and g67238 (n40301, n_6791, n_29978);
  not g67239 (n_29979, n40300);
  and g67240 (n40302, n_29979, n40301);
  not g67241 (n_29980, n40302);
  and g67242 (n40303, n40291, n_29980);
  and g67243 (n40304, n40224, n40248);
  not g67244 (n_29981, n40303);
  and g67245 (n40305, n_29981, n40304);
  and g67246 (n40306, n_28512, n39736);
  and g67247 (n40307, n_28511, n40071);
  not g67248 (n_29982, n40306);
  and g67249 (n40308, pi0219, n_29982);
  not g67250 (n_29983, n40307);
  and g67251 (n40309, n_29983, n40308);
  not g67252 (n_29984, n40309);
  and g67253 (n40310, n_4226, n_29984);
  and g67254 (n40311, n11384, n40310);
  not g67255 (n_29985, n40311);
  and g67256 (n40312, n_29924, n_29985);
  and g67257 (n40313, n_29794, n_29928);
  not g67258 (n_29986, n40313);
  and g67259 (n40314, n40063, n_29986);
  and g67260 (n40315, pi0212, n_29800);
  and g67261 (n40316, n_29794, n40215);
  not g67262 (n_29987, n40316);
  and g67263 (n40317, n40315, n_29987);
  not g67264 (n_29988, n40314);
  and g67265 (n40318, n_6791, n_29988);
  not g67266 (n_29989, n40317);
  and g67267 (n40319, n_29989, n40318);
  not g67268 (n_29990, n40312);
  not g67269 (n_29991, n40319);
  and g67270 (n40320, n_29990, n_29991);
  not g67271 (n_29992, n40320);
  and g67272 (n40321, n40244, n_29992);
  not g67273 (n_29993, n40305);
  and g67274 (n40322, pi1148, n_29993);
  not g67275 (n_29994, n40321);
  and g67276 (n40323, n_29994, n40322);
  not g67277 (n_29995, n40289);
  not g67278 (n_29996, n40323);
  and g67279 (n40324, n_29995, n_29996);
  not g67280 (n_29997, n40324);
  and g67281 (n40325, pi1149, n_29997);
  not g67282 (n_29998, n40267);
  not g67283 (n_29999, n40325);
  and g67284 (n40326, n_29998, n_29999);
  not g67285 (n_30000, n40326);
  and g67286 (n40327, n_26557, n_30000);
  not g67287 (n_30001, n40327);
  and g67288 (n40328, pi0209, n_30001);
  not g67289 (n_30002, n40206);
  and g67290 (n40329, n_30002, n40328);
  and g67291 (n40330, pi0200, n_29278);
  and g67292 (n40331, pi0199, pi1145);
  not g67293 (n_30003, n40331);
  and g67294 (n40332, n_7045, n_30003);
  and g67295 (n40333, n_7044, pi1146);
  not g67296 (n_30004, n40333);
  and g67297 (n40334, n40332, n_30004);
  not g67298 (n_30005, n40330);
  and g67299 (n40335, n38441, n_30005);
  not g67300 (n_30006, n40334);
  and g67301 (n40336, n_30006, n40335);
  not g67302 (n_30007, n40336);
  and g67303 (n40337, n_28828, n_30007);
  and g67304 (n40338, pi0200, n_30004);
  not g67305 (n_30008, n40338);
  and g67306 (n40339, n_234, n_30008);
  not g67307 (n_30009, n40332);
  and g67308 (n40340, n_30009, n40339);
  not g67309 (n_30010, n40340);
  and g67310 (n40341, n_6900, n_30010);
  not g67311 (n_30011, n40337);
  not g67312 (n_30012, n40341);
  and g67313 (n40342, n_30011, n_30012);
  and g67314 (n40343, n38413, n40342);
  not g67315 (n_30013, n40343);
  and g67316 (n40344, pi0219, n_30013);
  and g67317 (n40345, n_28511, n40342);
  not g67318 (n_30014, n40345);
  and g67319 (n40346, n_28512, n_30014);
  and g67320 (n40347, n38699, n_30003);
  not g67321 (n_30015, n40347);
  and g67322 (n40348, n40339, n_30015);
  and g67323 (n40349, n_25873, n40348);
  and g67324 (n40350, n40332, n40349);
  and g67325 (n40351, n_29958, n_30007);
  not g67326 (n_30016, n40349);
  and g67327 (n40352, n_30016, n40351);
  not g67328 (n_30017, n40352);
  and g67329 (n40353, pi0208, n_30017);
  not g67330 (n_30018, n40350);
  and g67331 (n40354, n_30018, n40353);
  and g67332 (n40355, n38449, n40340);
  not g67333 (n_30019, n40354);
  not g67334 (n_30020, n40355);
  and g67335 (n40356, n_30019, n_30020);
  not g67336 (n_30021, n40356);
  and g67337 (n40357, n_234, n_30021);
  and g67338 (n40358, n_7075, n_29346);
  not g67339 (n_30022, n40357);
  and g67340 (n40359, n_30022, n40358);
  not g67341 (n_30023, n40346);
  not g67342 (n_30024, n40359);
  and g67343 (n40360, n_30023, n_30024);
  not g67344 (n_30025, n40360);
  and g67345 (n40361, n40344, n_30025);
  not g67346 (n_30026, n40342);
  and g67347 (n40362, n_29928, n_30026);
  and g67348 (n40363, n_26565, n_30026);
  not g67349 (n_30027, n40363);
  and g67350 (n40364, n_26538, n_30027);
  not g67351 (n_30028, n40362);
  and g67352 (n40365, n_30028, n40364);
  not g67353 (n_30029, n40365);
  and g67354 (n40366, n_6791, n_30029);
  and g67355 (n40367, n40278, n_30022);
  and g67356 (n40368, n_26565, n40362);
  not g67357 (n_30030, n40368);
  and g67358 (n40369, pi0212, n_30030);
  not g67359 (n_30031, n40367);
  and g67360 (n40370, n_30031, n40369);
  not g67361 (n_30032, n40370);
  and g67362 (n40371, n40366, n_30032);
  not g67363 (n_30033, n40361);
  and g67364 (n40372, n_4226, n_30033);
  not g67365 (n_30034, n40371);
  and g67366 (n40373, n_30034, n40372);
  not g67367 (n_30035, n40373);
  and g67368 (n40374, n40244, n_30035);
  not g67369 (n_30036, n40348);
  and g67370 (n40375, n_6900, n_30036);
  not g67371 (n_30037, n40375);
  and g67372 (n40376, n_30011, n_30037);
  and g67373 (n40377, n_28512, n40376);
  not g67374 (n_30038, n40377);
  and g67375 (n40378, pi0219, n_30038);
  and g67376 (n40379, n38449, n40348);
  not g67377 (n_30039, n40353);
  not g67378 (n_30040, n40379);
  and g67379 (n40380, n_30039, n_30040);
  and g67380 (n40381, n_234, n40380);
  not g67381 (n_30041, n40381);
  and g67382 (n40382, n_7075, n_30041);
  and g67383 (n40383, n_29345, n40382);
  and g67384 (n40384, n_28511, n40383);
  not g67385 (n_30042, n40384);
  and g67386 (n40385, n40378, n_30042);
  not g67387 (n_30043, n40376);
  not g67388 (n_30044, n40382);
  and g67389 (n40386, n_30043, n_30044);
  and g67390 (n40387, n_26565, n_30043);
  not g67391 (n_30045, n40387);
  and g67392 (n40388, n_26538, n_30045);
  not g67393 (n_30046, n40386);
  and g67394 (n40389, n_30046, n40388);
  and g67395 (n40390, pi0211, n_30041);
  and g67396 (n40391, n_29345, n40390);
  and g67397 (n40392, n40278, n40380);
  and g67398 (n40393, n10484, n_30041);
  not g67399 (n_30047, n40392);
  not g67400 (n_30048, n40393);
  and g67401 (n40394, n_30047, n_30048);
  not g67402 (n_30049, n40391);
  not g67403 (n_30050, n40394);
  and g67404 (n40395, n_30049, n_30050);
  and g67405 (n40396, n_26565, n40236);
  and g67406 (n40397, n40380, n40396);
  not g67407 (n_30051, n40397);
  and g67408 (n40398, pi0212, n_30051);
  not g67409 (n_30052, n40395);
  and g67410 (n40399, n_30052, n40398);
  not g67411 (n_30053, n40389);
  and g67412 (n40400, n40366, n_30053);
  not g67413 (n_30054, n40399);
  and g67414 (n40401, n_30054, n40400);
  not g67415 (n_30055, n40385);
  and g67416 (n40402, n_4226, n_30055);
  not g67417 (n_30056, n40401);
  and g67418 (n40403, n_30056, n40402);
  not g67419 (n_30057, n40403);
  and g67420 (n40404, n40224, n_30057);
  not g67421 (n_30058, n40374);
  not g67422 (n_30059, n40404);
  and g67423 (n40405, n_30058, n_30059);
  and g67424 (n40406, n_26557, n40405);
  and g67425 (n40407, pi1147, n_29848);
  and g67426 (n40408, n_28511, n40382);
  not g67427 (n_30060, n40408);
  and g67428 (n40409, n40378, n_30060);
  not g67429 (n_30061, n40409);
  and g67430 (n40410, n_4226, n_30061);
  and g67431 (n40411, n_234, n40356);
  not g67432 (n_30062, n40411);
  and g67433 (n40412, pi0214, n_30062);
  not g67434 (n_30063, n40390);
  not g67435 (n_30064, n40412);
  and g67436 (n40413, n_30063, n_30064);
  not g67437 (n_30065, n40413);
  and g67438 (n40414, pi0212, n_30065);
  and g67439 (n40415, n_6791, n_30043);
  and g67440 (n40416, n_30048, n40415);
  not g67441 (n_30066, n40414);
  and g67442 (n40417, n_30066, n40416);
  not g67443 (n_30067, n40417);
  and g67444 (n40418, n40410, n_30067);
  not g67445 (n_30068, n40418);
  and g67446 (n40419, n40407, n_30068);
  and g67447 (n40420, n_30013, n40417);
  and g67448 (n40421, pi0219, n_30026);
  and g67449 (n40422, pi0214, n40386);
  not g67450 (n_30069, n40422);
  and g67451 (n40423, n_30062, n_30069);
  not g67452 (n_30070, n40423);
  and g67453 (n40424, pi0212, n_30070);
  and g67454 (n40425, n_26565, n40342);
  not g67455 (n_30071, n40425);
  and g67456 (n40426, n_26538, n_30071);
  and g67457 (n40427, n_30064, n40426);
  not g67458 (n_30072, n40424);
  not g67459 (n_30073, n40427);
  and g67460 (n40428, n_30072, n_30073);
  not g67461 (n_30074, n40428);
  and g67462 (n40429, n_6791, n_30074);
  not g67463 (n_30075, n40421);
  and g67464 (n40430, n_4226, n_30075);
  not g67465 (n_30076, n40429);
  and g67466 (n40431, n_30076, n40430);
  not g67467 (n_30077, n40420);
  and g67468 (n40432, n_30077, n40431);
  and g67469 (n40433, n_29810, n_29842);
  not g67470 (n_30078, n40432);
  and g67471 (n40434, n_30078, n40433);
  not g67472 (n_30079, n40419);
  and g67473 (n40435, n_29850, n_30079);
  not g67474 (n_30080, n40434);
  and g67475 (n40436, n_30080, n40435);
  not g67476 (n_30081, n40083);
  and g67477 (n40437, n_30081, n40415);
  not g67478 (n_30082, n40437);
  and g67479 (n40438, n40410, n_30082);
  and g67480 (n40439, pi1147, n_29815);
  not g67481 (n_30083, n40438);
  and g67482 (n40440, n_30083, n40439);
  and g67483 (n40441, n_29810, n_29807);
  not g67484 (n_30084, n40431);
  and g67485 (n40442, n_30084, n40441);
  not g67486 (n_30085, n40440);
  and g67487 (n40443, pi1149, n_30085);
  not g67488 (n_30086, n40442);
  and g67489 (n40444, n_30086, n40443);
  not g67490 (n_30087, n40444);
  and g67491 (n40445, pi1148, n_30087);
  not g67492 (n_30088, n40436);
  and g67493 (n40446, n_30088, n40445);
  and g67494 (n40447, n_29810, n_4226);
  and g67495 (n40448, n40342, n40447);
  and g67496 (n40449, pi0214, n_30043);
  and g67497 (n40450, n_30063, n40449);
  and g67498 (n40451, n_30044, n40387);
  not g67499 (n_30089, n40450);
  and g67500 (n40452, pi0212, n_30089);
  not g67501 (n_30090, n40451);
  and g67502 (n40453, n_30090, n40452);
  and g67503 (n40454, n_6791, n_30053);
  not g67504 (n_30091, n40453);
  and g67505 (n40455, n_30091, n40454);
  not g67506 (n_30092, n40455);
  and g67507 (n40456, n40418, n_30092);
  not g67508 (n_30093, n40456);
  and g67509 (n40457, n_29646, n_30093);
  not g67510 (n_30094, n40457);
  and g67511 (n40458, pi1147, n_30094);
  not g67512 (n_30095, n40448);
  not g67513 (n_30096, n40458);
  and g67514 (n40459, n_30095, n_30096);
  not g67515 (n_30097, n40459);
  and g67516 (n40460, n_29850, n_30097);
  and g67517 (n40461, n40410, n_30092);
  not g67518 (n_30098, n40461);
  and g67519 (n40462, n_29872, n_30098);
  not g67520 (n_30099, n40462);
  and g67521 (n40463, pi1147, n_30099);
  and g67522 (n40464, n_29810, n40207);
  not g67523 (n_30100, n40464);
  and g67524 (n40465, n_30095, n_30100);
  and g67525 (n40466, n16479, n40207);
  and g67526 (n40467, n40356, n40466);
  not g67527 (n_30101, n40465);
  not g67528 (n_30102, n40467);
  and g67529 (n40468, n_30101, n_30102);
  not g67530 (n_30103, n40463);
  not g67531 (n_30104, n40468);
  and g67532 (n40469, n_30103, n_30104);
  not g67533 (n_30105, n40469);
  and g67534 (n40470, pi1149, n_30105);
  not g67535 (n_30106, n40470);
  and g67536 (n40471, n_29904, n_30106);
  not g67537 (n_30107, n40460);
  and g67538 (n40472, n_30107, n40471);
  not g67539 (n_30108, n40446);
  and g67540 (n40473, pi0213, n_30108);
  not g67541 (n_30109, n40472);
  and g67542 (n40474, n_30109, n40473);
  not g67543 (n_30110, n40406);
  and g67544 (n40475, n_26372, n_30110);
  not g67545 (n_30111, n40474);
  and g67546 (n40476, n_30111, n40475);
  not g67547 (n_30112, n40329);
  not g67548 (n_30113, n40476);
  and g67549 (n40477, n_30112, n_30113);
  not g67550 (n_30114, n40477);
  and g67551 (n40478, pi0230, n_30114);
  and g67552 (n40479, n_28510, n_2307);
  not g67553 (n_30115, n40478);
  not g67554 (n_30116, n40479);
  and g67555 (po0397, n_30115, n_30116);
  not g67556 (n_30117, n39907);
  and g67557 (n40481, pi0213, n_30117);
  and g67558 (n40482, n39635, n39646);
  and g67559 (n40483, n38508, n39825);
  not g67560 (n_30118, n40483);
  and g67561 (n40484, n_29487, n_30118);
  not g67562 (n_30119, n40207);
  and g67563 (n40485, po1038, n_30119);
  not g67564 (n_30120, n40485);
  and g67565 (n40486, pi1151, n_30120);
  not g67566 (n_30121, n40484);
  and g67567 (n40487, n_30121, n40486);
  not g67568 (n_30122, n40482);
  not g67569 (n_30123, n40487);
  and g67570 (n40488, n_30122, n_30123);
  not g67571 (n_30124, n40488);
  and g67572 (n40489, n_28873, n_30124);
  and g67573 (n40490, n_29563, n40207);
  not g67574 (n_30125, n40490);
  and g67575 (n40491, n39872, n_30125);
  not g67576 (n_30126, n40491);
  and g67577 (n40492, pi1152, n_30126);
  not g67578 (n_30127, n40492);
  and g67579 (n40493, n_4226, n_30127);
  not g67580 (n_30128, n40493);
  and g67581 (n40494, n40486, n_30128);
  and g67582 (n40495, pi1152, n39635);
  and g67583 (n40496, n39737, n40495);
  not g67584 (n_30129, n40489);
  not g67585 (n_30130, n40496);
  and g67586 (n40497, n_30129, n_30130);
  not g67587 (n_30131, n40494);
  and g67588 (n40498, n_30131, n40497);
  not g67589 (n_30133, pi1150);
  not g67590 (n_30134, n40498);
  and g67591 (n40499, n_30133, n_30134);
  and g67592 (n40500, pi1151, n_29807);
  and g67593 (n40501, pi0219, n_29474);
  not g67594 (n_30135, n40501);
  and g67595 (n40502, n_4226, n_30135);
  not g67596 (n_30136, n40502);
  and g67597 (n40503, n_29847, n_30136);
  and g67598 (n40504, n39750, n_29658);
  not g67599 (n_30137, n40504);
  and g67600 (n40505, n_6791, n_30137);
  and g67601 (n40506, n_26565, n39755);
  not g67602 (n_30138, n40506);
  and g67603 (n40507, pi0212, n_30138);
  and g67604 (n40508, n_29649, n40507);
  not g67605 (n_30139, n40508);
  and g67606 (n40509, n40505, n_30139);
  not g67607 (n_30140, n40509);
  and g67608 (n40510, pi1152, n_30140);
  and g67609 (n40511, n_234, n_29508);
  and g67610 (n40512, n_26565, n39686);
  not g67611 (n_30141, n40512);
  and g67612 (n40513, pi0212, n_30141);
  and g67613 (n40514, n_29865, n40513);
  not g67614 (n_30142, n39664);
  not g67615 (n_30143, n40514);
  and g67616 (n40515, n_30142, n_30143);
  not g67617 (n_30144, n40511);
  not g67618 (n_30145, n40515);
  and g67619 (n40516, n_30144, n_30145);
  not g67620 (n_30146, n40516);
  and g67621 (n40517, n_6791, n_30146);
  and g67622 (n40518, n_28873, n_29954);
  not g67623 (n_30147, n40517);
  and g67624 (n40519, n_30147, n40518);
  not g67625 (n_30148, n40510);
  not g67626 (n_30149, n40519);
  and g67627 (n40520, n_30148, n_30149);
  not g67628 (n_30150, n40503);
  not g67629 (n_30151, n40520);
  and g67630 (n40521, n_30150, n_30151);
  not g67631 (n_30152, n40521);
  and g67632 (n40522, n40500, n_30152);
  and g67633 (n40523, n_29468, n_29842);
  and g67634 (n40524, n_26538, n_29470);
  and g67635 (n40525, n_29618, n40524);
  and g67636 (n40526, n_29634, n40525);
  not g67637 (n_30153, n40526);
  and g67638 (n40527, n_6791, n_30153);
  not g67639 (n_30154, n39638);
  and g67640 (n40528, pi0214, n_30154);
  and g67641 (n40529, n_7075, n39640);
  and g67642 (n40530, pi0212, n_29470);
  not g67643 (n_30155, n40529);
  and g67644 (n40531, n_30155, n40530);
  not g67645 (n_30156, n40528);
  and g67646 (n40532, n_30156, n40531);
  not g67647 (n_30157, n40532);
  and g67648 (n40533, n40527, n_30157);
  and g67649 (n40534, n_29474, n39834);
  and g67650 (n40535, n_234, n40534);
  not g67651 (n_30158, n40533);
  not g67652 (n_30159, n40535);
  and g67653 (n40536, n_30158, n_30159);
  and g67654 (n40537, n40502, n40536);
  not g67655 (n_30160, n40537);
  and g67656 (n40538, n_28873, n_30160);
  not g67657 (n_30161, n40536);
  and g67658 (n40539, n_29550, n_30161);
  not g67659 (n_30162, n40539);
  and g67660 (n40540, n39895, n_30162);
  not g67661 (n_30163, n40540);
  and g67662 (n40541, pi1152, n_30163);
  not g67663 (n_30164, n40538);
  not g67664 (n_30165, n40541);
  and g67665 (n40542, n_30164, n_30165);
  not g67666 (n_30166, n40542);
  and g67667 (n40543, n40523, n_30166);
  not g67668 (n_30167, n40543);
  and g67669 (n40544, pi1150, n_30167);
  not g67670 (n_30168, n40522);
  and g67671 (n40545, n_30168, n40544);
  not g67672 (n_30169, n40499);
  not g67673 (n_30170, n40545);
  and g67674 (n40546, n_30169, n_30170);
  not g67675 (n_30171, n40546);
  and g67676 (n40547, n_29850, n_30171);
  and g67677 (n40548, pi1151, n_29872);
  and g67678 (n40549, n_26565, n_29635);
  not g67679 (n_30172, n40549);
  and g67680 (n40550, n39849, n_30172);
  and g67681 (n40551, n_26538, n_29636);
  not g67682 (n_30173, n40550);
  not g67683 (n_30174, n40551);
  and g67684 (n40552, n_30173, n_30174);
  not g67685 (n_30175, n40552);
  and g67686 (n40553, n_6791, n_30175);
  and g67687 (n40554, n_28873, n39859);
  not g67688 (n_30176, n40553);
  and g67689 (n40555, n_30176, n40554);
  not g67690 (n_30177, n38783);
  and g67691 (n40556, n_30177, n_29563);
  and g67692 (n40557, pi0212, n39872);
  not g67693 (n_30178, n40556);
  and g67694 (n40558, n_30178, n40557);
  not g67695 (n_30179, n40558);
  and g67696 (n40559, n_29652, n_30179);
  not g67697 (n_30180, n40559);
  and g67698 (n40560, n_6791, n_30180);
  not g67699 (n_30181, n40560);
  and g67700 (n40561, pi1152, n_30181);
  and g67701 (n40562, n39879, n40561);
  not g67702 (n_30182, n40555);
  and g67703 (n40563, n40548, n_30182);
  not g67704 (n_30183, n40562);
  and g67705 (n40564, n_30183, n40563);
  and g67706 (n40565, n_29468, n_29646);
  and g67707 (n40566, n_29895, n_30136);
  not g67708 (n_30184, n40534);
  not g67709 (n_30185, n40566);
  and g67710 (n40567, n_30184, n_30185);
  and g67711 (n40568, n_28873, n40567);
  not g67712 (n_30186, n39895);
  and g67713 (n40569, n_30186, n40566);
  and g67714 (n40570, n_29550, n39834);
  not g67715 (n_30187, n40569);
  and g67716 (n40571, pi1152, n_30187);
  not g67717 (n_30188, n40570);
  and g67718 (n40572, n_30188, n40571);
  not g67719 (n_30189, n40568);
  and g67720 (n40573, n40565, n_30189);
  not g67721 (n_30190, n40572);
  and g67722 (n40574, n_30190, n40573);
  not g67723 (n_30191, n40574);
  and g67724 (n40575, n_30133, n_30191);
  not g67725 (n_30192, n40564);
  and g67726 (n40576, n_30192, n40575);
  and g67727 (n40577, n_29468, n_29848);
  and g67728 (n40578, n10843, n39724);
  and g67729 (n40579, n_29472, n_29619);
  and g67730 (n40580, n_7077, n_29550);
  not g67731 (n_30193, n40579);
  and g67732 (n40581, n_30193, n40580);
  not g67733 (n_30194, n40578);
  not g67734 (n_30195, n40581);
  and g67735 (n40582, n_30194, n_30195);
  not g67736 (n_30196, n40582);
  and g67737 (n40583, n_6791, n_30196);
  not g67738 (n_30197, n40583);
  and g67739 (n40584, n_30187, n_30197);
  not g67740 (n_30198, n40584);
  and g67741 (n40585, pi1152, n_30198);
  not g67742 (n_30199, n40567);
  and g67743 (n40586, n40538, n_30199);
  not g67744 (n_30200, n40585);
  not g67745 (n_30201, n40586);
  and g67746 (n40587, n_30200, n_30201);
  not g67747 (n_30202, n40587);
  and g67748 (n40588, n40577, n_30202);
  and g67749 (n40589, pi0212, n_29563);
  not g67750 (n_30203, n40589);
  and g67751 (n40590, n40505, n_30203);
  not g67752 (n_30204, n40590);
  and g67753 (n40591, pi1152, n_30204);
  and g67754 (n40592, n39879, n40591);
  and g67755 (n40593, pi1151, n_29815);
  and g67756 (n40594, n_29517, n_30144);
  not g67757 (n_30205, n40594);
  and g67758 (n40595, n_6791, n_30205);
  not g67759 (n_30206, n40595);
  and g67760 (n40596, n40554, n_30206);
  not g67761 (n_30207, n40596);
  and g67762 (n40597, n40593, n_30207);
  not g67763 (n_30208, n40592);
  and g67764 (n40598, n_30208, n40597);
  not g67765 (n_30209, n40588);
  and g67766 (n40599, pi1150, n_30209);
  not g67767 (n_30210, n40598);
  and g67768 (n40600, n_30210, n40599);
  not g67769 (n_30211, n40576);
  not g67770 (n_30212, n40600);
  and g67771 (n40601, n_30211, n_30212);
  not g67772 (n_30213, n40601);
  and g67773 (n40602, pi1149, n_30213);
  not g67774 (n_30214, n40547);
  not g67775 (n_30215, n40602);
  and g67776 (n40603, n_30214, n_30215);
  not g67777 (n_30216, n40603);
  and g67778 (n40604, n_26557, n_30216);
  not g67779 (n_30217, n40481);
  and g67780 (n40605, pi0209, n_30217);
  not g67781 (n_30218, n40604);
  and g67782 (n40606, n_30218, n40605);
  and g67783 (n40607, n_30133, pi1151);
  not g67784 (n_30219, n40143);
  and g67785 (n40608, n_30219, n40607);
  and g67786 (n40609, n_29843, n40523);
  and g67787 (n40610, n_29808, n40500);
  not g67788 (n_30220, n40610);
  and g67789 (n40611, pi1150, n_30220);
  not g67790 (n_30221, n40609);
  and g67791 (n40612, n_30221, n40611);
  not g67792 (n_30222, n40608);
  and g67793 (n40613, n_29850, n_30222);
  not g67794 (n_30223, n40612);
  and g67795 (n40614, n_30223, n40613);
  and g67796 (n40615, n40088, n40593);
  and g67797 (n40616, n_29468, n40134);
  not g67798 (n_30224, n40615);
  and g67799 (n40617, pi1150, n_30224);
  not g67800 (n_30225, n40616);
  and g67801 (n40618, n_30225, n40617);
  and g67802 (n40619, n_29900, n40565);
  and g67803 (n40620, n_29873, n40548);
  not g67804 (n_30226, n40619);
  and g67805 (n40621, n_30133, n_30226);
  not g67806 (n_30227, n40620);
  and g67807 (n40622, n_30227, n40621);
  not g67808 (n_30228, n40618);
  and g67809 (n40623, pi1149, n_30228);
  not g67810 (n_30229, n40622);
  and g67811 (n40624, n_30229, n40623);
  not g67812 (n_30230, n40614);
  not g67813 (n_30231, n40624);
  and g67814 (n40625, n_30230, n_30231);
  and g67815 (n40626, n_26557, n40625);
  not g67816 (n_30232, n40153);
  not g67817 (n_30233, n40157);
  and g67818 (n40627, n_30232, n_30233);
  and g67819 (n40628, n_28774, n39695);
  not g67820 (n_30234, n40628);
  and g67821 (n40629, n_29515, n_30234);
  and g67822 (n40630, n_29868, n40629);
  not g67823 (n_30235, n40627);
  not g67824 (n_30236, n40630);
  and g67825 (n40631, n_30235, n_30236);
  not g67826 (n_30237, n40631);
  and g67827 (n40632, n_6791, n_30237);
  not g67828 (n_30238, n40632);
  and g67829 (n40633, n40164, n_30238);
  not g67830 (n_30239, n40633);
  and g67831 (n40634, n39845, n_30239);
  and g67832 (n40635, pi0299, n39631);
  and g67833 (n40636, n_29886, n_30118);
  not g67834 (n_30240, n40636);
  and g67835 (n40637, n_4226, n_30240);
  not g67836 (n_30241, n40635);
  and g67837 (n40638, n_30241, n40637);
  not g67838 (n_30242, n40638);
  and g67839 (n40639, n39828, n_30242);
  not g67840 (n_30243, n40639);
  and g67841 (n40640, n_28873, n_30243);
  not g67842 (n_30244, n40634);
  and g67843 (n40641, n_30244, n40640);
  and g67844 (n40642, n_29863, n_29864);
  not g67847 (n_30245, n40642);
  not g67849 (n_30246, n40645);
  and g67850 (n40646, n40164, n_30246);
  not g67851 (n_30247, n40646);
  and g67852 (n40647, n39871, n_30247);
  and g67853 (n40648, n_30081, n_29886);
  and g67854 (n40649, n_29326, n39867);
  not g67855 (n_30248, n40648);
  not g67856 (n_30249, n40649);
  and g67857 (n40650, n_30248, n_30249);
  not g67858 (n_30250, n40650);
  and g67859 (n40651, n_6791, n_30250);
  and g67860 (n40652, pi0219, n_29886);
  not g67861 (n_30251, n40652);
  and g67862 (n40653, n_4226, n_30251);
  not g67863 (n_30252, n40651);
  and g67864 (n40654, n_30252, n40653);
  not g67865 (n_30253, n40654);
  and g67866 (n40655, n39893, n_30253);
  not g67867 (n_30254, n40655);
  and g67868 (n40656, pi1152, n_30254);
  not g67869 (n_30255, n40647);
  and g67870 (n40657, n_30255, n40656);
  not g67871 (n_30256, n40657);
  and g67872 (n40658, n_30133, n_30256);
  not g67873 (n_30257, n40641);
  and g67874 (n40659, n_30257, n40658);
  and g67875 (n40660, n_6791, n_29971);
  and g67876 (n40661, n_29977, n40660);
  and g67877 (n40662, n_11757, n40661);
  and g67878 (n40663, pi0299, n10485);
  not g67879 (n_30258, n40663);
  and g67880 (n40664, n_6791, n_30258);
  not g67881 (n_30259, n40664);
  and g67882 (n40665, n40195, n_30259);
  not g67883 (n_30260, n40665);
  and g67884 (n40666, n_29981, n_30260);
  not g67885 (n_30261, n40662);
  not g67886 (n_30262, n40666);
  and g67887 (n40667, n_30261, n_30262);
  not g67888 (n_30263, n40667);
  and g67889 (n40668, n39845, n_30263);
  and g67890 (n40669, pi1153, n40483);
  not g67891 (n_30264, n40669);
  and g67892 (n40670, n39828, n_30264);
  not g67893 (n_30265, n40670);
  and g67894 (n40671, n_28873, n_30265);
  and g67895 (n40672, n_29468, n_29847);
  not g67896 (n_30266, n40672);
  and g67897 (n40673, n_28873, n_30266);
  not g67898 (n_30267, n40671);
  not g67899 (n_30268, n40673);
  and g67900 (n40674, n_30267, n_30268);
  not g67901 (n_30269, n40668);
  not g67902 (n_30270, n40674);
  and g67903 (n40675, n_30269, n_30270);
  and g67904 (n40676, n_7075, n40661);
  not g67905 (n_30271, n40088);
  not g67906 (n_30272, n40676);
  and g67907 (n40677, n_30271, n_30272);
  not g67908 (n_30273, n40677);
  and g67909 (n40678, n39871, n_30273);
  and g67910 (n40679, n_30263, n40678);
  not g67911 (n_30274, n39768);
  and g67912 (n40680, n_4226, n_30274);
  and g67913 (n40681, n10843, n_29877);
  and g67914 (n40682, n_234, n39747);
  and g67915 (n40683, n_28519, n_30241);
  not g67916 (n_30275, n40682);
  and g67917 (n40684, n_30275, n40683);
  not g67918 (n_30276, n40681);
  and g67919 (n40685, n40230, n_30276);
  not g67920 (n_30277, n40684);
  and g67921 (n40686, n_30277, n40685);
  not g67922 (n_30278, n40686);
  and g67923 (n40687, n40680, n_30278);
  not g67924 (n_30279, n40687);
  and g67925 (n40688, n39893, n_30279);
  not g67926 (n_30280, n40688);
  and g67927 (n40689, pi1152, n_30280);
  not g67928 (n_30281, n40679);
  and g67929 (n40690, n_30281, n40689);
  not g67930 (n_30282, n40675);
  and g67931 (n40691, pi1150, n_30282);
  not g67932 (n_30283, n40690);
  and g67933 (n40692, n_30283, n40691);
  not g67934 (n_30284, n40692);
  and g67935 (n40693, pi1149, n_30284);
  not g67936 (n_30285, n40659);
  and g67937 (n40694, n_30285, n40693);
  not g67938 (n_30286, n39642);
  and g67939 (n40695, pi0219, n_30286);
  not g67940 (n_30287, n40695);
  and g67941 (n40696, n_4226, n_30287);
  and g67942 (n40697, n_29623, n40696);
  not g67943 (n_30288, n40697);
  and g67944 (n40698, n39845, n_30288);
  not g67945 (n_30289, n40698);
  and g67946 (n40699, n40671, n_30289);
  and g67947 (n40700, pi0299, n39864);
  and g67948 (n40701, n_29645, n40700);
  not g67949 (n_30290, n40701);
  and g67950 (n40702, n39893, n_30290);
  not g67951 (n_30291, n40531);
  and g67952 (n40703, n40527, n_30291);
  not g67953 (n_30292, n40703);
  and g67954 (n40704, n40696, n_30292);
  and g67955 (n40705, n39871, n_30288);
  not g67956 (n_30293, n40704);
  and g67957 (n40706, n_30293, n40705);
  not g67958 (n_30294, n40702);
  and g67959 (n40707, pi1152, n_30294);
  not g67960 (n_30295, n40706);
  and g67961 (n40708, n_30295, n40707);
  not g67962 (n_30296, n40699);
  and g67963 (n40709, n_30133, n_30296);
  not g67964 (n_30297, n40708);
  and g67965 (n40710, n_30297, n40709);
  and g67966 (n40711, n_29675, n40100);
  and g67967 (n40712, n_28774, n_29829);
  not g67968 (n_30298, n40712);
  and g67969 (n40713, n_7075, n_30298);
  and g67970 (n40714, n39909, n_29833);
  not g67971 (n_30299, n40713);
  and g67972 (n40715, n_30299, n40714);
  not g67973 (n_30300, n40711);
  not g67974 (n_30301, n40715);
  and g67975 (n40716, n_30300, n_30301);
  not g67976 (n_30302, n40716);
  and g67977 (n40717, n_4226, n_30302);
  not g67978 (n_30303, n40717);
  and g67979 (n40718, n39828, n_30303);
  and g67980 (n40719, pi0211, n_29800);
  and g67981 (n40720, n_28639, n38675);
  not g67982 (n_30304, n40720);
  and g67983 (n40721, n_29797, n_30304);
  and g67984 (n40722, n_7075, n_28774);
  not g67985 (n_30305, n40721);
  and g67986 (n40723, n_30305, n40722);
  not g67987 (n_30306, n40719);
  not g67988 (n_30307, n40723);
  and g67989 (n40724, n_30306, n_30307);
  and g67990 (n40725, n_29794, n_30306);
  and g67991 (n40726, pi0214, n40725);
  and g67992 (n40727, n40062, n_29802);
  not g67993 (n_30308, n40727);
  and g67994 (n40728, pi0212, n_30308);
  not g67995 (n_30309, n40726);
  and g67996 (n40729, n_30309, n40728);
  not g67997 (n_30310, n40724);
  and g67998 (n40730, n_30310, n40729);
  and g67999 (n40731, n_29801, n_30307);
  not g68000 (n_30311, n40731);
  and g68001 (n40732, n40063, n_30311);
  not g68002 (n_30312, n40732);
  and g68003 (n40733, n_6791, n_30312);
  not g68004 (n_30313, n40730);
  and g68005 (n40734, n_30313, n40733);
  not g68006 (n_30314, n40734);
  and g68007 (n40735, n40310, n_30314);
  not g68008 (n_30315, n40735);
  and g68009 (n40736, n39845, n_30315);
  not g68010 (n_30316, n40718);
  and g68011 (n40737, n_28873, n_30316);
  not g68012 (n_30317, n40736);
  and g68013 (n40738, n_30317, n40737);
  and g68014 (n40739, pi0214, n40724);
  not g68015 (n_30318, n40739);
  and g68016 (n40740, n40063, n_30318);
  and g68017 (n40741, n_26565, n40724);
  not g68018 (n_30319, n40741);
  and g68019 (n40742, n40315, n_30319);
  not g68020 (n_30320, n40740);
  and g68021 (n40743, n_6791, n_30320);
  not g68022 (n_30321, n40742);
  and g68023 (n40744, n_30321, n40743);
  not g68024 (n_30322, n40744);
  and g68025 (n40745, n40310, n_30322);
  not g68026 (n_30323, n40745);
  and g68027 (n40746, n39871, n_30323);
  and g68028 (n40747, n_29829, n_30241);
  and g68029 (n40748, pi0214, n40747);
  not g68030 (n_30324, n40748);
  and g68031 (n40749, n40108, n_30324);
  and g68032 (n40750, n_26565, n40747);
  not g68033 (n_30325, n40750);
  and g68034 (n40751, n40113, n_30325);
  not g68035 (n_30326, n40749);
  not g68036 (n_30327, n40751);
  and g68037 (n40752, n_30326, n_30327);
  not g68038 (n_30328, n40752);
  and g68039 (n40753, n_6791, n_30328);
  not g68040 (n_30329, n40753);
  and g68041 (n40754, n40123, n_30329);
  not g68042 (n_30330, n40754);
  and g68043 (n40755, n39893, n_30330);
  not g68044 (n_30331, n40746);
  and g68045 (n40756, pi1152, n_30331);
  not g68046 (n_30332, n40755);
  and g68047 (n40757, n_30332, n40756);
  not g68048 (n_30333, n40738);
  and g68049 (n40758, pi1150, n_30333);
  not g68050 (n_30334, n40757);
  and g68051 (n40759, n_30334, n40758);
  not g68052 (n_30335, n40710);
  and g68053 (n40760, n_29850, n_30335);
  not g68054 (n_30336, n40759);
  and g68055 (n40761, n_30336, n40760);
  not g68056 (n_30337, n40694);
  not g68057 (n_30338, n40761);
  and g68058 (n40762, n_30337, n_30338);
  not g68059 (n_30339, n40762);
  and g68060 (n40763, pi0213, n_30339);
  not g68061 (n_30340, n40626);
  and g68062 (n40764, n_26372, n_30340);
  not g68063 (n_30341, n40763);
  and g68064 (n40765, n_30341, n40764);
  not g68065 (n_30342, n40606);
  not g68066 (n_30343, n40765);
  and g68067 (n40766, n_30342, n_30343);
  not g68068 (n_30344, n40766);
  and g68069 (n40767, pi0230, n_30344);
  and g68070 (n40768, n_28510, n_1595);
  not g68071 (n_30345, n40767);
  not g68072 (n_30346, n40768);
  and g68073 (po0398, n_30345, n_30346);
  and g68074 (n40770, n_28510, n_2915);
  and g68075 (n40771, pi0219, n_28515);
  not g68076 (n_30347, n39414);
  and g68077 (n40772, pi0214, n_30347);
  and g68078 (n40773, n_26565, n_29911);
  not g68079 (n_30348, n40772);
  not g68080 (n_30349, n40773);
  and g68081 (n40774, n_30348, n_30349);
  not g68082 (n_30350, n40774);
  and g68083 (n40775, pi0212, n_30350);
  and g68084 (n40776, n_26538, n40212);
  not g68085 (n_30351, n40776);
  and g68086 (n40777, n_6791, n_30351);
  not g68087 (n_30352, n40775);
  and g68088 (n40778, n_30352, n40777);
  not g68089 (n_30353, n40771);
  and g68090 (n40779, n38416, n_30353);
  not g68091 (n_30354, n40778);
  and g68092 (n40780, n_30354, n40779);
  and g68093 (n40781, pi0199, pi1144);
  not g68094 (n_30355, n40781);
  and g68095 (n40782, n_7045, n_30355);
  and g68096 (n40783, n_30004, n40782);
  and g68097 (n40784, n_234, n_30005);
  not g68098 (n_30356, n40783);
  and g68099 (n40785, n_30356, n40784);
  and g68100 (n40786, n38826, n40785);
  not g68101 (n_30357, n40785);
  and g68102 (n40787, n_25873, n_30357);
  and g68103 (n40788, n_234, n_29279);
  and g68104 (n40789, n_29278, n40782);
  not g68105 (n_30358, n40789);
  and g68106 (n40790, n40788, n_30358);
  not g68107 (n_30359, n40790);
  and g68108 (n40791, pi0207, n_30359);
  not g68109 (n_30360, n40787);
  and g68110 (n40792, pi0208, n_30360);
  not g68111 (n_30361, n40791);
  and g68112 (n40793, n_30361, n40792);
  not g68113 (n_30362, n40786);
  not g68114 (n_30363, n40793);
  and g68115 (n40794, n_30362, n_30363);
  and g68116 (n40795, n_26565, n40794);
  not g68117 (n_30364, n40795);
  and g68118 (n40796, n_26538, n_30364);
  and g68119 (n40797, n38449, n40785);
  not g68120 (n_30365, n40797);
  and g68121 (n40798, n_29958, n_30365);
  and g68122 (n40799, n_30363, n40798);
  not g68123 (n_30366, n40799);
  and g68124 (n40800, n_7075, n_30366);
  and g68125 (n40801, n_29346, n_30365);
  and g68126 (n40802, n_30363, n40801);
  not g68127 (n_30367, n40802);
  and g68128 (n40803, pi0211, n_30367);
  not g68129 (n_30368, n40800);
  not g68130 (n_30369, n40803);
  and g68131 (n40804, n_30368, n_30369);
  and g68132 (n40805, pi0214, n40804);
  not g68133 (n_30370, n40805);
  and g68134 (n40806, n40796, n_30370);
  and g68135 (n40807, n_7075, n_30367);
  and g68136 (n40808, n_28654, n_30365);
  and g68137 (n40809, n_30363, n40808);
  not g68138 (n_30371, n40809);
  and g68139 (n40810, pi0211, n_30371);
  not g68140 (n_30372, n40807);
  and g68141 (n40811, pi0214, n_30372);
  not g68142 (n_30373, n40810);
  and g68143 (n40812, n_30373, n40811);
  and g68144 (n40813, n_26565, n40804);
  not g68145 (n_30374, n40812);
  and g68146 (n40814, pi0212, n_30374);
  not g68147 (n_30375, n40813);
  and g68148 (n40815, n_30375, n40814);
  not g68149 (n_30376, n40806);
  and g68150 (n40816, n_6791, n_30376);
  not g68151 (n_30377, n40815);
  and g68152 (n40817, n_30377, n40816);
  not g68153 (n_30378, n40794);
  and g68154 (n40818, n_28512, n_30378);
  not g68155 (n_30379, n40818);
  and g68156 (n40819, pi0219, n_30379);
  and g68157 (n40820, n38414, n_30371);
  not g68158 (n_30380, n40820);
  and g68159 (n40821, n40819, n_30380);
  not g68160 (n_30381, n40821);
  and g68161 (n40822, n_4226, n_30381);
  not g68162 (n_30382, n40817);
  and g68163 (n40823, n_30382, n40822);
  not g68164 (n_30383, n40780);
  not g68165 (n_30384, n40823);
  and g68166 (n40824, n_30383, n_30384);
  and g68167 (n40825, pi0213, n40824);
  and g68168 (n40826, n38413, n_30362);
  and g68169 (n40827, pi0211, n_30362);
  and g68170 (n40828, n38414, n_28720);
  and g68171 (n40829, n_30365, n40828);
  not g68172 (n_30385, n40827);
  not g68173 (n_30386, n40829);
  and g68174 (n40830, n_30385, n_30386);
  not g68175 (n_30387, n40830);
  and g68176 (n40831, pi0219, n_30387);
  and g68177 (n40832, n10843, n_28547);
  and g68178 (n40833, n_28543, n38608);
  not g68179 (n_30388, n40832);
  not g68180 (n_30389, n40833);
  and g68181 (n40834, n_30388, n_30389);
  and g68182 (n40835, n_6791, n_30365);
  not g68183 (n_30390, n40834);
  and g68184 (n40836, n_30390, n40835);
  not g68185 (n_30391, n40826);
  not g68186 (n_30392, n40836);
  and g68187 (n40837, n_30391, n_30392);
  not g68188 (n_30393, n40831);
  and g68189 (n40838, n_30393, n40837);
  not g68190 (n_30394, n40838);
  and g68191 (n40839, n_30363, n_30394);
  not g68192 (n_30395, n40839);
  and g68193 (n40840, n_4226, n_30395);
  and g68194 (n40841, n_26557, n_28560);
  not g68195 (n_30396, n40840);
  and g68196 (n40842, n_30396, n40841);
  not g68197 (n_30397, n40825);
  not g68198 (n_30398, n40842);
  and g68199 (n40843, n_30397, n_30398);
  not g68200 (n_30399, n40843);
  and g68201 (n40844, pi0209, n_30399);
  not g68202 (n_30400, n38476);
  and g68203 (n40845, n_26557, n_30400);
  and g68204 (n40846, pi0219, n38413);
  not g68205 (n_30401, n40846);
  and g68206 (n40847, n_30353, n_30401);
  and g68207 (n40848, n_30354, n40847);
  not g68208 (n_30402, n40848);
  and g68209 (n40849, pi0299, n_30402);
  not g68210 (n_30403, n40849);
  and g68211 (n40850, n_4226, n_30403);
  and g68212 (n40851, n_28555, n40850);
  not g68213 (n_30404, n40851);
  and g68214 (n40852, n_30383, n_30404);
  not g68215 (n_30405, n40852);
  and g68216 (n40853, pi0213, n_30405);
  not g68217 (n_30406, n40853);
  and g68218 (n40854, n_26372, n_30406);
  not g68219 (n_30407, n40845);
  and g68220 (n40855, n_30407, n40854);
  not g68221 (n_30408, n40844);
  not g68222 (n_30409, n40855);
  and g68223 (n40856, n_30408, n_30409);
  not g68224 (n_30410, n40856);
  and g68225 (n40857, pi0230, n_30410);
  not g68226 (n_30411, n40770);
  not g68227 (n_30412, n40857);
  and g68228 (po0399, n_30411, n_30412);
  and g68229 (n40859, pi0253, pi0254);
  and g68230 (n40860, pi0267, n40859);
  not g68231 (n_30417, pi0263);
  and g68232 (n40861, n_30417, n40860);
  and g68233 (n40862, n_60, n_76);
  not g68234 (n_30418, n40862);
  and g68235 (n40863, pi0314, n_30418);
  and g68236 (n40864, pi0802, n40863);
  and g68237 (n40865, pi0276, n40864);
  and g68238 (n40866, n_3128, n40865);
  and g68239 (n40867, pi0271, n40866);
  and g68240 (n40868, pi0273, n40867);
  and g68241 (n40869, pi0243, n40868);
  not g68242 (n_30423, n40865);
  and g68243 (n40870, n_3128, n_30423);
  not g68244 (n_30424, n40870);
  and g68245 (n40871, pi0271, n_30424);
  not g68246 (n_30425, n40871);
  and g68247 (n40872, n_3128, n_30425);
  not g68248 (n_30426, n40872);
  and g68249 (n40873, pi0273, n_30426);
  not g68250 (n_30427, n40873);
  and g68251 (n40874, n_3128, n_30427);
  not g68252 (n_30428, pi0243);
  and g68253 (n40875, n_30428, n40874);
  and g68254 (n40876, pi0243, n_3128);
  not g68255 (n_30429, n40876);
  and g68256 (n40877, n38478, n_30429);
  not g68257 (n_30430, n40866);
  and g68258 (n40878, n_30430, n40877);
  not g68259 (n_30431, n40869);
  not g68260 (n_30432, n40878);
  and g68261 (n40879, n_30431, n_30432);
  not g68262 (n_30433, n40875);
  and g68263 (n40880, n_30433, n40879);
  not g68264 (n_30434, n40880);
  and g68265 (n40881, pi0219, n_30434);
  and g68266 (n40882, n_28563, n_28569);
  and g68267 (n40883, pi1091, n40882);
  and g68268 (n40884, n_105, n40862);
  not g68269 (n_30435, n40884);
  and g68270 (n40885, pi0314, n_30435);
  and g68271 (n40886, pi0802, n40885);
  and g68272 (n40887, pi0276, n40886);
  and g68273 (n40888, n_3128, n40887);
  and g68274 (n40889, pi0271, n40888);
  and g68275 (n40890, pi0273, n40889);
  not g68276 (n_30436, n40890);
  and g68277 (n40891, n_30427, n_30436);
  and g68278 (n40892, n40876, n40891);
  and g68279 (n40893, n_30428, n40890);
  not g68286 (n_30440, n40881);
  not g68287 (n_30441, n40896);
  and g68288 (n40897, n_30440, n_30441);
  not g68289 (n_30442, n40897);
  and g68290 (n40898, n40861, n_30442);
  and g68291 (n40899, n_30428, n_3128);
  not g68292 (n_30443, n40882);
  and g68293 (n40900, n_6791, n_30443);
  and g68294 (n40901, pi1157, n38519);
  not g68295 (n_30444, n40900);
  not g68296 (n_30445, n40901);
  and g68297 (n40902, n_30444, n_30445);
  not g68298 (n_30446, n40902);
  and g68299 (n40903, pi1091, n_30446);
  not g68300 (n_30447, n40899);
  not g68301 (n_30448, n40903);
  and g68302 (n40904, n_30447, n_30448);
  not g68303 (n_30449, n40861);
  not g68304 (n_30450, n40904);
  and g68305 (n40905, n_30449, n_30450);
  not g68306 (n_30451, n40905);
  and g68307 (n40906, po1038, n_30451);
  not g68308 (n_30452, n40898);
  and g68309 (n40907, n_30452, n40906);
  and g68310 (n40908, pi0272, pi0283);
  and g68311 (n40909, pi0275, n40908);
  and g68312 (n40910, pi0268, n40909);
  and g68313 (n40911, n_234, pi1091);
  and g68314 (n40912, n38841, n40911);
  not g68315 (n_30457, n40912);
  and g68316 (n40913, n_30447, n_30457);
  not g68317 (n_30458, n40913);
  and g68318 (n40914, pi1156, n_30458);
  and g68319 (n40915, pi1091, n_28928);
  and g68320 (n40916, n39457, n40915);
  not g68321 (n_30459, n40914);
  not g68322 (n_30460, n40916);
  and g68323 (n40917, n_30459, n_30460);
  and g68324 (n40918, n_234, n38699);
  not g68325 (n_30461, n40918);
  and g68326 (n40919, pi1091, n_30461);
  not g68327 (n_30462, n40919);
  and g68328 (n40920, n_30429, n_30462);
  and g68329 (n40921, n_11768, n_30447);
  not g68330 (n_30463, n40921);
  and g68331 (n40922, n_30429, n_30463);
  and g68332 (n40923, n38568, n40922);
  not g68333 (n_30464, n40920);
  not g68334 (n_30465, n40923);
  and g68335 (n40924, n_30464, n_30465);
  not g68336 (n_30466, n40924);
  and g68337 (n40925, n_11794, n_30466);
  not g68338 (n_30467, n40925);
  and g68339 (n40926, n40917, n_30467);
  not g68340 (n_30468, n40926);
  and g68341 (n40927, pi1157, n_30468);
  not g68342 (n_30469, n40915);
  and g68343 (n40928, n_30469, n40922);
  not g68344 (n_30470, n40928);
  and g68345 (n40929, n_11794, n_30470);
  and g68346 (n40930, pi1155, n_30429);
  and g68347 (n40931, pi0199, pi1091);
  and g68348 (n40932, n_234, n40931);
  not g68349 (n_30471, n40932);
  and g68350 (n40933, n40930, n_30471);
  not g68351 (n_30472, n40933);
  and g68352 (n40934, pi1156, n_30472);
  and g68353 (n40935, n_11768, n_30429);
  and g68354 (n40936, n_28601, n40911);
  not g68355 (n_30473, n40936);
  and g68356 (n40937, n40935, n_30473);
  not g68357 (n_30474, n40937);
  and g68358 (n40938, n40934, n_30474);
  not g68359 (n_30475, n40929);
  and g68360 (n40939, n_11810, n_30475);
  not g68361 (n_30476, n40938);
  and g68362 (n40940, n_30476, n40939);
  not g68363 (n_30477, n40927);
  not g68364 (n_30478, n40940);
  and g68365 (n40941, n_30477, n_30478);
  not g68366 (n_30479, n40941);
  and g68367 (n40942, pi0211, n_30479);
  and g68368 (n40943, pi1091, n_7409);
  not g68369 (n_30480, n40943);
  and g68370 (n40944, n40935, n_30480);
  not g68371 (n_30481, n40944);
  and g68372 (n40945, n_30472, n_30481);
  and g68373 (n40946, pi0200, n_11794);
  and g68374 (n40947, n40911, n40946);
  not g68375 (n_30482, n40945);
  not g68376 (n_30483, n40947);
  and g68377 (n40948, n_30482, n_30483);
  not g68378 (n_30484, n40948);
  and g68379 (n40949, n_11810, n_30484);
  and g68380 (n40950, n40913, n40934);
  and g68381 (n40951, pi0200, pi1091);
  and g68382 (n40952, n_234, n40951);
  not g68383 (n_30485, n40952);
  and g68384 (n40953, n40930, n_30485);
  and g68385 (n40954, n_11768, n40920);
  not g68386 (n_30486, n40953);
  and g68387 (n40955, n_11794, n_30486);
  not g68388 (n_30487, n40954);
  and g68389 (n40956, n_30487, n40955);
  not g68390 (n_30488, n40950);
  not g68391 (n_30489, n40956);
  and g68392 (n40957, n_30488, n_30489);
  not g68393 (n_30490, n40957);
  and g68394 (n40958, pi1157, n_30490);
  not g68395 (n_30491, n40949);
  and g68396 (n40959, n_7075, n_30491);
  not g68397 (n_30492, n40958);
  and g68398 (n40960, n_30492, n40959);
  not g68399 (n_30493, n40942);
  not g68400 (n_30494, n40960);
  and g68401 (n40961, n_30493, n_30494);
  not g68402 (n_30495, n40961);
  and g68403 (n40962, n_6791, n_30495);
  and g68404 (n40963, n39369, n_30459);
  and g68405 (n40964, n_30467, n40963);
  and g68406 (n40965, pi0299, pi1091);
  not g68407 (n_30496, n40965);
  and g68408 (n40966, n40948, n_30496);
  not g68409 (n_30497, n40966);
  and g68410 (n40967, n_11810, n_30497);
  and g68411 (n40968, pi1091, n38700);
  not g68412 (n_30498, n40968);
  and g68413 (n40969, n40935, n_30498);
  not g68414 (n_30499, n40969);
  and g68415 (n40970, n_30486, n_30499);
  not g68416 (n_30500, n40970);
  and g68417 (n40971, n_11794, n_30500);
  not g68418 (n_30501, n40971);
  and g68419 (n40972, n38478, n_30501);
  and g68420 (n40973, n40917, n40972);
  not g68427 (n_30505, n40962);
  not g68428 (n_30506, n40976);
  and g68429 (n40977, n_30505, n_30506);
  not g68430 (n_30507, n40977);
  and g68431 (n40978, n_30449, n_30507);
  not g68432 (n_30508, n40874);
  and g68433 (n40979, pi0199, n_30508);
  and g68434 (n40980, n_3128, n40891);
  not g68435 (n_30509, n40980);
  and g68436 (n40981, n_7044, n_30509);
  not g68437 (n_30510, n40979);
  not g68438 (n_30511, n40981);
  and g68439 (n40982, n_30510, n_30511);
  not g68440 (n_30512, n40888);
  and g68441 (n40983, n_7045, n_30512);
  not g68442 (n_30513, n40982);
  not g68443 (n_30514, n40983);
  and g68444 (n40984, n_30513, n_30514);
  not g68445 (n_30515, n40984);
  and g68446 (n40985, n_234, n_30515);
  and g68447 (n40986, pi0299, n40874);
  and g68448 (n40987, n_30436, n40986);
  not g68449 (n_30516, n40985);
  not g68450 (n_30517, n40987);
  and g68451 (n40988, n_30516, n_30517);
  not g68452 (n_30518, n40988);
  and g68453 (n40989, n_30428, n_30518);
  and g68454 (n40990, n_7045, n_30508);
  and g68455 (n40991, n40888, n_30513);
  not g68456 (n_30519, n40991);
  and g68457 (n40992, n_234, n_30519);
  not g68458 (n_30520, n40990);
  and g68459 (n40993, n_30520, n40992);
  not g68460 (n_30521, n40868);
  and g68461 (n40994, pi0299, n_30521);
  not g68462 (n_30522, n40993);
  not g68463 (n_30523, n40994);
  and g68464 (n40995, n_30522, n_30523);
  and g68465 (n40996, pi0243, n40995);
  not g68466 (n_30524, n40989);
  not g68467 (n_30525, n40996);
  and g68468 (n40997, n_30524, n_30525);
  not g68469 (n_30526, n40997);
  and g68470 (n40998, pi1155, n_30526);
  and g68471 (n40999, n_30511, n40985);
  not g68472 (n_30527, n40986);
  not g68473 (n_30528, n40999);
  and g68474 (n41000, n_30527, n_30528);
  not g68475 (n_30529, n41000);
  and g68476 (n41001, n_30428, n_30529);
  and g68477 (n41002, n_30510, n40992);
  not g68478 (n_30530, n41002);
  and g68479 (n41003, n40995, n_30530);
  and g68480 (n41004, pi0243, n41003);
  not g68481 (n_30531, n41001);
  not g68482 (n_30532, n41004);
  and g68483 (n41005, n_30531, n_30532);
  not g68484 (n_30533, n40998);
  and g68485 (n41006, n_30533, n41005);
  not g68486 (n_30534, n41006);
  and g68487 (n41007, n_11794, n_30534);
  and g68488 (n41008, n_30520, n41002);
  not g68489 (n_30535, n41008);
  and g68490 (n41009, n_30527, n_30535);
  and g68491 (n41010, n_30428, n41009);
  and g68492 (n41011, n_30510, n40985);
  and g68493 (n41012, n_30511, n40993);
  not g68494 (n_30536, n41012);
  and g68495 (n41013, n_30523, n_30536);
  not g68496 (n_30537, n41011);
  and g68497 (n41014, n_30537, n41013);
  not g68498 (n_30538, n41014);
  and g68499 (n41015, pi0243, n_30538);
  not g68500 (n_30539, n41010);
  not g68501 (n_30540, n41015);
  and g68502 (n41016, n_30539, n_30540);
  and g68503 (n41017, n_11768, n_30531);
  and g68504 (n41018, pi1155, n_30524);
  and g68505 (n41019, pi0243, n41013);
  not g68506 (n_30541, n41019);
  and g68507 (n41020, n41018, n_30541);
  not g68508 (n_30542, n41017);
  not g68509 (n_30543, n41020);
  and g68510 (n41021, n_30542, n_30543);
  not g68511 (n_30544, n41016);
  not g68512 (n_30545, n41021);
  and g68513 (n41022, n_30544, n_30545);
  not g68514 (n_30546, n41022);
  and g68515 (n41023, pi1156, n_30546);
  not g68516 (n_30547, n41007);
  and g68517 (n41024, n39369, n_30547);
  not g68518 (n_30548, n41023);
  and g68519 (n41025, n_30548, n41024);
  and g68520 (n41026, n_30511, n40992);
  not g68521 (n_30549, n41026);
  and g68522 (n41027, n40996, n_30549);
  and g68523 (n41028, n_30527, n_30537);
  not g68524 (n_30550, n41028);
  and g68525 (n41029, n_30428, n_30550);
  not g68526 (n_30551, n41029);
  and g68527 (n41030, pi1155, n_30551);
  not g68528 (n_30552, n41027);
  and g68529 (n41031, n_30552, n41030);
  not g68530 (n_30553, n40992);
  and g68531 (n41032, n_30553, n_30523);
  not g68532 (n_30554, n41032);
  and g68533 (n41033, n40899, n_30554);
  not g68534 (n_30555, n41033);
  and g68535 (n41034, n_11768, n_30555);
  and g68536 (n41035, pi0243, n41032);
  not g68537 (n_30556, n41035);
  and g68538 (n41036, n41034, n_30556);
  not g68539 (n_30557, n41036);
  and g68540 (n41037, n_11794, n_30557);
  not g68541 (n_30558, n41031);
  and g68542 (n41038, n_30558, n41037);
  and g68543 (n41039, n_30523, n_30549);
  and g68544 (n41040, pi1155, n41039);
  and g68545 (n41041, n_30516, n41039);
  not g68546 (n_30559, n41040);
  not g68547 (n_30560, n41041);
  and g68548 (n41042, n_30559, n_30560);
  not g68549 (n_30561, n41042);
  and g68550 (n41043, pi0243, n_30561);
  and g68551 (n41044, pi0299, n_30436);
  not g68552 (n_30562, n41044);
  and g68553 (n41045, n_30522, n_30562);
  and g68554 (n41046, n_11768, n41045);
  and g68555 (n41047, n_30512, n41046);
  and g68556 (n41048, n_30527, n_30530);
  not g68557 (n_30563, n41048);
  and g68558 (n41049, n_30428, n_30563);
  not g68559 (n_30564, n41047);
  and g68560 (n41050, n_30564, n41049);
  not g68561 (n_30565, n41043);
  not g68562 (n_30566, n41050);
  and g68563 (n41051, n_30565, n_30566);
  not g68564 (n_30567, n41051);
  and g68565 (n41052, pi1156, n_30567);
  not g68566 (n_30568, n41038);
  and g68567 (n41053, n_11810, n_30568);
  not g68568 (n_30569, n41052);
  and g68569 (n41054, n_30569, n41053);
  and g68570 (n41055, n_30527, n_30522);
  not g68571 (n_30570, n41055);
  and g68572 (n41056, pi0243, n_30570);
  and g68573 (n41057, n_30523, n_30528);
  not g68574 (n_30571, n41057);
  and g68575 (n41058, n_30428, n_30571);
  and g68576 (n41059, pi0243, n_30530);
  not g68577 (n_30572, n41059);
  and g68578 (n41060, n_11768, n_30572);
  not g68579 (n_30573, n41058);
  and g68580 (n41061, n_30573, n41060);
  and g68581 (n41062, n_30516, n_30523);
  and g68582 (n41063, n_30428, pi1155);
  and g68583 (n41064, n41062, n41063);
  and g68590 (n41068, n_30538, n41056);
  not g68591 (n_30577, n41068);
  and g68592 (n41069, pi1155, n_30577);
  and g68593 (n41070, n41010, n41062);
  not g68594 (n_30578, n41070);
  and g68595 (n41071, n41069, n_30578);
  and g68596 (n41072, n_30535, n_30562);
  not g68597 (n_30579, n41072);
  and g68598 (n41073, n_30429, n_30579);
  not g68599 (n_30580, n41073);
  and g68600 (n41074, n_30531, n_30580);
  and g68601 (n41075, n_30544, n41074);
  not g68602 (n_30581, n41075);
  and g68603 (n41076, n_11768, n_30581);
  not g68604 (n_30582, n41071);
  not g68605 (n_30583, n41076);
  and g68606 (n41077, n_30582, n_30583);
  not g68607 (n_30584, n41077);
  and g68608 (n41078, pi1156, n_30584);
  not g68609 (n_30585, n41067);
  and g68610 (n41079, n38478, n_30585);
  not g68611 (n_30586, n41078);
  and g68612 (n41080, n_30586, n41079);
  not g68613 (n_30587, n41025);
  not g68614 (n_30588, n41054);
  and g68615 (n41081, n_30587, n_30588);
  not g68616 (n_30589, n41080);
  and g68617 (n41082, n_30589, n41081);
  not g68618 (n_30590, n41082);
  and g68619 (n41083, pi0219, n_30590);
  and g68620 (n41084, n_30553, n_30562);
  and g68621 (n41085, n_11768, n41084);
  not g68622 (n_30591, n41085);
  and g68623 (n41086, n_30542, n_30591);
  and g68624 (n41087, pi0243, n41045);
  and g68625 (n41088, n_30530, n41087);
  not g68626 (n_30592, n41086);
  not g68627 (n_30593, n41088);
  and g68628 (n41089, n_30592, n_30593);
  not g68629 (n_30594, n41089);
  and g68630 (n41090, n_11794, n_30594);
  and g68631 (n41091, n_30516, n_30562);
  and g68632 (n41092, n_30428, n41091);
  and g68633 (n41093, n_30517, n_30522);
  not g68634 (n_30595, n41093);
  and g68635 (n41094, pi0243, n_30595);
  not g68636 (n_30596, n41092);
  not g68637 (n_30597, n41094);
  and g68638 (n41095, n_30596, n_30597);
  and g68639 (n41096, n41090, n41095);
  and g68640 (n41097, n_30517, n_30536);
  and g68641 (n41098, pi1155, n41097);
  not g68642 (n_30598, n41069);
  not g68643 (n_30599, n41098);
  and g68644 (n41099, n_30598, n_30599);
  and g68645 (n41100, n_30535, n41092);
  not g68646 (n_30600, n41099);
  not g68647 (n_30601, n41100);
  and g68648 (n41101, n_30600, n_30601);
  and g68649 (n41102, n_30528, n_30535);
  and g68650 (n41103, n_30517, n41102);
  not g68651 (n_30602, n41103);
  and g68652 (n41104, n_30428, n_30602);
  and g68653 (n41105, n_30537, n_30562);
  and g68654 (n41106, pi0243, n_30536);
  and g68655 (n41107, n41105, n41106);
  not g68656 (n_30603, n41104);
  not g68657 (n_30604, n41107);
  and g68658 (n41108, n_30603, n_30604);
  not g68659 (n_30605, n41108);
  and g68660 (n41109, n_11768, n_30605);
  not g68661 (n_30606, n41101);
  not g68662 (n_30607, n41109);
  and g68663 (n41110, n_30606, n_30607);
  not g68664 (n_30608, n41110);
  and g68665 (n41111, pi1156, n_30608);
  not g68666 (n_30609, n41096);
  and g68667 (n41112, pi1157, n_30609);
  not g68668 (n_30610, n41111);
  and g68669 (n41113, n_30610, n41112);
  and g68670 (n41114, n_11768, n41093);
  not g68671 (n_30611, n41091);
  and g68672 (n41115, n_30611, n41114);
  and g68673 (n41116, n_30517, n_30549);
  not g68674 (n_30612, n41116);
  and g68675 (n41117, pi0243, n_30612);
  and g68676 (n41118, n_30530, n_30562);
  and g68677 (n41119, n_30428, n41118);
  not g68678 (n_30613, n41117);
  not g68679 (n_30614, n41119);
  and g68680 (n41120, n_30613, n_30614);
  and g68681 (n41121, pi1156, n_30564);
  and g68682 (n41122, n41120, n41121);
  not g68683 (n_30615, n41115);
  and g68684 (n41123, n_30615, n41122);
  and g68685 (n41124, pi0243, n41084);
  not g68686 (n_30616, n41034);
  and g68687 (n41125, n_30616, n_30591);
  not g68688 (n_30617, n41124);
  not g68689 (n_30618, n41125);
  and g68690 (n41126, n_30617, n_30618);
  not g68691 (n_30619, n41126);
  and g68692 (n41127, n_11794, n_30619);
  and g68693 (n41128, n41095, n41120);
  not g68694 (n_30620, n41128);
  and g68695 (n41129, pi1155, n_30620);
  not g68696 (n_30621, n41129);
  and g68697 (n41130, n41127, n_30621);
  not g68698 (n_30622, n41123);
  and g68699 (n41131, n_11810, n_30622);
  not g68700 (n_30623, n41130);
  and g68701 (n41132, n_30623, n41131);
  not g68702 (n_30624, n41132);
  and g68703 (n41133, n_7075, n_30624);
  not g68704 (n_30625, n41113);
  and g68705 (n41134, n_30625, n41133);
  not g68706 (n_30626, n41087);
  and g68707 (n41135, n41018, n_30626);
  and g68708 (n41136, n40930, n40979);
  not g68709 (n_30627, n41135);
  not g68710 (n_30628, n41136);
  and g68711 (n41137, n_30627, n_30628);
  and g68712 (n41138, n41127, n41137);
  not g68713 (n_30629, n41122);
  and g68714 (n41139, n_11810, n_30629);
  not g68715 (n_30630, n41138);
  and g68716 (n41140, n_30630, n41139);
  and g68717 (n41141, n41090, n_30627);
  and g68718 (n41142, n_30580, n41110);
  not g68719 (n_30631, n41142);
  and g68720 (n41143, pi1156, n_30631);
  not g68721 (n_30632, n41141);
  and g68722 (n41144, pi1157, n_30632);
  not g68723 (n_30633, n41143);
  and g68724 (n41145, n_30633, n41144);
  not g68725 (n_30634, n41140);
  and g68726 (n41146, pi0211, n_30634);
  not g68727 (n_30635, n41145);
  and g68728 (n41147, n_30635, n41146);
  not g68729 (n_30636, n41134);
  and g68730 (n41148, n_6791, n_30636);
  not g68731 (n_30637, n41147);
  and g68732 (n41149, n_30637, n41148);
  not g68733 (n_30638, n41083);
  and g68734 (n41150, n40861, n_30638);
  not g68735 (n_30639, n41149);
  and g68736 (n41151, n_30639, n41150);
  not g68737 (n_30640, n40978);
  and g68738 (n41152, n_4226, n_30640);
  not g68739 (n_30641, n41151);
  and g68740 (n41153, n_30641, n41152);
  not g68741 (n_30642, n40907);
  and g68742 (n41154, n_30642, n40910);
  not g68743 (n_30643, n41153);
  and g68744 (n41155, n_30643, n41154);
  and g68745 (n41156, n_4226, n40977);
  and g68746 (n41157, po1038, n40904);
  not g68747 (n_30644, n40910);
  not g68748 (n_30645, n41157);
  and g68749 (n41158, n_30644, n_30645);
  not g68750 (n_30646, n41156);
  and g68751 (n41159, n_30646, n41158);
  not g68752 (n_30647, n41159);
  and g68753 (n41160, n_28510, n_30647);
  not g68754 (n_30648, n41155);
  and g68755 (n41161, n_30648, n41160);
  and g68756 (n41162, n_25711, n_30446);
  not g68757 (n_30649, n39467);
  and g68758 (n41163, pi0199, n_30649);
  not g68764 (n_30652, n41162);
  and g68765 (n41167, pi0230, n_30652);
  not g68766 (n_30653, n41166);
  and g68767 (n41168, n_30653, n41167);
  not g68768 (n_30654, n41161);
  not g68769 (n_30655, n41168);
  and g68770 (po0400, n_30654, n_30655);
  and g68771 (n41170, n_28510, n_2688);
  not g68772 (n_30656, n40405);
  and g68773 (n41171, pi0213, n_30656);
  and g68774 (n41172, n_7075, n_28615);
  and g68775 (n41173, n_30022, n41172);
  not g68776 (n_30657, n41173);
  and g68777 (n41174, n_30023, n_30657);
  not g68778 (n_30658, n41174);
  and g68779 (n41175, n40344, n_30658);
  and g68780 (n41176, n_28653, n40390);
  not g68781 (n_30659, n40383);
  not g68782 (n_30660, n41176);
  and g68783 (n41177, n_30659, n_30660);
  not g68784 (n_30661, n41177);
  and g68785 (n41178, n_30062, n_30661);
  not g68786 (n_30662, n41178);
  and g68787 (n41179, pi0214, n_30662);
  not g68788 (n_30663, n41179);
  and g68789 (n41180, n40364, n_30663);
  and g68790 (n41181, n38420, n40293);
  and g68791 (n41182, n_26565, n41177);
  not g68792 (n_30664, n41181);
  and g68793 (n41183, pi0212, n_30664);
  not g68794 (n_30665, n41182);
  and g68795 (n41184, n_30665, n41183);
  and g68796 (n41185, n_30062, n41184);
  not g68797 (n_30666, n41180);
  and g68798 (n41186, n_6791, n_30666);
  not g68799 (n_30667, n41185);
  and g68800 (n41187, n_30667, n41186);
  not g68801 (n_30668, n41175);
  and g68802 (n41188, n40447, n_30668);
  not g68803 (n_30669, n41187);
  and g68804 (n41189, n_30669, n41188);
  and g68805 (n41190, pi0299, n39410);
  and g68806 (n41191, pi0214, n41177);
  not g68807 (n_30670, n41191);
  and g68808 (n41192, n40388, n_30670);
  and g68809 (n41193, n_30041, n41184);
  not g68810 (n_30671, n41192);
  and g68811 (n41194, n_6791, n_30671);
  not g68812 (n_30672, n41193);
  and g68813 (n41195, n_30672, n41194);
  not g68824 (n_30677, n41171);
  not g68825 (n_30678, n41201);
  and g68826 (n41202, n_30677, n_30678);
  not g68827 (n_30679, n41202);
  and g68828 (n41203, pi0209, n_30679);
  not g68829 (n_30680, n39427);
  and g68830 (n41204, n_26557, n_30680);
  and g68831 (n41205, n40244, n_29937);
  not g68832 (n_30681, n40224);
  not g68833 (n_30682, n41205);
  and g68834 (n41206, n_30681, n_30682);
  and g68835 (n41207, n_7077, n40236);
  and g68836 (n41208, n10843, n_29926);
  not g68837 (n_30683, n40246);
  and g68838 (n41209, n40244, n_30683);
  and g68845 (n41213, n_29289, n_29944);
  not g68846 (n_30687, n41212);
  and g68847 (n41214, n_30687, n41213);
  not g68848 (n_30688, n41214);
  and g68849 (n41215, n_4226, n_30688);
  not g68850 (n_30689, n41206);
  not g68851 (n_30690, n41215);
  and g68852 (n41216, n_30689, n_30690);
  not g68853 (n_30691, n41216);
  and g68854 (n41217, pi0213, n_30691);
  not g68855 (n_30692, n41204);
  and g68856 (n41218, n_26372, n_30692);
  not g68857 (n_30693, n41217);
  and g68858 (n41219, n_30693, n41218);
  not g68859 (n_30694, n41203);
  not g68860 (n_30695, n41219);
  and g68861 (n41220, n_30694, n_30695);
  not g68862 (n_30696, n41220);
  and g68863 (n41221, pi0230, n_30696);
  not g68864 (n_30697, n41170);
  not g68865 (n_30698, n41221);
  and g68866 (po0401, n_30697, n_30698);
  not g68867 (n_30699, n40824);
  and g68868 (n41223, n_26557, n_30699);
  and g68869 (n41224, pi1146, n39869);
  not g68870 (n_30700, n41224);
  and g68871 (n41225, n_29810, n_30700);
  and g68872 (n41226, n39865, n_29860);
  not g68873 (n_30701, n41226);
  and g68874 (n41227, n41225, n_30701);
  and g68875 (n41228, n_28511, n40800);
  not g68876 (n_30702, n41228);
  and g68877 (n41229, n40819, n_30702);
  not g68878 (n_30703, n41229);
  and g68879 (n41230, n_4226, n_30703);
  and g68880 (n41231, pi0214, n_29928);
  not g68881 (n_30704, n40804);
  and g68882 (n41232, n_234, n_30704);
  not g68883 (n_30705, n41232);
  and g68884 (n41233, n41231, n_30705);
  not g68885 (n_30706, n41233);
  and g68886 (n41234, pi0212, n_30706);
  and g68887 (n41235, n_234, n40802);
  not g68888 (n_30707, n41235);
  and g68889 (n41236, n_7075, n_30707);
  not g68890 (n_30708, n41236);
  and g68891 (n41237, n40794, n_30708);
  and g68892 (n41238, n_26565, n41237);
  not g68893 (n_30709, n41238);
  and g68894 (n41239, n41234, n_30709);
  not g68895 (n_30710, n41237);
  and g68896 (n41240, n40796, n_30710);
  not g68897 (n_30711, n41240);
  and g68898 (n41241, n_6791, n_30711);
  not g68899 (n_30712, n41239);
  and g68900 (n41242, n_30712, n41241);
  not g68901 (n_30713, n41242);
  and g68902 (n41243, n41230, n_30713);
  not g68903 (n_30714, n41243);
  and g68904 (n41244, n41227, n_30714);
  and g68905 (n41245, pi1147, n_29807);
  and g68906 (n41246, n_30700, n41245);
  and g68907 (n41247, pi0211, n_30366);
  not g68908 (n_30715, n41247);
  and g68909 (n41248, n_30708, n_30715);
  not g68910 (n_30716, n41248);
  and g68911 (n41249, pi0214, n_30716);
  and g68912 (n41250, n_26565, n_30707);
  not g68913 (n_30717, n41249);
  not g68914 (n_30718, n41250);
  and g68915 (n41251, n_30717, n_30718);
  not g68916 (n_30719, n41251);
  and g68917 (n41252, pi0212, n_30719);
  and g68918 (n41253, n40796, n_30707);
  not g68919 (n_30720, n41253);
  and g68920 (n41254, n_6791, n_30720);
  not g68921 (n_30721, n41252);
  and g68922 (n41255, n_30721, n41254);
  not g68923 (n_30722, n41255);
  and g68924 (n41256, n41230, n_30722);
  not g68925 (n_30723, n41256);
  and g68926 (n41257, n41246, n_30723);
  not g68927 (n_30724, n41244);
  and g68928 (n41258, pi1148, n_30724);
  not g68929 (n_30725, n41257);
  and g68930 (n41259, n_30725, n41258);
  not g68931 (n_30726, n40407);
  not g68932 (n_30727, n41246);
  and g68933 (n41260, n_30726, n_30727);
  and g68934 (n41261, n_8688, n40794);
  not g68935 (n_30728, n41261);
  and g68936 (n41262, n_26565, n_30728);
  not g68937 (n_30729, n41262);
  and g68938 (n41263, n_30717, n_30729);
  not g68939 (n_30730, n41263);
  and g68940 (n41264, pi0212, n_30730);
  and g68941 (n41265, n40796, n_30728);
  not g68942 (n_30731, n41265);
  and g68943 (n41266, n_6791, n_30731);
  not g68944 (n_30732, n41264);
  and g68945 (n41267, n_30732, n41266);
  not g68946 (n_30733, n41267);
  and g68947 (n41268, n41230, n_30733);
  not g68948 (n_30734, n41260);
  not g68949 (n_30735, n41268);
  and g68950 (n41269, n_30734, n_30735);
  and g68951 (n41270, n_30364, n41234);
  and g68952 (n41271, n_26538, n_30378);
  not g68953 (n_30736, n41271);
  and g68954 (n41272, n_6791, n_30736);
  not g68955 (n_30737, n41270);
  and g68956 (n41273, n_30737, n41272);
  not g68957 (n_30738, n41273);
  and g68958 (n41274, n41230, n_30738);
  not g68959 (n_30739, n41274);
  and g68960 (n41275, n41225, n_30739);
  not g68961 (n_30740, n41269);
  and g68962 (n41276, n_29904, n_30740);
  not g68963 (n_30741, n41275);
  and g68964 (n41277, n_30741, n41276);
  not g68965 (n_30742, n41259);
  not g68966 (n_30743, n41277);
  and g68967 (n41278, n_30742, n_30743);
  not g68968 (n_30744, n41278);
  and g68969 (n41279, pi0213, n_30744);
  not g68970 (n_30745, n41223);
  and g68971 (n41280, n_26372, n_30745);
  not g68972 (n_30746, n41279);
  and g68973 (n41281, n_30746, n41280);
  and g68974 (n41282, pi0199, pi1146);
  not g68975 (n_30747, n41282);
  and g68976 (n41283, n38699, n_30747);
  not g68977 (n_30748, n41283);
  and g68978 (n41284, n38550, n_30748);
  not g68979 (n_30749, n41284);
  and g68980 (n41285, n_6900, n_30749);
  and g68981 (n41286, n40339, n_30748);
  and g68982 (n41287, pi0207, n41286);
  not g68983 (n_30750, n41287);
  and g68984 (n41288, n_28828, n_30750);
  not g68985 (n_30751, n41285);
  not g68986 (n_30752, n41288);
  and g68987 (n41289, n_30751, n_30752);
  and g68988 (n41290, n_28512, n41289);
  not g68989 (n_30753, n41290);
  and g68990 (n41291, pi0219, n_30753);
  and g68991 (n41292, n38449, n41284);
  and g68992 (n41293, pi0208, n41286);
  and g68993 (n41294, n_7045, n_30747);
  not g68994 (n_30754, n41294);
  and g68995 (n41295, n38550, n_30754);
  and g68996 (n41296, n_25873, n41295);
  not g68997 (n_30755, n41296);
  and g68998 (n41297, n_29958, n_30755);
  and g68999 (n41298, n_30750, n41297);
  not g69000 (n_30756, n41298);
  and g69001 (n41299, pi0208, n_30756);
  and g69002 (n41300, n_234, n41299);
  not g69003 (n_30757, n41292);
  not g69004 (n_30758, n41293);
  and g69005 (n41301, n_30757, n_30758);
  not g69006 (n_30759, n41300);
  and g69007 (n41302, n_30759, n41301);
  and g69008 (n41303, n_29958, n41302);
  not g69009 (n_30760, n41303);
  and g69010 (n41304, n38414, n_30760);
  not g69011 (n_30761, n41304);
  and g69012 (n41305, n41291, n_30761);
  not g69013 (n_30762, n41289);
  and g69014 (n41306, n_26565, n_30762);
  not g69015 (n_30763, n41306);
  and g69016 (n41307, n_26538, n_30763);
  and g69017 (n41308, n_234, n41302);
  not g69018 (n_30764, n41308);
  and g69019 (n41309, n41307, n_30764);
  not g69020 (n_30765, n41309);
  and g69021 (n41310, n_6791, n_30765);
  and g69022 (n41311, pi0212, n_30764);
  and g69023 (n41312, n10484, n41303);
  not g69024 (n_30766, n41312);
  and g69025 (n41313, n41311, n_30766);
  not g69026 (n_30767, n41313);
  and g69027 (n41314, n41310, n_30767);
  not g69028 (n_30768, n41305);
  and g69029 (n41315, n_4226, n_30768);
  not g69030 (n_30769, n41314);
  and g69031 (n41316, n_30769, n41315);
  not g69032 (n_30770, n41316);
  and g69033 (n41317, n41246, n_30770);
  and g69034 (n41318, n_26242, n40234);
  and g69035 (n41319, n40339, n_30754);
  and g69036 (n41320, pi0207, n41319);
  and g69037 (n41321, pi1146, n_28724);
  not g69038 (n_30771, n41320);
  not g69039 (n_30772, n41321);
  and g69040 (n41322, n_30771, n_30772);
  not g69041 (n_30773, n41322);
  and g69042 (n41323, pi0208, n_30773);
  and g69043 (n41324, n_25873, n_30758);
  and g69044 (n41325, n39658, n_30748);
  not g69045 (n_30774, n41324);
  and g69046 (n41326, n_30774, n41325);
  not g69047 (n_30775, n41318);
  not g69048 (n_30776, n41323);
  and g69049 (n41327, n_30775, n_30776);
  not g69050 (n_30777, n41326);
  and g69051 (n41328, n_30777, n41327);
  not g69052 (n_30778, n41328);
  and g69053 (n41329, n_234, n_30778);
  not g69054 (n_30779, n41329);
  and g69055 (n41330, n_26565, n_30779);
  not g69056 (n_30780, n41330);
  and g69057 (n41331, n_26538, n_30780);
  and g69058 (n41332, n_6900, n_29484);
  not g69059 (n_30781, n41332);
  and g69060 (n41333, n41319, n_30781);
  not g69061 (n_30782, n41333);
  and g69062 (n41334, pi0211, n_30782);
  not g69063 (n_30783, n41319);
  and g69064 (n41335, n_234, n_30783);
  not g69065 (n_30784, n41335);
  and g69066 (n41336, n_30778, n_30784);
  not g69067 (n_30785, n41336);
  and g69068 (n41337, n_234, n_30785);
  and g69069 (n41338, n_7075, n41337);
  not g69070 (n_30786, n41334);
  not g69071 (n_30787, n41338);
  and g69072 (n41339, n_30786, n_30787);
  not g69073 (n_30788, n41339);
  and g69074 (n41340, n_30779, n_30788);
  not g69075 (n_30789, n41340);
  and g69076 (n41341, n41331, n_30789);
  not g69077 (n_30790, n41341);
  and g69078 (n41342, n_6791, n_30790);
  and g69079 (n41343, n41231, n_30779);
  and g69080 (n41344, n_26565, n41340);
  not g69081 (n_30791, n41344);
  and g69082 (n41345, pi0212, n_30791);
  not g69083 (n_30792, n41343);
  and g69084 (n41346, n_30792, n41345);
  not g69085 (n_30793, n41346);
  and g69086 (n41347, n41342, n_30793);
  and g69087 (n41348, n_28512, n41329);
  not g69088 (n_30794, n41348);
  and g69089 (n41349, pi0219, n_30794);
  and g69090 (n41350, n38414, n_30778);
  not g69091 (n_30795, n41350);
  and g69092 (n41351, n41349, n_30795);
  not g69093 (n_30796, n41351);
  and g69094 (n41352, n_4226, n_30796);
  not g69095 (n_30797, n41347);
  and g69096 (n41353, n_30797, n41352);
  not g69097 (n_30798, n41353);
  and g69098 (n41354, n41227, n_30798);
  not g69099 (n_30799, n41317);
  and g69100 (n41355, pi1148, n_30799);
  not g69101 (n_30800, n41354);
  and g69102 (n41356, n_30800, n41355);
  and g69103 (n41357, n_30258, n_30779);
  not g69104 (n_30801, n41357);
  and g69105 (n41358, n_30773, n_30801);
  not g69106 (n_30802, n41358);
  and g69107 (n41359, n_6791, n_30802);
  and g69108 (n41360, pi0219, n_30782);
  not g69109 (n_30803, n41360);
  and g69110 (n41361, n_28940, n_30803);
  and g69111 (n41362, n_28511, n_30786);
  and g69112 (n41363, n41336, n41362);
  not g69113 (n_30804, n41361);
  not g69114 (n_30805, n41363);
  and g69115 (n41364, n_30804, n_30805);
  not g69116 (n_30806, n41364);
  and g69117 (n41365, n_4226, n_30806);
  not g69118 (n_30807, n41359);
  and g69119 (n41366, n_30807, n41365);
  not g69120 (n_30808, n41366);
  and g69121 (n41367, n41225, n_30808);
  not g69122 (n_30809, n41295);
  and g69123 (n41368, n_6900, n_30809);
  not g69124 (n_30810, n41368);
  and g69125 (n41369, n_30752, n_30810);
  not g69126 (n_30811, n41369);
  and g69127 (n41370, n_8688, n_30811);
  not g69128 (n_30812, n41370);
  and g69129 (n41371, pi0214, n_30812);
  and g69130 (n41372, n_26565, n41369);
  not g69131 (n_30813, n41372);
  and g69132 (n41373, n_26538, n_30813);
  not g69133 (n_30814, n41371);
  and g69134 (n41374, n_30814, n41373);
  and g69135 (n41375, n_26565, n_30812);
  and g69136 (n41376, n38449, n41295);
  not g69137 (n_30815, n41376);
  and g69138 (n41377, n_30775, n_30815);
  not g69139 (n_30816, n41299);
  and g69140 (n41378, n_30816, n41377);
  and g69141 (n41379, n_234, n41378);
  not g69142 (n_30817, n41379);
  and g69143 (n41380, pi0214, n_30817);
  and g69144 (n41381, n_7075, n_30764);
  not g69145 (n_30818, n41381);
  and g69146 (n41382, n_30762, n_30818);
  not g69147 (n_30819, n41382);
  and g69148 (n41383, n41380, n_30819);
  not g69149 (n_30820, n41383);
  and g69150 (n41384, pi0212, n_30820);
  not g69151 (n_30821, n41375);
  and g69152 (n41385, n_30821, n41384);
  not g69153 (n_30822, n41374);
  not g69154 (n_30823, n41385);
  and g69155 (n41386, n_30822, n_30823);
  not g69156 (n_30824, n41386);
  and g69157 (n41387, n_6791, n_30824);
  and g69158 (n41388, n_803, n_30177);
  not g69159 (n_30825, n41388);
  and g69160 (n41389, n40299, n_30825);
  not g69161 (n_30826, n41389);
  and g69162 (n41390, n41387, n_30826);
  and g69163 (n41391, n_28511, n41369);
  not g69164 (n_30827, n41391);
  and g69165 (n41392, n_28512, n_30827);
  not g69166 (n_30828, n41378);
  not g69167 (n_30829, n41392);
  and g69168 (n41393, n_30828, n_30829);
  and g69169 (n41394, n_26538, n41372);
  not g69170 (n_30830, n41394);
  and g69171 (n41395, pi0219, n_30830);
  not g69172 (n_30831, n41393);
  and g69173 (n41396, n_30831, n41395);
  not g69174 (n_30832, n41396);
  and g69175 (n41397, n_4226, n_30832);
  not g69176 (n_30833, n41390);
  and g69177 (n41398, n_30833, n41397);
  not g69178 (n_30834, n41398);
  and g69179 (n41399, n_30734, n_30834);
  not g69180 (n_30835, n41367);
  and g69181 (n41400, n_29904, n_30835);
  not g69182 (n_30836, n41399);
  and g69183 (n41401, n_30836, n41400);
  not g69184 (n_30837, n41356);
  not g69185 (n_30838, n41401);
  and g69186 (n41402, n_30837, n_30838);
  not g69187 (n_30839, n41402);
  and g69188 (n41403, pi0213, n_30839);
  and g69189 (n41404, pi1147, n_4226);
  and g69190 (n41405, n_28654, n41302);
  not g69191 (n_30840, n41405);
  and g69192 (n41406, n38414, n_30840);
  not g69193 (n_30841, n41406);
  and g69194 (n41407, n41291, n_30841);
  and g69195 (n41408, n_29926, n41302);
  and g69196 (n41409, pi0214, n41408);
  not g69197 (n_30842, n41409);
  and g69198 (n41410, n41307, n_30842);
  and g69199 (n41411, pi0299, n_30350);
  not g69200 (n_30843, n41411);
  and g69201 (n41412, n41302, n_30843);
  not g69202 (n_30844, n41412);
  and g69203 (n41413, pi0212, n_30844);
  not g69204 (n_30845, n41413);
  and g69205 (n41414, n_6791, n_30845);
  not g69206 (n_30846, n41410);
  and g69207 (n41415, n_30846, n41414);
  not g69208 (n_30847, n41407);
  and g69209 (n41416, n41404, n_30847);
  not g69210 (n_30848, n41415);
  and g69211 (n41417, n_30848, n41416);
  and g69212 (n41418, n_234, n41328);
  not g69213 (n_30849, n41418);
  and g69214 (n41419, n38414, n_30849);
  and g69215 (n41420, n_28653, n41419);
  not g69216 (n_30850, n41420);
  and g69217 (n41421, n41349, n_30850);
  and g69218 (n41422, n_29926, n_30779);
  not g69219 (n_30851, n41422);
  and g69220 (n41423, n41331, n_30851);
  and g69221 (n41424, n_30779, n_30843);
  not g69222 (n_30852, n41424);
  and g69223 (n41425, pi0212, n_30852);
  not g69224 (n_30853, n41425);
  and g69225 (n41426, n_6791, n_30853);
  not g69226 (n_30854, n41423);
  and g69227 (n41427, n_30854, n41426);
  not g69228 (n_30855, n41421);
  and g69229 (n41428, n40447, n_30855);
  not g69230 (n_30856, n41427);
  and g69231 (n41429, n_30856, n41428);
  and g69237 (n41433, n_30817, n41413);
  not g69238 (n_30859, n41408);
  and g69239 (n41434, n41380, n_30859);
  not g69240 (n_30860, n41434);
  and g69241 (n41435, n_30813, n_30860);
  not g69242 (n_30861, n41435);
  and g69243 (n41436, n_26538, n_30861);
  not g69244 (n_30862, n41433);
  and g69245 (n41437, n_6791, n_30862);
  not g69246 (n_30863, n41436);
  and g69247 (n41438, n_30863, n41437);
  and g69248 (n41439, n_30817, n_30840);
  not g69249 (n_30864, n41439);
  and g69250 (n41440, n_7075, n_30864);
  not g69251 (n_30865, n41440);
  and g69252 (n41441, n_30829, n_30865);
  not g69253 (n_30866, n41441);
  and g69254 (n41442, n41395, n_30866);
  not g69255 (n_30867, n41438);
  and g69256 (n41443, n41404, n_30867);
  not g69257 (n_30868, n41442);
  and g69258 (n41444, n_30868, n41443);
  and g69259 (n41445, n_30784, n41425);
  and g69260 (n41446, n_26565, n41333);
  not g69261 (n_30869, n41337);
  and g69262 (n41447, pi0214, n_30869);
  and g69263 (n41448, n_30851, n41447);
  not g69264 (n_30870, n41446);
  not g69265 (n_30871, n41448);
  and g69266 (n41449, n_30870, n_30871);
  not g69267 (n_30872, n41449);
  and g69268 (n41450, n_26538, n_30872);
  not g69269 (n_30873, n41445);
  and g69270 (n41451, n_6791, n_30873);
  not g69271 (n_30874, n41450);
  and g69272 (n41452, n_30874, n41451);
  and g69273 (n41453, n_28653, n_30869);
  not g69274 (n_30875, n41453);
  and g69275 (n41454, n_7075, n_30875);
  not g69276 (n_30876, n41454);
  and g69277 (n41455, n41362, n_30876);
  not g69278 (n_30877, n41455);
  and g69279 (n41456, n_30804, n_30877);
  not g69280 (n_30878, n41456);
  and g69281 (n41457, n40447, n_30878);
  not g69282 (n_30879, n41452);
  and g69283 (n41458, n_30879, n41457);
  not g69289 (n_30882, n41432);
  and g69290 (n41462, n_26557, n_30882);
  not g69291 (n_30883, n41461);
  and g69292 (n41463, n_30883, n41462);
  not g69293 (n_30884, n41463);
  and g69294 (n41464, pi0209, n_30884);
  not g69295 (n_30885, n41403);
  and g69296 (n41465, n_30885, n41464);
  not g69297 (n_30886, n41281);
  not g69298 (n_30887, n41465);
  and g69299 (n41466, n_30886, n_30887);
  not g69300 (n_30888, n41466);
  and g69301 (n41467, pi0230, n_30888);
  and g69302 (n41468, n_28510, n_2498);
  not g69303 (n_30889, n41467);
  not g69304 (n_30890, n41468);
  and g69305 (po0402, n_30889, n_30890);
  and g69306 (n41470, n_30133, n40134);
  and g69307 (n41471, pi1150, n40089);
  not g69308 (n_30891, n41470);
  and g69309 (n41472, pi1149, n_30891);
  not g69310 (n_30892, n41471);
  and g69311 (n41473, n_30892, n41472);
  and g69312 (n41474, n_30133, n40200);
  and g69313 (n41475, pi1150, n40166);
  not g69314 (n_30893, n41474);
  and g69315 (n41476, n_29850, n_30893);
  not g69316 (n_30894, n41475);
  and g69317 (n41477, n_30894, n41476);
  not g69318 (n_30895, n41473);
  not g69319 (n_30896, n41477);
  and g69320 (n41478, n_30895, n_30896);
  not g69321 (n_30897, n41478);
  and g69322 (n41479, pi1148, n_30897);
  and g69323 (n41480, n_30133, n40125);
  and g69324 (n41481, pi1150, n40078);
  not g69325 (n_30898, n41481);
  and g69326 (n41482, pi1149, n_30898);
  not g69327 (n_30899, n41480);
  and g69328 (n41483, n_30899, n41482);
  and g69329 (n41484, n_29850, pi1150);
  and g69330 (n41485, n_30219, n41484);
  not g69331 (n_30900, n41483);
  not g69332 (n_30901, n41485);
  and g69333 (n41486, n_30900, n_30901);
  not g69334 (n_30902, n41486);
  and g69335 (n41487, n_29904, n_30902);
  not g69336 (n_30903, n41479);
  not g69337 (n_30904, n41487);
  and g69338 (n41488, n_30903, n_30904);
  not g69339 (n_30905, n41488);
  and g69340 (n41489, pi0213, n_30905);
  and g69341 (n41490, n_29888, n_29896);
  not g69342 (n_30906, n41490);
  and g69343 (n41491, n41227, n_30906);
  not g69344 (n_30907, n41227);
  and g69345 (n41492, n_30907, n_30727);
  and g69346 (n41493, pi0219, n_29958);
  not g69347 (n_30908, n41493);
  and g69348 (n41494, n40084, n_30908);
  and g69349 (n41495, n40127, n_29885);
  not g69350 (n_30909, n41494);
  not g69351 (n_30910, n41495);
  and g69352 (n41496, n_30909, n_30910);
  and g69353 (n41497, n_29898, n_29941);
  not g69354 (n_30911, n41497);
  and g69355 (n41498, n38423, n_30911);
  not g69356 (n_30912, n41498);
  and g69357 (n41499, n_30248, n_30912);
  not g69358 (n_30913, n41499);
  and g69359 (n41500, n_6791, n_30913);
  not g69360 (n_30914, n41496);
  not g69361 (n_30915, n41500);
  and g69362 (n41501, n_30914, n_30915);
  not g69363 (n_30916, n41492);
  not g69364 (n_30917, n41501);
  and g69365 (n41502, n_30916, n_30917);
  not g69366 (n_30918, n41491);
  and g69367 (n41503, n_30133, n_30918);
  not g69368 (n_30919, n41502);
  and g69369 (n41504, n_30919, n41503);
  and g69370 (n41505, n_29955, n_30909);
  and g69371 (n41506, n_26565, n39697);
  and g69372 (n41507, pi0214, n_29862);
  and g69373 (n41508, n_29960, n41507);
  not g69374 (n_30920, n41506);
  and g69375 (n41509, pi0212, n_30920);
  not g69376 (n_30921, n41508);
  and g69377 (n41510, n_30921, n41509);
  not g69378 (n_30922, n41510);
  and g69379 (n41511, n40156, n_30922);
  not g69380 (n_30923, n41505);
  not g69381 (n_30924, n41511);
  and g69382 (n41512, n_30923, n_30924);
  not g69383 (n_30925, n41512);
  and g69384 (n41513, n41227, n_30925);
  and g69385 (n41514, n_29961, n40513);
  and g69386 (n41515, n_26538, n_29486);
  not g69387 (n_30926, n41515);
  and g69388 (n41516, n_6791, n_30926);
  not g69389 (n_30927, n40525);
  and g69390 (n41517, n_30927, n41516);
  not g69391 (n_30928, n41514);
  and g69392 (n41518, n_30928, n41517);
  not g69393 (n_30929, n41518);
  and g69394 (n41519, n_30923, n_30929);
  not g69395 (n_30930, n41519);
  and g69396 (n41520, n41246, n_30930);
  not g69397 (n_30931, n41513);
  and g69398 (n41521, pi1150, n_30931);
  not g69399 (n_30932, n41520);
  and g69400 (n41522, n_30932, n41521);
  not g69401 (n_30933, n41504);
  not g69402 (n_30934, n41522);
  and g69403 (n41523, n_30933, n_30934);
  not g69404 (n_30935, n41523);
  and g69405 (n41524, pi1148, n_30935);
  and g69406 (n41525, pi1150, n39639);
  and g69407 (n41526, pi0299, n40093);
  not g69414 (n_30938, n40213);
  and g69415 (n41531, n_6791, n_30938);
  not g69416 (n_30939, n41531);
  and g69417 (n41532, n_30259, n_30939);
  and g69418 (n41533, n41494, n41532);
  not g69419 (n_30940, n41533);
  and g69420 (n41534, n41225, n_30940);
  and g69421 (n41535, n_30734, n_30909);
  not g69422 (n_30941, n41534);
  not g69423 (n_30942, n41535);
  and g69424 (n41536, n_30941, n_30942);
  and g69425 (n41537, pi1150, n40140);
  not g69426 (n_30943, n41536);
  not g69427 (n_30944, n41537);
  and g69428 (n41538, n_30943, n_30944);
  not g69429 (n_30945, n41530);
  and g69430 (n41539, n_29904, n_30945);
  not g69431 (n_30946, n41538);
  and g69432 (n41540, n_30946, n41539);
  not g69433 (n_30947, n41524);
  not g69434 (n_30948, n41540);
  and g69435 (n41541, n_30947, n_30948);
  not g69436 (n_30949, n41541);
  and g69437 (n41542, n_29850, n_30949);
  and g69438 (n41543, n_803, n40122);
  and g69439 (n41544, n40084, n_29829);
  not g69440 (n_30950, n40123);
  not g69441 (n_30951, n41544);
  and g69442 (n41545, n_30950, n_30951);
  and g69443 (n41546, n40213, n40293);
  not g69444 (n_30952, n41546);
  and g69445 (n41547, n_29824, n_30952);
  and g69446 (n41548, n40121, n41547);
  not g69447 (n_30953, n41543);
  not g69448 (n_30954, n41545);
  and g69449 (n41549, n_30953, n_30954);
  not g69450 (n_30955, n41548);
  and g69451 (n41550, n_30955, n41549);
  not g69452 (n_30956, n41550);
  and g69453 (n41551, n_30734, n_30956);
  not g69454 (n_30957, n40524);
  and g69455 (n41552, n_29826, n_30957);
  not g69456 (n_30958, n41552);
  and g69457 (n41553, n_6791, n_30958);
  not g69458 (n_30959, n41553);
  and g69459 (n41554, n_30954, n_30959);
  and g69460 (n41555, n_803, n_29824);
  not g69461 (n_30960, n41555);
  and g69462 (n41556, n41554, n_30960);
  not g69463 (n_30961, n41556);
  and g69464 (n41557, n41225, n_30961);
  not g69465 (n_30962, n41557);
  and g69466 (n41558, n_30133, n_30962);
  not g69467 (n_30963, n41551);
  and g69468 (n41559, n_30963, n41558);
  and g69469 (n41560, n_29985, n_30909);
  not g69470 (n_30964, n40725);
  and g69471 (n41561, n_29795, n_30964);
  and g69472 (n41562, n_26565, n40725);
  not g69473 (n_30965, n41562);
  and g69474 (n41563, n40074, n_30965);
  not g69475 (n_30966, n41563);
  and g69476 (n41564, n_6791, n_30966);
  not g69477 (n_30967, n41561);
  and g69478 (n41565, n_30967, n41564);
  and g69479 (n41566, n_26538, n41561);
  not g69480 (n_30968, n41566);
  and g69481 (n41567, n41564, n_30968);
  and g69482 (n41568, n_234, n39713);
  not g69487 (n_30970, n41560);
  not g69488 (n_30971, n41565);
  and g69489 (n41572, n_30970, n_30971);
  not g69490 (n_30972, n41571);
  and g69491 (n41573, n_30972, n41572);
  not g69492 (n_30973, n41573);
  and g69493 (n41574, n_29793, n_30973);
  and g69494 (n41575, n40063, n_29803);
  not g69495 (n_30974, n41575);
  and g69496 (n41576, n_6791, n_30974);
  not g69497 (n_30975, n40729);
  and g69498 (n41577, n_30975, n41576);
  not g69499 (n_30976, n41577);
  and g69500 (n41578, n40310, n_30976);
  not g69501 (n_30977, n41574);
  and g69502 (n41579, n_30977, n41578);
  not g69503 (n_30978, n41579);
  and g69504 (n41580, n41225, n_30978);
  and g69505 (n41581, n_30734, n_30973);
  not g69506 (n_30979, n41581);
  and g69507 (n41582, pi1150, n_30979);
  not g69508 (n_30980, n41580);
  and g69509 (n41583, n_30980, n41582);
  not g69510 (n_30981, n41583);
  and g69511 (n41584, n_29904, n_30981);
  not g69512 (n_30982, n41559);
  and g69513 (n41585, n_30982, n41584);
  and g69514 (n41586, n_29847, n_30909);
  and g69515 (n41587, n39747, n41231);
  not g69516 (n_30983, n41587);
  and g69517 (n41588, n40189, n_30983);
  and g69518 (n41589, n_29877, n40190);
  not g69519 (n_30984, n41589);
  and g69520 (n41590, n_29882, n_30984);
  not g69521 (n_30985, n41590);
  and g69522 (n41591, n_30907, n_30985);
  not g69523 (n_30986, n41588);
  and g69524 (n41592, n40192, n_30986);
  not g69525 (n_30987, n41591);
  and g69526 (n41593, n_30987, n41592);
  not g69527 (n_30988, n41586);
  not g69528 (n_30989, n41593);
  and g69529 (n41594, n_30988, n_30989);
  not g69530 (n_30990, n41594);
  and g69531 (n41595, n_30916, n_30990);
  not g69532 (n_30991, n41595);
  and g69533 (n41596, n_30133, n_30991);
  and g69534 (n41597, n_29981, n_30940);
  and g69535 (n41598, n41227, n41597);
  and g69536 (n41599, pi0214, n40292);
  not g69537 (n_30992, n41599);
  and g69538 (n41600, n40298, n_30992);
  not g69539 (n_30993, n40295);
  and g69540 (n41601, n_6791, n_30993);
  not g69541 (n_30994, n41600);
  and g69542 (n41602, n_30994, n41601);
  not g69543 (n_30995, n41602);
  and g69544 (n41603, n40291, n_30995);
  and g69545 (n41604, pi1146, n40085);
  not g69546 (n_30996, n41604);
  and g69547 (n41605, n41246, n_30996);
  not g69548 (n_30997, n41603);
  and g69549 (n41606, n_30997, n41605);
  not g69550 (n_30998, n41606);
  and g69551 (n41607, pi1150, n_30998);
  not g69552 (n_30999, n41598);
  and g69553 (n41608, n_30999, n41607);
  not g69554 (n_31000, n41608);
  and g69555 (n41609, pi1148, n_31000);
  not g69556 (n_31001, n41596);
  and g69557 (n41610, n_31001, n41609);
  not g69558 (n_31002, n41610);
  and g69559 (n41611, pi1149, n_31002);
  not g69560 (n_31003, n41585);
  and g69561 (n41612, n_31003, n41611);
  not g69562 (n_31004, n41542);
  not g69563 (n_31005, n41612);
  and g69564 (n41613, n_31004, n_31005);
  not g69565 (n_31006, n41613);
  and g69566 (n41614, n_26557, n_31006);
  not g69567 (n_31007, n41489);
  and g69568 (n41615, pi0209, n_31007);
  not g69569 (n_31008, n41614);
  and g69570 (n41616, n_31008, n41615);
  and g69571 (n41617, n_26557, n_30839);
  and g69572 (n41618, pi0219, n_30811);
  not g69573 (n_31009, n41618);
  and g69574 (n41619, n41404, n_31009);
  not g69575 (n_31010, n41387);
  and g69576 (n41620, n_31010, n41619);
  and g69577 (n41621, n_26538, n_30870);
  and g69578 (n41622, n_8688, n_30782);
  not g69579 (n_31011, n41622);
  and g69580 (n41623, pi0214, n_31011);
  not g69581 (n_31012, n41623);
  and g69582 (n41624, n41621, n_31012);
  and g69583 (n41625, n_26565, n_31011);
  and g69584 (n41626, pi0214, n41339);
  not g69585 (n_31013, n41626);
  and g69586 (n41627, pi0212, n_31013);
  not g69587 (n_31014, n41625);
  and g69588 (n41628, n_31014, n41627);
  not g69589 (n_31015, n41624);
  not g69590 (n_31016, n41628);
  and g69591 (n41629, n_31015, n_31016);
  not g69592 (n_31017, n41629);
  and g69593 (n41630, n_6791, n_31017);
  and g69594 (n41631, n40447, n_30803);
  not g69595 (n_31018, n41630);
  and g69596 (n41632, n_31018, n41631);
  not g69602 (n_31021, n41380);
  and g69603 (n41636, n41373, n_31021);
  and g69604 (n41637, n_26565, n_30817);
  not g69605 (n_31022, n41637);
  and g69606 (n41638, n41384, n_31022);
  not g69607 (n_31023, n41636);
  not g69608 (n_31024, n41638);
  and g69609 (n41639, n_31023, n_31024);
  not g69610 (n_31025, n41639);
  and g69611 (n41640, n_6791, n_31025);
  not g69612 (n_31026, n41640);
  and g69613 (n41641, n_31009, n_31026);
  not g69614 (n_31027, n41641);
  and g69615 (n41642, pi1147, n_31027);
  not g69616 (n_31028, n41447);
  and g69617 (n41643, n_31028, n41621);
  and g69618 (n41644, n_26565, n_30869);
  not g69619 (n_31029, n41644);
  and g69620 (n41645, n41627, n_31029);
  not g69621 (n_31030, n41643);
  not g69622 (n_31031, n41645);
  and g69623 (n41646, n_31030, n_31031);
  not g69624 (n_31032, n41646);
  and g69625 (n41647, n_6791, n_31032);
  not g69626 (n_31033, n41647);
  and g69627 (n41648, n_30803, n_31033);
  not g69628 (n_31034, n41648);
  and g69629 (n41649, n_29810, n_31034);
  not g69630 (n_31035, n41642);
  and g69631 (n41650, n_4226, n_31035);
  not g69632 (n_31036, n41649);
  and g69633 (n41651, n_31036, n41650);
  and g69634 (n41652, pi1150, n_29807);
  not g69635 (n_31037, n41651);
  and g69636 (n41653, n_31037, n41652);
  not g69637 (n_31038, n41635);
  not g69638 (n_31039, n41653);
  and g69639 (n41654, n_31038, n_31039);
  not g69640 (n_31040, n41654);
  and g69641 (n41655, pi1149, n_31040);
  and g69642 (n41656, pi1150, n40207);
  not g69643 (n_31041, n41656);
  and g69644 (n41657, n41333, n_31041);
  not g69645 (n_31042, n41657);
  and g69646 (n41658, n_29810, n_31042);
  and g69647 (n41659, pi1147, n_30811);
  not g69648 (n_31043, n41658);
  and g69649 (n41660, n_4226, n_31043);
  not g69650 (n_31044, n41659);
  and g69651 (n41661, n_31044, n41660);
  and g69652 (n41662, n_29810, n41336);
  not g69653 (n_31045, n41662);
  and g69654 (n41663, n16479, n_31045);
  not g69655 (n_31046, n41663);
  and g69656 (n41664, n41656, n_31046);
  not g69657 (n_31047, n41661);
  and g69658 (n41665, n_29850, n_31047);
  not g69659 (n_31048, n41664);
  and g69660 (n41666, n_31048, n41665);
  not g69661 (n_31049, n41655);
  not g69662 (n_31050, n41666);
  and g69663 (n41667, n_31049, n_31050);
  not g69664 (n_31051, n41667);
  and g69665 (n41668, n_29904, n_31051);
  and g69666 (n41669, n_28511, n41381);
  not g69667 (n_31052, n41669);
  and g69668 (n41670, n41291, n_31052);
  not g69669 (n_31053, n41670);
  and g69670 (n41671, n41404, n_31053);
  and g69671 (n41672, pi0214, n_8688);
  and g69672 (n41673, n41302, n41672);
  not g69673 (n_31054, n41673);
  and g69674 (n41674, pi0212, n_31054);
  and g69675 (n41675, n_30763, n41674);
  and g69676 (n41676, n_26538, n41289);
  not g69677 (n_31055, n41676);
  and g69678 (n41677, n_6791, n_31055);
  not g69679 (n_31056, n41675);
  and g69680 (n41678, n_31056, n41677);
  not g69681 (n_31057, n41678);
  and g69682 (n41679, n41671, n_31057);
  not g69683 (n_31058, n41419);
  and g69684 (n41680, n41349, n_31058);
  not g69685 (n_31059, n41680);
  and g69686 (n41681, n40447, n_31059);
  and g69687 (n41682, n_6791, n41357);
  not g69688 (n_31060, n41682);
  and g69689 (n41683, n41681, n_31060);
  and g69695 (n41687, n_30779, n41622);
  and g69696 (n41688, pi0214, n41687);
  not g69697 (n_31063, n41688);
  and g69698 (n41689, n41345, n_31063);
  not g69699 (n_31064, n41689);
  and g69700 (n41690, n41342, n_31064);
  not g69701 (n_31065, n41690);
  and g69702 (n41691, n41681, n_31065);
  and g69703 (n41692, n_26565, n41382);
  not g69704 (n_31066, n41692);
  and g69705 (n41693, n41674, n_31066);
  and g69706 (n41694, n41307, n_30819);
  not g69707 (n_31067, n41694);
  and g69708 (n41695, n_6791, n_31067);
  not g69709 (n_31068, n41693);
  and g69710 (n41696, n_31068, n41695);
  not g69711 (n_31069, n41696);
  and g69712 (n41697, n41671, n_31069);
  not g69718 (n_31072, n41686);
  and g69719 (n41701, n_29850, n_31072);
  not g69720 (n_31073, n41700);
  and g69721 (n41702, n_31073, n41701);
  and g69722 (n41703, pi0057, n38666);
  and g69723 (n41704, n_3232, n_28735);
  not g69724 (n_31074, n41311);
  and g69725 (n41705, n41310, n_31074);
  not g69726 (n_31075, n41705);
  and g69727 (n41706, n_31053, n_31075);
  and g69728 (n41707, n6305, n41706);
  not g69730 (n_31076, n41704);
  and g69734 (n41711, n6305, n_28696);
  and g69735 (n41712, n41348, n41711);
  and g69736 (n41713, n_28735, n_30849);
  not g69743 (n_31080, n41703);
  not g69744 (n_31081, n41717);
  and g69745 (n41718, n_31080, n_31081);
  not g69746 (n_31082, n41710);
  and g69747 (n41719, n_31082, n41718);
  not g69748 (n_31083, n41719);
  and g69749 (n41720, pi1150, n_31083);
  and g69750 (n41721, n41331, n_31063);
  and g69751 (n41722, n_31028, n41687);
  not g69752 (n_31084, n41722);
  and g69753 (n41723, pi0212, n_31084);
  not g69754 (n_31085, n41721);
  and g69755 (n41724, n_6791, n_31085);
  not g69756 (n_31086, n41723);
  and g69757 (n41725, n_31086, n41724);
  not g69758 (n_31087, n41725);
  and g69759 (n41726, n41681, n_31087);
  and g69760 (n41727, n_30272, n41404);
  and g69761 (n41728, n41706, n41727);
  not g69767 (n_31090, n41731);
  and g69768 (n41732, pi1149, n_31090);
  not g69769 (n_31091, n41720);
  and g69770 (n41733, n_31091, n41732);
  not g69771 (n_31092, n41733);
  and g69772 (n41734, pi1148, n_31092);
  not g69773 (n_31093, n41702);
  and g69774 (n41735, n_31093, n41734);
  not g69775 (n_31094, n41735);
  and g69776 (n41736, pi0213, n_31094);
  not g69777 (n_31095, n41668);
  and g69778 (n41737, n_31095, n41736);
  not g69779 (n_31096, n41617);
  and g69780 (n41738, n_26372, n_31096);
  not g69781 (n_31097, n41737);
  and g69782 (n41739, n_31097, n41738);
  not g69783 (n_31098, n41616);
  not g69784 (n_31099, n41739);
  and g69785 (n41740, n_31098, n_31099);
  not g69786 (n_31100, n41740);
  and g69787 (n41741, pi0230, n_31100);
  and g69788 (n41742, n_28510, n_2128);
  not g69789 (n_31101, n41741);
  not g69790 (n_31102, n41742);
  and g69791 (po0403, n_31101, n_31102);
  and g69792 (n41744, pi0213, n40625);
  and g69793 (n41745, pi1151, n_29848);
  and g69794 (n41746, n40310, n_30971);
  not g69795 (n_31103, n41746);
  and g69796 (n41747, n41745, n_31103);
  not g69797 (n_31104, n40119);
  and g69798 (n41748, n40104, n_31104);
  not g69799 (n_31105, n41748);
  and g69800 (n41749, n_30954, n_31105);
  not g69801 (n_31106, n41749);
  and g69802 (n41750, n_29848, n_31106);
  and g69803 (n41751, n_29468, n41750);
  not g69804 (n_31107, n41747);
  and g69805 (n41752, pi1147, n_31107);
  not g69806 (n_31108, n41751);
  and g69807 (n41753, n_31108, n41752);
  and g69808 (n41754, n_29810, n_30221);
  and g69809 (n41755, pi1151, n_29842);
  not g69810 (n_31109, n41567);
  and g69811 (n41756, n_29805, n_31109);
  not g69812 (n_31110, n41756);
  and g69813 (n41757, n41755, n_31110);
  not g69814 (n_31111, n41757);
  and g69815 (n41758, n41754, n_31111);
  not g69816 (n_31112, n41753);
  and g69817 (n41759, n_29850, n_31112);
  not g69818 (n_31113, n41758);
  and g69819 (n41760, n_31113, n41759);
  and g69820 (n41761, pi1147, n_30224);
  and g69821 (n41762, n_29815, n_29813);
  and g69822 (n41763, n40672, n41762);
  not g69823 (n_31114, n41763);
  and g69824 (n41764, n41761, n_31114);
  and g69825 (n41765, n_29468, n_29807);
  and g69826 (n41766, n40192, n_30984);
  not g69827 (n_31115, n41766);
  and g69828 (n41767, n40680, n_31115);
  and g69829 (n41768, n_29887, n40680);
  not g69830 (n_31116, n41767);
  not g69831 (n_31117, n41768);
  and g69832 (n41769, n_31116, n_31117);
  and g69833 (n41770, n41765, n41769);
  and g69834 (n41771, n40500, n_30997);
  not g69835 (n_31118, n41771);
  and g69836 (n41772, n_29810, n_31118);
  not g69837 (n_31119, n41770);
  and g69838 (n41773, n_31119, n41772);
  not g69839 (n_31120, n41764);
  and g69840 (n41774, pi1149, n_31120);
  not g69841 (n_31121, n41773);
  and g69842 (n41775, n_31121, n41774);
  not g69843 (n_31122, n41775);
  and g69844 (n41776, pi1150, n_31122);
  not g69845 (n_31123, n41760);
  and g69846 (n41777, n_31123, n41776);
  and g69847 (n41778, n_29821, n40141);
  not g69848 (n_31124, n41778);
  and g69849 (n41779, n_29468, n_31124);
  not g69850 (n_31125, n41779);
  and g69851 (n41780, n_29810, n_31125);
  and g69852 (n41781, n39830, n_30158);
  not g69853 (n_31126, n41781);
  and g69854 (n41782, n41755, n_31126);
  not g69855 (n_31127, n41782);
  and g69856 (n41783, n41780, n_31127);
  and g69857 (n41784, n_30293, n41745);
  and g69858 (n41785, n_29849, n40577);
  not g69859 (n_31128, n41785);
  and g69860 (n41786, pi1147, n_31128);
  not g69861 (n_31129, n41784);
  and g69862 (n41787, n_31129, n41786);
  not g69863 (n_31130, n41783);
  and g69864 (n41788, n_29850, n_31130);
  not g69865 (n_31131, n41787);
  and g69866 (n41789, n_31131, n41788);
  and g69867 (n41790, pi0212, n_29507);
  not g69868 (n_31132, n41790);
  and g69869 (n41791, n41517, n_31132);
  not g69870 (n_31133, n41791);
  and g69871 (n41792, n40164, n_31133);
  not g69872 (n_31134, n41792);
  and g69873 (n41793, n40593, n_31134);
  not g69874 (n_31135, n41793);
  and g69875 (n41794, pi1147, n_31135);
  and g69876 (n41795, n38423, n_29879);
  and g69877 (n41796, n_29898, n40653);
  not g69878 (n_31136, n41795);
  and g69879 (n41797, n_31136, n41796);
  and g69880 (n41798, n_29468, n_29815);
  not g69881 (n_31137, n41797);
  and g69882 (n41799, n_31137, n41798);
  not g69883 (n_31138, n40198);
  and g69884 (n41800, n_31138, n41799);
  not g69885 (n_31139, n41800);
  and g69886 (n41801, n41794, n_31139);
  and g69887 (n41802, n41765, n_31137);
  and g69888 (n41803, n_30143, n41517);
  not g69889 (n_31140, n41803);
  and g69890 (n41804, n40269, n_31140);
  not g69891 (n_31141, n41804);
  and g69892 (n41805, n_29807, n_31141);
  and g69893 (n41806, pi1151, n41805);
  not g69894 (n_31142, n41802);
  and g69895 (n41807, n_29810, n_31142);
  not g69896 (n_31143, n41806);
  and g69897 (n41808, n_31143, n41807);
  not g69898 (n_31144, n41808);
  and g69899 (n41809, pi1149, n_31144);
  not g69900 (n_31145, n41801);
  and g69901 (n41810, n_31145, n41809);
  not g69902 (n_31146, n41789);
  and g69903 (n41811, n_30133, n_31146);
  not g69904 (n_31147, n41810);
  and g69905 (n41812, n_31147, n41811);
  not g69906 (n_31148, n41777);
  not g69907 (n_31149, n41812);
  and g69908 (n41813, n_31148, n_31149);
  not g69909 (n_31150, n41813);
  and g69910 (n41814, pi1148, n_31150);
  and g69911 (n41815, n_29468, n_29938);
  not g69912 (n_31151, n41815);
  and g69913 (n41816, n_29810, n_31151);
  and g69914 (n41817, pi1151, n_29793);
  not g69915 (n_31152, n41817);
  and g69916 (n41818, n41816, n_31152);
  and g69917 (n41819, n_30976, n41746);
  not g69918 (n_31153, n41819);
  and g69919 (n41820, n39870, n_31153);
  not g69920 (n_31154, n41554);
  and g69921 (n41821, n_29646, n_31154);
  and g69922 (n41822, n_29468, n41821);
  not g69923 (n_31155, n41822);
  and g69924 (n41823, pi1147, n_31155);
  not g69925 (n_31156, n41820);
  and g69926 (n41824, n_31156, n41823);
  not g69927 (n_31157, n41818);
  and g69928 (n41825, pi1150, n_31157);
  not g69929 (n_31158, n41824);
  and g69930 (n41826, n_31158, n41825);
  and g69931 (n41827, n_29810, pi1151);
  and g69932 (n41828, n40140, n41827);
  and g69933 (n41829, n_29471, n40664);
  not g69934 (n_31159, n41829);
  and g69935 (n41830, n40696, n_31159);
  not g69936 (n_31160, n41830);
  and g69937 (n41831, n39870, n_31160);
  and g69938 (n41832, n40565, n_30260);
  not g69939 (n_31161, n41832);
  and g69940 (n41833, pi1147, n_31161);
  not g69941 (n_31162, n41831);
  and g69942 (n41834, n_31162, n41833);
  not g69943 (n_31163, n41828);
  and g69944 (n41835, n_30133, n_31163);
  not g69945 (n_31164, n41834);
  and g69946 (n41836, n_31164, n41835);
  not g69947 (n_31165, n41826);
  not g69948 (n_31166, n41836);
  and g69949 (n41837, n_31165, n_31166);
  not g69950 (n_31167, n41837);
  and g69951 (n41838, n_29850, n_31167);
  and g69952 (n41839, n_29468, n_29920);
  not g69953 (n_31168, n40637);
  and g69954 (n41840, n_31168, n41839);
  not g69955 (n_31169, n40159);
  and g69956 (n41841, n_31169, n40269);
  not g69957 (n_31170, n41841);
  and g69958 (n41842, n_29920, n_31170);
  and g69959 (n41843, pi1151, n41842);
  not g69960 (n_31171, n41840);
  and g69961 (n41844, n_29810, n_31171);
  not g69962 (n_31172, n41843);
  and g69963 (n41845, n_31172, n41844);
  and g69964 (n41846, pi1147, n_30227);
  and g69965 (n41847, n_29468, n_29872);
  and g69966 (n41848, n_31138, n41847);
  not g69967 (n_31173, n41848);
  and g69968 (n41849, n41846, n_31173);
  not g69969 (n_31174, n41845);
  and g69970 (n41850, n_30133, n_31174);
  not g69971 (n_31175, n41849);
  and g69972 (n41851, n_31175, n41850);
  and g69973 (n41852, n40548, n40666);
  not g69974 (n_31176, n41852);
  and g69975 (n41853, pi1147, n_31176);
  not g69976 (n_31177, n40197);
  and g69977 (n41854, n_29872, n_31177);
  and g69978 (n41855, n_29468, n41854);
  not g69979 (n_31178, n41855);
  and g69980 (n41856, n41853, n_31178);
  and g69981 (n41857, n_31116, n41839);
  and g69982 (n41858, pi1151, n_29920);
  and g69983 (n41859, n_29981, n41858);
  not g69984 (n_31179, n41859);
  and g69985 (n41860, n_29810, n_31179);
  not g69986 (n_31180, n41857);
  and g69987 (n41861, n_31180, n41860);
  not g69988 (n_31181, n41856);
  and g69989 (n41862, pi1150, n_31181);
  not g69990 (n_31182, n41861);
  and g69991 (n41863, n_31182, n41862);
  not g69992 (n_31183, n41851);
  not g69993 (n_31184, n41863);
  and g69994 (n41864, n_31183, n_31184);
  not g69995 (n_31185, n41864);
  and g69996 (n41865, pi1149, n_31185);
  not g69997 (n_31186, n41838);
  and g69998 (n41866, n_29904, n_31186);
  not g69999 (n_31187, n41865);
  and g70000 (n41867, n_31187, n41866);
  not g70001 (n_31188, n41814);
  not g70002 (n_31189, n41867);
  and g70003 (n41868, n_31188, n_31189);
  not g70004 (n_31190, n41868);
  and g70005 (n41869, n_26557, n_31190);
  not g70006 (n_31191, n41744);
  and g70007 (n41870, pi0209, n_31191);
  not g70008 (n_31192, n41869);
  and g70009 (n41871, n_31192, n41870);
  and g70010 (n41872, n_26557, n_29908);
  and g70011 (n41873, n_31116, n41858);
  and g70012 (n41874, pi1147, n_30266);
  not g70013 (n_31193, n41873);
  and g70014 (n41875, n_31193, n41874);
  and g70015 (n41876, n_4226, n_30300);
  not g70016 (n_31194, n40714);
  and g70017 (n41877, n_31194, n41876);
  not g70018 (n_31195, n41877);
  and g70019 (n41878, n_30120, n_31195);
  and g70020 (n41879, n41816, n41878);
  not g70021 (n_31196, n41879);
  and g70022 (n41880, n_30133, n_31196);
  not g70023 (n_31197, n41875);
  and g70024 (n41881, n_31197, n41880);
  and g70025 (n41882, n40500, n41769);
  and g70026 (n41883, n40523, n_31117);
  not g70027 (n_31198, n41883);
  and g70028 (n41884, pi1147, n_31198);
  not g70029 (n_31199, n41882);
  and g70030 (n41885, n_31199, n41884);
  and g70031 (n41886, n40116, n40123);
  not g70032 (n_31200, n41886);
  and g70033 (n41887, n40500, n_31200);
  not g70034 (n_31201, n41887);
  and g70035 (n41888, n41754, n_31201);
  not g70036 (n_31202, n41885);
  and g70037 (n41889, pi1150, n_31202);
  not g70038 (n_31203, n41888);
  and g70039 (n41890, n_31203, n41889);
  not g70040 (n_31204, n41881);
  not g70041 (n_31205, n41890);
  and g70042 (n41891, n_31204, n_31205);
  not g70043 (n_31206, n41891);
  and g70044 (n41892, n_29850, n_31206);
  and g70045 (n41893, n40565, n_31153);
  not g70046 (n_31207, n41578);
  and g70047 (n41894, n_29872, n_31207);
  and g70048 (n41895, pi1151, n41894);
  not g70049 (n_31208, n41895);
  and g70050 (n41896, n_29810, n_31208);
  not g70051 (n_31209, n41893);
  and g70052 (n41897, n_31209, n41896);
  and g70053 (n41898, n_29814, n41832);
  not g70054 (n_31210, n41898);
  and g70055 (n41899, n41853, n_31210);
  not g70056 (n_31211, n41899);
  and g70057 (n41900, n_30133, n_31211);
  not g70058 (n_31212, n41897);
  and g70059 (n41901, n_31212, n41900);
  and g70060 (n41902, n_29848, n_30273);
  and g70061 (n41903, n_29468, n41902);
  not g70062 (n_31213, n41903);
  and g70063 (n41904, n41761, n_31213);
  and g70064 (n41905, n40577, n_31103);
  not g70065 (n_31214, n40315);
  and g70066 (n41906, n40069, n_31214);
  not g70067 (n_31215, n41906);
  and g70068 (n41907, n40310, n_31215);
  not g70069 (n_31216, n41907);
  and g70070 (n41908, n40593, n_31216);
  not g70071 (n_31217, n41908);
  and g70072 (n41909, n_29810, n_31217);
  not g70073 (n_31218, n41905);
  and g70074 (n41910, n_31218, n41909);
  not g70075 (n_31219, n41904);
  and g70076 (n41911, pi1150, n_31219);
  not g70077 (n_31220, n41910);
  and g70078 (n41912, n_31220, n41911);
  not g70079 (n_31221, n41901);
  not g70080 (n_31222, n41912);
  and g70081 (n41913, n_31221, n_31222);
  not g70082 (n_31223, n41913);
  and g70083 (n41914, pi1149, n_31223);
  not g70084 (n_31224, n41914);
  and g70085 (n41915, pi1148, n_31224);
  not g70086 (n_31225, n41892);
  and g70087 (n41916, n_31225, n41915);
  and g70088 (n41917, n_25711, n39864);
  not g70089 (n_31226, n41917);
  and g70090 (n41918, pi1151, n_31226);
  not g70091 (n_31227, n41918);
  and g70092 (n41919, n41780, n_31227);
  and g70093 (n41920, n40500, n_31137);
  and g70094 (n41921, n40185, n40653);
  not g70095 (n_31228, n41921);
  and g70096 (n41922, n_29842, n_31228);
  and g70097 (n41923, n_29468, n41922);
  not g70098 (n_31229, n41920);
  and g70099 (n41924, pi1147, n_31229);
  not g70100 (n_31230, n41923);
  and g70101 (n41925, n_31230, n41924);
  not g70102 (n_31231, n41919);
  and g70103 (n41926, pi1150, n_31231);
  not g70104 (n_31232, n41925);
  and g70105 (n41927, n_31232, n41926);
  and g70106 (n41928, n40142, n41827);
  and g70107 (n41929, n_29920, n_31168);
  and g70108 (n41930, n_29468, n_30910);
  not g70109 (n_31233, n41930);
  and g70110 (n41931, pi1147, n_31233);
  not g70111 (n_31234, n41929);
  and g70112 (n41932, n_31234, n41931);
  not g70113 (n_31235, n41928);
  and g70114 (n41933, n_30133, n_31235);
  not g70115 (n_31236, n41932);
  and g70116 (n41934, n_31236, n41933);
  not g70117 (n_31237, n41927);
  not g70118 (n_31238, n41934);
  and g70119 (n41935, n_31237, n_31238);
  not g70120 (n_31239, n41935);
  and g70121 (n41936, n_29850, n_31239);
  and g70122 (n41937, n39642, n39830);
  and g70123 (n41938, n_7077, n41937);
  not g70124 (n_31240, n41938);
  and g70125 (n41939, n_31160, n_31240);
  and g70126 (n41940, n40548, n41939);
  and g70127 (n41941, n40565, n_31160);
  not g70128 (n_31241, n41941);
  and g70129 (n41942, n_29810, n_31241);
  not g70130 (n_31242, n41940);
  and g70131 (n41943, n_31242, n41942);
  and g70132 (n41944, n_6791, n_30291);
  and g70133 (n41945, n_30245, n41944);
  not g70134 (n_31243, n41945);
  and g70135 (n41946, n40164, n_31243);
  and g70136 (n41947, n_29871, n41946);
  not g70137 (n_31244, n41947);
  and g70138 (n41948, n40565, n_31244);
  not g70139 (n_31245, n41948);
  and g70140 (n41949, n41846, n_31245);
  not g70141 (n_31246, n41943);
  and g70142 (n41950, n_30133, n_31246);
  not g70143 (n_31247, n41949);
  and g70144 (n41951, n_31247, n41950);
  not g70145 (n_31248, n41937);
  and g70146 (n41952, n40593, n_31248);
  and g70147 (n41953, n_30293, n41952);
  and g70148 (n41954, n40577, n_30293);
  not g70149 (n_31249, n41953);
  and g70150 (n41955, n_29810, n_31249);
  not g70151 (n_31250, n41954);
  and g70152 (n41956, n_31250, n41955);
  not g70153 (n_31251, n41946);
  and g70154 (n41957, n_29848, n_31251);
  and g70155 (n41958, n_29468, n41957);
  not g70156 (n_31252, n41958);
  and g70157 (n41959, n41794, n_31252);
  not g70158 (n_31253, n41956);
  and g70159 (n41960, pi1150, n_31253);
  not g70160 (n_31254, n41959);
  and g70161 (n41961, n_31254, n41960);
  not g70162 (n_31255, n41951);
  not g70163 (n_31256, n41961);
  and g70164 (n41962, n_31255, n_31256);
  not g70165 (n_31257, n41962);
  and g70166 (n41963, pi1149, n_31257);
  not g70167 (n_31258, n41936);
  and g70168 (n41964, n_29904, n_31258);
  not g70169 (n_31259, n41963);
  and g70170 (n41965, n_31259, n41964);
  not g70171 (n_31260, n41916);
  not g70172 (n_31261, n41965);
  and g70173 (n41966, n_31260, n_31261);
  not g70174 (n_31262, n41966);
  and g70175 (n41967, pi0213, n_31262);
  not g70176 (n_31263, n41872);
  and g70177 (n41968, n_26372, n_31263);
  not g70178 (n_31264, n41967);
  and g70179 (n41969, n_31264, n41968);
  not g70180 (n_31265, n41871);
  not g70181 (n_31266, n41969);
  and g70182 (n41970, n_31265, n_31266);
  not g70183 (n_31267, n41970);
  and g70184 (n41971, pi0230, n_31267);
  and g70185 (n41972, n_28510, n_1955);
  not g70186 (n_31268, n41971);
  not g70187 (n_31269, n41972);
  and g70188 (po0404, n_31268, n_31269);
  and g70189 (n41974, n_29468, n_29858);
  and g70190 (n41975, n_29857, n41974);
  not g70191 (n_31270, n41975);
  and g70192 (n41976, pi1152, n_31270);
  and g70193 (n41977, n_30220, n41976);
  and g70194 (n41978, pi1151, n_28873);
  not g70195 (n_31271, n40125);
  and g70196 (n41979, n_31271, n41978);
  not g70197 (n_31272, n41977);
  and g70198 (n41980, n_30133, n_31272);
  not g70199 (n_31273, n41979);
  and g70200 (n41981, n_31273, n41980);
  and g70201 (n41982, pi1151, n40134);
  not g70202 (n_31274, n41982);
  and g70203 (n41983, n_28873, n_31274);
  and g70204 (n41984, n_30226, n41983);
  and g70205 (n41985, pi1152, n_30224);
  and g70206 (n41986, n_29873, n41847);
  not g70207 (n_31275, n41986);
  and g70208 (n41987, n41985, n_31275);
  not g70209 (n_31276, n41984);
  and g70210 (n41988, pi1150, n_31276);
  not g70211 (n_31277, n41987);
  and g70212 (n41989, n_31277, n41988);
  not g70213 (n_31278, n41981);
  not g70214 (n_31279, n41989);
  and g70215 (n41990, n_31278, n_31279);
  and g70216 (n41991, pi0213, n41990);
  and g70217 (n41992, pi1152, n_31250);
  and g70218 (n41993, n_31107, n41992);
  and g70219 (n41994, pi1151, n41750);
  and g70220 (n41995, n_28873, n_31128);
  not g70221 (n_31280, n41994);
  and g70222 (n41996, n_31280, n41995);
  not g70223 (n_31281, n41993);
  and g70224 (n41997, n_30133, n_31281);
  not g70225 (n_31282, n41996);
  and g70226 (n41998, n_31282, n41997);
  and g70227 (n41999, n_31134, n41798);
  not g70228 (n_31283, n41999);
  and g70229 (n42000, n41985, n_31283);
  and g70230 (n42001, pi1151, n_29847);
  and g70231 (n42002, n41762, n42001);
  not g70232 (n_31284, n42002);
  and g70233 (n42003, n_28873, n_31284);
  and g70234 (n42004, n_31139, n42003);
  not g70235 (n_31285, n42004);
  and g70236 (n42005, pi1150, n_31285);
  not g70237 (n_31286, n42000);
  and g70238 (n42006, n_31286, n42005);
  not g70239 (n_31287, n41998);
  and g70240 (n42007, pi1148, n_31287);
  not g70241 (n_31288, n42006);
  and g70242 (n42008, n_31288, n42007);
  and g70243 (n42009, n_29843, n41755);
  not g70244 (n_31289, n42009);
  and g70245 (n42010, n_28873, n_31289);
  and g70246 (n42011, n_31125, n42010);
  and g70247 (n42012, n40523, n_31126);
  not g70248 (n_31290, n42012);
  and g70249 (n42013, pi1152, n_31290);
  and g70250 (n42014, n_31111, n42013);
  not g70251 (n_31291, n42014);
  and g70252 (n42015, n_30133, n_31291);
  not g70253 (n_31292, n42011);
  and g70254 (n42016, n_31292, n42015);
  and g70255 (n42017, n_29468, n41805);
  and g70256 (n42018, pi1152, n_31118);
  not g70257 (n_31293, n42017);
  and g70258 (n42019, n_31293, n42018);
  and g70259 (n42020, n_28873, n_31142);
  and g70260 (n42021, n_31199, n42020);
  not g70261 (n_31294, n42019);
  and g70262 (n42022, pi1150, n_31294);
  not g70263 (n_31295, n42021);
  and g70264 (n42023, n_31295, n42022);
  not g70265 (n_31296, n42023);
  and g70266 (n42024, n_29904, n_31296);
  not g70267 (n_31297, n42016);
  and g70268 (n42025, n_31297, n42024);
  not g70269 (n_31298, n42008);
  not g70270 (n_31299, n42025);
  and g70271 (n42026, n_31298, n_31299);
  not g70272 (n_31300, n42026);
  and g70273 (n42027, pi1149, n_31300);
  and g70274 (n42028, n_28873, n_31171);
  and g70275 (n42029, n_31193, n42028);
  and g70276 (n42030, n_29468, n41842);
  and g70277 (n42031, pi1152, n_31179);
  not g70278 (n_31301, n42030);
  and g70279 (n42032, n_31301, n42031);
  not g70280 (n_31302, n42029);
  and g70281 (n42033, pi1150, n_31302);
  not g70282 (n_31303, n42032);
  and g70283 (n42034, n_31303, n42033);
  and g70284 (n42035, n40243, n41978);
  and g70285 (n42036, n_29468, n_29857);
  and g70286 (n42037, pi1152, n_31152);
  not g70287 (n_31304, n42036);
  and g70288 (n42038, n_31304, n42037);
  not g70289 (n_31305, n42035);
  and g70290 (n42039, n_30133, n_31305);
  not g70291 (n_31306, n42038);
  and g70292 (n42040, n_31306, n42039);
  not g70293 (n_31307, n42034);
  not g70294 (n_31308, n42040);
  and g70295 (n42041, n_31307, n_31308);
  not g70296 (n_31309, n42041);
  and g70297 (n42042, n_29904, n_31309);
  and g70298 (n42043, pi1152, n_31275);
  and g70299 (n42044, n_31176, n42043);
  and g70300 (n42045, pi1151, n41854);
  and g70301 (n42046, n_28873, n_31173);
  not g70302 (n_31310, n42045);
  and g70303 (n42047, n_31310, n42046);
  not g70304 (n_31311, n42044);
  not g70305 (n_31312, n42047);
  and g70306 (n42048, n_31311, n_31312);
  not g70307 (n_31313, n42048);
  and g70308 (n42049, pi1150, n_31313);
  and g70309 (n42050, pi1151, n41821);
  not g70310 (n_31314, n42050);
  and g70311 (n42051, n_31161, n_31314);
  not g70312 (n_31315, n42051);
  and g70313 (n42052, n_28873, n_31315);
  and g70314 (n42053, n_31156, n_31241);
  not g70315 (n_31316, n42053);
  and g70316 (n42054, pi1152, n_31316);
  not g70317 (n_31317, n42052);
  and g70318 (n42055, n_30133, n_31317);
  not g70319 (n_31318, n42054);
  and g70320 (n42056, n_31318, n42055);
  not g70321 (n_31319, n42056);
  and g70322 (n42057, pi1148, n_31319);
  not g70323 (n_31320, n42049);
  and g70324 (n42058, n_31320, n42057);
  not g70325 (n_31321, n42042);
  and g70326 (n42059, n_29850, n_31321);
  not g70327 (n_31322, n42058);
  and g70328 (n42060, n_31322, n42059);
  not g70329 (n_31323, n42027);
  not g70330 (n_31324, n42060);
  and g70331 (n42061, n_31323, n_31324);
  not g70332 (n_31325, n42061);
  and g70333 (n42062, n_26557, n_31325);
  not g70334 (n_31326, n41991);
  and g70335 (n42063, pi0209, n_31326);
  not g70336 (n_31327, n42062);
  and g70337 (n42064, n_31327, n42063);
  and g70338 (n42065, n_26557, n_30905);
  and g70339 (n42066, n41778, n41978);
  and g70340 (n42067, pi1152, n_31227);
  not g70341 (n_31328, n41974);
  and g70342 (n42068, n_31328, n42067);
  not g70343 (n_31329, n42066);
  and g70344 (n42069, n_30133, n_31329);
  not g70345 (n_31330, n42068);
  and g70346 (n42070, n_31330, n42069);
  and g70347 (n42071, n_28873, n_31241);
  and g70348 (n42072, n_31129, n42071);
  and g70349 (n42073, n41847, n41939);
  and g70350 (n42074, pi1152, n_31249);
  not g70351 (n_31331, n42073);
  and g70352 (n42075, n_31331, n42074);
  not g70353 (n_31332, n42072);
  and g70354 (n42076, pi1150, n_31332);
  not g70355 (n_31333, n42075);
  and g70356 (n42077, n_31333, n42076);
  not g70357 (n_31334, n42070);
  and g70358 (n42078, n_29850, n_31334);
  not g70359 (n_31335, n42077);
  and g70360 (n42079, n_31335, n42078);
  and g70361 (n42080, n_29468, n41894);
  and g70362 (n42081, pi1152, n_31217);
  not g70363 (n_31336, n42080);
  and g70364 (n42082, n_31336, n42081);
  and g70365 (n42083, n_28873, n_31107);
  and g70366 (n42084, n_31209, n42083);
  not g70367 (n_31337, n42082);
  and g70368 (n42085, pi1150, n_31337);
  not g70369 (n_31338, n42084);
  and g70370 (n42086, n_31338, n42085);
  and g70371 (n42087, n_31151, n42010);
  not g70372 (n_31339, n41878);
  and g70373 (n42088, n_29468, n_31339);
  not g70374 (n_31340, n42088);
  and g70375 (n42089, pi1152, n_31340);
  and g70376 (n42090, n_31201, n42089);
  not g70377 (n_31341, n42090);
  and g70378 (n42091, n_30133, n_31341);
  not g70379 (n_31342, n42087);
  and g70380 (n42092, n_31342, n42091);
  not g70381 (n_31343, n42086);
  and g70382 (n42093, pi1149, n_31343);
  not g70383 (n_31344, n42092);
  and g70384 (n42094, n_31344, n42093);
  not g70385 (n_31345, n42079);
  and g70386 (n42095, n_29904, n_31345);
  not g70387 (n_31346, n42094);
  and g70388 (n42096, n_31346, n42095);
  and g70389 (n42097, n41755, n_31117);
  not g70390 (n_31347, n42097);
  and g70391 (n42098, n40673, n_31347);
  and g70392 (n42099, pi1152, n_31180);
  and g70393 (n42100, n_31199, n42099);
  not g70394 (n_31348, n42098);
  and g70395 (n42101, n_30133, n_31348);
  not g70396 (n_31349, n42100);
  and g70397 (n42102, n_31349, n42101);
  and g70398 (n42103, pi1151, n41902);
  and g70399 (n42104, n_28873, n_31210);
  not g70400 (n_31350, n42103);
  and g70401 (n42105, n_31350, n42104);
  and g70402 (n42106, n40666, n41847);
  not g70403 (n_31351, n42106);
  and g70404 (n42107, n41985, n_31351);
  not g70405 (n_31352, n42105);
  and g70406 (n42108, pi1150, n_31352);
  not g70407 (n_31353, n42107);
  and g70408 (n42109, n_31353, n42108);
  not g70409 (n_31354, n42109);
  and g70410 (n42110, pi1149, n_31354);
  not g70411 (n_31355, n42102);
  and g70412 (n42111, n_31355, n42110);
  and g70413 (n42112, pi1151, n41922);
  and g70414 (n42113, n_28873, n_31233);
  not g70415 (n_31356, n42112);
  and g70416 (n42114, n_31356, n42113);
  and g70417 (n42115, pi1152, n_31171);
  and g70418 (n42116, n_31229, n42115);
  not g70419 (n_31357, n42116);
  and g70420 (n42117, n_30133, n_31357);
  not g70421 (n_31358, n42114);
  and g70422 (n42118, n_31358, n42117);
  and g70423 (n42119, n_31135, n42043);
  and g70424 (n42120, pi1151, n41957);
  and g70425 (n42121, n_28873, n_31245);
  not g70426 (n_31359, n42120);
  and g70427 (n42122, n_31359, n42121);
  not g70428 (n_31360, n42119);
  and g70429 (n42123, pi1150, n_31360);
  not g70430 (n_31361, n42122);
  and g70431 (n42124, n_31361, n42123);
  not g70432 (n_31362, n42118);
  and g70433 (n42125, n_29850, n_31362);
  not g70434 (n_31363, n42124);
  and g70435 (n42126, n_31363, n42125);
  not g70436 (n_31364, n42111);
  and g70437 (n42127, pi1148, n_31364);
  not g70438 (n_31365, n42126);
  and g70439 (n42128, n_31365, n42127);
  not g70440 (n_31366, n42096);
  and g70441 (n42129, pi0213, n_31366);
  not g70442 (n_31367, n42128);
  and g70443 (n42130, n_31367, n42129);
  not g70444 (n_31368, n42065);
  and g70445 (n42131, n_26372, n_31368);
  not g70446 (n_31369, n42130);
  and g70447 (n42132, n_31369, n42131);
  not g70448 (n_31370, n42064);
  not g70449 (n_31371, n42132);
  and g70450 (n42133, n_31370, n_31371);
  not g70451 (n_31372, n42133);
  and g70452 (n42134, pi0230, n_31372);
  and g70453 (n42135, n_28510, n_1774);
  not g70454 (n_31373, n42134);
  not g70455 (n_31374, n42135);
  and g70456 (po0405, n_31373, n_31374);
  and g70457 (n42137, n_26557, n41990);
  not g70458 (n_31375, n38886);
  and g70459 (n42138, pi0057, n_31375);
  and g70460 (n42139, n_3232, n38886);
  not g70461 (n_31376, n39738);
  and g70462 (n42140, n_31376, n39882);
  and g70463 (n42141, pi0299, n38883);
  not g70464 (n_31377, n42141);
  and g70465 (n42142, n_30275, n_31377);
  not g70466 (n_31378, n42142);
  and g70467 (n42143, n_26565, n_31378);
  not g70468 (n_31379, n42140);
  and g70469 (n42144, pi0212, n_31379);
  not g70470 (n_31380, n42143);
  and g70471 (n42145, n_31380, n42144);
  and g70472 (n42146, pi0214, n_31378);
  and g70473 (n42147, n_26538, n_29876);
  not g70474 (n_31381, n42146);
  and g70475 (n42148, n_31381, n42147);
  not g70476 (n_31382, n42145);
  and g70477 (n42149, n_6791, n_31382);
  not g70478 (n_31383, n42148);
  and g70479 (n42150, n_31383, n42149);
  and g70480 (n42151, n6305, n_30274);
  not g70481 (n_31384, n42150);
  and g70482 (n42152, n_31384, n42151);
  not g70484 (n_31385, n42139);
  and g70488 (n42156, n_29898, n_31377);
  and g70489 (n42157, n_29876, n42156);
  not g70490 (n_31387, n42157);
  and g70491 (n42158, n_26538, n_31387);
  and g70492 (n42159, n_26565, n42156);
  and g70493 (n42160, n_29634, n_29886);
  and g70494 (n42161, pi0214, n_30241);
  not g70495 (n_31388, n42160);
  and g70496 (n42162, n_31388, n42161);
  not g70497 (n_31389, n42162);
  and g70498 (n42163, pi0212, n_31389);
  not g70499 (n_31390, n42159);
  and g70500 (n42164, n_31390, n42163);
  not g70501 (n_31391, n42158);
  not g70502 (n_31392, n42164);
  and g70503 (n42165, n_31391, n_31392);
  not g70504 (n_31393, n42165);
  and g70505 (n42166, n_6791, n_31393);
  and g70506 (n42167, n6305, n_30251);
  not g70507 (n_31394, n42166);
  and g70508 (n42168, n_31394, n42167);
  not g70513 (n_31396, n42138);
  not g70514 (n_31397, n42155);
  and g70515 (n42172, n_31396, n_31397);
  not g70516 (n_31398, n42171);
  and g70517 (n42173, n_31398, n42172);
  not g70518 (n_31399, n42173);
  and g70519 (n42174, n_28873, n_31399);
  and g70520 (n42175, pi0299, n_28900);
  and g70521 (n42176, n_7077, n42175);
  not g70522 (n_31400, n42176);
  and g70523 (n42177, n_28902, n_31400);
  not g70524 (n_31401, n42177);
  and g70525 (n42178, n40083, n_31401);
  not g70526 (n_31402, n42178);
  and g70527 (n42179, n40660, n_31402);
  not g70528 (n_31403, n40291);
  and g70529 (n42180, n_29895, n_31403);
  not g70530 (n_31404, n42180);
  and g70531 (n42181, pi1151, n_31404);
  not g70532 (n_31405, n42179);
  and g70533 (n42182, n_31405, n42181);
  and g70534 (n42183, n40525, n_31377);
  and g70535 (n42184, n_29507, n_31377);
  not g70536 (n_31406, n42184);
  and g70537 (n42185, n_26565, n_31406);
  and g70538 (n42186, n40149, n_30234);
  not g70539 (n_31407, n42185);
  and g70540 (n42187, pi0212, n_31407);
  not g70541 (n_31408, n42186);
  and g70542 (n42188, n_31408, n42187);
  not g70543 (n_31409, n42183);
  and g70544 (n42189, n41516, n_31409);
  not g70545 (n_31410, n42188);
  and g70546 (n42190, n_31410, n42189);
  not g70547 (n_31411, n42190);
  and g70548 (n42191, n_29468, n_31411);
  and g70549 (n42192, n40164, n42191);
  not g70550 (n_31412, n42182);
  and g70551 (n42193, n38922, n_31412);
  not g70552 (n_31413, n42192);
  and g70553 (n42194, n_31413, n42193);
  not g70554 (n_31414, n42194);
  and g70555 (n42195, pi1150, n_31414);
  not g70556 (n_31415, n42174);
  and g70557 (n42196, n_31415, n42195);
  and g70558 (n42197, n_26538, n39736);
  not g70559 (n_31416, n42175);
  and g70560 (n42198, n40062, n_31416);
  not g70561 (n_31417, n42198);
  and g70562 (n42199, pi0212, n_31417);
  and g70563 (n42200, n_30318, n42199);
  and g70569 (n42204, n39694, n_29984);
  not g70570 (n_31420, n42203);
  and g70571 (n42205, n_31420, n42204);
  and g70572 (n42206, n_29468, n41830);
  and g70573 (n42207, n_31376, n_31400);
  and g70574 (n42208, n38885, n39635);
  not g70575 (n_31421, n42207);
  and g70576 (n42209, n_31421, n42208);
  not g70577 (n_31422, n42209);
  and g70583 (n42213, n10843, n40713);
  and g70584 (n42214, n39066, n_29824);
  and g70585 (n42215, n_28757, n40110);
  and g70586 (n42216, pi0211, n40712);
  not g70587 (n_31425, n42215);
  and g70588 (n42217, n38608, n_31425);
  not g70589 (n_31426, n42216);
  and g70590 (n42218, n_31426, n42217);
  not g70591 (n_31427, n42213);
  not g70592 (n_31428, n42214);
  and g70593 (n42219, n_31427, n_31428);
  not g70594 (n_31429, n42218);
  and g70595 (n42220, n_31429, n42219);
  not g70596 (n_31430, n42220);
  and g70597 (n42221, n_6791, n_31430);
  and g70598 (n42222, pi1151, n40123);
  not g70599 (n_31431, n42221);
  and g70600 (n42223, n_31431, n42222);
  and g70601 (n42224, n38888, n_31422);
  not g70602 (n_31432, n42223);
  and g70603 (n42225, n_31432, n42224);
  not g70604 (n_31433, n42212);
  and g70605 (n42226, n_30133, n_31433);
  not g70606 (n_31434, n42225);
  and g70607 (n42227, n_31434, n42226);
  not g70608 (n_31435, n42196);
  not g70609 (n_31436, n42227);
  and g70610 (n42228, n_31435, n_31436);
  not g70611 (n_31437, n42228);
  and g70612 (n42229, pi0213, n_31437);
  not g70613 (n_31438, n42229);
  and g70614 (n42230, n_26372, n_31438);
  not g70615 (n_31439, n42137);
  and g70616 (n42231, n_31439, n42230);
  and g70617 (n42232, pi0213, n39071);
  and g70618 (n42233, n_28788, n_29024);
  and g70619 (n42234, n38675, n_29158);
  and g70620 (n42235, pi0207, n_28774);
  not g70621 (n_31440, n39027);
  and g70622 (n42236, n_31440, n42235);
  and g70623 (n42237, n_25873, n39252);
  not g70624 (n_31441, n42236);
  and g70625 (n42238, pi0208, n_31441);
  not g70626 (n_31442, n42237);
  and g70627 (n42239, n_31442, n42238);
  not g70628 (n_31443, n42234);
  not g70629 (n_31444, n42239);
  and g70630 (n42240, n_31443, n_31444);
  not g70631 (n_31445, n42240);
  and g70632 (n42241, pi0211, n_31445);
  and g70633 (n42242, pi0214, n42241);
  not g70634 (n_31446, n42233);
  not g70635 (n_31447, n42242);
  and g70636 (n42243, n_31446, n_31447);
  not g70637 (n_31448, n42243);
  and g70638 (n42244, n_26538, n_31448);
  not g70639 (n_31449, n42244);
  and g70640 (n42245, n_6791, n_31449);
  and g70641 (n42246, n_7075, n42240);
  not g70642 (n_31450, n42246);
  and g70643 (n42247, n_29042, n_31450);
  not g70644 (n_31451, n42247);
  and g70645 (n42248, pi0214, n_31451);
  and g70646 (n42249, n_7075, n_29024);
  not g70647 (n_31452, n42249);
  and g70648 (n42250, n_26565, n_31452);
  not g70649 (n_31453, n42241);
  and g70650 (n42251, n_31453, n42250);
  not g70651 (n_31454, n42251);
  and g70652 (n42252, pi0212, n_31454);
  not g70653 (n_31455, n42248);
  and g70654 (n42253, n_31455, n42252);
  not g70655 (n_31456, n42253);
  and g70656 (n42254, n42245, n_31456);
  not g70657 (n_31457, n42254);
  and g70658 (n42255, n39031, n_31457);
  not g70659 (n_31458, n42255);
  and g70660 (n42256, n41755, n_31458);
  and g70661 (n42257, n_29024, n39073);
  not g70662 (n_31459, n41978);
  not g70663 (n_31460, n42257);
  and g70664 (n42258, n_31459, n_31460);
  not g70665 (n_31461, n42256);
  not g70666 (n_31462, n42258);
  and g70667 (n42259, n_31461, n_31462);
  and g70668 (n42260, n_28937, n_29675);
  not g70669 (n_31463, n38968);
  and g70670 (n42261, n_31463, n39909);
  not g70671 (n_31464, n42260);
  and g70672 (n42262, n_4226, n_31464);
  not g70673 (n_31465, n42261);
  and g70674 (n42263, n_31465, n42262);
  not g70675 (n_31466, n42263);
  and g70676 (n42264, n41839, n_31466);
  and g70677 (n42265, pi0214, n38953);
  not g70678 (n_31467, n42265);
  and g70679 (n42266, n39014, n_31467);
  not g70680 (n_31468, n42266);
  and g70681 (n42267, n_6791, n_31468);
  and g70682 (n42268, pi0214, n_31463);
  and g70683 (n42269, n_26565, n38953);
  not g70684 (n_31469, n42269);
  and g70685 (n42270, pi0212, n_31469);
  not g70686 (n_31470, n42268);
  and g70687 (n42271, n_31470, n42270);
  not g70688 (n_31471, n42271);
  and g70689 (n42272, n42267, n_31471);
  and g70690 (n42273, n_4226, n_28941);
  not g70691 (n_31472, n42272);
  and g70692 (n42274, n_31472, n42273);
  not g70693 (n_31473, n42274);
  and g70694 (n42275, n40500, n_31473);
  not g70695 (n_31474, n42264);
  and g70696 (n42276, pi1152, n_31474);
  not g70697 (n_31475, n42275);
  and g70698 (n42277, n_31475, n42276);
  not g70699 (n_31476, n42259);
  not g70700 (n_31477, n42277);
  and g70701 (n42278, n_31476, n_31477);
  not g70702 (n_31478, n42278);
  and g70703 (n42279, n_30133, n_31478);
  and g70704 (n42280, n_28511, n42247);
  and g70705 (n42281, pi0219, n_29043);
  not g70706 (n_31479, n42280);
  and g70707 (n42282, n_31479, n42281);
  not g70708 (n_31480, n42282);
  and g70709 (n42283, n_4226, n_31480);
  and g70710 (n42284, pi0212, n_31448);
  and g70711 (n42285, n_26538, n_29024);
  not g70712 (n_31481, n42285);
  and g70713 (n42286, n_6791, n_31481);
  not g70714 (n_31482, n42284);
  and g70715 (n42287, n_31482, n42286);
  not g70716 (n_31483, n42287);
  and g70717 (n42288, n42283, n_31483);
  not g70718 (n_31484, n42288);
  and g70719 (n42289, n40565, n_31484);
  and g70720 (n42290, pi0214, n42240);
  not g70721 (n_31485, n42290);
  and g70722 (n42291, n42252, n_31485);
  not g70723 (n_31486, n42291);
  and g70724 (n42292, n42245, n_31486);
  not g70725 (n_31487, n42292);
  and g70726 (n42293, n42283, n_31487);
  not g70727 (n_31488, n42293);
  and g70728 (n42294, n41745, n_31488);
  not g70729 (n_31489, n42289);
  and g70730 (n42295, n_28873, n_31489);
  not g70731 (n_31490, n42294);
  and g70732 (n42296, n_31490, n42295);
  and g70733 (n42297, pi0212, n_28960);
  not g70734 (n_31491, n42297);
  and g70735 (n42298, n42267, n_31491);
  not g70736 (n_31492, n42298);
  and g70737 (n42299, n38974, n_31492);
  not g70738 (n_31493, n42299);
  and g70739 (n42300, n40593, n_31493);
  and g70740 (n42301, n_28979, n_31470);
  not g70741 (n_31494, n42301);
  and g70742 (n42302, n_26538, n_31494);
  and g70743 (n42303, n_7075, n38966);
  not g70744 (n_31495, n42303);
  and g70745 (n42304, n_28962, n_31495);
  not g70746 (n_31496, n42304);
  and g70747 (n42305, pi0214, n_31496);
  and g70748 (n42306, n_26565, n38968);
  not g70749 (n_31497, n42305);
  and g70750 (n42307, pi0212, n_31497);
  not g70751 (n_31498, n42306);
  and g70752 (n42308, n_31498, n42307);
  not g70753 (n_31499, n42302);
  not g70754 (n_31500, n42308);
  and g70755 (n42309, n_31499, n_31500);
  not g70756 (n_31501, n42309);
  and g70757 (n42310, n_6791, n_31501);
  not g70758 (n_31502, n42310);
  and g70759 (n42311, n38974, n_31502);
  not g70760 (n_31503, n42311);
  and g70761 (n42312, n41847, n_31503);
  not g70762 (n_31504, n42300);
  and g70763 (n42313, pi1152, n_31504);
  not g70764 (n_31505, n42312);
  and g70765 (n42314, n_31505, n42313);
  not g70766 (n_31506, n42296);
  not g70767 (n_31507, n42314);
  and g70768 (n42315, n_31506, n_31507);
  not g70769 (n_31508, n42315);
  and g70770 (n42316, pi1150, n_31508);
  not g70771 (n_31509, n42279);
  not g70772 (n_31510, n42316);
  and g70773 (n42317, n_31509, n_31510);
  not g70774 (n_31511, n42317);
  and g70775 (n42318, n_26557, n_31511);
  not g70776 (n_31512, n42232);
  and g70777 (n42319, pi0209, n_31512);
  not g70778 (n_31513, n42318);
  and g70779 (n42320, n_31513, n42319);
  not g70780 (n_31514, n42231);
  not g70781 (n_31515, n42320);
  and g70782 (n42321, n_31514, n_31515);
  not g70783 (n_31516, n42321);
  and g70784 (n42322, pi0230, n_31516);
  and g70785 (n42323, n_28510, n_1415);
  not g70786 (n_31517, n42322);
  not g70787 (n_31518, n42323);
  and g70788 (po0406, n_31517, n_31518);
  and g70789 (n42325, n2531, n11513);
  not g70790 (n_31519, n42325);
  and g70791 (n42326, n_28494, n_31519);
  not g70792 (n_31520, n42326);
  and g70793 (n42327, n_171, n_31520);
  and g70794 (n42328, n7333, n8966);
  not g70795 (n_31521, n42327);
  not g70796 (n_31522, n42328);
  and g70797 (n42329, n_31521, n_31522);
  and g70802 (n42333, pi0897, n10809);
  not g70803 (n_31526, pi0476);
  and g70804 (n42334, n_31526, n11444);
  not g70805 (n_31527, n42333);
  not g70806 (n_31528, n42334);
  and g70807 (n42335, n_31527, n_31528);
  and g70808 (n42336, n_7045, pi1053);
  and g70809 (n42337, pi0200, pi1039);
  not g70810 (n_31531, n42336);
  and g70811 (n42338, n_7044, n_31531);
  not g70812 (n_31532, n42337);
  and g70813 (n42339, n_31532, n42338);
  not g70814 (n_31533, n42335);
  not g70815 (n_31534, n42339);
  and g70816 (n42340, n_31533, n_31534);
  and g70817 (n42341, pi0251, n42335);
  or g70818 (po0408, n42340, n42341);
  not g70819 (n_31536, n10983);
  and g70820 (n42343, n_31536, n11552);
  and g70821 (n42344, n_3120, n11552);
  and g70822 (n42345, n_3080, n_6604);
  and g70823 (n42346, pi1001, n42345);
  and g70824 (n42347, n6186, n42346);
  and g70825 (n42348, n_3130, n42347);
  and g70826 (n42349, n6380, n42348);
  not g70827 (n_31537, n42349);
  and g70828 (n42350, n_280, n_31537);
  and g70829 (n42351, pi1092, n_3206);
  not g70830 (n_31538, n42350);
  and g70831 (n42352, n_31538, n42351);
  not g70832 (n_31539, n42352);
  and g70833 (n42353, n6392, n_31539);
  and g70834 (n42354, n6391, n42352);
  not g70835 (n_31540, n42353);
  not g70836 (n_31541, n42354);
  and g70837 (n42355, n_31540, n_31541);
  and g70838 (n42356, n6198, n42355);
  not g70839 (n_31542, n42344);
  not g70840 (n_31543, n42356);
  and g70841 (n42357, n_31542, n_31543);
  not g70842 (n_31544, n42357);
  and g70843 (n42358, n6242, n_31544);
  and g70844 (n42359, n_3140, n42355);
  and g70845 (n42360, n6227, n11552);
  not g70846 (n_31545, n42359);
  not g70847 (n_31546, n42360);
  and g70848 (n42361, n_31545, n_31546);
  not g70849 (n_31547, n42361);
  and g70850 (n42362, n_3162, n_31547);
  not g70851 (n_31548, n42358);
  and g70852 (n42363, pi0299, n_31548);
  not g70853 (n_31549, n42362);
  and g70854 (n42364, n_31549, n42363);
  and g70855 (n42365, n6205, n_31544);
  and g70856 (n42366, n_3119, n_31547);
  not g70857 (n_31550, n42365);
  and g70858 (n42367, n_234, n_31550);
  not g70859 (n_31551, n42366);
  and g70860 (n42368, n_31551, n42367);
  not g70861 (n_31552, n42364);
  and g70862 (n42369, n10983, n_31552);
  not g70863 (n_31553, n42368);
  and g70864 (n42370, n_31553, n42369);
  not g70865 (n_31554, n42343);
  and g70866 (n42371, n_9495, n_31554);
  not g70867 (n_31555, n42370);
  and g70868 (n42372, n_31555, n42371);
  and g70869 (n42373, pi0057, n11551);
  not g70875 (n_31556, n42378);
  and g70876 (n42379, n_280, n_31556);
  and g70877 (n42380, n_796, pi1092);
  not g70878 (n_31557, n42379);
  and g70879 (n42381, n_31557, n42380);
  not g70880 (n_31558, n42373);
  and g70881 (n42382, n7643, n_31558);
  not g70882 (n_31559, n42381);
  and g70883 (n42383, n_31559, n42382);
  not g70884 (n_31560, n42372);
  not g70885 (n_31561, n42383);
  and g70886 (po0409, n_31560, n_31561);
  not g70887 (n_31562, n38508);
  and g70888 (n42385, n_8688, n_31562);
  and g70889 (n42386, n_28724, n42385);
  and g70890 (n42387, n_4226, n42386);
  and g70891 (n42388, pi0219, n40080);
  not g70892 (n_31563, n42387);
  not g70893 (n_31564, n42388);
  and g70894 (n42389, n_31563, n_31564);
  not g70895 (n_31565, n42389);
  and g70896 (n42390, pi1153, n_31565);
  not g70897 (n_31566, n42390);
  and g70898 (n42391, n_29468, n_31566);
  and g70899 (n42392, n10844, n38684);
  not g70900 (n_31567, n38570);
  and g70901 (n42393, pi0211, n_31567);
  not g70902 (n_31568, n42392);
  not g70903 (n_31569, n42393);
  and g70904 (n42394, n_31568, n_31569);
  and g70905 (n42395, n_28608, n_28620);
  not g70906 (n_31570, n42395);
  and g70907 (n42396, n38519, n_31570);
  not g70908 (n_31571, n42396);
  and g70909 (n42397, n_4226, n_31571);
  and g70910 (n42398, n42394, n42397);
  not g70911 (n_31572, n11446);
  and g70912 (n42399, n_31572, n39281);
  not g70913 (n_31573, n42399);
  and g70914 (n42400, pi1151, n_31573);
  not g70915 (n_31574, n42398);
  and g70916 (n42401, n_31574, n42400);
  not g70917 (n_31575, n42391);
  not g70918 (n_31576, n42401);
  and g70919 (n42402, n_31575, n_31576);
  not g70920 (n_31577, n42402);
  and g70921 (n42403, n_28873, n_31577);
  and g70922 (n42404, n38519, n39783);
  and g70927 (n42408, n_7385, n_31562);
  and g70928 (n42409, n_28945, n_29634);
  not g70929 (n_31579, n42409);
  and g70930 (n42410, pi1153, n_31579);
  and g70931 (n42411, pi1151, n42408);
  not g70932 (n_31580, n42410);
  and g70933 (n42412, n_31580, n42411);
  not g70934 (n_31581, n42412);
  and g70935 (n42413, n_4226, n_31581);
  not g70936 (n_31582, n42407);
  and g70937 (n42414, n_31582, n42413);
  and g70938 (n42415, n_29468, n10844);
  not g70939 (n_31583, n42415);
  and g70940 (n42416, n_29182, n_31583);
  and g70941 (n42417, po1038, n42416);
  not g70942 (n_31584, n42417);
  and g70943 (n42418, pi1152, n_31584);
  not g70944 (n_31585, n42414);
  and g70945 (n42419, n_31585, n42418);
  not g70946 (n_31586, n42403);
  not g70947 (n_31587, n42419);
  and g70948 (n42420, n_31586, n_31587);
  not g70949 (n_31588, n42420);
  and g70950 (n42421, pi0230, n_31588);
  not g70951 (n_31589, pi0253);
  and g70952 (n42422, n_31589, n_3128);
  not g70953 (n_31590, n42422);
  and g70954 (n42423, po1038, n_31590);
  and g70955 (n42424, pi0211, pi1091);
  and g70956 (n42425, pi1091, n_11757);
  and g70957 (n42426, pi0219, n42425);
  not g70958 (n_31591, n42424);
  not g70959 (n_31592, n42426);
  and g70960 (n42427, n_31591, n_31592);
  and g70961 (n42428, n42423, n42427);
  not g70962 (n_31593, n42394);
  and g70963 (n42429, pi1091, n_31593);
  and g70964 (n42430, n_11757, n_30469);
  and g70965 (n42431, pi1153, n_30485);
  not g70966 (n_31594, n42431);
  and g70967 (n42432, n38519, n_31594);
  not g70968 (n_31595, n42430);
  and g70969 (n42433, n_31595, n42432);
  not g70970 (n_31596, n42429);
  not g70971 (n_31597, n42433);
  and g70972 (n42434, n_31596, n_31597);
  not g70973 (n_31598, n42434);
  and g70974 (n42435, pi0253, n_31598);
  not g70975 (n_31599, n13064);
  and g70976 (n42436, n_31599, n_31580);
  not g70977 (n_31600, n42436);
  and g70978 (n42437, pi1091, n_31600);
  not g70979 (n_31601, n42437);
  and g70980 (n42438, n_31589, n_31601);
  not g70981 (n_31602, n42438);
  and g70982 (n42439, n_4226, n_31602);
  not g70983 (n_31603, n42435);
  and g70984 (n42440, n_31603, n42439);
  not g70985 (n_31604, n42428);
  and g70986 (n42441, pi1151, n_31604);
  not g70987 (n_31605, n42440);
  and g70988 (n42442, n_31605, n42441);
  and g70989 (n42443, pi0253, n_3128);
  and g70990 (n42444, pi0219, pi1091);
  and g70991 (n42445, n_28578, n42444);
  not g70992 (n_31606, n42445);
  and g70993 (n42446, n42423, n_31606);
  and g70994 (n42447, pi0219, n42446);
  and g70995 (n42448, pi1091, pi1153);
  and g70996 (n42449, n42387, n42448);
  not g70997 (n_31607, n42443);
  not g71003 (n_31610, n42442);
  not g71004 (n_31611, n42452);
  and g71005 (n42453, n_31610, n_31611);
  not g71006 (n_31612, n42453);
  and g71007 (n42454, n_28873, n_31612);
  and g71008 (n42455, n_7075, pi1091);
  and g71009 (n42456, n_6791, n42455);
  not g71010 (n_31613, n42456);
  and g71011 (n42457, n42446, n_31613);
  and g71012 (n42458, n11446, n40911);
  and g71013 (n42459, n_28715, n42458);
  and g71014 (n42460, n_11757, n_30480);
  and g71015 (n42461, n_28629, n40911);
  not g71016 (n_31614, n42461);
  and g71017 (n42462, pi1153, n_31614);
  not g71018 (n_31615, n42462);
  and g71019 (n42463, n38519, n_31615);
  not g71020 (n_31616, n42460);
  and g71021 (n42464, n_31616, n42463);
  not g71022 (n_31617, n42459);
  and g71023 (n42465, pi0253, n_31617);
  not g71024 (n_31618, n42464);
  and g71025 (n42466, n_31618, n42465);
  and g71026 (n42467, pi1091, n39783);
  and g71027 (n42468, pi1091, n38545);
  and g71028 (n42469, n38958, n42468);
  not g71029 (n_31619, n42469);
  and g71030 (n42470, n38519, n_31619);
  not g71031 (n_31620, n42467);
  and g71032 (n42471, n_31620, n42470);
  and g71033 (n42472, pi1091, n38688);
  and g71034 (n42473, pi0211, n_30496);
  not g71035 (n_31621, n42472);
  and g71036 (n42474, n_31621, n42473);
  not g71037 (n_31622, n42471);
  and g71038 (n42475, n_31589, n_31622);
  not g71039 (n_31623, n42474);
  and g71040 (n42476, n_31623, n42475);
  not g71041 (n_31624, n42466);
  not g71042 (n_31625, n42476);
  and g71043 (n42477, n_31624, n_31625);
  not g71044 (n_31626, n38519);
  and g71045 (n42478, n_31572, n_31626);
  and g71046 (n42479, n_31607, n42478);
  and g71047 (n42480, n_31621, n42479);
  not g71048 (n_31627, n42480);
  and g71049 (n42481, n39635, n_31627);
  not g71050 (n_31628, n42477);
  and g71051 (n42482, n_31628, n42481);
  and g71052 (n42483, n42409, n_31607);
  not g71053 (n_31629, n42425);
  not g71054 (n_31630, n42483);
  and g71055 (n42484, n_31629, n_31630);
  not g71056 (n_31631, n42484);
  and g71057 (n42485, n42408, n_31631);
  and g71058 (n42486, n_4226, n_31590);
  not g71059 (n_31632, n42485);
  and g71060 (n42487, n_31632, n42486);
  not g71061 (n_31633, n42446);
  not g71062 (n_31634, n42487);
  and g71063 (n42488, n_31633, n_31634);
  not g71064 (n_31635, n42488);
  and g71065 (n42489, pi1151, n_31635);
  not g71072 (n_31639, n42492);
  and g71073 (n42493, n_30644, n_31639);
  not g71074 (n_31640, n42454);
  and g71075 (n42494, n_31640, n42493);
  and g71076 (n42495, n40988, n41072);
  not g71077 (n_31641, n42495);
  and g71078 (n42496, pi1153, n_31641);
  not g71079 (n_31642, n41118);
  and g71080 (n42497, n_11757, n_31642);
  not g71081 (n_31643, n42497);
  and g71082 (n42498, n_6791, n_31643);
  not g71083 (n_31644, n42496);
  and g71084 (n42499, n_31644, n42498);
  and g71085 (n42500, n_11757, n_30563);
  and g71086 (n42501, n_30517, n_30537);
  and g71087 (n42502, n_7075, n41044);
  not g71088 (n_31645, n42502);
  and g71089 (n42503, n42501, n_31645);
  and g71090 (n42504, n41000, n_30535);
  and g71091 (n42505, n42503, n42504);
  not g71092 (n_31646, n42505);
  and g71093 (n42506, pi1153, n_31646);
  not g71094 (n_31647, n42500);
  and g71095 (n42507, pi0219, n_31647);
  not g71096 (n_31648, n42506);
  and g71097 (n42508, n_31648, n42507);
  not g71098 (n_31649, n42499);
  and g71099 (n42509, pi0253, n_31649);
  not g71100 (n_31650, n42508);
  and g71101 (n42510, n_31650, n42509);
  and g71102 (n42511, n_30522, n41048);
  and g71103 (n42512, n_7075, n42511);
  not g71104 (n_31651, n41013);
  not g71105 (n_31652, n42512);
  and g71106 (n42513, n_31651, n_31652);
  not g71107 (n_31653, n42513);
  and g71108 (n42514, pi1153, n_31653);
  not g71109 (n_31654, n41039);
  not g71110 (n_31655, n42514);
  and g71111 (n42515, n_31654, n_31655);
  and g71112 (n42516, pi0219, n42515);
  and g71113 (n42517, n_11757, n41116);
  and g71114 (n42518, pi1153, n41097);
  not g71115 (n_31656, n42517);
  and g71116 (n42519, n_6791, n_31656);
  not g71117 (n_31657, n42518);
  and g71118 (n42520, n_31657, n42519);
  not g71119 (n_31658, n42520);
  and g71120 (n42521, n_31589, n_31658);
  not g71121 (n_31659, n42516);
  and g71122 (n42522, n_31659, n42521);
  not g71123 (n_31660, n42510);
  not g71124 (n_31661, n42522);
  and g71125 (n42523, n_31660, n_31661);
  not g71126 (n_31662, n42523);
  and g71127 (n42524, n_4226, n_31662);
  and g71128 (n42525, n_6791, n_30509);
  and g71129 (n42526, n_7075, n_30436);
  not g71130 (n_31663, n42526);
  and g71131 (n42527, n42525, n_31663);
  not g71132 (n_31664, n42527);
  and g71133 (n42528, n_6791, n_31664);
  and g71134 (n42529, po1038, n42528);
  and g71135 (n42530, n_30508, n42529);
  and g71136 (n42531, n_30521, n_31606);
  not g71137 (n_31665, n42525);
  and g71138 (n42532, n_31665, n42531);
  not g71139 (n_31666, n42532);
  and g71140 (n42533, pi0253, n_31666);
  and g71141 (n42534, n_6791, n_30436);
  and g71142 (n42535, pi0211, n40868);
  and g71143 (n42536, n_7075, n_30508);
  not g71144 (n_31667, n42535);
  and g71145 (n42537, pi0219, n_31667);
  not g71146 (n_31668, n42536);
  and g71147 (n42538, n_31668, n42537);
  not g71148 (n_31669, n42534);
  and g71149 (n42539, n_31606, n_31669);
  not g71150 (n_31670, n42538);
  and g71151 (n42540, n_31670, n42539);
  not g71152 (n_31671, n42540);
  and g71153 (n42541, n_31589, n_31671);
  not g71154 (n_31672, n42533);
  and g71155 (n42542, po1038, n_31672);
  not g71156 (n_31673, n42541);
  and g71157 (n42543, n_31673, n42542);
  not g71158 (n_31674, n42530);
  and g71159 (n42544, pi1151, n_31674);
  not g71160 (n_31675, n42543);
  and g71161 (n42545, n_31675, n42544);
  not g71162 (n_31676, n42524);
  and g71163 (n42546, n_31676, n42545);
  and g71164 (n42547, n_30579, n_31652);
  not g71165 (n_31677, n42547);
  and g71166 (n42548, n42525, n_31677);
  and g71167 (n42549, n_30517, n_30528);
  not g71168 (n_31678, n42549);
  and g71169 (n42550, n_11757, n_31678);
  not g71170 (n_31679, n41102);
  not g71171 (n_31680, n42550);
  and g71172 (n42551, n_31679, n_31680);
  not g71173 (n_31681, n42551);
  and g71174 (n42552, n42548, n_31681);
  and g71175 (n42553, pi0219, n41009);
  and g71176 (n42554, n_30571, n42506);
  not g71177 (n_31682, n42554);
  and g71178 (n42555, n42553, n_31682);
  not g71179 (n_31683, n42552);
  not g71180 (n_31684, n42555);
  and g71181 (n42556, n_31683, n_31684);
  not g71182 (n_31685, n42556);
  and g71183 (n42557, pi0253, n_31685);
  and g71184 (n42558, n_30536, n42503);
  and g71185 (n42559, n_31680, n42558);
  not g71186 (n_31686, n42559);
  and g71187 (n42560, n_6791, n_31686);
  and g71188 (n42561, pi0219, n41011);
  not g71189 (n_31687, n42560);
  not g71190 (n_31688, n42561);
  and g71191 (n42562, n_31687, n_31688);
  and g71192 (n42563, n_31659, n42562);
  not g71193 (n_31689, n42563);
  and g71194 (n42564, n_31589, n_31689);
  not g71195 (n_31690, n42557);
  and g71196 (n42565, n_4226, n_31690);
  not g71197 (n_31691, n42564);
  and g71198 (n42566, n_31691, n42565);
  not g71199 (n_31692, n42566);
  and g71200 (n42567, n_29468, n_31692);
  not g71201 (n_31693, n42546);
  not g71202 (n_31694, n42567);
  and g71203 (n42568, n_31693, n_31694);
  and g71204 (n42569, n42534, n_31668);
  not g71205 (n_31695, n42569);
  and g71206 (n42570, n42525, n_31695);
  and g71207 (n42571, pi0219, n_30508);
  not g71208 (n_31696, n42571);
  and g71209 (n42572, po1038, n_31696);
  not g71210 (n_31697, n42570);
  and g71211 (n42573, n_31697, n42572);
  and g71212 (n42574, n_30508, n42573);
  not g71213 (n_31698, n42574);
  and g71214 (n42575, n_31675, n_31698);
  not g71215 (n_31699, n42568);
  and g71216 (n42576, n_31699, n42575);
  not g71217 (n_31700, n42576);
  and g71218 (n42577, pi1152, n_31700);
  not g71219 (n_31701, n42515);
  and g71220 (n42578, pi0219, n_31701);
  and g71221 (n42579, n_31658, n42548);
  not g71222 (n_31702, n42578);
  not g71223 (n_31703, n42579);
  and g71224 (n42580, n_31702, n_31703);
  not g71225 (n_31704, n42580);
  and g71226 (n42581, n_30522, n_31704);
  not g71227 (n_31705, n42581);
  and g71228 (n42582, n_31589, n_31705);
  and g71229 (n42583, pi1153, n_30518);
  and g71230 (n42584, n42503, n42525);
  not g71231 (n_31706, n42583);
  and g71232 (n42585, n_31706, n42584);
  and g71233 (n42586, n_11757, n_30550);
  not g71234 (n_31707, n41062);
  and g71235 (n42587, n_31707, n_31646);
  and g71236 (n42588, pi1153, n42587);
  not g71237 (n_31708, n42586);
  and g71238 (n42589, pi0219, n_31708);
  not g71239 (n_31709, n42588);
  and g71240 (n42590, n_31709, n42589);
  not g71241 (n_31710, n42585);
  not g71242 (n_31711, n42590);
  and g71243 (n42591, n_31710, n_31711);
  not g71244 (n_31712, n42591);
  and g71245 (n42592, pi0253, n_31712);
  not g71246 (n_31713, n42592);
  and g71247 (n42593, n_4226, n_31713);
  not g71248 (n_31714, n42582);
  and g71249 (n42594, n_31714, n42593);
  not g71250 (n_31715, n42594);
  and g71251 (n42595, n42545, n_31715);
  and g71252 (n42596, n_3128, n_31654);
  not g71253 (n_31716, n42596);
  and g71254 (n42597, n_11757, n_31716);
  and g71255 (n42598, n_30571, n_31646);
  and g71256 (n42599, n_6791, n42549);
  not g71257 (n_31717, n42597);
  not g71258 (n_31718, n42599);
  and g71259 (n42600, n_31717, n_31718);
  and g71260 (n42601, n42598, n42600);
  not g71261 (n_31719, n42601);
  and g71262 (n42602, pi0253, n_31719);
  and g71263 (n42603, n_30530, n42578);
  not g71264 (n_31720, n41084);
  and g71265 (n42604, n_11757, n_31720);
  not g71266 (n_31721, n42604);
  and g71267 (n42605, n_30522, n_31721);
  and g71268 (n42606, n_6791, n41118);
  and g71269 (n42607, n42605, n42606);
  not g71270 (n_31722, n42607);
  and g71271 (n42608, n_31589, n_31722);
  not g71272 (n_31723, n42603);
  and g71273 (n42609, n_31723, n42608);
  not g71274 (n_31724, n42602);
  and g71275 (n42610, n_4226, n_31724);
  not g71276 (n_31725, n42609);
  and g71277 (n42611, n_31725, n42610);
  and g71278 (n42612, n_29468, n_31675);
  not g71279 (n_31726, n42611);
  and g71280 (n42613, n_31726, n42612);
  not g71281 (n_31727, n42613);
  and g71282 (n42614, n_28873, n_31727);
  not g71283 (n_31728, n42595);
  and g71284 (n42615, n_31728, n42614);
  not g71285 (n_31729, n42577);
  not g71286 (n_31730, n42615);
  and g71287 (n42616, n_31729, n_31730);
  not g71288 (n_31731, n42616);
  and g71289 (n42617, n40910, n_31731);
  not g71290 (n_31732, n42494);
  and g71291 (n42618, n_28510, n_31732);
  not g71292 (n_31733, n42617);
  and g71293 (n42619, n_31733, n42618);
  not g71294 (n_31734, n42421);
  not g71295 (n_31735, n42619);
  and g71296 (po0410, n_31734, n_31735);
  and g71297 (n42621, n_6791, n_28870);
  not g71298 (n_31736, n42621);
  and g71299 (n42622, n_29079, n_31736);
  and g71300 (n42623, po1038, n42622);
  and g71301 (n42624, pi1154, n38977);
  not g71302 (n_31737, n42624);
  and g71303 (n42625, n_28991, n_31737);
  not g71304 (n_31738, n42625);
  and g71305 (n42626, n11446, n_31738);
  and g71306 (n42627, pi0299, n38519);
  and g71307 (n42628, n_31572, n38959);
  not g71308 (n_31739, n42627);
  not g71309 (n_31740, n42628);
  and g71310 (n42629, n_31739, n_31740);
  not g71311 (n_31741, n42629);
  and g71312 (n42630, n_28918, n_31741);
  not g71313 (n_31742, n42626);
  not g71314 (n_31743, n42630);
  and g71315 (n42631, n_31742, n_31743);
  not g71316 (n_31744, n42631);
  and g71317 (n42632, n_4226, n_31744);
  not g71318 (n_31745, n42623);
  and g71319 (n42633, n_28873, n_31745);
  not g71320 (n_31746, n42632);
  and g71321 (n42634, n_31746, n42633);
  and g71322 (n42635, n11446, n_28870);
  not g71323 (n_31747, n42635);
  and g71324 (n42636, n40028, n_31747);
  and g71325 (n42637, n_7045, pi1154);
  not g71326 (n_31748, n42637);
  and g71327 (n42638, n11373, n_31748);
  and g71328 (n42639, n38976, n_29634);
  not g71329 (n_31749, n42638);
  not g71330 (n_31750, n42639);
  and g71331 (n42640, n_31749, n_31750);
  not g71332 (n_31751, n42640);
  and g71333 (n42641, n_6791, n_31751);
  and g71334 (n42642, n_28619, n_28946);
  not g71335 (n_31752, n42642);
  and g71336 (n42643, n38488, n_31752);
  and g71337 (n42644, n_11413, n_28986);
  not g71338 (n_31753, n42644);
  and g71339 (n42645, n_28919, n_31753);
  not g71340 (n_31754, n42643);
  and g71341 (n42646, n_31754, n42645);
  not g71342 (n_31755, n42646);
  and g71343 (n42647, pi0219, n_31755);
  not g71344 (n_31756, n42641);
  and g71345 (n42648, n_4226, n_31756);
  not g71346 (n_31757, n42647);
  and g71347 (n42649, n_31757, n42648);
  not g71348 (n_31758, n42636);
  and g71349 (n42650, pi1152, n_31758);
  not g71350 (n_31759, n42649);
  and g71351 (n42651, n_31759, n42650);
  not g71352 (n_31760, n42634);
  not g71353 (n_31761, n42651);
  and g71354 (n42652, n_31760, n_31761);
  not g71355 (n_31762, n42652);
  and g71356 (n42653, pi0230, n_31762);
  not g71357 (n_31763, pi0254);
  and g71358 (n42654, n_31763, n_3128);
  not g71359 (n_31764, n42622);
  and g71360 (n42655, pi1091, n_31764);
  not g71361 (n_31765, n42654);
  and g71362 (n42656, po1038, n_31765);
  not g71363 (n_31766, n42655);
  and g71364 (n42657, n_31766, n42656);
  and g71365 (n42658, po1038, n42456);
  not g71366 (n_31767, n42657);
  not g71367 (n_31768, n42658);
  and g71368 (n42659, n_31767, n_31768);
  and g71369 (n42660, pi1153, n_30471);
  not g71370 (n_31769, n42660);
  and g71371 (n42661, n_11413, n_31769);
  and g71372 (n42662, n_7075, n38683);
  and g71373 (n42663, n_31595, n42661);
  not g71374 (n_31770, n42662);
  and g71375 (n42664, n_31770, n42663);
  not g71379 (n_31771, n42664);
  not g71380 (n_31772, n42667);
  and g71381 (n42668, n_31771, n_31772);
  not g71382 (n_31773, n42668);
  and g71383 (n42669, n_6791, n_31773);
  and g71384 (n42670, pi1154, n42455);
  not g71385 (n_31774, n42444);
  not g71386 (n_31775, n42670);
  and g71387 (n42671, n_31774, n_31775);
  not g71388 (n_31776, n42671);
  and g71389 (n42672, n_31755, n_31776);
  not g71390 (n_31777, n42669);
  not g71391 (n_31778, n42672);
  and g71392 (n42673, n_31777, n_31778);
  not g71393 (n_31779, n42673);
  and g71394 (n42674, pi0254, n_31779);
  and g71395 (n42675, pi1154, n_31579);
  and g71396 (n42676, pi0219, n_28986);
  not g71397 (n_31780, n42675);
  and g71398 (n42677, n_31780, n42676);
  not g71399 (n_31781, n42677);
  and g71400 (n42678, n_31756, n_31781);
  not g71401 (n_31782, n42678);
  and g71402 (n42679, n_31763, n_31782);
  not g71403 (n_31783, n42679);
  and g71404 (n42680, n_31765, n_31783);
  not g71405 (n_31784, n42674);
  and g71406 (n42681, n_31784, n42680);
  and g71407 (n42682, n_4226, n42681);
  and g71408 (n42683, pi1152, n42659);
  not g71409 (n_31785, n42682);
  and g71410 (n42684, n_31785, n42683);
  and g71411 (n42685, n40918, n42425);
  not g71412 (n_31786, n42685);
  and g71413 (n42686, n_31620, n_31786);
  not g71414 (n_31787, n42661);
  and g71415 (n42687, pi0211, n_31787);
  not g71416 (n_31788, n42686);
  and g71417 (n42688, n_31788, n42687);
  and g71418 (n42689, n11445, n42448);
  not g71419 (n_31789, n42689);
  and g71420 (n42690, n_11413, n_31789);
  and g71421 (n42691, pi1091, n38959);
  not g71422 (n_31790, n42691);
  and g71423 (n42692, pi1154, n_31790);
  not g71424 (n_31791, n42690);
  and g71425 (n42693, n_7075, n_31791);
  not g71426 (n_31792, n42692);
  and g71427 (n42694, n_31792, n42693);
  not g71428 (n_31793, n42688);
  not g71429 (n_31794, n42694);
  and g71430 (n42695, n_31793, n_31794);
  not g71431 (n_31795, n42695);
  and g71432 (n42696, n_6791, n_31795);
  and g71433 (n42697, pi0211, n42692);
  and g71434 (n42698, pi1091, n39666);
  not g71435 (n_31796, n42698);
  and g71436 (n42699, n38495, n_31796);
  and g71437 (n42700, n_31620, n42699);
  not g71443 (n_31799, n42696);
  not g71444 (n_31800, n42703);
  and g71445 (n42704, n_31799, n_31800);
  not g71446 (n_31801, n42704);
  and g71447 (n42705, n_31763, n_31801);
  and g71448 (n42706, n_11757, n_30462);
  not g71449 (n_31802, n42706);
  and g71450 (n42707, n_31615, n_31802);
  and g71451 (n42708, pi1091, n_11413);
  and g71452 (n42709, n38533, n42708);
  not g71453 (n_31803, n42707);
  not g71454 (n_31804, n42709);
  and g71455 (n42710, n_31803, n_31804);
  not g71456 (n_31805, n42710);
  and g71457 (n42711, n11446, n_31805);
  and g71458 (n42712, pi1091, n_31572);
  and g71459 (n42713, n_28916, n42712);
  not g71460 (n_31806, n42713);
  and g71461 (n42714, n_11413, n_31806);
  and g71462 (n42715, n40968, n42463);
  and g71463 (n42716, pi1091, n_29326);
  not g71464 (n_31807, n42716);
  and g71465 (n42717, n_31803, n_31807);
  not g71466 (n_31808, n42717);
  and g71467 (n42718, n42478, n_31808);
  not g71468 (n_31809, n42715);
  and g71469 (n42719, pi1154, n_31809);
  not g71470 (n_31810, n42718);
  and g71471 (n42720, n_31810, n42719);
  not g71472 (n_31811, n42714);
  not g71473 (n_31812, n42720);
  and g71474 (n42721, n_31811, n_31812);
  not g71475 (n_31813, n42711);
  and g71476 (n42722, pi0254, n_31813);
  not g71477 (n_31814, n42721);
  and g71478 (n42723, n_31814, n42722);
  not g71479 (n_31815, n42705);
  not g71480 (n_31816, n42723);
  and g71481 (n42724, n_31815, n_31816);
  not g71482 (n_31817, n42724);
  and g71483 (n42725, n_4226, n_31817);
  and g71484 (n42726, n_28873, n_31767);
  not g71485 (n_31818, n42725);
  and g71486 (n42727, n_31818, n42726);
  not g71487 (n_31819, n42684);
  and g71488 (n42728, n_30644, n_31819);
  not g71489 (n_31820, n42727);
  and g71490 (n42729, n_31820, n42728);
  and g71491 (n42730, pi1091, n39145);
  and g71492 (n42731, n_7075, n_30430);
  not g71493 (n_31821, n42731);
  and g71494 (n42732, n42571, n_31821);
  and g71495 (n42733, n_6791, n40890);
  not g71496 (n_31822, n42732);
  not g71497 (n_31823, n42733);
  and g71498 (n42734, n_31822, n_31823);
  and g71499 (n42735, n11446, n42425);
  not g71502 (n_31825, n42730);
  not g71505 (n_31826, n42448);
  and g71506 (n42739, n_31826, n42569);
  not g71511 (n_31828, n42738);
  and g71512 (n42743, pi0253, n_31828);
  not g71513 (n_31829, n42742);
  and g71514 (n42744, n_31829, n42743);
  and g71515 (n42745, pi0253, po1038);
  not g71516 (n_31830, n42745);
  and g71517 (n42746, n42659, n_31830);
  not g71518 (n_31831, n42744);
  not g71519 (n_31832, n42746);
  and g71520 (n42747, n_31831, n_31832);
  not g71521 (n_31833, n42681);
  and g71522 (n42748, n_31589, n_31833);
  and g71523 (n42749, pi1154, n_30516);
  and g71524 (n42750, n42503, n42749);
  and g71525 (n42751, n_31644, n42750);
  and g71526 (n42752, n_11757, n42559);
  not g71527 (n_31834, n42752);
  and g71528 (n42753, n_31642, n_31834);
  not g71529 (n_31835, n42753);
  and g71530 (n42754, n_11413, n_31835);
  not g71531 (n_31836, n42751);
  and g71532 (n42755, pi0254, n_31836);
  not g71533 (n_31837, n42754);
  and g71534 (n42756, n_31837, n42755);
  and g71535 (n42757, pi0211, n41044);
  not g71536 (n_31838, n42757);
  and g71537 (n42758, n_30522, n_31838);
  not g71538 (n_31839, n42758);
  and g71539 (n42759, n_11757, n_31839);
  and g71540 (n42760, n_30536, n41028);
  and g71541 (n42761, pi1154, n42760);
  not g71542 (n_31840, n42761);
  and g71543 (n42762, n_30612, n_31840);
  not g71544 (n_31841, n42759);
  and g71545 (n42763, n_31763, n_31841);
  not g71546 (n_31842, n42762);
  and g71547 (n42764, n_31842, n42763);
  not g71548 (n_31843, n42756);
  not g71549 (n_31844, n42764);
  and g71550 (n42765, n_31843, n_31844);
  not g71551 (n_31845, n42765);
  and g71552 (n42766, n_6791, n_31845);
  and g71553 (n42767, pi1154, n_31648);
  not g71554 (n_31846, n42587);
  and g71555 (n42768, n_31846, n42767);
  and g71556 (n42769, pi1153, n_30563);
  and g71557 (n42770, n_11413, n_31708);
  not g71558 (n_31847, n42769);
  and g71559 (n42771, n_31847, n42770);
  not g71560 (n_31848, n42771);
  and g71561 (n42772, pi0254, n_31848);
  not g71562 (n_31849, n42768);
  and g71563 (n42773, n_31849, n42772);
  and g71564 (n42774, n_31647, n42760);
  not g71565 (n_31850, n42774);
  and g71566 (n42775, n38495, n_31850);
  and g71567 (n42776, n_30520, n42775);
  and g71568 (n42777, n_11757, n_30554);
  not g71569 (n_31851, n42777);
  and g71570 (n42778, n41041, n_31851);
  not g71571 (n_31852, n42778);
  and g71572 (n42779, n_11413, n_31852);
  and g71573 (n42780, n_30522, n41039);
  not g71574 (n_31853, n42780);
  and g71575 (n42781, n42779, n_31853);
  and g71576 (n42782, pi1153, n41013);
  not g71577 (n_31854, n40995);
  and g71578 (n42783, n38488, n_31854);
  not g71579 (n_31855, n42782);
  and g71580 (n42784, n_31855, n42783);
  not g71587 (n_31859, n42773);
  not g71588 (n_31860, n42787);
  and g71589 (n42788, n_31859, n_31860);
  not g71590 (n_31861, n42788);
  and g71591 (n42789, pi0219, n_31861);
  not g71592 (n_31862, n42789);
  and g71593 (n42790, pi0253, n_31862);
  not g71594 (n_31863, n42766);
  and g71595 (n42791, n_31863, n42790);
  not g71596 (n_31864, n42748);
  and g71597 (n42792, n_4226, n_31864);
  not g71598 (n_31865, n42791);
  and g71599 (n42793, n_31865, n42792);
  not g71600 (n_31866, n42747);
  and g71601 (n42794, pi1152, n_31866);
  not g71602 (n_31867, n42793);
  and g71603 (n42795, n_31867, n42794);
  and g71604 (n42796, n_31767, n_31830);
  and g71605 (n42797, n_31697, n42738);
  not g71606 (n_31868, n42528);
  and g71607 (n42798, n_31868, n42742);
  not g71608 (n_31869, n42797);
  and g71609 (n42799, pi0253, n_31869);
  not g71610 (n_31870, n42798);
  and g71611 (n42800, n_31870, n42799);
  not g71612 (n_31871, n42796);
  not g71613 (n_31872, n42800);
  and g71614 (n42801, n_31871, n_31872);
  and g71615 (n42802, n_31589, n42724);
  and g71616 (n42803, n38495, n_30571);
  and g71617 (n42804, n_11757, n41000);
  not g71618 (n_31873, n41003);
  and g71619 (n42805, n_11413, n_31873);
  not g71620 (n_31874, n42805);
  and g71621 (n42806, n_11413, n_31874);
  not g71622 (n_31875, n42504);
  not g71623 (n_31876, n42804);
  and g71624 (n42807, n_31875, n_31876);
  not g71625 (n_31877, n42806);
  and g71626 (n42808, n_31877, n42807);
  not g71627 (n_31878, n42803);
  and g71628 (n42809, pi0219, n_31878);
  not g71629 (n_31879, n42808);
  and g71630 (n42810, n_31879, n42809);
  and g71631 (n42811, pi1154, n40999);
  and g71632 (n42812, n42547, n_31876);
  not g71633 (n_31880, n42811);
  and g71634 (n42813, n_6791, n_31880);
  not g71635 (n_31881, n42812);
  and g71636 (n42814, n_31881, n42813);
  not g71637 (n_31882, n42810);
  not g71638 (n_31883, n42814);
  and g71639 (n42815, n_31882, n_31883);
  not g71640 (n_31884, n42815);
  and g71641 (n42816, pi0254, n_31884);
  and g71642 (n42817, n41014, n_31647);
  not g71643 (n_31885, n42817);
  and g71644 (n42818, n38488, n_31885);
  and g71651 (n42822, pi1154, n41011);
  not g71652 (n_31889, n42822);
  and g71653 (n42823, n_30562, n_31889);
  not g71654 (n_31890, n42823);
  and g71655 (n42824, n_7075, n_31890);
  and g71656 (n42825, n_30516, n41116);
  and g71657 (n42826, n_31721, n42825);
  not g71658 (n_31891, n42826);
  and g71659 (n42827, n_11413, n_31891);
  and g71660 (n42828, n_30522, n41118);
  not g71661 (n_31892, n42828);
  and g71662 (n42829, pi1154, n_31892);
  and g71663 (n42830, n_31891, n42829);
  not g71670 (n_31896, n42833);
  and g71671 (n42834, n_31763, n_31896);
  not g71672 (n_31897, n42821);
  and g71673 (n42835, n_31897, n42834);
  not g71674 (n_31898, n42816);
  not g71675 (n_31899, n42835);
  and g71676 (n42836, n_31898, n_31899);
  not g71677 (n_31900, n42836);
  and g71678 (n42837, pi0253, n_31900);
  not g71679 (n_31901, n42802);
  and g71680 (n42838, n_4226, n_31901);
  not g71681 (n_31902, n42837);
  and g71682 (n42839, n_31902, n42838);
  not g71683 (n_31903, n42801);
  and g71684 (n42840, n_28873, n_31903);
  not g71685 (n_31904, n42839);
  and g71686 (n42841, n_31904, n42840);
  not g71687 (n_31905, n42841);
  and g71688 (n42842, n40910, n_31905);
  not g71689 (n_31906, n42795);
  and g71690 (n42843, n_31906, n42842);
  not g71691 (n_31907, n42729);
  and g71692 (n42844, n_28510, n_31907);
  not g71693 (n_31908, n42843);
  and g71694 (n42845, n_31908, n42844);
  not g71695 (n_31909, n42653);
  not g71696 (n_31910, n42845);
  and g71697 (po0411, n_31909, n_31910);
  and g71698 (n42847, n_7045, pi1049);
  and g71699 (n42848, pi0200, pi1036);
  not g71700 (n_31913, n42847);
  not g71701 (n_31914, n42848);
  and g71702 (n42849, n_31913, n_31914);
  and g71703 (n42850, n_31533, n42849);
  not g71704 (n_31916, pi0255);
  and g71705 (n42851, n_31916, n42335);
  not g71706 (n_31917, n42850);
  not g71707 (n_31918, n42851);
  and g71708 (po0412, n_31917, n_31918);
  and g71709 (n42853, n_7045, pi1048);
  and g71710 (n42854, pi0200, pi1070);
  not g71711 (n_31921, n42853);
  not g71712 (n_31922, n42854);
  and g71713 (n42855, n_31921, n_31922);
  and g71714 (n42856, n_31533, n42855);
  not g71715 (n_31924, pi0256);
  and g71716 (n42857, n_31924, n42335);
  not g71717 (n_31925, n42856);
  not g71718 (n_31926, n42857);
  and g71719 (po0413, n_31925, n_31926);
  and g71720 (n42859, n_7045, pi1084);
  and g71721 (n42860, pi0200, pi1065);
  not g71722 (n_31929, n42859);
  not g71723 (n_31930, n42860);
  and g71724 (n42861, n_31929, n_31930);
  and g71725 (n42862, n_31533, n42861);
  not g71726 (n_31932, pi0257);
  and g71727 (n42863, n_31932, n42335);
  not g71728 (n_31933, n42862);
  not g71729 (n_31934, n42863);
  and g71730 (po0414, n_31933, n_31934);
  and g71731 (n42865, n_7045, pi1072);
  and g71732 (n42866, pi0200, pi1062);
  not g71733 (n_31937, n42865);
  not g71734 (n_31938, n42866);
  and g71735 (n42867, n_31937, n_31938);
  and g71736 (n42868, n_31533, n42867);
  not g71737 (n_31940, pi0258);
  and g71738 (n42869, n_31940, n42335);
  not g71739 (n_31941, n42868);
  not g71740 (n_31942, n42869);
  and g71741 (po0415, n_31941, n_31942);
  and g71742 (n42871, n_7045, pi1059);
  and g71743 (n42872, pi0200, pi1069);
  not g71744 (n_31945, n42871);
  not g71745 (n_31946, n42872);
  and g71746 (n42873, n_31945, n_31946);
  and g71747 (n42874, n_31533, n42873);
  not g71748 (n_31948, pi0259);
  and g71749 (n42875, n_31948, n42335);
  not g71750 (n_31949, n42874);
  not g71751 (n_31950, n42875);
  and g71752 (po0416, n_31949, n_31950);
  and g71753 (n42877, n_7045, pi1044);
  and g71754 (n42878, pi0200, pi1067);
  not g71755 (n_31953, n42877);
  and g71756 (n42879, n_7044, n_31953);
  not g71757 (n_31954, n42878);
  and g71758 (n42880, n_31954, n42879);
  not g71759 (n_31955, n42880);
  and g71760 (n42881, n_31533, n_31955);
  and g71761 (n42882, pi0260, n42335);
  or g71762 (po0417, n42881, n42882);
  and g71763 (n42884, n_7045, pi1037);
  and g71764 (n42885, pi0200, pi1040);
  not g71765 (n_31959, n42884);
  and g71766 (n42886, n_7044, n_31959);
  not g71767 (n_31960, n42885);
  and g71768 (n42887, n_31960, n42886);
  not g71769 (n_31961, n42887);
  and g71770 (n42888, n_31533, n_31961);
  and g71771 (n42889, pi0261, n42335);
  or g71772 (po0418, n42888, n42889);
  and g71773 (n42891, pi1093, pi1142);
  and g71774 (n42892, n_1323, n_3206);
  not g71775 (n_31963, n42891);
  not g71776 (n_31964, n42892);
  and g71777 (n42893, n_31963, n_31964);
  not g71778 (n_31965, n42893);
  and g71779 (n42894, n_188, n_31965);
  not g71780 (n_31967, pi0123);
  and g71781 (n42895, n_31967, n_1311);
  and g71782 (n42896, pi0123, pi0262);
  not g71783 (n_31968, n42895);
  and g71784 (n42897, pi0228, n_31968);
  not g71785 (n_31969, n42896);
  and g71786 (n42898, n_31969, n42897);
  not g71787 (n_31970, n42894);
  not g71788 (n_31971, n42898);
  and g71789 (n42899, n_31970, n_31971);
  and g71790 (n42900, n_188, n_3206);
  and g71791 (n42901, pi0123, pi0228);
  not g71792 (n_31972, n42900);
  not g71793 (n_31973, n42901);
  and g71794 (n42902, n_31972, n_31973);
  not g71795 (n_31974, n42902);
  and g71796 (n42903, n_1323, n_31974);
  not g71797 (n_31975, n40700);
  not g71798 (n_31976, n42903);
  and g71799 (n42904, n_31975, n_31976);
  and g71800 (n42905, pi0199, n42902);
  not g71801 (n_31977, n42905);
  and g71802 (n42906, n38441, n_31977);
  not g71803 (n_31978, n42906);
  and g71804 (n42907, n42904, n_31978);
  not g71805 (n_31979, n42899);
  not g71806 (n_31980, n42907);
  and g71807 (n42908, n_31979, n_31980);
  and g71808 (n42909, n_25873, n42903);
  not g71809 (n_31981, n42909);
  and g71810 (n42910, n_26242, n_31981);
  not g71811 (n_31982, n42910);
  and g71812 (n42911, n_31975, n_31982);
  not g71813 (n_31983, n42908);
  not g71814 (n_31984, n42911);
  and g71815 (n42912, n_31983, n_31984);
  and g71816 (n42913, n_29527, n42902);
  not g71817 (n_31985, n42913);
  and g71818 (n42914, n_234, n_31985);
  and g71819 (n42915, n_31979, n42914);
  not g71820 (n_31986, n42904);
  and g71821 (n42916, pi0299, n_31986);
  not g71822 (n_31987, n42915);
  and g71823 (n42917, pi0208, n_31987);
  not g71824 (n_31988, n42916);
  and g71825 (n42918, n_31988, n42917);
  not g71826 (n_31989, n42918);
  and g71827 (n42919, n_4226, n_31989);
  not g71828 (n_31990, n42912);
  and g71829 (n42920, n_31990, n42919);
  not g71830 (n_31991, n39864);
  and g71831 (n42921, n_31991, n42902);
  and g71832 (n42922, po1038, n_31979);
  not g71833 (n_31992, n42921);
  and g71834 (n42923, n_31992, n42922);
  or g71835 (po0419, n42920, n42923);
  not g71836 (n_31993, n42708);
  and g71837 (n42925, n_30469, n_31993);
  and g71838 (n42926, n_11794, n_28628);
  not g71839 (n_31994, n42925);
  and g71840 (n42927, n_31994, n42926);
  and g71841 (n42928, pi1155, n_28953);
  not g71842 (n_31995, n42928);
  and g71843 (n42929, n40952, n_31995);
  and g71844 (n42930, n_11413, n42716);
  not g71845 (n_31996, n42929);
  not g71846 (n_31997, n42930);
  and g71847 (n42931, n_31996, n_31997);
  and g71848 (n42932, n_30496, n42931);
  not g71849 (n_31998, n42932);
  and g71850 (n42933, n38479, n_31998);
  and g71851 (n42934, n_11413, n_28727);
  and g71852 (n42935, n38545, n_28636);
  not g71853 (n_31999, n42935);
  and g71854 (n42936, pi1154, n_31999);
  not g71866 (n_32005, n42931);
  and g71867 (n42943, n_7075, n_32005);
  not g71868 (n_32006, n39111);
  and g71869 (n42944, n38568, n_32006);
  not g71870 (n_32007, n42944);
  and g71871 (n42945, n42424, n_32007);
  and g71872 (n42946, n_28773, n42945);
  not g71873 (n_32008, n42943);
  not g71874 (n_32009, n42946);
  and g71875 (n42947, n_32008, n_32009);
  not g71876 (n_32010, n42947);
  and g71877 (n42948, pi1156, n_32010);
  and g71878 (n42949, n_28773, n_31994);
  and g71879 (n42950, pi0211, n42949);
  and g71880 (n42951, n_28628, n_28967);
  and g71881 (n42952, n42455, n42951);
  not g71882 (n_32011, n42950);
  not g71883 (n_32012, n42952);
  and g71884 (n42953, n_32011, n_32012);
  not g71885 (n_32013, n42953);
  and g71886 (n42954, n_11794, n_32013);
  not g71887 (n_32014, n42954);
  and g71888 (n42955, n_6791, n_32014);
  not g71889 (n_32015, n42948);
  and g71890 (n42956, n_32015, n42955);
  not g71891 (n_32016, n42942);
  not g71892 (n_32017, n42956);
  and g71893 (n42957, n_32016, n_32017);
  not g71894 (n_32018, n42957);
  and g71895 (n42958, n_30417, n_32018);
  and g71896 (n42959, n_11413, n38646);
  and g71897 (n42960, pi1154, n_28637);
  not g71898 (n_32019, n42960);
  and g71899 (n42961, pi1156, n_32019);
  not g71900 (n_32020, n42961);
  and g71901 (n42962, n_234, n_32020);
  not g71902 (n_32021, n42959);
  and g71903 (n42963, n_29634, n_32021);
  not g71904 (n_32022, n42962);
  and g71905 (n42964, n_32022, n42963);
  not g71906 (n_32023, n42964);
  and g71907 (n42965, pi1156, n_32023);
  not g71908 (n_32024, n42951);
  and g71909 (n42966, n_32024, n42962);
  not g71910 (n_32025, n42966);
  and g71911 (n42967, pi0219, n_32025);
  not g71912 (n_32026, n42965);
  and g71913 (n42968, n_32026, n42967);
  and g71914 (n42969, n_28680, n39499);
  not g71915 (n_32027, n42969);
  and g71916 (n42970, n_28967, n_32027);
  not g71917 (n_32028, n42970);
  and g71918 (n42971, n_7075, n_32028);
  and g71919 (n42972, n_11794, n42949);
  and g71920 (n42973, n_28945, n_28640);
  not g71921 (n_32029, n42973);
  and g71922 (n42974, pi1154, n_32029);
  and g71923 (n42975, n_28609, n42934);
  not g71924 (n_32030, n42974);
  and g71925 (n42976, pi1156, n_32030);
  not g71926 (n_32031, n42975);
  and g71927 (n42977, n_32031, n42976);
  not g71928 (n_32032, n42972);
  and g71929 (n42978, pi0211, n_32032);
  not g71930 (n_32033, n42977);
  and g71931 (n42979, n_32033, n42978);
  not g71932 (n_32034, n42971);
  and g71933 (n42980, n_6791, n_32034);
  not g71934 (n_32035, n42979);
  and g71935 (n42981, n_32035, n42980);
  not g71941 (n_32038, n42958);
  not g71942 (n_32039, n42984);
  and g71943 (n42985, n_32038, n_32039);
  and g71944 (n42986, n_4226, n42985);
  and g71945 (n42987, pi0219, n_28566);
  and g71946 (n42988, n_6791, n_28567);
  and g71947 (n42989, n_28577, n42988);
  not g71948 (n_32040, n42987);
  not g71949 (n_32041, n42989);
  and g71950 (n42990, n_32040, n_32041);
  not g71951 (n_32042, n42990);
  and g71952 (n42991, pi1091, n_32042);
  and g71953 (n42992, pi0263, n_3128);
  not g71954 (n_32043, n42991);
  not g71955 (n_32044, n42992);
  and g71956 (n42993, n_32043, n_32044);
  not g71957 (n_32045, n42993);
  and g71958 (n42994, po1038, n_32045);
  not g71959 (n_32046, n42994);
  and g71960 (n42995, n_30644, n_32046);
  not g71961 (n_32047, n42986);
  and g71962 (n42996, n_32047, n42995);
  and g71963 (n42997, pi1091, n42987);
  and g71964 (n42998, pi0211, n40874);
  and g71965 (n42999, n_7075, n_31993);
  not g71966 (n_32048, n42999);
  and g71967 (n43000, n_28567, n_32048);
  not g71968 (n_32049, n42998);
  and g71969 (n43001, n_32049, n43000);
  not g71970 (n_32050, n43001);
  and g71971 (n43002, n_30436, n_32050);
  not g71972 (n_32051, n43002);
  and g71973 (n43003, n_6791, n_32051);
  and g71974 (n43004, n_30417, n_31822);
  not g71975 (n_32052, n43003);
  and g71976 (n43005, n_32052, n43004);
  and g71977 (n43006, n_28567, n_31775);
  not g71978 (n_32053, n43006);
  and g71979 (n43007, n_32049, n_32053);
  not g71980 (n_32054, n43007);
  and g71981 (n43008, n42534, n_32054);
  and g71982 (n43009, pi0263, n_31670);
  not g71983 (n_32055, n43008);
  and g71984 (n43010, n_32055, n43009);
  not g71985 (n_32056, n43005);
  not g71986 (n_32057, n43010);
  and g71987 (n43011, n_32056, n_32057);
  not g71988 (n_32058, n42997);
  and g71989 (n43012, n40860, n_32058);
  not g71990 (n_32059, n43011);
  and g71991 (n43013, n_32059, n43012);
  not g71992 (n_32060, n40860);
  and g71993 (n43014, n_32060, n42993);
  not g71994 (n_32061, n43014);
  and g71995 (n43015, po1038, n_32061);
  not g71996 (n_32062, n43013);
  and g71997 (n43016, n_32062, n43015);
  not g71998 (n_32063, n42985);
  and g71999 (n43017, n_32060, n_32063);
  and g72000 (n43018, pi1155, n_31642);
  not g72001 (n_32064, n43018);
  and g72002 (n43019, pi1154, n_32064);
  and g72003 (n43020, n41105, n43019);
  and g72004 (n43021, n_11768, n42596);
  not g72005 (n_32065, n41009);
  and g72006 (n43022, pi1155, n_32065);
  not g72007 (n_32066, n43022);
  and g72008 (n43023, n_11413, n_32066);
  not g72009 (n_32067, n43021);
  and g72010 (n43024, n_32067, n43023);
  and g72011 (n43025, n_30612, n43021);
  and g72012 (n43026, pi1155, n_30579);
  not g72013 (n_32068, n43026);
  and g72014 (n43027, n_11413, n_32068);
  not g72015 (n_32069, n43025);
  and g72016 (n43028, n_32069, n43027);
  not g72017 (n_32070, n43028);
  and g72018 (n43029, n_11794, n_32070);
  not g72019 (n_32071, n43020);
  not g72020 (n_32072, n43024);
  and g72021 (n43030, n_32071, n_32072);
  and g72022 (n43031, n43029, n43030);
  and g72023 (n43032, n_11768, n41000);
  and g72024 (n43033, n_30562, n41102);
  not g72025 (n_32073, n43032);
  not g72026 (n_32074, n43033);
  and g72027 (n43034, n_32073, n_32074);
  not g72028 (n_32075, n43034);
  and g72029 (n43035, n_11413, n_32075);
  not g72030 (n_32076, n43035);
  and g72031 (n43036, pi1156, n_32076);
  and g72032 (n43037, n41000, n43023);
  and g72033 (n43038, n_30514, n43020);
  not g72034 (n_32077, n43037);
  not g72035 (n_32078, n43038);
  and g72036 (n43039, n_32077, n_32078);
  and g72037 (n43040, n43036, n43039);
  not g72038 (n_32079, n43031);
  and g72039 (n43041, n_7075, n_32079);
  not g72040 (n_32080, n43040);
  and g72041 (n43042, n_32080, n43041);
  and g72042 (n43043, n40988, n43019);
  not g72043 (n_32081, n43043);
  and g72044 (n43044, n43036, n_32081);
  and g72045 (n43045, n42501, n43019);
  not g72046 (n_32082, n43045);
  and g72047 (n43046, n43029, n_32082);
  not g72048 (n_32083, n43044);
  and g72049 (n43047, pi0211, n_32083);
  not g72050 (n_32084, n43046);
  and g72051 (n43048, n_32084, n43047);
  not g72052 (n_32085, n43042);
  and g72053 (n43049, n_6791, n_32085);
  not g72054 (n_32086, n43048);
  and g72055 (n43050, n_32086, n43049);
  and g72056 (n43051, pi1155, n41008);
  and g72057 (n43052, pi1154, n41028);
  not g72058 (n_32087, n43051);
  and g72059 (n43053, n_32087, n43052);
  and g72060 (n43054, n_30516, n43053);
  not g72061 (n_32088, n43054);
  and g72062 (n43055, n_32077, n_32088);
  not g72063 (n_32089, n43055);
  and g72064 (n43056, n38479, n_32089);
  not g72065 (n_32090, n43053);
  and g72066 (n43057, n_32072, n_32090);
  not g72067 (n_32091, n43057);
  and g72068 (n43058, n_11794, n_32091);
  and g72069 (n43059, n_11413, n41039);
  not g72070 (n_32092, n43059);
  and g72071 (n43060, n_31707, n_32092);
  and g72072 (n43061, n38483, n_32087);
  not g72073 (n_32093, n43060);
  and g72074 (n43062, n_32093, n43061);
  not g72081 (n_32097, n43065);
  and g72082 (n43066, n_30417, n_32097);
  not g72083 (n_32098, n43050);
  and g72084 (n43067, n_32098, n43066);
  and g72085 (n43068, n_30559, n_30570);
  not g72086 (n_32099, n43068);
  and g72087 (n43069, pi1154, n_32099);
  not g72088 (n_32100, n42760);
  and g72089 (n43070, pi1155, n_32100);
  not g72090 (n_32101, n42511);
  and g72091 (n43071, n_11768, n_32101);
  not g72092 (n_32102, n43070);
  and g72093 (n43072, n_11413, n_32102);
  not g72094 (n_32103, n43071);
  and g72095 (n43073, n_32103, n43072);
  not g72096 (n_32104, n43069);
  and g72097 (n43074, n38483, n_32104);
  not g72098 (n_32105, n43073);
  and g72099 (n43075, n_32105, n43074);
  and g72100 (n43076, n_30538, n_31889);
  not g72101 (n_32106, n43076);
  and g72102 (n43077, n_32099, n_32106);
  not g72103 (n_32107, n43077);
  and g72104 (n43078, n38479, n_32107);
  and g72105 (n43079, n_30549, n43077);
  not g72106 (n_32108, n43079);
  and g72107 (n43080, n_11794, n_32108);
  and g72114 (n43084, pi1154, n_30599);
  not g72115 (n_32112, n41046);
  and g72116 (n43085, n_32112, n43084);
  and g72117 (n43086, n_11413, n_30591);
  and g72118 (n43087, pi1155, n42825);
  not g72119 (n_32113, n43087);
  and g72120 (n43088, n43086, n_32113);
  not g72121 (n_32114, n41114);
  and g72122 (n43089, n_32114, n43084);
  and g72123 (n43090, n_11794, n_31880);
  not g72124 (n_32115, n43089);
  and g72125 (n43091, n_32115, n43090);
  not g72126 (n_32116, n43091);
  and g72127 (n43092, n_11794, n_32116);
  not g72128 (n_32117, n43088);
  not g72129 (n_32118, n43092);
  and g72130 (n43093, n_32117, n_32118);
  and g72131 (n43094, pi1156, n42828);
  not g72132 (n_32119, n43093);
  not g72133 (n_32120, n43094);
  and g72134 (n43095, n_32119, n_32120);
  not g72135 (n_32121, n43085);
  not g72136 (n_32122, n43095);
  and g72137 (n43096, n_32121, n_32122);
  not g72138 (n_32123, n43096);
  and g72139 (n43097, pi0211, n_32123);
  and g72140 (n43098, n_30549, n41091);
  and g72141 (n43099, pi1155, n43098);
  not g72142 (n_32124, n43099);
  and g72143 (n43100, n43086, n_32124);
  and g72144 (n43101, n_31892, n43100);
  not g72145 (n_32125, n43101);
  and g72146 (n43102, pi1156, n_32125);
  and g72147 (n43103, n_32115, n43102);
  not g72148 (n_32126, n43100);
  and g72149 (n43104, n43091, n_32126);
  not g72150 (n_32127, n43103);
  and g72151 (n43105, n_7075, n_32127);
  not g72152 (n_32128, n43104);
  and g72153 (n43106, n_32128, n43105);
  not g72154 (n_32129, n43106);
  and g72155 (n43107, n_6791, n_32129);
  not g72156 (n_32130, n43097);
  and g72157 (n43108, n_32130, n43107);
  not g72158 (n_32131, n43083);
  and g72159 (n43109, pi0263, n_32131);
  not g72160 (n_32132, n43108);
  and g72161 (n43110, n_32132, n43109);
  not g72162 (n_32133, n43067);
  and g72163 (n43111, n40860, n_32133);
  not g72164 (n_32134, n43110);
  and g72165 (n43112, n_32134, n43111);
  not g72166 (n_32135, n43017);
  and g72167 (n43113, n_4226, n_32135);
  not g72168 (n_32136, n43112);
  and g72169 (n43114, n_32136, n43113);
  not g72170 (n_32137, n43016);
  and g72171 (n43115, n40910, n_32137);
  not g72172 (n_32138, n43114);
  and g72173 (n43116, n_32138, n43115);
  not g72174 (n_32139, n42996);
  and g72175 (n43117, n_28510, n_32139);
  not g72176 (n_32140, n43116);
  and g72177 (n43118, n_32140, n43117);
  and g72178 (n43119, po1038, n42990);
  and g72179 (n43120, n_28679, n38649);
  not g72180 (n_32141, n43120);
  and g72181 (n43121, n_11794, n_32141);
  not g72182 (n_32142, n39112);
  and g72183 (n43122, n38592, n_32142);
  not g72184 (n_32143, n43121);
  and g72185 (n43123, n_32143, n43122);
  and g72186 (n43124, pi1156, n39854);
  not g72187 (n_32144, n43124);
  and g72188 (n43125, pi0219, n_32144);
  not g72189 (n_32145, n43123);
  and g72190 (n43126, n_32145, n43125);
  and g72191 (n43127, n_28743, n_32145);
  not g72192 (n_32146, n43127);
  and g72193 (n43128, pi0211, n_32146);
  not g72194 (n_32147, n43128);
  and g72195 (n43129, n42980, n_32147);
  not g72196 (n_32148, n43126);
  and g72197 (n43130, n_4226, n_32148);
  not g72198 (n_32149, n43129);
  and g72199 (n43131, n_32149, n43130);
  not g72200 (n_32150, n43119);
  and g72201 (n43132, pi0230, n_32150);
  not g72202 (n_32151, n43131);
  and g72203 (n43133, n_32151, n43132);
  not g72204 (n_32152, n43118);
  not g72205 (n_32153, n43133);
  and g72206 (po0420, n_32152, n_32153);
  and g72207 (n43135, pi1091, pi1143);
  and g72208 (n43136, n_7045, n43135);
  not g72209 (n_32155, pi0796);
  and g72210 (n43137, n_32155, n40863);
  not g72211 (n_32156, n40863);
  and g72212 (n43138, pi0264, n_32156);
  not g72213 (n_32157, n43137);
  and g72214 (n43139, n_3128, n_32157);
  not g72215 (n_32158, n43138);
  and g72216 (n43140, n_32158, n43139);
  not g72217 (n_32159, n43136);
  and g72218 (n43141, pi0199, n_32159);
  not g72219 (n_32160, n43140);
  and g72220 (n43142, n_32160, n43141);
  and g72221 (n43143, pi1091, pi1141);
  and g72222 (n43144, n_32155, n40885);
  not g72223 (n_32161, n40885);
  and g72224 (n43145, pi0264, n_32161);
  not g72225 (n_32162, n43144);
  and g72226 (n43146, n_3128, n_32162);
  not g72227 (n_32163, n43145);
  and g72228 (n43147, n_32163, n43146);
  not g72229 (n_32164, n43143);
  not g72230 (n_32165, n43147);
  and g72231 (n43148, n_32164, n_32165);
  not g72232 (n_32166, n43148);
  and g72233 (n43149, n_7045, n_32166);
  and g72234 (n43150, pi1091, pi1142);
  not g72235 (n_32167, n43150);
  and g72236 (n43151, n_32165, n_32167);
  not g72237 (n_32168, n43151);
  and g72238 (n43152, pi0200, n_32168);
  not g72239 (n_32169, n43149);
  and g72240 (n43153, n_7044, n_32169);
  not g72241 (n_32170, n43152);
  and g72242 (n43154, n_32170, n43153);
  not g72243 (n_32171, n43142);
  and g72244 (n43155, n16479, n_32171);
  not g72245 (n_32172, n43154);
  and g72246 (n43156, n_32172, n43155);
  not g72247 (n_32173, n42455);
  and g72248 (n43157, pi0219, n_32173);
  not g72249 (n_32174, n43157);
  and g72250 (n43158, n_29299, n_32174);
  not g72251 (n_32175, n43158);
  and g72252 (n43159, n_32160, n_32175);
  and g72253 (n43160, n_7075, n_32166);
  and g72254 (n43161, pi0211, n_32168);
  not g72255 (n_32176, n43160);
  and g72256 (n43162, n_6791, n_32176);
  not g72257 (n_32177, n43161);
  and g72258 (n43163, n_32177, n43162);
  not g72259 (n_32178, n43159);
  and g72260 (n43164, n_25711, n_32178);
  not g72261 (n_32179, n43163);
  and g72262 (n43165, n_32179, n43164);
  not g72263 (n_32180, n43156);
  not g72264 (n_32181, n43165);
  and g72265 (n43166, n_32180, n_32181);
  not g72266 (n_32182, n43166);
  and g72267 (n43167, n_28510, n_32182);
  and g72268 (n43168, n_7075, pi1141);
  and g72269 (n43169, n_6791, n_28545);
  not g72270 (n_32183, n43168);
  and g72271 (n43170, n_32183, n43169);
  not g72272 (n_32184, n43170);
  and g72273 (n43171, n_29299, n_32184);
  not g72274 (n_32185, n43171);
  and g72275 (n43172, n_25711, n_32185);
  and g72276 (n43173, n_7044, pi1141);
  not g72277 (n_32186, n43173);
  and g72278 (n43174, n39388, n_32186);
  not g72279 (n_32187, n43174);
  and g72280 (n43175, n_28534, n_32187);
  not g72281 (n_32188, n43175);
  and g72282 (n43176, n16479, n_32188);
  not g72283 (n_32189, n43172);
  and g72284 (n43177, pi0230, n_32189);
  not g72285 (n_32190, n43176);
  and g72286 (n43178, n_32190, n43177);
  or g72287 (po0421, n43167, n43178);
  and g72288 (n43180, pi1091, pi1144);
  and g72289 (n43181, n_7045, n43180);
  not g72290 (n_32192, pi0819);
  and g72291 (n43182, n_32192, n40863);
  and g72292 (n43183, pi0265, n_32156);
  not g72293 (n_32193, n43182);
  and g72294 (n43184, n_3128, n_32193);
  not g72295 (n_32194, n43183);
  and g72296 (n43185, n_32194, n43184);
  not g72297 (n_32195, n43181);
  and g72298 (n43186, pi0199, n_32195);
  not g72299 (n_32196, n43185);
  and g72300 (n43187, n_32196, n43186);
  and g72301 (n43188, n_32192, n40885);
  and g72302 (n43189, pi0265, n_32161);
  not g72303 (n_32197, n43188);
  and g72304 (n43190, n_3128, n_32197);
  not g72305 (n_32198, n43189);
  and g72306 (n43191, n_32198, n43190);
  not g72307 (n_32199, n43191);
  and g72308 (n43192, n_32167, n_32199);
  not g72309 (n_32200, n43192);
  and g72310 (n43193, n_7045, n_32200);
  not g72311 (n_32201, n43135);
  and g72312 (n43194, n_32201, n_32199);
  not g72313 (n_32202, n43194);
  and g72314 (n43195, pi0200, n_32202);
  not g72315 (n_32203, n43193);
  and g72316 (n43196, n_7044, n_32203);
  not g72317 (n_32204, n43195);
  and g72318 (n43197, n_32204, n43196);
  not g72319 (n_32205, n43187);
  and g72320 (n43198, n16479, n_32205);
  not g72321 (n_32206, n43197);
  and g72322 (n43199, n_32206, n43198);
  and g72323 (n43200, n_30353, n_32174);
  not g72324 (n_32207, n43200);
  and g72325 (n43201, n_32196, n_32207);
  and g72326 (n43202, n_7075, n_32200);
  and g72327 (n43203, pi0211, n_32202);
  not g72328 (n_32208, n43202);
  and g72329 (n43204, n_6791, n_32208);
  not g72330 (n_32209, n43203);
  and g72331 (n43205, n_32209, n43204);
  not g72332 (n_32210, n43201);
  and g72333 (n43206, n_25711, n_32210);
  not g72334 (n_32211, n43205);
  and g72335 (n43207, n_32211, n43206);
  not g72336 (n_32212, n43199);
  not g72337 (n_32213, n43207);
  and g72338 (n43208, n_32212, n_32213);
  not g72339 (n_32214, n43208);
  and g72340 (n43209, n_28510, n_32214);
  and g72341 (n43210, n_7075, pi1142);
  and g72342 (n43211, n_6791, n_28514);
  not g72343 (n_32215, n43210);
  and g72344 (n43212, n_32215, n43211);
  not g72345 (n_32216, n43212);
  and g72346 (n43213, n_30353, n_32216);
  not g72347 (n_32217, n43213);
  and g72348 (n43214, n_25711, n_32217);
  and g72349 (n43215, n_28533, n40782);
  not g72350 (n_32218, n43215);
  and g72351 (n43216, n_28530, n_32218);
  not g72352 (n_32219, n43216);
  and g72353 (n43217, n16479, n_32219);
  not g72354 (n_32220, n43214);
  and g72355 (n43218, pi0230, n_32220);
  not g72356 (n_32221, n43217);
  and g72357 (n43219, n_32221, n43218);
  or g72358 (po0422, n43209, n43219);
  and g72359 (n43221, n_7075, pi1136);
  not g72360 (n_32222, n43221);
  and g72361 (n43222, pi0219, n_32222);
  and g72362 (n43223, pi0211, n_2581);
  not g72363 (n_32223, n43222);
  not g72364 (n_32224, n43223);
  and g72365 (n43224, n_32223, n_32224);
  and g72366 (n43225, n_7076, n43224);
  and g72367 (n43226, po1038, n43225);
  and g72368 (n43227, pi0299, n43225);
  and g72369 (n43228, n_7044, pi1135);
  not g72370 (n_32225, n43228);
  and g72371 (n43229, pi0200, n_32225);
  and g72372 (n43230, pi0199, pi1136);
  not g72373 (n_32226, n43230);
  and g72374 (n43231, n_7045, n_32226);
  not g72375 (n_32227, n43229);
  and g72376 (n43232, n_234, n_32227);
  not g72377 (n_32228, n43231);
  and g72378 (n43233, n_32228, n43232);
  not g72379 (n_32229, n43227);
  not g72380 (n_32230, n43233);
  and g72381 (n43234, n_32229, n_32230);
  not g72382 (n_32231, n43234);
  and g72383 (n43235, n_4226, n_32231);
  not g72384 (n_32232, n43226);
  and g72385 (n43236, pi0230, n_32232);
  not g72386 (n_32233, n43235);
  and g72387 (n43237, n_32233, n43236);
  and g72388 (n43238, n_32174, n_32223);
  and g72389 (n43239, n_2416, n_32156);
  not g72390 (n_32235, pi0948);
  and g72391 (n43240, n_32235, n40863);
  not g72392 (n_32236, n43239);
  and g72393 (n43241, n_3128, n_32236);
  not g72394 (n_32237, n43240);
  and g72395 (n43242, n_32237, n43241);
  not g72396 (n_32238, n43238);
  not g72397 (n_32239, n43242);
  and g72398 (n43243, n_32238, n_32239);
  not g72399 (n_32240, n43243);
  and g72400 (n43244, n_25711, n_32240);
  and g72401 (n43245, n_2416, n_32161);
  and g72402 (n43246, n_32235, n40885);
  not g72403 (n_32241, n43245);
  and g72404 (n43247, n_3128, n_32241);
  not g72405 (n_32242, n43246);
  and g72406 (n43248, n_32242, n43247);
  not g72407 (n_32243, n43248);
  and g72408 (n43249, n_6791, n_32243);
  and g72409 (n43250, pi1135, n42424);
  not g72410 (n_32244, n43250);
  and g72411 (n43251, n43249, n_32244);
  not g72412 (n_32245, n43251);
  and g72413 (n43252, n43244, n_32245);
  and g72414 (n43253, n_7044, n_32243);
  and g72415 (n43254, pi1091, pi1136);
  and g72416 (n43255, pi0199, n_32239);
  not g72417 (n_32246, n43254);
  and g72418 (n43256, n_32246, n43255);
  not g72419 (n_32247, n43253);
  not g72420 (n_32248, n43256);
  and g72421 (n43257, n_32247, n_32248);
  and g72422 (n43258, n_7045, n43257);
  and g72423 (n43259, pi1091, pi1135);
  not g72424 (n_32249, n43259);
  and g72425 (n43260, n43253, n_32249);
  not g72426 (n_32250, n43255);
  and g72427 (n43261, pi0200, n_32250);
  not g72428 (n_32251, n43260);
  and g72429 (n43262, n_32251, n43261);
  not g72430 (n_32252, n43258);
  not g72431 (n_32253, n43262);
  and g72432 (n43263, n_32252, n_32253);
  not g72433 (n_32254, n43263);
  and g72434 (n43264, n16479, n_32254);
  not g72435 (n_32255, n43252);
  and g72436 (n43265, n_28510, n_32255);
  not g72437 (n_32256, n43264);
  and g72438 (n43266, n_32256, n43265);
  not g72439 (n_32257, n43237);
  not g72440 (n_32258, n43266);
  and g72441 (n43267, n_32257, n_32258);
  not g72442 (n_32259, n43267);
  and g72443 (n43268, n_2921, n_32259);
  and g72444 (n43269, n38699, n_32226);
  not g72445 (n_32260, n43269);
  and g72446 (n43270, n_32227, n_32260);
  and g72447 (n43271, n16479, n43270);
  and g72448 (n43272, n_25711, n43224);
  not g72449 (n_32261, n43271);
  and g72450 (n43273, pi0230, n_32261);
  not g72451 (n_32262, n43272);
  and g72452 (n43274, n_32262, n43273);
  and g72453 (n43275, pi1091, n_32224);
  not g72454 (n_32263, n43275);
  and g72455 (n43276, n43249, n_32263);
  not g72456 (n_32264, n43276);
  and g72457 (n43277, n43244, n_32264);
  and g72458 (n43278, n_7044, pi1091);
  not g72459 (n_32265, n43257);
  not g72460 (n_32266, n43278);
  and g72461 (n43279, n_32265, n_32266);
  not g72462 (n_32267, n43279);
  and g72463 (n43280, n_7045, n_32267);
  not g72464 (n_32268, n43280);
  and g72465 (n43281, n_32253, n_32268);
  not g72466 (n_32269, n43281);
  and g72467 (n43282, n16479, n_32269);
  not g72468 (n_32270, n43277);
  and g72469 (n43283, n_28510, n_32270);
  not g72470 (n_32271, n43282);
  and g72471 (n43284, n_32271, n43283);
  not g72472 (n_32272, n43274);
  not g72473 (n_32273, n43284);
  and g72474 (n43285, n_32272, n_32273);
  not g72475 (n_32274, n43285);
  and g72476 (n43286, pi1134, n_32274);
  not g72477 (n_32275, n43268);
  not g72478 (n_32276, n43286);
  and g72479 (po0423, n_32275, n_32276);
  and g72480 (n43288, pi1155, n_31594);
  and g72481 (n43289, n_31802, n43288);
  and g72482 (n43290, n_11768, n_31440);
  and g72483 (n43291, pi1091, n43290);
  not g72484 (n_32277, n43289);
  not g72485 (n_32278, n43291);
  and g72486 (n43292, n_32277, n_32278);
  not g72487 (n_32279, n43292);
  and g72488 (n43293, n_11413, n_32279);
  and g72489 (n43294, n42716, n43288);
  and g72490 (n43295, n_11768, n_31769);
  and g72491 (n43296, n_31616, n43295);
  not g72492 (n_32280, n43294);
  not g72493 (n_32281, n43296);
  and g72494 (n43297, n_32280, n_32281);
  not g72495 (n_32282, n43297);
  and g72496 (n43298, pi1154, n_32282);
  not g72497 (n_32283, n43293);
  and g72498 (n43299, n_6791, n_32283);
  not g72499 (n_32284, n43298);
  and g72500 (n43300, n_32284, n43299);
  and g72501 (n43301, pi1153, n38955);
  not g72502 (n_32285, n43301);
  and g72503 (n43302, n42708, n_32285);
  and g72504 (n43303, n_29492, n43302);
  and g72505 (n43304, pi1091, n42928);
  and g72506 (n43305, n_31595, n43304);
  not g72507 (n_32286, n43305);
  and g72508 (n43306, pi1154, n_32286);
  and g72509 (n43307, n_234, n38946);
  not g72510 (n_32287, n43307);
  and g72511 (n43308, pi1091, n_32287);
  and g72512 (n43309, n43306, n43308);
  not g72513 (n_32288, n43303);
  and g72514 (n43310, pi0219, n_32288);
  not g72515 (n_32289, n43309);
  and g72516 (n43311, n_32289, n43310);
  not g72517 (n_32290, n43300);
  not g72518 (n_32291, n43311);
  and g72519 (n43312, n_32290, n_32291);
  not g72520 (n_32292, n43312);
  and g72521 (n43313, n_7075, n_32292);
  and g72522 (n43314, pi1155, n38963);
  not g72523 (n_32293, n43314);
  and g72524 (n43315, pi1154, n_32293);
  and g72525 (n43316, n_11768, n_29535);
  not g72526 (n_32294, n43316);
  and g72527 (n43317, n_28725, n_32294);
  not g72528 (n_32295, n43317);
  and g72529 (n43318, n_8689, n_32295);
  and g72530 (n43319, pi1091, n43315);
  not g72531 (n_32296, n43318);
  and g72532 (n43320, n_32296, n43319);
  and g72533 (n43321, n_28726, n_30462);
  not g72534 (n_32297, n43321);
  and g72535 (n43322, n43302, n_32297);
  not g72536 (n_32298, n43322);
  and g72537 (n43323, pi0211, n_32298);
  not g72538 (n_32299, n43320);
  and g72539 (n43324, n_32299, n43323);
  not g72540 (n_32300, n43313);
  not g72541 (n_32301, n43324);
  and g72542 (n43325, n_32300, n_32301);
  not g72543 (n_32302, n43325);
  and g72544 (n43326, pi0267, n_32302);
  and g72545 (n43327, n38568, n42448);
  not g72546 (n_32303, n43327);
  and g72547 (n43328, n_31786, n_32303);
  not g72548 (n_32304, n43290);
  not g72549 (n_32305, n43328);
  and g72550 (n43329, n_32304, n_32305);
  and g72551 (n43330, pi0211, n_11413);
  not g72552 (n_32306, n43329);
  and g72553 (n43331, n_32306, n43330);
  and g72554 (n43332, pi1091, n_11768);
  and g72555 (n43333, n_29535, n43332);
  not g72556 (n_32307, n43333);
  and g72557 (n43334, n38488, n_32307);
  and g72558 (n43335, n_32286, n43334);
  and g72559 (n43336, n_11413, n38545);
  not g72560 (n_32308, n43336);
  and g72561 (n43337, n_28701, n_32308);
  and g72562 (n43338, n_28710, n43337);
  and g72563 (n43339, pi1091, n43338);
  not g72564 (n_32309, n43339);
  and g72565 (n43340, n_7075, n_32309);
  not g72566 (n_32310, n43335);
  and g72567 (n43341, n_6791, n_32310);
  not g72568 (n_32311, n43340);
  and g72569 (n43342, n_32311, n43341);
  and g72570 (n43343, n43307, n43332);
  not g72571 (n_32312, n43343);
  and g72572 (n43344, n43306, n_32312);
  and g72573 (n43345, n42928, n43315);
  not g72574 (n_32313, n43344);
  not g72575 (n_32314, n43345);
  and g72576 (n43346, n_32313, n_32314);
  not g72577 (n_32315, n43346);
  and g72578 (n43347, pi0211, n_32315);
  and g72579 (n43348, pi1154, n_32313);
  and g72580 (n43349, n_28726, n42708);
  and g72581 (n43350, n_29490, n43349);
  not g72582 (n_32316, n43350);
  and g72583 (n43351, n_7075, n_32316);
  not g72584 (n_32317, n43348);
  and g72585 (n43352, n_32317, n43351);
  not g72586 (n_32318, n43347);
  and g72587 (n43353, pi0219, n_32318);
  not g72588 (n_32319, n43352);
  and g72589 (n43354, n_32319, n43353);
  not g72590 (n_32320, n43342);
  not g72591 (n_32321, n43354);
  and g72592 (n43355, n_32320, n_32321);
  not g72593 (n_32322, pi0267);
  not g72594 (n_32323, n43331);
  and g72595 (n43356, n_32322, n_32323);
  not g72596 (n_32324, n43355);
  and g72597 (n43357, n_32324, n43356);
  not g72598 (n_32325, n43326);
  not g72599 (n_32326, n43357);
  and g72600 (n43358, n_32325, n_32326);
  and g72601 (n43359, n_4226, n43358);
  and g72602 (n43360, n_6791, n_28570);
  and g72603 (n43361, n_28578, n43360);
  not g72604 (n_32327, n43361);
  and g72605 (n43362, n_29089, n_32327);
  not g72606 (n_32328, n43362);
  and g72607 (n43363, pi1091, n_32328);
  and g72608 (n43364, n_32322, n_3128);
  not g72609 (n_32329, n43363);
  not g72610 (n_32330, n43364);
  and g72611 (n43365, n_32329, n_32330);
  not g72612 (n_32331, n43365);
  and g72613 (n43366, po1038, n_32331);
  not g72614 (n_32332, n43366);
  and g72615 (n43367, n_30644, n_32332);
  not g72616 (n_32333, n43359);
  and g72617 (n43368, n_32333, n43367);
  and g72618 (n43369, n_32322, n_30509);
  and g72619 (n43370, n_31670, n43369);
  and g72620 (n43371, pi0267, n42734);
  not g72621 (n_32334, n43370);
  and g72622 (n43372, n40859, n_32334);
  not g72623 (n_32335, n43371);
  and g72624 (n43373, n_32335, n43372);
  not g72625 (n_32336, n40859);
  and g72626 (n43374, n_32336, n43364);
  not g72627 (n_32337, n43374);
  and g72628 (n43375, n_32329, n_32337);
  not g72629 (n_32338, n43373);
  and g72630 (n43376, n_32338, n43375);
  not g72631 (n_32339, n43376);
  and g72632 (n43377, po1038, n_32339);
  not g72633 (n_32340, n43358);
  and g72634 (n43378, n_32336, n_32340);
  and g72635 (n43379, n_31851, n42780);
  not g72636 (n_32341, n43379);
  and g72637 (n43380, n42805, n_32341);
  not g72641 (n_32342, n43380);
  not g72642 (n_32343, n43383);
  and g72643 (n43384, n_32342, n_32343);
  not g72644 (n_32344, n43384);
  and g72645 (n43385, pi0211, n_32344);
  and g72646 (n43386, pi1153, n41055);
  not g72648 (n_32345, n43386);
  and g72651 (n43390, n41039, n42749);
  not g72652 (n_32346, n43390);
  and g72653 (n43391, n_11768, n_32346);
  and g72654 (n43392, n_32341, n43391);
  and g72661 (n43396, pi1155, n_31706);
  and g72662 (n43397, n41008, n_32092);
  not g72663 (n_32350, n43397);
  and g72664 (n43398, n43396, n_32350);
  not g72665 (n_32351, n42598);
  and g72666 (n43399, n_32351, n43398);
  not g72667 (n_32352, n42501);
  and g72668 (n43400, n_32352, n_31656);
  not g72669 (n_32353, n43400);
  and g72670 (n43401, n41009, n_32353);
  not g72671 (n_32354, n43401);
  and g72672 (n43402, pi1154, n_32354);
  and g72673 (n43403, n_11413, n_30550);
  and g72674 (n43404, n_31717, n43403);
  not g72675 (n_32355, n43404);
  and g72676 (n43405, n_11768, n_32355);
  not g72677 (n_32356, n43402);
  and g72678 (n43406, n_32356, n43405);
  not g72679 (n_32357, n43399);
  and g72680 (n43407, pi0267, n_32357);
  not g72681 (n_32358, n43406);
  and g72682 (n43408, n_32358, n43407);
  not g72683 (n_32359, n43395);
  not g72684 (n_32360, n43408);
  and g72685 (n43409, n_32359, n_32360);
  not g72686 (n_32361, n43409);
  and g72687 (n43410, pi0219, n_32361);
  not g72688 (n_32362, n42825);
  and g72689 (n43411, n_11768, n_32362);
  and g72690 (n43412, n_32341, n43411);
  and g72691 (n43413, n41072, n_32354);
  not g72692 (n_32363, n43413);
  and g72693 (n43414, n43070, n_32363);
  not g72694 (n_32364, n43414);
  and g72695 (n43415, pi1154, n_32364);
  and g72696 (n43416, n_11413, n_31643);
  not g72697 (n_32365, n43416);
  and g72698 (n43417, pi1155, n_32365);
  not g72699 (n_32366, n43417);
  and g72700 (n43418, n41045, n_32366);
  not g72701 (n_32367, n43415);
  not g72702 (n_32368, n43418);
  and g72703 (n43419, n_32367, n_32368);
  not g72704 (n_32369, n43412);
  and g72705 (n43420, pi0211, n_32369);
  not g72706 (n_32370, n43419);
  and g72707 (n43421, n_32370, n43420);
  and g72708 (n43422, n_31892, n_32345);
  not g72709 (n_32371, n43422);
  and g72710 (n43423, pi1155, n_32371);
  and g72711 (n43424, pi1153, n_30612);
  not g72712 (n_32372, n43424);
  and g72713 (n43425, n_11768, n_32372);
  and g72714 (n43426, n42605, n43425);
  not g72715 (n_32373, n43423);
  and g72716 (n43427, n_11413, n_32373);
  not g72717 (n_32374, n43426);
  and g72718 (n43428, n_32374, n43427);
  not g72719 (n_32375, n43098);
  and g72720 (n43429, n_11757, n_32375);
  not g72721 (n_32376, n43429);
  and g72722 (n43430, n43425, n_32376);
  not g72727 (n_32378, n43428);
  and g72728 (n43434, n_7075, n_32378);
  not g72729 (n_32379, n43433);
  and g72730 (n43435, n_32379, n43434);
  not g72731 (n_32380, n43435);
  and g72732 (n43436, n_32322, n_32380);
  not g72733 (n_32381, n43421);
  and g72734 (n43437, n_32381, n43436);
  and g72735 (n43438, n_11757, n41093);
  not g72736 (n_32382, n43438);
  and g72737 (n43439, n_31642, n_32382);
  and g72738 (n43440, n_11768, n41072);
  not g72739 (n_32383, n43439);
  and g72740 (n43441, n_32383, n43440);
  and g72741 (n43442, n43033, n43396);
  not g72742 (n_32384, n43441);
  and g72743 (n43443, pi1154, n_32384);
  not g72744 (n_32385, n43442);
  and g72745 (n43444, n_32385, n43443);
  and g72746 (n43445, n_11413, n_31656);
  not g72747 (n_32386, n41105);
  and g72748 (n43446, n_32386, n43445);
  not g72749 (n_32387, n43446);
  and g72750 (n43447, n_11768, n_32387);
  and g72751 (n43448, n_30518, n43445);
  not g72752 (n_32388, n43447);
  and g72753 (n43449, n_32388, n43448);
  not g72754 (n_32389, n43444);
  not g72755 (n_32390, n43449);
  and g72756 (n43450, n_32389, n_32390);
  not g72757 (n_32391, n43450);
  and g72758 (n43451, pi0211, n_32391);
  and g72759 (n43452, pi1154, n43439);
  not g72760 (n_32392, n43452);
  and g72761 (n43453, n43447, n_32392);
  and g72762 (n43454, pi1154, n41008);
  and g72763 (n43455, n_30611, n_31876);
  not g72764 (n_32393, n43454);
  and g72765 (n43456, pi1155, n_32393);
  not g72766 (n_32394, n43455);
  and g72767 (n43457, n_32394, n43456);
  not g72768 (n_32395, n43457);
  and g72769 (n43458, n_7075, n_32395);
  not g72770 (n_32396, n43453);
  and g72771 (n43459, n_32396, n43458);
  not g72772 (n_32397, n43459);
  and g72773 (n43460, pi0267, n_32397);
  not g72774 (n_32398, n43451);
  and g72775 (n43461, n_32398, n43460);
  not g72776 (n_32399, n43461);
  and g72777 (n43462, n_6791, n_32399);
  not g72778 (n_32400, n43437);
  and g72779 (n43463, n_32400, n43462);
  not g72780 (n_32401, n43410);
  not g72781 (n_32402, n43463);
  and g72782 (n43464, n_32401, n_32402);
  not g72783 (n_32403, n43464);
  and g72784 (n43465, n40859, n_32403);
  not g72785 (n_32404, n43378);
  and g72786 (n43466, n_4226, n_32404);
  not g72787 (n_32405, n43465);
  and g72788 (n43467, n_32405, n43466);
  not g72789 (n_32406, n43377);
  and g72790 (n43468, n40910, n_32406);
  not g72791 (n_32407, n43467);
  and g72792 (n43469, n_32407, n43468);
  not g72793 (n_32408, n43368);
  and g72794 (n43470, n_28510, n_32408);
  not g72795 (n_32409, n43469);
  and g72796 (n43471, n_32409, n43470);
  and g72797 (n43472, pi0219, n_28934);
  and g72798 (n43473, n_11768, n43301);
  not g72799 (n_32410, n43473);
  and g72800 (n43474, n_11413, n_32410);
  not g72801 (n_32411, n43474);
  and g72802 (n43475, n_29535, n_32411);
  and g72803 (n43476, pi1155, n39665);
  not g72804 (n_32412, n43475);
  not g72805 (n_32413, n43476);
  and g72806 (n43477, n_32412, n_32413);
  not g72807 (n_32414, n43472);
  not g72808 (n_32415, n43477);
  and g72809 (n43478, n_32414, n_32415);
  not g72810 (n_32416, n43478);
  and g72811 (n43479, pi0211, n_32416);
  and g72812 (n43480, n_7044, pi1154);
  not g72813 (n_32417, n43480);
  and g72814 (n43481, pi0200, n_32417);
  and g72815 (n43482, n_28749, n_28933);
  not g72816 (n_32418, n43481);
  and g72817 (n43483, n_32418, n43482);
  not g72818 (n_32419, n43483);
  and g72819 (n43484, n_28743, n_32419);
  not g72820 (n_32420, n43484);
  and g72821 (n43485, pi0219, n_32420);
  and g72822 (n43486, n_6791, n43338);
  not g72823 (n_32421, n43486);
  and g72824 (n43487, n_7075, n_32421);
  not g72825 (n_32422, n43485);
  and g72826 (n43488, n_32422, n43487);
  not g72827 (n_32423, n43488);
  and g72828 (n43489, n_4226, n_32423);
  not g72829 (n_32424, n43479);
  and g72830 (n43490, n_32424, n43489);
  and g72831 (n43491, po1038, n43362);
  not g72832 (n_32425, n43491);
  and g72833 (n43492, pi0230, n_32425);
  not g72834 (n_32426, n43490);
  and g72835 (n43493, n_32426, n43492);
  not g72836 (n_32427, n43471);
  not g72837 (n_32428, n43493);
  and g72838 (po0424, n_32427, n_32428);
  and g72839 (n43495, pi0268, pi1152);
  and g72840 (n43496, n_7075, n_25711);
  and g72841 (n43497, n_4226, n38568);
  not g72842 (n_32429, n43496);
  not g72843 (n_32430, n43497);
  and g72844 (n43498, n_32429, n_32430);
  and g72845 (n43499, n_29468, n43498);
  and g72846 (n43500, n_7044, n16479);
  not g72847 (n_32431, n40141);
  not g72848 (n_32432, n43500);
  and g72849 (n43501, n_32431, n_32432);
  not g72850 (n_32433, n43498);
  and g72851 (n43502, pi1152, n_32433);
  not g72852 (n_32434, n43502);
  and g72853 (n43503, n43501, n_32434);
  not g72854 (n_32435, n43499);
  and g72855 (n43504, pi1150, n_32435);
  not g72856 (n_32436, n43503);
  and g72857 (n43505, n_32436, n43504);
  not g72858 (n_32437, n43495);
  and g72859 (n43506, n_32437, n43505);
  and g72860 (n43507, n_29468, n42389);
  and g72861 (n43508, n_4226, n_7411);
  and g72862 (n43509, po1038, n11446);
  not g72863 (n_32438, n43508);
  not g72864 (n_32439, n43509);
  and g72865 (n43510, n_32438, n_32439);
  not g72866 (n_32440, n43510);
  and g72867 (n43511, pi1151, n_32440);
  not g72868 (n_32441, n43511);
  and g72869 (n43512, n_28873, n_32441);
  and g72870 (n43513, n_25711, n42478);
  and g72871 (n43514, n_4226, n38581);
  not g72872 (n_32442, n43513);
  not g72873 (n_32443, n43514);
  and g72874 (n43515, n_32442, n_32443);
  not g72875 (n_32444, n43515);
  and g72876 (n43516, pi1151, n_32444);
  and g72877 (n43517, pi1152, n43516);
  not g72884 (n_32448, n43506);
  not g72885 (n_32449, n43520);
  and g72886 (n43521, n_32448, n_32449);
  not g72887 (n_32450, n43521);
  and g72888 (n43522, pi1091, n_32450);
  and g72889 (n43523, pi1152, n43505);
  not g72890 (n_32451, n43523);
  and g72891 (n43524, pi1091, n_32451);
  not g72892 (n_32452, n43524);
  and g72893 (n43525, pi0268, n_32452);
  not g72894 (n_32453, n43522);
  not g72895 (n_32454, n43525);
  and g72896 (n43526, n_32453, n_32454);
  not g72897 (n_32455, n40909);
  not g72898 (n_32456, n43526);
  and g72899 (n43527, n_32455, n_32456);
  and g72900 (n43528, n_31664, n42572);
  and g72901 (n43529, n_30536, n42584);
  and g72902 (n43530, pi0219, n_31653);
  and g72903 (n43531, n_30537, n43530);
  not g72904 (n_32457, n43529);
  not g72905 (n_32458, n43531);
  and g72906 (n43532, n_32457, n_32458);
  and g72907 (n43533, n_4226, n_31646);
  and g72908 (n43534, n43532, n43533);
  not g72909 (n_32459, n43528);
  not g72910 (n_32460, n43534);
  and g72911 (n43535, n_32459, n_32460);
  not g72912 (n_32461, n43535);
  and g72913 (n43536, n_29468, n_32461);
  not g72914 (n_32462, n42606);
  and g72915 (n43537, n_4226, n_32462);
  and g72916 (n43538, pi0219, n41048);
  not g72917 (n_32463, n43538);
  and g72918 (n43539, n43537, n_32463);
  and g72919 (n43540, n42572, n_31823);
  not g72920 (n_32464, n43539);
  not g72921 (n_32465, n43540);
  and g72922 (n43541, n_32464, n_32465);
  not g72923 (n_32466, n43541);
  and g72924 (n43542, pi1151, n_32466);
  not g72925 (n_32467, n43536);
  not g72926 (n_32468, n43542);
  and g72927 (n43543, n_32467, n_32468);
  not g72928 (n_32469, n43543);
  and g72929 (n43544, pi0268, n_32469);
  and g72930 (n43545, po1038, n_31670);
  and g72931 (n43546, n_31695, n43545);
  and g72932 (n43547, po1038, n_31822);
  and g72933 (n43548, n_31665, n43547);
  not g72934 (n_32470, n43548);
  and g72935 (n43549, n43546, n_32470);
  and g72936 (n43550, pi0219, n_30523);
  not g72937 (n_32471, n42548);
  not g72938 (n_32472, n43550);
  and g72939 (n43551, n_32471, n_32472);
  not g72940 (n_32473, n43551);
  and g72941 (n43552, n_30522, n_32473);
  and g72942 (n43553, n_4226, n_30549);
  and g72943 (n43554, n43552, n43553);
  not g72944 (n_32474, n43549);
  not g72945 (n_32475, n43554);
  and g72946 (n43555, n_32474, n_32475);
  and g72947 (n43556, n_29468, n43555);
  and g72948 (n43557, n_30508, n_32466);
  and g72949 (n43558, pi0219, po1038);
  and g72950 (n43559, n_30521, n43558);
  and g72951 (n43560, n_30554, n43537);
  not g72952 (n_32476, n43559);
  and g72953 (n43561, n_31669, n_32476);
  not g72954 (n_32477, n43560);
  and g72955 (n43562, n_32477, n43561);
  not g72956 (n_32478, n43557);
  not g72957 (n_32479, n43562);
  and g72958 (n43563, n_32478, n_32479);
  and g72959 (n43564, pi1151, n43563);
  not g72960 (n_32480, pi0268);
  not g72961 (n_32481, n43564);
  and g72962 (n43565, n_32480, n_32481);
  not g72963 (n_32482, n43556);
  and g72964 (n43566, n_32482, n43565);
  not g72965 (n_32483, n43544);
  not g72966 (n_32484, n43566);
  and g72967 (n43567, n_32483, n_32484);
  not g72968 (n_32485, n43567);
  and g72969 (n43568, n_28873, n_32485);
  and g72970 (n43569, n_31664, n43547);
  and g72971 (n43570, n_31707, n_31718);
  not g72972 (n_32486, n43532);
  not g72973 (n_32487, n43570);
  and g72974 (n43571, n_32486, n_32487);
  not g72975 (n_32488, n43571);
  and g72976 (n43572, n_4226, n_32488);
  and g72977 (n43573, n_30521, n_31846);
  not g72978 (n_32489, n43573);
  and g72979 (n43574, n43572, n_32489);
  not g72980 (n_32490, n43569);
  not g72981 (n_32491, n43574);
  and g72982 (n43575, n_32490, n_32491);
  not g72983 (n_32492, n43575);
  and g72984 (n43576, n_29468, n_32492);
  and g72985 (n43577, n_30424, n43533);
  and g72986 (n43578, n_31823, n43547);
  not g72987 (n_32493, n43578);
  and g72988 (n43579, n_32464, n_32493);
  not g72989 (n_32494, n43577);
  and g72990 (n43580, n_32494, n43579);
  not g72991 (n_32495, n43580);
  and g72992 (n43581, pi1151, n_32495);
  not g72993 (n_32496, n43581);
  and g72994 (n43582, pi0268, n_32496);
  not g72995 (n_32497, n43576);
  and g72996 (n43583, n_32497, n43582);
  not g72997 (n_32498, n43552);
  and g72998 (n43584, n_31652, n_32498);
  not g72999 (n_32499, n43584);
  and g73000 (n43585, n_4226, n_32499);
  not g73001 (n_32500, n43546);
  not g73002 (n_32501, n43585);
  and g73003 (n43586, n_32500, n_32501);
  not g73004 (n_32502, n43586);
  and g73005 (n43587, n_29468, n_32502);
  and g73006 (n43588, n_31868, n43545);
  and g73007 (n43589, n_6791, n41097);
  not g73008 (n_32503, n43530);
  not g73009 (n_32504, n43589);
  and g73010 (n43590, n_32503, n_32504);
  not g73011 (n_32505, n43590);
  and g73012 (n43591, n_4226, n_32505);
  not g73013 (n_32506, n43588);
  and g73014 (n43592, n_32474, n_32506);
  not g73015 (n_32507, n43591);
  and g73016 (n43593, n_32507, n43592);
  not g73017 (n_32508, n43593);
  and g73018 (n43594, pi1151, n_32508);
  not g73019 (n_32509, n43594);
  and g73020 (n43595, n_32480, n_32509);
  not g73021 (n_32510, n43587);
  and g73022 (n43596, n_32510, n43595);
  not g73023 (n_32511, n43596);
  and g73024 (n43597, pi1152, n_32511);
  not g73025 (n_32512, n43583);
  and g73026 (n43598, n_32512, n43597);
  not g73027 (n_32513, n43568);
  not g73028 (n_32514, n43598);
  and g73029 (n43599, n_32513, n_32514);
  not g73030 (n_32515, n43599);
  and g73031 (n43600, pi1150, n_32515);
  and g73032 (n43601, n_31669, n43545);
  not g73033 (n_32516, n41045);
  and g73034 (n43602, n_6791, n_32516);
  not g73035 (n_32517, n43602);
  and g73036 (n43603, n_30530, n_32517);
  and g73037 (n43604, n43591, n43603);
  not g73038 (n_32518, n43601);
  not g73039 (n_32519, n43604);
  and g73040 (n43605, n_32518, n_32519);
  not g73041 (n_32520, n43605);
  and g73042 (n43606, n_29468, n_32520);
  and g73043 (n43607, n_4226, n_32486);
  not g73044 (n_32521, n43607);
  and g73045 (n43608, n_32506, n_32521);
  not g73046 (n_32522, n43608);
  and g73047 (n43609, pi1151, n_32522);
  not g73048 (n_32523, n43606);
  and g73049 (n43610, pi1152, n_32523);
  not g73050 (n_32524, n43609);
  and g73051 (n43611, n_32524, n43610);
  and g73052 (n43612, n_29468, n43562);
  not g73053 (n_32525, n42529);
  and g73054 (n43613, n_32525, n_32476);
  not g73055 (n_32526, n43572);
  and g73056 (n43614, n_32526, n43613);
  and g73057 (n43615, pi1151, n43614);
  not g73058 (n_32527, n43612);
  and g73059 (n43616, n_28873, n_32527);
  not g73060 (n_32528, n43615);
  and g73061 (n43617, n_32528, n43616);
  not g73062 (n_32529, n43611);
  not g73063 (n_32530, n43617);
  and g73064 (n43618, n_32529, n_32530);
  not g73065 (n_32531, n43618);
  and g73066 (n43619, n_32480, n_32531);
  and g73067 (n43620, pi0219, n_32351);
  and g73068 (n43621, n_4226, n_31718);
  not g73069 (n_32532, n43620);
  and g73070 (n43622, n_32532, n43621);
  not g73071 (n_32533, n43622);
  and g73072 (n43623, n_32470, n_32533);
  and g73073 (n43624, n_29468, n43623);
  and g73074 (n43625, n_31697, n43547);
  and g73075 (n43626, n_32471, n_32532);
  not g73076 (n_32534, n43626);
  and g73077 (n43627, n41102, n_32534);
  not g73078 (n_32535, n43627);
  and g73079 (n43628, n_4226, n_32535);
  not g73080 (n_32536, n43625);
  not g73081 (n_32537, n43628);
  and g73082 (n43629, n_32536, n_32537);
  and g73083 (n43630, pi1151, n43629);
  not g73084 (n_32538, n43624);
  and g73085 (n43631, pi1152, n_32538);
  not g73086 (n_32539, n43630);
  and g73087 (n43632, n_32539, n43631);
  and g73088 (n43633, n40874, n_32466);
  not g73089 (n_32540, n43633);
  and g73090 (n43634, n_29468, n_32540);
  not g73091 (n_32541, n42553);
  and g73092 (n43635, n_4226, n_32541);
  and g73093 (n43636, n_32471, n43635);
  not g73094 (n_32542, n42573);
  not g73095 (n_32543, n43636);
  and g73096 (n43637, n_32542, n_32543);
  and g73097 (n43638, pi1151, n43637);
  not g73098 (n_32544, n43634);
  and g73099 (n43639, n_28873, n_32544);
  not g73100 (n_32545, n43638);
  and g73101 (n43640, n_32545, n43639);
  not g73102 (n_32546, n43640);
  and g73103 (n43641, pi0268, n_32546);
  not g73104 (n_32547, n43632);
  and g73105 (n43642, n_32547, n43641);
  not g73106 (n_32548, n43642);
  and g73107 (n43643, n_30133, n_32548);
  not g73108 (n_32549, n43619);
  and g73109 (n43644, n_32549, n43643);
  not g73110 (n_32550, n43600);
  not g73111 (n_32551, n43644);
  and g73112 (n43645, n_32550, n_32551);
  not g73113 (n_32552, n43645);
  and g73114 (n43646, n40909, n_32552);
  not g73115 (n_32553, n43527);
  and g73116 (n43647, n_28510, n_32553);
  not g73117 (n_32554, n43646);
  and g73118 (n43648, n_32554, n43647);
  not g73119 (n_32555, n43505);
  and g73120 (n43649, pi0230, n_32555);
  and g73121 (n43650, n_32449, n43649);
  not g73122 (n_32556, n43648);
  not g73123 (n_32557, n43650);
  and g73124 (po0425, n_32556, n_32557);
  and g73125 (n43652, n_7044, pi1137);
  not g73126 (n_32558, n43652);
  and g73127 (n43653, pi0200, n_32558);
  and g73128 (n43654, pi0199, pi1138);
  and g73129 (n43655, n_7044, pi1136);
  not g73130 (n_32559, n43654);
  and g73131 (n43656, n_7045, n_32559);
  not g73132 (n_32560, n43655);
  and g73133 (n43657, n_32560, n43656);
  not g73134 (n_32561, n43653);
  not g73135 (n_32562, n43657);
  and g73136 (n43658, n_32561, n_32562);
  not g73137 (n_32563, n43658);
  and g73138 (n43659, n16479, n_32563);
  and g73139 (n43660, n_7075, pi1138);
  and g73140 (n43661, pi0219, n43660);
  and g73141 (n43662, pi0211, pi1137);
  not g73142 (n_32564, n43662);
  and g73143 (n43663, n_32222, n_32564);
  not g73144 (n_32565, n43663);
  and g73145 (n43664, n_6791, n_32565);
  not g73146 (n_32566, n43661);
  not g73147 (n_32567, n43664);
  and g73148 (n43665, n_32566, n_32567);
  and g73149 (n43666, n_25711, n43665);
  not g73150 (n_32568, n43659);
  not g73151 (n_32569, n43666);
  and g73152 (n43667, n_32568, n_32569);
  not g73153 (n_32570, n43667);
  and g73154 (n43668, pi0230, n_32570);
  and g73155 (n43669, n_7045, n43254);
  and g73156 (n43670, pi1137, n40951);
  not g73157 (n_32571, n43669);
  not g73158 (n_32572, n43670);
  and g73159 (n43671, n_32571, n_32572);
  and g73160 (n43672, n43500, n43671);
  and g73161 (n43673, pi1091, n_32565);
  not g73162 (n_32573, n43673);
  and g73163 (n43674, n40141, n_32573);
  not g73164 (n_32574, n43672);
  not g73165 (n_32575, n43674);
  and g73166 (n43675, n_32574, n_32575);
  not g73167 (n_32577, pi0817);
  and g73168 (n43676, n_32577, n40885);
  and g73169 (n43677, pi0269, n_32161);
  not g73170 (n_32578, n43676);
  and g73171 (n43678, n_3128, n_32578);
  not g73172 (n_32579, n43677);
  and g73173 (n43679, n_32579, n43678);
  not g73174 (n_32580, n43675);
  not g73175 (n_32581, n43679);
  and g73176 (n43680, n_32580, n_32581);
  and g73177 (n43681, n_32577, n40863);
  and g73178 (n43682, pi0269, n_32156);
  not g73179 (n_32582, n43681);
  and g73180 (n43683, n_3128, n_32582);
  not g73181 (n_32583, n43682);
  and g73182 (n43684, n_32583, n43683);
  and g73183 (n43685, pi1138, n42455);
  and g73184 (n43686, pi0219, n_25711);
  not g73185 (n_32584, n43685);
  and g73186 (n43687, n_32584, n43686);
  and g73187 (n43688, n_7045, pi1091);
  and g73188 (n43689, pi1138, n43688);
  not g73189 (n_32585, n43689);
  and g73190 (n43690, pi0199, n_32585);
  and g73191 (n43691, n16479, n43690);
  not g73192 (n_32586, n43687);
  not g73193 (n_32587, n43691);
  and g73194 (n43692, n_32586, n_32587);
  not g73195 (n_32588, n43684);
  not g73196 (n_32589, n43692);
  and g73197 (n43693, n_32588, n_32589);
  not g73198 (n_32590, n43680);
  not g73199 (n_32591, n43693);
  and g73200 (n43694, n_32590, n_32591);
  not g73201 (n_32592, n43694);
  and g73202 (n43695, n_28510, n_32592);
  not g73203 (n_32593, n43668);
  not g73204 (n_32594, n43695);
  and g73205 (po0426, n_32593, n_32594);
  not g73206 (n_32596, pi0805);
  and g73207 (n43697, n_32596, n40863);
  and g73208 (n43698, pi0270, n_32156);
  not g73209 (n_32597, n43697);
  and g73210 (n43699, n_3128, n_32597);
  not g73211 (n_32598, n43698);
  and g73212 (n43700, n_32598, n43699);
  and g73213 (n43701, n42455, n43168);
  not g73214 (n_32599, n43701);
  and g73215 (n43702, n43686, n_32599);
  and g73216 (n43703, n_7045, n43143);
  not g73217 (n_32600, n43703);
  and g73218 (n43704, pi0199, n_32600);
  and g73219 (n43705, n16479, n43704);
  not g73220 (n_32601, n43702);
  not g73221 (n_32602, n43705);
  and g73222 (n43706, n_32601, n_32602);
  not g73223 (n_32603, n43700);
  not g73224 (n_32604, n43706);
  and g73225 (n43707, n_32603, n_32604);
  and g73226 (n43708, n_32596, n40885);
  and g73227 (n43709, pi0270, n_32161);
  not g73228 (n_32605, n43708);
  and g73229 (n43710, n_3128, n_32605);
  not g73230 (n_32606, n43709);
  and g73231 (n43711, n_32606, n43710);
  and g73232 (n43712, n_7075, pi1139);
  and g73233 (n43713, pi0211, pi1140);
  not g73234 (n_32607, n43712);
  not g73235 (n_32608, n43713);
  and g73236 (n43714, n_32607, n_32608);
  not g73237 (n_32609, n43714);
  and g73238 (n43715, pi1091, n_32609);
  not g73239 (n_32610, n43715);
  and g73240 (n43716, n40141, n_32610);
  and g73241 (n43717, pi1091, pi1140);
  and g73242 (n43718, pi0200, n43717);
  and g73243 (n43719, pi1139, n43688);
  not g73244 (n_32611, n43718);
  not g73245 (n_32612, n43719);
  and g73246 (n43720, n_32611, n_32612);
  and g73247 (n43721, n43500, n43720);
  not g73248 (n_32613, n43716);
  not g73249 (n_32614, n43721);
  and g73250 (n43722, n_32613, n_32614);
  not g73251 (n_32615, n43711);
  not g73252 (n_32616, n43722);
  and g73253 (n43723, n_32615, n_32616);
  not g73254 (n_32617, n43707);
  and g73255 (n43724, n_28510, n_32617);
  not g73256 (n_32618, n43723);
  and g73257 (n43725, n_32618, n43724);
  and g73258 (n43726, pi0219, n_32183);
  and g73259 (n43727, n_6791, n43714);
  not g73260 (n_32619, n43726);
  not g73261 (n_32620, n43727);
  and g73262 (n43728, n_32619, n_32620);
  not g73263 (n_32621, n43728);
  and g73264 (n43729, n_25711, n_32621);
  and g73265 (n43730, n_7044, pi1140);
  not g73266 (n_32622, n43730);
  and g73267 (n43731, pi0200, n_32622);
  and g73268 (n43732, pi0199, pi1141);
  and g73269 (n43733, n_7044, pi1139);
  not g73270 (n_32623, n43732);
  and g73271 (n43734, n_7045, n_32623);
  not g73272 (n_32624, n43733);
  and g73273 (n43735, n_32624, n43734);
  not g73274 (n_32625, n43731);
  not g73275 (n_32626, n43735);
  and g73276 (n43736, n_32625, n_32626);
  not g73277 (n_32627, n43736);
  and g73278 (n43737, n16479, n_32627);
  not g73279 (n_32628, n43729);
  and g73280 (n43738, pi0230, n_32628);
  not g73281 (n_32629, n43737);
  and g73282 (n43739, n_32629, n43738);
  or g73283 (po0427, n43725, n43739);
  and g73284 (n43741, n_7075, pi1147);
  and g73285 (n43742, n42444, n43741);
  not g73286 (n_32630, pi0271);
  and g73287 (n43743, n_32630, n_30430);
  not g73288 (n_32631, n43743);
  and g73289 (n43744, n_30425, n_32631);
  not g73290 (n_32632, n43744);
  and g73291 (n43745, pi0219, n_32632);
  not g73292 (n_32633, n40887);
  and g73293 (n43746, n_3128, n_32633);
  not g73294 (n_32634, n43746);
  and g73295 (n43747, pi0271, n_32634);
  and g73296 (n43748, n_32630, n_30512);
  not g73297 (n_32635, n43747);
  not g73298 (n_32636, n43748);
  and g73299 (n43749, n_32635, n_32636);
  and g73300 (n43750, pi1091, pi1146);
  not g73301 (n_32637, n43749);
  not g73302 (n_32638, n43750);
  and g73303 (n43751, n_32637, n_32638);
  and g73304 (n43752, n_7075, n43750);
  not g73305 (n_32639, n43751);
  not g73306 (n_32640, n43752);
  and g73307 (n43753, n_32639, n_32640);
  and g73308 (n43754, pi1091, n39412);
  not g73309 (n_32641, n43754);
  and g73310 (n43755, n_6791, n_32641);
  not g73311 (n_32642, n43753);
  and g73312 (n43756, n_32642, n43755);
  not g73313 (n_32643, n43745);
  not g73314 (n_32644, n43756);
  and g73315 (n43757, n_32643, n_32644);
  not g73316 (n_32645, n43742);
  and g73317 (n43758, n_25711, n_32645);
  not g73318 (n_32646, n43757);
  and g73319 (n43759, n_32646, n43758);
  and g73320 (n43760, pi0199, n_32632);
  and g73321 (n43761, n_7044, n43751);
  not g73322 (n_32647, n43760);
  not g73323 (n_32648, n43761);
  and g73324 (n43762, n_32647, n_32648);
  not g73325 (n_32649, n43762);
  and g73326 (n43763, pi0200, n_32649);
  and g73327 (n43764, pi1147, n40931);
  and g73328 (n43765, pi1091, pi1145);
  not g73329 (n_32650, n43765);
  and g73330 (n43766, n_7044, n_32650);
  and g73331 (n43767, n_32637, n43766);
  not g73332 (n_32651, n43767);
  and g73333 (n43768, n_32647, n_32651);
  not g73334 (n_32652, n43764);
  and g73335 (n43769, n_7045, n_32652);
  not g73336 (n_32653, n43768);
  and g73337 (n43770, n_32653, n43769);
  not g73338 (n_32654, n43763);
  not g73339 (n_32655, n43770);
  and g73340 (n43771, n_32654, n_32655);
  not g73341 (n_32656, n43771);
  and g73342 (n43772, n16479, n_32656);
  not g73343 (n_32657, n43759);
  not g73344 (n_32658, n43772);
  and g73345 (n43773, n_32657, n_32658);
  not g73346 (n_32659, n43773);
  and g73347 (n43774, n_28510, n_32659);
  and g73348 (n43775, pi1147, n42386);
  and g73349 (n43776, n_29922, n_29928);
  not g73350 (n_32660, n43776);
  and g73351 (n43777, n_6791, n_32660);
  and g73352 (n43778, n_7045, n_29278);
  not g73353 (n_32661, n43778);
  and g73354 (n43779, n40339, n_32661);
  not g73355 (n_32662, n43775);
  not g73356 (n_32663, n43777);
  and g73357 (n43780, n_32662, n_32663);
  not g73358 (n_32664, n43779);
  and g73359 (n43781, n_32664, n43780);
  not g73360 (n_32665, n43781);
  and g73361 (n43782, n_4226, n_32665);
  not g73362 (n_32666, n43741);
  and g73363 (n43783, pi0219, n_32666);
  and g73364 (n43784, n_29294, n41531);
  not g73365 (n_32667, n43783);
  not g73366 (n_32668, n43784);
  and g73367 (n43785, n_32667, n_32668);
  and g73368 (n43786, po1038, n43785);
  not g73369 (n_32669, n43786);
  and g73370 (n43787, pi0230, n_32669);
  not g73371 (n_32670, n43782);
  and g73372 (n43788, n_32670, n43787);
  not g73373 (n_32671, n43774);
  not g73374 (n_32672, n43788);
  and g73375 (po0428, n_32671, n_32672);
  and g73376 (n43790, po1038, n10844);
  not g73377 (n_32673, n13065);
  not g73378 (n_32674, n43790);
  and g73379 (n43791, n_32673, n_32674);
  and g73380 (n43792, n_30133, n43791);
  not g73381 (n_32675, n43792);
  and g73382 (n43793, n_32433, n_32675);
  not g73383 (n_32676, n43793);
  and g73384 (n43794, n_29850, n_32676);
  and g73385 (n43795, pi1149, n_30133);
  not g73386 (n_32677, n43795);
  and g73387 (n43796, n_32433, n_32677);
  not g73388 (n_32678, n43796);
  and g73389 (n43797, n43501, n_32678);
  not g73390 (n_32679, n43794);
  not g73391 (n_32680, n43797);
  and g73392 (n43798, n_32679, n_32680);
  not g73393 (n_32681, n43798);
  and g73394 (n43799, pi1091, n_32681);
  not g73395 (n_32682, n43799);
  and g73396 (n43800, pi1148, n_32682);
  and g73397 (n43801, pi1150, n_31565);
  not g73398 (n_32683, n43801);
  and g73399 (n43802, n_29850, n_32683);
  and g73400 (n43803, pi1091, n43802);
  and g73401 (n43804, n_25711, n42712);
  and g73402 (n43805, n_4226, n40936);
  not g73403 (n_32684, n43804);
  not g73404 (n_32685, n43805);
  and g73405 (n43806, n_32684, n_32685);
  and g73406 (n43807, n_30133, n43806);
  and g73407 (n43808, pi1091, n_32444);
  not g73408 (n_32686, n43808);
  and g73409 (n43809, pi1150, n_32686);
  not g73410 (n_32687, n43807);
  and g73411 (n43810, pi1149, n_32687);
  not g73412 (n_32688, n43809);
  and g73413 (n43811, n_32688, n43810);
  not g73414 (n_32689, n43803);
  and g73415 (n43812, n_29904, n_32689);
  not g73416 (n_32690, n43811);
  and g73417 (n43813, n_32690, n43812);
  not g73418 (n_32691, pi0283);
  not g73419 (n_32692, n43800);
  and g73420 (n43814, n_32691, n_32692);
  not g73421 (n_32693, n43813);
  and g73422 (n43815, n_32693, n43814);
  and g73423 (n43816, n_30133, n_32540);
  and g73424 (n43817, pi1150, n43623);
  not g73425 (n_32694, n43816);
  and g73426 (n43818, n_29850, n_32694);
  not g73427 (n_32695, n43817);
  and g73428 (n43819, n_32695, n43818);
  and g73429 (n43820, pi1150, n43629);
  and g73430 (n43821, n_30133, n43637);
  not g73431 (n_32696, n43821);
  and g73432 (n43822, pi1149, n_32696);
  not g73433 (n_32697, n43820);
  and g73434 (n43823, n_32697, n43822);
  not g73435 (n_32698, n43819);
  not g73436 (n_32699, n43823);
  and g73437 (n43824, n_32698, n_32699);
  not g73438 (n_32700, n43824);
  and g73439 (n43825, n_29904, n_32700);
  and g73440 (n43826, n_30133, n43541);
  and g73441 (n43827, pi1150, n43580);
  not g73442 (n_32701, n43826);
  and g73443 (n43828, pi1149, n_32701);
  not g73444 (n_32702, n43827);
  and g73445 (n43829, n_32702, n43828);
  and g73446 (n43830, n_30133, n43535);
  and g73447 (n43831, pi1150, n43575);
  not g73448 (n_32703, n43830);
  and g73449 (n43832, n_29850, n_32703);
  not g73450 (n_32704, n43831);
  and g73451 (n43833, n_32704, n43832);
  not g73452 (n_32705, n43829);
  not g73453 (n_32706, n43833);
  and g73454 (n43834, n_32705, n_32706);
  not g73455 (n_32707, n43834);
  and g73456 (n43835, pi1148, n_32707);
  not g73457 (n_32708, n43825);
  and g73458 (n43836, pi0283, n_32708);
  not g73459 (n_32709, n43835);
  and g73460 (n43837, n_32709, n43836);
  not g73461 (n_32710, n43815);
  and g73462 (n43838, pi0272, n_32710);
  not g73463 (n_32711, n43837);
  and g73464 (n43839, n_32711, n43838);
  not g73465 (n_32712, n43563);
  and g73466 (n43840, n_30133, n_32712);
  and g73467 (n43841, pi1150, n_32508);
  not g73468 (n_32713, n43840);
  and g73469 (n43842, pi1149, n_32713);
  not g73470 (n_32714, n43841);
  and g73471 (n43843, n_32714, n43842);
  and g73472 (n43844, pi1150, n_32502);
  not g73473 (n_32715, n43555);
  and g73474 (n43845, n_30133, n_32715);
  not g73475 (n_32716, n43845);
  and g73476 (n43846, n_29850, n_32716);
  not g73477 (n_32717, n43844);
  and g73478 (n43847, n_32717, n43846);
  not g73479 (n_32718, n43843);
  not g73480 (n_32719, n43847);
  and g73481 (n43848, n_32718, n_32719);
  not g73482 (n_32720, n43848);
  and g73483 (n43849, pi1148, n_32720);
  and g73484 (n43850, pi1150, n43605);
  and g73485 (n43851, n_30133, n_32479);
  not g73486 (n_32721, n43851);
  and g73487 (n43852, n_29850, n_32721);
  not g73488 (n_32722, n43850);
  and g73489 (n43853, n_32722, n43852);
  not g73490 (n_32723, n43614);
  and g73491 (n43854, n_30133, n_32723);
  and g73492 (n43855, pi1150, n43608);
  not g73493 (n_32724, n43855);
  and g73494 (n43856, pi1149, n_32724);
  not g73495 (n_32725, n43854);
  and g73496 (n43857, n_32725, n43856);
  not g73497 (n_32726, n43853);
  and g73498 (n43858, n_29904, n_32726);
  not g73499 (n_32727, n43857);
  and g73500 (n43859, n_32727, n43858);
  not g73501 (n_32728, n43849);
  not g73502 (n_32729, n43859);
  and g73503 (n43860, n_32728, n_32729);
  not g73504 (n_32730, n43860);
  and g73505 (n43861, pi0283, n_32730);
  and g73506 (n43862, n_4226, n38550);
  not g73507 (n_32731, n43862);
  and g73508 (n43863, n_32431, n_32731);
  and g73509 (n43864, n_32429, n43863);
  not g73510 (n_32732, n43864);
  and g73511 (n43865, pi1150, n_32732);
  not g73512 (n_32733, n43865);
  and g73513 (n43866, pi1149, n_32733);
  and g73514 (n43867, n43501, n43866);
  and g73515 (n43868, pi1148, n_32679);
  not g73516 (n_32734, n43867);
  and g73517 (n43869, n_32734, n43868);
  and g73518 (n43870, pi1091, n43869);
  not g73519 (n_32735, n43802);
  and g73520 (n43871, n_29904, n_32735);
  and g73521 (n43872, n_30133, n_32440);
  and g73522 (n43873, pi1150, n43515);
  not g73523 (n_32736, n43872);
  and g73524 (n43874, pi1149, n_32736);
  not g73525 (n_32737, n43873);
  and g73526 (n43875, n_32737, n43874);
  not g73527 (n_32738, n43875);
  and g73528 (n43876, pi1091, n_32738);
  and g73529 (n43877, n43871, n43876);
  not g73530 (n_32739, n43877);
  and g73531 (n43878, n_32691, n_32739);
  not g73532 (n_32740, n43870);
  and g73533 (n43879, n_32740, n43878);
  not g73534 (n_32741, pi0272);
  not g73535 (n_32742, n43879);
  and g73536 (n43880, n_32741, n_32742);
  not g73537 (n_32743, n43861);
  and g73538 (n43881, n_32743, n43880);
  not g73539 (n_32744, n43839);
  and g73540 (n43882, n_28510, n_32744);
  not g73541 (n_32745, n43881);
  and g73542 (n43883, n_32745, n43882);
  and g73543 (n43884, pi1149, n_32444);
  not g73544 (n_32746, n43866);
  not g73545 (n_32747, n43884);
  and g73546 (n43885, n_32746, n_32747);
  not g73547 (n_32748, n43885);
  and g73548 (n43886, n_32736, n_32748);
  not g73549 (n_32749, n43886);
  and g73550 (n43887, n43871, n_32749);
  not g73551 (n_32750, n43869);
  and g73552 (n43888, pi0230, n_32750);
  not g73553 (n_32751, n43887);
  and g73554 (n43889, n_32751, n43888);
  not g73555 (n_32752, n43883);
  not g73556 (n_32753, n43889);
  and g73557 (po0429, n_32752, n_32753);
  not g73558 (n_32754, pi0273);
  not g73559 (n_32755, n40867);
  and g73560 (n43891, n_32754, n_32755);
  not g73561 (n_32756, n43891);
  and g73562 (n43892, n_30427, n_32756);
  not g73563 (n_32757, n43892);
  and g73564 (n43893, pi0219, n_32757);
  not g73565 (n_32758, n40889);
  and g73566 (n43894, n_32754, n_32758);
  not g73567 (n_32759, n43894);
  and g73568 (n43895, n40891, n_32759);
  and g73569 (n43896, n_6791, n_32640);
  not g73570 (n_32760, n43895);
  and g73571 (n43897, n_32760, n43896);
  not g73572 (n_32761, n43893);
  not g73573 (n_32762, n43897);
  and g73574 (n43898, n_32761, n_32762);
  and g73575 (n43899, po1038, n43898);
  and g73576 (n43900, pi0299, n43898);
  and g73577 (n43901, pi0199, n_32757);
  and g73578 (n43902, n_7045, n43750);
  not g73579 (n_32763, n43902);
  and g73580 (n43903, n_7044, n_32763);
  and g73581 (n43904, n_32760, n43903);
  not g73582 (n_32764, n43901);
  and g73583 (n43905, n_234, n_32764);
  not g73584 (n_32765, n43904);
  and g73585 (n43906, n_32765, n43905);
  not g73586 (n_32766, n43900);
  not g73587 (n_32767, n43906);
  and g73588 (n43907, n_32766, n_32767);
  and g73589 (n43908, n_7410, n_30560);
  not g73590 (n_32768, n43908);
  and g73591 (n43909, pi1091, n_32768);
  not g73592 (n_32769, n43909);
  and g73593 (n43910, n43907, n_32769);
  not g73594 (n_32770, n43910);
  and g73595 (n43911, n_4226, n_32770);
  and g73596 (n43912, pi1091, n42573);
  not g73597 (n_32771, n43911);
  not g73598 (n_32772, n43912);
  and g73599 (n43913, n_32771, n_32772);
  not g73600 (n_32773, n43913);
  and g73601 (n43914, pi1147, n_32773);
  not g73602 (n_32774, n43907);
  and g73603 (n43915, n40447, n_32774);
  not g73604 (n_32775, n43915);
  and g73605 (n43916, n_29904, n_32775);
  and g73606 (n43917, pi1091, n38519);
  not g73607 (n_32776, n43898);
  not g73608 (n_32777, n43917);
  and g73609 (n43918, n_32776, n_32777);
  not g73610 (n_32778, n43918);
  and g73611 (n43919, pi0299, n_32778);
  and g73612 (n43920, n40932, n_32654);
  not g73613 (n_32779, n43920);
  and g73614 (n43921, n_32767, n_32779);
  not g73615 (n_32780, n43919);
  and g73616 (n43922, n_32780, n43921);
  not g73617 (n_32781, n43922);
  and g73618 (n43923, n_4226, n_32781);
  and g73619 (n43924, n40080, n42444);
  not g73620 (n_32782, n43924);
  and g73621 (n43925, pi1148, n_32782);
  not g73622 (n_32783, n43923);
  and g73623 (n43926, n_32783, n43925);
  not g73624 (n_32784, n43916);
  not g73625 (n_32785, n43926);
  and g73626 (n43927, n_32784, n_32785);
  not g73627 (n_32786, n43899);
  not g73628 (n_32787, n43927);
  and g73629 (n43928, n_32786, n_32787);
  not g73630 (n_32788, n43914);
  and g73631 (n43929, n_32788, n43928);
  not g73632 (n_32789, n43929);
  and g73633 (n43930, n_28510, n_32789);
  not g73634 (n_32790, n41404);
  and g73635 (n43931, pi1146, n_32790);
  not g73636 (n_32791, n43791);
  and g73637 (n43932, n_32791, n43931);
  and g73638 (n43933, n_7075, n_29958);
  not g73639 (n_32792, n43933);
  and g73640 (n43934, n40141, n_32792);
  and g73641 (n43935, n_803, n10809);
  not g73642 (n_32793, n43935);
  and g73643 (n43936, n43500, n_32793);
  not g73644 (n_32794, n43934);
  not g73645 (n_32795, n43936);
  and g73646 (n43937, n_32794, n_32795);
  not g73647 (n_32796, n43937);
  and g73648 (n43938, pi1147, n_32796);
  not g73649 (n_32797, n43932);
  and g73650 (n43939, n_29904, n_32797);
  not g73651 (n_32798, n43938);
  and g73652 (n43940, n_32798, n43939);
  and g73653 (n43941, n_7044, pi1147);
  not g73654 (n_32799, n43941);
  and g73655 (n43942, pi0200, n_32799);
  not g73656 (n_32800, n43942);
  and g73657 (n43943, n_32793, n_32800);
  and g73658 (n43944, n16479, n43943);
  and g73659 (n43945, n_803, n10844);
  and g73660 (n43946, pi1147, n40141);
  not g73661 (n_32801, n43946);
  and g73662 (n43947, n_32429, n_32801);
  not g73663 (n_32802, n43945);
  not g73664 (n_32803, n43947);
  and g73665 (n43948, n_32802, n_32803);
  not g73666 (n_32804, n43944);
  and g73667 (n43949, pi1148, n_32804);
  not g73668 (n_32805, n43948);
  and g73669 (n43950, n_32805, n43949);
  not g73670 (n_32806, n43940);
  and g73671 (n43951, pi0230, n_32806);
  not g73672 (n_32807, n43950);
  and g73673 (n43952, n_32807, n43951);
  or g73674 (po0430, n43930, n43952);
  and g73675 (n43954, n_7045, n43765);
  not g73676 (n_32809, pi0659);
  and g73677 (n43955, n_32809, n40863);
  and g73678 (n43956, pi0274, n_32156);
  not g73679 (n_32810, n43955);
  and g73680 (n43957, n_3128, n_32810);
  not g73681 (n_32811, n43956);
  and g73682 (n43958, n_32811, n43957);
  not g73683 (n_32812, n43954);
  and g73684 (n43959, pi0199, n_32812);
  not g73685 (n_32813, n43958);
  and g73686 (n43960, n_32813, n43959);
  and g73687 (n43961, n_32809, n40885);
  and g73688 (n43962, pi0274, n_32161);
  not g73689 (n_32814, n43961);
  and g73690 (n43963, n_3128, n_32814);
  not g73691 (n_32815, n43962);
  and g73692 (n43964, n_32815, n43963);
  not g73693 (n_32816, n43180);
  not g73694 (n_32817, n43964);
  and g73695 (n43965, n_32816, n_32817);
  not g73696 (n_32818, n43965);
  and g73697 (n43966, pi0200, n_32818);
  and g73698 (n43967, n_32201, n_32817);
  not g73699 (n_32819, n43967);
  and g73700 (n43968, n_7045, n_32819);
  not g73701 (n_32820, n43966);
  and g73702 (n43969, n_7044, n_32820);
  not g73703 (n_32821, n43968);
  and g73704 (n43970, n_32821, n43969);
  not g73705 (n_32822, n43960);
  and g73706 (n43971, n16479, n_32822);
  not g73707 (n_32823, n43970);
  and g73708 (n43972, n_32823, n43971);
  and g73709 (n43973, pi0211, n_32818);
  and g73710 (n43974, n_7075, n_32819);
  not g73711 (n_32824, n43973);
  and g73712 (n43975, n_6791, n_32824);
  not g73713 (n_32825, n43974);
  and g73714 (n43976, n_32825, n43975);
  and g73715 (n43977, pi0219, n_32641);
  and g73716 (n43978, n_32813, n43977);
  not g73717 (n_32826, n43978);
  and g73718 (n43979, n_25711, n_32826);
  not g73719 (n_32827, n43976);
  and g73720 (n43980, n_32827, n43979);
  not g73721 (n_32828, n43972);
  and g73722 (n43981, n_28510, n_32828);
  not g73723 (n_32829, n43980);
  and g73724 (n43982, n_32829, n43981);
  and g73725 (n43983, n_31562, n_29922);
  and g73726 (n43984, n_6791, n_28544);
  and g73727 (n43985, n_29295, n43984);
  not g73728 (n_32830, n43983);
  not g73729 (n_32831, n43985);
  and g73730 (n43986, n_32830, n_32831);
  and g73731 (n43987, n_28528, n40332);
  not g73732 (n_32832, n43987);
  and g73733 (n43988, n40788, n_32832);
  not g73734 (n_32833, n43986);
  not g73735 (n_32834, n43988);
  and g73736 (n43989, n_32833, n_32834);
  not g73737 (n_32835, n43989);
  and g73738 (n43990, n_4226, n_32835);
  and g73739 (n43991, n_29919, n_32831);
  not g73740 (n_32836, n43990);
  and g73741 (n43992, pi0230, n_32836);
  not g73742 (n_32837, n43991);
  and g73743 (n43993, n_32837, n43992);
  not g73744 (n_32838, n43982);
  not g73745 (n_32839, n43993);
  and g73746 (po0431, n_32838, n_32839);
  and g73747 (n43995, pi1151, n_32433);
  and g73748 (n43996, pi1149, n43501);
  not g73749 (n_32840, n43995);
  and g73750 (n43997, n_32840, n43996);
  and g73751 (n43998, n_29850, n43516);
  not g73752 (n_32841, n43997);
  not g73753 (n_32842, n43998);
  and g73754 (n43999, n_32841, n_32842);
  not g73755 (n_32843, n43999);
  and g73756 (n44000, pi1150, n_32843);
  and g73757 (n44001, n_29468, n43791);
  and g73758 (n44002, pi1149, n_32433);
  not g73759 (n_32844, n44001);
  and g73760 (n44003, n_32844, n44002);
  and g73761 (n44004, n_29850, pi1151);
  and g73762 (n44005, n_31565, n44004);
  not g73763 (n_32845, n44005);
  and g73764 (n44006, n_30133, n_32845);
  not g73765 (n_32846, n44003);
  and g73766 (n44007, n_32846, n44006);
  not g73767 (n_32847, n44000);
  not g73768 (n_32848, n44007);
  and g73769 (n44008, n_32847, n_32848);
  not g73770 (n_32849, n44008);
  and g73771 (n44009, pi1091, n_32849);
  and g73772 (n44010, n_29468, n41484);
  not g73773 (n_32850, n43806);
  and g73774 (n44011, n_32850, n44010);
  not g73775 (n_32851, n44009);
  not g73776 (n_32852, n44011);
  and g73777 (n44012, n_32851, n_32852);
  not g73778 (n_32853, n44012);
  and g73779 (n44013, pi0275, n_32853);
  and g73780 (n44014, n43498, n43795);
  and g73781 (n44015, n40607, n_31565);
  and g73782 (n44016, n_29468, n43510);
  not g73783 (n_32854, n44016);
  and g73784 (n44017, pi1150, n_32854);
  not g73785 (n_32855, n43516);
  and g73786 (n44018, n_32855, n44017);
  not g73787 (n_32856, n44015);
  and g73788 (n44019, n_29850, n_32856);
  not g73789 (n_32857, n44018);
  and g73790 (n44020, n_32857, n44019);
  not g73791 (n_32858, n44014);
  and g73792 (n44021, n_32841, n_32858);
  not g73793 (n_32859, n44020);
  and g73794 (n44022, n_32859, n44021);
  and g73795 (n44023, pi1091, n44022);
  not g73796 (n_32860, pi0275);
  not g73797 (n_32861, n44023);
  and g73798 (n44024, n_32860, n_32861);
  not g73799 (n_32862, n40908);
  not g73800 (n_32863, n44024);
  and g73801 (n44025, n_32862, n_32863);
  not g73802 (n_32864, n44013);
  and g73803 (n44026, n_32864, n44025);
  and g73804 (n44027, n_30133, n43605);
  and g73805 (n44028, pi1151, n_32724);
  not g73806 (n_32865, n44027);
  and g73807 (n44029, n_32865, n44028);
  and g73808 (n44030, pi1150, n_32723);
  and g73809 (n44031, n_29468, n_32721);
  not g73810 (n_32866, n44030);
  and g73811 (n44032, n_32866, n44031);
  not g73812 (n_32867, n44029);
  not g73813 (n_32868, n44032);
  and g73814 (n44033, n_32867, n_32868);
  not g73815 (n_32869, n44033);
  and g73816 (n44034, n_32860, n_32869);
  and g73817 (n44035, pi1150, n43637);
  not g73818 (n_32870, n44035);
  and g73819 (n44036, n_32694, n_32870);
  not g73820 (n_32871, n44036);
  and g73821 (n44037, n_29468, n_32871);
  and g73822 (n44038, n_30133, n43623);
  not g73823 (n_32872, n44038);
  and g73824 (n44039, n_32697, n_32872);
  not g73825 (n_32873, n44039);
  and g73826 (n44040, pi1151, n_32873);
  not g73827 (n_32874, n44037);
  and g73828 (n44041, pi0275, n_32874);
  not g73829 (n_32875, n44040);
  and g73830 (n44042, n_32875, n44041);
  not g73831 (n_32876, n44042);
  and g73832 (n44043, n_29850, n_32876);
  not g73833 (n_32877, n44034);
  and g73834 (n44044, n_32877, n44043);
  and g73835 (n44045, pi1150, n_32712);
  not g73836 (n_32878, n44045);
  and g73837 (n44046, n_29468, n_32878);
  and g73838 (n44047, n_32716, n44046);
  and g73839 (n44048, n_30133, n_32502);
  and g73840 (n44049, pi1151, n_32714);
  not g73841 (n_32879, n44048);
  and g73842 (n44050, n_32879, n44049);
  not g73843 (n_32880, n44047);
  and g73844 (n44051, n_32860, n_32880);
  not g73845 (n_32881, n44050);
  and g73846 (n44052, n_32881, n44051);
  and g73847 (n44053, pi1151, n_32492);
  and g73848 (n44054, n_30133, n_32467);
  not g73849 (n_32882, n44053);
  and g73850 (n44055, n_32882, n44054);
  and g73851 (n44056, n_29468, n_32466);
  not g73852 (n_32883, n44056);
  and g73853 (n44057, pi1150, n_32883);
  and g73854 (n44058, n_32496, n44057);
  not g73855 (n_32884, n44058);
  and g73856 (n44059, pi0275, n_32884);
  not g73857 (n_32885, n44055);
  and g73858 (n44060, n_32885, n44059);
  not g73859 (n_32886, n44052);
  and g73860 (n44061, pi1149, n_32886);
  not g73861 (n_32887, n44060);
  and g73862 (n44062, n_32887, n44061);
  not g73863 (n_32888, n44044);
  and g73864 (n44063, n40908, n_32888);
  not g73865 (n_32889, n44062);
  and g73866 (n44064, n_32889, n44063);
  not g73867 (n_32890, n44026);
  not g73868 (n_32891, n44064);
  and g73869 (n44065, n_32890, n_32891);
  not g73870 (n_32892, n44065);
  and g73871 (n44066, n_28510, n_32892);
  and g73872 (n44067, pi0230, n44022);
  or g73873 (po0432, n44066, n44067);
  not g73874 (n_32893, n40886);
  and g73875 (n44069, n_930, n_32893);
  not g73876 (n_32894, n44069);
  and g73877 (n44070, n43746, n_32894);
  and g73878 (n44071, n_28515, n_29910);
  not g73879 (n_32895, n44071);
  and g73880 (n44072, pi1091, n_32895);
  not g73881 (n_32896, n44072);
  and g73882 (n44073, n40141, n_32896);
  and g73883 (n44074, pi1145, n40951);
  not g73884 (n_32897, n44074);
  and g73885 (n44075, n_32195, n_32897);
  and g73886 (n44076, n43500, n44075);
  not g73887 (n_32898, n44073);
  not g73888 (n_32899, n44076);
  and g73889 (n44077, n_32898, n_32899);
  not g73890 (n_32900, n44070);
  not g73891 (n_32901, n44077);
  and g73892 (n44078, n_32900, n_32901);
  not g73893 (n_32902, n40864);
  and g73894 (n44079, n_930, n_32902);
  not g73895 (n_32903, n44079);
  and g73896 (n44080, n40870, n_32903);
  and g73897 (n44081, n43686, n_32640);
  and g73898 (n44082, pi0199, n_32763);
  and g73899 (n44083, n16479, n44082);
  not g73900 (n_32904, n44081);
  not g73901 (n_32905, n44083);
  and g73902 (n44084, n_32904, n_32905);
  not g73903 (n_32906, n44080);
  not g73904 (n_32907, n44084);
  and g73905 (n44085, n_32906, n_32907);
  not g73906 (n_32908, n44078);
  and g73907 (n44086, n_28510, n_32908);
  not g73908 (n_32909, n44085);
  and g73909 (n44087, n_32909, n44086);
  and g73910 (n44088, n_28527, n41294);
  not g73911 (n_32910, n44088);
  and g73912 (n44089, n_30005, n_32910);
  not g73913 (n_32911, n44089);
  and g73914 (n44090, n16479, n_32911);
  and g73915 (n44091, n_6791, n_32895);
  and g73916 (n44092, pi1146, n38519);
  not g73917 (n_32912, n44091);
  not g73918 (n_32913, n44092);
  and g73919 (n44093, n_32912, n_32913);
  and g73920 (n44094, n_25711, n44093);
  not g73921 (n_32914, n44090);
  and g73922 (n44095, pi0230, n_32914);
  not g73923 (n_32915, n44094);
  and g73924 (n44096, n_32915, n44095);
  or g73925 (po0433, n44087, n44096);
  and g73926 (n44098, n_7045, n43150);
  not g73927 (n_32917, pi0820);
  and g73928 (n44099, n_32917, n40863);
  and g73929 (n44100, pi0277, n_32156);
  not g73930 (n_32918, n44099);
  and g73931 (n44101, n_3128, n_32918);
  not g73932 (n_32919, n44100);
  and g73933 (n44102, n_32919, n44101);
  not g73934 (n_32920, n44098);
  and g73935 (n44103, pi0199, n_32920);
  not g73936 (n_32921, n44102);
  and g73937 (n44104, n_32921, n44103);
  and g73938 (n44105, n_32917, n40885);
  and g73939 (n44106, pi0277, n_32161);
  not g73940 (n_32922, n44105);
  and g73941 (n44107, n_3128, n_32922);
  not g73942 (n_32923, n44106);
  and g73943 (n44108, n_32923, n44107);
  not g73944 (n_32924, n43717);
  not g73945 (n_32925, n44108);
  and g73946 (n44109, n_32924, n_32925);
  not g73947 (n_32926, n44109);
  and g73948 (n44110, n_7045, n_32926);
  and g73949 (n44111, n_32164, n_32925);
  not g73950 (n_32927, n44111);
  and g73951 (n44112, pi0200, n_32927);
  not g73952 (n_32928, n44110);
  and g73953 (n44113, n_7044, n_32928);
  not g73954 (n_32929, n44112);
  and g73955 (n44114, n_32929, n44113);
  not g73956 (n_32930, n44104);
  and g73957 (n44115, n16479, n_32930);
  not g73958 (n_32931, n44114);
  and g73959 (n44116, n_32931, n44115);
  and g73960 (n44117, pi0219, n_32215);
  not g73961 (n_32932, n44117);
  and g73962 (n44118, n_32174, n_32932);
  not g73963 (n_32933, n44118);
  and g73964 (n44119, n_32921, n_32933);
  and g73965 (n44120, n_7075, n_32926);
  and g73966 (n44121, pi0211, n_32927);
  not g73967 (n_32934, n44120);
  and g73968 (n44122, n_6791, n_32934);
  not g73969 (n_32935, n44121);
  and g73970 (n44123, n_32935, n44122);
  not g73971 (n_32936, n44119);
  and g73972 (n44124, n_25711, n_32936);
  not g73973 (n_32937, n44123);
  and g73974 (n44125, n_32937, n44124);
  not g73975 (n_32938, n44116);
  not g73976 (n_32939, n44125);
  and g73977 (n44126, n_32938, n_32939);
  not g73978 (n_32940, n44126);
  and g73979 (n44127, n_28510, n_32940);
  and g73980 (n44128, pi0211, pi1141);
  and g73981 (n44129, n_7075, pi1140);
  not g73982 (n_32941, n44128);
  and g73983 (n44130, n_6791, n_32941);
  not g73984 (n_32942, n44129);
  and g73985 (n44131, n_32942, n44130);
  not g73986 (n_32943, n44131);
  and g73987 (n44132, n_32932, n_32943);
  not g73988 (n_32944, n44132);
  and g73989 (n44133, n_25711, n_32944);
  and g73990 (n44134, n38433, n_32622);
  and g73991 (n44135, pi0200, n_32186);
  not g73992 (n_32945, n44134);
  not g73993 (n_32946, n44135);
  and g73994 (n44136, n_32945, n_32946);
  not g73995 (n_32947, n44136);
  and g73996 (n44137, n16479, n_32947);
  not g73997 (n_32948, n44133);
  and g73998 (n44138, pi0230, n_32948);
  not g73999 (n_32949, n44137);
  and g74000 (n44139, n_32949, n44138);
  or g74001 (po0434, n44127, n44139);
  not g74002 (po1130, pi0278);
  and g74003 (n44141, po1130, n_32156);
  not g74004 (n_32952, pi0976);
  and g74005 (n44142, n_32952, n40863);
  not g74006 (n_32953, n44141);
  and g74007 (n44143, n_3128, n_32953);
  not g74008 (n_32954, n44142);
  and g74009 (n44144, n_32954, n44143);
  not g74010 (n_32955, n44144);
  and g74011 (n44145, pi0199, n_32955);
  not g74012 (n_32957, pi1132);
  and g74013 (n44146, pi1091, n_32957);
  and g74014 (n44147, pi0976, n40885);
  and g74015 (n44148, pi0278, n_32161);
  not g74016 (n_32958, n44147);
  and g74017 (n44149, n_3128, n_32958);
  not g74018 (n_32959, n44148);
  and g74019 (n44150, n_32959, n44149);
  not g74020 (n_32960, n44146);
  not g74021 (n_32961, n44150);
  and g74022 (n44151, n_32960, n_32961);
  not g74023 (n_32962, n44151);
  and g74024 (n44152, n_7044, n_32962);
  not g74025 (n_32963, n44145);
  not g74026 (n_32964, n44152);
  and g74027 (n44153, n_32963, n_32964);
  not g74028 (n_32965, n44153);
  and g74029 (n44154, n_7045, n_32965);
  not g74030 (n_32967, pi1133);
  and g74031 (n44155, pi1091, n_32967);
  not g74032 (n_32968, n44155);
  and g74033 (n44156, n_32961, n_32968);
  not g74034 (n_32969, n44156);
  and g74035 (n44157, n_7044, n_32969);
  not g74036 (n_32970, n44157);
  and g74037 (n44158, n_32963, n_32970);
  not g74038 (n_32971, n44158);
  and g74039 (n44159, pi0200, n_32971);
  not g74040 (n_32972, n44159);
  and g74041 (n44160, n_234, n_32972);
  not g74042 (n_32973, n44154);
  and g74043 (n44161, n_32973, n44160);
  and g74044 (n44162, pi0219, n_32955);
  and g74045 (n44163, pi0211, n_32967);
  and g74046 (n44164, n_7075, n_32957);
  not g74047 (n_32974, n44163);
  not g74048 (n_32975, n44164);
  and g74049 (n44165, n_32974, n_32975);
  not g74050 (n_32976, n44165);
  and g74051 (n44166, pi1091, n_32976);
  not g74052 (n_32977, n44166);
  and g74053 (n44167, n_32961, n_32977);
  not g74054 (n_32978, n44167);
  and g74055 (n44168, n_6791, n_32978);
  not g74056 (n_32979, n44162);
  not g74057 (n_32980, n44168);
  and g74058 (n44169, n_32979, n_32980);
  and g74059 (n44170, pi0299, n44169);
  not g74060 (n_32981, n44161);
  not g74061 (n_32982, n44170);
  and g74062 (n44171, n_32981, n_32982);
  not g74063 (n_32983, n44171);
  and g74064 (n44172, n_4226, n_32983);
  and g74065 (n44173, po1038, n44169);
  not g74066 (n_32984, n44173);
  and g74067 (n44174, n_28510, n_32984);
  not g74068 (n_32985, n44172);
  and g74069 (n44175, n_32985, n44174);
  and g74070 (n44176, n39374, n44165);
  and g74071 (n44177, n_7044, pi1132);
  not g74072 (n_32986, n44177);
  and g74073 (n44178, n_7045, n_32986);
  and g74074 (n44179, n_7044, pi1133);
  not g74075 (n_32987, n44179);
  and g74076 (n44180, pi0200, n_32987);
  not g74077 (n_32988, n44180);
  and g74078 (n44181, n_234, n_32988);
  not g74079 (n_32989, n44178);
  and g74080 (n44182, n_32989, n44181);
  and g74081 (n44183, n38508, n44165);
  not g74082 (n_32990, n44182);
  not g74083 (n_32991, n44183);
  and g74084 (n44184, n_32990, n_32991);
  not g74085 (n_32992, n44184);
  and g74086 (n44185, n_4226, n_32992);
  not g74087 (n_32993, n44176);
  and g74088 (n44186, pi0230, n_32993);
  not g74089 (n_32994, n44185);
  and g74090 (n44187, n_32994, n44186);
  not g74091 (n_32995, n44175);
  not g74092 (n_32996, n44187);
  and g74093 (n44188, n_32995, n_32996);
  not g74094 (n_32997, n44188);
  and g74095 (n44189, n_2921, n_32997);
  and g74096 (n44190, n10809, n_32986);
  not g74097 (n_32998, n44190);
  and g74098 (n44191, n44181, n_32998);
  and g74099 (n44192, n_31739, n_32991);
  not g74100 (n_32999, n44191);
  and g74101 (n44193, n_32999, n44192);
  not g74102 (n_33000, n44193);
  and g74103 (n44194, n_4226, n_33000);
  and g74104 (n44195, n_6791, n_32976);
  not g74105 (n_33001, n44195);
  and g74106 (n44196, n_29812, n_33001);
  not g74107 (n_33002, n44194);
  and g74108 (n44197, pi0230, n_33002);
  not g74109 (n_33003, n44196);
  and g74110 (n44198, n_33003, n44197);
  not g74111 (n_33004, n40931);
  and g74112 (n44199, n_33004, n44154);
  not g74113 (n_33005, n44199);
  and g74114 (n44200, n44160, n_33005);
  and g74115 (n44201, n13062, n42455);
  not g74116 (n_33006, n44201);
  and g74117 (n44202, n_32982, n_33006);
  not g74118 (n_33007, n44200);
  and g74119 (n44203, n_33007, n44202);
  not g74120 (n_33008, n44203);
  and g74121 (n44204, n_4226, n_33008);
  and g74122 (n44205, n_32782, n44174);
  not g74123 (n_33009, n44204);
  and g74124 (n44206, n_33009, n44205);
  not g74125 (n_33010, n44198);
  not g74126 (n_33011, n44206);
  and g74127 (n44207, n_33010, n_33011);
  not g74128 (n_33012, n44207);
  and g74129 (n44208, pi1134, n_33012);
  not g74130 (n_33013, n44189);
  not g74131 (n_33014, n44208);
  and g74132 (po0435, n_33013, n_33014);
  and g74133 (n44210, n_2611, n_32156);
  not g74134 (n_33016, pi0958);
  and g74135 (n44211, n_33016, n40863);
  not g74136 (n_33017, n44210);
  and g74137 (n44212, n_3128, n_33017);
  not g74138 (n_33018, n44211);
  and g74139 (n44213, n_33018, n44212);
  and g74140 (n44214, pi1135, n43688);
  not g74141 (n_33019, n44213);
  not g74142 (n_33020, n44214);
  and g74143 (n44215, n_33019, n_33020);
  not g74144 (n_33021, n44215);
  and g74145 (n44216, pi0199, n_33021);
  and g74146 (n44217, pi0958, n40885);
  and g74147 (n44218, pi0279, n_32161);
  not g74148 (n_33022, n44217);
  and g74149 (n44219, n_3128, n_33022);
  not g74150 (n_33023, n44218);
  and g74151 (n44220, n_33023, n44219);
  and g74152 (n44221, n_32967, n43688);
  not g74153 (n_33024, n44221);
  and g74154 (n44222, n_7044, n_33024);
  not g74155 (n_33025, n44220);
  and g74156 (n44223, n_33025, n44222);
  not g74157 (n_33026, n44216);
  not g74158 (n_33027, n44223);
  and g74159 (n44224, n_33026, n_33027);
  not g74160 (n_33028, n44224);
  and g74161 (n44225, n16479, n_33028);
  not g74162 (n_33029, n40951);
  and g74163 (n44226, n_33029, n44225);
  and g74164 (n44227, n_31591, n_32968);
  and g74165 (n44228, n_33025, n44227);
  not g74166 (n_33030, n44228);
  and g74167 (n44229, n_6791, n_33030);
  and g74168 (n44230, pi1135, n42455);
  not g74169 (n_33031, n44230);
  and g74170 (n44231, pi0219, n_33031);
  and g74171 (n44232, n_33019, n44231);
  not g74172 (n_33032, n44232);
  and g74173 (n44233, n_25711, n_33032);
  not g74174 (n_33033, n44229);
  and g74175 (n44234, n_33033, n44233);
  not g74176 (n_33034, n44234);
  and g74177 (n44235, n_28510, n_33034);
  not g74178 (n_33035, n44226);
  and g74179 (n44236, n_33035, n44235);
  and g74180 (n44237, pi1135, n38519);
  and g74181 (n44238, n_7075, n_32967);
  not g74182 (n_33036, n44238);
  and g74183 (n44239, n_6791, n_33036);
  and g74184 (n44240, n_7075, n44239);
  not g74185 (n_33037, n44237);
  not g74186 (n_33038, n44240);
  and g74187 (n44241, n_33037, n_33038);
  not g74188 (n_33039, n44241);
  and g74189 (n44242, po1038, n_33039);
  and g74190 (n44243, pi0199, pi1135);
  not g74191 (n_33040, n44243);
  and g74192 (n44244, n_32987, n_33040);
  not g74193 (n_33041, n44244);
  and g74194 (n44245, n38568, n_33041);
  and g74195 (n44246, pi0299, n_33039);
  not g74196 (n_33042, n44245);
  not g74197 (n_33043, n44246);
  and g74198 (n44247, n_33042, n_33043);
  not g74199 (n_33044, n44247);
  and g74200 (n44248, n_4226, n_33044);
  not g74201 (n_33045, n44242);
  and g74202 (n44249, pi0230, n_33045);
  not g74203 (n_33046, n44248);
  and g74204 (n44250, n_33046, n44249);
  not g74205 (n_33047, n44236);
  not g74206 (n_33048, n44250);
  and g74207 (n44251, n_33047, n_33048);
  not g74208 (n_33049, n44251);
  and g74209 (n44252, n_2921, n_33049);
  and g74210 (n44253, n_32967, n10809);
  and g74211 (n44254, n_7045, pi1135);
  not g74212 (n_33050, n44254);
  and g74213 (n44255, pi0199, n_33050);
  not g74214 (n_33051, n44253);
  not g74215 (n_33052, n44255);
  and g74216 (n44256, n_33051, n_33052);
  not g74217 (n_33053, n44256);
  and g74218 (n44257, n16479, n_33053);
  not g74219 (n_33054, n44239);
  and g74220 (n44258, n_33037, n_33054);
  and g74221 (n44259, n_25711, n44258);
  not g74222 (n_33055, n44257);
  not g74223 (n_33056, n44259);
  and g74224 (n44260, n_33055, n_33056);
  not g74225 (n_33057, n44260);
  and g74226 (n44261, pi0230, n_33057);
  and g74227 (n44262, pi1091, n_33036);
  and g74228 (n44263, n40141, n44262);
  not g74229 (n_33058, n44225);
  not g74230 (n_33059, n44263);
  and g74231 (n44264, n_33058, n_33059);
  and g74232 (n44265, n44235, n44264);
  not g74233 (n_33060, n44261);
  not g74234 (n_33061, n44265);
  and g74235 (n44266, n_33060, n_33061);
  not g74236 (n_33062, n44266);
  and g74237 (n44267, pi1134, n_33062);
  not g74238 (n_33063, n44252);
  not g74239 (n_33064, n44267);
  and g74240 (po0436, n_33063, n_33064);
  and g74241 (n44269, n_7075, pi1135);
  and g74242 (n44270, pi0211, pi1136);
  not g74243 (n_33065, n44269);
  not g74244 (n_33066, n44270);
  and g74245 (n44271, n_33065, n_33066);
  and g74246 (n44272, pi1091, n44271);
  not g74247 (n_33067, pi0280);
  and g74248 (n44273, n_33067, n_32161);
  and g74249 (n44274, pi0914, n40885);
  not g74250 (n_33069, n44273);
  and g74251 (n44275, n_3128, n_33069);
  not g74252 (n_33070, n44274);
  and g74253 (n44276, n_33070, n44275);
  not g74254 (n_33071, n44272);
  not g74255 (n_33072, n44276);
  and g74256 (n44277, n_33071, n_33072);
  not g74257 (n_33073, n44277);
  and g74258 (n44278, n_6791, n_33073);
  and g74259 (n44279, n_7075, pi1137);
  not g74260 (n_33074, n44279);
  and g74261 (n44280, pi0219, n_33074);
  not g74262 (n_33075, n44280);
  and g74263 (n44281, n_32174, n_33075);
  not g74264 (n_33076, pi0914);
  and g74265 (n44282, n_33076, n40863);
  and g74266 (n44283, pi0280, n_32156);
  not g74267 (n_33077, n44282);
  and g74268 (n44284, n_3128, n_33077);
  not g74269 (n_33078, n44283);
  and g74270 (n44285, n_33078, n44284);
  not g74271 (n_33079, n44281);
  not g74272 (n_33080, n44285);
  and g74273 (n44286, n_33079, n_33080);
  not g74274 (n_33081, n44278);
  not g74275 (n_33082, n44286);
  and g74276 (n44287, n_33081, n_33082);
  not g74277 (n_33083, n44287);
  and g74278 (n44288, n_25711, n_33083);
  and g74279 (n44289, pi1137, n43688);
  not g74280 (n_33084, n44289);
  and g74281 (n44290, n_33080, n_33084);
  not g74282 (n_33085, n44290);
  and g74283 (n44291, pi0199, n_33085);
  and g74284 (n44292, pi0200, pi1136);
  and g74285 (n44293, pi1091, n_33050);
  not g74286 (n_33086, n44292);
  and g74287 (n44294, n_33086, n44293);
  not g74288 (n_33087, n44294);
  and g74289 (n44295, n_7044, n_33087);
  and g74290 (n44296, n_33072, n44295);
  not g74291 (n_33088, n44291);
  and g74292 (n44297, n16479, n_33088);
  not g74293 (n_33089, n44296);
  and g74294 (n44298, n_33089, n44297);
  not g74295 (n_33090, n44288);
  not g74296 (n_33091, n44298);
  and g74297 (n44299, n_33090, n_33091);
  not g74298 (n_33092, n44299);
  and g74299 (n44300, n_28510, n_33092);
  and g74300 (n44301, pi0200, n_32560);
  and g74301 (n44302, pi0199, pi1137);
  and g74302 (n44303, n_7045, n_32225);
  not g74303 (n_33093, n44302);
  and g74304 (n44304, n_33093, n44303);
  not g74305 (n_33094, n44301);
  not g74306 (n_33095, n44304);
  and g74307 (n44305, n_33094, n_33095);
  and g74308 (n44306, n16479, n44305);
  and g74309 (n44307, n_6791, n44271);
  not g74310 (n_33096, n44307);
  and g74311 (n44308, n_33075, n_33096);
  and g74312 (n44309, n_25711, n44308);
  not g74313 (n_33097, n44306);
  and g74314 (n44310, pi0230, n_33097);
  not g74315 (n_33098, n44309);
  and g74316 (n44311, n_33098, n44310);
  not g74317 (n_33099, n44300);
  not g74318 (n_33100, n44311);
  and g74319 (po0437, n_33099, n_33100);
  and g74320 (n44313, n_7044, pi1138);
  not g74321 (n_33101, n44313);
  and g74322 (n44314, pi0200, n_33101);
  and g74323 (n44315, pi0199, pi1139);
  and g74324 (n44316, n_7045, n_32558);
  not g74325 (n_33102, n44315);
  and g74326 (n44317, n_33102, n44316);
  not g74327 (n_33103, n44314);
  not g74328 (n_33104, n44317);
  and g74329 (n44318, n_33103, n_33104);
  not g74330 (n_33105, n44318);
  and g74331 (n44319, n16479, n_33105);
  and g74332 (n44320, pi0219, n43712);
  and g74333 (n44321, pi0211, pi1138);
  not g74334 (n_33106, n44321);
  and g74335 (n44322, n_33074, n_33106);
  not g74336 (n_33107, n44322);
  and g74337 (n44323, n_6791, n_33107);
  not g74338 (n_33108, n44320);
  not g74339 (n_33109, n44323);
  and g74340 (n44324, n_33108, n_33109);
  and g74341 (n44325, n_25711, n44324);
  not g74342 (n_33110, n44319);
  not g74343 (n_33111, n44325);
  and g74344 (n44326, n_33110, n_33111);
  not g74345 (n_33112, n44326);
  and g74346 (n44327, pi0230, n_33112);
  not g74347 (n_33114, pi0830);
  and g74348 (n44328, n_33114, n40885);
  and g74349 (n44329, pi0281, n_32161);
  not g74350 (n_33115, n44328);
  and g74351 (n44330, n_3128, n_33115);
  not g74352 (n_33116, n44329);
  and g74353 (n44331, n_33116, n44330);
  and g74354 (n44332, pi1091, n_33107);
  not g74355 (n_33117, n44332);
  and g74356 (n44333, n40141, n_33117);
  and g74357 (n44334, pi1138, n40951);
  not g74358 (n_33118, n44334);
  and g74359 (n44335, n_33084, n_33118);
  and g74360 (n44336, n43500, n44335);
  not g74361 (n_33119, n44333);
  not g74362 (n_33120, n44336);
  and g74363 (n44337, n_33119, n_33120);
  not g74364 (n_33121, n44331);
  not g74365 (n_33122, n44337);
  and g74366 (n44338, n_33121, n_33122);
  and g74367 (n44339, n_33114, n40863);
  and g74368 (n44340, pi0281, n_32156);
  not g74369 (n_33123, n44339);
  and g74370 (n44341, n_3128, n_33123);
  not g74371 (n_33124, n44340);
  and g74372 (n44342, n_33124, n44341);
  and g74373 (n44343, pi1139, n42455);
  not g74374 (n_33125, n44343);
  and g74375 (n44344, n43686, n_33125);
  and g74376 (n44345, pi0199, n_32612);
  and g74377 (n44346, n16479, n44345);
  not g74378 (n_33126, n44344);
  not g74379 (n_33127, n44346);
  and g74380 (n44347, n_33126, n_33127);
  not g74381 (n_33128, n44342);
  not g74382 (n_33129, n44347);
  and g74383 (n44348, n_33128, n_33129);
  not g74384 (n_33130, n44338);
  not g74385 (n_33131, n44348);
  and g74386 (n44349, n_33130, n_33131);
  not g74387 (n_33132, n44349);
  and g74388 (n44350, n_28510, n_33132);
  not g74389 (n_33133, n44327);
  not g74390 (n_33134, n44350);
  and g74391 (po0438, n_33133, n_33134);
  and g74392 (n44352, pi0200, n_32624);
  and g74393 (n44353, pi0199, pi1140);
  and g74394 (n44354, n_7045, n_33101);
  not g74395 (n_33135, n44353);
  and g74396 (n44355, n_33135, n44354);
  not g74397 (n_33136, n44352);
  not g74398 (n_33137, n44355);
  and g74399 (n44356, n_33136, n_33137);
  not g74400 (n_33138, n44356);
  and g74401 (n44357, n16479, n_33138);
  and g74402 (n44358, pi0219, n44129);
  and g74403 (n44359, pi0211, pi1139);
  not g74404 (n_33139, n43660);
  not g74405 (n_33140, n44359);
  and g74406 (n44360, n_33139, n_33140);
  not g74407 (n_33141, n44360);
  and g74408 (n44361, n_6791, n_33141);
  not g74409 (n_33142, n44358);
  not g74410 (n_33143, n44361);
  and g74411 (n44362, n_33142, n_33143);
  and g74412 (n44363, n_25711, n44362);
  not g74413 (n_33144, n44357);
  not g74414 (n_33145, n44363);
  and g74415 (n44364, n_33144, n_33145);
  not g74416 (n_33146, n44364);
  and g74417 (n44365, pi0230, n_33146);
  not g74418 (n_33148, pi0836);
  and g74419 (n44366, n_33148, n40885);
  and g74420 (n44367, pi0282, n_32161);
  not g74421 (n_33149, n44366);
  and g74422 (n44368, n_3128, n_33149);
  not g74423 (n_33150, n44367);
  and g74424 (n44369, n_33150, n44368);
  and g74425 (n44370, pi1091, n_33141);
  not g74426 (n_33151, n44370);
  and g74427 (n44371, n40141, n_33151);
  and g74428 (n44372, pi1139, n40951);
  not g74429 (n_33152, n44372);
  and g74430 (n44373, n_32585, n_33152);
  and g74431 (n44374, n43500, n44373);
  not g74432 (n_33153, n44371);
  not g74433 (n_33154, n44374);
  and g74434 (n44375, n_33153, n_33154);
  not g74435 (n_33155, n44369);
  not g74436 (n_33156, n44375);
  and g74437 (n44376, n_33155, n_33156);
  and g74438 (n44377, n_33148, n40863);
  and g74439 (n44378, pi0282, n_32156);
  not g74440 (n_33157, n44377);
  and g74441 (n44379, n_3128, n_33157);
  not g74442 (n_33158, n44378);
  and g74443 (n44380, n_33158, n44379);
  and g74444 (n44381, pi1140, n42455);
  not g74445 (n_33159, n44381);
  and g74446 (n44382, n43686, n_33159);
  and g74447 (n44383, n_7045, n43717);
  not g74448 (n_33160, n44383);
  and g74449 (n44384, pi0199, n_33160);
  and g74450 (n44385, n16479, n44384);
  not g74451 (n_33161, n44382);
  not g74452 (n_33162, n44385);
  and g74453 (n44386, n_33161, n_33162);
  not g74454 (n_33163, n44380);
  not g74455 (n_33164, n44386);
  and g74456 (n44387, n_33163, n_33164);
  not g74457 (n_33165, n44376);
  not g74458 (n_33166, n44387);
  and g74459 (n44388, n_33165, n_33166);
  not g74460 (n_33167, n44388);
  and g74461 (n44389, n_28510, n_33167);
  not g74462 (n_33168, n44365);
  not g74463 (n_33169, n44389);
  and g74464 (po0439, n_33168, n_33169);
  and g74465 (n44391, pi1147, n_32791);
  and g74466 (n44392, pi1149, n_31565);
  not g74467 (n_33170, n44391);
  not g74468 (n_33171, n44392);
  and g74469 (n44393, n_33170, n_33171);
  not g74470 (n_33172, n44393);
  and g74471 (n44394, n_29904, n_33172);
  and g74472 (n44395, n43884, n_33170);
  not g74473 (n_33173, n43501);
  and g74474 (n44396, pi1147, n_33173);
  and g74475 (n44397, n_29850, n43510);
  not g74476 (n_33174, n44396);
  and g74477 (n44398, n_33174, n44397);
  not g74478 (n_33175, n44395);
  and g74479 (n44399, pi1148, n_33175);
  not g74480 (n_33176, n44398);
  and g74481 (n44400, n_33176, n44399);
  not g74482 (n_33177, n44394);
  and g74483 (n44401, pi0230, n_33177);
  not g74484 (n_33178, n44400);
  and g74485 (n44402, n_33178, n44401);
  and g74486 (n44403, n_29810, n43637);
  and g74487 (n44404, pi1147, n43541);
  not g74488 (n_33179, n44404);
  and g74489 (n44405, pi1148, n_33179);
  not g74490 (n_33180, n44403);
  and g74491 (n44406, n_33180, n44405);
  and g74492 (n44407, pi1147, n43535);
  and g74493 (n44408, n_29810, n_32540);
  not g74494 (n_33181, n44408);
  and g74495 (n44409, n_29904, n_33181);
  not g74496 (n_33182, n44407);
  and g74497 (n44410, n_33182, n44409);
  not g74498 (n_33183, n44406);
  and g74499 (n44411, n_29850, n_33183);
  not g74500 (n_33184, n44410);
  and g74501 (n44412, n_33184, n44411);
  and g74502 (n44413, n_29810, n43629);
  and g74503 (n44414, pi1147, n43580);
  not g74504 (n_33185, n44414);
  and g74505 (n44415, pi1148, n_33185);
  not g74506 (n_33186, n44413);
  and g74507 (n44416, n_33186, n44415);
  and g74508 (n44417, n_29810, n43623);
  and g74509 (n44418, pi1147, n43575);
  not g74510 (n_33187, n44417);
  and g74511 (n44419, n_29904, n_33187);
  not g74512 (n_33188, n44418);
  and g74513 (n44420, n_33188, n44419);
  not g74514 (n_33189, n44416);
  and g74515 (n44421, pi1149, n_33189);
  not g74516 (n_33190, n44420);
  and g74517 (n44422, n_33190, n44421);
  not g74518 (n_33191, n44412);
  and g74519 (n44423, pi0283, n_33191);
  not g74520 (n_33192, n44422);
  and g74521 (n44424, n_33192, n44423);
  and g74522 (n44425, n_29810, n43605);
  and g74523 (n44426, pi1147, n43586);
  not g74524 (n_33193, n44425);
  and g74525 (n44427, pi1149, n_33193);
  not g74526 (n_33194, n44426);
  and g74527 (n44428, n_33194, n44427);
  and g74528 (n44429, n_29810, n_32479);
  and g74529 (n44430, pi1147, n43555);
  not g74530 (n_33195, n44429);
  and g74531 (n44431, n_29850, n_33195);
  not g74532 (n_33196, n44430);
  and g74533 (n44432, n_33196, n44431);
  not g74534 (n_33197, n44432);
  and g74535 (n44433, n_29904, n_33197);
  not g74536 (n_33198, n44428);
  and g74537 (n44434, n_33198, n44433);
  and g74538 (n44435, n_29810, n43608);
  and g74539 (n44436, pi1147, n43593);
  not g74540 (n_33199, n44436);
  and g74541 (n44437, pi1149, n_33199);
  not g74542 (n_33200, n44435);
  and g74543 (n44438, n_33200, n44437);
  and g74544 (n44439, pi1147, n43563);
  and g74545 (n44440, n_29810, n_32723);
  not g74546 (n_33201, n44439);
  and g74547 (n44441, n_29850, n_33201);
  not g74548 (n_33202, n44440);
  and g74549 (n44442, n_33202, n44441);
  not g74550 (n_33203, n44438);
  and g74551 (n44443, pi1148, n_33203);
  not g74552 (n_33204, n44442);
  and g74553 (n44444, n_33204, n44443);
  not g74554 (n_33205, n44434);
  and g74555 (n44445, n_32691, n_33205);
  not g74556 (n_33206, n44444);
  and g74557 (n44446, n_33206, n44445);
  not g74558 (n_33207, n44424);
  and g74559 (n44447, n_28510, n_33207);
  not g74560 (n_33208, n44446);
  and g74561 (n44448, n_33208, n44447);
  not g74562 (n_33209, n44402);
  not g74563 (n_33210, n44448);
  and g74564 (po0440, n_33209, n_33210);
  and g74565 (n44450, n_1170, n_31974);
  and g74566 (n44451, pi1143, n42902);
  and g74567 (n44452, n_30219, n44451);
  or g74568 (po0441, n44450, n44452);
  and g74569 (n44454, n2572, n_6724);
  and g74570 (n44455, n_8134, n44454);
  and g74571 (n44456, pi0286, n44455);
  and g74572 (n44457, pi0288, pi0289);
  and g74573 (n44458, n44456, n44457);
  and g74574 (n44459, pi0285, n44458);
  and g74575 (n44460, pi0285, n44454);
  not g74576 (n_33211, n44458);
  not g74577 (n_33212, n44460);
  and g74578 (n44461, n_33211, n_33212);
  not g74579 (n_33213, n44459);
  and g74580 (n44462, n_4226, n_33213);
  not g74581 (n_33214, n44461);
  and g74582 (n44463, n_33214, n44462);
  and g74583 (n44464, n_4226, n44458);
  and g74584 (n44465, n_4086, n7420);
  and g74585 (n44466, n_4090, n44465);
  and g74586 (n44467, n_4088, n44466);
  not g74587 (n_33215, n44467);
  and g74588 (n44468, pi0285, n_33215);
  not g74589 (n_33216, n44464);
  and g74590 (n44469, n_33216, n44468);
  not g74591 (n_33217, n44463);
  not g74592 (n_33218, n44469);
  and g74593 (n44470, n_33217, n_33218);
  not g74594 (n_33220, pi0793);
  not g74595 (n_33221, n44470);
  and g74596 (po0442, n_33220, n_33221);
  not g74597 (n_33222, n7424);
  and g74598 (n44472, n_4090, n_33222);
  and g74599 (n44473, n7420, n44472);
  not g74600 (n_33223, n44473);
  and g74601 (n44474, pi0286, n_33223);
  and g74602 (n44475, n_4086, n44473);
  not g74603 (n_33224, n44474);
  and g74604 (n44476, po1038, n_33224);
  not g74605 (n_33225, n44475);
  and g74606 (n44477, n_33225, n44476);
  not g74607 (n_33226, n44454);
  and g74608 (n44478, n7420, n_33226);
  not g74609 (n_33227, n44478);
  and g74610 (n44479, pi0286, n_33227);
  and g74611 (n44480, n_33226, n44465);
  not g74612 (n_33228, n44479);
  not g74613 (n_33229, n44480);
  and g74614 (n44481, n_33228, n_33229);
  not g74615 (n_33230, n44481);
  and g74616 (n44482, n44472, n_33230);
  not g74617 (n_33231, n44455);
  and g74618 (n44483, n_4086, n_33231);
  not g74619 (n_33232, n44456);
  and g74620 (n44484, pi0288, n_33232);
  not g74621 (n_33233, n44483);
  and g74622 (n44485, n_33233, n44484);
  not g74623 (n_33234, n44482);
  and g74624 (n44486, n_4226, n_33234);
  not g74625 (n_33235, n44485);
  and g74626 (n44487, n_33235, n44486);
  not g74627 (n_33236, n44477);
  and g74628 (n44488, n_33220, n_33236);
  not g74629 (n_33237, n44487);
  and g74630 (po0443, n_33237, n44488);
  and g74631 (n44490, n_3084, pi0457);
  not g74632 (n_33239, n44490);
  and g74633 (po0444, n_4, n_33239);
  and g74634 (n44492, pi0288, n_8134);
  not g74635 (n_33240, n44492);
  and g74636 (n44493, n_33223, n_33240);
  and g74637 (po0637, n_4226, n44454);
  not g74638 (n_33241, n44493);
  and g74639 (n44495, n_33241, po0637);
  not g74640 (n_33243, po0637);
  and g74641 (n44496, n44493, n_33243);
  not g74642 (n_33244, n44495);
  and g74643 (n44497, n_33220, n_33244);
  not g74644 (n_33245, n44496);
  and g74645 (po0445, n_33245, n44497);
  not g74646 (n_33246, n44466);
  and g74647 (n44499, pi0289, n_33246);
  and g74648 (n44500, pi0285, n_4088);
  and g74649 (n44501, n44466, n44500);
  not g74650 (n_33247, n44499);
  and g74651 (n44502, po1038, n_33247);
  not g74652 (n_33248, n44501);
  and g74653 (n44503, n_33248, n44502);
  and g74654 (n44504, n_4088, n44484);
  and g74655 (n44505, n44480, n44500);
  and g74656 (n44506, pi0289, n_33229);
  not g74657 (n_33249, n44505);
  and g74658 (n44507, n_4090, n_33249);
  not g74659 (n_33250, n44506);
  and g74660 (n44508, n_33250, n44507);
  not g74661 (n_33251, n44504);
  and g74662 (n44509, n_33211, n_33251);
  not g74663 (n_33252, n44508);
  and g74664 (n44510, n_33252, n44509);
  not g74665 (n_33253, n44510);
  and g74666 (n44511, n_4226, n_33253);
  not g74667 (n_33254, n44503);
  and g74668 (n44512, n_33220, n_33254);
  not g74669 (n_33255, n44511);
  and g74670 (po0446, n_33255, n44512);
  not g74671 (n_33257, pi0290);
  and g74672 (n44514, n_33257, pi0476);
  not g74673 (n_33258, pi1048);
  and g74674 (n44515, n_31526, n_33258);
  not g74675 (n_33259, n44514);
  not g74676 (n_33260, n44515);
  and g74677 (po0447, n_33259, n_33260);
  not g74678 (n_33262, pi0291);
  and g74679 (n44517, n_33262, pi0476);
  not g74680 (n_33263, pi1049);
  and g74681 (n44518, n_31526, n_33263);
  not g74682 (n_33264, n44517);
  not g74683 (n_33265, n44518);
  and g74684 (po0448, n_33264, n_33265);
  not g74685 (n_33267, pi0292);
  and g74686 (n44520, n_33267, pi0476);
  not g74687 (n_33268, pi1084);
  and g74688 (n44521, n_31526, n_33268);
  not g74689 (n_33269, n44520);
  not g74690 (n_33270, n44521);
  and g74691 (po0449, n_33269, n_33270);
  not g74692 (n_33272, pi0293);
  and g74693 (n44523, n_33272, pi0476);
  not g74694 (n_33273, pi1059);
  and g74695 (n44524, n_31526, n_33273);
  not g74696 (n_33274, n44523);
  not g74697 (n_33275, n44524);
  and g74698 (po0450, n_33274, n_33275);
  not g74699 (n_33277, pi0294);
  and g74700 (n44526, n_33277, pi0476);
  not g74701 (n_33278, pi1072);
  and g74702 (n44527, n_31526, n_33278);
  not g74703 (n_33279, n44526);
  not g74704 (n_33280, n44527);
  and g74705 (po0451, n_33279, n_33280);
  not g74706 (n_33282, pi0295);
  and g74707 (n44529, n_33282, pi0476);
  not g74708 (n_33283, pi1053);
  and g74709 (n44530, n_31526, n_33283);
  not g74710 (n_33284, n44529);
  not g74711 (n_33285, n44530);
  and g74712 (po0452, n_33284, n_33285);
  not g74713 (n_33287, pi0296);
  and g74714 (n44532, n_33287, pi0476);
  not g74715 (n_33288, pi1037);
  and g74716 (n44533, n_31526, n_33288);
  not g74717 (n_33289, n44532);
  not g74718 (n_33290, n44533);
  and g74719 (po0453, n_33289, n_33290);
  not g74720 (n_33292, pi0297);
  and g74721 (n44535, n_33292, pi0476);
  not g74722 (n_33293, pi1044);
  and g74723 (n44536, n_31526, n_33293);
  not g74724 (n_33294, n44535);
  not g74725 (n_33295, n44536);
  and g74726 (po0454, n_33294, n_33295);
  not g74727 (n_33297, pi0478);
  and g74728 (n44538, n_33297, pi1044);
  and g74729 (n44539, pi0298, pi0478);
  or g74730 (po0455, n44538, n44539);
  and g74731 (n44541, pi0054, n2521);
  and g74732 (n44542, n_167, n13153);
  and g74733 (n44543, n13411, n44542);
  not g74734 (n_33299, n44541);
  not g74735 (n_33300, n44543);
  and g74736 (n44544, n_33299, n_33300);
  and g74737 (n44545, n2621, n8880);
  not g74738 (n_33301, n44544);
  and g74739 (n44546, n_33301, n44545);
  not g74740 (n_33302, n44546);
  and g74741 (n44547, n_162, n_33302);
  not g74742 (n_33303, n44547);
  and g74743 (po0456, n_7337, n_33303);
  and g74744 (n44549, pi0057, n_792);
  and g74745 (n44550, n10068, n44549);
  not g74746 (n_33305, pi0312);
  and g74747 (n44551, n_33305, n44550);
  not g74748 (n_33307, n44551);
  and g74749 (n44552, pi0300, n_33307);
  not g74750 (n_33308, pi0300);
  and g74751 (n44553, n_33308, n44551);
  not g74752 (n_33309, n44553);
  and g74753 (n44554, n_176, n_33309);
  not g74754 (n_33310, n44554);
  or g74755 (po0457, n44552, n_33310);
  not g74756 (n_33312, pi0301);
  and g74757 (n44556, n_33312, n44554);
  and g74758 (n44557, n_176, pi0301);
  and g74759 (n44558, n44553, n44557);
  or g74760 (po0458, n44556, n44558);
  and g74761 (n44560, n5836, n_4226);
  and g74762 (n44561, n_226, n_223);
  not g74763 (n_33314, n44561);
  and g74764 (n44562, pi0937, n_33314);
  and g74765 (n44563, pi0273, n3351);
  not g74766 (n_33315, n44562);
  not g74767 (n_33316, n44563);
  and g74768 (n44564, n_33315, n_33316);
  and g74769 (n44565, n44560, n44564);
  and g74770 (n44566, n_9349, n44565);
  and g74771 (n44567, n3449, n_25711);
  not g74772 (n_33317, n44565);
  not g74773 (n_33318, n44567);
  and g74774 (n44568, n_33317, n_33318);
  not g74775 (n_33319, n44568);
  and g74776 (n44569, pi0237, n_33319);
  and g74777 (n44570, n5780, n_25711);
  not g74778 (n_33320, n44560);
  not g74779 (n_33321, n44570);
  and g74780 (n44571, n_33320, n_33321);
  and g74781 (n44572, n_29904, n44571);
  and g74782 (n44573, n_36, n3310);
  and g74783 (n44574, n_32754, n44573);
  and g74784 (n44575, pi0833, n7570);
  not g74785 (n_33322, pi0937);
  and g74786 (n44576, n_33322, n44575);
  not g74787 (n_33323, n44574);
  not g74788 (n_33324, n44576);
  and g74789 (n44577, n_33323, n_33324);
  not g74790 (n_33325, n44577);
  and g74791 (n44578, n_25711, n_33325);
  and g74799 (n44582, n_33297, pi1049);
  and g74800 (n44583, pi0303, pi0478);
  or g74801 (po0460, n44582, n44583);
  and g74802 (n44585, n_33297, pi1048);
  and g74803 (n44586, pi0304, pi0478);
  or g74804 (po0461, n44585, n44586);
  and g74805 (n44588, n_33297, pi1084);
  and g74806 (n44589, pi0305, pi0478);
  or g74807 (po0462, n44588, n44589);
  and g74808 (n44591, n_33297, pi1059);
  and g74809 (n44592, pi0306, pi0478);
  or g74810 (po0463, n44591, n44592);
  and g74811 (n44594, n_33297, pi1053);
  and g74812 (n44595, pi0307, pi0478);
  or g74813 (po0464, n44594, n44595);
  and g74814 (n44597, n_33297, pi1037);
  and g74815 (n44598, pi0308, pi0478);
  or g74816 (po0465, n44597, n44598);
  and g74817 (n44600, n_33297, pi1072);
  and g74818 (n44601, pi0309, pi0478);
  or g74819 (po0466, n44600, n44601);
  and g74820 (n44603, pi1147, n44571);
  not g74821 (n_33338, pi0934);
  and g74822 (n44604, pi0222, n_33338);
  and g74823 (n44605, n_32630, n3351);
  not g74824 (n_33339, n44604);
  not g74825 (n_33340, n44605);
  and g74826 (n44606, n_33339, n_33340);
  and g74827 (n44607, n44560, n44606);
  and g74828 (n44608, n_9350, n44570);
  not g74829 (n_33341, n2526);
  and g74830 (n44609, pi0934, n_33341);
  and g74831 (n44610, pi0271, n3310);
  not g74832 (n_33342, n44609);
  not g74833 (n_33343, n44610);
  and g74834 (n44611, n_33342, n_33343);
  not g74835 (n_33344, n44611);
  and g74836 (n44612, n44608, n_33344);
  not g74837 (n_33345, n44607);
  and g74838 (n44613, n_33318, n_33345);
  not g74839 (n_33346, n44612);
  and g74840 (n44614, n_33346, n44613);
  not g74841 (n_33347, n44603);
  and g74842 (n44615, n_33347, n44614);
  not g74843 (n_33348, n44615);
  and g74844 (n44616, n_25720, n_33348);
  and g74845 (n44617, n2604, n16479);
  not g74846 (n_33349, n44606);
  and g74847 (n44618, n44560, n_33349);
  and g74848 (n44619, n44570, n44611);
  not g74849 (n_33350, n44617);
  and g74855 (n44623, n_9349, n44560);
  not g74856 (n_33353, n44608);
  not g74857 (n_33354, n44623);
  and g74858 (n44624, n_33353, n_33354);
  not g74859 (n_33355, n44624);
  and g74860 (n44625, n_29810, n_33355);
  not g74861 (n_33356, n44614);
  and g74862 (n44626, n_33356, n44625);
  not g74863 (n_33357, n44622);
  not g74864 (n_33358, n44626);
  and g74865 (n44627, n_33357, n_33358);
  not g74866 (n_33359, n44627);
  and g74867 (n44628, pi0233, n_33359);
  or g74868 (po0467, n44616, n44628);
  not g74869 (n_33361, pi0311);
  and g74870 (n44630, n_176, n_33361);
  not g74871 (n_33362, n44558);
  not g74872 (n_33363, n44630);
  and g74873 (n44631, n_33362, n_33363);
  and g74874 (n44632, n_33361, n44558);
  not g74875 (n_33364, n44631);
  not g74876 (n_33365, n44632);
  and g74877 (po0468, n_33364, n_33365);
  not g74878 (n_33366, n44550);
  and g74879 (n44634, pi0312, n_33366);
  not g74880 (n_33367, n44634);
  and g74881 (n44635, n_33307, n_33367);
  not g74882 (n_33368, n44635);
  and g74883 (po0469, n_176, n_33368);
  not g74884 (n_33369, n10388);
  not g74885 (n_33370, n13446);
  and g74886 (n44637, n_33369, n_33370);
  not g74887 (n_33371, n13453);
  and g74888 (n44638, po0740, n_33371);
  not g74889 (n_33372, n44638);
  and g74890 (n44639, n10166, n_33372);
  not g74891 (n_33373, n44639);
  or g74892 (po0634, n44637, n_33373);
  and g74893 (n44641, po1110, po0634);
  and g74894 (n44642, pi0313, pi0954);
  not g74895 (n_33376, n44641);
  not g74896 (n_33377, n44642);
  and g74897 (po0470, n_33376, n_33377);
  and g74898 (n44644, n6323, n8880);
  not g74899 (n_33378, n44644);
  and g74900 (n44645, n14440, n_33378);
  and g74901 (n44646, pi0039, n_10353);
  and g74902 (n44647, n_162, n_9763);
  not g74903 (n_33379, n44646);
  and g74904 (n44648, n2608, n_33379);
  not g74905 (n_33380, n44647);
  and g74906 (n44649, n_33380, n44648);
  not g74907 (n_33381, n44649);
  and g74908 (n44650, n_10963, n_33381);
  and g74909 (n44651, n2534, n10163);
  not g74910 (n_33382, n44650);
  and g74911 (n44652, n_33382, n44651);
  not g74912 (n_33383, n44645);
  not g74913 (n_33384, n44652);
  and g74914 (n44653, n_33383, n_33384);
  and g74915 (n44654, n14432, n14433);
  not g74916 (n_33385, n44653);
  and g74917 (po0471, n_33385, n44654);
  not g74918 (n_33387, pi0340);
  and g74919 (n44656, n_33387, n44454);
  and g74920 (n44657, n_4226, n44656);
  not g74921 (n_33388, n44657);
  and g74922 (n44658, pi0315, n_33388);
  and g74923 (n44659, pi1080, n44657);
  or g74924 (po0472, n44658, n44659);
  and g74925 (n44661, pi0316, n_33388);
  and g74926 (n44662, pi1047, n44657);
  or g74927 (po0473, n44661, n44662);
  not g74928 (n_33392, pi0330);
  and g74929 (n44664, n_33392, po0637);
  not g74930 (n_33393, n44664);
  and g74931 (n44665, pi0317, n_33393);
  and g74932 (n44666, pi1078, n44664);
  or g74933 (po0474, n44665, n44666);
  not g74934 (n_33396, pi0341);
  and g74935 (n44668, n_33396, n44454);
  and g74936 (n44669, n_4226, n44668);
  not g74937 (n_33397, n44669);
  and g74938 (n44670, pi0318, n_33397);
  and g74939 (n44671, pi1074, n44669);
  or g74940 (po0475, n44670, n44671);
  and g74941 (n44673, pi0319, n_33397);
  and g74942 (n44674, pi1072, n44669);
  or g74943 (po0476, n44673, n44674);
  and g74944 (n44676, pi0320, n_33388);
  and g74945 (n44677, pi1048, n44657);
  or g74946 (po0477, n44676, n44677);
  and g74947 (n44679, pi0321, n_33388);
  and g74948 (n44680, pi1058, n44657);
  or g74949 (po0478, n44679, n44680);
  and g74950 (n44682, pi0322, n_33388);
  and g74951 (n44683, pi1051, n44657);
  or g74952 (po0479, n44682, n44683);
  and g74953 (n44685, pi0323, n_33388);
  and g74954 (n44686, pi1065, n44657);
  or g74955 (po0480, n44685, n44686);
  and g74956 (n44688, pi0324, n_33397);
  and g74957 (n44689, pi1086, n44669);
  or g74958 (po0481, n44688, n44689);
  and g74959 (n44691, pi0325, n_33397);
  and g74960 (n44692, pi1063, n44669);
  or g74961 (po0482, n44691, n44692);
  and g74962 (n44694, pi0326, n_33397);
  and g74963 (n44695, pi1057, n44669);
  or g74964 (po0483, n44694, n44695);
  and g74965 (n44697, pi0327, n_33388);
  and g74966 (n44698, pi1040, n44657);
  or g74967 (po0484, n44697, n44698);
  and g74968 (n44700, pi0328, n_33397);
  and g74969 (n44701, pi1058, n44669);
  or g74970 (po0485, n44700, n44701);
  and g74971 (n44703, pi0329, n_33397);
  and g74972 (n44704, pi1043, n44669);
  or g74973 (po0486, n44703, n44704);
  and g74974 (n44706, pi1092, n_28380);
  and g74975 (n44707, po1038, n44706);
  and g74976 (n44708, n_33392, n44707);
  and g74977 (n44709, n_4226, n44706);
  and g74978 (n44710, n_33392, n_33226);
  not g74979 (n_33405, n44656);
  not g74980 (n_33406, n44710);
  and g74981 (n44711, n_33405, n_33406);
  not g74982 (n_33407, n44711);
  and g74983 (n44712, n44709, n_33407);
  or g74984 (po0487, n44708, n44712);
  not g74985 (n_33409, pi0331);
  and g74986 (n44714, n_33409, n44707);
  and g74987 (n44715, n_33409, n_33226);
  not g74988 (n_33410, n44668);
  not g74989 (n_33411, n44715);
  and g74990 (n44716, n_33410, n_33411);
  not g74991 (n_33412, n44716);
  and g74992 (n44717, n44709, n_33412);
  or g74993 (po0488, n44714, n44717);
  and g74994 (n44719, n11002, n13166);
  not g74995 (n_33413, n11002);
  not g74996 (n_33414, n13102);
  and g74997 (n44720, n_33413, n_33414);
  not g74998 (n_33415, n44720);
  and g74999 (n44721, n7445, n_33415);
  not g75000 (n_33416, n44721);
  and g75001 (n44722, n_139, n_33416);
  and g75002 (n44723, pi0332, n9117);
  not g75003 (n_33417, n44722);
  and g75004 (n44724, n_33417, n44723);
  not g75005 (n_33418, n44719);
  not g75006 (n_33419, n44724);
  and g75007 (n44725, n_33418, n_33419);
  not g75008 (n_33420, n44725);
  and g75009 (n44726, n_162, n_33420);
  and g75010 (n44727, pi0039, n10368);
  not g75011 (n_33421, n44727);
  and g75012 (n44728, n_161, n_33421);
  not g75013 (n_33422, n44726);
  and g75014 (n44729, n_33422, n44728);
  not g75015 (n_33423, n44729);
  and g75016 (po0489, n38269, n_33423);
  and g75017 (n44731, pi0333, n_33397);
  and g75018 (n44732, pi1040, n44669);
  or g75019 (po0490, n44731, n44732);
  and g75020 (n44734, pi0334, n_33397);
  and g75021 (n44735, pi1065, n44669);
  or g75022 (po0491, n44734, n44735);
  and g75023 (n44737, pi0335, n_33397);
  and g75024 (n44738, pi1069, n44669);
  or g75025 (po0492, n44737, n44738);
  and g75026 (n44740, pi0336, n_33393);
  and g75027 (n44741, pi1070, n44664);
  or g75028 (po0493, n44740, n44741);
  and g75029 (n44743, pi0337, n_33393);
  and g75030 (n44744, pi1044, n44664);
  or g75031 (po0494, n44743, n44744);
  and g75032 (n44746, pi0338, n_33393);
  and g75033 (n44747, pi1072, n44664);
  or g75034 (po0495, n44746, n44747);
  and g75035 (n44749, pi0339, n_33393);
  and g75036 (n44750, pi1086, n44664);
  or g75037 (po0496, n44749, n44750);
  and g75038 (n44752, pi0340, n44707);
  and g75039 (n44753, n_33387, n_33226);
  and g75040 (n44754, n_33409, n44454);
  not g75041 (n_33424, n44753);
  and g75042 (n44755, n44709, n_33424);
  not g75043 (n_33425, n44754);
  and g75044 (n44756, n_33425, n44755);
  not g75045 (n_33426, n44752);
  not g75046 (n_33427, n44756);
  and g75047 (po0497, n_33426, n_33427);
  and g75048 (n44758, n_33396, n_33243);
  not g75049 (n_33428, n44758);
  and g75050 (n44759, n_33393, n_33428);
  not g75051 (n_33429, n44759);
  and g75052 (po0498, n44706, n_33429);
  and g75053 (n44761, pi0342, n_33388);
  and g75054 (n44762, pi1049, n44657);
  or g75055 (po0499, n44761, n44762);
  and g75056 (n44764, pi0343, n_33388);
  and g75057 (n44765, pi1062, n44657);
  or g75058 (po0500, n44764, n44765);
  and g75059 (n44767, pi0344, n_33388);
  and g75060 (n44768, pi1069, n44657);
  or g75061 (po0501, n44767, n44768);
  and g75062 (n44770, pi0345, n_33388);
  and g75063 (n44771, pi1039, n44657);
  or g75064 (po0502, n44770, n44771);
  and g75065 (n44773, pi0346, n_33388);
  and g75066 (n44774, pi1067, n44657);
  or g75067 (po0503, n44773, n44774);
  and g75068 (n44776, pi0347, n_33388);
  and g75069 (n44777, pi1055, n44657);
  or g75070 (po0504, n44776, n44777);
  and g75071 (n44779, pi0348, n_33388);
  and g75072 (n44780, pi1087, n44657);
  or g75073 (po0505, n44779, n44780);
  and g75074 (n44782, pi0349, n_33388);
  and g75075 (n44783, pi1043, n44657);
  or g75076 (po0506, n44782, n44783);
  and g75077 (n44785, pi0350, n_33388);
  and g75078 (n44786, pi1035, n44657);
  or g75079 (po0507, n44785, n44786);
  and g75080 (n44788, pi0351, n_33388);
  and g75081 (n44789, pi1079, n44657);
  or g75082 (po0508, n44788, n44789);
  and g75083 (n44791, pi0352, n_33388);
  and g75084 (n44792, pi1078, n44657);
  or g75085 (po0509, n44791, n44792);
  and g75086 (n44794, pi0353, n_33388);
  and g75087 (n44795, pi1063, n44657);
  or g75088 (po0510, n44794, n44795);
  and g75089 (n44797, pi0354, n_33388);
  and g75090 (n44798, pi1045, n44657);
  or g75091 (po0511, n44797, n44798);
  and g75092 (n44800, pi0355, n_33388);
  and g75093 (n44801, pi1084, n44657);
  or g75094 (po0512, n44800, n44801);
  and g75095 (n44803, pi0356, n_33388);
  and g75096 (n44804, pi1081, n44657);
  or g75097 (po0513, n44803, n44804);
  and g75098 (n44806, pi0357, n_33388);
  and g75099 (n44807, pi1076, n44657);
  or g75100 (po0514, n44806, n44807);
  and g75101 (n44809, pi0358, n_33388);
  and g75102 (n44810, pi1071, n44657);
  or g75103 (po0515, n44809, n44810);
  and g75104 (n44812, pi0359, n_33388);
  and g75105 (n44813, pi1068, n44657);
  or g75106 (po0516, n44812, n44813);
  and g75107 (n44815, pi0360, n_33388);
  and g75108 (n44816, pi1042, n44657);
  or g75109 (po0517, n44815, n44816);
  and g75110 (n44818, pi0361, n_33388);
  and g75111 (n44819, pi1059, n44657);
  or g75112 (po0518, n44818, n44819);
  and g75113 (n44821, pi0362, n_33388);
  and g75114 (n44822, pi1070, n44657);
  or g75115 (po0519, n44821, n44822);
  and g75116 (n44824, pi0363, n_33393);
  and g75117 (n44825, pi1049, n44664);
  or g75118 (po0520, n44824, n44825);
  and g75119 (n44827, pi0364, n_33393);
  and g75120 (n44828, pi1062, n44664);
  or g75121 (po0521, n44827, n44828);
  and g75122 (n44830, pi0365, n_33393);
  and g75123 (n44831, pi1065, n44664);
  or g75124 (po0522, n44830, n44831);
  and g75125 (n44833, pi0366, n_33393);
  and g75126 (n44834, pi1069, n44664);
  or g75127 (po0523, n44833, n44834);
  and g75128 (n44836, pi0367, n_33393);
  and g75129 (n44837, pi1039, n44664);
  or g75130 (po0524, n44836, n44837);
  and g75131 (n44839, pi0368, n_33393);
  and g75132 (n44840, pi1067, n44664);
  or g75133 (po0525, n44839, n44840);
  and g75134 (n44842, pi0369, n_33393);
  and g75135 (n44843, pi1080, n44664);
  or g75136 (po0526, n44842, n44843);
  and g75137 (n44845, pi0370, n_33393);
  and g75138 (n44846, pi1055, n44664);
  or g75139 (po0527, n44845, n44846);
  and g75140 (n44848, pi0371, n_33393);
  and g75141 (n44849, pi1051, n44664);
  or g75142 (po0528, n44848, n44849);
  and g75143 (n44851, pi0372, n_33393);
  and g75144 (n44852, pi1048, n44664);
  or g75145 (po0529, n44851, n44852);
  and g75146 (n44854, pi0373, n_33393);
  and g75147 (n44855, pi1087, n44664);
  or g75148 (po0530, n44854, n44855);
  and g75149 (n44857, pi0374, n_33393);
  and g75150 (n44858, pi1035, n44664);
  or g75151 (po0531, n44857, n44858);
  and g75152 (n44860, pi0375, n_33393);
  and g75153 (n44861, pi1047, n44664);
  or g75154 (po0532, n44860, n44861);
  and g75155 (n44863, pi0376, n_33393);
  and g75156 (n44864, pi1079, n44664);
  or g75157 (po0533, n44863, n44864);
  and g75158 (n44866, pi0377, n_33393);
  and g75159 (n44867, pi1074, n44664);
  or g75160 (po0534, n44866, n44867);
  and g75161 (n44869, pi0378, n_33393);
  and g75162 (n44870, pi1063, n44664);
  or g75163 (po0535, n44869, n44870);
  and g75164 (n44872, pi0379, n_33393);
  and g75165 (n44873, pi1045, n44664);
  or g75166 (po0536, n44872, n44873);
  and g75167 (n44875, pi0380, n_33393);
  and g75168 (n44876, pi1084, n44664);
  or g75169 (po0537, n44875, n44876);
  and g75170 (n44878, pi0381, n_33393);
  and g75171 (n44879, pi1081, n44664);
  or g75172 (po0538, n44878, n44879);
  and g75173 (n44881, pi0382, n_33393);
  and g75174 (n44882, pi1076, n44664);
  or g75175 (po0539, n44881, n44882);
  and g75176 (n44884, pi0383, n_33393);
  and g75177 (n44885, pi1071, n44664);
  or g75178 (po0540, n44884, n44885);
  and g75179 (n44887, pi0384, n_33393);
  and g75180 (n44888, pi1068, n44664);
  or g75181 (po0541, n44887, n44888);
  and g75182 (n44890, pi0385, n_33393);
  and g75183 (n44891, pi1042, n44664);
  or g75184 (po0542, n44890, n44891);
  and g75185 (n44893, pi0386, n_33393);
  and g75186 (n44894, pi1059, n44664);
  or g75187 (po0543, n44893, n44894);
  and g75188 (n44896, pi0387, n_33393);
  and g75189 (n44897, pi1053, n44664);
  or g75190 (po0544, n44896, n44897);
  and g75191 (n44899, pi0388, n_33393);
  and g75192 (n44900, pi1037, n44664);
  or g75193 (po0545, n44899, n44900);
  and g75194 (n44902, pi0389, n_33393);
  and g75195 (n44903, pi1036, n44664);
  or g75196 (po0546, n44902, n44903);
  and g75197 (n44905, pi0390, n_33397);
  and g75198 (n44906, pi1049, n44669);
  or g75199 (po0547, n44905, n44906);
  and g75200 (n44908, pi0391, n_33397);
  and g75201 (n44909, pi1062, n44669);
  or g75202 (po0548, n44908, n44909);
  and g75203 (n44911, pi0392, n_33397);
  and g75204 (n44912, pi1039, n44669);
  or g75205 (po0549, n44911, n44912);
  and g75206 (n44914, pi0393, n_33397);
  and g75207 (n44915, pi1067, n44669);
  or g75208 (po0550, n44914, n44915);
  and g75209 (n44917, pi0394, n_33397);
  and g75210 (n44918, pi1080, n44669);
  or g75211 (po0551, n44917, n44918);
  and g75212 (n44920, pi0395, n_33397);
  and g75213 (n44921, pi1055, n44669);
  or g75214 (po0552, n44920, n44921);
  and g75215 (n44923, pi0396, n_33397);
  and g75216 (n44924, pi1051, n44669);
  or g75217 (po0553, n44923, n44924);
  and g75218 (n44926, pi0397, n_33397);
  and g75219 (n44927, pi1048, n44669);
  or g75220 (po0554, n44926, n44927);
  and g75221 (n44929, pi0398, n_33397);
  and g75222 (n44930, pi1087, n44669);
  or g75223 (po0555, n44929, n44930);
  and g75224 (n44932, pi0399, n_33397);
  and g75225 (n44933, pi1047, n44669);
  or g75226 (po0556, n44932, n44933);
  and g75227 (n44935, pi0400, n_33397);
  and g75228 (n44936, pi1035, n44669);
  or g75229 (po0557, n44935, n44936);
  and g75230 (n44938, pi0401, n_33397);
  and g75231 (n44939, pi1079, n44669);
  or g75232 (po0558, n44938, n44939);
  and g75233 (n44941, pi0402, n_33397);
  and g75234 (n44942, pi1078, n44669);
  or g75235 (po0559, n44941, n44942);
  and g75236 (n44944, pi0403, n_33397);
  and g75237 (n44945, pi1045, n44669);
  or g75238 (po0560, n44944, n44945);
  and g75239 (n44947, pi0404, n_33397);
  and g75240 (n44948, pi1084, n44669);
  or g75241 (po0561, n44947, n44948);
  and g75242 (n44950, pi0405, n_33397);
  and g75243 (n44951, pi1081, n44669);
  or g75244 (po0562, n44950, n44951);
  and g75245 (n44953, pi0406, n_33397);
  and g75246 (n44954, pi1076, n44669);
  or g75247 (po0563, n44953, n44954);
  and g75248 (n44956, pi0407, n_33397);
  and g75249 (n44957, pi1071, n44669);
  or g75250 (po0564, n44956, n44957);
  and g75251 (n44959, pi0408, n_33397);
  and g75252 (n44960, pi1068, n44669);
  or g75253 (po0565, n44959, n44960);
  and g75254 (n44962, pi0409, n_33397);
  and g75255 (n44963, pi1042, n44669);
  or g75256 (po0566, n44962, n44963);
  and g75257 (n44965, pi0410, n_33397);
  and g75258 (n44966, pi1059, n44669);
  or g75259 (po0567, n44965, n44966);
  and g75260 (n44968, pi0411, n_33397);
  and g75261 (n44969, pi1053, n44669);
  or g75262 (po0568, n44968, n44969);
  and g75263 (n44971, pi0412, n_33397);
  and g75264 (n44972, pi1037, n44669);
  or g75265 (po0569, n44971, n44972);
  and g75266 (n44974, pi0413, n_33397);
  and g75267 (n44975, pi1036, n44669);
  or g75268 (po0570, n44974, n44975);
  and g75269 (n44977, n_4226, n44754);
  not g75270 (n_33440, n44977);
  and g75271 (n44978, pi0414, n_33440);
  and g75272 (n44979, pi1049, n44977);
  or g75273 (po0571, n44978, n44979);
  and g75274 (n44981, pi0415, n_33440);
  and g75275 (n44982, pi1062, n44977);
  or g75276 (po0572, n44981, n44982);
  and g75277 (n44984, pi0416, n_33440);
  and g75278 (n44985, pi1069, n44977);
  or g75279 (po0573, n44984, n44985);
  and g75280 (n44987, pi0417, n_33440);
  and g75281 (n44988, pi1039, n44977);
  or g75282 (po0574, n44987, n44988);
  and g75283 (n44990, pi0418, n_33440);
  and g75284 (n44991, pi1067, n44977);
  or g75285 (po0575, n44990, n44991);
  and g75286 (n44993, pi0419, n_33440);
  and g75287 (n44994, pi1080, n44977);
  or g75288 (po0576, n44993, n44994);
  and g75289 (n44996, pi0420, n_33440);
  and g75290 (n44997, pi1055, n44977);
  or g75291 (po0577, n44996, n44997);
  and g75292 (n44999, pi0421, n_33440);
  and g75293 (n45000, pi1051, n44977);
  or g75294 (po0578, n44999, n45000);
  and g75295 (n45002, pi0422, n_33440);
  and g75296 (n45003, pi1048, n44977);
  or g75297 (po0579, n45002, n45003);
  and g75298 (n45005, pi0423, n_33440);
  and g75299 (n45006, pi1087, n44977);
  or g75300 (po0580, n45005, n45006);
  and g75301 (n45008, pi0424, n_33440);
  and g75302 (n45009, pi1047, n44977);
  or g75303 (po0581, n45008, n45009);
  and g75304 (n45011, pi0425, n_33440);
  and g75305 (n45012, pi1035, n44977);
  or g75306 (po0582, n45011, n45012);
  and g75307 (n45014, pi0426, n_33440);
  and g75308 (n45015, pi1079, n44977);
  or g75309 (po0583, n45014, n45015);
  and g75310 (n45017, pi0427, n_33440);
  and g75311 (n45018, pi1078, n44977);
  or g75312 (po0584, n45017, n45018);
  and g75313 (n45020, pi0428, n_33440);
  and g75314 (n45021, pi1045, n44977);
  or g75315 (po0585, n45020, n45021);
  and g75316 (n45023, pi0429, n_33440);
  and g75317 (n45024, pi1084, n44977);
  or g75318 (po0586, n45023, n45024);
  and g75319 (n45026, pi0430, n_33440);
  and g75320 (n45027, pi1076, n44977);
  or g75321 (po0587, n45026, n45027);
  and g75322 (n45029, pi0431, n_33440);
  and g75323 (n45030, pi1071, n44977);
  or g75324 (po0588, n45029, n45030);
  and g75325 (n45032, pi0432, n_33440);
  and g75326 (n45033, pi1068, n44977);
  or g75327 (po0589, n45032, n45033);
  and g75328 (n45035, pi0433, n_33440);
  and g75329 (n45036, pi1042, n44977);
  or g75330 (po0590, n45035, n45036);
  and g75331 (n45038, pi0434, n_33440);
  and g75332 (n45039, pi1059, n44977);
  or g75333 (po0591, n45038, n45039);
  and g75334 (n45041, pi0435, n_33440);
  and g75335 (n45042, pi1053, n44977);
  or g75336 (po0592, n45041, n45042);
  and g75337 (n45044, pi0436, n_33440);
  and g75338 (n45045, pi1037, n44977);
  or g75339 (po0593, n45044, n45045);
  and g75340 (n45047, pi0437, n_33440);
  and g75341 (n45048, pi1070, n44977);
  or g75342 (po0594, n45047, n45048);
  and g75343 (n45050, pi0438, n_33440);
  and g75344 (n45051, pi1036, n44977);
  or g75345 (po0595, n45050, n45051);
  and g75346 (n45053, pi0439, n_33393);
  and g75347 (n45054, pi1057, n44664);
  or g75348 (po0596, n45053, n45054);
  and g75349 (n45056, pi0440, n_33393);
  and g75350 (n45057, pi1043, n44664);
  or g75351 (po0597, n45056, n45057);
  and g75352 (n45059, pi0441, n_33388);
  and g75353 (n45060, pi1044, n44657);
  or g75354 (po0598, n45059, n45060);
  and g75355 (n45062, pi0442, n_33393);
  and g75356 (n45063, pi1058, n44664);
  or g75357 (po0599, n45062, n45063);
  and g75358 (n45065, pi0443, n_33440);
  and g75359 (n45066, pi1044, n44977);
  or g75360 (po0600, n45065, n45066);
  and g75361 (n45068, pi0444, n_33440);
  and g75362 (n45069, pi1072, n44977);
  or g75363 (po0601, n45068, n45069);
  and g75364 (n45071, pi0445, n_33440);
  and g75365 (n45072, pi1081, n44977);
  or g75366 (po0602, n45071, n45072);
  and g75367 (n45074, pi0446, n_33440);
  and g75368 (n45075, pi1086, n44977);
  or g75369 (po0603, n45074, n45075);
  and g75370 (n45077, pi0447, n_33393);
  and g75371 (n45078, pi1040, n44664);
  or g75372 (po0604, n45077, n45078);
  and g75373 (n45080, pi0448, n_33440);
  and g75374 (n45081, pi1074, n44977);
  or g75375 (po0605, n45080, n45081);
  and g75376 (n45083, pi0449, n_33440);
  and g75377 (n45084, pi1057, n44977);
  or g75378 (po0606, n45083, n45084);
  and g75379 (n45086, pi0450, n_33388);
  and g75380 (n45087, pi1036, n44657);
  or g75381 (po0607, n45086, n45087);
  and g75382 (n45089, pi0451, n_33440);
  and g75383 (n45090, pi1063, n44977);
  or g75384 (po0608, n45089, n45090);
  and g75385 (n45092, pi0452, n_33388);
  and g75386 (n45093, pi1053, n44657);
  or g75387 (po0609, n45092, n45093);
  and g75388 (n45095, pi0453, n_33440);
  and g75389 (n45096, pi1040, n44977);
  or g75390 (po0610, n45095, n45096);
  and g75391 (n45098, pi0454, n_33440);
  and g75392 (n45099, pi1043, n44977);
  or g75393 (po0611, n45098, n45099);
  and g75394 (n45101, pi0455, n_33388);
  and g75395 (n45102, pi1037, n44657);
  or g75396 (po0612, n45101, n45102);
  and g75397 (n45104, pi0456, n_33397);
  and g75398 (n45105, pi1044, n44669);
  or g75399 (po0613, n45104, n45105);
  and g75400 (n45107, pi0594, pi0600);
  and g75401 (n45108, pi0597, n45107);
  and g75402 (n45109, pi0601, n45108);
  not g75403 (n_33447, pi0804);
  not g75404 (n_33448, pi0810);
  and g75405 (n45110, n_33447, n_33448);
  not g75406 (n_33450, pi0595);
  and g75407 (n45111, n_33450, n45110);
  not g75408 (n_33452, pi0599);
  and g75409 (n45112, n_33452, pi0810);
  not g75410 (n_33454, n45112);
  and g75411 (n45113, pi0596, n_33454);
  not g75412 (n_33455, n45113);
  and g75413 (n45114, pi0804, n_33455);
  and g75414 (n45115, pi0595, pi0815);
  not g75415 (n_33457, n45114);
  and g75416 (n45116, n_33457, n45115);
  not g75417 (n_33458, n45111);
  not g75418 (n_33459, n45116);
  and g75419 (n45117, n_33458, n_33459);
  not g75420 (n_33460, n45117);
  and g75421 (n45118, n45109, n_33460);
  and g75422 (n45119, pi0600, n_33448);
  not g75423 (n_33461, n45119);
  and g75424 (n45120, pi0804, n_33461);
  not g75425 (n_33462, pi0601);
  not g75426 (n_33463, n45110);
  and g75427 (n45121, n_33462, n_33463);
  not g75428 (n_33464, pi0815);
  not g75429 (n_33465, n45120);
  and g75430 (n45122, n_33464, n_33465);
  not g75431 (n_33466, n45121);
  and g75432 (n45123, n_33466, n45122);
  not g75433 (n_33467, n45118);
  not g75434 (n_33468, n45123);
  and g75435 (n45124, n_33467, n_33468);
  not g75436 (n_33470, n45124);
  and g75437 (n45125, pi0605, n_33470);
  and g75438 (n45126, pi0990, n45107);
  and g75439 (n45127, n_33464, n45120);
  and g75440 (n45128, n45126, n45127);
  not g75441 (n_33472, n45125);
  not g75442 (n_33473, n45128);
  and g75443 (n45129, n_33472, n_33473);
  not g75444 (n_33475, n45129);
  and g75445 (po0614, pi0821, n_33475);
  and g75446 (n45131, pi0458, n_33388);
  and g75447 (n45132, pi1072, n44657);
  or g75448 (po0615, n45131, n45132);
  and g75449 (n45134, pi0459, n_33440);
  and g75450 (n45135, pi1058, n44977);
  or g75451 (po0616, n45134, n45135);
  and g75452 (n45137, pi0460, n_33388);
  and g75453 (n45138, pi1086, n44657);
  or g75454 (po0617, n45137, n45138);
  and g75455 (n45140, pi0461, n_33388);
  and g75456 (n45141, pi1057, n44657);
  or g75457 (po0618, n45140, n45141);
  and g75458 (n45143, pi0462, n_33388);
  and g75459 (n45144, pi1074, n44657);
  or g75460 (po0619, n45143, n45144);
  and g75461 (n45146, pi0463, n_33397);
  and g75462 (n45147, pi1070, n44669);
  or g75463 (po0620, n45146, n45147);
  and g75464 (n45149, pi0464, n_33440);
  and g75465 (n45150, pi1065, n44977);
  or g75466 (po0621, n45149, n45150);
  and g75467 (n45152, n_234, n44561);
  not g75468 (n_33476, n11423);
  not g75469 (n_33477, n45152);
  and g75470 (n45153, n_33476, n_33477);
  not g75471 (n_33478, n11396);
  not g75472 (n_33479, n11399);
  and g75473 (n45154, n_33478, n_33479);
  not g75474 (n_33480, n45154);
  and g75475 (n45155, n_30428, n_33480);
  and g75476 (n45156, n_30428, pi1157);
  not g75477 (n_33481, n45153);
  not g75478 (n_33482, n45156);
  and g75479 (n45157, n_33481, n_33482);
  not g75480 (n_33483, n45155);
  and g75481 (n45158, n_33483, n45157);
  not g75482 (n_33484, n3471);
  not g75483 (n_33485, n11424);
  and g75484 (n45159, n_33484, n_33485);
  and g75485 (n45160, pi0926, n45156);
  not g75486 (n_33487, n45159);
  and g75487 (n45161, n_33487, n45160);
  not g75488 (n_33488, n5836);
  not g75489 (n_33489, n5854);
  and g75490 (n45162, n_33488, n_33489);
  not g75491 (n_33490, n45162);
  and g75492 (n45163, pi0926, n_33490);
  and g75493 (n45164, pi1157, n45162);
  not g75494 (n_33491, n45163);
  and g75495 (n45165, n_33483, n_33491);
  not g75496 (n_33492, n45164);
  and g75497 (n45166, n_33492, n45165);
  not g75498 (n_33493, n45158);
  not g75499 (n_33494, n45161);
  and g75500 (n45167, n_33493, n_33494);
  not g75501 (n_33495, n45166);
  and g75502 (n45168, n_33495, n45167);
  not g75503 (n_33496, n45168);
  and g75504 (n45169, n_4226, n_33496);
  and g75505 (n45170, n_30428, n44573);
  and g75506 (n45171, pi0926, n44575);
  not g75507 (n_33497, n5780);
  and g75508 (n45172, pi1157, n_33497);
  not g75515 (n_33501, n45169);
  not g75516 (n_33502, n45175);
  and g75517 (po0622, n_33501, n_33502);
  not g75518 (n_33503, n44573);
  and g75519 (n45177, po1038, n_33503);
  and g75520 (n45178, n_4226, n45154);
  not g75521 (n_33504, n45177);
  not g75522 (n_33505, n45178);
  and g75523 (n45179, n_33504, n_33505);
  not g75524 (n_33507, pi0943);
  not g75525 (n_33508, n45179);
  and g75526 (n45180, n_33507, n_33508);
  not g75527 (n_33509, n44571);
  and g75528 (n45181, n_33509, n45180);
  and g75529 (n45182, pi0943, n44624);
  not g75530 (n_33510, n45180);
  not g75531 (n_33511, n45182);
  and g75532 (n45183, n_33510, n_33511);
  not g75533 (n_33512, n45183);
  and g75534 (n45184, n_29468, n_33512);
  and g75535 (n45185, n_4226, n_33481);
  and g75536 (n45186, n2526, po1038);
  not g75537 (n_33513, n45185);
  not g75538 (n_33514, n45186);
  and g75539 (n45187, n_33513, n_33514);
  not g75540 (n_33515, n45187);
  and g75541 (n45188, n_32860, n_33515);
  and g75542 (n45189, n_33318, n_33350);
  and g75543 (n45190, pi0943, pi1151);
  not g75544 (n_33516, n45189);
  and g75545 (n45191, n_33516, n45190);
  and g75553 (n45195, pi0040, n_3084);
  and g75554 (n45196, n42346, n45195);
  and g75555 (n45197, po0950, n45196);
  not g75556 (n_33521, n10165);
  not g75557 (n_33522, n45197);
  and g75558 (n45198, n_33521, n_33522);
  not g75559 (n_33523, n13381);
  and g75560 (n45199, n_53, n_33523);
  not g75566 (n_33525, n45203);
  and g75567 (n45204, n45196, n_33525);
  not g75568 (n_33526, n45196);
  and g75569 (n45205, n_33526, n45203);
  not g75570 (n_33527, n45204);
  not g75571 (n_33528, n45205);
  and g75572 (n45206, n_33527, n_33528);
  not g75573 (n_33529, n45206);
  and g75574 (n45207, n7490, n_33529);
  and g75575 (n45208, n_7462, n_33529);
  and g75576 (n45209, n6277, n45203);
  not g75577 (n_33530, n45208);
  not g75578 (n_33531, n45209);
  and g75579 (n45210, n_33530, n_33531);
  not g75580 (n_33532, n45210);
  and g75581 (n45211, n_4126, n_33532);
  not g75582 (n_33533, n45207);
  and g75583 (n45212, pi1091, n_33533);
  not g75584 (n_33534, n45211);
  and g75585 (n45213, n_33534, n45212);
  and g75586 (n45214, n_3206, n_33532);
  and g75587 (n45215, n_7196, n_33529);
  and g75588 (n45216, n7417, n45203);
  not g75589 (n_33535, n45215);
  not g75590 (n_33536, n45216);
  and g75591 (n45217, n_33535, n_33536);
  not g75592 (n_33537, n45217);
  and g75593 (n45218, pi1093, n_33537);
  not g75594 (n_33538, n45214);
  and g75595 (n45219, n_3128, n_33538);
  not g75596 (n_33539, n45218);
  and g75597 (n45220, n_33539, n45219);
  not g75598 (n_33540, n45213);
  not g75599 (n_33541, n45220);
  and g75600 (n45221, n_33540, n_33541);
  and g75601 (n45222, n2610, n44644);
  not g75602 (n_33542, n45221);
  and g75603 (n45223, n_33542, n45222);
  not g75604 (n_33543, n45198);
  not g75605 (n_33544, n45223);
  and g75606 (po0624, n_33543, n_33544);
  and g75607 (n45225, n10200, n11337);
  not g75611 (n_33545, n45228);
  and g75612 (n45229, pi0468, n_33545);
  or g75613 (po0625, n45225, n45229);
  and g75614 (n45231, n_30417, n_33480);
  and g75615 (n45232, n_30417, pi1156);
  not g75616 (n_33546, n45232);
  and g75617 (n45233, n_33481, n_33546);
  not g75618 (n_33547, n45231);
  and g75619 (n45234, n_33547, n45233);
  and g75620 (n45235, pi0942, n45232);
  and g75621 (n45236, n_33487, n45235);
  and g75622 (n45237, pi0942, n_33490);
  and g75623 (n45238, pi1156, n45162);
  not g75624 (n_33549, n45237);
  and g75625 (n45239, n_33547, n_33549);
  not g75626 (n_33550, n45238);
  and g75627 (n45240, n_33550, n45239);
  not g75628 (n_33551, n45234);
  not g75629 (n_33552, n45236);
  and g75630 (n45241, n_33551, n_33552);
  not g75631 (n_33553, n45240);
  and g75632 (n45242, n_33553, n45241);
  not g75633 (n_33554, n45242);
  and g75634 (n45243, n_4226, n_33554);
  and g75635 (n45244, pi1156, n_33497);
  and g75636 (n45245, pi0942, n44575);
  and g75637 (n45246, n_30417, n44573);
  not g75644 (n_33558, n45243);
  not g75645 (n_33559, n45249);
  and g75646 (po0626, n_33558, n_33559);
  and g75647 (n45251, pi0267, n_33480);
  and g75648 (n45252, pi0267, pi1155);
  not g75649 (n_33560, n45252);
  and g75650 (n45253, n_33481, n_33560);
  not g75651 (n_33561, n45251);
  and g75652 (n45254, n_33561, n45253);
  and g75653 (n45255, pi0925, n45252);
  and g75654 (n45256, n_33487, n45255);
  and g75655 (n45257, pi0925, n_33490);
  and g75656 (n45258, pi1155, n45162);
  not g75657 (n_33563, n45257);
  and g75658 (n45259, n_33561, n_33563);
  not g75659 (n_33564, n45258);
  and g75660 (n45260, n_33564, n45259);
  not g75661 (n_33565, n45254);
  not g75662 (n_33566, n45256);
  and g75663 (n45261, n_33565, n_33566);
  not g75664 (n_33567, n45260);
  and g75665 (n45262, n_33567, n45261);
  not g75666 (n_33568, n45262);
  and g75667 (n45263, n_4226, n_33568);
  and g75668 (n45264, pi1155, n_33497);
  and g75669 (n45265, pi0925, n44575);
  and g75670 (n45266, pi0267, n44573);
  not g75677 (n_33572, n45263);
  not g75678 (n_33573, n45269);
  and g75679 (po0627, n_33572, n_33573);
  and g75680 (n45271, pi0253, n_33480);
  and g75681 (n45272, pi0253, pi1153);
  not g75682 (n_33574, n45272);
  and g75683 (n45273, n_33481, n_33574);
  not g75684 (n_33575, n45271);
  and g75685 (n45274, n_33575, n45273);
  and g75686 (n45275, pi0941, n45272);
  and g75687 (n45276, n_33487, n45275);
  and g75688 (n45277, pi0941, n_33490);
  and g75689 (n45278, pi1153, n45162);
  not g75690 (n_33577, n45277);
  and g75691 (n45279, n_33575, n_33577);
  not g75692 (n_33578, n45278);
  and g75693 (n45280, n_33578, n45279);
  not g75694 (n_33579, n45274);
  not g75695 (n_33580, n45276);
  and g75696 (n45281, n_33579, n_33580);
  not g75697 (n_33581, n45280);
  and g75698 (n45282, n_33581, n45281);
  not g75699 (n_33582, n45282);
  and g75700 (n45283, n_4226, n_33582);
  and g75701 (n45284, pi1153, n_33497);
  and g75702 (n45285, pi0941, n44575);
  and g75703 (n45286, pi0253, n44573);
  not g75710 (n_33586, n45283);
  not g75711 (n_33587, n45289);
  and g75712 (po0628, n_33586, n_33587);
  and g75713 (n45291, pi0254, n_33480);
  and g75714 (n45292, pi0254, pi1154);
  not g75715 (n_33588, n45292);
  and g75716 (n45293, n_33481, n_33588);
  not g75717 (n_33589, n45291);
  and g75718 (n45294, n_33589, n45293);
  and g75719 (n45295, pi0923, n45292);
  and g75720 (n45296, n_33487, n45295);
  and g75721 (n45297, pi0923, n_33490);
  and g75722 (n45298, pi1154, n45162);
  not g75723 (n_33591, n45297);
  and g75724 (n45299, n_33589, n_33591);
  not g75725 (n_33592, n45298);
  and g75726 (n45300, n_33592, n45299);
  not g75727 (n_33593, n45294);
  not g75728 (n_33594, n45296);
  and g75729 (n45301, n_33593, n_33594);
  not g75730 (n_33595, n45300);
  and g75731 (n45302, n_33595, n45301);
  not g75732 (n_33596, n45302);
  and g75733 (n45303, n_4226, n_33596);
  and g75734 (n45304, pi1154, n_33497);
  and g75735 (n45305, pi0923, n44575);
  and g75736 (n45306, pi0254, n44573);
  not g75743 (n_33600, n45303);
  not g75744 (n_33601, n45309);
  and g75745 (po0629, n_33600, n_33601);
  not g75746 (n_33603, pi0922);
  and g75747 (n45311, n_33603, n_33508);
  and g75748 (n45312, n_33509, n45311);
  and g75749 (n45313, pi0922, n44624);
  not g75750 (n_33604, n45311);
  not g75751 (n_33605, n45313);
  and g75752 (n45314, n_33604, n_33605);
  not g75753 (n_33606, n45314);
  and g75754 (n45315, n_28873, n_33606);
  and g75755 (n45316, n_32480, n_33515);
  and g75756 (n45317, pi0922, pi1152);
  and g75757 (n45318, n_33516, n45317);
  not g75765 (n_33612, pi0931);
  and g75766 (n45322, n_33612, n_33508);
  and g75767 (n45323, n_33509, n45322);
  and g75768 (n45324, pi0931, n44624);
  not g75769 (n_33613, n45322);
  not g75770 (n_33614, n45324);
  and g75771 (n45325, n_33613, n_33614);
  not g75772 (n_33615, n45325);
  and g75773 (n45326, n_30133, n_33615);
  and g75774 (n45327, n_32741, n_33515);
  and g75775 (n45328, pi0931, pi1150);
  and g75776 (n45329, n_33516, n45328);
  not g75784 (n_33621, pi0936);
  and g75785 (n45333, n_33621, n_33508);
  and g75786 (n45334, n_33509, n45333);
  and g75787 (n45335, pi0936, n44624);
  not g75788 (n_33622, n45333);
  not g75789 (n_33623, n45335);
  and g75790 (n45336, n_33622, n_33623);
  not g75791 (n_33624, n45336);
  and g75792 (n45337, n_29850, n_33624);
  and g75793 (n45338, n_32691, n_33515);
  and g75794 (n45339, pi0936, pi1149);
  and g75795 (n45340, n_33516, n45339);
  and g75803 (n45344, pi0071, n43509);
  and g75804 (n45345, pi0071, n_7411);
  and g75805 (n45346, n11448, n13052);
  and g75806 (n45347, n10150, n_7411);
  and g75807 (n45348, n10147, n45347);
  not g75808 (n_33629, n45346);
  not g75809 (n_33630, n45348);
  and g75810 (n45349, n_33629, n_33630);
  not g75815 (n_33632, n45345);
  not g75816 (n_33633, n45352);
  and g75817 (n45353, n_33632, n_33633);
  not g75818 (n_33634, n45353);
  and g75819 (n45354, n_4226, n_33634);
  or g75820 (po0633, n45344, n45354);
  and g75821 (po0635, pi0071, n_32791);
  and g75822 (n45357, pi0481, n_25717);
  and g75823 (n45358, pi0248, n34775);
  or g75824 (po0638, n45357, n45358);
  and g75825 (n45360, pi0482, n_25737);
  and g75826 (n45361, pi0249, n34791);
  or g75827 (po0639, n45360, n45361);
  and g75828 (n45363, pi0483, n_25845);
  and g75829 (n45364, pi0242, n34915);
  or g75830 (po0640, n45363, n45364);
  and g75831 (n45366, pi0484, n_25845);
  and g75832 (n45367, pi0249, n34915);
  or g75833 (po0641, n45366, n45367);
  and g75834 (n45369, pi0485, n_26758);
  and g75835 (n45370, pi0234, n36111);
  or g75836 (po0642, n45369, n45370);
  and g75837 (n45372, pi0486, n_26758);
  and g75838 (n45373, pi0244, n36111);
  or g75839 (po0643, n45372, n45373);
  and g75840 (n45375, pi0487, n_25717);
  and g75841 (n45376, pi0246, n34775);
  or g75842 (po0644, n45375, n45376);
  and g75843 (n45378, pi0488, n_25717);
  and g75844 (n45379, n_906, n34775);
  not g75845 (n_33643, n45378);
  not g75846 (n_33644, n45379);
  and g75847 (po0645, n_33643, n_33644);
  and g75848 (n45381, pi0489, n_26758);
  and g75849 (n45382, pi0242, n36111);
  or g75850 (po0646, n45381, n45382);
  and g75851 (n45384, pi0490, n_25845);
  and g75852 (n45385, pi0241, n34915);
  or g75853 (po0647, n45384, n45385);
  and g75854 (n45387, pi0491, n_25845);
  and g75855 (n45388, pi0238, n34915);
  or g75856 (po0648, n45387, n45388);
  and g75857 (n45390, pi0492, n_25845);
  and g75858 (n45391, pi0240, n34915);
  or g75859 (po0649, n45390, n45391);
  and g75860 (n45393, pi0493, n_25845);
  and g75861 (n45394, pi0244, n34915);
  or g75862 (po0650, n45393, n45394);
  and g75863 (n45396, pi0494, n_25845);
  and g75864 (n45397, n_906, n34915);
  not g75865 (n_33651, n45396);
  not g75866 (n_33652, n45397);
  and g75867 (po0651, n_33651, n_33652);
  and g75868 (n45399, pi0495, n_25845);
  and g75869 (n45400, pi0235, n34915);
  or g75870 (po0652, n45399, n45400);
  and g75871 (n45402, pi0496, n_25836);
  and g75872 (n45403, pi0249, n34907);
  or g75873 (po0653, n45402, n45403);
  and g75874 (n45405, pi0497, n_25836);
  and g75875 (n45406, n_906, n34907);
  not g75876 (n_33656, n45405);
  not g75877 (n_33657, n45406);
  and g75878 (po0654, n_33656, n_33657);
  and g75879 (n45408, pi0498, n_25737);
  and g75880 (n45409, pi0238, n34791);
  or g75881 (po0655, n45408, n45409);
  and g75882 (n45411, pi0499, n_25836);
  and g75883 (n45412, pi0246, n34907);
  or g75884 (po0656, n45411, n45412);
  and g75885 (n45414, pi0500, n_25836);
  and g75886 (n45415, pi0241, n34907);
  or g75887 (po0657, n45414, n45415);
  and g75888 (n45417, pi0501, n_25836);
  and g75889 (n45418, pi0248, n34907);
  or g75890 (po0658, n45417, n45418);
  and g75891 (n45420, pi0502, n_25836);
  and g75892 (n45421, pi0247, n34907);
  or g75893 (po0659, n45420, n45421);
  and g75894 (n45423, pi0503, n_25836);
  and g75895 (n45424, pi0245, n34907);
  or g75896 (po0660, n45423, n45424);
  and g75897 (n45426, pi0504, n_25828);
  and g75898 (n45427, pi0242, n34900);
  or g75899 (po0661, n45426, n45427);
  not g75900 (n_33665, n6326);
  and g75901 (n45429, n_33665, n16479);
  not g75902 (n_33666, n45429);
  and g75903 (n45430, n_25826, n_33666);
  and g75904 (n45431, n_148, n45430);
  and g75905 (n45432, n34907, n45431);
  not g75906 (n_33668, n45432);
  and g75907 (n45433, pi0505, n_33668);
  and g75908 (n45434, pi0234, n34899);
  not g75909 (n_33669, pi0505);
  and g75910 (n45435, n_33669, n34778);
  and g75911 (n45436, n45434, n45435);
  or g75912 (po0662, n45433, n45436);
  and g75913 (n45438, pi0506, n_25828);
  and g75914 (n45439, pi0241, n34900);
  or g75915 (po0663, n45438, n45439);
  and g75916 (n45441, pi0507, n_25828);
  and g75917 (n45442, pi0238, n34900);
  or g75918 (po0664, n45441, n45442);
  and g75919 (n45444, pi0508, n_25828);
  and g75920 (n45445, pi0247, n34900);
  or g75921 (po0665, n45444, n45445);
  and g75922 (n45447, pi0509, n_25828);
  and g75923 (n45448, pi0245, n34900);
  or g75924 (po0666, n45447, n45448);
  and g75925 (n45450, pi0510, n_25717);
  and g75926 (n45451, pi0242, n34775);
  or g75927 (po0667, n45450, n45451);
  and g75928 (n45453, n6584, n_4226);
  not g75929 (n_33675, n45453);
  and g75930 (n45454, n_25714, n_33675);
  and g75931 (n45455, n_148, n45454);
  not g75932 (n_33676, n45455);
  and g75933 (n45456, n34775, n_33676);
  and g75934 (n45457, pi0511, n_25717);
  or g75935 (po0668, n45456, n45457);
  and g75936 (n45459, pi0512, n_25717);
  and g75937 (n45460, pi0235, n34775);
  or g75938 (po0669, n45459, n45460);
  and g75939 (n45462, pi0513, n_25717);
  and g75940 (n45463, pi0244, n34775);
  or g75941 (po0670, n45462, n45463);
  and g75942 (n45465, pi0514, n_25717);
  and g75943 (n45466, pi0245, n34775);
  or g75944 (po0671, n45465, n45466);
  and g75945 (n45468, pi0515, n_25717);
  and g75946 (n45469, pi0240, n34775);
  or g75947 (po0672, n45468, n45469);
  and g75948 (n45471, pi0516, n_25717);
  and g75949 (n45472, pi0247, n34775);
  or g75950 (po0673, n45471, n45472);
  and g75951 (n45474, pi0517, n_25717);
  and g75952 (n45475, pi0238, n34775);
  or g75953 (po0674, n45474, n45475);
  and g75954 (n45477, n34783, n45455);
  not g75955 (n_33685, n45477);
  and g75956 (n45478, pi0518, n_33685);
  and g75957 (n45479, pi0234, n34774);
  not g75958 (n_33686, pi0518);
  and g75959 (n45480, n_33686, n34778);
  and g75960 (n45481, n45479, n45480);
  or g75961 (po0675, n45478, n45481);
  and g75962 (n45483, pi0519, n_25727);
  and g75963 (n45484, n_906, n34783);
  not g75964 (n_33688, n45483);
  not g75965 (n_33689, n45484);
  and g75966 (po0676, n_33688, n_33689);
  and g75967 (n45486, pi0520, n_25727);
  and g75968 (n45487, pi0246, n34783);
  or g75969 (po0677, n45486, n45487);
  and g75970 (n45489, pi0521, n_25727);
  and g75971 (n45490, pi0248, n34783);
  or g75972 (po0678, n45489, n45490);
  and g75973 (n45492, pi0522, n_25727);
  and g75974 (n45493, pi0238, n34783);
  or g75975 (po0679, n45492, n45493);
  and g75976 (n45495, n36139, n45455);
  not g75977 (n_33694, n45495);
  and g75978 (n45496, pi0523, n_33694);
  not g75979 (n_33695, pi0523);
  and g75980 (n45497, n_33695, n34910);
  and g75981 (n45498, n45479, n45497);
  or g75982 (po0680, n45496, n45498);
  and g75983 (n45500, pi0524, n_26778);
  and g75984 (n45501, n_906, n36139);
  not g75985 (n_33697, n45500);
  not g75986 (n_33698, n45501);
  and g75987 (po0681, n_33697, n_33698);
  and g75988 (n45503, pi0525, n_26778);
  and g75989 (n45504, pi0245, n36139);
  or g75990 (po0682, n45503, n45504);
  and g75991 (n45506, pi0526, n_26778);
  and g75992 (n45507, pi0246, n36139);
  or g75993 (po0683, n45506, n45507);
  and g75994 (n45509, pi0527, n_26778);
  and g75995 (n45510, pi0247, n36139);
  or g75996 (po0684, n45509, n45510);
  and g75997 (n45512, pi0528, n_26778);
  and g75998 (n45513, pi0249, n36139);
  or g75999 (po0685, n45512, n45513);
  and g76000 (n45515, pi0529, n_26778);
  and g76001 (n45516, pi0238, n36139);
  or g76002 (po0686, n45515, n45516);
  and g76003 (n45518, pi0530, n_26778);
  and g76004 (n45519, pi0240, n36139);
  or g76005 (po0687, n45518, n45519);
  and g76006 (n45521, pi0531, n_25737);
  and g76007 (n45522, pi0235, n34791);
  or g76008 (po0688, n45521, n45522);
  and g76009 (n45524, pi0532, n_25737);
  and g76010 (n45525, pi0247, n34791);
  or g76011 (po0689, n45524, n45525);
  and g76012 (n45527, pi0533, n_25828);
  and g76013 (n45528, pi0235, n34900);
  or g76014 (po0690, n45527, n45528);
  and g76015 (n45530, pi0534, n_25828);
  and g76016 (n45531, n_906, n34900);
  not g76017 (n_33709, n45530);
  not g76018 (n_33710, n45531);
  and g76019 (po0691, n_33709, n_33710);
  and g76020 (n45533, pi0535, n_25828);
  and g76021 (n45534, pi0240, n34900);
  or g76022 (po0692, n45533, n45534);
  and g76023 (n45536, pi0536, n_25828);
  and g76024 (n45537, pi0246, n34900);
  or g76025 (po0693, n45536, n45537);
  and g76026 (n45539, pi0537, n_25828);
  and g76027 (n45540, pi0248, n34900);
  or g76028 (po0694, n45539, n45540);
  and g76029 (n45542, pi0538, n_25828);
  and g76030 (n45543, pi0249, n34900);
  or g76031 (po0695, n45542, n45543);
  and g76032 (n45545, pi0539, n_25836);
  and g76033 (n45546, pi0242, n34907);
  or g76034 (po0696, n45545, n45546);
  and g76035 (n45548, pi0540, n_25836);
  and g76036 (n45549, pi0235, n34907);
  or g76037 (po0697, n45548, n45549);
  and g76038 (n45551, pi0541, n_25836);
  and g76039 (n45552, pi0244, n34907);
  or g76040 (po0698, n45551, n45552);
  and g76041 (n45554, pi0542, n_25836);
  and g76042 (n45555, pi0240, n34907);
  or g76043 (po0699, n45554, n45555);
  and g76044 (n45557, pi0543, n_25836);
  and g76045 (n45558, pi0238, n34907);
  or g76046 (po0700, n45557, n45558);
  and g76047 (n45560, n34915, n45431);
  not g76048 (n_33721, n45560);
  and g76049 (n45561, pi0544, n_33721);
  not g76050 (n_33722, pi0544);
  and g76051 (n45562, n_33722, n34910);
  and g76052 (n45563, n45434, n45562);
  or g76053 (po0701, n45561, n45563);
  and g76054 (n45565, pi0545, n_25845);
  and g76055 (n45566, pi0245, n34915);
  or g76056 (po0702, n45565, n45566);
  and g76057 (n45568, pi0546, n_25845);
  and g76058 (n45569, pi0246, n34915);
  or g76059 (po0703, n45568, n45569);
  and g76060 (n45571, pi0547, n_25845);
  and g76061 (n45572, pi0247, n34915);
  or g76062 (po0704, n45571, n45572);
  and g76063 (n45574, pi0548, n_25845);
  and g76064 (n45575, pi0248, n34915);
  or g76065 (po0705, n45574, n45575);
  and g76066 (n45577, pi0549, n_26758);
  and g76067 (n45578, pi0235, n36111);
  or g76068 (po0706, n45577, n45578);
  and g76069 (n45580, pi0550, n_26758);
  and g76070 (n45581, n_906, n36111);
  not g76071 (n_33729, n45580);
  not g76072 (n_33730, n45581);
  and g76073 (po0707, n_33729, n_33730);
  and g76074 (n45583, pi0551, n_26758);
  and g76075 (n45584, pi0240, n36111);
  or g76076 (po0708, n45583, n45584);
  and g76077 (n45586, pi0552, n_26758);
  and g76078 (n45587, pi0247, n36111);
  or g76079 (po0709, n45586, n45587);
  and g76080 (n45589, pi0553, n_26758);
  and g76081 (n45590, pi0241, n36111);
  or g76082 (po0710, n45589, n45590);
  and g76083 (n45592, pi0554, n_26758);
  and g76084 (n45593, pi0248, n36111);
  or g76085 (po0711, n45592, n45593);
  and g76086 (n45595, pi0555, n_26758);
  and g76087 (n45596, pi0249, n36111);
  or g76088 (po0712, n45595, n45596);
  and g76089 (n45598, pi0556, n_25737);
  and g76090 (n45599, pi0242, n34791);
  or g76091 (po0713, n45598, n45599);
  and g76092 (n45601, n34900, n45431);
  not g76093 (n_33738, n45601);
  and g76094 (n45602, pi0557, n_33738);
  not g76095 (n_33739, pi0557);
  and g76096 (n45603, n_33739, n34583);
  and g76097 (n45604, n45434, n45603);
  or g76098 (po0714, n45602, n45604);
  and g76099 (n45606, pi0558, n_25828);
  and g76100 (n45607, pi0244, n34900);
  or g76101 (po0715, n45606, n45607);
  and g76102 (n45609, pi0559, n_25717);
  and g76103 (n45610, pi0241, n34775);
  or g76104 (po0716, n45609, n45610);
  and g76105 (n45612, pi0560, n_25737);
  and g76106 (n45613, pi0240, n34791);
  or g76107 (po0717, n45612, n45613);
  and g76108 (n45615, pi0561, n_25727);
  and g76109 (n45616, pi0247, n34783);
  or g76110 (po0718, n45615, n45616);
  and g76111 (n45618, pi0562, n_25737);
  and g76112 (n45619, pi0241, n34791);
  or g76113 (po0719, n45618, n45619);
  and g76114 (n45621, pi0563, n_26758);
  and g76115 (n45622, pi0246, n36111);
  or g76116 (po0720, n45621, n45622);
  and g76117 (n45624, pi0564, n_25737);
  and g76118 (n45625, pi0246, n34791);
  or g76119 (po0721, n45624, n45625);
  and g76120 (n45627, pi0565, n_25737);
  and g76121 (n45628, pi0248, n34791);
  or g76122 (po0722, n45627, n45628);
  and g76123 (n45630, pi0566, n_25737);
  and g76124 (n45631, pi0244, n34791);
  or g76125 (po0723, n45630, n45631);
  and g76126 (n45633, n_4112, pi1092);
  and g76127 (n45634, n_3206, n45633);
  not g76132 (n_33749, n45634);
  and g76133 (n45639, n_12315, n_33749);
  not g76134 (n_33750, n45638);
  and g76135 (n45640, n_33750, n45639);
  and g76136 (n45641, n_11821, n45638);
  not g76137 (n_33751, n45641);
  and g76138 (n45642, n_33749, n_33751);
  not g76139 (n_33752, n45642);
  and g76140 (n45643, n_11405, n_33752);
  and g76141 (n45644, pi0619, n45638);
  not g76142 (n_33753, n45644);
  and g76143 (n45645, n_33749, n_33753);
  not g76144 (n_33754, n45645);
  and g76145 (n45646, pi1159, n_33754);
  not g76146 (n_33755, n45643);
  and g76147 (n45647, pi0789, n_33755);
  not g76148 (n_33756, n45646);
  and g76149 (n45648, n_33756, n45647);
  not g76150 (n_33757, n45640);
  not g76151 (n_33758, n45648);
  and g76152 (n45649, n_33757, n_33758);
  and g76153 (n45650, pi0680, n16826);
  and g76154 (n45651, n_13449, n45650);
  not g76155 (n_33759, n45651);
  and g76156 (n45652, n_33749, n_33759);
  not g76157 (n_33760, n45652);
  and g76158 (n45653, n19150, n_33760);
  and g76159 (n45654, n_11409, n45648);
  not g76160 (n_33761, n45654);
  and g76161 (n45655, n45653, n_33761);
  not g76162 (n_33762, n45649);
  not g76163 (n_33763, n45655);
  and g76164 (n45656, n_33762, n_33763);
  not g76165 (n_33764, n45656);
  and g76166 (n45657, n17970, n_33764);
  and g76167 (n45658, n35357, n45649);
  and g76168 (n45659, n_11780, n45653);
  and g76169 (n45660, pi0641, n45659);
  not g76170 (n_33765, n45660);
  and g76171 (n45661, n_33749, n_33765);
  not g76172 (n_33766, n45661);
  and g76173 (n45662, n17865, n_33766);
  and g76174 (n45663, n_11395, n45659);
  not g76175 (n_33767, n45663);
  and g76176 (n45664, n_33749, n_33767);
  not g76177 (n_33768, n45664);
  and g76178 (n45665, n17866, n_33768);
  not g76179 (n_33769, n45662);
  not g76180 (n_33770, n45665);
  and g76181 (n45666, n_33769, n_33770);
  not g76182 (n_33771, n45658);
  and g76183 (n45667, n_33771, n45666);
  not g76184 (n_33772, n45667);
  and g76185 (n45668, pi0788, n_33772);
  not g76186 (n_33773, n45657);
  not g76187 (n_33774, n45668);
  and g76188 (n45669, n_33773, n_33774);
  not g76189 (n_33775, n45669);
  and g76190 (n45670, n_14638, n_33775);
  and g76191 (n45671, n19151, n_33760);
  and g76192 (n45672, pi0628, n45671);
  not g76193 (n_33776, n45672);
  and g76194 (n45673, n_33749, n_33776);
  not g76195 (n_33777, n45673);
  and g76196 (n45674, pi1156, n_33777);
  and g76197 (n45675, n_12524, n45649);
  and g76198 (n45676, n17969, n45634);
  not g76199 (n_33778, n45675);
  not g76200 (n_33779, n45676);
  and g76201 (n45677, n_33778, n_33779);
  not g76202 (n_33780, n45677);
  and g76203 (n45678, n17854, n_33780);
  not g76204 (n_33781, n45674);
  and g76205 (n45679, n_12354, n_33781);
  not g76206 (n_33782, n45678);
  and g76207 (n45680, n_33782, n45679);
  and g76208 (n45681, n_11789, n45671);
  not g76209 (n_33783, n45681);
  and g76210 (n45682, n_33749, n_33783);
  not g76211 (n_33784, n45682);
  and g76212 (n45683, n_11794, n_33784);
  and g76213 (n45684, n17853, n_33780);
  not g76214 (n_33785, n45683);
  and g76215 (n45685, pi0629, n_33785);
  not g76216 (n_33786, n45684);
  and g76217 (n45686, n_33786, n45685);
  not g76218 (n_33787, n45680);
  and g76219 (n45687, pi0792, n_33787);
  not g76220 (n_33788, n45686);
  and g76221 (n45688, n_33788, n45687);
  not g76222 (n_33789, n45670);
  not g76223 (n_33790, n45688);
  and g76224 (n45689, n_33789, n_33790);
  not g76225 (n_33791, n45689);
  and g76226 (n45690, n_11806, n_33791);
  and g76227 (n45691, n_12368, n_33780);
  and g76228 (n45692, n17779, n45634);
  not g76229 (n_33792, n45691);
  not g76230 (n_33793, n45692);
  and g76231 (n45693, n_33792, n_33793);
  not g76232 (n_33794, n45693);
  and g76233 (n45694, pi0647, n_33794);
  not g76234 (n_33795, n45694);
  and g76235 (n45695, n_11810, n_33795);
  not g76236 (n_33796, n45690);
  and g76237 (n45696, n_33796, n45695);
  and g76238 (n45697, n_13453, n45671);
  and g76239 (n45698, pi0647, n45697);
  and g76240 (n45699, pi1157, n_33749);
  not g76241 (n_33797, n45698);
  and g76242 (n45700, n_33797, n45699);
  not g76243 (n_33798, n45700);
  and g76244 (n45701, n_12375, n_33798);
  not g76245 (n_33799, n45696);
  and g76246 (n45702, n_33799, n45701);
  and g76247 (n45703, pi0647, n_33791);
  and g76248 (n45704, n_11806, n_33794);
  not g76249 (n_33800, n45704);
  and g76250 (n45705, pi1157, n_33800);
  not g76251 (n_33801, n45703);
  and g76252 (n45706, n_33801, n45705);
  and g76253 (n45707, n_11806, n45697);
  and g76254 (n45708, n_11810, n_33749);
  not g76255 (n_33802, n45707);
  and g76256 (n45709, n_33802, n45708);
  not g76257 (n_33803, n45709);
  and g76258 (n45710, pi0630, n_33803);
  not g76259 (n_33804, n45706);
  and g76260 (n45711, n_33804, n45710);
  not g76261 (n_33805, n45702);
  not g76262 (n_33806, n45711);
  and g76263 (n45712, n_33805, n_33806);
  not g76264 (n_33807, n45712);
  and g76265 (n45713, pi0787, n_33807);
  and g76266 (n45714, n_11803, n_33791);
  not g76267 (n_33808, n45713);
  not g76268 (n_33809, n45714);
  and g76269 (n45715, n_33808, n_33809);
  not g76270 (n_33810, n45715);
  and g76271 (n45716, n_12411, n_33810);
  and g76272 (n45717, n_13598, n45697);
  not g76273 (n_33811, n45717);
  and g76274 (n45718, n_33749, n_33811);
  not g76275 (n_33812, n45718);
  and g76276 (n45719, pi0644, n_33812);
  and g76277 (n45720, n_11819, n_33810);
  not g76278 (n_33813, n45719);
  and g76279 (n45721, n_12395, n_33813);
  not g76280 (n_33814, n45720);
  and g76281 (n45722, n_33814, n45721);
  and g76282 (n45723, n_12392, n45691);
  and g76283 (n45724, n_11819, n45723);
  and g76284 (n45725, pi0715, n_33749);
  not g76285 (n_33815, n45724);
  and g76286 (n45726, n_33815, n45725);
  not g76287 (n_33816, n45722);
  not g76288 (n_33817, n45726);
  and g76289 (n45727, n_33816, n_33817);
  not g76290 (n_33818, n45727);
  and g76291 (n45728, n_12405, n_33818);
  and g76292 (n45729, pi0644, n45723);
  not g76293 (n_33819, n45729);
  and g76294 (n45730, n_33749, n_33819);
  not g76295 (n_33820, n45730);
  and g76296 (n45731, n_12395, n_33820);
  and g76297 (n45732, n_11819, n45718);
  and g76298 (n45733, pi0644, n45715);
  not g76299 (n_33821, n45732);
  and g76300 (n45734, pi0715, n_33821);
  not g76301 (n_33822, n45733);
  and g76302 (n45735, n_33822, n45734);
  not g76303 (n_33823, n45731);
  and g76304 (n45736, pi1160, n_33823);
  not g76305 (n_33824, n45735);
  and g76306 (n45737, n_33824, n45736);
  not g76307 (n_33825, n45737);
  and g76308 (n45738, pi0790, n_33825);
  not g76309 (n_33826, n45728);
  and g76310 (n45739, n_33826, n45738);
  not g76311 (n_33827, n45716);
  not g76312 (n_33828, n45739);
  and g76313 (n45740, n_33827, n_33828);
  not g76314 (n_33829, n45740);
  and g76315 (n45741, pi0230, n_33829);
  and g76316 (n45742, n_28510, n45633);
  or g76317 (po0724, n45741, n45742);
  and g76318 (n45744, pi0568, n_25737);
  and g76319 (n45745, pi0245, n34791);
  or g76320 (po0725, n45744, n45745);
  and g76321 (n45747, pi0569, n_25737);
  and g76322 (n45748, n_906, n34791);
  not g76323 (n_33832, n45747);
  not g76324 (n_33833, n45748);
  and g76325 (po0726, n_33832, n_33833);
  and g76326 (n45750, n34791, n45455);
  not g76327 (n_33835, n45750);
  and g76328 (n45751, pi0570, n_33835);
  not g76329 (n_33836, pi0570);
  and g76330 (n45752, n_33836, n34786);
  and g76331 (n45753, n45479, n45752);
  or g76332 (po0727, n45751, n45753);
  and g76333 (n45755, pi0571, n_26778);
  and g76334 (n45756, pi0241, n36139);
  or g76335 (po0728, n45755, n45756);
  and g76336 (n45758, pi0572, n_26778);
  and g76337 (n45759, pi0244, n36139);
  or g76338 (po0729, n45758, n45759);
  and g76339 (n45761, pi0573, n_26778);
  and g76340 (n45762, pi0242, n36139);
  or g76341 (po0730, n45761, n45762);
  and g76342 (n45764, pi0574, n_25727);
  and g76343 (n45765, pi0241, n34783);
  or g76344 (po0731, n45764, n45765);
  and g76345 (n45767, pi0575, n_26778);
  and g76346 (n45768, pi0235, n36139);
  or g76347 (po0732, n45767, n45768);
  and g76348 (n45770, pi0576, n_26778);
  and g76349 (n45771, pi0248, n36139);
  or g76350 (po0733, n45770, n45771);
  and g76351 (n45773, pi0577, n_26758);
  and g76352 (n45774, pi0238, n36111);
  or g76353 (po0734, n45773, n45774);
  and g76354 (n45776, pi0578, n_25727);
  and g76355 (n45777, pi0249, n34783);
  or g76356 (po0735, n45776, n45777);
  and g76357 (n45779, pi0579, n_25717);
  and g76358 (n45780, pi0249, n34775);
  or g76359 (po0736, n45779, n45780);
  and g76360 (n45782, pi0580, n_26758);
  and g76361 (n45783, pi0245, n36111);
  or g76362 (po0737, n45782, n45783);
  and g76363 (n45785, pi0581, n_25727);
  and g76364 (n45786, pi0235, n34783);
  or g76365 (po0738, n45785, n45786);
  and g76366 (n45788, pi0582, n_25727);
  and g76367 (n45789, pi0240, n34783);
  or g76368 (po0739, n45788, n45789);
  and g76369 (n45791, pi0584, n_25727);
  and g76370 (n45792, pi0245, n34783);
  or g76371 (po0741, n45791, n45792);
  and g76372 (n45794, pi0585, n_25727);
  and g76373 (n45795, pi0244, n34783);
  or g76374 (po0742, n45794, n45795);
  and g76375 (n45797, pi0586, n_25727);
  and g76376 (n45798, pi0242, n34783);
  or g76377 (po0743, n45797, n45798);
  and g76378 (n45800, n_28510, pi0587);
  or g76384 (po0744, n45800, n45805);
  and g76385 (n45807, n_31967, n12373);
  not g76386 (n_33852, n45807);
  and g76387 (n45808, n_4832, n_33852);
  and g76388 (n45809, n_4628, n45807);
  not g76389 (n_33853, n45808);
  and g76390 (n45810, n44706, n_33853);
  not g76391 (n_33854, n45809);
  and g76392 (po0745, n_33854, n45810);
  and g76393 (n45812, n_25822, n45430);
  and g76394 (n45813, n_25709, n45454);
  not g76395 (n_33855, n45812);
  and g76396 (n45814, pi0233, n_33855);
  not g76397 (n_33856, n45813);
  and g76398 (n45815, n_33856, n45814);
  and g76399 (n45816, n_25834, n45430);
  and g76400 (n45817, n_25725, n45454);
  not g76401 (n_33857, n45816);
  and g76402 (n45818, n_25720, n_33857);
  not g76403 (n_33858, n45817);
  and g76404 (n45819, n_33858, n45818);
  not g76405 (n_33859, n45815);
  not g76406 (n_33860, n45819);
  and g76407 (n45820, n_33859, n_33860);
  not g76408 (n_33861, n45820);
  and g76409 (n45821, pi0237, n_33861);
  and g76410 (n45822, n_25843, n45430);
  and g76411 (n45823, n_26776, n45454);
  not g76412 (n_33862, n45822);
  and g76413 (n45824, pi0233, n_33862);
  not g76414 (n_33863, n45823);
  and g76415 (n45825, n_33863, n45824);
  and g76416 (n45826, n_26756, n45430);
  and g76417 (n45827, n_25735, n45454);
  not g76418 (n_33864, n45826);
  and g76419 (n45828, n_25720, n_33864);
  not g76420 (n_33865, n45827);
  and g76421 (n45829, n_33865, n45828);
  not g76422 (n_33866, n45825);
  not g76423 (n_33867, n45829);
  and g76424 (n45830, n_33866, n_33867);
  not g76425 (n_33868, n45830);
  and g76426 (n45831, n_25730, n_33868);
  not g76427 (n_33869, n45821);
  not g76428 (n_33870, n45831);
  and g76429 (po0746, n_33869, n_33870);
  and g76430 (n45833, pi0588, n45807);
  and g76431 (n45834, pi0590, n_33852);
  not g76432 (n_33871, n45833);
  and g76433 (n45835, n44706, n_33871);
  not g76434 (n_33872, n45835);
  or g76435 (po0747, n45834, n_33872);
  and g76436 (n45837, n_4628, n_33852);
  and g76437 (n45838, n_4239, n45807);
  not g76438 (n_33873, n45837);
  and g76439 (n45839, n44706, n_33873);
  not g76440 (n_33874, n45838);
  and g76441 (po0748, n_33874, n45839);
  and g76442 (n45841, n_4239, n_33852);
  and g76443 (n45842, n_4423, n45807);
  not g76444 (n_33875, n45841);
  and g76445 (n45843, n44706, n_33875);
  not g76446 (n_33876, n45842);
  and g76447 (po0749, n_33876, n45843);
  and g76448 (n45845, pi0234, n45454);
  not g76449 (n_33877, n45845);
  and g76450 (n45846, pi0518, n_33877);
  not g76451 (n_33878, pi0520);
  and g76452 (n45847, pi0246, n_33878);
  and g76453 (n45848, n_2128, pi0520);
  not g76454 (n_33879, pi0578);
  and g76455 (n45849, pi0249, n_33879);
  and g76456 (n45850, n_1415, pi0578);
  not g76457 (n_33880, pi0521);
  and g76458 (n45851, pi0248, n_33880);
  and g76459 (n45852, n_1774, pi0521);
  and g76460 (n45853, pi0241, pi0574);
  not g76461 (n_33881, pi0574);
  and g76462 (n45854, n_1595, n_33881);
  not g76463 (n_33882, n45853);
  not g76464 (n_33883, n45854);
  and g76465 (n45855, n_33882, n_33883);
  and g76466 (n45856, n_33686, n_33676);
  and g76484 (n45865, pi0582, n45864);
  not g76485 (n_33893, n45865);
  and g76486 (n45866, pi0240, n_33893);
  not g76487 (n_33894, pi0582);
  and g76488 (n45867, n_33894, n45864);
  not g76489 (n_33895, n45867);
  and g76490 (n45868, n_2307, n_33895);
  not g76491 (n_33896, n45866);
  not g76492 (n_33897, n45868);
  and g76493 (n45869, n_33896, n_33897);
  and g76494 (n45870, n_906, pi0519);
  not g76495 (n_33898, pi0519);
  and g76496 (n45871, pi0239, n_33898);
  not g76497 (n_33899, n45870);
  not g76498 (n_33900, n45871);
  and g76499 (n45872, n_33899, n_33900);
  not g76500 (n_33901, n45872);
  and g76501 (n45873, n45869, n_33901);
  and g76502 (n45874, pi0242, pi0586);
  not g76503 (n_33902, pi0586);
  and g76504 (n45875, n_2915, n_33902);
  not g76505 (n_33903, n45874);
  not g76506 (n_33904, n45875);
  and g76507 (n45876, n_33903, n_33904);
  not g76508 (n_33905, n45876);
  and g76509 (n45877, n45873, n_33905);
  and g76510 (n45878, pi0235, pi0581);
  not g76511 (n_33906, pi0581);
  and g76512 (n45879, n_1106, n_33906);
  not g76513 (n_33907, n45878);
  not g76514 (n_33908, n45879);
  and g76515 (n45880, n_33907, n_33908);
  not g76516 (n_33909, n45880);
  and g76517 (n45881, n45877, n_33909);
  and g76518 (n45882, pi0585, n45881);
  not g76519 (n_33910, n45882);
  and g76520 (n45883, pi0244, n_33910);
  not g76521 (n_33911, pi0585);
  and g76522 (n45884, n_33911, n45881);
  not g76523 (n_33912, n45884);
  and g76524 (n45885, n_2688, n_33912);
  not g76525 (n_33913, n45883);
  not g76526 (n_33914, n45885);
  and g76527 (n45886, n_33913, n_33914);
  and g76528 (n45887, pi0584, n45886);
  not g76529 (n_33915, n45887);
  and g76530 (n45888, pi0245, n_33915);
  not g76531 (n_33916, pi0584);
  and g76532 (n45889, n_33916, n45886);
  not g76533 (n_33917, n45889);
  and g76534 (n45890, n_2498, n_33917);
  not g76535 (n_33918, n45888);
  not g76536 (n_33919, n45890);
  and g76537 (n45891, n_33918, n_33919);
  not g76538 (n_33920, pi0561);
  and g76539 (n45892, n_1955, n_33920);
  and g76540 (n45893, pi0247, pi0561);
  not g76541 (n_33921, n45892);
  not g76542 (n_33922, n45893);
  and g76543 (n45894, n_33921, n_33922);
  not g76544 (n_33923, n45894);
  and g76545 (n45895, n45891, n_33923);
  and g76546 (n45896, pi0238, n45895);
  and g76547 (n45897, pi0240, pi0542);
  not g76548 (n_33924, pi0542);
  and g76549 (n45898, n_2307, n_33924);
  not g76550 (n_33925, n45897);
  not g76551 (n_33926, n45898);
  and g76552 (n45899, n_33925, n_33926);
  not g76553 (n_33927, pi0501);
  and g76554 (n45900, n_1774, n_33927);
  and g76555 (n45901, pi0248, pi0501);
  not g76556 (n_33928, n45900);
  not g76557 (n_33929, n45901);
  and g76558 (n45902, n_33928, n_33929);
  and g76559 (n45903, pi0234, n45430);
  not g76560 (n_33930, n45903);
  and g76561 (n45904, pi0505, n_33930);
  not g76562 (n_33931, n45431);
  and g76563 (n45905, n_33669, n_33931);
  not g76564 (n_33932, pi0496);
  and g76565 (n45906, pi0249, n_33932);
  and g76566 (n45907, n_1415, pi0496);
  not g76567 (n_33933, pi0499);
  and g76568 (n45908, n_2128, n_33933);
  and g76569 (n45909, pi0246, pi0499);
  not g76570 (n_33934, n45908);
  not g76571 (n_33935, n45909);
  and g76572 (n45910, n_33934, n_33935);
  not g76584 (n_33942, pi0500);
  and g76585 (n45916, n_1595, n_33942);
  and g76586 (n45917, pi0241, pi0500);
  not g76587 (n_33943, n45916);
  not g76588 (n_33944, n45917);
  and g76589 (n45918, n_33943, n_33944);
  not g76590 (n_33945, n45918);
  and g76591 (n45919, n45915, n_33945);
  not g76592 (n_33946, n45899);
  and g76593 (n45920, n_33946, n45919);
  and g76594 (n45921, pi0497, n45920);
  not g76595 (n_33947, n45921);
  and g76596 (n45922, n_906, n_33947);
  not g76597 (n_33948, pi0497);
  and g76598 (n45923, n_33948, n45920);
  not g76599 (n_33949, n45923);
  and g76600 (n45924, pi0239, n_33949);
  not g76601 (n_33950, n45922);
  not g76602 (n_33951, n45924);
  and g76603 (n45925, n_33950, n_33951);
  and g76604 (n45926, pi0539, n45925);
  not g76605 (n_33952, n45926);
  and g76606 (n45927, pi0242, n_33952);
  not g76607 (n_33953, pi0539);
  and g76608 (n45928, n_33953, n45925);
  not g76609 (n_33954, n45928);
  and g76610 (n45929, n_2915, n_33954);
  not g76611 (n_33955, n45927);
  not g76612 (n_33956, n45929);
  and g76613 (n45930, n_33955, n_33956);
  and g76614 (n45931, pi0540, n45930);
  not g76615 (n_33957, n45931);
  and g76616 (n45932, pi0235, n_33957);
  not g76617 (n_33958, pi0540);
  and g76618 (n45933, n_33958, n45930);
  not g76619 (n_33959, n45933);
  and g76620 (n45934, n_1106, n_33959);
  not g76621 (n_33960, n45932);
  not g76622 (n_33961, n45934);
  and g76623 (n45935, n_33960, n_33961);
  and g76624 (n45936, pi0244, pi0541);
  not g76625 (n_33962, pi0541);
  and g76626 (n45937, n_2688, n_33962);
  not g76627 (n_33963, n45936);
  not g76628 (n_33964, n45937);
  and g76629 (n45938, n_33963, n_33964);
  not g76630 (n_33965, n45938);
  and g76631 (n45939, n45935, n_33965);
  and g76632 (n45940, pi0245, pi0503);
  not g76633 (n_33966, pi0503);
  and g76634 (n45941, n_2498, n_33966);
  not g76635 (n_33967, n45940);
  not g76636 (n_33968, n45941);
  and g76637 (n45942, n_33967, n_33968);
  not g76638 (n_33969, n45942);
  and g76639 (n45943, n45939, n_33969);
  not g76640 (n_33970, pi0502);
  and g76641 (n45944, n_33970, n45943);
  not g76642 (n_33971, n45944);
  and g76643 (n45945, n_1955, n_33971);
  and g76644 (n45946, pi0502, n45943);
  not g76645 (n_33972, n45946);
  and g76646 (n45947, pi0247, n_33972);
  not g76647 (n_33973, n45945);
  not g76648 (n_33974, n45947);
  and g76649 (n45948, n_33973, n_33974);
  and g76650 (n45949, n_1226, n45948);
  not g76651 (n_33975, n45896);
  and g76652 (n45950, pi0522, n_33975);
  not g76653 (n_33976, n45949);
  and g76654 (n45951, n_33976, n45950);
  and g76655 (n45952, n_33921, n_33973);
  not g76656 (n_33977, n45891);
  and g76657 (n45953, pi0502, n_33977);
  and g76658 (n45954, n_33942, n45919);
  and g76659 (n45955, n45915, n45917);
  not g76660 (n_33978, n45864);
  not g76661 (n_33979, n45955);
  and g76662 (n45956, n_33978, n_33979);
  not g76663 (n_33980, n45954);
  and g76664 (n45957, n_33980, n45956);
  not g76665 (n_33981, n45957);
  and g76666 (n45958, n_33894, n_33981);
  and g76667 (n45959, pi0582, n45919);
  not g76668 (n_33982, n45959);
  and g76669 (n45960, n_2307, n_33982);
  not g76670 (n_33983, n45958);
  and g76671 (n45961, n_33983, n45960);
  not g76672 (n_33984, n45961);
  and g76673 (n45962, n_33896, n_33984);
  not g76674 (n_33985, n45962);
  and g76675 (n45963, n_33924, n_33985);
  and g76676 (n45964, pi0582, n_33981);
  and g76677 (n45965, n_33894, n45919);
  not g76678 (n_33986, n45965);
  and g76679 (n45966, pi0240, n_33986);
  not g76680 (n_33987, n45964);
  and g76681 (n45967, n_33987, n45966);
  not g76682 (n_33988, n45967);
  and g76683 (n45968, n_33897, n_33988);
  not g76684 (n_33989, n45968);
  and g76685 (n45969, pi0542, n_33989);
  not g76686 (n_33990, n45963);
  not g76687 (n_33991, n45969);
  and g76688 (n45970, n_33990, n_33991);
  and g76689 (n45971, n_33948, n45970);
  and g76690 (n45972, pi0497, n45869);
  not g76691 (n_33992, n45972);
  and g76692 (n45973, pi0239, n_33992);
  not g76693 (n_33993, n45971);
  and g76694 (n45974, n_33993, n45973);
  not g76695 (n_33994, n45974);
  and g76696 (n45975, n_33950, n_33994);
  not g76697 (n_33995, n45975);
  and g76698 (n45976, n_33898, n_33995);
  and g76699 (n45977, pi0497, n45970);
  and g76700 (n45978, n_33948, n45869);
  not g76701 (n_33996, n45978);
  and g76702 (n45979, n_906, n_33996);
  not g76703 (n_33997, n45977);
  and g76704 (n45980, n_33997, n45979);
  not g76705 (n_33998, n45980);
  and g76706 (n45981, n_33951, n_33998);
  not g76707 (n_33999, n45981);
  and g76708 (n45982, pi0519, n_33999);
  not g76709 (n_34000, n45976);
  not g76710 (n_34001, n45982);
  and g76711 (n45983, n_34000, n_34001);
  and g76712 (n45984, n_33953, n45983);
  and g76713 (n45985, pi0539, n45873);
  not g76714 (n_34002, n45985);
  and g76715 (n45986, n_2915, n_34002);
  not g76716 (n_34003, n45984);
  and g76717 (n45987, n_34003, n45986);
  not g76718 (n_34004, n45987);
  and g76719 (n45988, n_33955, n_34004);
  not g76720 (n_34005, n45988);
  and g76721 (n45989, n_33902, n_34005);
  and g76722 (n45990, pi0539, n45983);
  and g76723 (n45991, n_33953, n45873);
  not g76724 (n_34006, n45991);
  and g76725 (n45992, pi0242, n_34006);
  not g76726 (n_34007, n45990);
  and g76727 (n45993, n_34007, n45992);
  not g76728 (n_34008, n45993);
  and g76729 (n45994, n_33956, n_34008);
  not g76730 (n_34009, n45994);
  and g76731 (n45995, pi0586, n_34009);
  not g76732 (n_34010, n45989);
  not g76733 (n_34011, n45995);
  and g76734 (n45996, n_34010, n_34011);
  and g76735 (n45997, n_33958, n45996);
  and g76736 (n45998, pi0540, n45877);
  not g76737 (n_34012, n45998);
  and g76738 (n45999, n_1106, n_34012);
  not g76739 (n_34013, n45997);
  and g76740 (n46000, n_34013, n45999);
  not g76741 (n_34014, n46000);
  and g76742 (n46001, n_33960, n_34014);
  not g76743 (n_34015, n46001);
  and g76744 (n46002, n_33906, n_34015);
  and g76745 (n46003, pi0540, n45996);
  and g76746 (n46004, n_33958, n45877);
  not g76747 (n_34016, n46004);
  and g76748 (n46005, pi0235, n_34016);
  not g76749 (n_34017, n46003);
  and g76750 (n46006, n_34017, n46005);
  not g76751 (n_34018, n46006);
  and g76752 (n46007, n_33961, n_34018);
  not g76753 (n_34019, n46007);
  and g76754 (n46008, pi0581, n_34019);
  not g76755 (n_34020, n46002);
  not g76756 (n_34021, n46008);
  and g76757 (n46009, n_34020, n_34021);
  and g76758 (n46010, n_33911, n46009);
  and g76759 (n46011, pi0585, n45935);
  not g76760 (n_34022, n46011);
  and g76761 (n46012, n_2688, n_34022);
  not g76762 (n_34023, n46010);
  and g76763 (n46013, n_34023, n46012);
  not g76764 (n_34024, n46013);
  and g76765 (n46014, n_33913, n_34024);
  not g76766 (n_34025, n46014);
  and g76767 (n46015, n_33962, n_34025);
  and g76768 (n46016, pi0585, n46009);
  and g76769 (n46017, n_33911, n45935);
  not g76770 (n_34026, n46017);
  and g76771 (n46018, pi0244, n_34026);
  not g76772 (n_34027, n46016);
  and g76773 (n46019, n_34027, n46018);
  not g76774 (n_34028, n46019);
  and g76775 (n46020, n_33914, n_34028);
  not g76776 (n_34029, n46020);
  and g76777 (n46021, pi0541, n_34029);
  not g76778 (n_34030, n46015);
  not g76779 (n_34031, n46021);
  and g76780 (n46022, n_34030, n_34031);
  and g76781 (n46023, n_33916, n46022);
  and g76782 (n46024, pi0584, n45939);
  not g76783 (n_34032, n46024);
  and g76784 (n46025, n_2498, n_34032);
  not g76785 (n_34033, n46023);
  and g76786 (n46026, n_34033, n46025);
  not g76787 (n_34034, n46026);
  and g76788 (n46027, n_33918, n_34034);
  not g76789 (n_34035, n46027);
  and g76790 (n46028, n_33966, n_34035);
  and g76791 (n46029, pi0584, n46022);
  and g76792 (n46030, n_33916, n45939);
  not g76793 (n_34036, n46030);
  and g76794 (n46031, pi0245, n_34036);
  not g76795 (n_34037, n46029);
  and g76796 (n46032, n_34037, n46031);
  not g76797 (n_34038, n46032);
  and g76798 (n46033, n_33919, n_34038);
  not g76799 (n_34039, n46033);
  and g76800 (n46034, pi0503, n_34039);
  not g76801 (n_34040, n46028);
  not g76802 (n_34041, n46034);
  and g76803 (n46035, n_34040, n_34041);
  not g76804 (n_34042, n46035);
  and g76805 (n46036, n_33970, n_34042);
  not g76806 (n_34043, n45953);
  and g76807 (n46037, n_33920, n_34043);
  not g76808 (n_34044, n46036);
  and g76809 (n46038, n_34044, n46037);
  not g76810 (n_34045, n45952);
  not g76811 (n_34046, n46038);
  and g76812 (n46039, n_34045, n_34046);
  and g76813 (n46040, n_33922, n_33974);
  and g76814 (n46041, n_33970, n_33977);
  and g76815 (n46042, pi0502, n_34042);
  not g76816 (n_34047, n46041);
  and g76817 (n46043, pi0561, n_34047);
  not g76818 (n_34048, n46042);
  and g76819 (n46044, n_34048, n46043);
  not g76820 (n_34049, n46040);
  not g76821 (n_34050, n46044);
  and g76822 (n46045, n_34049, n_34050);
  not g76823 (n_34051, n46039);
  not g76824 (n_34052, n46045);
  and g76825 (n46046, n_34051, n_34052);
  and g76826 (n46047, n_1226, n46046);
  not g76827 (n_34053, pi0522);
  not g76828 (n_34054, n46047);
  and g76829 (n46048, n_34053, n_34054);
  not g76830 (n_34055, pi0543);
  not g76831 (n_34056, n45951);
  and g76832 (n46049, n_34055, n_34056);
  not g76833 (n_34057, n46048);
  and g76834 (n46050, n_34057, n46049);
  and g76835 (n46051, n_1226, n45895);
  and g76836 (n46052, pi0238, n45948);
  not g76837 (n_34058, n46051);
  and g76838 (n46053, n_34053, n_34058);
  not g76839 (n_34059, n46052);
  and g76840 (n46054, n_34059, n46053);
  and g76841 (n46055, pi0238, n46046);
  not g76842 (n_34060, n46055);
  and g76843 (n46056, pi0522, n_34060);
  not g76844 (n_34061, n46054);
  and g76845 (n46057, pi0543, n_34061);
  not g76846 (n_34062, n46056);
  and g76847 (n46058, n_34062, n46057);
  not g76848 (n_34063, n46050);
  not g76849 (n_34064, n46058);
  and g76850 (n46059, n_34063, n_34064);
  not g76851 (n_34065, n46059);
  and g76852 (n46060, n_25720, n_34065);
  and g76853 (n46061, pi0246, pi0536);
  not g76854 (n_34066, pi0536);
  and g76855 (n46062, n_2128, n_34066);
  not g76856 (n_34067, n46061);
  not g76857 (n_34068, n46062);
  and g76858 (n46063, n_34067, n_34068);
  and g76859 (n46064, n_33739, n_33931);
  and g76860 (n46065, pi0557, n_33930);
  not g76861 (n_34069, n46063);
  not g76862 (n_34070, n46064);
  and g76863 (n46066, n_34069, n_34070);
  not g76864 (n_34071, n46065);
  and g76865 (n46067, n_34071, n46066);
  not g76866 (n_34072, pi0538);
  and g76867 (n46068, n_34072, n46067);
  not g76868 (n_34073, n46068);
  and g76869 (n46069, n_1415, n_34073);
  and g76870 (n46070, pi0538, n46067);
  not g76871 (n_34074, n46070);
  and g76872 (n46071, pi0249, n_34074);
  not g76873 (n_34075, n46069);
  not g76874 (n_34076, n46071);
  and g76875 (n46072, n_34075, n_34076);
  not g76876 (n_34077, pi0537);
  and g76877 (n46073, n_34077, n46072);
  not g76878 (n_34078, n46073);
  and g76879 (n46074, n_1774, n_34078);
  and g76880 (n46075, pi0537, n46072);
  not g76881 (n_34079, n46075);
  and g76882 (n46076, pi0248, n_34079);
  not g76883 (n_34080, n46074);
  not g76884 (n_34081, n46076);
  and g76885 (n46077, n_34080, n_34081);
  and g76886 (n46078, pi0241, pi0506);
  not g76887 (n_34082, pi0506);
  and g76888 (n46079, n_1595, n_34082);
  not g76889 (n_34083, n46078);
  not g76890 (n_34084, n46079);
  and g76891 (n46080, n_34083, n_34084);
  not g76892 (n_34085, n46080);
  and g76893 (n46081, n46077, n_34085);
  and g76894 (n46082, pi0240, pi0535);
  not g76895 (n_34086, pi0535);
  and g76896 (n46083, n_2307, n_34086);
  not g76897 (n_34087, n46082);
  not g76898 (n_34088, n46083);
  and g76899 (n46084, n_34087, n_34088);
  not g76900 (n_34089, n46084);
  and g76901 (n46085, n46081, n_34089);
  and g76902 (n46086, pi0534, n46085);
  not g76903 (n_34090, n46086);
  and g76904 (n46087, n_906, n_34090);
  not g76905 (n_34091, pi0534);
  and g76906 (n46088, n_34091, n46085);
  not g76907 (n_34092, n46088);
  and g76908 (n46089, pi0239, n_34092);
  not g76909 (n_34093, n46087);
  not g76910 (n_34094, n46089);
  and g76911 (n46090, n_34093, n_34094);
  and g76912 (n46091, pi0504, n46090);
  not g76913 (n_34095, n46091);
  and g76914 (n46092, pi0242, n_34095);
  not g76915 (n_34096, pi0504);
  and g76916 (n46093, n_34096, n46090);
  not g76917 (n_34097, n46093);
  and g76918 (n46094, n_2915, n_34097);
  not g76919 (n_34098, n46092);
  not g76920 (n_34099, n46094);
  and g76921 (n46095, n_34098, n_34099);
  and g76922 (n46096, pi0533, n46095);
  not g76923 (n_34100, n46096);
  and g76924 (n46097, pi0235, n_34100);
  not g76925 (n_34101, pi0533);
  and g76926 (n46098, n_34101, n46095);
  not g76927 (n_34102, n46098);
  and g76928 (n46099, n_1106, n_34102);
  not g76929 (n_34103, n46097);
  not g76930 (n_34104, n46099);
  and g76931 (n46100, n_34103, n_34104);
  and g76932 (n46101, pi0558, n46100);
  not g76933 (n_34105, n46101);
  and g76934 (n46102, pi0244, n_34105);
  not g76935 (n_34106, pi0558);
  and g76936 (n46103, n_34106, n46100);
  not g76937 (n_34107, n46103);
  and g76938 (n46104, n_2688, n_34107);
  not g76939 (n_34108, n46102);
  not g76940 (n_34109, n46104);
  and g76941 (n46105, n_34108, n_34109);
  and g76942 (n46106, pi0509, n46105);
  not g76943 (n_34110, n46106);
  and g76944 (n46107, pi0245, n_34110);
  not g76945 (n_34111, pi0509);
  and g76946 (n46108, n_34111, n46105);
  not g76947 (n_34112, n46108);
  and g76948 (n46109, n_2498, n_34112);
  not g76949 (n_34113, n46107);
  not g76950 (n_34114, n46109);
  and g76951 (n46110, n_34113, n_34114);
  and g76952 (n46111, pi0508, n46110);
  not g76953 (n_34115, n46111);
  and g76954 (n46112, pi0247, n_34115);
  not g76955 (n_34116, pi0508);
  and g76956 (n46113, n_34116, n46110);
  not g76957 (n_34117, n46113);
  and g76958 (n46114, n_1955, n_34117);
  not g76959 (n_34118, n46112);
  not g76960 (n_34119, n46114);
  and g76961 (n46115, n_34118, n_34119);
  and g76962 (n46116, n_1226, n46115);
  and g76963 (n46117, pi0248, pi0481);
  not g76964 (n_34120, pi0481);
  and g76965 (n46118, n_1774, n_34120);
  not g76966 (n_34121, n46117);
  not g76967 (n_34122, n46118);
  and g76968 (n46119, n_34121, n_34122);
  and g76969 (n46120, pi0246, pi0487);
  not g76970 (n_34123, pi0487);
  and g76971 (n46121, n_2128, n_34123);
  not g76972 (n_34124, n46120);
  not g76973 (n_34125, n46121);
  and g76974 (n46122, n_34124, n_34125);
  not g76975 (n_34126, pi0511);
  and g76976 (n46123, n_34126, n_33676);
  and g76977 (n46124, pi0511, n_33877);
  not g76978 (n_34127, n46122);
  not g76979 (n_34128, n46123);
  and g76980 (n46125, n_34127, n_34128);
  not g76981 (n_34129, n46124);
  and g76982 (n46126, n_34129, n46125);
  not g76983 (n_34130, pi0579);
  and g76984 (n46127, n_1415, n_34130);
  and g76985 (n46128, pi0249, pi0579);
  not g76986 (n_34131, n46127);
  not g76987 (n_34132, n46128);
  and g76988 (n46129, n_34131, n_34132);
  not g76989 (n_34133, n46129);
  and g76990 (n46130, n46126, n_34133);
  not g76991 (n_34134, n46119);
  and g76992 (n46131, n_34134, n46130);
  and g76993 (n46132, pi0559, n46131);
  not g76994 (n_34135, n46132);
  and g76995 (n46133, pi0241, n_34135);
  not g76996 (n_34136, pi0559);
  and g76997 (n46134, n_34136, n46131);
  not g76998 (n_34137, n46134);
  and g76999 (n46135, n_1595, n_34137);
  not g77000 (n_34138, n46133);
  not g77001 (n_34139, n46135);
  and g77002 (n46136, n_34138, n_34139);
  and g77003 (n46137, pi0515, n46136);
  not g77004 (n_34140, n46137);
  and g77005 (n46138, pi0240, n_34140);
  not g77006 (n_34141, pi0515);
  and g77007 (n46139, n_34141, n46136);
  not g77008 (n_34142, n46139);
  and g77009 (n46140, n_2307, n_34142);
  not g77010 (n_34143, n46138);
  not g77011 (n_34144, n46140);
  and g77012 (n46141, n_34143, n_34144);
  and g77013 (n46142, n_906, pi0488);
  not g77014 (n_34145, pi0488);
  and g77015 (n46143, pi0239, n_34145);
  not g77016 (n_34146, n46142);
  not g77017 (n_34147, n46143);
  and g77018 (n46144, n_34146, n_34147);
  not g77019 (n_34148, n46144);
  and g77020 (n46145, n46141, n_34148);
  and g77021 (n46146, pi0242, pi0510);
  not g77022 (n_34149, pi0510);
  and g77023 (n46147, n_2915, n_34149);
  not g77024 (n_34150, n46146);
  not g77025 (n_34151, n46147);
  and g77026 (n46148, n_34150, n_34151);
  not g77027 (n_34152, n46148);
  and g77028 (n46149, n46145, n_34152);
  and g77029 (n46150, pi0235, pi0512);
  not g77030 (n_34153, pi0512);
  and g77031 (n46151, n_1106, n_34153);
  not g77032 (n_34154, n46150);
  not g77033 (n_34155, n46151);
  and g77034 (n46152, n_34154, n_34155);
  not g77035 (n_34156, n46152);
  and g77036 (n46153, n46149, n_34156);
  and g77037 (n46154, pi0244, pi0513);
  not g77038 (n_34157, pi0513);
  and g77039 (n46155, n_2688, n_34157);
  not g77040 (n_34158, n46154);
  not g77041 (n_34159, n46155);
  and g77042 (n46156, n_34158, n_34159);
  not g77043 (n_34160, n46156);
  and g77044 (n46157, n46153, n_34160);
  and g77045 (n46158, pi0245, pi0514);
  not g77046 (n_34161, pi0514);
  and g77047 (n46159, n_2498, n_34161);
  not g77048 (n_34162, n46158);
  not g77049 (n_34163, n46159);
  and g77050 (n46160, n_34162, n_34163);
  not g77051 (n_34164, n46160);
  and g77052 (n46161, n46157, n_34164);
  and g77053 (n46162, pi0247, pi0516);
  not g77054 (n_34165, pi0516);
  and g77055 (n46163, n_1955, n_34165);
  not g77056 (n_34166, n46162);
  not g77057 (n_34167, n46163);
  and g77058 (n46164, n_34166, n_34167);
  not g77059 (n_34168, n46164);
  and g77060 (n46165, n46161, n_34168);
  and g77061 (n46166, pi0238, n46165);
  not g77062 (n_34169, n46166);
  and g77063 (n46167, pi0517, n_34169);
  not g77064 (n_34170, n46116);
  and g77065 (n46168, n_34170, n46167);
  not g77066 (n_34171, n46130);
  and g77067 (n46169, n_34130, n_34171);
  and g77068 (n46170, n_34075, n46126);
  not g77069 (n_34172, n46170);
  and g77070 (n46171, pi0579, n_34172);
  not g77071 (n_34173, n46169);
  not g77072 (n_34174, n46171);
  and g77073 (n46172, n_34173, n_34174);
  not g77074 (n_34175, n46072);
  not g77075 (n_34176, n46172);
  and g77076 (n46173, n_34175, n_34176);
  not g77077 (n_34177, n46173);
  and g77078 (n46174, n_34077, n_34177);
  and g77079 (n46175, pi0537, n46130);
  not g77080 (n_34178, n46175);
  and g77081 (n46176, n_1774, n_34178);
  not g77082 (n_34179, n46174);
  and g77083 (n46177, n_34179, n46176);
  not g77084 (n_34180, n46177);
  and g77085 (n46178, n_34081, n_34180);
  not g77086 (n_34181, n46178);
  and g77087 (n46179, n_34120, n_34181);
  and g77088 (n46180, pi0537, n_34177);
  and g77089 (n46181, n_34077, n46130);
  not g77090 (n_34182, n46181);
  and g77091 (n46182, pi0248, n_34182);
  not g77092 (n_34183, n46180);
  and g77093 (n46183, n_34183, n46182);
  not g77094 (n_34184, n46183);
  and g77095 (n46184, n_34080, n_34184);
  not g77096 (n_34185, n46184);
  and g77097 (n46185, pi0481, n_34185);
  not g77098 (n_34186, n46179);
  not g77099 (n_34187, n46185);
  and g77100 (n46186, n_34186, n_34187);
  and g77101 (n46187, n_34136, n46186);
  and g77102 (n46188, pi0559, n46077);
  not g77103 (n_34188, n46188);
  and g77104 (n46189, n_1595, n_34188);
  not g77105 (n_34189, n46187);
  and g77106 (n46190, n_34189, n46189);
  not g77107 (n_34190, n46190);
  and g77108 (n46191, n_34138, n_34190);
  not g77109 (n_34191, n46191);
  and g77110 (n46192, n_34082, n_34191);
  and g77111 (n46193, pi0559, n46186);
  and g77112 (n46194, n_34136, n46077);
  not g77113 (n_34192, n46194);
  and g77114 (n46195, pi0241, n_34192);
  not g77115 (n_34193, n46193);
  and g77116 (n46196, n_34193, n46195);
  not g77117 (n_34194, n46196);
  and g77118 (n46197, n_34139, n_34194);
  not g77119 (n_34195, n46197);
  and g77120 (n46198, pi0506, n_34195);
  not g77121 (n_34196, n46192);
  not g77122 (n_34197, n46198);
  and g77123 (n46199, n_34196, n_34197);
  and g77124 (n46200, n_34141, n46199);
  and g77125 (n46201, pi0515, n46081);
  not g77126 (n_34198, n46201);
  and g77127 (n46202, n_2307, n_34198);
  not g77128 (n_34199, n46200);
  and g77129 (n46203, n_34199, n46202);
  not g77130 (n_34200, n46203);
  and g77131 (n46204, n_34143, n_34200);
  not g77132 (n_34201, n46204);
  and g77133 (n46205, n_34086, n_34201);
  and g77134 (n46206, pi0515, n46199);
  and g77135 (n46207, n_34141, n46081);
  not g77136 (n_34202, n46207);
  and g77137 (n46208, pi0240, n_34202);
  not g77138 (n_34203, n46206);
  and g77139 (n46209, n_34203, n46208);
  not g77140 (n_34204, n46209);
  and g77141 (n46210, n_34144, n_34204);
  not g77142 (n_34205, n46210);
  and g77143 (n46211, pi0535, n_34205);
  not g77144 (n_34206, n46205);
  not g77145 (n_34207, n46211);
  and g77146 (n46212, n_34206, n_34207);
  and g77147 (n46213, n_34091, n46212);
  and g77148 (n46214, pi0534, n46141);
  not g77149 (n_34208, n46214);
  and g77150 (n46215, pi0239, n_34208);
  not g77151 (n_34209, n46213);
  and g77152 (n46216, n_34209, n46215);
  not g77153 (n_34210, n46216);
  and g77154 (n46217, n_34093, n_34210);
  not g77155 (n_34211, n46217);
  and g77156 (n46218, n_34145, n_34211);
  and g77157 (n46219, pi0534, n46212);
  and g77158 (n46220, n_34091, n46141);
  not g77159 (n_34212, n46220);
  and g77160 (n46221, n_906, n_34212);
  not g77161 (n_34213, n46219);
  and g77162 (n46222, n_34213, n46221);
  not g77163 (n_34214, n46222);
  and g77164 (n46223, n_34094, n_34214);
  not g77165 (n_34215, n46223);
  and g77166 (n46224, pi0488, n_34215);
  not g77167 (n_34216, n46218);
  not g77168 (n_34217, n46224);
  and g77169 (n46225, n_34216, n_34217);
  and g77170 (n46226, n_34096, n46225);
  and g77171 (n46227, pi0504, n46145);
  not g77172 (n_34218, n46227);
  and g77173 (n46228, n_2915, n_34218);
  not g77174 (n_34219, n46226);
  and g77175 (n46229, n_34219, n46228);
  not g77176 (n_34220, n46229);
  and g77177 (n46230, n_34098, n_34220);
  not g77178 (n_34221, n46230);
  and g77179 (n46231, n_34149, n_34221);
  and g77180 (n46232, pi0504, n46225);
  and g77181 (n46233, n_34096, n46145);
  not g77182 (n_34222, n46233);
  and g77183 (n46234, pi0242, n_34222);
  not g77184 (n_34223, n46232);
  and g77185 (n46235, n_34223, n46234);
  not g77186 (n_34224, n46235);
  and g77187 (n46236, n_34099, n_34224);
  not g77188 (n_34225, n46236);
  and g77189 (n46237, pi0510, n_34225);
  not g77190 (n_34226, n46231);
  not g77191 (n_34227, n46237);
  and g77192 (n46238, n_34226, n_34227);
  and g77193 (n46239, n_34101, n46238);
  and g77194 (n46240, pi0533, n46149);
  not g77195 (n_34228, n46240);
  and g77196 (n46241, n_1106, n_34228);
  not g77197 (n_34229, n46239);
  and g77198 (n46242, n_34229, n46241);
  not g77199 (n_34230, n46242);
  and g77200 (n46243, n_34103, n_34230);
  not g77201 (n_34231, n46243);
  and g77202 (n46244, n_34153, n_34231);
  and g77203 (n46245, pi0533, n46238);
  and g77204 (n46246, n_34101, n46149);
  not g77205 (n_34232, n46246);
  and g77206 (n46247, pi0235, n_34232);
  not g77207 (n_34233, n46245);
  and g77208 (n46248, n_34233, n46247);
  not g77209 (n_34234, n46248);
  and g77210 (n46249, n_34104, n_34234);
  not g77211 (n_34235, n46249);
  and g77212 (n46250, pi0512, n_34235);
  not g77213 (n_34236, n46244);
  not g77214 (n_34237, n46250);
  and g77215 (n46251, n_34236, n_34237);
  and g77216 (n46252, n_34106, n46251);
  and g77217 (n46253, pi0558, n46153);
  not g77218 (n_34238, n46253);
  and g77219 (n46254, n_2688, n_34238);
  not g77220 (n_34239, n46252);
  and g77221 (n46255, n_34239, n46254);
  not g77222 (n_34240, n46255);
  and g77223 (n46256, n_34108, n_34240);
  not g77224 (n_34241, n46256);
  and g77225 (n46257, n_34157, n_34241);
  and g77226 (n46258, pi0558, n46251);
  and g77227 (n46259, n_34106, n46153);
  not g77228 (n_34242, n46259);
  and g77229 (n46260, pi0244, n_34242);
  not g77230 (n_34243, n46258);
  and g77231 (n46261, n_34243, n46260);
  not g77232 (n_34244, n46261);
  and g77233 (n46262, n_34109, n_34244);
  not g77234 (n_34245, n46262);
  and g77235 (n46263, pi0513, n_34245);
  not g77236 (n_34246, n46257);
  not g77237 (n_34247, n46263);
  and g77238 (n46264, n_34246, n_34247);
  and g77239 (n46265, n_34111, n46264);
  and g77240 (n46266, pi0509, n46157);
  not g77241 (n_34248, n46266);
  and g77242 (n46267, n_2498, n_34248);
  not g77243 (n_34249, n46265);
  and g77244 (n46268, n_34249, n46267);
  not g77245 (n_34250, n46268);
  and g77246 (n46269, n_34113, n_34250);
  not g77247 (n_34251, n46269);
  and g77248 (n46270, n_34161, n_34251);
  and g77249 (n46271, pi0509, n46264);
  and g77250 (n46272, n_34111, n46157);
  not g77251 (n_34252, n46272);
  and g77252 (n46273, pi0245, n_34252);
  not g77253 (n_34253, n46271);
  and g77254 (n46274, n_34253, n46273);
  not g77255 (n_34254, n46274);
  and g77256 (n46275, n_34114, n_34254);
  not g77257 (n_34255, n46275);
  and g77258 (n46276, pi0514, n_34255);
  not g77259 (n_34256, n46270);
  not g77260 (n_34257, n46276);
  and g77261 (n46277, n_34256, n_34257);
  and g77262 (n46278, n_34116, n46277);
  and g77263 (n46279, pi0508, n46161);
  not g77264 (n_34258, n46279);
  and g77265 (n46280, n_1955, n_34258);
  not g77266 (n_34259, n46278);
  and g77267 (n46281, n_34259, n46280);
  not g77268 (n_34260, n46281);
  and g77269 (n46282, n_34118, n_34260);
  not g77270 (n_34261, n46282);
  and g77271 (n46283, n_34165, n_34261);
  and g77272 (n46284, pi0508, n46277);
  and g77273 (n46285, n_34116, n46161);
  not g77274 (n_34262, n46285);
  and g77275 (n46286, pi0247, n_34262);
  not g77276 (n_34263, n46284);
  and g77277 (n46287, n_34263, n46286);
  not g77278 (n_34264, n46287);
  and g77279 (n46288, n_34119, n_34264);
  not g77280 (n_34265, n46288);
  and g77281 (n46289, pi0516, n_34265);
  not g77282 (n_34266, n46283);
  not g77283 (n_34267, n46289);
  and g77284 (n46290, n_34266, n_34267);
  and g77285 (n46291, n_1226, n46290);
  not g77286 (n_34268, pi0517);
  not g77287 (n_34269, n46291);
  and g77288 (n46292, n_34268, n_34269);
  not g77289 (n_34270, pi0507);
  not g77290 (n_34271, n46168);
  and g77291 (n46293, n_34270, n_34271);
  not g77292 (n_34272, n46292);
  and g77293 (n46294, n_34272, n46293);
  and g77294 (n46295, pi0238, n46115);
  and g77295 (n46296, n_1226, n46165);
  not g77296 (n_34273, n46296);
  and g77297 (n46297, n_34268, n_34273);
  not g77298 (n_34274, n46295);
  and g77299 (n46298, n_34274, n46297);
  and g77300 (n46299, pi0238, n46290);
  not g77301 (n_34275, n46299);
  and g77302 (n46300, pi0517, n_34275);
  not g77303 (n_34276, n46298);
  and g77304 (n46301, pi0507, n_34276);
  not g77305 (n_34277, n46300);
  and g77306 (n46302, n_34277, n46301);
  not g77307 (n_34278, n46294);
  not g77308 (n_34279, n46302);
  and g77309 (n46303, n_34278, n_34279);
  not g77310 (n_34280, n46303);
  and g77311 (n46304, pi0233, n_34280);
  not g77312 (n_34281, n46060);
  and g77313 (n46305, pi0237, n_34281);
  not g77314 (n_34282, n46304);
  and g77315 (n46306, n_34282, n46305);
  not g77316 (n_34283, pi0492);
  and g77317 (n46307, n_2307, n_34283);
  and g77318 (n46308, pi0240, pi0492);
  not g77319 (n_34284, n46307);
  not g77320 (n_34285, n46308);
  and g77321 (n46309, n_34284, n_34285);
  and g77322 (n46310, pi0241, pi0490);
  not g77323 (n_34286, pi0490);
  and g77324 (n46311, n_1595, n_34286);
  not g77325 (n_34287, n46310);
  not g77326 (n_34288, n46311);
  and g77327 (n46312, n_34287, n_34288);
  and g77328 (n46313, pi0248, pi0548);
  not g77329 (n_34289, pi0548);
  and g77330 (n46314, n_1774, n_34289);
  not g77331 (n_34290, n46313);
  not g77332 (n_34291, n46314);
  and g77333 (n46315, n_34290, n_34291);
  and g77334 (n46316, pi0249, pi0484);
  not g77335 (n_34292, pi0484);
  and g77336 (n46317, n_1415, n_34292);
  not g77337 (n_34293, n46316);
  not g77338 (n_34294, n46317);
  and g77339 (n46318, n_34293, n_34294);
  and g77340 (n46319, pi0246, pi0546);
  not g77341 (n_34295, pi0546);
  and g77342 (n46320, n_2128, n_34295);
  not g77343 (n_34296, n46319);
  not g77344 (n_34297, n46320);
  and g77345 (n46321, n_34296, n_34297);
  and g77346 (n46322, n_33722, n_33931);
  and g77347 (n46323, pi0544, n_33930);
  not g77357 (n_34303, n46312);
  and g77358 (n46328, n_34303, n46327);
  not g77359 (n_34304, n46309);
  and g77360 (n46329, n_34304, n46328);
  and g77361 (n46330, pi0494, n46329);
  not g77362 (n_34305, n46330);
  and g77363 (n46331, n_906, n_34305);
  not g77364 (n_34306, pi0494);
  and g77365 (n46332, n_34306, n46329);
  not g77366 (n_34307, n46332);
  and g77367 (n46333, pi0239, n_34307);
  not g77368 (n_34308, n46331);
  not g77369 (n_34309, n46333);
  and g77370 (n46334, n_34308, n_34309);
  and g77371 (n46335, pi0483, n46334);
  not g77372 (n_34310, n46335);
  and g77373 (n46336, pi0242, n_34310);
  not g77374 (n_34311, pi0483);
  and g77375 (n46337, n_34311, n46334);
  not g77376 (n_34312, n46337);
  and g77377 (n46338, n_2915, n_34312);
  not g77378 (n_34313, n46336);
  not g77379 (n_34314, n46338);
  and g77380 (n46339, n_34313, n_34314);
  and g77381 (n46340, pi0495, n46339);
  not g77382 (n_34315, n46340);
  and g77383 (n46341, pi0235, n_34315);
  not g77384 (n_34316, pi0495);
  and g77385 (n46342, n_34316, n46339);
  not g77386 (n_34317, n46342);
  and g77387 (n46343, n_1106, n_34317);
  not g77388 (n_34318, n46341);
  not g77389 (n_34319, n46343);
  and g77390 (n46344, n_34318, n_34319);
  and g77391 (n46345, pi0244, pi0493);
  not g77392 (n_34320, pi0493);
  and g77393 (n46346, n_2688, n_34320);
  not g77394 (n_34321, n46345);
  not g77395 (n_34322, n46346);
  and g77396 (n46347, n_34321, n_34322);
  not g77397 (n_34323, n46347);
  and g77398 (n46348, n46344, n_34323);
  and g77399 (n46349, pi0545, n46348);
  not g77400 (n_34324, n46349);
  and g77401 (n46350, pi0245, n_34324);
  not g77402 (n_34325, pi0545);
  and g77403 (n46351, n_34325, n46348);
  not g77404 (n_34326, n46351);
  and g77405 (n46352, n_2498, n_34326);
  not g77406 (n_34327, n46350);
  not g77407 (n_34328, n46352);
  and g77408 (n46353, n_34327, n_34328);
  and g77409 (n46354, pi0547, n46353);
  not g77410 (n_34329, n46354);
  and g77411 (n46355, pi0247, n_34329);
  not g77412 (n_34330, pi0547);
  and g77413 (n46356, n_34330, n46353);
  not g77414 (n_34331, n46356);
  and g77415 (n46357, n_1955, n_34331);
  not g77416 (n_34332, n46355);
  not g77417 (n_34333, n46357);
  and g77418 (n46358, n_34332, n_34333);
  and g77419 (n46359, n_1226, n46358);
  and g77420 (n46360, pi0523, n_33877);
  and g77421 (n46361, pi0248, pi0576);
  not g77422 (n_34334, pi0576);
  and g77423 (n46362, n_1774, n_34334);
  not g77424 (n_34335, n46361);
  not g77425 (n_34336, n46362);
  and g77426 (n46363, n_34335, n_34336);
  and g77427 (n46364, pi0249, pi0528);
  not g77428 (n_34337, pi0528);
  and g77429 (n46365, n_1415, n_34337);
  not g77430 (n_34338, n46364);
  not g77431 (n_34339, n46365);
  and g77432 (n46366, n_34338, n_34339);
  and g77433 (n46367, pi0246, pi0526);
  not g77434 (n_34340, pi0526);
  and g77435 (n46368, n_2128, n_34340);
  not g77436 (n_34341, n46367);
  not g77437 (n_34342, n46368);
  and g77438 (n46369, n_34341, n_34342);
  and g77439 (n46370, n_33695, n_33676);
  and g77449 (n46375, pi0571, n46374);
  not g77450 (n_34348, n46375);
  and g77451 (n46376, pi0241, n_34348);
  not g77452 (n_34349, pi0571);
  and g77453 (n46377, n_34349, n46374);
  not g77454 (n_34350, n46377);
  and g77455 (n46378, n_1595, n_34350);
  not g77456 (n_34351, n46376);
  not g77457 (n_34352, n46378);
  and g77458 (n46379, n_34351, n_34352);
  not g77459 (n_34353, pi0530);
  and g77460 (n46380, n_34353, n46379);
  not g77461 (n_34354, n46380);
  and g77462 (n46381, n_2307, n_34354);
  and g77463 (n46382, pi0530, n46379);
  not g77464 (n_34355, n46382);
  and g77465 (n46383, pi0240, n_34355);
  not g77466 (n_34356, n46381);
  not g77467 (n_34357, n46383);
  and g77468 (n46384, n_34356, n_34357);
  and g77469 (n46385, n_906, pi0524);
  not g77470 (n_34358, pi0524);
  and g77471 (n46386, pi0239, n_34358);
  not g77472 (n_34359, n46385);
  not g77473 (n_34360, n46386);
  and g77474 (n46387, n_34359, n_34360);
  not g77475 (n_34361, n46387);
  and g77476 (n46388, n46384, n_34361);
  and g77477 (n46389, pi0242, pi0573);
  not g77478 (n_34362, pi0573);
  and g77479 (n46390, n_2915, n_34362);
  not g77480 (n_34363, n46389);
  not g77481 (n_34364, n46390);
  and g77482 (n46391, n_34363, n_34364);
  not g77483 (n_34365, n46391);
  and g77484 (n46392, n46388, n_34365);
  and g77485 (n46393, pi0235, pi0575);
  not g77486 (n_34366, pi0575);
  and g77487 (n46394, n_1106, n_34366);
  not g77488 (n_34367, n46393);
  not g77489 (n_34368, n46394);
  and g77490 (n46395, n_34367, n_34368);
  not g77491 (n_34369, n46395);
  and g77492 (n46396, n46392, n_34369);
  and g77493 (n46397, pi0572, n46396);
  not g77494 (n_34370, n46397);
  and g77495 (n46398, pi0244, n_34370);
  not g77496 (n_34371, pi0572);
  and g77497 (n46399, n_34371, n46396);
  not g77498 (n_34372, n46399);
  and g77499 (n46400, n_2688, n_34372);
  not g77500 (n_34373, n46398);
  not g77501 (n_34374, n46400);
  and g77502 (n46401, n_34373, n_34374);
  and g77503 (n46402, pi0245, pi0525);
  not g77504 (n_34375, pi0525);
  and g77505 (n46403, n_2498, n_34375);
  not g77506 (n_34376, n46402);
  not g77507 (n_34377, n46403);
  and g77508 (n46404, n_34376, n_34377);
  not g77509 (n_34378, n46404);
  and g77510 (n46405, n46401, n_34378);
  and g77511 (n46406, pi0247, pi0527);
  not g77512 (n_34379, pi0527);
  and g77513 (n46407, n_1955, n_34379);
  not g77514 (n_34380, n46406);
  not g77515 (n_34381, n46407);
  and g77516 (n46408, n_34380, n_34381);
  not g77517 (n_34382, n46408);
  and g77518 (n46409, n46405, n_34382);
  and g77519 (n46410, pi0238, n46409);
  not g77520 (n_34383, n46410);
  and g77521 (n46411, pi0529, n_34383);
  not g77522 (n_34384, n46359);
  and g77523 (n46412, n_34384, n46411);
  and g77524 (n46413, n_34284, n_34356);
  not g77525 (n_34385, n46328);
  and g77526 (n46414, pi0530, n_34385);
  not g77527 (n_34386, n46327);
  and g77528 (n46415, n_1595, n_34386);
  and g77529 (n46416, n_34350, n46415);
  not g77530 (n_34387, n46416);
  and g77531 (n46417, n_34351, n_34387);
  not g77532 (n_34388, n46417);
  and g77533 (n46418, n_34286, n_34388);
  and g77534 (n46419, pi0241, n_34386);
  and g77535 (n46420, n_34348, n46419);
  not g77536 (n_34389, n46420);
  and g77537 (n46421, n_34352, n_34389);
  not g77538 (n_34390, n46421);
  and g77539 (n46422, pi0490, n_34390);
  not g77540 (n_34391, n46418);
  not g77541 (n_34392, n46422);
  and g77542 (n46423, n_34391, n_34392);
  not g77543 (n_34393, n46423);
  and g77544 (n46424, n_34353, n_34393);
  not g77545 (n_34394, n46414);
  and g77546 (n46425, n_34283, n_34394);
  not g77547 (n_34395, n46424);
  and g77548 (n46426, n_34395, n46425);
  not g77549 (n_34396, n46413);
  not g77550 (n_34397, n46426);
  and g77551 (n46427, n_34396, n_34397);
  and g77552 (n46428, n_34285, n_34357);
  and g77553 (n46429, n_34353, n_34385);
  and g77554 (n46430, pi0530, n_34393);
  not g77555 (n_34398, n46429);
  and g77556 (n46431, pi0492, n_34398);
  not g77557 (n_34399, n46430);
  and g77558 (n46432, n_34399, n46431);
  not g77559 (n_34400, n46428);
  not g77560 (n_34401, n46432);
  and g77561 (n46433, n_34400, n_34401);
  not g77562 (n_34402, n46427);
  not g77563 (n_34403, n46433);
  and g77564 (n46434, n_34402, n_34403);
  and g77565 (n46435, n_34306, n46434);
  and g77566 (n46436, pi0494, n46384);
  not g77567 (n_34404, n46436);
  and g77568 (n46437, pi0239, n_34404);
  not g77569 (n_34405, n46435);
  and g77570 (n46438, n_34405, n46437);
  not g77571 (n_34406, n46438);
  and g77572 (n46439, n_34308, n_34406);
  not g77573 (n_34407, n46439);
  and g77574 (n46440, n_34358, n_34407);
  and g77575 (n46441, pi0494, n46434);
  and g77576 (n46442, n_34306, n46384);
  not g77577 (n_34408, n46442);
  and g77578 (n46443, n_906, n_34408);
  not g77579 (n_34409, n46441);
  and g77580 (n46444, n_34409, n46443);
  not g77581 (n_34410, n46444);
  and g77582 (n46445, n_34309, n_34410);
  not g77583 (n_34411, n46445);
  and g77584 (n46446, pi0524, n_34411);
  not g77585 (n_34412, n46440);
  not g77586 (n_34413, n46446);
  and g77587 (n46447, n_34412, n_34413);
  and g77588 (n46448, n_34311, n46447);
  and g77589 (n46449, pi0483, n46388);
  not g77590 (n_34414, n46449);
  and g77591 (n46450, n_2915, n_34414);
  not g77592 (n_34415, n46448);
  and g77593 (n46451, n_34415, n46450);
  not g77594 (n_34416, n46451);
  and g77595 (n46452, n_34313, n_34416);
  not g77596 (n_34417, n46452);
  and g77597 (n46453, n_34362, n_34417);
  and g77598 (n46454, pi0483, n46447);
  and g77599 (n46455, n_34311, n46388);
  not g77600 (n_34418, n46455);
  and g77601 (n46456, pi0242, n_34418);
  not g77602 (n_34419, n46454);
  and g77603 (n46457, n_34419, n46456);
  not g77604 (n_34420, n46457);
  and g77605 (n46458, n_34314, n_34420);
  not g77606 (n_34421, n46458);
  and g77607 (n46459, pi0573, n_34421);
  not g77608 (n_34422, n46453);
  not g77609 (n_34423, n46459);
  and g77610 (n46460, n_34422, n_34423);
  and g77611 (n46461, n_34316, n46460);
  and g77612 (n46462, pi0495, n46392);
  not g77613 (n_34424, n46462);
  and g77614 (n46463, n_1106, n_34424);
  not g77615 (n_34425, n46461);
  and g77616 (n46464, n_34425, n46463);
  not g77617 (n_34426, n46464);
  and g77618 (n46465, n_34318, n_34426);
  not g77619 (n_34427, n46465);
  and g77620 (n46466, n_34366, n_34427);
  and g77621 (n46467, pi0495, n46460);
  and g77622 (n46468, n_34316, n46392);
  not g77623 (n_34428, n46468);
  and g77624 (n46469, pi0235, n_34428);
  not g77625 (n_34429, n46467);
  and g77626 (n46470, n_34429, n46469);
  not g77627 (n_34430, n46470);
  and g77628 (n46471, n_34319, n_34430);
  not g77629 (n_34431, n46471);
  and g77630 (n46472, pi0575, n_34431);
  not g77631 (n_34432, n46466);
  not g77632 (n_34433, n46472);
  and g77633 (n46473, n_34432, n_34433);
  and g77634 (n46474, n_34371, n46473);
  and g77635 (n46475, pi0572, n46344);
  not g77636 (n_34434, n46475);
  and g77637 (n46476, n_2688, n_34434);
  not g77638 (n_34435, n46474);
  and g77639 (n46477, n_34435, n46476);
  not g77640 (n_34436, n46477);
  and g77641 (n46478, n_34373, n_34436);
  not g77642 (n_34437, n46478);
  and g77643 (n46479, n_34320, n_34437);
  and g77644 (n46480, pi0572, n46473);
  and g77645 (n46481, n_34371, n46344);
  not g77646 (n_34438, n46481);
  and g77647 (n46482, pi0244, n_34438);
  not g77648 (n_34439, n46480);
  and g77649 (n46483, n_34439, n46482);
  not g77650 (n_34440, n46483);
  and g77651 (n46484, n_34374, n_34440);
  not g77652 (n_34441, n46484);
  and g77653 (n46485, pi0493, n_34441);
  not g77654 (n_34442, n46479);
  not g77655 (n_34443, n46485);
  and g77656 (n46486, n_34442, n_34443);
  and g77657 (n46487, n_34325, n46486);
  and g77658 (n46488, pi0545, n46401);
  not g77659 (n_34444, n46488);
  and g77660 (n46489, n_2498, n_34444);
  not g77661 (n_34445, n46487);
  and g77662 (n46490, n_34445, n46489);
  not g77663 (n_34446, n46490);
  and g77664 (n46491, n_34327, n_34446);
  not g77665 (n_34447, n46491);
  and g77666 (n46492, n_34375, n_34447);
  and g77667 (n46493, pi0545, n46486);
  and g77668 (n46494, n_34325, n46401);
  not g77669 (n_34448, n46494);
  and g77670 (n46495, pi0245, n_34448);
  not g77671 (n_34449, n46493);
  and g77672 (n46496, n_34449, n46495);
  not g77673 (n_34450, n46496);
  and g77674 (n46497, n_34328, n_34450);
  not g77675 (n_34451, n46497);
  and g77676 (n46498, pi0525, n_34451);
  not g77677 (n_34452, n46492);
  not g77678 (n_34453, n46498);
  and g77679 (n46499, n_34452, n_34453);
  and g77680 (n46500, n_34330, n46499);
  and g77681 (n46501, pi0547, n46405);
  not g77682 (n_34454, n46501);
  and g77683 (n46502, n_1955, n_34454);
  not g77684 (n_34455, n46500);
  and g77685 (n46503, n_34455, n46502);
  not g77686 (n_34456, n46503);
  and g77687 (n46504, n_34332, n_34456);
  not g77688 (n_34457, n46504);
  and g77689 (n46505, n_34379, n_34457);
  and g77690 (n46506, pi0547, n46499);
  and g77691 (n46507, n_34330, n46405);
  not g77692 (n_34458, n46507);
  and g77693 (n46508, pi0247, n_34458);
  not g77694 (n_34459, n46506);
  and g77695 (n46509, n_34459, n46508);
  not g77696 (n_34460, n46509);
  and g77697 (n46510, n_34333, n_34460);
  not g77698 (n_34461, n46510);
  and g77699 (n46511, pi0527, n_34461);
  not g77700 (n_34462, n46505);
  not g77701 (n_34463, n46511);
  and g77702 (n46512, n_34462, n_34463);
  and g77703 (n46513, n_1226, n46512);
  not g77704 (n_34464, pi0529);
  not g77705 (n_34465, n46513);
  and g77706 (n46514, n_34464, n_34465);
  not g77707 (n_34466, pi0491);
  not g77708 (n_34467, n46412);
  and g77709 (n46515, n_34466, n_34467);
  not g77710 (n_34468, n46514);
  and g77711 (n46516, n_34468, n46515);
  and g77712 (n46517, pi0238, n46358);
  and g77713 (n46518, n_1226, n46409);
  not g77714 (n_34469, n46518);
  and g77715 (n46519, n_34464, n_34469);
  not g77716 (n_34470, n46517);
  and g77717 (n46520, n_34470, n46519);
  and g77718 (n46521, pi0238, n46512);
  not g77719 (n_34471, n46521);
  and g77720 (n46522, pi0529, n_34471);
  not g77721 (n_34472, n46520);
  and g77722 (n46523, pi0491, n_34472);
  not g77723 (n_34473, n46522);
  and g77724 (n46524, n_34473, n46523);
  not g77725 (n_34474, n46516);
  not g77726 (n_34475, n46524);
  and g77727 (n46525, n_34474, n_34475);
  not g77728 (n_34476, n46525);
  and g77729 (n46526, pi0233, n_34476);
  and g77730 (n46527, pi0485, n_33930);
  and g77731 (n46528, pi0240, pi0551);
  not g77732 (n_34477, pi0551);
  and g77733 (n46529, n_2307, n_34477);
  not g77734 (n_34478, n46528);
  not g77735 (n_34479, n46529);
  and g77736 (n46530, n_34478, n_34479);
  not g77737 (n_34480, pi0555);
  and g77738 (n46531, pi0249, n_34480);
  and g77739 (n46532, n_1415, pi0555);
  not g77740 (n_34481, pi0553);
  and g77741 (n46533, pi0241, n_34481);
  and g77742 (n46534, n_1595, pi0553);
  not g77743 (n_34482, pi0554);
  and g77744 (n46535, pi0248, n_34482);
  and g77745 (n46536, n_1774, pi0554);
  and g77746 (n46537, n_2128, pi0563);
  not g77747 (n_34483, pi0563);
  and g77748 (n46538, pi0246, n_34483);
  not g77749 (n_34484, pi0485);
  and g77750 (n46539, n_34484, n_33931);
  and g77772 (n46550, pi0550, n46549);
  not g77773 (n_34496, n46550);
  and g77774 (n46551, n_906, n_34496);
  not g77775 (n_34497, pi0550);
  and g77776 (n46552, n_34497, n46549);
  not g77777 (n_34498, n46552);
  and g77778 (n46553, pi0239, n_34498);
  not g77779 (n_34499, n46551);
  not g77780 (n_34500, n46553);
  and g77781 (n46554, n_34499, n_34500);
  not g77782 (n_34501, pi0489);
  and g77783 (n46555, n_34501, n46554);
  not g77784 (n_34502, n46555);
  and g77785 (n46556, n_2915, n_34502);
  and g77786 (n46557, pi0489, n46554);
  not g77787 (n_34503, n46557);
  and g77788 (n46558, pi0242, n_34503);
  not g77789 (n_34504, n46556);
  not g77790 (n_34505, n46558);
  and g77791 (n46559, n_34504, n_34505);
  and g77792 (n46560, pi0549, n46559);
  not g77793 (n_34506, n46560);
  and g77794 (n46561, pi0235, n_34506);
  not g77795 (n_34507, pi0549);
  and g77796 (n46562, n_34507, n46559);
  not g77797 (n_34508, n46562);
  and g77798 (n46563, n_1106, n_34508);
  not g77799 (n_34509, n46561);
  not g77800 (n_34510, n46563);
  and g77801 (n46564, n_34509, n_34510);
  and g77802 (n46565, pi0486, n46564);
  not g77803 (n_34511, n46565);
  and g77804 (n46566, pi0244, n_34511);
  not g77805 (n_34512, pi0486);
  and g77806 (n46567, n_34512, n46564);
  not g77807 (n_34513, n46567);
  and g77808 (n46568, n_2688, n_34513);
  not g77809 (n_34514, n46566);
  not g77810 (n_34515, n46568);
  and g77811 (n46569, n_34514, n_34515);
  and g77812 (n46570, pi0245, pi0580);
  not g77813 (n_34516, pi0580);
  and g77814 (n46571, n_2498, n_34516);
  not g77815 (n_34517, n46570);
  not g77816 (n_34518, n46571);
  and g77817 (n46572, n_34517, n_34518);
  not g77818 (n_34519, n46572);
  and g77819 (n46573, n46569, n_34519);
  and g77820 (n46574, pi0552, n46573);
  not g77821 (n_34520, n46574);
  and g77822 (n46575, pi0247, n_34520);
  not g77823 (n_34521, pi0552);
  and g77824 (n46576, n_34521, n46573);
  not g77825 (n_34522, n46576);
  and g77826 (n46577, n_1955, n_34522);
  not g77827 (n_34523, n46575);
  not g77828 (n_34524, n46577);
  and g77829 (n46578, n_34523, n_34524);
  and g77830 (n46579, pi0238, n46578);
  not g77831 (n_34525, pi0556);
  and g77832 (n46580, n_2915, n_34525);
  and g77833 (n46581, pi0242, pi0556);
  not g77834 (n_34526, n46580);
  not g77835 (n_34527, n46581);
  and g77836 (n46582, n_34526, n_34527);
  not g77837 (n_34528, pi0564);
  and g77838 (n46583, pi0246, n_34528);
  and g77839 (n46584, pi0570, n_33877);
  and g77840 (n46585, n_2128, pi0564);
  not g77841 (n_34529, pi0482);
  and g77842 (n46586, pi0249, n_34529);
  and g77843 (n46587, n_1415, pi0482);
  and g77844 (n46588, pi0241, pi0562);
  not g77845 (n_34530, pi0562);
  and g77846 (n46589, n_1595, n_34530);
  not g77847 (n_34531, n46588);
  not g77848 (n_34532, n46589);
  and g77849 (n46590, n_34531, n_34532);
  and g77850 (n46591, n_33836, n_33676);
  not g77862 (n_34539, pi0565);
  and g77863 (n46597, pi0248, n_34539);
  and g77864 (n46598, n_1774, pi0565);
  not g77865 (n_34540, n46597);
  not g77866 (n_34541, n46598);
  and g77867 (n46599, n_34540, n_34541);
  and g77868 (n46600, pi0240, pi0560);
  not g77869 (n_34542, pi0560);
  and g77870 (n46601, n_2307, n_34542);
  not g77871 (n_34543, n46600);
  not g77872 (n_34544, n46601);
  and g77873 (n46602, n_34543, n_34544);
  not g77874 (n_34545, n46583);
  not g77879 (n_34547, n46605);
  and g77880 (n46606, n_2307, n_34547);
  not g77884 (n_34548, n46609);
  and g77885 (n46610, pi0240, n_34548);
  not g77886 (n_34549, n46606);
  not g77887 (n_34550, n46610);
  and g77888 (n46611, n_34549, n_34550);
  and g77889 (n46612, n_906, pi0569);
  not g77890 (n_34551, pi0569);
  and g77891 (n46613, pi0239, n_34551);
  not g77892 (n_34552, n46612);
  not g77893 (n_34553, n46613);
  and g77894 (n46614, n_34552, n_34553);
  not g77895 (n_34554, n46614);
  and g77896 (n46615, n46611, n_34554);
  not g77897 (n_34555, n46582);
  and g77898 (n46616, n_34555, n46615);
  and g77899 (n46617, pi0235, pi0531);
  not g77900 (n_34556, pi0531);
  and g77901 (n46618, n_1106, n_34556);
  not g77902 (n_34557, n46617);
  not g77903 (n_34558, n46618);
  and g77904 (n46619, n_34557, n_34558);
  not g77905 (n_34559, n46619);
  and g77906 (n46620, n46616, n_34559);
  and g77907 (n46621, pi0244, pi0566);
  not g77908 (n_34560, pi0566);
  and g77909 (n46622, n_2688, n_34560);
  not g77910 (n_34561, n46621);
  not g77911 (n_34562, n46622);
  and g77912 (n46623, n_34561, n_34562);
  not g77913 (n_34563, n46623);
  and g77914 (n46624, n46620, n_34563);
  and g77915 (n46625, pi0568, n46624);
  not g77916 (n_34564, n46625);
  and g77917 (n46626, pi0245, n_34564);
  not g77918 (n_34565, pi0568);
  and g77919 (n46627, n_34565, n46624);
  not g77920 (n_34566, n46627);
  and g77921 (n46628, n_2498, n_34566);
  not g77922 (n_34567, n46626);
  not g77923 (n_34568, n46628);
  and g77924 (n46629, n_34567, n_34568);
  and g77925 (n46630, pi0247, pi0532);
  not g77926 (n_34569, pi0532);
  and g77927 (n46631, n_1955, n_34569);
  not g77928 (n_34570, n46630);
  not g77929 (n_34571, n46631);
  and g77930 (n46632, n_34570, n_34571);
  not g77931 (n_34572, n46632);
  and g77932 (n46633, n46629, n_34572);
  and g77933 (n46634, n_1226, n46633);
  not g77934 (n_34573, n46634);
  and g77935 (n46635, pi0577, n_34573);
  not g77936 (n_34574, n46579);
  and g77937 (n46636, n_34574, n46635);
  and g77938 (n46637, n_34504, n_34526);
  not g77939 (n_34575, n46615);
  and g77940 (n46638, pi0489, n_34575);
  and g77941 (n46639, n46605, n46613);
  and g77942 (n46640, pi0569, n_34500);
  and g77943 (n46641, n46611, n46640);
  not g77944 (n_34576, n46554);
  not g77945 (n_34577, n46639);
  and g77946 (n46642, n_34576, n_34577);
  not g77947 (n_34578, n46641);
  and g77948 (n46643, n_34578, n46642);
  and g77949 (n46644, n_34501, n46643);
  not g77950 (n_34579, n46638);
  and g77951 (n46645, n_34525, n_34579);
  not g77952 (n_34580, n46644);
  and g77953 (n46646, n_34580, n46645);
  not g77954 (n_34581, n46637);
  not g77955 (n_34582, n46646);
  and g77956 (n46647, n_34581, n_34582);
  and g77957 (n46648, n_34505, n_34527);
  and g77958 (n46649, n_34501, n_34575);
  and g77959 (n46650, pi0489, n46643);
  not g77960 (n_34583, n46649);
  and g77961 (n46651, pi0556, n_34583);
  not g77962 (n_34584, n46650);
  and g77963 (n46652, n_34584, n46651);
  not g77964 (n_34585, n46648);
  not g77965 (n_34586, n46652);
  and g77966 (n46653, n_34585, n_34586);
  not g77967 (n_34587, n46647);
  not g77968 (n_34588, n46653);
  and g77969 (n46654, n_34587, n_34588);
  and g77970 (n46655, n_34507, n46654);
  and g77971 (n46656, pi0549, n46616);
  not g77972 (n_34589, n46656);
  and g77973 (n46657, n_1106, n_34589);
  not g77974 (n_34590, n46655);
  and g77975 (n46658, n_34590, n46657);
  not g77976 (n_34591, n46658);
  and g77977 (n46659, n_34509, n_34591);
  not g77978 (n_34592, n46659);
  and g77979 (n46660, n_34556, n_34592);
  and g77980 (n46661, pi0549, n46654);
  and g77981 (n46662, n_34507, n46616);
  not g77982 (n_34593, n46662);
  and g77983 (n46663, pi0235, n_34593);
  not g77984 (n_34594, n46661);
  and g77985 (n46664, n_34594, n46663);
  not g77986 (n_34595, n46664);
  and g77987 (n46665, n_34510, n_34595);
  not g77988 (n_34596, n46665);
  and g77989 (n46666, pi0531, n_34596);
  not g77990 (n_34597, n46660);
  not g77991 (n_34598, n46666);
  and g77992 (n46667, n_34597, n_34598);
  and g77993 (n46668, n_34512, n46667);
  and g77994 (n46669, pi0486, n46620);
  not g77995 (n_34599, n46669);
  and g77996 (n46670, n_2688, n_34599);
  not g77997 (n_34600, n46668);
  and g77998 (n46671, n_34600, n46670);
  not g77999 (n_34601, n46671);
  and g78000 (n46672, n_34514, n_34601);
  not g78001 (n_34602, n46672);
  and g78002 (n46673, n_34560, n_34602);
  and g78003 (n46674, pi0486, n46667);
  and g78004 (n46675, n_34512, n46620);
  not g78005 (n_34603, n46675);
  and g78006 (n46676, pi0244, n_34603);
  not g78007 (n_34604, n46674);
  and g78008 (n46677, n_34604, n46676);
  not g78009 (n_34605, n46677);
  and g78010 (n46678, n_34515, n_34605);
  not g78011 (n_34606, n46678);
  and g78012 (n46679, pi0566, n_34606);
  not g78013 (n_34607, n46673);
  not g78014 (n_34608, n46679);
  and g78015 (n46680, n_34607, n_34608);
  and g78016 (n46681, n_34565, n46680);
  and g78017 (n46682, pi0568, n46569);
  not g78018 (n_34609, n46682);
  and g78019 (n46683, n_2498, n_34609);
  not g78020 (n_34610, n46681);
  and g78021 (n46684, n_34610, n46683);
  not g78022 (n_34611, n46684);
  and g78023 (n46685, n_34567, n_34611);
  not g78024 (n_34612, n46685);
  and g78025 (n46686, n_34516, n_34612);
  and g78026 (n46687, pi0568, n46680);
  and g78027 (n46688, n_34565, n46569);
  not g78028 (n_34613, n46688);
  and g78029 (n46689, pi0245, n_34613);
  not g78030 (n_34614, n46687);
  and g78031 (n46690, n_34614, n46689);
  not g78032 (n_34615, n46690);
  and g78033 (n46691, n_34568, n_34615);
  not g78034 (n_34616, n46691);
  and g78035 (n46692, pi0580, n_34616);
  not g78036 (n_34617, n46686);
  not g78037 (n_34618, n46692);
  and g78038 (n46693, n_34617, n_34618);
  and g78039 (n46694, n_34521, n46693);
  and g78040 (n46695, pi0552, n46629);
  not g78041 (n_34619, n46695);
  and g78042 (n46696, n_1955, n_34619);
  not g78043 (n_34620, n46694);
  and g78044 (n46697, n_34620, n46696);
  not g78045 (n_34621, n46697);
  and g78046 (n46698, n_34523, n_34621);
  not g78047 (n_34622, n46698);
  and g78048 (n46699, n_34569, n_34622);
  and g78049 (n46700, pi0552, n46693);
  and g78050 (n46701, n_34521, n46629);
  not g78051 (n_34623, n46701);
  and g78052 (n46702, pi0247, n_34623);
  not g78053 (n_34624, n46700);
  and g78054 (n46703, n_34624, n46702);
  not g78055 (n_34625, n46703);
  and g78056 (n46704, n_34524, n_34625);
  not g78057 (n_34626, n46704);
  and g78058 (n46705, pi0532, n_34626);
  not g78059 (n_34627, n46699);
  not g78060 (n_34628, n46705);
  and g78061 (n46706, n_34627, n_34628);
  and g78062 (n46707, n_1226, n46706);
  not g78063 (n_34629, pi0577);
  not g78064 (n_34630, n46707);
  and g78065 (n46708, n_34629, n_34630);
  not g78066 (n_34631, pi0498);
  not g78067 (n_34632, n46636);
  and g78068 (n46709, n_34631, n_34632);
  not g78069 (n_34633, n46708);
  and g78070 (n46710, n_34633, n46709);
  and g78071 (n46711, n_1226, n46578);
  and g78072 (n46712, pi0238, n46633);
  not g78073 (n_34634, n46712);
  and g78074 (n46713, n_34629, n_34634);
  not g78075 (n_34635, n46711);
  and g78076 (n46714, n_34635, n46713);
  and g78077 (n46715, pi0238, n46706);
  not g78078 (n_34636, n46715);
  and g78079 (n46716, pi0577, n_34636);
  not g78080 (n_34637, n46714);
  and g78081 (n46717, pi0498, n_34637);
  not g78082 (n_34638, n46716);
  and g78083 (n46718, n_34638, n46717);
  not g78084 (n_34639, n46710);
  not g78085 (n_34640, n46718);
  and g78086 (n46719, n_34639, n_34640);
  not g78087 (n_34641, n46719);
  and g78088 (n46720, n_25720, n_34641);
  not g78089 (n_34642, n46720);
  and g78090 (n46721, n_25730, n_34642);
  not g78091 (n_34643, n46526);
  and g78092 (n46722, n_34643, n46721);
  not g78093 (n_34644, n46306);
  not g78094 (n_34645, n46722);
  and g78095 (po0750, n_34644, n_34645);
  not g78096 (n_34647, pi0806);
  and g78097 (n46724, n_34647, n45126);
  and g78098 (n46725, n_4, n_34647);
  and g78099 (n46726, pi0990, n46725);
  and g78100 (n46727, pi0600, n46726);
  and g78101 (n46728, n_4, pi0594);
  not g78102 (n_34648, n46727);
  not g78103 (n_34649, n46728);
  and g78104 (n46729, n_34648, n_34649);
  not g78105 (n_34650, n46724);
  not g78106 (n_34651, n46729);
  and g78107 (po0751, n_34650, n_34651);
  and g78108 (n46731, pi0605, n_34647);
  and g78109 (n46732, n45109, n46731);
  not g78110 (n_34652, n46732);
  and g78111 (n46733, n_33450, n_34652);
  and g78112 (n46734, pi0595, n46732);
  not g78113 (n_34653, n46733);
  and g78114 (n46735, n_4, n_34653);
  not g78115 (n_34654, n46734);
  and g78116 (po0752, n_34654, n46735);
  and g78117 (n46737, n_4, pi0596);
  and g78118 (n46738, pi0595, n45108);
  and g78119 (n46739, n46726, n46738);
  not g78120 (n_34655, n46737);
  not g78121 (n_34656, n46739);
  and g78122 (n46740, n_34655, n_34656);
  and g78123 (n46741, pi0596, n46739);
  not g78124 (n_34657, n46740);
  not g78125 (n_34658, n46741);
  and g78126 (po0753, n_34657, n_34658);
  not g78127 (n_34659, pi0597);
  and g78128 (n46743, n_34659, n_34650);
  and g78129 (n46744, pi0597, n46724);
  not g78130 (n_34660, n46743);
  and g78131 (n46745, n_4, n_34660);
  not g78132 (n_34661, n46744);
  and g78133 (po0754, n_34661, n46745);
  not g78134 (n_34663, pi0882);
  and g78135 (n46747, n_34663, n_4226);
  and g78136 (n46748, pi0947, n46747);
  not g78137 (n_34665, n46748);
  and g78138 (n46749, pi0598, n_34665);
  and g78139 (n46750, pi0740, pi0780);
  and g78140 (n46751, n6192, n46750);
  or g78141 (po0755, n46749, n46751);
  and g78142 (n46753, n_4, pi0599);
  not g78143 (n_34668, n46753);
  and g78144 (n46754, n_34658, n_34668);
  and g78145 (n46755, pi0599, n46741);
  not g78146 (n_34669, n46754);
  not g78147 (n_34670, n46755);
  and g78148 (po0756, n_34669, n_34670);
  and g78149 (n46757, n_4, pi0600);
  not g78150 (n_34671, n46726);
  not g78151 (n_34672, n46757);
  and g78152 (n46758, n_34671, n_34672);
  not g78153 (n_34673, n46758);
  and g78154 (po0757, n_34648, n_34673);
  not g78155 (n_34675, pi0989);
  and g78156 (n46760, n_34647, n_34675);
  and g78157 (n46761, n_33462, pi0806);
  not g78158 (n_34676, n46760);
  and g78159 (n46762, n_4, n_34676);
  not g78160 (n_34677, n46761);
  and g78161 (po0758, n_34677, n46762);
  and g78162 (n46764, n_28510, pi0602);
  and g78163 (n46765, n_12395, n_12405);
  and g78164 (n46766, pi0715, pi1160);
  not g78165 (n_34678, n46765);
  and g78166 (n46767, pi0790, n_34678);
  not g78167 (n_34679, n46766);
  and g78168 (n46768, n_34679, n46767);
  or g78177 (po0759, n46764, n46774);
  and g78178 (n46776, pi0871, pi0966);
  and g78179 (n46777, pi0872, pi0966);
  not g78180 (n_34686, pi1100);
  and g78181 (n46778, pi0832, n_34686);
  not g78182 (n_34688, pi0980);
  and g78183 (n46779, n_34688, pi1038);
  and g78184 (n46780, pi1060, n46779);
  not g78185 (n_34693, pi1061);
  and g78186 (n46781, pi0952, n_34693);
  and g78187 (n46782, n46780, n46781);
  and g78188 (n46783, n46778, n46782);
  and g78189 (po0897, pi0832, n46782);
  not g78190 (n_34695, po0897);
  and g78191 (n46785, n_11512, n_34695);
  not g78192 (n_34696, pi0966);
  not g78193 (n_34697, n46783);
  and g78194 (n46786, n_34696, n_34697);
  not g78195 (n_34698, n46785);
  and g78196 (n46787, n_34698, n46786);
  not g78197 (n_34699, n46776);
  not g78198 (n_34700, n46777);
  and g78199 (n46788, n_34699, n_34700);
  not g78200 (n_34701, n46788);
  or g78201 (po0760, n46787, n_34701);
  and g78202 (n46790, pi0823, n16657);
  not g78203 (n_34704, pi0779);
  and g78204 (n46791, n_34704, n46790);
  and g78205 (n46792, n_234, pi0983);
  and g78206 (n46793, pi0907, n46792);
  not g78207 (n_34707, n46793);
  and g78208 (n46794, pi0604, n_34707);
  not g78209 (n_34708, n46790);
  and g78210 (n46795, n_34708, n46794);
  or g78211 (po0761, n46791, n46795);
  not g78212 (n_34709, pi0605);
  not g78213 (n_34710, n46725);
  and g78214 (n46797, n_34709, n_34710);
  not g78215 (n_34711, n46731);
  and g78216 (n46798, n_4, n_34711);
  not g78217 (n_34712, n46797);
  and g78218 (po0762, n_34712, n46798);
  and g78219 (n46800, n_25343, n_34695);
  not g78220 (n_34714, pi1104);
  and g78221 (n46801, n_34714, po0897);
  not g78222 (n_34715, n46800);
  not g78223 (n_34716, n46801);
  and g78224 (n46802, n_34715, n_34716);
  not g78225 (n_34717, n46802);
  and g78226 (n46803, n_34696, n_34717);
  not g78227 (n_34719, pi0837);
  and g78228 (n46804, n_34719, pi0966);
  not g78229 (n_34720, n46803);
  not g78230 (n_34721, n46804);
  and g78231 (po0763, n_34720, n_34721);
  and g78232 (n46806, n_26264, n_34695);
  not g78233 (n_34723, pi1107);
  and g78234 (n46807, n_34723, po0897);
  not g78235 (n_34724, n46806);
  and g78236 (n46808, n_34696, n_34724);
  not g78237 (n_34725, n46807);
  and g78238 (po0764, n_34725, n46808);
  and g78239 (n46810, n_11823, n_34695);
  not g78240 (n_34727, pi1116);
  and g78241 (n46811, n_34727, po0897);
  not g78242 (n_34728, n46810);
  and g78243 (n46812, n_34696, n_34728);
  not g78244 (n_34729, n46811);
  and g78245 (po0765, n_34729, n46812);
  and g78246 (n46814, n_11971, n_34695);
  not g78247 (n_34731, pi1118);
  and g78248 (n46815, n_34731, po0897);
  not g78249 (n_34732, n46814);
  and g78250 (n46816, n_34696, n_34732);
  not g78251 (n_34733, n46815);
  and g78252 (po0766, n_34733, n46816);
  not g78253 (n_34735, pi0610);
  and g78254 (n46818, n_34735, n_34695);
  not g78255 (n_34737, pi1113);
  and g78256 (n46819, n_34737, po0897);
  not g78257 (n_34738, n46818);
  and g78258 (n46820, n_34696, n_34738);
  not g78259 (n_34739, n46819);
  and g78260 (po0767, n_34739, n46820);
  not g78261 (n_34741, pi0611);
  and g78262 (n46822, n_34741, n_34695);
  not g78263 (n_34743, pi1114);
  and g78264 (n46823, n_34743, po0897);
  not g78265 (n_34744, n46822);
  and g78266 (n46824, n_34696, n_34744);
  not g78267 (n_34745, n46823);
  and g78268 (po0768, n_34745, n46824);
  and g78269 (n46826, n_26742, n_34695);
  not g78270 (n_34747, pi1111);
  and g78271 (n46827, n_34747, po0897);
  not g78272 (n_34748, n46826);
  and g78273 (n46828, n_34696, n_34748);
  not g78274 (n_34749, n46827);
  and g78275 (po0769, n_34749, n46828);
  not g78276 (n_34751, pi0613);
  and g78277 (n46830, n_34751, n_34695);
  not g78278 (n_34753, pi1115);
  and g78279 (n46831, n_34753, po0897);
  not g78280 (n_34754, n46830);
  and g78281 (n46832, n_34696, n_34754);
  not g78282 (n_34755, n46831);
  and g78283 (po0770, n_34755, n46832);
  and g78284 (n46834, n_3090, n_34695);
  not g78285 (n_34757, pi1102);
  and g78286 (n46835, n_34757, po0897);
  not g78287 (n_34758, n46834);
  and g78288 (n46836, n_34696, n_34758);
  not g78289 (n_34759, n46835);
  and g78290 (n46837, n_34759, n46836);
  or g78291 (po0771, n46776, n46837);
  and g78292 (n46839, pi0907, n46747);
  not g78293 (n_34761, pi0615);
  not g78294 (n_34762, n46839);
  and g78295 (n46840, n_34761, n_34762);
  and g78296 (n46841, pi0779, pi0797);
  and g78297 (n46842, n6195, n46841);
  or g78298 (po0772, n46840, n46842);
  and g78299 (n46844, n_3091, n_34695);
  not g78300 (n_34765, pi1101);
  and g78301 (n46845, n_34765, po0897);
  not g78302 (n_34766, n46844);
  and g78303 (n46846, n_34696, n_34766);
  not g78304 (n_34767, n46845);
  and g78305 (n46847, n_34767, n46846);
  or g78306 (po0773, n46777, n46847);
  and g78307 (n46849, n_25117, n_34695);
  not g78308 (n_34769, pi1105);
  and g78309 (n46850, n_34769, po0897);
  not g78310 (n_34770, n46849);
  not g78311 (n_34771, n46850);
  and g78312 (n46851, n_34770, n_34771);
  not g78313 (n_34772, n46851);
  and g78314 (n46852, n_34696, n_34772);
  not g78315 (n_34774, pi0850);
  and g78316 (n46853, n_34774, pi0966);
  not g78317 (n_34775, n46852);
  not g78318 (n_34776, n46853);
  and g78319 (po0774, n_34775, n_34776);
  and g78320 (n46855, n_11984, n_34695);
  not g78321 (n_34778, pi1117);
  and g78322 (n46856, n_34778, po0897);
  not g78323 (n_34779, n46855);
  and g78324 (n46857, n_34696, n_34779);
  not g78325 (n_34780, n46856);
  and g78326 (po0775, n_34780, n46857);
  and g78327 (n46859, n_11821, n_34695);
  not g78328 (n_34782, pi1122);
  and g78329 (n46860, n_34782, po0897);
  not g78330 (n_34783, n46859);
  and g78331 (n46861, n_34696, n_34783);
  not g78332 (n_34784, n46860);
  and g78333 (po0776, n_34784, n46861);
  not g78334 (n_34786, pi0620);
  and g78335 (n46863, n_34786, n_34695);
  not g78336 (n_34788, pi1112);
  and g78337 (n46864, n_34788, po0897);
  not g78338 (n_34789, n46863);
  and g78339 (n46865, n_34696, n_34789);
  not g78340 (n_34790, n46864);
  and g78341 (po0777, n_34790, n46865);
  and g78342 (n46867, n_12038, n_34695);
  not g78343 (n_34792, pi1108);
  and g78344 (n46868, n_34792, po0897);
  not g78345 (n_34793, n46867);
  and g78346 (n46869, n_34696, n_34793);
  not g78347 (n_34794, n46868);
  and g78348 (po0778, n_34794, n46869);
  and g78349 (n46871, n_26336, n_34695);
  not g78350 (n_34796, pi1109);
  and g78351 (n46872, n_34796, po0897);
  not g78352 (n_34797, n46871);
  and g78353 (n46873, n_34696, n_34797);
  not g78354 (n_34798, n46872);
  and g78355 (po0779, n_34798, n46873);
  and g78356 (n46875, n_25938, n_34695);
  not g78357 (n_34800, pi1106);
  and g78358 (n46876, n_34800, po0897);
  not g78359 (n_34801, n46875);
  and g78360 (n46877, n_34696, n_34801);
  not g78361 (n_34802, n46876);
  and g78362 (po0780, n_34802, n46877);
  and g78363 (n46879, pi0831, n17167);
  not g78364 (n_34804, pi0780);
  and g78365 (n46880, n_34804, n46879);
  and g78366 (n46881, pi0947, n46792);
  not g78367 (n_34806, n46881);
  and g78368 (n46882, pi0624, n_34806);
  not g78369 (n_34807, n46879);
  and g78370 (n46883, n_34807, n46882);
  or g78371 (po0781, n46880, n46883);
  not g78378 (n_34815, pi0953);
  and g78379 (po0954, n_34815, n46888);
  not g78380 (n_34817, po0954);
  and g78381 (n46890, n_11753, n_34817);
  and g78382 (n46891, n_34727, po0954);
  not g78383 (n_34819, pi0962);
  not g78384 (n_34820, n46890);
  and g78385 (n46892, n_34819, n_34820);
  not g78386 (n_34821, n46891);
  and g78387 (po0782, n_34821, n46892);
  and g78388 (n46894, n_12320, n_34695);
  not g78389 (n_34823, pi1121);
  and g78390 (n46895, n_34823, po0897);
  not g78391 (n_34824, n46894);
  and g78392 (n46896, n_34696, n_34824);
  not g78393 (n_34825, n46895);
  and g78394 (po0783, n_34825, n46896);
  and g78395 (n46898, n_11412, n_34817);
  and g78396 (n46899, n_34778, po0954);
  not g78397 (n_34826, n46898);
  and g78398 (n46900, n_34819, n_34826);
  not g78399 (n_34827, n46899);
  and g78400 (po0784, n_34827, n46900);
  and g78401 (n46902, n_11789, n_34817);
  not g78402 (n_34829, pi1119);
  and g78403 (n46903, n_34829, po0954);
  not g78404 (n_34830, n46902);
  and g78405 (n46904, n_34819, n_34830);
  not g78406 (n_34831, n46903);
  and g78407 (po0785, n_34831, n46904);
  and g78408 (n46906, n_12354, n_34695);
  and g78409 (n46907, n_34829, po0897);
  not g78410 (n_34832, n46906);
  and g78411 (n46908, n_34696, n_34832);
  not g78412 (n_34833, n46907);
  and g78413 (po0786, n_34833, n46908);
  and g78414 (n46910, n_12375, n_34695);
  not g78415 (n_34835, pi1120);
  and g78416 (n46911, n_34835, po0897);
  not g78417 (n_34836, n46910);
  and g78418 (n46912, n_34696, n_34836);
  not g78419 (n_34837, n46911);
  and g78420 (po0787, n_34837, n46912);
  and g78421 (n46914, n_34737, po0954);
  and g78422 (n46915, pi0631, n_34817);
  not g78423 (n_34839, n46914);
  and g78424 (n46916, n_34819, n_34839);
  not g78425 (n_34840, n46915);
  and g78426 (po0788, n_34840, n46916);
  and g78427 (n46918, n_34753, po0954);
  and g78428 (n46919, pi0632, n_34817);
  not g78429 (n_34842, n46918);
  and g78430 (n46920, n_34819, n_34842);
  not g78431 (n_34843, n46919);
  and g78432 (po0789, n_34843, n46920);
  and g78433 (n46922, n_24918, n_34695);
  not g78434 (n_34845, pi1110);
  and g78435 (n46923, n_34845, po0897);
  not g78436 (n_34846, n46922);
  and g78437 (n46924, n_34696, n_34846);
  not g78438 (n_34847, n46923);
  and g78439 (po0790, n_34847, n46924);
  and g78440 (n46926, n_24930, n_34817);
  and g78441 (n46927, n_34845, po0954);
  not g78442 (n_34848, n46926);
  and g78443 (n46928, n_34819, n_34848);
  not g78444 (n_34849, n46927);
  and g78445 (po0791, n_34849, n46928);
  and g78446 (n46930, n_34788, po0954);
  and g78447 (n46931, pi0635, n_34817);
  not g78448 (n_34851, n46930);
  and g78449 (n46932, n_34819, n_34851);
  not g78450 (n_34852, n46931);
  and g78451 (po0792, n_34852, n46932);
  not g78452 (n_34854, pi0636);
  and g78453 (n46934, n_34854, n_34695);
  not g78454 (n_34856, pi1127);
  and g78455 (n46935, n_34856, po0897);
  not g78456 (n_34857, n46934);
  and g78457 (n46936, n_34696, n_34857);
  not g78458 (n_34858, n46935);
  and g78459 (po0793, n_34858, n46936);
  and g78460 (n46938, n_25155, n_34817);
  and g78461 (n46939, n_34769, po0954);
  not g78462 (n_34859, n46938);
  and g78463 (n46940, n_34819, n_34859);
  not g78464 (n_34860, n46939);
  and g78465 (po0794, n_34860, n46940);
  and g78466 (n46942, n_26247, n_34817);
  and g78467 (n46943, n_34723, po0954);
  not g78468 (n_34861, n46942);
  and g78469 (n46944, n_34819, n_34861);
  not g78470 (n_34862, n46943);
  and g78471 (po0795, n_34862, n46944);
  and g78472 (n46946, n_26303, n_34817);
  and g78473 (n46947, n_34796, po0954);
  not g78474 (n_34863, n46946);
  and g78475 (n46948, n_34819, n_34863);
  not g78476 (n_34864, n46947);
  and g78477 (po0796, n_34864, n46948);
  not g78478 (n_34866, pi0640);
  and g78479 (n46950, n_34866, n_34695);
  not g78480 (n_34868, pi1128);
  and g78481 (n46951, n_34868, po0897);
  not g78482 (n_34869, n46950);
  and g78483 (n46952, n_34696, n_34869);
  not g78484 (n_34870, n46951);
  and g78485 (po0797, n_34870, n46952);
  and g78486 (n46954, n_11395, n_34817);
  and g78487 (n46955, n_34823, po0954);
  not g78488 (n_34871, n46954);
  and g78489 (n46956, n_34819, n_34871);
  not g78490 (n_34872, n46955);
  and g78491 (po0798, n_34872, n46956);
  and g78492 (n46958, n_3087, n_34695);
  not g78493 (n_34874, pi1103);
  and g78494 (n46959, n_34874, po0897);
  not g78495 (n_34875, n46958);
  and g78496 (n46960, n_34696, n_34875);
  not g78497 (n_34876, n46959);
  and g78498 (po0799, n_34876, n46960);
  and g78499 (n46962, n_25400, n_34817);
  and g78500 (n46963, n_34714, po0954);
  not g78501 (n_34877, n46962);
  and g78502 (n46964, n_34819, n_34877);
  not g78503 (n_34878, n46963);
  and g78504 (po0800, n_34878, n46964);
  and g78505 (n46966, n_11819, n_34695);
  not g78506 (n_34880, pi1123);
  and g78507 (n46967, n_34880, po0897);
  not g78508 (n_34881, n46966);
  and g78509 (n46968, n_34696, n_34881);
  not g78510 (n_34882, n46967);
  and g78511 (po0801, n_34882, n46968);
  not g78512 (n_34884, pi0645);
  and g78513 (n46970, n_34884, n_34695);
  not g78514 (n_34886, pi1125);
  and g78515 (n46971, n_34886, po0897);
  not g78516 (n_34887, n46970);
  and g78517 (n46972, n_34696, n_34887);
  not g78518 (n_34888, n46971);
  and g78519 (po0802, n_34888, n46972);
  and g78520 (n46974, n_34743, po0954);
  and g78521 (n46975, pi0646, n_34817);
  not g78522 (n_34890, n46974);
  and g78523 (n46976, n_34819, n_34890);
  not g78524 (n_34891, n46975);
  and g78525 (po0803, n_34891, n46976);
  and g78526 (n46978, n_11806, n_34817);
  and g78527 (n46979, n_34835, po0954);
  not g78528 (n_34892, n46978);
  and g78529 (n46980, n_34819, n_34892);
  not g78530 (n_34893, n46979);
  and g78531 (po0804, n_34893, n46980);
  and g78532 (n46982, n_11403, n_34817);
  and g78533 (n46983, n_34782, po0954);
  not g78534 (n_34894, n46982);
  and g78535 (n46984, n_34819, n_34894);
  not g78536 (n_34895, n46983);
  and g78537 (po0805, n_34895, n46984);
  not g78538 (n_34897, pi1126);
  and g78539 (n46986, n_34897, po0954);
  and g78540 (n46987, pi0649, n_34817);
  not g78541 (n_34899, n46986);
  and g78542 (n46988, n_34819, n_34899);
  not g78543 (n_34900, n46987);
  and g78544 (po0806, n_34900, n46988);
  and g78545 (n46990, n_34856, po0954);
  and g78546 (n46991, pi0650, n_34817);
  not g78547 (n_34902, n46990);
  and g78548 (n46992, n_34819, n_34902);
  not g78549 (n_34903, n46991);
  and g78550 (po0807, n_34903, n46992);
  not g78551 (n_34905, pi0651);
  and g78552 (n46994, n_34905, n_34695);
  not g78553 (n_34907, pi1130);
  and g78554 (n46995, n_34907, po0897);
  not g78555 (n_34908, n46994);
  and g78556 (n46996, n_34696, n_34908);
  not g78557 (n_34909, n46995);
  and g78558 (po0808, n_34909, n46996);
  not g78559 (n_34911, pi0652);
  and g78560 (n46998, n_34911, n_34695);
  not g78561 (n_34913, pi1131);
  and g78562 (n46999, n_34913, po0897);
  not g78563 (n_34914, n46998);
  and g78564 (n47000, n_34696, n_34914);
  not g78565 (n_34915, n46999);
  and g78566 (po0809, n_34915, n47000);
  not g78567 (n_34917, pi0653);
  and g78568 (n47002, n_34917, n_34695);
  not g78569 (n_34919, pi1129);
  and g78570 (n47003, n_34919, po0897);
  not g78571 (n_34920, n47002);
  and g78572 (n47004, n_34696, n_34920);
  not g78573 (n_34921, n47003);
  and g78574 (po0810, n_34921, n47004);
  and g78575 (n47006, n_34907, po0954);
  and g78576 (n47007, pi0654, n_34817);
  not g78577 (n_34923, n47006);
  and g78578 (n47008, n_34819, n_34923);
  not g78579 (n_34924, n47007);
  and g78580 (po0811, n_34924, n47008);
  not g78581 (n_34926, pi1124);
  and g78582 (n47010, n_34926, po0954);
  and g78583 (n47011, pi0655, n_34817);
  not g78584 (n_34928, n47010);
  and g78585 (n47012, n_34819, n_34928);
  not g78586 (n_34929, n47011);
  and g78587 (po0812, n_34929, n47012);
  not g78588 (n_34931, pi0656);
  and g78589 (n47014, n_34931, n_34695);
  and g78590 (n47015, n_34897, po0897);
  not g78591 (n_34932, n47014);
  and g78592 (n47016, n_34696, n_34932);
  not g78593 (n_34933, n47015);
  and g78594 (po0813, n_34933, n47016);
  and g78595 (n47018, n_34913, po0954);
  and g78596 (n47019, pi0657, n_34817);
  not g78597 (n_34935, n47018);
  and g78598 (n47020, n_34819, n_34935);
  not g78599 (n_34936, n47019);
  and g78600 (po0814, n_34936, n47020);
  not g78601 (n_34938, pi0658);
  and g78602 (n47022, n_34938, n_34695);
  and g78603 (n47023, n_34926, po0897);
  not g78604 (n_34939, n47022);
  and g78605 (n47024, n_34696, n_34939);
  not g78606 (n_34940, n47023);
  and g78607 (po0815, n_34940, n47024);
  and g78608 (n47026, pi0266, pi0992);
  and g78609 (n47027, n_33067, n47026);
  not g78610 (n_34942, pi0269);
  and g78611 (n47028, n_34942, n47027);
  not g78612 (n_34943, pi0281);
  and g78613 (n47029, n_34943, n47028);
  not g78614 (n_34944, pi0270);
  not g78615 (n_34945, pi0277);
  and g78616 (n47030, n_34944, n_34945);
  not g78617 (n_34946, pi0282);
  and g78618 (n47031, n_34946, n47030);
  and g78619 (n47032, n47029, n47031);
  not g78620 (n_34947, pi0264);
  and g78621 (n47033, n_34947, n47032);
  not g78622 (n_34948, pi0265);
  and g78623 (n47034, n_34948, n47033);
  not g78624 (n_34949, pi0274);
  and g78625 (po0959, n_34949, n47034);
  not g78626 (n_34950, n47034);
  and g78627 (n47036, pi0274, n_34950);
  not g78628 (n_34952, po0959);
  not g78629 (n_34953, n47036);
  and g78630 (po0816, n_34952, n_34953);
  and g78631 (n47038, n_11767, n_34817);
  and g78632 (n47039, n_34731, po0954);
  not g78633 (n_34954, n47038);
  and g78634 (n47040, n_34819, n_34954);
  not g78635 (n_34955, n47039);
  and g78636 (po0817, n_34955, n47040);
  and g78637 (n47042, n_3096, n_34817);
  and g78638 (n47043, n_34765, po0954);
  not g78639 (n_34956, n47042);
  and g78640 (n47044, n_34819, n_34956);
  not g78641 (n_34957, n47043);
  and g78642 (po0818, n_34957, n47044);
  and g78643 (n47046, n_3093, n_34817);
  and g78644 (n47047, n_34757, po0954);
  not g78645 (n_34958, n47046);
  and g78646 (n47048, n_34819, n_34958);
  not g78647 (n_34959, n47047);
  and g78648 (po0819, n_34959, n47048);
  and g78649 (n47050, n_223, n_219);
  and g78650 (n47051, n_7044, n_31932);
  not g78651 (n_34960, pi1065);
  and g78652 (n47052, pi0199, n_34960);
  not g78653 (n_34961, n47050);
  not g78654 (n_34962, n47051);
  and g78655 (n47053, n_34961, n_34962);
  not g78656 (n_34963, n47052);
  and g78657 (n47054, n_34963, n47053);
  and g78658 (n47055, n_4239, n8041);
  and g78659 (n47056, pi0464, n47055);
  not g78660 (n_34964, n47056);
  and g78661 (n47057, pi0588, n_34964);
  and g78662 (n47058, n_4628, pi0592);
  and g78663 (n47059, pi0365, n47058);
  and g78664 (n47060, pi0334, pi0591);
  and g78665 (n47061, n_4239, n47060);
  not g78666 (n_34965, n47059);
  not g78667 (n_34966, n47061);
  and g78668 (n47062, n_34965, n_34966);
  not g78669 (n_34967, n47062);
  and g78670 (n47063, n_4423, n_34967);
  and g78671 (n47064, pi0590, n_4628);
  and g78672 (n47065, n_4239, n47064);
  and g78673 (n47066, pi0323, n47065);
  not g78674 (n_34968, n47066);
  and g78675 (n47067, n_4832, n_34968);
  not g78676 (n_34969, n47063);
  and g78677 (n47068, n_34969, n47067);
  not g78678 (n_34970, n47057);
  and g78679 (n47069, n47050, n_34970);
  not g78680 (n_34971, n47068);
  and g78681 (n47070, n_34971, n47069);
  not g78682 (n_34972, n47054);
  not g78683 (n_34973, n47070);
  and g78684 (n47071, n_34972, n_34973);
  not g78685 (n_34974, n47071);
  and g78686 (n47072, n7643, n_34974);
  and g78687 (n47073, n_2209, n_2030);
  and g78688 (n47074, n_2921, n47073);
  not g78689 (n_34976, pi0784);
  and g78690 (n47075, n_34976, n_2388);
  and g78691 (n47076, n_24930, pi1136);
  not g78692 (n_34977, n47075);
  and g78693 (n47077, pi1135, n_34977);
  not g78694 (n_34978, n47076);
  and g78695 (n47078, n_34978, n47077);
  and g78696 (n47079, n_33464, n_2388);
  and g78697 (n47080, n_24918, pi1136);
  not g78698 (n_34979, n47079);
  and g78699 (n47081, n_2581, n_34979);
  not g78700 (n_34980, n47080);
  and g78701 (n47082, n_34980, n47081);
  not g78702 (n_34981, n47078);
  not g78703 (n_34982, n47082);
  and g78704 (n47083, n_34981, n_34982);
  not g78705 (n_34983, n47083);
  and g78706 (n47084, n47074, n_34983);
  and g78707 (n47085, pi1135, n47073);
  not g78708 (n_34984, n47085);
  and g78709 (n47086, pi1136, n_34984);
  and g78710 (n47087, n_15271, n47086);
  not g78711 (n_34986, pi0855);
  and g78712 (n47088, n_34986, n_2388);
  and g78713 (n47089, n_15317, pi1135);
  and g78714 (n47090, pi1135, n_2388);
  and g78715 (n47091, pi1134, n47073);
  not g78716 (n_34987, n47090);
  and g78717 (n47092, n_34987, n47091);
  not g78724 (n_34991, n47084);
  not g78725 (n_34992, n47095);
  and g78726 (n47096, n_34991, n_34992);
  not g78727 (n_34993, n47096);
  and g78728 (n47097, n_9495, n_34993);
  or g78729 (po0820, n47072, n47097);
  and g78730 (n47099, pi0429, n47055);
  not g78731 (n_34994, n47099);
  and g78732 (n47100, pi0588, n_34994);
  and g78733 (n47101, n_4423, pi0591);
  and g78734 (n47102, pi0404, n47101);
  and g78735 (n47103, n_4423, pi0592);
  not g78736 (n_34995, n47103);
  and g78737 (n47104, n_4832, n_34995);
  not g78738 (n_34996, n47102);
  and g78739 (n47105, n_34996, n47104);
  and g78740 (n47106, pi0380, n_4628);
  not g78741 (n_34997, n47106);
  and g78742 (n47107, pi0592, n_34997);
  not g78743 (n_34998, n47105);
  not g78744 (n_34999, n47107);
  and g78745 (n47108, n_34998, n_34999);
  and g78746 (n47109, pi0355, n47065);
  not g78747 (n_35000, n47108);
  not g78748 (n_35001, n47109);
  and g78749 (n47110, n_35000, n_35001);
  not g78750 (n_35002, n47100);
  and g78751 (n47111, n47050, n_35002);
  not g78752 (n_35003, n47110);
  and g78753 (n47112, n_35003, n47111);
  and g78754 (n47113, n_7044, n_33267);
  and g78755 (n47114, pi0199, n_33268);
  not g78756 (n_35004, n47113);
  and g78757 (n47115, n_34961, n_35004);
  not g78758 (n_35005, n47114);
  and g78759 (n47116, n_35005, n47115);
  not g78760 (n_35006, n47112);
  not g78761 (n_35007, n47116);
  and g78762 (n47117, n_35006, n_35007);
  not g78763 (n_35008, n47117);
  and g78764 (n47118, n7643, n_35008);
  and g78765 (n47119, n_2581, n_2388);
  and g78766 (n47120, pi0872, n47119);
  and g78767 (n47121, n_15864, n_2581);
  and g78768 (n47122, n_15870, pi1135);
  not g78769 (n_35009, n47121);
  and g78770 (n47123, pi1136, n_35009);
  not g78771 (n_35010, n47122);
  and g78772 (n47124, n_35010, n47123);
  not g78773 (n_35011, n47120);
  and g78774 (n47125, pi1134, n_35011);
  not g78775 (n_35012, n47124);
  and g78776 (n47126, n_35012, n47125);
  and g78777 (n47127, n_9495, n47073);
  and g78778 (n47128, pi0614, n_2581);
  and g78779 (n47129, pi0662, pi1135);
  not g78780 (n_35013, n47128);
  and g78781 (n47130, pi1136, n_35013);
  not g78782 (n_35014, n47129);
  and g78783 (n47131, n_35014, n47130);
  and g78784 (n47132, pi0811, n_2581);
  and g78785 (n47133, pi0785, pi1135);
  not g78786 (n_35016, n47132);
  and g78787 (n47134, n_2388, n_35016);
  not g78788 (n_35017, n47133);
  and g78789 (n47135, n_35017, n47134);
  not g78790 (n_35018, n47131);
  not g78791 (n_35019, n47135);
  and g78792 (n47136, n_35018, n_35019);
  not g78793 (n_35020, n47136);
  and g78794 (n47137, n_2921, n_35020);
  not g78795 (n_35021, n47126);
  and g78796 (n47138, n_35021, n47127);
  not g78797 (n_35022, n47137);
  and g78798 (n47139, n_35022, n47138);
  or g78799 (po0821, n47118, n47139);
  and g78800 (n47141, n_12032, n_34817);
  and g78801 (n47142, n_34792, po0954);
  not g78802 (n_35023, n47141);
  and g78803 (n47143, n_34819, n_35023);
  not g78804 (n_35024, n47142);
  and g78805 (po0822, n_35024, n47143);
  and g78806 (n47145, n_26264, n_2581);
  and g78807 (n47146, n_26247, pi1135);
  not g78808 (n_35025, n47145);
  and g78809 (n47147, pi1136, n_35025);
  not g78810 (n_35026, n47146);
  and g78811 (n47148, n_35026, n47147);
  and g78812 (n47149, n_12411, pi1135);
  and g78813 (n47150, pi0799, n_2581);
  not g78814 (n_35028, n47149);
  and g78815 (n47151, n_2388, n_35028);
  not g78816 (n_35029, n47150);
  and g78817 (n47152, n_35029, n47151);
  not g78818 (n_35030, n47148);
  not g78819 (n_35031, n47152);
  and g78820 (n47153, n_35030, n_35031);
  not g78821 (n_35032, n47153);
  and g78822 (n47154, n47074, n_35032);
  and g78823 (n47155, n_16132, n47086);
  and g78824 (n47156, n_16177, pi1135);
  not g78825 (n_35034, pi0873);
  and g78826 (n47157, n_35034, n_2388);
  not g78833 (n_35038, n47154);
  not g78834 (n_35039, n47160);
  and g78835 (n47161, n_35038, n_35039);
  not g78836 (n_35040, n47161);
  and g78837 (n47162, n_9495, n_35040);
  and g78838 (n47163, n_7044, n_33292);
  and g78839 (n47164, pi0199, n_33293);
  not g78840 (n_35041, n47163);
  and g78841 (n47165, n_34961, n_35041);
  not g78842 (n_35042, n47164);
  and g78843 (n47166, n_35042, n47165);
  and g78844 (n47167, pi0443, n47055);
  not g78845 (n_35043, n47167);
  and g78846 (n47168, pi0588, n_35043);
  and g78847 (n47169, pi0456, n47101);
  not g78848 (n_35044, n47169);
  and g78849 (n47170, n47104, n_35044);
  and g78850 (n47171, pi0337, n_4628);
  not g78851 (n_35045, n47171);
  and g78852 (n47172, pi0592, n_35045);
  not g78853 (n_35046, n47170);
  not g78854 (n_35047, n47172);
  and g78855 (n47173, n_35046, n_35047);
  and g78856 (n47174, pi0441, n47065);
  not g78857 (n_35048, n47173);
  not g78858 (n_35049, n47174);
  and g78859 (n47175, n_35048, n_35049);
  not g78860 (n_35050, n47168);
  and g78861 (n47176, n47050, n_35050);
  not g78862 (n_35051, n47175);
  and g78863 (n47177, n_35051, n47176);
  not g78864 (n_35052, n47166);
  not g78865 (n_35053, n47177);
  and g78866 (n47178, n_35052, n_35053);
  not g78867 (n_35054, n47178);
  and g78868 (n47179, n7643, n_35054);
  or g78869 (po0823, n47162, n47179);
  and g78870 (n47181, pi0444, n47055);
  not g78871 (n_35055, n47181);
  and g78872 (n47182, pi0588, n_35055);
  and g78873 (n47183, pi0319, n47101);
  not g78874 (n_35056, n47183);
  and g78875 (n47184, n47104, n_35056);
  and g78876 (n47185, pi0338, n_4628);
  not g78877 (n_35057, n47185);
  and g78878 (n47186, pi0592, n_35057);
  not g78879 (n_35058, n47184);
  not g78880 (n_35059, n47186);
  and g78881 (n47187, n_35058, n_35059);
  and g78882 (n47188, pi0458, n47065);
  not g78883 (n_35060, n47187);
  not g78884 (n_35061, n47188);
  and g78885 (n47189, n_35060, n_35061);
  not g78886 (n_35062, n47182);
  and g78887 (n47190, n47050, n_35062);
  not g78888 (n_35063, n47189);
  and g78889 (n47191, n_35063, n47190);
  and g78890 (n47192, n_7044, n_33277);
  and g78891 (n47193, pi0199, n_33278);
  not g78892 (n_35064, n47192);
  and g78893 (n47194, n_34961, n_35064);
  not g78894 (n_35065, n47193);
  and g78895 (n47195, n_35065, n47194);
  not g78896 (n_35066, n47191);
  not g78897 (n_35067, n47195);
  and g78898 (n47196, n_35066, n_35067);
  not g78899 (n_35068, n47196);
  and g78900 (n47197, n7643, n_35068);
  and g78901 (n47198, pi0871, n47119);
  and g78902 (n47199, n_15951, n_2581);
  and g78903 (n47200, n_15996, pi1135);
  not g78904 (n_35069, n47199);
  and g78905 (n47201, pi1136, n_35069);
  not g78906 (n_35070, n47200);
  and g78907 (n47202, n_35070, n47201);
  not g78908 (n_35071, n47198);
  and g78909 (n47203, pi1134, n_35071);
  not g78910 (n_35072, n47202);
  and g78911 (n47204, n_35072, n47203);
  and g78912 (n47205, pi0792, n_2388);
  and g78913 (n47206, pi0681, pi1136);
  not g78914 (n_35073, n47205);
  and g78915 (n47207, pi1135, n_35073);
  not g78916 (n_35074, n47206);
  and g78917 (n47208, n_35074, n47207);
  not g78918 (n_35076, pi0809);
  and g78919 (n47209, n_35076, n_2388);
  and g78920 (n47210, pi0642, pi1136);
  not g78921 (n_35077, n47209);
  and g78922 (n47211, n_2581, n_35077);
  not g78923 (n_35078, n47210);
  and g78924 (n47212, n_35078, n47211);
  not g78925 (n_35079, n47208);
  not g78926 (n_35080, n47212);
  and g78927 (n47213, n_35079, n_35080);
  not g78928 (n_35081, n47213);
  and g78929 (n47214, n_2921, n_35081);
  not g78930 (n_35082, n47204);
  and g78931 (n47215, n47127, n_35082);
  not g78932 (n_35083, n47214);
  and g78933 (n47216, n_35083, n47215);
  or g78934 (po0824, n47197, n47216);
  and g78935 (n47218, n_11512, n_2581);
  and g78936 (n47219, n_11502, pi1135);
  not g78937 (n_35084, n47218);
  and g78938 (n47220, pi1136, n_35084);
  not g78939 (n_35085, n47219);
  and g78940 (n47221, n_35085, n47220);
  not g78941 (n_35087, pi0981);
  and g78942 (n47222, n_35087, n_2581);
  and g78943 (n47223, n_11749, pi1135);
  not g78944 (n_35088, n47222);
  and g78945 (n47224, n_2388, n_35088);
  not g78946 (n_35089, n47223);
  and g78947 (n47225, n_35089, n47224);
  not g78948 (n_35090, n47221);
  not g78949 (n_35091, n47225);
  and g78950 (n47226, n_35090, n_35091);
  not g78951 (n_35092, n47226);
  and g78952 (n47227, n47074, n_35092);
  and g78953 (n47228, n_15215, n47086);
  and g78954 (n47229, n_15254, pi1135);
  and g78955 (n47230, n_34719, n_2388);
  not g78962 (n_35096, n47227);
  not g78963 (n_35097, n47233);
  and g78964 (n47234, n_35096, n_35097);
  not g78965 (n_35098, n47234);
  and g78966 (n47235, n_9495, n_35098);
  and g78967 (n47236, n_7044, n_33262);
  and g78968 (n47237, pi0199, n_33263);
  not g78969 (n_35099, n47236);
  and g78970 (n47238, n_34961, n_35099);
  not g78971 (n_35100, n47237);
  and g78972 (n47239, n_35100, n47238);
  and g78973 (n47240, pi0414, n47055);
  not g78974 (n_35101, n47240);
  and g78975 (n47241, pi0588, n_35101);
  and g78976 (n47242, pi0390, n47101);
  not g78977 (n_35102, n47242);
  and g78978 (n47243, n47104, n_35102);
  and g78979 (n47244, pi0363, n_4628);
  not g78980 (n_35103, n47244);
  and g78981 (n47245, pi0592, n_35103);
  not g78982 (n_35104, n47243);
  not g78983 (n_35105, n47245);
  and g78984 (n47246, n_35104, n_35105);
  and g78985 (n47247, pi0342, n47065);
  not g78986 (n_35106, n47246);
  not g78987 (n_35107, n47247);
  and g78988 (n47248, n_35106, n_35107);
  not g78989 (n_35108, n47241);
  and g78990 (n47249, n47050, n_35108);
  not g78991 (n_35109, n47248);
  and g78992 (n47250, n_35109, n47249);
  not g78993 (n_35110, n47239);
  not g78994 (n_35111, n47250);
  and g78995 (n47251, n_35110, n_35111);
  not g78996 (n_35112, n47251);
  and g78997 (n47252, n7643, n_35112);
  or g78998 (po0825, n47235, n47252);
  and g78999 (n47254, n_34886, po0954);
  and g79000 (n47255, pi0669, n_34817);
  not g79001 (n_35114, n47254);
  and g79002 (n47256, n_34819, n_35114);
  not g79003 (n_35115, n47255);
  and g79004 (po0826, n_35115, n47256);
  and g79005 (n47258, n_7044, n_31940);
  not g79006 (n_35116, pi1062);
  and g79007 (n47259, pi0199, n_35116);
  not g79008 (n_35117, n47258);
  and g79009 (n47260, n_34961, n_35117);
  not g79010 (n_35118, n47259);
  and g79011 (n47261, n_35118, n47260);
  and g79012 (n47262, pi0415, n47055);
  not g79013 (n_35119, n47262);
  and g79014 (n47263, pi0588, n_35119);
  and g79015 (n47264, pi0364, n47058);
  and g79016 (n47265, pi0391, pi0591);
  and g79017 (n47266, n_4239, n47265);
  not g79018 (n_35120, n47264);
  not g79019 (n_35121, n47266);
  and g79020 (n47267, n_35120, n_35121);
  not g79021 (n_35122, n47267);
  and g79022 (n47268, n_4423, n_35122);
  and g79023 (n47269, pi0343, n47065);
  not g79024 (n_35123, n47269);
  and g79025 (n47270, n_4832, n_35123);
  not g79026 (n_35124, n47268);
  and g79027 (n47271, n_35124, n47270);
  not g79028 (n_35125, n47263);
  and g79029 (n47272, n47050, n_35125);
  not g79030 (n_35126, n47271);
  and g79031 (n47273, n_35126, n47272);
  not g79032 (n_35127, n47261);
  not g79033 (n_35128, n47273);
  and g79034 (n47274, n_35127, n_35128);
  not g79035 (n_35129, n47274);
  and g79036 (n47275, n7643, n_35129);
  and g79037 (n47276, pi0723, pi1135);
  not g79038 (n_35131, pi0852);
  and g79039 (n47277, n_35131, n_2388);
  and g79040 (n47278, pi0745, n47086);
  and g79047 (n47282, pi0695, pi1135);
  and g79048 (n47283, pi1136, n47073);
  and g79049 (n47284, n_26742, n_2581);
  not g79055 (n_35137, n47281);
  not g79056 (n_35138, n47287);
  and g79057 (n47288, n_35137, n_35138);
  not g79058 (n_35139, n47288);
  and g79059 (n47289, n_9495, n_35139);
  or g79060 (po0827, n47275, n47289);
  not g79061 (n_35140, pi0261);
  and g79062 (n47291, n_7044, n_35140);
  not g79063 (n_35141, pi1040);
  and g79064 (n47292, pi0199, n_35141);
  not g79065 (n_35142, n47291);
  and g79066 (n47293, n_34961, n_35142);
  not g79067 (n_35143, n47292);
  and g79068 (n47294, n_35143, n47293);
  and g79069 (n47295, pi0453, n47055);
  not g79070 (n_35144, n47295);
  and g79071 (n47296, pi0588, n_35144);
  and g79072 (n47297, pi0447, n47058);
  and g79073 (n47298, pi0333, pi0591);
  and g79074 (n47299, n_4239, n47298);
  not g79075 (n_35145, n47297);
  not g79076 (n_35146, n47299);
  and g79077 (n47300, n_35145, n_35146);
  not g79078 (n_35147, n47300);
  and g79079 (n47301, n_4423, n_35147);
  and g79080 (n47302, pi0327, n47065);
  not g79081 (n_35148, n47302);
  and g79082 (n47303, n_4832, n_35148);
  not g79083 (n_35149, n47301);
  and g79084 (n47304, n_35149, n47303);
  not g79085 (n_35150, n47296);
  and g79086 (n47305, n47050, n_35150);
  not g79087 (n_35151, n47304);
  and g79088 (n47306, n_35151, n47305);
  not g79089 (n_35152, n47294);
  not g79090 (n_35153, n47306);
  and g79091 (n47307, n_35152, n_35153);
  not g79092 (n_35154, n47307);
  and g79093 (n47308, n7643, n_35154);
  and g79094 (n47309, pi0724, pi1135);
  not g79095 (n_35156, pi0865);
  and g79096 (n47310, n_35156, n_2388);
  and g79097 (n47311, pi0741, n47086);
  and g79104 (n47315, pi0646, pi1135);
  and g79105 (n47316, n_34741, n_2581);
  not g79111 (n_35162, n47314);
  not g79112 (n_35163, n47319);
  and g79113 (n47320, n_35162, n_35163);
  not g79114 (n_35164, n47320);
  and g79115 (n47321, n_9495, n_35164);
  or g79116 (po0828, n47308, n47321);
  and g79117 (n47323, n_3091, n_2581);
  and g79118 (n47324, n_3096, pi1135);
  not g79119 (n_35165, n47323);
  and g79120 (n47325, pi1136, n_35165);
  not g79121 (n_35166, n47324);
  and g79122 (n47326, n_35166, n47325);
  not g79123 (n_35168, pi0808);
  and g79124 (n47327, n_35168, n_2581);
  and g79125 (n47328, n_11981, pi1135);
  not g79126 (n_35169, n47327);
  and g79127 (n47329, n_2388, n_35169);
  not g79128 (n_35170, n47328);
  and g79129 (n47330, n_35170, n47329);
  not g79130 (n_35171, n47326);
  not g79131 (n_35172, n47330);
  and g79132 (n47331, n_35171, n_35172);
  not g79133 (n_35173, n47331);
  and g79134 (n47332, n47074, n_35173);
  and g79135 (n47333, n_14083, n47086);
  and g79136 (n47334, n_14126, pi1135);
  and g79137 (n47335, n_34774, n_2388);
  not g79144 (n_35177, n47332);
  not g79145 (n_35178, n47338);
  and g79146 (n47339, n_35177, n_35178);
  not g79147 (n_35179, n47339);
  and g79148 (n47340, n_9495, n_35179);
  and g79149 (n47341, n_7044, n_33257);
  and g79150 (n47342, pi0199, n_33258);
  not g79151 (n_35180, n47341);
  and g79152 (n47343, n_34961, n_35180);
  not g79153 (n_35181, n47342);
  and g79154 (n47344, n_35181, n47343);
  and g79155 (n47345, pi0422, n47055);
  not g79156 (n_35182, n47345);
  and g79157 (n47346, pi0588, n_35182);
  and g79158 (n47347, pi0397, n47101);
  not g79159 (n_35183, n47347);
  and g79160 (n47348, n47104, n_35183);
  and g79161 (n47349, pi0372, n_4628);
  not g79162 (n_35184, n47349);
  and g79163 (n47350, pi0592, n_35184);
  not g79164 (n_35185, n47348);
  not g79165 (n_35186, n47350);
  and g79166 (n47351, n_35185, n_35186);
  and g79167 (n47352, pi0320, n47065);
  not g79168 (n_35187, n47351);
  not g79169 (n_35188, n47352);
  and g79170 (n47353, n_35187, n_35188);
  not g79171 (n_35189, n47346);
  and g79172 (n47354, n47050, n_35189);
  not g79173 (n_35190, n47353);
  and g79174 (n47355, n_35190, n47354);
  not g79175 (n_35191, n47344);
  not g79176 (n_35192, n47355);
  and g79177 (n47356, n_35191, n_35192);
  not g79178 (n_35193, n47356);
  and g79179 (n47357, n7643, n_35193);
  or g79180 (po0829, n47340, n47357);
  and g79181 (n47359, n_25117, n_2581);
  and g79182 (n47360, n_25155, pi1135);
  not g79183 (n_35194, n47359);
  and g79184 (n47361, pi1136, n_35194);
  not g79185 (n_35195, n47360);
  and g79186 (n47362, n_35195, n47361);
  and g79187 (n47363, n_12318, pi1135);
  and g79188 (n47364, pi0814, n_2581);
  not g79189 (n_35197, n47363);
  and g79190 (n47365, n_2388, n_35197);
  not g79191 (n_35198, n47364);
  and g79192 (n47366, n_35198, n47365);
  not g79193 (n_35199, n47362);
  not g79194 (n_35200, n47366);
  and g79195 (n47367, n_35199, n_35200);
  not g79196 (n_35201, n47367);
  and g79197 (n47368, n47074, n_35201);
  and g79198 (n47369, n_12661, n47086);
  and g79199 (n47370, n_12614, pi1135);
  not g79200 (n_35203, pi0866);
  and g79201 (n47371, n_35203, n_2388);
  not g79208 (n_35207, n47368);
  not g79209 (n_35208, n47374);
  and g79210 (n47375, n_35207, n_35208);
  not g79211 (n_35209, n47375);
  and g79212 (n47376, n_9495, n_35209);
  and g79213 (n47377, n_7044, n_33282);
  and g79214 (n47378, pi0199, n_33283);
  not g79215 (n_35210, n47377);
  and g79216 (n47379, n_34961, n_35210);
  not g79217 (n_35211, n47378);
  and g79218 (n47380, n_35211, n47379);
  and g79219 (n47381, pi0435, n47055);
  not g79220 (n_35212, n47381);
  and g79221 (n47382, pi0588, n_35212);
  and g79222 (n47383, pi0411, n47101);
  not g79223 (n_35213, n47383);
  and g79224 (n47384, n47104, n_35213);
  and g79225 (n47385, pi0387, n_4628);
  not g79226 (n_35214, n47385);
  and g79227 (n47386, pi0592, n_35214);
  not g79228 (n_35215, n47384);
  not g79229 (n_35216, n47386);
  and g79230 (n47387, n_35215, n_35216);
  and g79231 (n47388, pi0452, n47065);
  not g79232 (n_35217, n47387);
  not g79233 (n_35218, n47388);
  and g79234 (n47389, n_35217, n_35218);
  not g79235 (n_35219, n47382);
  and g79236 (n47390, n47050, n_35219);
  not g79237 (n_35220, n47389);
  and g79238 (n47391, n_35220, n47390);
  not g79239 (n_35221, n47380);
  not g79240 (n_35222, n47391);
  and g79241 (n47392, n_35221, n_35222);
  not g79242 (n_35223, n47392);
  and g79243 (n47393, n7643, n_35223);
  or g79244 (po0830, n47376, n47393);
  and g79245 (n47395, n_7044, n_31924);
  not g79246 (n_35224, pi1070);
  and g79247 (n47396, pi0199, n_35224);
  not g79248 (n_35225, n47395);
  and g79249 (n47397, n_34961, n_35225);
  not g79250 (n_35226, n47396);
  and g79251 (n47398, n_35226, n47397);
  and g79252 (n47399, pi0437, n47055);
  not g79253 (n_35227, n47399);
  and g79254 (n47400, pi0588, n_35227);
  and g79255 (n47401, pi0336, n47058);
  and g79256 (n47402, pi0463, pi0591);
  and g79257 (n47403, n_4239, n47402);
  not g79258 (n_35228, n47401);
  not g79259 (n_35229, n47403);
  and g79260 (n47404, n_35228, n_35229);
  not g79261 (n_35230, n47404);
  and g79262 (n47405, n_4423, n_35230);
  and g79263 (n47406, pi0362, n47065);
  not g79264 (n_35231, n47406);
  and g79265 (n47407, n_4832, n_35231);
  not g79266 (n_35232, n47405);
  and g79267 (n47408, n_35232, n47407);
  not g79268 (n_35233, n47400);
  and g79269 (n47409, n47050, n_35233);
  not g79270 (n_35234, n47408);
  and g79271 (n47410, n_35234, n47409);
  not g79272 (n_35235, n47398);
  not g79273 (n_35236, n47410);
  and g79274 (n47411, n_35235, n_35236);
  not g79275 (n_35237, n47411);
  and g79276 (n47412, n7643, n_35237);
  and g79277 (n47413, pi0859, n47119);
  and g79278 (n47414, n_13140, n_2581);
  and g79279 (n47415, n_13045, pi1135);
  not g79280 (n_35239, n47414);
  and g79281 (n47416, pi1136, n_35239);
  not g79282 (n_35240, n47415);
  and g79283 (n47417, n_35240, n47416);
  not g79284 (n_35241, n47413);
  and g79285 (n47418, pi1134, n_35241);
  not g79286 (n_35242, n47417);
  and g79287 (n47419, n_35242, n47418);
  and g79288 (n47420, pi0622, n_2581);
  and g79289 (n47421, pi0639, pi1135);
  not g79290 (n_35243, n47420);
  and g79291 (n47422, pi1136, n_35243);
  not g79292 (n_35244, n47421);
  and g79293 (n47423, n_35244, n47422);
  and g79294 (n47424, pi0804, n_2581);
  and g79295 (n47425, pi0783, pi1135);
  not g79296 (n_35246, n47424);
  and g79297 (n47426, n_2388, n_35246);
  not g79298 (n_35247, n47425);
  and g79299 (n47427, n_35247, n47426);
  not g79300 (n_35248, n47423);
  not g79301 (n_35249, n47427);
  and g79302 (n47428, n_35248, n_35249);
  not g79303 (n_35250, n47428);
  and g79304 (n47429, n_2921, n_35250);
  not g79305 (n_35251, n47419);
  and g79306 (n47430, n47127, n_35251);
  not g79307 (n_35252, n47429);
  and g79308 (n47431, n_35252, n47430);
  or g79309 (po0831, n47412, n47431);
  and g79310 (n47433, pi0876, n47119);
  and g79311 (n47434, n_16089, n_2581);
  and g79312 (n47435, n_16117, pi1135);
  not g79313 (n_35254, n47434);
  and g79314 (n47436, pi1136, n_35254);
  not g79315 (n_35255, n47435);
  and g79316 (n47437, n_35255, n47436);
  not g79317 (n_35256, n47433);
  not g79318 (n_35257, n47437);
  and g79319 (n47438, n_35256, n_35257);
  not g79320 (n_35258, n47438);
  and g79321 (n47439, n47091, n_35258);
  and g79322 (n47440, n_25938, n47086);
  and g79323 (n47441, pi0789, n47090);
  and g79324 (n47442, n_25879, pi1135);
  not g79325 (n_35259, n47442);
  and g79326 (n47443, pi1136, n_35259);
  not g79327 (n_35261, pi0803);
  and g79328 (n47444, n_35261, n_2581);
  not g79329 (n_35262, n47441);
  not g79330 (n_35263, n47444);
  and g79331 (n47445, n_35262, n_35263);
  not g79332 (n_35264, n47443);
  and g79333 (n47446, n_35264, n47445);
  not g79334 (n_35265, n47440);
  and g79335 (n47447, n47074, n_35265);
  not g79336 (n_35266, n47446);
  and g79337 (n47448, n_35266, n47447);
  not g79338 (n_35267, n47439);
  not g79339 (n_35268, n47448);
  and g79340 (n47449, n_35267, n_35268);
  not g79341 (n_35269, n47449);
  and g79342 (n47450, n_9495, n_35269);
  and g79343 (n47451, n_7044, n_33287);
  and g79344 (n47452, pi0199, n_33288);
  not g79345 (n_35270, n47451);
  and g79346 (n47453, n_34961, n_35270);
  not g79347 (n_35271, n47452);
  and g79348 (n47454, n_35271, n47453);
  and g79349 (n47455, pi0436, n47055);
  not g79350 (n_35272, n47455);
  and g79351 (n47456, pi0588, n_35272);
  and g79352 (n47457, pi0412, n47101);
  not g79353 (n_35273, n47457);
  and g79354 (n47458, n47104, n_35273);
  and g79355 (n47459, pi0388, n_4628);
  not g79356 (n_35274, n47459);
  and g79357 (n47460, pi0592, n_35274);
  not g79358 (n_35275, n47458);
  not g79359 (n_35276, n47460);
  and g79360 (n47461, n_35275, n_35276);
  and g79361 (n47462, pi0455, n47065);
  not g79362 (n_35277, n47461);
  not g79363 (n_35278, n47462);
  and g79364 (n47463, n_35277, n_35278);
  not g79365 (n_35279, n47456);
  and g79366 (n47464, n47050, n_35279);
  not g79367 (n_35280, n47463);
  and g79368 (n47465, n_35280, n47464);
  not g79369 (n_35281, n47454);
  not g79370 (n_35282, n47465);
  and g79371 (n47466, n_35281, n_35282);
  not g79372 (n_35283, n47466);
  and g79373 (n47467, n7643, n_35283);
  or g79374 (po0832, n47450, n47467);
  and g79375 (n47469, n_25343, n_2581);
  and g79376 (n47470, n_25400, pi1135);
  not g79377 (n_35284, n47469);
  and g79378 (n47471, pi1136, n_35284);
  not g79379 (n_35285, n47470);
  and g79380 (n47472, n_35285, n47471);
  and g79381 (n47473, n_11803, pi1135);
  and g79382 (n47474, pi0812, n_2581);
  not g79383 (n_35287, n47473);
  and g79384 (n47475, n_2388, n_35287);
  not g79385 (n_35288, n47474);
  and g79386 (n47476, n_35288, n47475);
  not g79387 (n_35289, n47472);
  not g79388 (n_35290, n47476);
  and g79389 (n47477, n_35289, n_35290);
  not g79390 (n_35291, n47477);
  and g79391 (n47478, n47074, n_35291);
  and g79392 (n47479, n_16011, n47086);
  and g79393 (n47480, n_16056, pi1135);
  not g79394 (n_35293, pi0881);
  and g79395 (n47481, n_35293, n_2388);
  not g79402 (n_35297, n47478);
  not g79403 (n_35298, n47484);
  and g79404 (n47485, n_35297, n_35298);
  not g79405 (n_35299, n47485);
  and g79406 (n47486, n_9495, n_35299);
  and g79407 (n47487, n_7044, n_33272);
  and g79408 (n47488, pi0199, n_33273);
  not g79409 (n_35300, n47487);
  and g79410 (n47489, n_34961, n_35300);
  not g79411 (n_35301, n47488);
  and g79412 (n47490, n_35301, n47489);
  and g79413 (n47491, pi0434, n47055);
  not g79414 (n_35302, n47491);
  and g79415 (n47492, pi0588, n_35302);
  and g79416 (n47493, pi0410, n47101);
  not g79417 (n_35303, n47493);
  and g79418 (n47494, n47104, n_35303);
  and g79419 (n47495, pi0386, n_4628);
  not g79420 (n_35304, n47495);
  and g79421 (n47496, pi0592, n_35304);
  not g79422 (n_35305, n47494);
  not g79423 (n_35306, n47496);
  and g79424 (n47497, n_35305, n_35306);
  and g79425 (n47498, pi0361, n47065);
  not g79426 (n_35307, n47497);
  not g79427 (n_35308, n47498);
  and g79428 (n47499, n_35307, n_35308);
  not g79429 (n_35309, n47492);
  and g79430 (n47500, n47050, n_35309);
  not g79431 (n_35310, n47499);
  and g79432 (n47501, n_35310, n47500);
  not g79433 (n_35311, n47490);
  not g79434 (n_35312, n47501);
  and g79435 (n47502, n_35311, n_35312);
  not g79436 (n_35313, n47502);
  and g79437 (n47503, n7643, n_35313);
  or g79438 (po0833, n47486, n47503);
  and g79439 (n47505, n_7044, n_31948);
  not g79440 (n_35314, pi1069);
  and g79441 (n47506, pi0199, n_35314);
  not g79442 (n_35315, n47505);
  and g79443 (n47507, n_34961, n_35315);
  not g79444 (n_35316, n47506);
  and g79445 (n47508, n_35316, n47507);
  and g79446 (n47509, pi0416, n47055);
  not g79447 (n_35317, n47509);
  and g79448 (n47510, pi0588, n_35317);
  and g79449 (n47511, pi0366, n47058);
  and g79450 (n47512, pi0335, pi0591);
  and g79451 (n47513, n_4239, n47512);
  not g79452 (n_35318, n47511);
  not g79453 (n_35319, n47513);
  and g79454 (n47514, n_35318, n_35319);
  not g79455 (n_35320, n47514);
  and g79456 (n47515, n_4423, n_35320);
  and g79457 (n47516, pi0344, n47065);
  not g79458 (n_35321, n47516);
  and g79459 (n47517, n_4832, n_35321);
  not g79460 (n_35322, n47515);
  and g79461 (n47518, n_35322, n47517);
  not g79462 (n_35323, n47510);
  and g79463 (n47519, n47050, n_35323);
  not g79464 (n_35324, n47518);
  and g79465 (n47520, n_35324, n47519);
  not g79466 (n_35325, n47508);
  not g79467 (n_35326, n47520);
  and g79468 (n47521, n_35325, n_35326);
  not g79469 (n_35327, n47521);
  and g79470 (n47522, n7643, n_35327);
  and g79471 (n47523, pi0704, pi1135);
  not g79472 (n_35329, pi0870);
  and g79473 (n47524, n_35329, n_2388);
  and g79474 (n47525, pi0742, n47086);
  and g79481 (n47529, pi0635, pi1135);
  and g79482 (n47530, n_34786, n_2581);
  not g79488 (n_35335, n47528);
  not g79489 (n_35336, n47533);
  and g79490 (n47534, n_35335, n_35336);
  not g79491 (n_35337, n47534);
  and g79492 (n47535, n_9495, n_35337);
  or g79493 (po0834, n47522, n47535);
  not g79494 (n_35338, pi0260);
  and g79495 (n47537, n_7044, n_35338);
  not g79496 (n_35339, pi1067);
  and g79497 (n47538, pi0199, n_35339);
  not g79498 (n_35340, n47537);
  and g79499 (n47539, n_34961, n_35340);
  not g79500 (n_35341, n47538);
  and g79501 (n47540, n_35341, n47539);
  and g79502 (n47541, pi0418, n47055);
  not g79503 (n_35342, n47541);
  and g79504 (n47542, pi0588, n_35342);
  and g79505 (n47543, pi0368, n47058);
  and g79506 (n47544, pi0393, pi0591);
  and g79507 (n47545, n_4239, n47544);
  not g79508 (n_35343, n47543);
  not g79509 (n_35344, n47545);
  and g79510 (n47546, n_35343, n_35344);
  not g79511 (n_35345, n47546);
  and g79512 (n47547, n_4423, n_35345);
  and g79513 (n47548, pi0346, n47065);
  not g79514 (n_35346, n47548);
  and g79515 (n47549, n_4832, n_35346);
  not g79516 (n_35347, n47547);
  and g79517 (n47550, n_35347, n47549);
  not g79518 (n_35348, n47542);
  and g79519 (n47551, n47050, n_35348);
  not g79520 (n_35349, n47550);
  and g79521 (n47552, n_35349, n47551);
  not g79522 (n_35350, n47540);
  not g79523 (n_35351, n47552);
  and g79524 (n47553, n_35350, n_35351);
  not g79525 (n_35352, n47553);
  and g79526 (n47554, n7643, n_35352);
  and g79527 (n47555, pi0688, pi1135);
  not g79528 (n_35354, pi0856);
  and g79529 (n47556, n_35354, n_2388);
  and g79530 (n47557, pi0760, n47086);
  and g79537 (n47561, pi0632, pi1135);
  and g79538 (n47562, n_34751, n_2581);
  not g79544 (n_35360, n47560);
  not g79545 (n_35361, n47565);
  and g79546 (n47566, n_35360, n_35361);
  not g79547 (n_35362, n47566);
  and g79548 (n47567, n_9495, n_35362);
  or g79549 (po0835, n47554, n47567);
  and g79550 (n47569, n_7044, n_31916);
  not g79551 (n_35363, pi1036);
  and g79552 (n47570, pi0199, n_35363);
  not g79553 (n_35364, n47569);
  and g79554 (n47571, n_34961, n_35364);
  not g79555 (n_35365, n47570);
  and g79556 (n47572, n_35365, n47571);
  and g79557 (n47573, pi0438, n47055);
  not g79558 (n_35366, n47573);
  and g79559 (n47574, pi0588, n_35366);
  and g79560 (n47575, pi0389, n47058);
  and g79561 (n47576, pi0413, pi0591);
  and g79562 (n47577, n_4239, n47576);
  not g79563 (n_35367, n47575);
  not g79564 (n_35368, n47577);
  and g79565 (n47578, n_35367, n_35368);
  not g79566 (n_35369, n47578);
  and g79567 (n47579, n_4423, n_35369);
  and g79568 (n47580, pi0450, n47065);
  not g79569 (n_35370, n47580);
  and g79570 (n47581, n_4832, n_35370);
  not g79571 (n_35371, n47579);
  and g79572 (n47582, n_35371, n47581);
  not g79573 (n_35372, n47574);
  and g79574 (n47583, n47050, n_35372);
  not g79575 (n_35373, n47582);
  and g79576 (n47584, n_35373, n47583);
  not g79577 (n_35374, n47572);
  not g79578 (n_35375, n47584);
  and g79579 (n47585, n_35374, n_35375);
  not g79580 (n_35376, n47585);
  and g79581 (n47586, n7643, n_35376);
  not g79582 (n_35378, pi0791);
  and g79583 (n47587, n_35378, n_2388);
  and g79584 (n47588, n_12032, pi1136);
  not g79585 (n_35379, n47587);
  and g79586 (n47589, pi1135, n_35379);
  not g79587 (n_35380, n47588);
  and g79588 (n47590, n_35380, n47589);
  and g79589 (n47591, n_33448, n_2388);
  and g79590 (n47592, n_12038, pi1136);
  not g79591 (n_35381, n47591);
  and g79592 (n47593, n_2581, n_35381);
  not g79593 (n_35382, n47592);
  and g79594 (n47594, n_35382, n47593);
  not g79595 (n_35383, n47590);
  not g79596 (n_35384, n47594);
  and g79597 (n47595, n_35383, n_35384);
  not g79598 (n_35385, n47595);
  and g79599 (n47596, n47074, n_35385);
  and g79600 (n47597, n_16204, n47086);
  not g79601 (n_35387, pi0874);
  and g79602 (n47598, n_35387, n_2388);
  and g79603 (n47599, n_16236, pi1135);
  not g79610 (n_35391, n47596);
  not g79611 (n_35392, n47602);
  and g79612 (n47603, n_35391, n_35392);
  not g79613 (n_35393, n47603);
  and g79614 (n47604, n_9495, n_35393);
  or g79615 (po0836, n47586, n47604);
  and g79616 (n47606, n_11502, n_34817);
  and g79617 (n47607, n_34686, po0954);
  not g79618 (n_35394, n47606);
  and g79619 (n47608, n_34819, n_35394);
  not g79620 (n_35395, n47607);
  and g79621 (po0837, n_35395, n47608);
  and g79622 (n47610, n_3098, n_34817);
  and g79623 (n47611, n_34874, po0954);
  not g79624 (n_35396, n47610);
  and g79625 (n47612, n_34819, n_35396);
  not g79626 (n_35397, n47611);
  and g79627 (po0838, n_35397, n47612);
  not g79628 (n_35398, pi0251);
  and g79629 (n47614, n_7044, n_35398);
  not g79630 (n_35399, pi1039);
  and g79631 (n47615, pi0199, n_35399);
  not g79632 (n_35400, n47614);
  and g79633 (n47616, n_34961, n_35400);
  not g79634 (n_35401, n47615);
  and g79635 (n47617, n_35401, n47616);
  and g79636 (n47618, pi0417, n47055);
  not g79637 (n_35402, n47618);
  and g79638 (n47619, pi0588, n_35402);
  and g79639 (n47620, pi0367, n47058);
  and g79640 (n47621, pi0392, pi0591);
  and g79641 (n47622, n_4239, n47621);
  not g79642 (n_35403, n47620);
  not g79643 (n_35404, n47622);
  and g79644 (n47623, n_35403, n_35404);
  not g79645 (n_35405, n47623);
  and g79646 (n47624, n_4423, n_35405);
  and g79647 (n47625, pi0345, n47065);
  not g79648 (n_35406, n47625);
  and g79649 (n47626, n_4832, n_35406);
  not g79650 (n_35407, n47624);
  and g79651 (n47627, n_35407, n47626);
  not g79652 (n_35408, n47619);
  and g79653 (n47628, n47050, n_35408);
  not g79654 (n_35409, n47627);
  and g79655 (n47629, n_35409, n47628);
  not g79656 (n_35410, n47617);
  not g79657 (n_35411, n47629);
  and g79658 (n47630, n_35410, n_35411);
  not g79659 (n_35412, n47630);
  and g79660 (n47631, n7643, n_35412);
  and g79661 (n47632, pi0686, pi1135);
  not g79662 (n_35414, pi0848);
  and g79663 (n47633, n_35414, n_2388);
  and g79664 (n47634, pi0757, n47086);
  and g79671 (n47638, pi0631, pi1135);
  and g79672 (n47639, n_34735, n_2581);
  not g79678 (n_35420, n47637);
  not g79679 (n_35421, n47642);
  and g79680 (n47643, n_35420, n_35421);
  not g79681 (n_35422, n47643);
  and g79682 (n47644, n_9495, n_35422);
  or g79683 (po0839, n47631, n47644);
  and g79684 (po0980, pi0953, n46888);
  and g79685 (n47647, n_34907, po0980);
  not g79686 (n_35425, po0980);
  and g79687 (n47648, pi0684, n_35425);
  not g79688 (n_35426, n47647);
  and g79689 (n47649, n_34819, n_35426);
  not g79690 (n_35427, n47648);
  and g79691 (po0841, n_35427, n47649);
  and g79692 (n47651, pi0590, n_4239);
  and g79693 (n47652, pi0357, n47651);
  and g79694 (n47653, pi0382, n47103);
  not g79695 (n_35428, n47652);
  not g79696 (n_35429, n47653);
  and g79697 (n47654, n_35428, n_35429);
  not g79698 (n_35430, n47654);
  and g79699 (n47655, n_4628, n_35430);
  and g79700 (n47656, pi0406, n_4239);
  and g79701 (n47657, n47101, n47656);
  not g79702 (n_35431, n47655);
  not g79703 (n_35432, n47657);
  and g79704 (n47658, n_35431, n_35432);
  not g79705 (n_35433, n47658);
  and g79706 (n47659, n_4832, n_35433);
  and g79707 (n47660, n_4628, n_4239);
  and g79708 (n47661, pi0588, n_4423);
  and g79709 (n47662, pi0430, n47660);
  and g79710 (n47663, n47661, n47662);
  not g79711 (n_35434, n47659);
  not g79712 (n_35435, n47663);
  and g79713 (n47664, n_35434, n_35435);
  not g79714 (n_35436, n47664);
  and g79715 (n47665, n47050, n_35436);
  not g79716 (n_35437, pi1076);
  and g79717 (n47666, pi0199, n_35437);
  not g79718 (n_35438, n47666);
  and g79719 (n47667, n_34961, n_35438);
  and g79720 (n47668, n_31955, n47667);
  not g79721 (n_35439, n47665);
  not g79722 (n_35440, n47668);
  and g79723 (n47669, n_35439, n_35440);
  not g79724 (n_35441, n47669);
  and g79725 (n47670, n7643, n_35441);
  and g79726 (n47671, pi0860, n47119);
  and g79727 (n47672, pi0744, n_2581);
  and g79728 (n47673, pi0728, pi1135);
  not g79729 (n_35445, n47672);
  and g79730 (n47674, pi1136, n_35445);
  not g79731 (n_35446, n47673);
  and g79732 (n47675, n_35446, n47674);
  not g79733 (n_35447, n47671);
  not g79734 (n_35448, n47675);
  and g79735 (n47676, n_35447, n_35448);
  not g79736 (n_35449, n47676);
  and g79737 (n47677, n47091, n_35449);
  not g79738 (n_35450, n47073);
  and g79739 (n47678, pi1136, n_35450);
  not g79740 (n_35451, n47678);
  and g79741 (n47679, n_2921, n_35451);
  and g79742 (n47680, n_34911, n_2581);
  and g79743 (n47681, pi0657, pi1135);
  not g79744 (n_35452, n47680);
  and g79745 (n47682, pi1136, n_35452);
  not g79746 (n_35453, n47681);
  and g79747 (n47683, n_35453, n47682);
  and g79748 (n47684, pi0813, n47073);
  and g79749 (n47685, n47119, n47684);
  not g79750 (n_35455, n47683);
  not g79751 (n_35456, n47685);
  and g79752 (n47686, n_35455, n_35456);
  not g79753 (n_35457, n47686);
  and g79754 (n47687, n47679, n_35457);
  not g79755 (n_35458, n47677);
  not g79756 (n_35459, n47687);
  and g79757 (n47688, n_35458, n_35459);
  not g79758 (n_35460, n47688);
  and g79759 (n47689, n_9495, n_35460);
  or g79760 (po0842, n47670, n47689);
  and g79761 (n47691, n_34737, po0980);
  and g79762 (n47692, pi0686, n_35425);
  not g79763 (n_35461, n47691);
  and g79764 (n47693, n_34819, n_35461);
  not g79765 (n_35462, n47692);
  and g79766 (po0843, n_35462, n47693);
  and g79767 (n47695, n_13620, n_35425);
  and g79768 (n47696, n_34856, po0980);
  not g79769 (n_35463, n47695);
  and g79770 (n47697, n_34819, n_35463);
  not g79771 (n_35464, n47696);
  and g79772 (po0844, n_35464, n47697);
  and g79773 (n47699, n_34753, po0980);
  and g79774 (n47700, pi0688, n_35425);
  not g79775 (n_35465, n47699);
  and g79776 (n47701, n_34819, n_35465);
  not g79777 (n_35466, n47700);
  and g79778 (po0845, n_35466, n47701);
  and g79779 (n47703, pi0351, n47651);
  and g79780 (n47704, pi0376, n47103);
  not g79781 (n_35467, n47703);
  not g79782 (n_35468, n47704);
  and g79783 (n47705, n_35467, n_35468);
  not g79784 (n_35469, n47705);
  and g79785 (n47706, n_4628, n_35469);
  and g79786 (n47707, pi0401, n_4239);
  and g79787 (n47708, n47101, n47707);
  not g79788 (n_35470, n47706);
  not g79789 (n_35471, n47708);
  and g79790 (n47709, n_35470, n_35471);
  not g79791 (n_35472, n47709);
  and g79792 (n47710, n_4832, n_35472);
  and g79793 (n47711, pi0426, n47660);
  and g79794 (n47712, n47661, n47711);
  not g79795 (n_35473, n47710);
  not g79796 (n_35474, n47712);
  and g79797 (n47713, n_35473, n_35474);
  not g79798 (n_35475, n47713);
  and g79799 (n47714, n47050, n_35475);
  not g79800 (n_35476, pi1079);
  and g79801 (n47715, pi0199, n_35476);
  and g79802 (n47716, n_7044, n42849);
  not g79803 (n_35477, n47715);
  and g79804 (n47717, n_34961, n_35477);
  not g79805 (n_35478, n47716);
  and g79806 (n47718, n_35478, n47717);
  not g79807 (n_35479, n47714);
  not g79808 (n_35480, n47718);
  and g79809 (n47719, n_35479, n_35480);
  not g79810 (n_35481, n47719);
  and g79811 (n47720, n7643, n_35481);
  and g79812 (n47721, pi0798, n47119);
  and g79813 (n47722, n_34938, n_2581);
  and g79814 (n47723, pi0655, pi1135);
  not g79815 (n_35483, n47722);
  and g79816 (n47724, pi1136, n_35483);
  not g79817 (n_35484, n47723);
  and g79818 (n47725, n_35484, n47724);
  not g79819 (n_35485, n47721);
  not g79820 (n_35486, n47725);
  and g79821 (n47726, n_35485, n_35486);
  not g79822 (n_35487, n47726);
  and g79823 (n47727, n47074, n_35487);
  and g79824 (n47728, pi0752, n47086);
  and g79825 (n47729, n_15798, pi1135);
  not g79826 (n_35489, pi0843);
  and g79827 (n47730, n_35489, n_2388);
  not g79834 (n_35493, n47727);
  not g79835 (n_35494, n47733);
  and g79836 (n47734, n_35493, n_35494);
  not g79837 (n_35495, n47734);
  and g79838 (n47735, n_9495, n_35495);
  or g79839 (po0846, n47720, n47735);
  and g79840 (n47737, n_16236, n_35425);
  and g79841 (n47738, n_34792, po0980);
  not g79842 (n_35496, n47737);
  and g79843 (n47739, n_34819, n_35496);
  not g79844 (n_35497, n47738);
  and g79845 (po0847, n_35497, n47739);
  and g79846 (n47741, n_16177, n_35425);
  and g79847 (n47742, n_34723, po0980);
  not g79848 (n_35498, n47741);
  and g79849 (n47743, n_34819, n_35498);
  not g79850 (n_35499, n47742);
  and g79851 (po0848, n_35499, n47743);
  and g79852 (n47745, pi0352, n47651);
  and g79853 (n47746, pi0317, n47103);
  not g79854 (n_35500, n47745);
  not g79855 (n_35501, n47746);
  and g79856 (n47747, n_35500, n_35501);
  not g79857 (n_35502, n47747);
  and g79858 (n47748, n_4628, n_35502);
  and g79859 (n47749, pi0402, n_4239);
  and g79860 (n47750, n47101, n47749);
  not g79861 (n_35503, n47748);
  not g79862 (n_35504, n47750);
  and g79863 (n47751, n_35503, n_35504);
  not g79864 (n_35505, n47751);
  and g79865 (n47752, n_4832, n_35505);
  and g79866 (n47753, pi0427, n47660);
  and g79867 (n47754, n47661, n47753);
  not g79868 (n_35506, n47752);
  not g79869 (n_35507, n47754);
  and g79870 (n47755, n_35506, n_35507);
  not g79871 (n_35508, n47755);
  and g79872 (n47756, n47050, n_35508);
  not g79873 (n_35509, pi1078);
  and g79874 (n47757, pi0199, n_35509);
  and g79875 (n47758, n_7044, n42861);
  not g79876 (n_35510, n47757);
  and g79877 (n47759, n_34961, n_35510);
  not g79878 (n_35511, n47758);
  and g79879 (n47760, n_35511, n47759);
  not g79880 (n_35512, n47756);
  not g79881 (n_35513, n47760);
  and g79882 (n47761, n_35512, n_35513);
  not g79883 (n_35514, n47761);
  and g79884 (n47762, n7643, n_35514);
  and g79885 (n47763, pi0844, n47119);
  and g79886 (n47764, n_14917, pi1135);
  and g79887 (n47765, pi0770, n_2581);
  not g79888 (n_35516, n47764);
  and g79889 (n47766, pi1136, n_35516);
  not g79890 (n_35517, n47765);
  and g79891 (n47767, n_35517, n47766);
  not g79892 (n_35518, n47763);
  and g79893 (n47768, pi1134, n_35518);
  not g79894 (n_35519, n47767);
  and g79895 (n47769, n_35519, n47768);
  and g79896 (n47770, pi0801, n47119);
  and g79897 (n47771, n_34931, n_2581);
  and g79898 (n47772, pi0649, pi1135);
  not g79899 (n_35521, n47771);
  and g79900 (n47773, pi1136, n_35521);
  not g79901 (n_35522, n47772);
  and g79902 (n47774, n_35522, n47773);
  not g79903 (n_35523, n47770);
  and g79904 (n47775, n_2921, n_35523);
  not g79905 (n_35524, n47774);
  and g79906 (n47776, n_35524, n47775);
  not g79907 (n_35525, n47769);
  and g79908 (n47777, n47127, n_35525);
  not g79909 (n_35526, n47776);
  and g79910 (n47778, n_35526, n47777);
  or g79911 (po0849, n47762, n47778);
  and g79912 (n47780, n_34919, po0954);
  and g79913 (n47781, pi0693, n_34817);
  not g79914 (n_35528, n47780);
  and g79915 (n47782, n_34819, n_35528);
  not g79916 (n_35529, n47781);
  and g79917 (po0850, n_35529, n47782);
  and g79918 (n47784, n_34868, po0980);
  and g79919 (n47785, pi0694, n_35425);
  not g79920 (n_35531, n47784);
  and g79921 (n47786, n_34819, n_35531);
  not g79922 (n_35532, n47785);
  and g79923 (po0851, n_35532, n47786);
  and g79924 (n47788, n_34747, po0954);
  and g79925 (n47789, pi0695, n_34817);
  not g79926 (n_35533, n47788);
  and g79927 (n47790, n_34819, n_35533);
  not g79928 (n_35534, n47789);
  and g79929 (po0852, n_35534, n47790);
  and g79930 (n47792, n_15254, n_35425);
  and g79931 (n47793, n_34686, po0980);
  not g79932 (n_35535, n47792);
  and g79933 (n47794, n_34819, n_35535);
  not g79934 (n_35536, n47793);
  and g79935 (po0853, n_35536, n47794);
  and g79936 (n47796, n_34919, po0980);
  and g79937 (n47797, pi0697, n_35425);
  not g79938 (n_35538, n47796);
  and g79939 (n47798, n_34819, n_35538);
  not g79940 (n_35539, n47797);
  and g79941 (po0854, n_35539, n47798);
  and g79942 (n47800, n_34727, po0980);
  and g79943 (n47801, pi0698, n_35425);
  not g79944 (n_35540, n47800);
  and g79945 (n47802, n_34819, n_35540);
  not g79946 (n_35541, n47801);
  and g79947 (po0855, n_35541, n47802);
  and g79948 (n47804, n_15996, n_35425);
  and g79949 (n47805, n_34874, po0980);
  not g79950 (n_35542, n47804);
  and g79951 (n47806, n_34819, n_35542);
  not g79952 (n_35543, n47805);
  and g79953 (po0856, n_35543, n47806);
  and g79954 (n47808, n_15317, n_35425);
  and g79955 (n47809, n_34845, po0980);
  not g79956 (n_35544, n47808);
  and g79957 (n47810, n_34819, n_35544);
  not g79958 (n_35545, n47809);
  and g79959 (po0857, n_35545, n47810);
  and g79960 (n47812, n_34880, po0980);
  and g79961 (n47813, pi0701, n_35425);
  not g79962 (n_35546, n47812);
  and g79963 (n47814, n_34819, n_35546);
  not g79964 (n_35547, n47813);
  and g79965 (po0858, n_35547, n47814);
  and g79966 (n47816, n_34778, po0980);
  and g79967 (n47817, pi0702, n_35425);
  not g79968 (n_35548, n47816);
  and g79969 (n47818, n_34819, n_35548);
  not g79970 (n_35549, n47817);
  and g79971 (po0859, n_35549, n47818);
  and g79972 (n47820, n_15798, n_35425);
  and g79973 (n47821, n_34926, po0980);
  not g79974 (n_35550, n47820);
  and g79975 (n47822, n_34819, n_35550);
  not g79976 (n_35551, n47821);
  and g79977 (po0860, n_35551, n47822);
  and g79978 (n47824, n_34788, po0980);
  and g79979 (n47825, pi0704, n_35425);
  not g79980 (n_35552, n47824);
  and g79981 (n47826, n_34819, n_35552);
  not g79982 (n_35553, n47825);
  and g79983 (po0861, n_35553, n47826);
  and g79984 (n47828, n_15924, n_35425);
  and g79985 (n47829, n_34886, po0980);
  not g79986 (n_35554, n47828);
  and g79987 (n47830, n_34819, n_35554);
  not g79988 (n_35555, n47829);
  and g79989 (po0862, n_35555, n47830);
  and g79990 (n47832, n_12614, n_35425);
  and g79991 (n47833, n_34769, po0980);
  not g79992 (n_35556, n47832);
  and g79993 (n47834, n_34819, n_35556);
  not g79994 (n_35557, n47833);
  and g79995 (po0863, n_35557, n47834);
  and g79996 (n47836, pi0370, n47058);
  and g79997 (n47837, pi0395, pi0591);
  and g79998 (n47838, n_4239, n47837);
  not g79999 (n_35558, n47836);
  not g80000 (n_35559, n47838);
  and g80001 (n47839, n_35558, n_35559);
  not g80002 (n_35560, n47839);
  and g80003 (n47840, n_4423, n_35560);
  and g80004 (n47841, pi0347, n47065);
  not g80005 (n_35561, n47840);
  not g80006 (n_35562, n47841);
  and g80007 (n47842, n_35561, n_35562);
  and g80008 (n47843, n_4832, n47050);
  not g80009 (n_35563, n47842);
  and g80010 (n47844, n_35563, n47843);
  not g80011 (n_35564, pi1055);
  and g80012 (n47845, pi0199, n_35564);
  not g80013 (n_35565, pi0304);
  and g80014 (n47846, n_7045, n_35565);
  and g80015 (n47847, pi0200, n_33258);
  not g80016 (n_35566, n47846);
  not g80017 (n_35567, n47847);
  and g80018 (n47848, n_35566, n_35567);
  not g80019 (n_35568, n47848);
  and g80020 (n47849, n_7044, n_35568);
  not g80021 (n_35569, n47845);
  and g80022 (n47850, n_34961, n_35569);
  not g80023 (n_35570, n47849);
  and g80024 (n47851, n_35570, n47850);
  and g80025 (n47852, n47050, n47055);
  and g80026 (n47853, pi0420, pi0588);
  and g80027 (n47854, n47852, n47853);
  not g80028 (n_35571, n47851);
  not g80029 (n_35572, n47854);
  and g80030 (n47855, n_35571, n_35572);
  not g80031 (n_35573, n47844);
  and g80032 (n47856, n_35573, n47855);
  not g80033 (n_35574, n47856);
  and g80034 (n47857, n7643, n_35574);
  and g80035 (n47858, n_11412, pi1135);
  and g80036 (n47859, n_11984, n_2581);
  and g80042 (n47863, pi0702, pi1135);
  not g80043 (n_35578, pi0847);
  and g80044 (n47864, n_35578, n_2388);
  and g80045 (n47865, pi0753, n47086);
  not g80052 (n_35582, n47862);
  not g80053 (n_35583, n47868);
  and g80054 (n47869, n_35582, n_35583);
  not g80055 (n_35584, n47869);
  and g80056 (n47870, n_9495, n_35584);
  or g80057 (po0864, n47857, n47870);
  and g80058 (n47872, n47050, n47660);
  and g80059 (n47873, pi0459, n47661);
  and g80060 (n47874, n47872, n47873);
  and g80061 (n47875, n47050, n47058);
  and g80062 (n47876, pi0442, n47875);
  and g80063 (n47877, n_4239, n47050);
  and g80064 (n47878, pi0328, pi0591);
  and g80065 (n47879, n47877, n47878);
  not g80066 (n_35585, n47876);
  not g80067 (n_35586, n47879);
  and g80068 (n47880, n_35585, n_35586);
  not g80069 (n_35587, n47880);
  and g80070 (n47881, n_4423, n_35587);
  and g80071 (n47882, pi0321, n47050);
  and g80072 (n47883, n47065, n47882);
  not g80073 (n_35588, n47881);
  not g80074 (n_35589, n47883);
  and g80075 (n47884, n_35588, n_35589);
  not g80076 (n_35590, n47884);
  and g80077 (n47885, n_4832, n_35590);
  not g80078 (n_35591, pi1058);
  and g80079 (n47886, pi0199, n_35591);
  not g80080 (n_35592, pi0305);
  and g80081 (n47887, n_7045, n_35592);
  and g80082 (n47888, pi0200, n_33268);
  not g80083 (n_35593, n47887);
  not g80084 (n_35594, n47888);
  and g80085 (n47889, n_35593, n_35594);
  not g80086 (n_35595, n47889);
  and g80087 (n47890, n_7044, n_35595);
  not g80088 (n_35596, n47886);
  and g80089 (n47891, n_34961, n_35596);
  not g80090 (n_35597, n47890);
  and g80091 (n47892, n_35597, n47891);
  and g80098 (n47896, n_11971, n_2581);
  and g80099 (n47897, n_11767, pi1135);
  and g80105 (n47901, n47073, n_34987);
  and g80106 (n47902, pi0709, pi1135);
  not g80107 (n_35604, pi0857);
  and g80108 (n47903, n_35604, n_2388);
  and g80109 (n47904, pi0754, n47086);
  not g80117 (n_35608, n47900);
  and g80118 (n47909, n_9495, n_35608);
  not g80119 (n_35609, n47908);
  and g80120 (n47910, n_35609, n47909);
  not g80121 (n_35610, n47895);
  not g80122 (n_35611, n47910);
  and g80123 (po0865, n_35610, n_35611);
  and g80124 (n47912, n_34731, po0980);
  and g80125 (n47913, pi0709, n_35425);
  not g80126 (n_35612, n47912);
  and g80127 (n47914, n_34819, n_35612);
  not g80128 (n_35613, n47913);
  and g80129 (po0866, n_35613, n47914);
  and g80130 (n47916, n_25879, n_34817);
  and g80131 (n47917, n_34800, po0954);
  not g80132 (n_35614, n47916);
  and g80133 (n47918, n_34819, n_35614);
  not g80134 (n_35615, n47917);
  and g80135 (po0867, n_35615, n47918);
  and g80136 (n47920, pi0373, n47058);
  and g80137 (n47921, pi0398, pi0591);
  and g80138 (n47922, n_4239, n47921);
  not g80139 (n_35616, n47920);
  not g80140 (n_35617, n47922);
  and g80141 (n47923, n_35616, n_35617);
  not g80142 (n_35618, n47923);
  and g80143 (n47924, n_4423, n_35618);
  and g80144 (n47925, pi0348, n47065);
  not g80145 (n_35619, n47924);
  not g80146 (n_35620, n47925);
  and g80147 (n47926, n_35619, n_35620);
  not g80148 (n_35621, n47926);
  and g80149 (n47927, n47843, n_35621);
  not g80150 (n_35622, pi1087);
  and g80151 (n47928, pi0199, n_35622);
  not g80152 (n_35623, pi0306);
  and g80153 (n47929, n_7045, n_35623);
  and g80154 (n47930, pi0200, n_33273);
  not g80155 (n_35624, n47929);
  not g80156 (n_35625, n47930);
  and g80157 (n47931, n_35624, n_35625);
  not g80158 (n_35626, n47931);
  and g80159 (n47932, n_7044, n_35626);
  not g80160 (n_35627, n47928);
  and g80161 (n47933, n_34961, n_35627);
  not g80162 (n_35628, n47932);
  and g80163 (n47934, n_35628, n47933);
  and g80164 (n47935, pi0423, pi0588);
  and g80165 (n47936, n47852, n47935);
  not g80166 (n_35629, n47934);
  not g80167 (n_35630, n47936);
  and g80168 (n47937, n_35629, n_35630);
  not g80169 (n_35631, n47927);
  and g80170 (n47938, n_35631, n47937);
  not g80171 (n_35632, n47938);
  and g80172 (n47939, n7643, n_35632);
  and g80173 (n47940, n_11806, pi1135);
  and g80174 (n47941, n_12375, n_2581);
  and g80180 (n47945, pi0725, pi1135);
  not g80181 (n_35636, pi0858);
  and g80182 (n47946, n_35636, n_2388);
  and g80183 (n47947, pi0755, n47086);
  not g80190 (n_35640, n47944);
  not g80191 (n_35641, n47950);
  and g80192 (n47951, n_35640, n_35641);
  not g80193 (n_35642, n47951);
  and g80194 (n47952, n_9495, n_35642);
  or g80195 (po0868, n47939, n47952);
  and g80196 (n47954, pi0701, pi1135);
  not g80197 (n_35644, pi0842);
  and g80198 (n47955, n_35644, n_2388);
  and g80199 (n47956, pi0751, n47086);
  and g80207 (n47961, n_12395, pi1135);
  and g80208 (n47962, n_11819, n_2581);
  not g80214 (n_35650, n47960);
  not g80215 (n_35651, n47965);
  and g80216 (n47966, n_35650, n_35651);
  not g80217 (n_35652, n47966);
  and g80218 (n47967, n_9495, n_35652);
  and g80219 (n47968, pi0199, pi1035);
  and g80220 (n47969, pi0298, n10809);
  and g80221 (n47970, pi1044, n11444);
  and g80228 (n47974, pi0425, n47660);
  and g80229 (n47975, n47661, n47974);
  and g80230 (n47976, pi0374, n47058);
  and g80231 (n47977, pi0400, pi0591);
  and g80232 (n47978, n_4239, n47977);
  not g80233 (n_35656, n47976);
  not g80234 (n_35657, n47978);
  and g80235 (n47979, n_35656, n_35657);
  not g80236 (n_35658, n47979);
  and g80237 (n47980, n_4423, n_35658);
  and g80238 (n47981, pi0350, n47065);
  not g80239 (n_35659, n47980);
  not g80240 (n_35660, n47981);
  and g80241 (n47982, n_35659, n_35660);
  not g80242 (n_35661, n47982);
  and g80243 (n47983, n_4832, n_35661);
  not g80244 (n_35662, n47975);
  and g80245 (n47984, n47050, n_35662);
  not g80246 (n_35663, n47983);
  and g80247 (n47985, n_35663, n47984);
  not g80248 (n_35664, n47973);
  and g80249 (n47986, n7643, n_35664);
  not g80250 (n_35665, n47985);
  and g80251 (n47987, n_35665, n47986);
  or g80252 (po0869, n47967, n47987);
  and g80253 (n47989, pi0371, n47058);
  and g80254 (n47990, pi0396, pi0591);
  and g80255 (n47991, n_4239, n47990);
  not g80256 (n_35666, n47989);
  not g80257 (n_35667, n47991);
  and g80258 (n47992, n_35666, n_35667);
  not g80259 (n_35668, n47992);
  and g80260 (n47993, n_4423, n_35668);
  and g80261 (n47994, pi0322, n47065);
  not g80262 (n_35669, n47993);
  not g80263 (n_35670, n47994);
  and g80264 (n47995, n_35669, n_35670);
  not g80265 (n_35671, n47995);
  and g80266 (n47996, n47843, n_35671);
  not g80267 (n_35672, pi1051);
  and g80268 (n47997, pi0199, n_35672);
  not g80269 (n_35673, pi0309);
  and g80270 (n47998, n_7045, n_35673);
  and g80271 (n47999, pi0200, n_33278);
  not g80272 (n_35674, n47998);
  not g80273 (n_35675, n47999);
  and g80274 (n48000, n_35674, n_35675);
  not g80275 (n_35676, n48000);
  and g80276 (n48001, n_7044, n_35676);
  not g80277 (n_35677, n47997);
  and g80278 (n48002, n_34961, n_35677);
  not g80279 (n_35678, n48001);
  and g80280 (n48003, n_35678, n48002);
  and g80281 (n48004, pi0421, pi0588);
  and g80282 (n48005, n47852, n48004);
  not g80283 (n_35679, n48003);
  not g80284 (n_35680, n48005);
  and g80285 (n48006, n_35679, n_35680);
  not g80286 (n_35681, n47996);
  and g80287 (n48007, n_35681, n48006);
  not g80288 (n_35682, n48007);
  and g80289 (n48008, n7643, n_35682);
  and g80290 (n48009, n_11789, pi1135);
  and g80291 (n48010, n_12354, n_2581);
  and g80297 (n48014, pi0734, pi1135);
  not g80298 (n_35686, pi0854);
  and g80299 (n48015, n_35686, n_2388);
  and g80300 (n48016, pi0756, n47086);
  not g80307 (n_35690, n48013);
  not g80308 (n_35691, n48019);
  and g80309 (n48020, n_35690, n_35691);
  not g80310 (n_35692, n48020);
  and g80311 (n48021, n_9495, n_35692);
  or g80312 (po0870, n48008, n48021);
  and g80313 (n48023, pi0461, n47651);
  and g80314 (n48024, pi0439, n47103);
  not g80315 (n_35693, n48023);
  not g80316 (n_35694, n48024);
  and g80317 (n48025, n_35693, n_35694);
  not g80318 (n_35695, n48025);
  and g80319 (n48026, n_4628, n_35695);
  and g80320 (n48027, pi0326, n_4239);
  and g80321 (n48028, n47101, n48027);
  not g80322 (n_35696, n48026);
  not g80323 (n_35697, n48028);
  and g80324 (n48029, n_35696, n_35697);
  not g80325 (n_35698, n48029);
  and g80326 (n48030, n_4832, n_35698);
  and g80327 (n48031, pi0449, n47660);
  and g80328 (n48032, n47661, n48031);
  not g80329 (n_35699, n48030);
  not g80330 (n_35700, n48032);
  and g80331 (n48033, n_35699, n_35700);
  not g80332 (n_35701, n48033);
  and g80333 (n48034, n47050, n_35701);
  not g80334 (n_35702, pi1057);
  and g80335 (n48035, pi0199, n_35702);
  not g80336 (n_35703, n48035);
  and g80337 (n48036, n_34961, n_35703);
  and g80338 (n48037, n_31534, n48036);
  not g80339 (n_35704, n48034);
  not g80340 (n_35705, n48037);
  and g80341 (n48038, n_35704, n_35705);
  not g80342 (n_35706, n48038);
  and g80343 (n48039, n7643, n_35706);
  and g80344 (n48040, pi0867, n47119);
  and g80345 (n48041, pi0762, n_2581);
  and g80346 (n48042, pi0697, pi1135);
  not g80347 (n_35709, n48041);
  and g80348 (n48043, pi1136, n_35709);
  not g80349 (n_35710, n48042);
  and g80350 (n48044, n_35710, n48043);
  not g80351 (n_35711, n48040);
  not g80352 (n_35712, n48044);
  and g80353 (n48045, n_35711, n_35712);
  not g80354 (n_35713, n48045);
  and g80355 (n48046, n47091, n_35713);
  and g80356 (n48047, n_34917, n_2581);
  and g80357 (n48048, pi0693, pi1135);
  not g80358 (n_35714, n48047);
  and g80359 (n48049, pi1136, n_35714);
  not g80360 (n_35715, n48048);
  and g80361 (n48050, n_35715, n48049);
  and g80362 (n48051, pi0816, n47073);
  and g80363 (n48052, n47119, n48051);
  not g80364 (n_35717, n48050);
  not g80365 (n_35718, n48052);
  and g80366 (n48053, n_35717, n_35718);
  not g80367 (n_35719, n48053);
  and g80368 (n48054, n47679, n_35719);
  not g80369 (n_35720, n48046);
  not g80370 (n_35721, n48054);
  and g80371 (n48055, n_35720, n_35721);
  not g80372 (n_35722, n48055);
  and g80373 (n48056, n_9495, n_35722);
  or g80374 (po0871, n48039, n48056);
  and g80375 (n48058, n_12395, n_34817);
  and g80376 (n48059, n_34880, po0954);
  not g80377 (n_35723, n48058);
  and g80378 (n48060, n_34819, n_35723);
  not g80379 (n_35724, n48059);
  and g80380 (po0872, n_35724, n48060);
  and g80381 (n48062, pi0454, n47661);
  and g80382 (n48063, n47872, n48062);
  and g80383 (n48064, pi0440, n47875);
  and g80384 (n48065, pi0329, pi0591);
  and g80385 (n48066, n47877, n48065);
  not g80386 (n_35725, n48064);
  not g80387 (n_35726, n48066);
  and g80388 (n48067, n_35725, n_35726);
  not g80389 (n_35727, n48067);
  and g80390 (n48068, n_4423, n_35727);
  and g80391 (n48069, pi0349, n47050);
  and g80392 (n48070, n47065, n48069);
  not g80393 (n_35728, n48068);
  not g80394 (n_35729, n48070);
  and g80395 (n48071, n_35728, n_35729);
  not g80396 (n_35730, n48071);
  and g80397 (n48072, n_4832, n_35730);
  not g80398 (n_35731, pi1043);
  and g80399 (n48073, pi0199, n_35731);
  not g80400 (n_35732, pi0307);
  and g80401 (n48074, n_7045, n_35732);
  and g80402 (n48075, pi0200, n_33283);
  not g80403 (n_35733, n48074);
  not g80404 (n_35734, n48075);
  and g80405 (n48076, n_35733, n_35734);
  not g80406 (n_35735, n48076);
  and g80407 (n48077, n_7044, n_35735);
  not g80408 (n_35736, n48073);
  and g80409 (n48078, n_34961, n_35736);
  not g80410 (n_35737, n48077);
  and g80411 (n48079, n_35737, n48078);
  and g80418 (n48083, n_12320, n_2581);
  and g80419 (n48084, n_11395, pi1135);
  and g80425 (n48088, pi0738, pi1135);
  not g80426 (n_35744, pi0845);
  and g80427 (n48089, n_35744, n_2388);
  and g80428 (n48090, pi0761, n47086);
  not g80436 (n_35748, n48087);
  and g80437 (n48095, n_9495, n_35748);
  not g80438 (n_35749, n48094);
  and g80439 (n48096, n_35749, n48095);
  not g80440 (n_35750, n48082);
  not g80441 (n_35751, n48096);
  and g80442 (po0873, n_35750, n_35751);
  and g80443 (n48098, pi0318, pi0591);
  and g80444 (n48099, n_4239, n48098);
  and g80445 (n48100, n_4628, n8468);
  not g80446 (n_35752, n48099);
  not g80447 (n_35753, n48100);
  and g80448 (n48101, n_35752, n_35753);
  not g80449 (n_35754, n48101);
  and g80450 (n48102, n_4423, n_35754);
  and g80451 (n48103, pi0462, n47065);
  not g80452 (n_35755, n48102);
  not g80453 (n_35756, n48103);
  and g80454 (n48104, n_35755, n_35756);
  not g80455 (n_35757, n48104);
  and g80456 (n48105, n47843, n_35757);
  not g80457 (n_35758, pi1074);
  and g80458 (n48106, pi0199, n_35758);
  and g80459 (n48107, n_7044, n42855);
  not g80460 (n_35759, n48106);
  and g80461 (n48108, n_34961, n_35759);
  not g80462 (n_35760, n48107);
  and g80463 (n48109, n_35760, n48108);
  and g80464 (n48110, pi0448, pi0588);
  and g80465 (n48111, n47852, n48110);
  not g80466 (n_35761, n48109);
  not g80467 (n_35762, n48111);
  and g80468 (n48112, n_35761, n_35762);
  not g80469 (n_35763, n48105);
  and g80470 (n48113, n_35763, n48112);
  not g80471 (n_35764, n48113);
  and g80472 (n48114, n7643, n_35764);
  and g80473 (n48115, n_15924, pi1135);
  and g80474 (n48116, pi0768, n47086);
  not g80475 (n_35766, pi0839);
  and g80476 (n48117, n_35766, n_2388);
  and g80484 (n48122, pi0800, n47119);
  and g80485 (n48123, n_34884, n_2581);
  and g80486 (n48124, pi0669, pi1135);
  not g80487 (n_35771, n48123);
  and g80488 (n48125, pi1136, n_35771);
  not g80489 (n_35772, n48124);
  and g80490 (n48126, n_35772, n48125);
  not g80491 (n_35773, n48122);
  not g80492 (n_35774, n48126);
  and g80493 (n48127, n_35773, n_35774);
  not g80494 (n_35775, n48127);
  and g80495 (n48128, n47074, n_35775);
  not g80496 (n_35776, n48121);
  not g80497 (n_35777, n48128);
  and g80498 (n48129, n_35776, n_35777);
  not g80499 (n_35778, n48129);
  and g80500 (n48130, n_9495, n_35778);
  or g80501 (po0874, n48114, n48130);
  and g80502 (n48132, pi0419, n47661);
  and g80503 (n48133, n47872, n48132);
  and g80504 (n48134, pi0369, n47875);
  and g80505 (n48135, pi0394, pi0591);
  and g80506 (n48136, n47877, n48135);
  not g80507 (n_35779, n48134);
  not g80508 (n_35780, n48136);
  and g80509 (n48137, n_35779, n_35780);
  not g80510 (n_35781, n48137);
  and g80511 (n48138, n_4423, n_35781);
  and g80512 (n48139, pi0315, n47050);
  and g80513 (n48140, n47065, n48139);
  not g80514 (n_35782, n48138);
  not g80515 (n_35783, n48140);
  and g80516 (n48141, n_35782, n_35783);
  not g80517 (n_35784, n48141);
  and g80518 (n48142, n_4832, n_35784);
  not g80519 (n_35785, pi1080);
  and g80520 (n48143, pi0199, n_35785);
  not g80521 (n_35786, pi0303);
  and g80522 (n48144, n_7045, n_35786);
  and g80523 (n48145, pi0200, n_33263);
  not g80524 (n_35787, n48144);
  not g80525 (n_35788, n48145);
  and g80526 (n48146, n_35787, n_35788);
  not g80527 (n_35789, n48146);
  and g80528 (n48147, n_7044, n_35789);
  not g80529 (n_35790, n48143);
  and g80530 (n48148, n_34961, n_35790);
  not g80531 (n_35791, n48147);
  and g80532 (n48149, n_35791, n48148);
  and g80539 (n48153, n_11823, n_2581);
  and g80540 (n48154, n_11753, pi1135);
  and g80546 (n48158, pi0698, pi1135);
  not g80547 (n_35798, pi0853);
  and g80548 (n48159, n_35798, n_2388);
  and g80549 (n48160, pi0767, n47086);
  not g80557 (n_35802, n48157);
  and g80558 (n48165, n_9495, n_35802);
  not g80559 (n_35803, n48164);
  and g80560 (n48166, n_35803, n48165);
  not g80561 (n_35804, n48152);
  not g80562 (n_35805, n48166);
  and g80563 (po0875, n_35804, n_35805);
  and g80564 (n48168, pi0378, n47058);
  and g80565 (n48169, pi0325, pi0591);
  and g80566 (n48170, n_4239, n48169);
  not g80567 (n_35806, n48168);
  not g80568 (n_35807, n48170);
  and g80569 (n48171, n_35806, n_35807);
  not g80570 (n_35808, n48171);
  and g80571 (n48172, n_4423, n_35808);
  and g80572 (n48173, pi0353, n47065);
  not g80573 (n_35809, n48172);
  not g80574 (n_35810, n48173);
  and g80575 (n48174, n_35809, n_35810);
  not g80576 (n_35811, n48174);
  and g80577 (n48175, n47843, n_35811);
  not g80578 (n_35812, pi1063);
  and g80579 (n48176, pi0199, n_35812);
  and g80580 (n48177, n_7044, n42867);
  not g80581 (n_35813, n48176);
  and g80582 (n48178, n_34961, n_35813);
  not g80583 (n_35814, n48177);
  and g80584 (n48179, n_35814, n48178);
  and g80585 (n48180, pi0451, pi0588);
  and g80586 (n48181, n47852, n48180);
  not g80587 (n_35815, n48179);
  not g80588 (n_35816, n48181);
  and g80589 (n48182, n_35815, n_35816);
  not g80590 (n_35817, n48175);
  and g80591 (n48183, n_35817, n48182);
  not g80592 (n_35818, n48183);
  and g80593 (n48184, n7643, n_35818);
  and g80594 (n48185, n_13620, pi1135);
  and g80595 (n48186, pi0774, n47086);
  not g80596 (n_35820, pi0868);
  and g80597 (n48187, n_35820, n_2388);
  and g80605 (n48192, pi0807, n47119);
  and g80606 (n48193, n_34854, n_2581);
  and g80607 (n48194, pi0650, pi1135);
  not g80608 (n_35825, n48193);
  and g80609 (n48195, pi1136, n_35825);
  not g80610 (n_35826, n48194);
  and g80611 (n48196, n_35826, n48195);
  not g80612 (n_35827, n48192);
  not g80613 (n_35828, n48196);
  and g80614 (n48197, n_35827, n_35828);
  not g80615 (n_35829, n48197);
  and g80616 (n48198, n47074, n_35829);
  not g80617 (n_35830, n48191);
  not g80618 (n_35831, n48198);
  and g80619 (n48199, n_35830, n_35831);
  not g80620 (n_35832, n48199);
  and g80621 (n48200, n_9495, n_35832);
  or g80622 (po0876, n48184, n48200);
  and g80623 (n48202, pi0356, n47651);
  and g80624 (n48203, pi0381, n47103);
  not g80625 (n_35833, n48202);
  not g80626 (n_35834, n48203);
  and g80627 (n48204, n_35833, n_35834);
  not g80628 (n_35835, n48204);
  and g80629 (n48205, n_4628, n_35835);
  and g80630 (n48206, pi0405, n_4239);
  and g80631 (n48207, n47101, n48206);
  not g80632 (n_35836, n48205);
  not g80633 (n_35837, n48207);
  and g80634 (n48208, n_35836, n_35837);
  not g80635 (n_35838, n48208);
  and g80636 (n48209, n_4832, n_35838);
  and g80637 (n48210, pi0445, n47660);
  and g80638 (n48211, n47661, n48210);
  not g80639 (n_35839, n48209);
  not g80640 (n_35840, n48211);
  and g80641 (n48212, n_35839, n_35840);
  not g80642 (n_35841, n48212);
  and g80643 (n48213, n47050, n_35841);
  not g80644 (n_35842, pi1081);
  and g80645 (n48214, pi0199, n_35842);
  not g80646 (n_35843, n48214);
  and g80647 (n48215, n_34961, n_35843);
  and g80648 (n48216, n_31961, n48215);
  not g80649 (n_35844, n48213);
  not g80650 (n_35845, n48216);
  and g80651 (n48217, n_35844, n_35845);
  not g80652 (n_35846, n48217);
  and g80653 (n48218, n7643, n_35846);
  and g80654 (n48219, pi0880, n47119);
  and g80655 (n48220, pi0750, n_2581);
  and g80656 (n48221, pi0684, pi1135);
  not g80657 (n_35849, n48220);
  and g80658 (n48222, pi1136, n_35849);
  not g80659 (n_35850, n48221);
  and g80660 (n48223, n_35850, n48222);
  not g80661 (n_35851, n48219);
  not g80662 (n_35852, n48223);
  and g80663 (n48224, n_35851, n_35852);
  not g80664 (n_35853, n48224);
  and g80665 (n48225, n47091, n_35853);
  and g80666 (n48226, n_34905, n_2581);
  and g80667 (n48227, pi0654, pi1135);
  not g80668 (n_35854, n48226);
  and g80669 (n48228, pi1136, n_35854);
  not g80670 (n_35855, n48227);
  and g80671 (n48229, n_35855, n48228);
  and g80672 (n48230, pi0794, n47073);
  and g80673 (n48231, n47119, n48230);
  not g80674 (n_35857, n48229);
  not g80675 (n_35858, n48231);
  and g80676 (n48232, n_35857, n_35858);
  not g80677 (n_35859, n48232);
  and g80678 (n48233, n47679, n_35859);
  not g80679 (n_35860, n48225);
  not g80680 (n_35861, n48233);
  and g80681 (n48234, n_35860, n_35861);
  not g80682 (n_35862, n48234);
  and g80683 (n48235, n_9495, n_35862);
  or g80684 (po0877, n48218, n48235);
  not g80685 (n_35865, pi0775);
  and g80686 (n48237, pi0721, n_35865);
  and g80687 (n48238, pi0721, pi0813);
  not g80688 (n_35867, pi0773);
  not g80689 (n_35868, pi0801);
  and g80690 (n48239, n_35867, n_35868);
  and g80691 (n48240, pi0773, pi0801);
  not g80692 (n_35869, n48239);
  not g80693 (n_35870, n48240);
  and g80694 (n48241, n_35869, n_35870);
  not g80695 (n_35872, pi0771);
  not g80696 (n_35873, pi0800);
  and g80697 (n48242, n_35872, n_35873);
  and g80698 (n48243, pi0771, pi0800);
  not g80699 (n_35874, n48242);
  not g80700 (n_35875, n48243);
  and g80701 (n48244, n_35874, n_35875);
  not g80702 (n_35877, pi0769);
  not g80703 (n_35878, pi0794);
  and g80704 (n48245, n_35877, n_35878);
  and g80705 (n48246, pi0769, pi0794);
  not g80706 (n_35879, n48245);
  not g80707 (n_35880, n48246);
  and g80708 (n48247, n_35879, n_35880);
  not g80709 (n_35882, pi0765);
  not g80710 (n_35883, pi0798);
  and g80711 (n48248, n_35882, n_35883);
  and g80712 (n48249, pi0765, pi0798);
  not g80713 (n_35884, n48248);
  not g80714 (n_35885, n48249);
  and g80715 (n48250, n_35884, n_35885);
  not g80716 (n_35886, n48250);
  and g80717 (n48251, pi0807, n_35886);
  and g80718 (n48252, pi0747, n48251);
  not g80719 (n_35888, pi0747);
  not g80720 (n_35889, pi0807);
  and g80721 (n48253, n_35888, n_35889);
  and g80722 (n48254, n_35886, n48253);
  not g80723 (n_35890, n48252);
  not g80724 (n_35891, n48254);
  and g80725 (n48255, n_35890, n_35891);
  not g80726 (n_35892, n48247);
  not g80727 (n_35893, n48255);
  and g80728 (n48256, n_35892, n_35893);
  not g80729 (n_35894, n48244);
  and g80730 (n48257, n_35894, n48256);
  not g80731 (n_35895, n48241);
  and g80732 (n48258, n_35895, n48257);
  and g80733 (n48259, n48238, n48258);
  not g80734 (n_35896, pi0816);
  and g80735 (n48260, n_35865, n_35896);
  and g80736 (n48261, pi0775, pi0816);
  not g80737 (n_35897, n48260);
  not g80738 (n_35898, n48261);
  and g80739 (n48262, n_35897, n_35898);
  not g80740 (n_35899, n48262);
  and g80741 (n48263, n48259, n_35899);
  not g80742 (n_35900, n48263);
  and g80743 (n48264, n48237, n_35900);
  and g80744 (n48265, pi0747, pi0773);
  and g80745 (n48266, pi0769, n48265);
  and g80746 (n48267, pi0721, n48266);
  not g80747 (n_35901, pi0721);
  not g80748 (n_35902, n48266);
  and g80749 (n48268, n_35901, n_35902);
  not g80750 (n_35903, n48267);
  and g80751 (n48269, pi0775, n_35903);
  not g80752 (n_35904, n48268);
  and g80753 (n48270, n_35904, n48269);
  and g80754 (n48271, n_35894, n48251);
  not g80755 (n_35905, pi0813);
  and g80756 (n48272, n_35901, n_35905);
  not g80760 (n_35906, n48259);
  not g80761 (n_35907, n48275);
  and g80762 (n48276, n_35906, n_35907);
  not g80763 (n_35908, n48276);
  and g80764 (n48277, pi0816, n_35908);
  not g80765 (n_35909, n48277);
  and g80766 (n48278, n48270, n_35909);
  not g80767 (n_35911, n48278);
  and g80768 (n48279, pi0795, n_35911);
  not g80769 (n_35913, pi0945);
  and g80770 (n48280, n_35913, pi0988);
  and g80771 (n48281, pi0731, n48280);
  not g80772 (n_35916, n48237);
  not g80773 (n_35917, n48270);
  and g80774 (n48282, n_35916, n_35917);
  not g80775 (n_35918, n48282);
  and g80776 (n48283, n48281, n_35918);
  not g80777 (n_35919, n48279);
  and g80778 (n48284, n_35919, n48283);
  not g80779 (n_35920, pi0731);
  not g80780 (n_35921, pi0795);
  and g80781 (n48285, n_35920, n_35921);
  and g80782 (n48286, pi0731, pi0795);
  not g80783 (n_35922, n48285);
  not g80784 (n_35923, n48286);
  and g80785 (n48287, n_35922, n_35923);
  not g80786 (n_35924, n48287);
  and g80787 (n48288, n48263, n_35924);
  not g80788 (n_35925, n48281);
  and g80789 (n48289, pi0721, n_35925);
  not g80790 (n_35926, n48288);
  and g80791 (n48290, n_35926, n48289);
  not g80792 (n_35927, n48264);
  not g80793 (n_35928, n48290);
  and g80794 (n48291, n_35927, n_35928);
  not g80795 (n_35929, n48291);
  or g80796 (po0878, n48284, n_35929);
  and g80797 (n48293, pi0379, n47058);
  and g80798 (n48294, pi0403, pi0591);
  and g80799 (n48295, n_4239, n48294);
  not g80800 (n_35930, n48293);
  not g80801 (n_35931, n48295);
  and g80802 (n48296, n_35930, n_35931);
  not g80803 (n_35932, n48296);
  and g80804 (n48297, n_4423, n_35932);
  and g80805 (n48298, pi0354, n47065);
  not g80806 (n_35933, n48297);
  not g80807 (n_35934, n48298);
  and g80808 (n48299, n_35933, n_35934);
  not g80809 (n_35935, n48299);
  and g80810 (n48300, n47843, n_35935);
  not g80811 (n_35936, pi1045);
  and g80812 (n48301, pi0199, n_35936);
  and g80813 (n48302, n_7044, n42873);
  not g80814 (n_35937, n48301);
  and g80815 (n48303, n_34961, n_35937);
  not g80816 (n_35938, n48302);
  and g80817 (n48304, n_35938, n48303);
  and g80818 (n48305, pi0428, pi0588);
  and g80819 (n48306, n47852, n48305);
  not g80820 (n_35939, n48304);
  not g80821 (n_35940, n48306);
  and g80822 (n48307, n_35939, n_35940);
  not g80823 (n_35941, n48300);
  and g80824 (n48308, n_35941, n48307);
  not g80825 (n_35942, n48308);
  and g80826 (n48309, n7643, n_35942);
  and g80827 (n48310, n_35921, n_2921);
  not g80828 (n_35944, pi0851);
  and g80829 (n48311, n_35944, pi1134);
  not g80830 (n_35945, n48310);
  and g80831 (n48312, n_2388, n_35945);
  not g80832 (n_35946, n48311);
  and g80833 (n48313, n_35946, n48312);
  and g80834 (n48314, n_34866, n_2921);
  and g80835 (n48315, pi0776, pi1134);
  not g80836 (n_35948, n48314);
  and g80837 (n48316, pi1136, n_35948);
  not g80838 (n_35949, n48315);
  and g80839 (n48317, n_35949, n48316);
  not g80840 (n_35950, n48313);
  not g80841 (n_35951, n48317);
  and g80842 (n48318, n_35950, n_35951);
  not g80843 (n_35952, n48318);
  and g80844 (n48319, n_2581, n_35952);
  and g80845 (n48320, pi0694, pi1134);
  and g80846 (n48321, pi0732, n_2921);
  not g80852 (n_35956, n48319);
  not g80853 (n_35957, n48324);
  and g80854 (n48325, n_35956, n_35957);
  not g80855 (n_35958, n48325);
  and g80856 (n48326, n47127, n_35958);
  or g80857 (po0879, n48309, n48326);
  and g80858 (n48328, n_34747, po0980);
  and g80859 (n48329, pi0723, n_35425);
  not g80860 (n_35959, n48328);
  and g80861 (n48330, n_34819, n_35959);
  not g80862 (n_35960, n48329);
  and g80863 (po0880, n_35960, n48330);
  and g80864 (n48332, n_34743, po0980);
  and g80865 (n48333, pi0724, n_35425);
  not g80866 (n_35961, n48332);
  and g80867 (n48334, n_34819, n_35961);
  not g80868 (n_35962, n48333);
  and g80869 (po0881, n_35962, n48334);
  and g80870 (n48336, n_34835, po0980);
  and g80871 (n48337, pi0725, n_35425);
  not g80872 (n_35963, n48336);
  and g80873 (n48338, n_34819, n_35963);
  not g80874 (n_35964, n48337);
  and g80875 (po0882, n_35964, n48338);
  and g80876 (n48340, n_14917, n_35425);
  and g80877 (n48341, n_34897, po0980);
  not g80878 (n_35965, n48340);
  and g80879 (n48342, n_34819, n_35965);
  not g80880 (n_35966, n48341);
  and g80881 (po0883, n_35966, n48342);
  and g80882 (n48344, n_15870, n_35425);
  and g80883 (n48345, n_34757, po0980);
  not g80884 (n_35967, n48344);
  and g80885 (n48346, n_34819, n_35967);
  not g80886 (n_35968, n48345);
  and g80887 (po0884, n_35968, n48346);
  and g80888 (n48348, n_34913, po0980);
  and g80889 (n48349, pi0728, n_35425);
  not g80890 (n_35969, n48348);
  and g80891 (n48350, n_34819, n_35969);
  not g80892 (n_35970, n48349);
  and g80893 (po0885, n_35970, n48350);
  and g80894 (n48352, n_16056, n_35425);
  and g80895 (n48353, n_34714, po0980);
  not g80896 (n_35971, n48352);
  and g80897 (n48354, n_34819, n_35971);
  not g80898 (n_35972, n48353);
  and g80899 (po0886, n_35972, n48354);
  and g80900 (n48356, n_16117, n_35425);
  and g80901 (n48357, n_34800, po0980);
  not g80902 (n_35973, n48356);
  and g80903 (n48358, n_34819, n_35973);
  not g80904 (n_35974, n48357);
  and g80905 (po0887, n_35974, n48358);
  not g80906 (n_35975, n48238);
  not g80907 (n_35976, n48272);
  and g80908 (n48360, n_35975, n_35976);
  not g80909 (n_35977, n48360);
  and g80910 (n48361, n48258, n_35977);
  and g80911 (n48362, pi0795, n_35899);
  and g80912 (n48363, n48361, n48362);
  not g80913 (n_35978, n48265);
  not g80914 (n_35979, n48363);
  and g80915 (n48364, n_35978, n_35979);
  not g80916 (n_35980, n48364);
  and g80917 (n48365, n48281, n_35980);
  and g80918 (n48366, pi0731, n_35979);
  and g80919 (n48367, n_35899, n_35977);
  not g80924 (n_35981, n48371);
  and g80925 (n48372, n48265, n_35981);
  not g80926 (n_35982, n48372);
  and g80927 (n48373, n_35920, n_35982);
  not g80928 (n_35983, n48373);
  and g80929 (n48374, n48280, n_35983);
  not g80930 (n_35984, n48366);
  not g80931 (n_35985, n48374);
  and g80932 (n48375, n_35984, n_35985);
  not g80933 (n_35986, n48365);
  not g80934 (n_35987, n48375);
  and g80935 (po0888, n_35986, n_35987);
  and g80936 (n48377, n_34868, po0954);
  and g80937 (n48378, pi0732, n_34817);
  not g80938 (n_35988, n48377);
  and g80939 (n48379, n_34819, n_35988);
  not g80940 (n_35989, n48378);
  and g80941 (po0889, n_35989, n48379);
  and g80942 (n48381, pi0424, n47661);
  and g80943 (n48382, n47872, n48381);
  and g80944 (n48383, pi0375, n47875);
  and g80945 (n48384, pi0399, pi0591);
  and g80946 (n48385, n47877, n48384);
  not g80947 (n_35990, n48383);
  not g80948 (n_35991, n48385);
  and g80949 (n48386, n_35990, n_35991);
  not g80950 (n_35992, n48386);
  and g80951 (n48387, n_4423, n_35992);
  and g80952 (n48388, pi0316, n47050);
  and g80953 (n48389, n47065, n48388);
  not g80954 (n_35993, n48387);
  not g80955 (n_35994, n48389);
  and g80956 (n48390, n_35993, n_35994);
  not g80957 (n_35995, n48390);
  and g80958 (n48391, n_4832, n_35995);
  not g80959 (n_35996, pi1047);
  and g80960 (n48392, pi0199, n_35996);
  not g80961 (n_35997, pi0308);
  and g80962 (n48393, n_7045, n_35997);
  and g80963 (n48394, pi0200, n_33288);
  not g80964 (n_35998, n48393);
  not g80965 (n_35999, n48394);
  and g80966 (n48395, n_35998, n_35999);
  not g80967 (n_36000, n48395);
  and g80968 (n48396, n_7044, n_36000);
  not g80969 (n_36001, n48392);
  and g80970 (n48397, n_34961, n_36001);
  not g80971 (n_36002, n48396);
  and g80972 (n48398, n_36002, n48397);
  and g80979 (n48402, n_11821, n_2581);
  and g80980 (n48403, n_11403, pi1135);
  and g80986 (n48407, pi0737, pi1135);
  not g80987 (n_36009, pi0838);
  and g80988 (n48408, n_36009, n_2388);
  and g80989 (n48409, pi0777, n47086);
  not g80997 (n_36013, n48406);
  and g80998 (n48414, n_9495, n_36013);
  not g80999 (n_36014, n48413);
  and g81000 (n48415, n_36014, n48414);
  not g81001 (n_36015, n48401);
  not g81002 (n_36016, n48415);
  and g81003 (po0890, n_36015, n_36016);
  and g81004 (n48417, n_34829, po0980);
  and g81005 (n48418, pi0734, n_35425);
  not g81006 (n_36017, n48417);
  and g81007 (n48419, n_34819, n_36017);
  not g81008 (n_36018, n48418);
  and g81009 (po0891, n_36018, n48419);
  and g81010 (n48421, n_13045, n_35425);
  and g81011 (n48422, n_34796, po0980);
  not g81012 (n_36019, n48421);
  and g81013 (n48423, n_34819, n_36019);
  not g81014 (n_36020, n48422);
  and g81015 (po0892, n_36020, n48423);
  and g81016 (n48425, n_14126, n_35425);
  and g81017 (n48426, n_34765, po0980);
  not g81018 (n_36021, n48425);
  and g81019 (n48427, n_34819, n_36021);
  not g81020 (n_36022, n48426);
  and g81021 (po0893, n_36022, n48427);
  and g81022 (n48429, n_34782, po0980);
  and g81023 (n48430, pi0737, n_35425);
  not g81024 (n_36023, n48429);
  and g81025 (n48431, n_34819, n_36023);
  not g81026 (n_36024, n48430);
  and g81027 (po0894, n_36024, n48431);
  and g81028 (n48433, n_34823, po0980);
  and g81029 (n48434, pi0738, n_35425);
  not g81030 (n_36025, n48433);
  and g81031 (n48435, n_34819, n_36025);
  not g81032 (n_36026, n48434);
  and g81033 (po0895, n_36026, n48435);
  not g81034 (n_36027, pi0952);
  and g81035 (n48437, n_36027, n_34693);
  and g81036 (n48438, n46780, n48437);
  and g81037 (po0988, pi0832, n48438);
  and g81038 (n48440, pi1108, po0988);
  not g81039 (n_36029, po0988);
  and g81040 (n48441, pi0739, n_36029);
  not g81041 (n_36030, n48440);
  and g81042 (n48442, n_34696, n_36030);
  not g81043 (n_36031, n48442);
  or g81044 (po0896, n48441, n_36031);
  and g81045 (n48444, n_15412, n_36029);
  and g81046 (n48445, pi1114, po0988);
  not g81047 (n_36032, n48444);
  and g81048 (n48446, n_34696, n_36032);
  not g81049 (n_36033, n48446);
  or g81050 (po0898, n48445, n_36033);
  and g81051 (n48448, n_15327, n_36029);
  and g81052 (n48449, pi1112, po0988);
  not g81053 (n_36034, n48448);
  and g81054 (n48450, n_34696, n_36034);
  not g81055 (n_36035, n48450);
  or g81056 (po0899, n48449, n_36035);
  and g81057 (n48452, pi1109, po0988);
  and g81058 (n48453, pi0743, n_36029);
  not g81059 (n_36036, n48452);
  and g81060 (n48454, n_34696, n_36036);
  not g81061 (n_36037, n48454);
  or g81062 (po0900, n48453, n_36037);
  not g81063 (n_36038, pi0744);
  and g81064 (n48456, n_36038, n_36029);
  and g81065 (n48457, pi1131, po0988);
  not g81066 (n_36039, n48456);
  and g81067 (n48458, n_34696, n_36039);
  not g81068 (n_36040, n48458);
  or g81069 (po0901, n48457, n_36040);
  and g81070 (n48460, n_15125, n_36029);
  and g81071 (n48461, pi1111, po0988);
  not g81072 (n_36041, n48460);
  and g81073 (n48462, n_34696, n_36041);
  not g81074 (n_36042, n48462);
  or g81075 (po0902, n48461, n_36042);
  and g81076 (n48464, pi1104, po0988);
  and g81077 (n48465, pi0746, n_36029);
  not g81078 (n_36043, n48464);
  and g81079 (n48466, n_34696, n_36043);
  not g81080 (n_36044, n48466);
  or g81081 (po0903, n48465, n_36044);
  and g81082 (n48468, pi0773, n48280);
  not g81083 (n_36045, n48468);
  and g81084 (n48469, n_35888, n_36045);
  and g81085 (n48470, n48265, n48280);
  and g81086 (n48471, n_35924, n48367);
  and g81087 (n48472, pi0801, n48254);
  and g81088 (n48473, n_35895, n_36045);
  and g81089 (n48474, n48251, n48473);
  not g81090 (n_36046, n48472);
  not g81091 (n_36047, n48474);
  and g81092 (n48475, n_36046, n_36047);
  not g81097 (n_36049, n48469);
  not g81098 (n_36050, n48470);
  and g81099 (n48479, n_36049, n_36050);
  not g81100 (n_36051, n48478);
  and g81101 (po0904, n_36051, n48479);
  and g81102 (n48481, pi1106, po0988);
  and g81103 (n48482, pi0748, n_36029);
  not g81104 (n_36052, n48481);
  and g81105 (n48483, n_34696, n_36052);
  not g81106 (n_36053, n48483);
  or g81107 (po0905, n48482, n_36053);
  and g81108 (n48485, pi1105, po0988);
  and g81109 (n48486, pi0749, n_36029);
  not g81110 (n_36054, n48485);
  and g81111 (n48487, n_34696, n_36054);
  not g81112 (n_36055, n48487);
  or g81113 (po0906, n48486, n_36055);
  not g81114 (n_36056, pi0750);
  and g81115 (n48489, n_36056, n_36029);
  and g81116 (n48490, pi1130, po0988);
  not g81117 (n_36057, n48489);
  and g81118 (n48491, n_34696, n_36057);
  not g81119 (n_36058, n48491);
  or g81120 (po0907, n48490, n_36058);
  and g81121 (n48493, n_15080, n_36029);
  and g81122 (n48494, pi1123, po0988);
  not g81123 (n_36059, n48493);
  and g81124 (n48495, n_34696, n_36059);
  not g81125 (n_36060, n48495);
  or g81126 (po0908, n48494, n_36060);
  and g81127 (n48497, n_15776, n_36029);
  and g81128 (n48498, pi1124, po0988);
  not g81129 (n_36061, n48497);
  and g81130 (n48499, n_34696, n_36061);
  not g81131 (n_36062, n48499);
  or g81132 (po0909, n48498, n_36062);
  and g81133 (n48501, n_15488, n_36029);
  and g81134 (n48502, pi1117, po0988);
  not g81135 (n_36063, n48501);
  and g81136 (n48503, n_34696, n_36063);
  not g81137 (n_36064, n48503);
  or g81138 (po0910, n48502, n_36064);
  and g81139 (n48505, n_15533, n_36029);
  and g81140 (n48506, pi1118, po0988);
  not g81141 (n_36065, n48505);
  and g81142 (n48507, n_34696, n_36065);
  not g81143 (n_36066, n48507);
  or g81144 (po0911, n48506, n_36066);
  and g81145 (n48509, n_15034, n_36029);
  and g81146 (n48510, pi1120, po0988);
  not g81147 (n_36067, n48509);
  and g81148 (n48511, n_34696, n_36067);
  not g81149 (n_36068, n48511);
  or g81150 (po0912, n48510, n_36068);
  and g81151 (n48513, n_15578, n_36029);
  and g81152 (n48514, pi1119, po0988);
  not g81153 (n_36069, n48513);
  and g81154 (n48515, n_34696, n_36069);
  not g81155 (n_36070, n48515);
  or g81156 (po0913, n48514, n_36070);
  and g81157 (n48517, n_15373, n_36029);
  and g81158 (n48518, pi1113, po0988);
  not g81159 (n_36071, n48517);
  and g81160 (n48519, n_34696, n_36071);
  not g81161 (n_36072, n48519);
  or g81162 (po0914, n48518, n_36072);
  and g81163 (n48521, pi1101, po0988);
  and g81164 (n48522, pi0758, n_36029);
  not g81165 (n_36073, n48521);
  and g81166 (n48523, n_34696, n_36073);
  not g81167 (n_36074, n48523);
  or g81168 (po0915, n48522, n_36074);
  and g81169 (n48525, n_15215, n_36029);
  and g81170 (n48526, n46778, n48438);
  not g81171 (n_36075, n48525);
  not g81172 (n_36076, n48526);
  and g81173 (n48527, n_36075, n_36076);
  or g81174 (po0916, pi0966, n48527);
  and g81175 (n48529, n_15442, n_36029);
  and g81176 (n48530, pi1115, po0988);
  not g81177 (n_36077, n48529);
  and g81178 (n48531, n_34696, n_36077);
  not g81179 (n_36078, n48531);
  or g81180 (po0917, n48530, n_36078);
  and g81181 (n48533, n_11912, n_36029);
  and g81182 (n48534, pi1121, po0988);
  not g81183 (n_36079, n48533);
  and g81184 (n48535, n_34696, n_36079);
  not g81185 (n_36080, n48535);
  or g81186 (po0918, n48534, n_36080);
  not g81187 (n_36081, pi0762);
  and g81188 (n48537, n_36081, n_36029);
  and g81189 (n48538, pi1129, po0988);
  not g81190 (n_36082, n48537);
  and g81191 (n48539, n_34696, n_36082);
  not g81192 (n_36083, n48539);
  or g81193 (po0919, n48538, n_36083);
  and g81194 (n48541, pi1103, po0988);
  and g81195 (n48542, pi0763, n_36029);
  not g81196 (n_36084, n48541);
  and g81197 (n48543, n_34696, n_36084);
  not g81198 (n_36085, n48543);
  or g81199 (po0920, n48542, n_36085);
  and g81200 (n48545, pi1107, po0988);
  and g81201 (n48546, pi0764, n_36029);
  not g81202 (n_36086, n48545);
  and g81203 (n48547, n_34696, n_36086);
  not g81204 (n_36087, n48547);
  or g81205 (po0921, n48546, n_36087);
  and g81206 (po0978, n48258, n48471);
  not g81207 (n_36089, po0978);
  and g81208 (n48550, pi0765, n_36089);
  not g81209 (n_36090, n48550);
  and g81210 (n48551, pi0945, n_36090);
  and g81211 (n48552, n_35906, n_35976);
  not g81215 (n_36091, n48555);
  and g81216 (n48556, n48239, n_36091);
  not g81217 (n_36092, n48556);
  and g81218 (n48557, n_35870, n_36092);
  not g81219 (n_36093, n48557);
  and g81220 (n48558, n48257, n_36093);
  not g81221 (n_36094, n48558);
  and g81222 (n48559, n_35901, n_36094);
  not g81223 (n_36095, n48559);
  and g81224 (n48560, n48260, n_36095);
  not g81225 (n_36096, n48552);
  and g81226 (n48561, n_36096, n48560);
  and g81227 (n48562, n48261, n48361);
  not g81228 (n_36097, n48562);
  and g81229 (n48563, n_35882, n_36097);
  not g81230 (n_36098, n48561);
  and g81231 (n48564, n_36098, n48563);
  not g81232 (n_36099, n48564);
  and g81233 (n48565, n_35921, n_36099);
  not g81234 (n_36100, n48565);
  and g81235 (n48566, n_35920, n_36100);
  and g81236 (n48567, n_35921, n48566);
  not g81237 (n_36101, n48567);
  and g81238 (n48568, pi0765, n_36101);
  not g81239 (n_36102, n48566);
  and g81240 (n48569, n_35984, n_36102);
  not g81241 (n_36103, n48568);
  not g81242 (n_36104, n48569);
  and g81243 (n48570, n_36103, n_36104);
  not g81244 (n_36105, n48570);
  and g81245 (n48571, n_35913, n_36105);
  not g81246 (n_36106, n48551);
  not g81247 (n_36107, n48571);
  and g81248 (po0922, n_36106, n_36107);
  and g81249 (n48573, pi1110, po0988);
  and g81250 (n48574, pi0766, n_36029);
  not g81251 (n_36108, n48573);
  and g81252 (n48575, n_34696, n_36108);
  not g81253 (n_36109, n48575);
  or g81254 (po0923, n48574, n_36109);
  and g81255 (n48577, n_14479, n_36029);
  and g81256 (n48578, pi1116, po0988);
  not g81257 (n_36110, n48577);
  and g81258 (n48579, n_34696, n_36110);
  not g81259 (n_36111, n48579);
  or g81260 (po0924, n48578, n_36111);
  and g81261 (n48581, n_15911, n_36029);
  and g81262 (n48582, pi1125, po0988);
  not g81263 (n_36112, n48581);
  and g81264 (n48583, n_34696, n_36112);
  not g81265 (n_36113, n48583);
  or g81266 (po0925, n48582, n_36113);
  and g81271 (n48589, n_35865, n48588);
  not g81272 (n_36114, n48589);
  and g81273 (n48590, n_36097, n_36114);
  not g81274 (n_36115, n48590);
  and g81275 (n48591, pi0795, n_36115);
  and g81276 (n48592, pi0775, n48265);
  not g81277 (n_36116, n48592);
  and g81278 (n48593, pi0769, n_36116);
  and g81279 (n48594, n_35877, n48592);
  not g81280 (n_36117, n48593);
  not g81281 (n_36118, n48594);
  and g81282 (n48595, n_36117, n_36118);
  not g81283 (n_36119, n48595);
  and g81284 (n48596, n48281, n_36119);
  not g81285 (n_36120, n48591);
  and g81286 (n48597, n_36120, n48596);
  and g81287 (n48598, n_35924, n48588);
  and g81288 (n48599, pi0769, n_35925);
  not g81289 (n_36121, n48598);
  and g81290 (n48600, n_36121, n48599);
  or g81291 (po0926, n48597, n48600);
  and g81292 (n48602, n_14875, n_36029);
  and g81293 (n48603, pi1126, po0988);
  not g81294 (n_36122, n48602);
  and g81295 (n48604, n_34696, n_36122);
  not g81296 (n_36123, n48604);
  or g81297 (po0927, n48603, n_36123);
  not g81298 (n_36124, n48560);
  and g81299 (n48606, n_35898, n_36124);
  not g81300 (n_36125, n48606);
  and g81301 (n48607, n48285, n_36125);
  and g81302 (n48608, n_35899, n48286);
  not g81303 (n_36126, n48607);
  not g81304 (n_36127, n48608);
  and g81305 (n48609, n_36126, n_36127);
  not g81306 (n_36128, n48609);
  and g81307 (po0963, n48361, n_36128);
  and g81308 (n48611, n_35913, pi0987);
  not g81309 (n_36131, po0963);
  and g81310 (n48612, n_36131, n48611);
  and g81311 (n48613, pi0771, pi0945);
  and g81312 (n48614, n_36089, n48613);
  or g81313 (po0928, n48612, n48614);
  and g81314 (n48616, pi1102, po0988);
  and g81315 (n48617, pi0772, n_36029);
  not g81316 (n_36132, n48616);
  and g81317 (n48618, n_34696, n_36132);
  not g81318 (n_36133, n48618);
  or g81319 (po0929, n48617, n_36133);
  and g81320 (n48620, n_35868, n48257);
  and g81321 (n48621, po0963, n48620);
  not g81322 (n_36134, n48621);
  and g81323 (n48622, n48280, n_36134);
  not g81324 (n_36135, n48471);
  and g81325 (n48623, pi0801, n_36135);
  not g81326 (n_36136, n48623);
  and g81327 (n48624, n48258, n_36136);
  not g81328 (n_36137, n48624);
  and g81329 (n48625, pi0773, n_36137);
  not g81330 (n_36138, n48622);
  not g81331 (n_36139, n48625);
  and g81332 (n48626, n_36138, n_36139);
  not g81333 (n_36140, n48626);
  and g81334 (po0930, n_36045, n_36140);
  and g81335 (n48628, n_13676, n_36029);
  and g81336 (n48629, pi1127, po0988);
  not g81337 (n_36141, n48628);
  and g81338 (n48630, n_34696, n_36141);
  not g81339 (n_36142, n48630);
  or g81340 (po0931, n48629, n_36142);
  and g81341 (n48632, pi0775, n_36089);
  and g81342 (n48633, pi0731, n_35913);
  and g81343 (n48634, pi0765, pi0771);
  and g81344 (n48635, n48265, n48634);
  not g81350 (n_36143, n48640);
  and g81351 (n48641, n48635, n_36143);
  not g81352 (n_36144, n48641);
  and g81353 (n48642, n_35865, n_36144);
  not g81354 (n_36145, n48642);
  and g81355 (n48643, n48633, n_36145);
  not g81356 (n_36146, n48632);
  not g81357 (n_36147, n48643);
  and g81358 (n48644, n_36146, n_36147);
  not g81359 (n_36148, n48635);
  and g81360 (n48645, n_35979, n_36148);
  and g81361 (n48646, pi0775, n48633);
  not g81362 (n_36149, n48645);
  and g81363 (n48647, n_36149, n48646);
  not g81364 (n_36150, n48644);
  not g81365 (n_36151, n48647);
  and g81366 (po0932, n_36150, n_36151);
  not g81367 (n_36152, pi0776);
  and g81368 (n48649, n_36152, n_36029);
  and g81369 (n48650, pi1128, po0988);
  not g81370 (n_36153, n48649);
  and g81371 (n48651, n_34696, n_36153);
  not g81372 (n_36154, n48651);
  or g81373 (po0933, n48650, n_36154);
  and g81374 (n48653, n_15730, n_36029);
  and g81375 (n48654, pi1122, po0988);
  not g81376 (n_36155, n48653);
  and g81377 (n48655, n_34696, n_36155);
  not g81378 (n_36156, n48655);
  or g81379 (po0934, n48654, n_36156);
  not g81386 (n_36164, pi0968);
  and g81387 (n48661, n_36164, n48660);
  not g81388 (n_36165, n48661);
  and g81389 (n48662, pi0778, n_36165);
  and g81390 (n48663, pi1100, n48661);
  or g81391 (po0935, n48662, n48663);
  or g81392 (po0936, n_34704, n46839);
  or g81393 (po0937, n_34804, n46748);
  and g81394 (n48667, pi0781, n_36165);
  and g81395 (n48668, pi1101, n48661);
  or g81396 (po0938, n48667, n48668);
  not g81397 (n_36166, n42345);
  not g81398 (n_36167, n46792);
  and g81399 (n48670, n_36166, n_36167);
  not g81400 (n_36168, n48670);
  or g81401 (po0939, n46747, n_36168);
  and g81402 (n48672, pi0783, n_36165);
  and g81403 (n48673, pi1109, n48661);
  or g81404 (po0940, n48672, n48673);
  and g81405 (n48675, pi0784, n_36165);
  and g81406 (n48676, pi1110, n48661);
  or g81407 (po0941, n48675, n48676);
  and g81408 (n48678, pi0785, n_36165);
  and g81409 (n48679, pi1102, n48661);
  or g81410 (po0942, n48678, n48679);
  and g81411 (n48681, pi0024, po1110);
  and g81412 (n48682, pi0786, pi0954);
  not g81413 (n_36169, n48681);
  not g81414 (n_36170, n48682);
  and g81415 (po0943, n_36169, n_36170);
  and g81416 (n48684, pi0787, n_36165);
  and g81417 (n48685, pi1104, n48661);
  or g81418 (po0944, n48684, n48685);
  and g81419 (n48687, pi0788, n_36165);
  and g81420 (n48688, pi1105, n48661);
  or g81421 (po0945, n48687, n48688);
  and g81422 (n48690, pi0789, n_36165);
  and g81423 (n48691, pi1106, n48661);
  or g81424 (po0946, n48690, n48691);
  and g81425 (n48693, pi0790, n_36165);
  and g81426 (n48694, pi1107, n48661);
  or g81427 (po0947, n48693, n48694);
  and g81428 (n48696, pi0791, n_36165);
  and g81429 (n48697, pi1108, n48661);
  or g81430 (po0948, n48696, n48697);
  and g81431 (n48699, pi0792, n_36165);
  and g81432 (n48700, pi1103, n48661);
  or g81433 (po0949, n48699, n48700);
  and g81434 (n48702, pi0968, n48660);
  not g81435 (n_36171, n48702);
  and g81436 (n48703, pi0794, n_36171);
  and g81437 (n48704, pi1130, n48702);
  or g81438 (po0951, n48703, n48704);
  and g81439 (n48706, pi0795, n_36171);
  and g81440 (n48707, pi1128, n48702);
  or g81441 (po0952, n48706, n48707);
  and g81446 (n48713, n_34943, n48712);
  and g81447 (n48714, n47031, n48713);
  not g81448 (n_36172, n48714);
  and g81449 (n48715, pi0264, n_36172);
  and g81450 (n48716, n_34947, n48714);
  not g81451 (n_36173, n48715);
  not g81452 (n_36174, n48716);
  and g81453 (po0953, n_36173, n_36174);
  and g81454 (n48718, pi0798, n_36171);
  and g81455 (n48719, pi1124, n48702);
  or g81456 (po0955, n48718, n48719);
  and g81457 (n48721, pi0799, n_36171);
  and g81458 (n48722, n_34723, n48702);
  not g81459 (n_36175, n48721);
  not g81460 (n_36176, n48722);
  and g81461 (po0956, n_36175, n_36176);
  and g81462 (n48724, pi0800, n_36171);
  and g81463 (n48725, pi1125, n48702);
  or g81464 (po0957, n48724, n48725);
  and g81465 (n48727, pi0801, n_36171);
  and g81466 (n48728, pi1126, n48702);
  or g81467 (po0958, n48727, n48728);
  and g81468 (n48730, pi0803, n_36171);
  and g81469 (n48731, n_34800, n48702);
  not g81470 (n_36177, n48730);
  not g81471 (n_36178, n48731);
  and g81472 (po0960, n_36177, n_36178);
  and g81473 (n48733, pi0804, n_36171);
  and g81474 (n48734, pi1109, n48702);
  or g81475 (po0961, n48733, n48734);
  and g81476 (n48736, n_34946, n47029);
  and g81477 (n48737, n_34944, n48736);
  not g81478 (n_36179, n48736);
  and g81479 (n48738, pi0270, n_36179);
  not g81480 (n_36180, n48737);
  not g81481 (n_36181, n48738);
  and g81482 (po0962, n_36180, n_36181);
  and g81483 (n48740, pi0807, n_36171);
  and g81484 (n48741, pi1127, n48702);
  or g81485 (po0964, n48740, n48741);
  and g81486 (n48743, pi0808, n_36171);
  and g81487 (n48744, pi1101, n48702);
  or g81488 (po0965, n48743, n48744);
  and g81489 (n48746, pi0809, n_36171);
  and g81490 (n48747, n_34874, n48702);
  not g81491 (n_36182, n48746);
  not g81492 (n_36183, n48747);
  and g81493 (po0966, n_36182, n_36183);
  and g81494 (n48749, pi0810, n_36171);
  and g81495 (n48750, pi1108, n48702);
  or g81496 (po0967, n48749, n48750);
  and g81497 (n48752, pi0811, n_36171);
  and g81498 (n48753, pi1102, n48702);
  or g81499 (po0968, n48752, n48753);
  and g81500 (n48755, pi0812, n_36171);
  and g81501 (n48756, n_34714, n48702);
  not g81502 (n_36184, n48755);
  not g81503 (n_36185, n48756);
  and g81504 (po0969, n_36184, n_36185);
  and g81505 (n48758, pi0813, n_36171);
  and g81506 (n48759, pi1131, n48702);
  or g81507 (po0970, n48758, n48759);
  and g81508 (n48761, pi0814, n_36171);
  and g81509 (n48762, n_34769, n48702);
  not g81510 (n_36186, n48761);
  not g81511 (n_36187, n48762);
  and g81512 (po0971, n_36186, n_36187);
  and g81513 (n48764, pi0815, n_36171);
  and g81514 (n48765, pi1110, n48702);
  or g81515 (po0972, n48764, n48765);
  and g81516 (n48767, pi0816, n_36171);
  and g81517 (n48768, pi1129, n48702);
  or g81518 (po0973, n48767, n48768);
  not g81519 (n_36188, n47027);
  and g81520 (n48770, pi0269, n_36188);
  not g81521 (n_36189, n47028);
  not g81522 (n_36190, n48770);
  and g81523 (po0974, n_36189, n_36190);
  and g81524 (n48772, n7643, n14172);
  or g81525 (po0975, n14025, n48772);
  not g81526 (n_36191, n47033);
  and g81527 (n48774, pi0265, n_36191);
  not g81528 (n_36192, n48774);
  and g81529 (po0976, n_34950, n_36192);
  and g81530 (n48776, pi0277, n_36180);
  not g81531 (n_36193, n47032);
  not g81532 (n_36194, n48776);
  and g81533 (po0977, n_36193, n_36194);
  not g81534 (n_36196, pi0811);
  not g81535 (n_36197, pi0893);
  and g81536 (po0979, n_36196, n_36197);
  not g81537 (n_36198, pi0982);
  and g81538 (n48779, n_36198, n_6537);
  and g81539 (n48780, n7626, n7643);
  not g81540 (n_36199, n48779);
  not g81541 (n_36200, n48780);
  and g81542 (n48781, n_36199, n_36200);
  not g81543 (n_36201, n48781);
  and g81544 (po0981, n2932, n_36201);
  and g81545 (n48783, pi0123, n2604);
  not g81546 (n_36202, n48783);
  and g81547 (n48784, pi1131, n_36202);
  and g81548 (n48785, pi1127, n_36202);
  not g81549 (n_36203, n48784);
  not g81550 (n_36204, n48785);
  and g81551 (n48786, n_36203, n_36204);
  not g81552 (po1147, pi0825);
  and g81553 (n48787, po1147, n48783);
  not g81554 (n_36207, n48787);
  and g81555 (n48788, n48786, n_36207);
  and g81556 (n48789, pi1131, n48785);
  not g81557 (n_36208, n48788);
  not g81558 (n_36209, n48789);
  and g81559 (n48790, n_36208, n_36209);
  and g81560 (n48791, pi1124, n_34907);
  and g81561 (n48792, n_34926, pi1130);
  not g81562 (n_36210, n48791);
  not g81563 (n_36211, n48792);
  and g81564 (n48793, n_36210, n_36211);
  and g81565 (n48794, n_34868, n_34919);
  and g81566 (n48795, pi1128, pi1129);
  not g81567 (n_36212, n48794);
  not g81568 (n_36213, n48795);
  and g81569 (n48796, n_36212, n_36213);
  and g81570 (n48797, n_34886, n_34897);
  and g81571 (n48798, pi1125, pi1126);
  not g81572 (n_36214, n48797);
  not g81573 (n_36215, n48798);
  and g81574 (n48799, n_36214, n_36215);
  not g81575 (n_36216, n48799);
  and g81576 (n48800, n48796, n_36216);
  not g81577 (n_36217, n48796);
  and g81578 (n48801, n_36217, n48799);
  not g81579 (n_36218, n48800);
  not g81580 (n_36219, n48801);
  and g81581 (n48802, n_36218, n_36219);
  and g81582 (n48803, n48793, n48802);
  not g81583 (n_36220, n48793);
  not g81584 (n_36221, n48802);
  and g81585 (n48804, n_36220, n_36221);
  not g81586 (n_36222, n48803);
  not g81587 (n_36223, n48804);
  and g81588 (n48805, n_36222, n_36223);
  not g81589 (n_36224, n48790);
  not g81590 (n_36225, n48805);
  and g81591 (n48806, n_36224, n_36225);
  and g81592 (n48807, pi0825, n48783);
  not g81593 (n_36226, n48807);
  and g81594 (n48808, n48786, n_36226);
  and g81595 (n48809, n_36209, n48805);
  not g81596 (n_36227, n48808);
  and g81597 (n48810, n_36227, n48809);
  not g81598 (n_36228, n48806);
  not g81599 (n_36229, n48810);
  and g81600 (po0982, n_36228, n_36229);
  and g81601 (n48812, pi1123, n_36202);
  and g81602 (n48813, pi1122, n_36202);
  not g81603 (n_36230, n48812);
  not g81604 (n_36231, n48813);
  and g81605 (n48814, n_36230, n_36231);
  not g81606 (po1148, pi0826);
  and g81607 (n48815, po1148, n48783);
  not g81608 (n_36234, n48815);
  and g81609 (n48816, n48814, n_36234);
  and g81610 (n48817, pi1123, n48813);
  not g81611 (n_36235, n48816);
  not g81612 (n_36236, n48817);
  and g81613 (n48818, n_36235, n_36236);
  and g81614 (n48819, pi1118, n_34829);
  and g81615 (n48820, n_34731, pi1119);
  not g81616 (n_36237, n48819);
  not g81617 (n_36238, n48820);
  and g81618 (n48821, n_36237, n_36238);
  and g81619 (n48822, n_34835, n_34823);
  and g81620 (n48823, pi1120, pi1121);
  not g81621 (n_36239, n48822);
  not g81622 (n_36240, n48823);
  and g81623 (n48824, n_36239, n_36240);
  and g81624 (n48825, n_34727, n_34778);
  and g81625 (n48826, pi1116, pi1117);
  not g81626 (n_36241, n48825);
  not g81627 (n_36242, n48826);
  and g81628 (n48827, n_36241, n_36242);
  not g81629 (n_36243, n48827);
  and g81630 (n48828, n48824, n_36243);
  not g81631 (n_36244, n48824);
  and g81632 (n48829, n_36244, n48827);
  not g81633 (n_36245, n48828);
  not g81634 (n_36246, n48829);
  and g81635 (n48830, n_36245, n_36246);
  and g81636 (n48831, n48821, n48830);
  not g81637 (n_36247, n48821);
  not g81638 (n_36248, n48830);
  and g81639 (n48832, n_36247, n_36248);
  not g81640 (n_36249, n48831);
  not g81641 (n_36250, n48832);
  and g81642 (n48833, n_36249, n_36250);
  not g81643 (n_36251, n48818);
  not g81644 (n_36252, n48833);
  and g81645 (n48834, n_36251, n_36252);
  and g81646 (n48835, pi0826, n48783);
  not g81647 (n_36253, n48835);
  and g81648 (n48836, n48814, n_36253);
  and g81649 (n48837, n_36236, n48833);
  not g81650 (n_36254, n48836);
  and g81651 (n48838, n_36254, n48837);
  not g81652 (n_36255, n48834);
  not g81653 (n_36256, n48838);
  and g81654 (po0983, n_36255, n_36256);
  and g81655 (n48840, pi1100, n_36202);
  and g81656 (n48841, pi1107, n_36202);
  not g81657 (n_36257, n48840);
  not g81658 (n_36258, n48841);
  and g81659 (n48842, n_36257, n_36258);
  not g81660 (po1178, pi0827);
  and g81661 (n48843, po1178, n48783);
  not g81662 (n_36261, n48843);
  and g81663 (n48844, n48842, n_36261);
  and g81664 (n48845, pi1100, n48841);
  not g81665 (n_36262, n48844);
  not g81666 (n_36263, n48845);
  and g81667 (n48846, n_36262, n_36263);
  and g81668 (n48847, pi1103, n_34769);
  and g81669 (n48848, n_34874, pi1105);
  not g81670 (n_36264, n48847);
  not g81671 (n_36265, n48848);
  and g81672 (n48849, n_36264, n_36265);
  and g81673 (n48850, n_34765, n_34757);
  and g81674 (n48851, pi1101, pi1102);
  not g81675 (n_36266, n48850);
  not g81676 (n_36267, n48851);
  and g81677 (n48852, n_36266, n_36267);
  and g81678 (n48853, n_34714, n_34800);
  and g81679 (n48854, pi1104, pi1106);
  not g81680 (n_36268, n48853);
  not g81681 (n_36269, n48854);
  and g81682 (n48855, n_36268, n_36269);
  not g81683 (n_36270, n48855);
  and g81684 (n48856, n48852, n_36270);
  not g81685 (n_36271, n48852);
  and g81686 (n48857, n_36271, n48855);
  not g81687 (n_36272, n48856);
  not g81688 (n_36273, n48857);
  and g81689 (n48858, n_36272, n_36273);
  and g81690 (n48859, n48849, n48858);
  not g81691 (n_36274, n48849);
  not g81692 (n_36275, n48858);
  and g81693 (n48860, n_36274, n_36275);
  not g81694 (n_36276, n48859);
  not g81695 (n_36277, n48860);
  and g81696 (n48861, n_36276, n_36277);
  not g81697 (n_36278, n48846);
  not g81698 (n_36279, n48861);
  and g81699 (n48862, n_36278, n_36279);
  and g81700 (n48863, pi0827, n48783);
  not g81701 (n_36280, n48863);
  and g81702 (n48864, n48842, n_36280);
  and g81703 (n48865, n_36263, n48861);
  not g81704 (n_36281, n48864);
  and g81705 (n48866, n_36281, n48865);
  not g81706 (n_36282, n48862);
  not g81707 (n_36283, n48866);
  and g81708 (po0984, n_36282, n_36283);
  and g81709 (n48868, pi1115, n_36202);
  and g81710 (n48869, pi1114, n_36202);
  not g81711 (n_36284, n48868);
  not g81712 (n_36285, n48869);
  and g81713 (n48870, n_36284, n_36285);
  not g81714 (po1182, pi0828);
  and g81715 (n48871, po1182, n48783);
  not g81716 (n_36288, n48871);
  and g81717 (n48872, n48870, n_36288);
  and g81718 (n48873, pi1115, n48869);
  not g81719 (n_36289, n48872);
  not g81720 (n_36290, n48873);
  and g81721 (n48874, n_36289, n_36290);
  and g81722 (n48875, pi1110, n_34747);
  and g81723 (n48876, n_34845, pi1111);
  not g81724 (n_36291, n48875);
  not g81725 (n_36292, n48876);
  and g81726 (n48877, n_36291, n_36292);
  and g81727 (n48878, n_34788, n_34737);
  and g81728 (n48879, pi1112, pi1113);
  not g81729 (n_36293, n48878);
  not g81730 (n_36294, n48879);
  and g81731 (n48880, n_36293, n_36294);
  and g81732 (n48881, n_34792, n_34796);
  and g81733 (n48882, pi1108, pi1109);
  not g81734 (n_36295, n48881);
  not g81735 (n_36296, n48882);
  and g81736 (n48883, n_36295, n_36296);
  not g81737 (n_36297, n48883);
  and g81738 (n48884, n48880, n_36297);
  not g81739 (n_36298, n48880);
  and g81740 (n48885, n_36298, n48883);
  not g81741 (n_36299, n48884);
  not g81742 (n_36300, n48885);
  and g81743 (n48886, n_36299, n_36300);
  and g81744 (n48887, n48877, n48886);
  not g81745 (n_36301, n48877);
  not g81746 (n_36302, n48886);
  and g81747 (n48888, n_36301, n_36302);
  not g81748 (n_36303, n48887);
  not g81749 (n_36304, n48888);
  and g81750 (n48889, n_36303, n_36304);
  not g81751 (n_36305, n48874);
  not g81752 (n_36306, n48889);
  and g81753 (n48890, n_36305, n_36306);
  and g81754 (n48891, pi0828, n48783);
  not g81755 (n_36307, n48891);
  and g81756 (n48892, n48870, n_36307);
  and g81757 (n48893, n_36290, n48889);
  not g81758 (n_36308, n48892);
  and g81759 (n48894, n_36308, n48893);
  not g81760 (n_36309, n48890);
  not g81761 (n_36310, n48894);
  and g81762 (po0985, n_36309, n_36310);
  and g81763 (n48896, n2930, n7643);
  not g81764 (n_36311, n48896);
  and g81765 (n48897, pi0951, n_36311);
  not g81766 (n_36312, n48897);
  and g81767 (po0986, pi1092, n_36312);
  not g81768 (n_36313, n48712);
  and g81769 (n48899, pi0281, n_36313);
  not g81770 (n_36314, n48713);
  not g81771 (n_36315, n48899);
  and g81772 (po0987, n_36314, n_36315);
  and g81776 (n48904, pi0833, n_12418);
  or g81777 (po0990, n16887, n48904);
  and g81778 (po0991, pi0946, n2926);
  not g81779 (n_36317, n47029);
  and g81780 (n48907, pi0282, n_36317);
  not g81781 (n_36318, n48907);
  and g81782 (po0992, n_36179, n_36318);
  not g81783 (n_36320, pi0955);
  and g81784 (n48909, n_36320, pi1049);
  and g81785 (n48910, pi0837, pi0955);
  or g81786 (po0993, n48909, n48910);
  and g81787 (n48912, n_36320, pi1047);
  and g81788 (n48913, pi0838, pi0955);
  or g81789 (po0994, n48912, n48913);
  and g81790 (n48915, n_36320, pi1074);
  and g81791 (n48916, pi0839, pi0955);
  or g81792 (po0995, n48915, n48916);
  and g81793 (n48918, pi0840, n_12418);
  and g81794 (n48919, pi1196, n2926);
  or g81795 (po0996, n48918, n48919);
  and g81796 (po0997, n_5681, n8979);
  and g81797 (n48922, n_36320, pi1035);
  and g81798 (n48923, pi0842, pi0955);
  or g81799 (po0998, n48922, n48923);
  and g81800 (n48925, n_36320, pi1079);
  and g81801 (n48926, pi0843, pi0955);
  or g81802 (po0999, n48925, n48926);
  and g81803 (n48928, n_36320, pi1078);
  and g81804 (n48929, pi0844, pi0955);
  or g81805 (po1000, n48928, n48929);
  and g81806 (n48931, n_36320, pi1043);
  and g81807 (n48932, pi0845, pi0955);
  or g81808 (po1001, n48931, n48932);
  and g81809 (n48934, pi0846, n_31974);
  and g81810 (n48935, pi1134, n42902);
  or g81811 (po1002, n48934, n48935);
  and g81812 (n48937, n_36320, pi1055);
  and g81813 (n48938, pi0847, pi0955);
  or g81814 (po1003, n48937, n48938);
  and g81815 (n48940, n_36320, pi1039);
  and g81816 (n48941, pi0848, pi0955);
  or g81817 (po1004, n48940, n48941);
  and g81818 (n48943, pi0849, n_12418);
  and g81819 (n48944, pi1198, n2926);
  or g81820 (po1005, n48943, n48944);
  and g81821 (n48946, n_36320, pi1048);
  and g81822 (n48947, pi0850, pi0955);
  or g81823 (po1006, n48946, n48947);
  and g81824 (n48949, n_36320, pi1045);
  and g81825 (n48950, pi0851, pi0955);
  or g81826 (po1007, n48949, n48950);
  and g81827 (n48952, n_36320, pi1062);
  and g81828 (n48953, pi0852, pi0955);
  or g81829 (po1008, n48952, n48953);
  and g81830 (n48955, n_36320, pi1080);
  and g81831 (n48956, pi0853, pi0955);
  or g81832 (po1009, n48955, n48956);
  and g81833 (n48958, n_36320, pi1051);
  and g81834 (n48959, pi0854, pi0955);
  or g81835 (po1010, n48958, n48959);
  and g81836 (n48961, n_36320, pi1065);
  and g81837 (n48962, pi0855, pi0955);
  or g81838 (po1011, n48961, n48962);
  and g81839 (n48964, n_36320, pi1067);
  and g81840 (n48965, pi0856, pi0955);
  or g81841 (po1012, n48964, n48965);
  and g81842 (n48967, n_36320, pi1058);
  and g81843 (n48968, pi0857, pi0955);
  or g81844 (po1013, n48967, n48968);
  and g81845 (n48970, n_36320, pi1087);
  and g81846 (n48971, pi0858, pi0955);
  or g81847 (po1014, n48970, n48971);
  and g81848 (n48973, n_36320, pi1070);
  and g81849 (n48974, pi0859, pi0955);
  or g81850 (po1015, n48973, n48974);
  and g81851 (n48976, n_36320, pi1076);
  and g81852 (n48977, pi0860, pi0955);
  or g81853 (po1016, n48976, n48977);
  and g81854 (n48979, pi1093, pi1141);
  and g81855 (n48980, pi0861, n_3206);
  not g81856 (n_36323, n48979);
  not g81857 (n_36324, n48980);
  and g81858 (n48981, n_36323, n_36324);
  not g81859 (n_36325, n48981);
  and g81860 (n48982, n_188, n_36325);
  and g81861 (n48983, n_31967, n_1496);
  and g81862 (n48984, pi0123, n_1506);
  not g81863 (n_36326, n48983);
  and g81864 (n48985, pi0228, n_36326);
  not g81865 (n_36327, n48984);
  and g81866 (n48986, n_36327, n48985);
  or g81867 (po1017, n48982, n48986);
  and g81868 (n48988, pi0862, n_31974);
  and g81869 (n48989, pi1139, n42902);
  or g81870 (po1018, n48988, n48989);
  and g81871 (n48991, pi0863, n_12418);
  and g81872 (n48992, pi1199, n2926);
  or g81873 (po1019, n48991, n48992);
  and g81874 (n48994, pi0864, n_12418);
  and g81875 (n48995, pi1197, n2926);
  or g81876 (po1020, n48994, n48995);
  and g81877 (n48997, n_36320, pi1040);
  and g81878 (n48998, pi0865, pi0955);
  or g81879 (po1021, n48997, n48998);
  and g81880 (n49000, n_36320, pi1053);
  and g81881 (n49001, pi0866, pi0955);
  or g81882 (po1022, n49000, n49001);
  and g81883 (n49003, n_36320, pi1057);
  and g81884 (n49004, pi0867, pi0955);
  or g81885 (po1023, n49003, n49004);
  and g81886 (n49006, n_36320, pi1063);
  and g81887 (n49007, pi0868, pi0955);
  or g81888 (po1024, n49006, n49007);
  and g81889 (n49009, pi1093, pi1140);
  and g81890 (n49010, pi0869, n_3206);
  not g81891 (n_36330, n49009);
  not g81892 (n_36331, n49010);
  and g81893 (n49011, n_36330, n_36331);
  not g81894 (n_36332, n49011);
  and g81895 (n49012, n_188, n_36332);
  and g81896 (n49013, n_31967, n_1676);
  and g81897 (n49014, pi0123, n_1686);
  not g81898 (n_36333, n49013);
  and g81899 (n49015, pi0228, n_36333);
  not g81900 (n_36334, n49014);
  and g81901 (n49016, n_36334, n49015);
  or g81902 (po1025, n49012, n49016);
  and g81903 (n49018, n_36320, pi1069);
  and g81904 (n49019, pi0870, pi0955);
  or g81905 (po1026, n49018, n49019);
  and g81906 (n49021, n_36320, pi1072);
  and g81907 (n49022, pi0871, pi0955);
  or g81908 (po1027, n49021, n49022);
  and g81909 (n49024, n_36320, pi1084);
  and g81910 (n49025, pi0872, pi0955);
  or g81911 (po1028, n49024, n49025);
  and g81912 (n49027, n_36320, pi1044);
  and g81913 (n49028, pi0873, pi0955);
  or g81914 (po1029, n49027, n49028);
  and g81915 (n49030, n_36320, pi1036);
  and g81916 (n49031, pi0874, pi0955);
  or g81917 (po1030, n49030, n49031);
  and g81918 (n49033, pi1093, n_2388);
  and g81919 (n49034, n_2398, n_3206);
  not g81920 (n_36335, n49033);
  not g81921 (n_36336, n49034);
  and g81922 (n49035, n_36335, n_36336);
  not g81923 (n_36337, n49035);
  and g81924 (n49036, n_188, n_36337);
  and g81925 (n49037, n_31967, pi1136);
  and g81926 (n49038, pi0123, pi0875);
  not g81927 (n_36338, n49037);
  and g81928 (n49039, pi0228, n_36338);
  not g81929 (n_36339, n49038);
  and g81930 (n49040, n_36339, n49039);
  not g81931 (n_36340, n49036);
  not g81932 (n_36341, n49040);
  and g81933 (po1031, n_36340, n_36341);
  and g81934 (n49042, n_36320, pi1037);
  and g81935 (n49043, pi0876, pi0955);
  or g81936 (po1032, n49042, n49043);
  and g81937 (n49045, pi1093, pi1138);
  and g81938 (n49046, pi0877, n_3206);
  not g81939 (n_36342, n49045);
  not g81940 (n_36343, n49046);
  and g81941 (n49047, n_36342, n_36343);
  not g81942 (n_36344, n49047);
  and g81943 (n49048, n_188, n_36344);
  and g81944 (n49049, n_31967, n_2030);
  and g81945 (n49050, pi0123, n_2040);
  not g81946 (n_36345, n49049);
  and g81947 (n49051, pi0228, n_36345);
  not g81948 (n_36346, n49050);
  and g81949 (n49052, n_36346, n49051);
  or g81950 (po1033, n49048, n49052);
  and g81951 (n49054, pi1093, pi1137);
  and g81952 (n49055, pi0878, n_3206);
  not g81953 (n_36347, n49054);
  not g81954 (n_36348, n49055);
  and g81955 (n49056, n_36347, n_36348);
  not g81956 (n_36349, n49056);
  and g81957 (n49057, n_188, n_36349);
  and g81958 (n49058, n_31967, n_2209);
  and g81959 (n49059, pi0123, n_2219);
  not g81960 (n_36350, n49058);
  and g81961 (n49060, pi0228, n_36350);
  not g81962 (n_36351, n49059);
  and g81963 (n49061, n_36351, n49060);
  or g81964 (po1034, n49057, n49061);
  and g81965 (n49063, pi1093, pi1135);
  and g81966 (n49064, pi0879, n_3206);
  not g81967 (n_36352, n49063);
  not g81968 (n_36353, n49064);
  and g81969 (n49065, n_36352, n_36353);
  not g81970 (n_36354, n49065);
  and g81971 (n49066, n_188, n_36354);
  and g81972 (n49067, n_31967, n_2581);
  and g81973 (n49068, pi0123, n_2591);
  not g81974 (n_36355, n49067);
  and g81975 (n49069, pi0228, n_36355);
  not g81976 (n_36356, n49068);
  and g81977 (n49070, n_36356, n49069);
  or g81978 (po1035, n49066, n49070);
  and g81979 (n49072, n_36320, pi1081);
  and g81980 (n49073, pi0880, pi0955);
  or g81981 (po1036, n49072, n49073);
  and g81982 (n49075, n_36320, pi1059);
  and g81983 (n49076, pi0881, pi0955);
  or g81984 (po1037, n49075, n49076);
  not g81985 (po1163, pi0883);
  and g81986 (n49078, po1163, n48783);
  or g81987 (po1039, n48841, n49078);
  and g81988 (n49080, pi1124, n_36202);
  not g81989 (po1180, pi0884);
  and g81990 (n49081, po1180, n48783);
  or g81991 (po1040, n49080, n49081);
  and g81992 (n49083, pi1125, n_36202);
  not g81993 (po1172, pi0885);
  and g81994 (n49084, po1172, n48783);
  or g81995 (po1041, n49083, n49084);
  and g81996 (n49086, pi1109, n_36202);
  not g81997 (po1166, pi0886);
  and g81998 (n49087, po1166, n48783);
  or g81999 (po1042, n49086, n49087);
  not g82000 (po1179, pi0887);
  and g82001 (n49089, po1179, n48783);
  or g82002 (po1043, n48840, n49089);
  and g82003 (n49091, pi1120, n_36202);
  not g82004 (po1164, pi0888);
  and g82005 (n49092, po1164, n48783);
  or g82006 (po1044, n49091, n49092);
  and g82007 (n49094, pi1103, n_36202);
  not g82008 (po1170, pi0889);
  and g82009 (n49095, po1170, n48783);
  or g82010 (po1045, n49094, n49095);
  and g82011 (n49097, pi1126, n_36202);
  not g82012 (po1153, pi0890);
  and g82013 (n49098, po1153, n48783);
  or g82014 (po1046, n49097, n49098);
  and g82015 (n49100, pi1116, n_36202);
  not g82016 (po1160, pi0891);
  and g82017 (n49101, po1160, n48783);
  or g82018 (po1047, n49100, n49101);
  and g82019 (n49103, pi1101, n_36202);
  not g82020 (po1183, pi0892);
  and g82021 (n49104, po1183, n48783);
  or g82022 (po1048, n49103, n49104);
  and g82023 (n49106, pi1119, n_36202);
  not g82024 (po1150, pi0894);
  and g82025 (n49107, po1150, n48783);
  or g82026 (po1050, n49106, n49107);
  and g82027 (n49109, pi1113, n_36202);
  not g82028 (po1168, pi0895);
  and g82029 (n49110, po1168, n48783);
  or g82030 (po1051, n49109, n49110);
  and g82031 (n49112, pi1118, n_36202);
  not g82032 (po1156, pi0896);
  and g82033 (n49113, po1156, n48783);
  or g82034 (po1052, n49112, n49113);
  and g82035 (n49115, pi1129, n_36202);
  not g82036 (po1176, pi0898);
  and g82037 (n49116, po1176, n48783);
  or g82038 (po1054, n49115, n49116);
  not g82039 (po1174, pi0899);
  and g82040 (n49118, po1174, n48783);
  or g82041 (po1055, n48868, n49118);
  and g82042 (n49120, pi1110, n_36202);
  not g82043 (po1171, pi0900);
  and g82044 (n49121, po1171, n48783);
  or g82045 (po1056, n49120, n49121);
  and g82046 (n49123, pi1111, n_36202);
  not g82047 (po1161, pi0902);
  and g82048 (n49124, po1161, n48783);
  or g82049 (po1058, n49123, n49124);
  and g82050 (n49126, pi1121, n_36202);
  not g82051 (po1162, pi0903);
  and g82052 (n49127, po1162, n48783);
  or g82053 (po1059, n49126, n49127);
  not g82054 (po1173, pi0904);
  and g82055 (n49129, po1173, n48783);
  or g82056 (po1060, n48785, n49129);
  not g82057 (po1151, pi0905);
  and g82058 (n49131, po1151, n48783);
  or g82059 (po1061, n48784, n49131);
  and g82060 (n49133, pi1128, n_36202);
  not g82061 (po1155, pi0906);
  and g82062 (n49134, po1155, n48783);
  or g82063 (po1062, n49133, n49134);
  not g82064 (n_36400, pi0782);
  and g82065 (n49136, n_36400, n_3148);
  not g82066 (n_36401, pi0624);
  and g82067 (n49137, n_36401, n_3080);
  not g82068 (n_36402, pi0598);
  and g82069 (n49138, n_36402, pi0979);
  not g82070 (n_36403, n49137);
  and g82071 (n49139, pi0782, n_36403);
  not g82072 (n_36404, n49138);
  and g82073 (n49140, n_36404, n49139);
  not g82074 (n_36405, pi0604);
  and g82075 (n49141, n_36405, n_3080);
  and g82076 (n49142, pi0615, pi0979);
  not g82077 (n_36406, n49141);
  not g82078 (n_36407, n49142);
  and g82079 (n49143, n_36406, n_36407);
  not g82080 (n_36408, n49143);
  and g82081 (n49144, pi0782, n_36408);
  not g82082 (n_36409, n49136);
  not g82083 (n_36410, n49140);
  and g82084 (n49145, n_36409, n_36410);
  not g82085 (n_36411, n49144);
  and g82086 (po1063, n_36411, n49145);
  not g82087 (po1159, pi0908);
  and g82088 (n49147, po1159, n48783);
  or g82089 (po1064, n48813, n49147);
  and g82090 (n49149, pi1105, n_36202);
  not g82091 (po1157, pi0909);
  and g82092 (n49150, po1157, n48783);
  or g82093 (po1065, n49149, n49150);
  and g82094 (n49152, pi1117, n_36202);
  not g82095 (po1181, pi0910);
  and g82096 (n49153, po1181, n48783);
  or g82097 (po1066, n49152, n49153);
  and g82098 (n49155, pi1130, n_36202);
  not g82099 (po1158, pi0911);
  and g82100 (n49156, po1158, n48783);
  or g82101 (po1067, n49155, n49156);
  not g82102 (po1167, pi0912);
  and g82103 (n49158, po1167, n48783);
  or g82104 (po1068, n48869, n49158);
  and g82105 (n49160, pi1106, n_36202);
  not g82106 (po1149, pi0913);
  and g82107 (n49161, po1149, n48783);
  or g82108 (po1069, n49160, n49161);
  not g82109 (n_36424, n47026);
  and g82110 (n49163, pi0280, n_36424);
  not g82111 (n_36425, n49163);
  and g82112 (po1070, n_36188, n_36425);
  and g82113 (n49165, pi1108, n_36202);
  not g82114 (po1146, pi0915);
  and g82115 (n49166, po1146, n48783);
  or g82116 (po1071, n49165, n49166);
  not g82117 (po1169, pi0916);
  and g82118 (n49168, po1169, n48783);
  or g82119 (po1072, n48812, n49168);
  and g82120 (n49170, pi1112, n_36202);
  not g82121 (po1177, pi0917);
  and g82122 (n49171, po1177, n48783);
  or g82123 (po1073, n49170, n49171);
  and g82124 (n49173, pi1104, n_36202);
  not g82125 (po1175, pi0918);
  and g82126 (n49174, po1175, n48783);
  or g82127 (po1074, n49173, n49174);
  and g82128 (n49176, pi1102, n_36202);
  not g82129 (po1165, pi0919);
  and g82130 (n49177, po1165, n48783);
  or g82131 (po1075, n49176, n49177);
  and g82132 (n49179, pi1093, pi1139);
  and g82133 (n49180, pi0920, n_3206);
  or g82134 (po1076, n49179, n49180);
  and g82135 (n49182, pi0921, n_3206);
  or g82136 (po1077, n49009, n49182);
  and g82137 (n49184, n_33603, n_3206);
  and g82138 (n49185, pi1093, n_28873);
  not g82139 (n_36436, n49184);
  not g82140 (n_36437, n49185);
  and g82141 (po1078, n_36436, n_36437);
  not g82142 (n_36438, pi0923);
  and g82143 (n49187, n_36438, n_3206);
  and g82144 (n49188, pi1093, n_11413);
  not g82145 (n_36439, n49187);
  not g82146 (n_36440, n49188);
  and g82147 (po1079, n_36439, n_36440);
  not g82151 (n_36441, pi0925);
  and g82152 (n49193, n_36441, n_3206);
  and g82153 (n49194, pi1093, n_11768);
  not g82154 (n_36442, n49193);
  not g82155 (n_36443, n49194);
  and g82156 (po1081, n_36442, n_36443);
  not g82157 (n_36444, pi0926);
  and g82158 (n49196, n_36444, n_3206);
  and g82159 (n49197, pi1093, n_11810);
  not g82160 (n_36445, n49196);
  not g82161 (n_36446, n49197);
  and g82162 (po1082, n_36445, n_36446);
  and g82163 (n49199, n_988, n_3206);
  and g82164 (n49200, pi1093, n_986);
  not g82165 (n_36447, n49199);
  not g82166 (n_36448, n49200);
  and g82167 (po1083, n_36447, n_36448);
  and g82168 (n49202, n_2390, n_3206);
  not g82169 (n_36449, n49202);
  and g82170 (po1084, n_36335, n_36449);
  and g82171 (n49204, n_228, n_3206);
  and g82172 (n49205, pi1093, n_5);
  not g82173 (n_36450, n49204);
  not g82174 (n_36451, n49205);
  and g82175 (po1085, n_36450, n_36451);
  and g82176 (n49207, n_2773, n_3206);
  and g82177 (n49208, pi1093, n_2921);
  not g82178 (n_36452, n49207);
  not g82179 (n_36453, n49208);
  and g82180 (po1086, n_36452, n_36453);
  and g82181 (n49210, n_33612, n_3206);
  and g82182 (n49211, pi1093, n_30133);
  not g82183 (n_36454, n49210);
  not g82184 (n_36455, n49211);
  and g82185 (po1087, n_36454, n_36455);
  and g82186 (n49213, pi0932, n_3206);
  or g82187 (po1088, n42891, n49213);
  and g82188 (n49215, pi0933, n_3206);
  or g82189 (po1089, n49054, n49215);
  and g82190 (n49217, n_33338, n_3206);
  and g82191 (n49218, pi1093, n_29810);
  not g82192 (n_36456, n49217);
  not g82193 (n_36457, n49218);
  and g82194 (po1090, n_36456, n_36457);
  and g82195 (n49220, pi0935, n_3206);
  or g82196 (po1091, n48979, n49220);
  and g82197 (n49222, n_33621, n_3206);
  and g82198 (n49223, pi1093, n_29850);
  not g82199 (n_36458, n49222);
  not g82200 (n_36459, n49223);
  and g82201 (po1092, n_36458, n_36459);
  and g82202 (n49225, n_33322, n_3206);
  and g82203 (n49226, pi1093, n_29904);
  not g82204 (n_36460, n49225);
  not g82205 (n_36461, n49226);
  and g82206 (po1093, n_36460, n_36461);
  and g82207 (n49228, pi0938, n_3206);
  or g82208 (po1094, n49063, n49228);
  and g82209 (n49230, n_805, n_3206);
  and g82210 (n49231, pi1093, n_803);
  not g82211 (n_36462, n49230);
  not g82212 (n_36463, n49231);
  and g82213 (po1095, n_36462, n_36463);
  and g82214 (n49233, pi0940, n_3206);
  or g82215 (po1096, n49045, n49233);
  not g82216 (n_36464, pi0941);
  and g82217 (n49235, n_36464, n_3206);
  and g82218 (n49236, pi1093, n_11757);
  not g82219 (n_36465, n49235);
  not g82220 (n_36466, n49236);
  and g82221 (po1097, n_36465, n_36466);
  not g82222 (n_36467, pi0942);
  and g82223 (n49238, n_36467, n_3206);
  and g82224 (n49239, pi1093, n_11794);
  not g82225 (n_36468, n49238);
  not g82226 (n_36469, n49239);
  and g82227 (po1098, n_36468, n_36469);
  and g82228 (n49241, n_33507, n_3206);
  and g82229 (n49242, pi1093, n_29468);
  not g82230 (n_36470, n49241);
  not g82231 (n_36471, n49242);
  and g82232 (po1099, n_36470, n_36471);
  and g82233 (n49244, pi1093, pi1143);
  and g82234 (n49245, pi0944, n_3206);
  or g82235 (po1100, n49244, n49245);
  and g82236 (po1102, pi0230, n2926);
  and g82237 (n49248, n_36400, pi0947);
  or g82238 (po1103, n49140, n49248);
  not g82239 (n_36472, pi0992);
  and g82240 (n49250, n_2416, n_36472);
  not g82241 (n_36473, n49250);
  and g82242 (po1104, n_36424, n_36473);
  not g82243 (n_36474, pi0313);
  and g82244 (n49252, n_36474, po1110);
  and g82245 (n49253, pi0949, pi0954);
  or g82246 (po1105, n49252, n49253);
  and g82247 (po1107, n_4214, n14271);
  and g82248 (n49256, pi0957, pi1092);
  or g82249 (po1112, pi0031, n49256);
  and g82250 (po1115, n_36400, pi0960);
  and g82251 (po1116, n_28510, pi0961);
  and g82252 (po1118, n_36400, pi0963);
  and g82253 (po1122, n_28510, pi0967);
  and g82254 (po1124, n_28510, pi0969);
  and g82255 (po1125, n_36400, pi0970);
  and g82256 (po1126, n_28510, pi0971);
  and g82257 (po1127, n_36400, pi0972);
  and g82258 (po1128, n_28510, pi0974);
  and g82259 (po1129, n_36400, pi0975);
  and g82260 (po1131, n_28510, pi0977);
  and g82261 (po1132, n_36400, pi0978);
  or g82262 (po1133, pi0598, n_34761);
  and g82263 (po1135, pi0824, pi1092);
  or g82264 (po1137, pi0604, pi0624);
  not g82265 (po0170, pi1090);
  and g82266 (n2652, n_37592, n2549, n_272, n_280);
  not g82267 (n_37592, n2649);
  and g82268 (n3092, n_37593, n_37594, pi0210, pi0234);
  not g82269 (n_37593, n3089);
  not g82270 (n_37594, n3085);
  nor g82271 (n_37596, n3053, n3055);
  and g82272 (n3059, n_37595, n_271, n_148, n_37596);
  not g82273 (n_37595, n3054);
  and g82274 (n_37597, n2916, n2705);
  and g82275 (n2920, pi0225, n_130, n_143, n_37597);
  and g82276 (n2942, n_37598, n2937, n2935, n2938);
  not g82277 (n_37598, n2939);
  and g82278 (n_37599, n3394, n3334);
  and g82279 (n3398, n3382, n_162, n3383, n_37599);
  and g82280 (n3421, n3418, n3334, n_20, n_188);
  and g82281 (n3659, n_37600, n_37601, pi0235, n3328);
  not g82282 (n_37600, n3656);
  not g82283 (n_37601, n3570);
  and g82284 (n3708, n_37602, n_37603, n_1106, n3328);
  not g82285 (n_37602, n3705);
  not g82286 (n_37603, n3665);
  and g82287 (n3938, n_37604, n_37605, pi0238, n3328);
  not g82288 (n_37604, n3935);
  not g82289 (n_37605, n3865);
  and g82290 (n3853, n_37606, n_37607, n_1226, n3328);
  not g82291 (n_37606, n3850);
  not g82292 (n_37607, n3746);
  and g82293 (n4304, n_37608, n_37609, n_1595, n3328);
  not g82294 (n_37608, n4301);
  not g82295 (n_37609, n4202);
  and g82296 (n4388, n_37610, n_37611, pi0241, n3328);
  not g82297 (n_37610, n4385);
  not g82298 (n_37611, n4316);
  and g82299 (n4527, n_37612, n_37613, n_1774, n3328);
  not g82300 (n_37612, n4524);
  not g82301 (n_37613, n4425);
  and g82302 (n4611, n_37614, n_37615, pi0248, n3328);
  not g82303 (n_37614, n4608);
  not g82304 (n_37615, n4539);
  and g82305 (n4740, n_37616, n_37617, pi0299, n_1861);
  not g82306 (n_37616, n4737);
  not g82307 (n_37617, n4728);
  and g82308 (n4981, n_37618, n_37619, n_2128, n3328);
  not g82309 (n_37618, n4978);
  not g82310 (n_37619, n4879);
  and g82311 (n5065, n_37620, n_37621, pi0246, n3328);
  not g82312 (n_37620, n5062);
  not g82313 (n_37621, n4993);
  and g82314 (n5204, n_37622, n_37623, n_2307, n3328);
  not g82315 (n_37622, n5201);
  not g82316 (n_37623, n5102);
  and g82317 (n5288, n_37624, n_37625, pi0240, n3328);
  not g82318 (n_37624, n5285);
  not g82319 (n_37625, n5216);
  nor g82320 (n_37626, pi0969, pi0971);
  nor g82321 (n_37627, pi0974, pi0977);
  nor g82322 (n_37628, pi0961, pi0967);
  and g82323 (n_37629, n_3105, n_3106);
  and g82324 (n6205, n_37626, n_37627, n_37628, n_37629);
  nor g82325 (n_37632, pi0960, pi0963);
  nor g82326 (n_37633, pi0970, pi0972);
  and g82327 (n6241, n_37630, n_37631, n_37632, n_37633);
  not g82328 (n_37630, pi0975);
  not g82329 (n_37631, pi0978);
  and g82330 (n6373, n_37634, n_37635, n_188, n_3235);
  not g82331 (n_37634, n6370);
  not g82332 (n_37635, n6369);
  and g82333 (n6527, pi0145, pi0180, pi0181, pi0182);
  and g82334 (n6628, n_37636, n_37637, n_37638, n_188);
  not g82335 (n_37636, n6624);
  not g82336 (n_37637, n6625);
  not g82337 (n_37638, n6623);
  and g82338 (n7326, n_37639, n_37640, n_37641, pi0232);
  not g82339 (n_37639, n7323);
  not g82340 (n_37640, n7320);
  not g82341 (n_37641, n7321);
  and g82342 (n7320, n_37642, n_3586, n_234, n_3399);
  not g82343 (n_37642, n7317);
  and g82344 (n7617, n_37643, n7612, n6384, n7519);
  not g82345 (n_37643, n7542);
  nor g82346 (n_37645, n8401, n8409);
  and g82347 (n8414, n_37644, pi1199, n8410, n_37645);
  not g82348 (n_37644, n8406);
  and g82349 (n8422, n_37646, n_37647, pi1196, n8410);
  not g82350 (n_37646, n8419);
  not g82351 (n_37647, n8416);
  and g82352 (n_37648, n2772, n6491);
  and g82353 (n7526, n_123, n_127, pi0097, n_37648);
  and g82354 (n_37649, n8963, n_5662);
  and g82355 (n8971, n_5661, n_186, n8967, n_37649);
  nor g82356 (n_37650, n8937, n8933);
  and g82357 (n_37651, n_5637, n8938);
  and g82358 (n8943, n_186, n7445, n_37650, n_37651);
  and g82359 (n_37652, n2479, pi0076, n_91);
  and g82360 (n_37653, n8909, n8920);
  and g82361 (n_37654, n8914, n8922);
  and g82362 (n_37655, n8912, n8919);
  and g82363 (n8930, n_37652, n_37653, n_37654, n_37655);
  and g82364 (n8919, n8916, n8915, n_72, n_85);
  and g82365 (n9215, n6135, n9212, n_164, n9208);
  and g82366 (n9345, n_37656, n_37657, pi0039, n_5920);
  not g82367 (n_37656, n9341);
  not g82368 (n_37657, n9342);
  and g82369 (n9181, n_37658, n_37659, n_37660, pi0299);
  not g82370 (n_37658, n9171);
  not g82371 (n_37659, n9178);
  not g82372 (n_37660, n9160);
  and g82373 (n9171, n_37661, n_37662, pi0149, n6197);
  not g82374 (n_37661, n9164);
  not g82375 (n_37662, n9168);
  and g82376 (n9621, n_37663, n_37664, n_6121, n9603);
  not g82377 (n_37663, n9618);
  not g82378 (n_37664, n9610);
  and g82379 (n_37665, n2477, n9083);
  and g82380 (n_37666, n9080, n9076);
  and g82381 (n9088, pi0073, n_94, n_37665, n_37666);
  and g82382 (n_37667, n6222, n9208);
  and g82383 (n9870, n9159, n_174, pi0162, n_37667);
  and g82384 (n10032, n_37668, n_37669, n_172, n_6342);
  not g82385 (n_37668, n10003);
  not g82386 (n_37669, n10029);
  and g82387 (n9923, n_37670, n_37671, n_6224, n_6121);
  not g82388 (n_37670, n9920);
  not g82389 (n_37671, n9916);
  and g82390 (n9808, n_37672, n_37673, n_37674, pi0299);
  not g82391 (n_37672, n9805);
  not g82392 (n_37673, n9802);
  not g82393 (n_37674, n9799);
  and g82394 (n10143, n_37675, n_37676, n2529, n8879);
  not g82395 (n_37675, n10140);
  not g82396 (n_37676, n10072);
  and g82397 (n10130, n_37677, n_37678, n_162, n_164);
  not g82398 (n_37677, n10126);
  not g82399 (n_37678, n10127);
  and g82400 (n10126, n_37679, n_37680, n_37681, n_161);
  not g82401 (n_37679, n10105);
  not g82402 (n_37680, n10123);
  not g82403 (n_37681, n10120);
  and g82404 (n10120, n_37682, n_37683, n2518, n10097);
  not g82405 (n_37682, n10115);
  not g82406 (n_37683, n10117);
  and g82407 (n10102, n7432, n8895, pi0032, n_131);
  and g82408 (n_37684, n10153, n10151);
  and g82409 (n10157, n10152, pi0036, n_61, n_37684);
  and g82410 (n10150, n9081, n2487, n_56, n2462);
  and g82411 (n_37686, n_37685, n10169);
  not g82412 (n_37685, n10183);
  and g82413 (n_37687, n10186, n2465);
  and g82414 (n10191, n_162, n_3052, n_37686, n_37687);
  and g82415 (n_37688, n10174, n9080);
  and g82416 (n_37689, n10171, n_79);
  and g82417 (n_37690, n_56, pi0089);
  and g82418 (n_37691, n_94, n_91);
  and g82419 (n10181, n_37688, n_37689, n_37690, n_37691);
  and g82420 (n10232, n_37692, n6382, po0740, n10201);
  not g82421 (n_37692, n10229);
  and g82422 (n10269, n_37693, n_37694, n2500, n2700);
  not g82423 (n_37693, n10266);
  not g82424 (n_37694, n10239);
  and g82425 (n10259, n10244, n10256, n_122, n10243);
  and g82426 (n_37695, n10174, n9078, n8910);
  and g82427 (n_37696, n8914, n10247, n10170);
  and g82428 (n_37697, pi0048, n_83);
  and g82429 (n_37698, n_90, n_94);
  and g82430 (n10256, n_37695, n_37696, n_37697, n_37698);
  and g82431 (n_37699, n2490, n2501);
  and g82432 (n_37700, n6170, n2464);
  and g82434 (n10286, pi0102, n_37699, n_37700, n2938);
  and g82435 (n10482, n_37702, po1038, n_134, n_6665);
  not g82436 (n_37702, n10479);
  and g82437 (n10470, n_37703, n_37704, n_37705, n_172);
  not g82438 (n_37703, n10467);
  not g82439 (n_37704, n10367);
  not g82440 (n_37705, n10354);
  and g82441 (n10353, n_37706, n_37707, n_6664, pi0087);
  not g82442 (n_37706, n10350);
  not g82443 (n_37707, n10340);
  and g82444 (n10394, n_37708, n_37709, n6479, n10391);
  not g82445 (n_37708, n10386);
  not g82446 (n_37709, n10390);
  and g82447 (n10384, n_37710, n10378, n_108, n10377);
  not g82448 (n_37710, n10381);
  and g82449 (n10695, n_37711, n_37712, n_37713, n_172);
  not g82450 (n_37711, n10692);
  not g82451 (n_37712, n10686);
  not g82452 (n_37713, n10688);
  and g82453 (n10595, n_37714, n_37715, pi0228, n_6840);
  not g82454 (n_37714, n10577);
  not g82455 (n_37715, n10592);
  and g82456 (n10866, n_37716, n_37717, n_37718, n_172);
  not g82457 (n_37716, n10863);
  not g82458 (n_37717, n10854);
  not g82459 (n_37718, n10856);
  and g82460 (n10891, n_37719, n_37720, n_37721, n_172);
  not g82461 (n_37719, n10888);
  not g82462 (n_37720, n10881);
  not g82463 (n_37721, n10882);
  and g82464 (n10801, n_37722, n_37723, n_37724, n_172);
  not g82465 (n_37722, n10798);
  not g82466 (n_37723, n10771);
  not g82467 (n_37724, n10773);
  and g82468 (n10833, n_37725, n_37726, n_37727, n_172);
  not g82469 (n_37725, n10830);
  not g82470 (n_37726, n10823);
  not g82471 (n_37727, n10824);
  and g82472 (n10968, n_37728, n_37729, n_37730, n_172);
  not g82473 (n_37728, n10965);
  not g82474 (n_37729, n10947);
  not g82475 (n_37730, n10939);
  and g82476 (n_37731, n8935, n10989, n10172);
  and g82477 (n_37732, n10987, n10247, n8912);
  and g82478 (n_37733, pi0061, n_94, n_60);
  and g82479 (n_37734, n_81, n7438, n8915);
  and g82480 (n11000, n_37731, n_37732, n_37733, n_37734);
  and g82481 (po0205, n_37735, n_37736, n_37737, n10165);
  not g82482 (n_37735, n11038);
  not g82483 (n_37736, n11042);
  not g82484 (n_37737, n11047);
  and g82485 (n11017, n_37738, n11012, n_47, n11014);
  not g82486 (n_37738, n11011);
  and g82487 (n_37739, n11006, n10171);
  and g82488 (n11010, n2805, n_91, pi0104, n_37739);
  and g82489 (n_37740, n10185, n10165);
  and g82490 (po0206, n10256, n_138, n11052, n_37740);
  and g82491 (po0207, n_37741, n_37742, n7363, n_4226);
  not g82492 (n_37741, n11072);
  not g82493 (n_37742, n11071);
  and g82494 (n_37743, n11006, n11061);
  and g82495 (n_37744, n11057, n10987);
  and g82496 (n11066, n_87, pi0049, n_37743, n_37744);
  and g82497 (n11085, n_37745, n_37746, n10162, n11080);
  not g82498 (n_37745, n11077);
  not g82499 (n_37746, n11082);
  and g82500 (n_37748, n_37747, n8901);
  not g82501 (n_37747, n11080);
  and g82502 (n11090, n11086, pi0024, n_43, n_37748);
  and g82503 (n11255, n_37749, n_37750, n_37751, n_4226);
  not g82504 (n_37749, n11252);
  not g82505 (n_37750, n11201);
  not g82506 (n_37751, n11203);
  and g82507 (n11250, n_37752, n_37753, n7429, n_6900);
  not g82508 (n_37752, n11240);
  not g82509 (n_37753, n11247);
  and g82510 (n11197, n_37754, n_37755, n_37756, pi0075);
  not g82511 (n_37754, n11192);
  not g82512 (n_37755, n11193);
  not g82513 (n_37756, n11194);
  and g82514 (n11238, n_37757, n_37758, n_37759, n_172);
  not g82515 (n_37757, n11233);
  not g82516 (n_37758, n11235);
  not g82517 (n_37759, n11179);
  and g82518 (po0211, n_37760, n_880, n10200, n_7337);
  not g82519 (n_37760, n11269);
  and g82520 (n11267, n2721, n2717, pi0053, n2720);
  and g82521 (n11287, n11282, n11284, n2611, n2706);
  and g82522 (n_37761, n11057, n10989, pi0106);
  and g82523 (n_37762, n_117, n_76);
  and g82524 (n_37763, n2479, n8913);
  and g82525 (n_37764, n8919, n11059);
  and g82526 (n11281, n_37761, n_37762, n_37763, n_37764);
  and g82527 (n_37765, n2476, n11061);
  and g82528 (n11299, n2487, pi0045, n2479, n_37765);
  and g82529 (n_37766, n6380, n6182);
  and g82530 (n11337, n_3082, pi0039, n_3080, n_37766);
  and g82531 (n11340, n2718, n11273, n_162, n11264);
  and g82532 (po0223, n_37767, n_37768, n10200, n11369);
  not g82533 (n_37767, n10223);
  not g82534 (n_37768, n10217);
  and g82535 (n11382, n11379, n11374, n2609, n11373);
  and g82536 (n11379, n2489, n11376, pi0081, n_53);
  and g82537 (n_37769, n2484, n11376);
  and g82538 (n_37770, n10165, n11102);
  and g82539 (po0225, pi0083, n_61, n_37769, n_37770);
  and g82540 (n_37772, n_37771, n6438);
  not g82541 (n_37771, n11405);
  and g82542 (n11409, n2465, n_105, n_3310, n_37772);
  and g82543 (n_37773, n2485, n10150);
  and g82544 (n11413, n7438, pi0071, pi0314, n_37773);
  and g82545 (n11430, n_37774, n_7402, n_3281, n6381);
  not g82546 (n_37774, pi0593);
  and g82547 (n_37776, n_37775, n11443);
  not g82548 (n_37775, n11441);
  and g82549 (n11452, n10162, pi0314, n_7411, n_37776);
  and g82550 (n11455, n11438, n11376, n11012, n11448);
  and g82551 (n11463, n2870, n11460, n6388, n9141);
  nor g82552 (n_37777, n11489, n11491);
  and g82553 (n_37778, n7456, n_7437);
  and g82554 (n_37779, n3373, n7429);
  and g82555 (n11497, n_5636, n_37777, n_37778, n_37779);
  and g82556 (n11875, n11746, n11872, n_174, n2609);
  and g82557 (n11733, n2509, n11730, n2518, n2609);
  and g82558 (n11987, n_37780, n_37781, n_37782, pi0039);
  not g82559 (n_37780, n11984);
  not g82560 (n_37781, n11975);
  not g82561 (n_37782, n11940);
  nor g82562 (n_37783, n12136, n12140);
  and g82563 (n12144, n11765, n_7715, n_7617, n_37783);
  and g82564 (n11760, n_37784, n11746, n_3119, n9051);
  not g82565 (n_37784, n11757);
  nor g82566 (n_37785, n11825, n11828);
  and g82567 (n11832, n_7688, pi0182, pi0184, n_37785);
  and g82568 (n11787, n_37786, n_37787, n_143, n_7591);
  not g82569 (n_37786, n11783);
  not g82570 (n_37787, n11784);
  nor g82571 (n_37788, n12073, n12070);
  and g82572 (n12077, n_7835, n_7697, n6197, n_37788);
  and g82573 (n11818, n_37789, n_37790, n_143, pi0163);
  not g82574 (n_37789, n11812);
  not g82575 (n_37790, n11815);
  and g82576 (n11845, n_37791, n_37792, n_7715, pi0184);
  not g82577 (n_37791, n11842);
  not g82578 (n_37792, n11841);
  and g82579 (n12028, n_37793, n_37794, pi0182, n_7617);
  not g82580 (n_37793, n12025);
  not g82581 (n_37794, n12024);
  and g82582 (n12011, n_37795, n_37796, n_7844, n6197);
  not g82583 (n_37795, n12006);
  not g82584 (n_37796, n12008);
  and g82585 (n11959, n_37797, n_37798, n_7636, n_3119);
  not g82586 (n_37797, n11956);
  not g82587 (n_37798, n11951);
  and g82588 (n13024, n_37799, n_37800, n_7977, n_4226);
  not g82589 (n_37799, n13021);
  not g82590 (n_37800, n12744);
  and g82591 (n12366, n_37801, n_37802, n_7977, po1038);
  not g82592 (n_37801, n12363);
  not g82593 (n_37802, n12184);
  nor g82594 (n_37803, n12381, n2704);
  and g82595 (n12385, n12378, n2962, n_3052, n_37803);
  and g82596 (n_37804, n2800, n11439);
  and g82597 (n_37805, n11014, n2480);
  and g82598 (n13036, pi0068, n_105, n_37804, n_37805);
  and g82599 (n13043, n2482, n2468, pi0066, n_69);
  and g82600 (n13096, n_37806, n_37807, n2572, n_6537);
  not g82601 (n_37806, n13088);
  not g82602 (n_37807, n13093);
  and g82603 (n_37808, n2870, n11460);
  and g82604 (n_37809, n13080, n2572);
  and g82605 (n13085, n_3206, n2519, n_37808, n_37809);
  and g82606 (po0247, n_37810, n_37811, n2520, n10165);
  not g82607 (n_37810, n13106);
  not g82608 (n_37811, n13105);
  and g82609 (n13102, n10181, n8935, n2465, n8921);
  and g82610 (po0248, n_37812, n_4093, n_466, n11326);
  not g82611 (n_37812, n13111);
  and g82612 (n_37813, n2756, n11086);
  and g82613 (n13122, n_494, pi0024, n2938, n_37813);
  and g82614 (n_37815, n_37814, n2916);
  not g82615 (n_37814, n13181);
  and g82616 (n13186, n2961, pi0096, n2510, n_37815);
  and g82617 (n13193, n_3284, n_7402, pi0039, pi0593);
  and g82618 (n13198, n_37816, n11486, n_135, n10193);
  not g82619 (n_37816, n13195);
  and g82620 (po0256, n_37817, n10164, pi0314, pi1050);
  not g82621 (n_37817, n13202);
  and g82622 (n13270, n_37818, n_37819, n_37820, n_172);
  not g82623 (n_37818, n13258);
  not g82624 (n_37819, n13267);
  not g82625 (n_37820, n13241);
  and g82626 (n13211, n10296, n_234, n_134, pi0174);
  and g82627 (n13293, n_37821, n6285, n_171, n2609);
  not g82628 (n_37821, n13290);
  and g82629 (n13296, n_5662, po0840, n_4119, n8967);
  and g82630 (n13368, n_37822, n_37823, n_37824, n_172);
  not g82631 (n_37822, n13356);
  not g82632 (n_37823, n13365);
  not g82633 (n_37824, n13335);
  and g82634 (n13402, n_37825, n_37826, n_4117, n_6537);
  not g82635 (n_37825, n13399);
  not g82636 (n_37826, n13394);
  and g82637 (n13398, n_37827, n10378, n_108, n11043);
  not g82638 (n_37827, n13395);
  and g82639 (n13429, n_37828, n_37829, n7446, n_6630);
  not g82640 (n_37828, n13425);
  not g82641 (n_37829, n13426);
  and g82642 (n_37830, n2801, n11105);
  and g82643 (n_37831, n2499, n12374);
  and g82644 (n_37832, pi0111, n_94);
  and g82645 (n13446, n_112, n_37830, n_37831, n_37832);
  and g82646 (n13548, n_37833, n_37834, n_37835, n_172);
  not g82647 (n_37833, n13545);
  not g82648 (n_37834, n13537);
  not g82649 (n_37835, n13531);
  and g82650 (n13590, n_37836, n_37837, n_37838, n_172);
  not g82651 (n_37836, n13587);
  not g82652 (n_37837, n13582);
  not g82653 (n_37838, n13576);
  and g82654 (n13633, n_37839, n_37840, n_172, n_9054);
  not g82655 (n_37839, n13622);
  not g82656 (n_37840, n13630);
  and g82657 (n13847, n_37841, n_37842, n_9119, n_824);
  not g82658 (n_37841, n13844);
  not g82659 (n_37842, n13843);
  and g82660 (n_37844, n_37843, n2521);
  not g82661 (n_37843, n13948);
  and g82662 (n_37845, n_9327, n8965);
  and g82663 (n13953, n_174, n8989, n_37844, n_37845);
  and g82664 (n13820, n_37846, n_37847, pi0190, n13815);
  not g82665 (n_37846, n13817);
  not g82666 (n_37847, n13814);
  and g82667 (n13995, n_37848, n2936, n_127, n2928);
  not g82668 (n_37848, n13992);
  and g82669 (n_37849, n2703, n7478, n10324);
  and g82670 (n_37850, n2962, n2506);
  and g82671 (n_37851, n_131, n_4081);
  and g82672 (n_37852, n2925, n8894);
  and g82673 (n14192, n_37849, n_37850, n_37851, n_37852);
  and g82674 (n14138, n_37853, n_37854, n7602, n7551);
  not g82675 (n_37853, n14134);
  not g82676 (n_37854, n14135);
  and g82677 (n14131, n_37855, n_37856, n7602, n7570);
  not g82678 (n_37855, n14127);
  not g82679 (n_37856, n14128);
  and g82680 (n14274, n_37857, n14271, pi0122, n14170);
  not g82681 (n_37857, n14252);
  and g82682 (n14268, n_37858, n10416, n_134, pi0950);
  not g82683 (n_37858, n14265);
  and g82684 (n14741, n_37859, n_37860, n_9722, n_9945);
  not g82685 (n_37859, n14733);
  not g82686 (n_37860, n14466);
  and g82687 (n14843, n_37861, n_37862, n14437, n_9945);
  not g82688 (n_37861, n14840);
  not g82689 (n_37862, n14742);
  and g82690 (n14784, n_37863, n_37864, n_37865, n10478);
  not g82691 (n_37863, n14773);
  not g82692 (n_37864, n14781);
  not g82693 (n_37865, n14760);
  and g82694 (n14723, n_37866, n_37867, n_37868, pi0232);
  not g82695 (n_37866, n14720);
  not g82696 (n_37867, n14698);
  not g82697 (n_37868, n14710);
  and g82698 (n14490, n14487, n9253, n_42, n14476);
  and g82699 (n14483, n14480, n2495, n_51, pi0077);
  and g82700 (n14857, n_37869, po1057, pi0110, n10075);
  not g82701 (n_37869, n10976);
  and g82702 (n15134, n_37870, n_37871, n14912, n_10233);
  not g82703 (n_37870, n15131);
  not g82704 (n_37871, n14931);
  and g82705 (n15311, n_37872, n_37873, n_10071, n_10233);
  not g82706 (n_37872, n15308);
  not g82707 (n_37873, n15135);
  and g82708 (n15207, n_37874, n_37875, pi0299, n9766);
  not g82709 (n_37874, n15204);
  not g82710 (n_37875, n15194);
  and g82711 (n15229, n_37876, n_37877, pi0299, n9760);
  not g82712 (n_37876, n15226);
  not g82713 (n_37877, n15214);
  and g82714 (n15194, n_37878, n_37879, n_37880, pi0197);
  not g82715 (n_37878, n15191);
  not g82716 (n_37879, n15190);
  not g82717 (n_37880, n15185);
  and g82718 (n15046, n_37881, n_37882, pi0152, pi0197);
  not g82719 (n_37881, n15040);
  not g82720 (n_37882, n15043);
  and g82721 (n15596, n_37883, n_37884, n_37885, n2535);
  not g82722 (n_37883, n15593);
  not g82723 (n_37884, n15328);
  not g82724 (n_37885, n15334);
  nor g82725 (n15587, n15584, n15526, n15543, n15567);
  nor g82726 (n15460, n15457, n15399, n15418, n15437);
  and g82727 (n15445, n_37886, n_37887, n_37888, pi0157);
  not g82728 (n_37886, n15441);
  not g82729 (n_37887, n15438);
  not g82730 (n_37888, n15442);
  and g82731 (n15408, n_37889, n_37890, n_9765, pi0181);
  not g82732 (n_37889, n15403);
  not g82733 (n_37890, n15405);
  and g82734 (n15435, n_37891, n_37892, n_37893, n_5686);
  not g82735 (n_37891, n15428);
  not g82736 (n_37892, n15432);
  not g82737 (n_37893, n15427);
  and g82738 (n15524, n_37894, n_37895, n_266, n_10372);
  not g82739 (n_37894, n15521);
  not g82740 (n_37895, n15520);
  and g82741 (n15541, n_37896, n_37897, n_5686, n_10372);
  not g82742 (n_37896, n15538);
  not g82743 (n_37897, n15537);
  and g82744 (n15687, n_37898, n_345, n_162, pi0129);
  not g82745 (n_37898, n15684);
  and g82746 (n15718, n_37899, n_37900, n2521, n8967);
  not g82747 (n_37899, n15715);
  not g82748 (n_37900, n15714);
  and g82749 (n15870, n_37901, n_37902, n_37903, po1038);
  not g82750 (n_37901, n15867);
  not g82751 (n_37902, n15864);
  not g82752 (n_37903, n15861);
  and g82753 (n15781, n_37904, n_37905, n_37906, pi0299);
  not g82754 (n_37904, n15773);
  not g82755 (n_37905, n15778);
  not g82756 (n_37906, n15766);
  and g82757 (n15778, n_37907, n_37908, n_6224, n9036);
  not g82758 (n_37907, n15774);
  not g82759 (n_37908, n15775);
  and g82760 (n15802, n_37909, n_37910, pi0162, pi0216);
  not g82761 (n_37909, n15799);
  not g82762 (n_37910, n15797);
  and g82763 (n16011, n_37911, n_37912, n15888, n_10905);
  not g82764 (n_37911, n16008);
  not g82765 (n_37912, n15901);
  and g82766 (n16092, n_37913, n_37914, n_10817, n_10905);
  not g82767 (n_37913, n16089);
  not g82768 (n_37914, n16012);
  and g82769 (n16089, n_37915, n_10903, n2535, n_10963);
  not g82770 (n_37915, n16086);
  and g82771 (n16082, n_37916, n_37917, n_37918, pi0232);
  not g82772 (n_37916, n16079);
  not g82773 (n_37917, n16060);
  not g82774 (n_37918, n16056);
  and g82775 (n15953, n_37919, n_37920, n_37921, pi0232);
  not g82776 (n_37919, n15950);
  not g82777 (n_37920, n15929);
  not g82778 (n_37921, n15937);
  and g82779 (n16146, n_37922, n_37923, n_37924, n11374);
  not g82780 (n_37922, n16143);
  not g82781 (n_37923, n16126);
  not g82782 (n_37924, n16136);
  and g82783 (n16143, n_37925, n_37926, n_162, n_5742);
  not g82784 (n_37925, n16140);
  not g82785 (n_37926, n16139);
  and g82786 (n16126, n_37927, n_37928, n_162, pi0176);
  not g82787 (n_37927, n16123);
  not g82788 (n_37928, n16120);
  and g82789 (n16261, n_37929, n_37930, pi0164, n_11086);
  not g82790 (n_37929, n16258);
  not g82791 (n_37930, n16254);
  and g82792 (n16245, n_37931, n_37932, n_5727, n_11086);
  not g82793 (n_37931, n16242);
  not g82794 (n_37932, n16232);
  and g82795 (n16188, n_37933, n_37934, pi0164, pi0216);
  not g82796 (n_37933, n16185);
  not g82797 (n_37934, n16184);
  and g82798 (n16549, n_37935, n_37936, n_37937, pi0232);
  not g82799 (n_37935, n16545);
  not g82800 (n_37936, n16540);
  not g82801 (n_37937, n16546);
  and g82802 (n16581, n_37938, n_37939, n_37940, n_7429);
  not g82803 (n_37938, n16577);
  not g82804 (n_37939, n16576);
  not g82805 (n_37940, n16578);
  and g82806 (n16607, n_37941, n_37942, n_37943, pi0232);
  not g82807 (n_37941, n16603);
  not g82808 (n_37942, n16599);
  not g82809 (n_37943, n16604);
  and g82810 (n17036, n_37944, n_11726, n_11725, n_36);
  not g82811 (n_37944, n17026);
  and g82812 (n17343, n17328, n_11925, n_3087, n_11552);
  and g82813 (n19481, n_37945, n_37946, pi0774, n_13711);
  not g82814 (n_37945, n19478);
  not g82815 (n_37946, n19469);
  and g82816 (n20033, n_37947, n_14098, pi0736, n_13711);
  not g82817 (n_37947, n20030);
  and g82818 (n21233, n_37948, n_37949, pi0755, n_14960);
  not g82819 (n_37948, n21229);
  not g82820 (n_37949, n21230);
  and g82821 (n21902, n_37950, n_37951, pi0756, n_14960);
  not g82822 (n_37950, n21899);
  not g82823 (n_37951, n21898);
  and g82824 (n22110, n_37952, n_37953, pi0777, n_14960);
  not g82825 (n_37952, n22106);
  not g82826 (n_37953, n22107);
  and g82827 (n22162, n_37954, n_37955, n_37956, n_15798);
  not g82828 (n_37954, n22159);
  not g82829 (n_37955, n22156);
  not g82830 (n_37956, n22154);
  and g82831 (n22202, n_37957, n_37958, n_37959, n_13620);
  not g82832 (n_37957, n22199);
  not g82833 (n_37958, n22196);
  not g82834 (n_37959, n22194);
  and g82835 (n23365, n_37960, n_16686, pi0696, n_13711);
  not g82836 (n_37960, n23362);
  and g82837 (n23975, n_37961, n_37962, n_37963, n_15272);
  not g82838 (n_37961, n23968);
  not g82839 (n_37962, n23972);
  not g82840 (n_37963, n23970);
  and g82841 (n25662, n19439, n_13679, n_7636, n_15412);
  nor g82842 (n26341, n26333, n26338, n26329, n26336);
  nor g82843 (n26818, n26810, n26815, n26806, n26813);
  nor g82844 (n28708, n28700, n28705, n28696, n28703);
  and g82845 (n29016, n_37964, n_37965, pi0752, n_13711);
  not g82846 (n_37964, n29013);
  not g82847 (n_37965, n29012);
  and g82848 (n29491, n_37966, n_37967, pi0770, n_13711);
  not g82849 (n_37966, n29488);
  not g82850 (n_37967, n29487);
  and g82851 (n29966, n_37968, n_37969, pi0768, n_13711);
  not g82852 (n_37968, n29963);
  not g82853 (n_37969, n29962);
  and g82854 (n30483, n_37970, n_22302, pi0727, n_13711);
  not g82855 (n_37970, n30480);
  and g82856 (n31088, n_37971, n_37972, n_37973, n_15952);
  not g82857 (n_37971, n31081);
  not g82858 (n_37972, n31085);
  not g82859 (n_37973, n31083);
  and g82860 (n31565, n_37974, n_37975, n_37976, n_16012);
  not g82861 (n_37974, n31558);
  not g82862 (n_37975, n31562);
  not g82863 (n_37976, n31560);
  and g82864 (n32042, n_37977, n_37978, n_37979, n_16133);
  not g82865 (n_37977, n32035);
  not g82866 (n_37978, n32039);
  not g82867 (n_37979, n32037);
  and g82868 (n33211, n_37980, n_37981, n_37982, n10200);
  not g82869 (n_37980, n33206);
  not g82870 (n_37981, n33208);
  not g82871 (n_37982, n33197);
  and g82872 (n33203, n_37983, n_37984, n_37985, n_7429);
  not g82873 (n_37983, n33199);
  not g82874 (n_37984, n33198);
  not g82875 (n_37985, n33200);
  and g82876 (n33231, n_37986, n_37987, n_37988, pi0232);
  not g82877 (n_37986, n33227);
  not g82878 (n_37987, n33223);
  not g82879 (n_37988, n33228);
  and g82880 (n33416, n_37989, n_37990, n2571, n10982);
  not g82881 (n_37989, n33413);
  not g82882 (n_37990, n33401);
  and g82883 (n33787, n_37991, n_37992, n_24770, pi0603);
  not g82884 (n_37991, n33784);
  not g82885 (n_37992, n33779);
  and g82886 (n33767, n_37993, n33580, n_24724, pi0633);
  not g82887 (n_37993, n33764);
  and g82888 (n33862, n_37994, n_37995, n_37996, n_24970);
  not g82889 (n_37994, n33858);
  not g82890 (n_37995, n33857);
  not g82891 (n_37996, n33859);
  and g82892 (n34084, n_37997, n_37998, n_25117, n_13709);
  not g82893 (n_37997, n34079);
  not g82894 (n_37998, n34081);
  nor g82895 (n_38000, n34456, n34450);
  and g82896 (n34460, n_37999, pi0606, n2571, n_38000);
  not g82897 (n_37999, n34452);
  and g82898 (n34692, n_38001, n_38002, n_234, n_3446);
  not g82899 (n_38001, n34689);
  not g82900 (n_38002, n34687);
  and g82901 (n35227, n_38003, n_38004, pi0619, n_11403);
  not g82902 (n_38003, n35224);
  not g82903 (n_38004, n35223);
  and g82904 (n35222, n_38005, n_38006, n_11821, pi0648);
  not g82905 (n_38005, n35219);
  not g82906 (n_38006, n35218);
  and g82907 (n35643, n_38007, n_38008, n_38009, pi0209);
  not g82908 (n_38007, n35640);
  not g82909 (n_38008, n35601);
  not g82910 (n_38009, n35580);
  and g82911 (n35909, n_38010, n_38011, n_26602, n_223);
  not g82912 (n_38010, n35906);
  not g82913 (n_38011, n35889);
  and g82914 (n36075, n_38012, n_26587, pi0216, n_26654);
  not g82915 (n_38012, n36072);
  and g82916 (n36052, n_38013, n_38014, n_26602, n_223);
  not g82917 (n_38013, n36049);
  not g82918 (n_38014, n36003);
  and g82919 (n36042, n_26695, n_26694, n_3119, n_26654);
  and g82920 (n36236, n_26587, n_26833, pi0221, n_26781);
  and g82921 (n36219, n_38015, n_38016, pi0223, n_26781);
  not g82922 (n_38015, n36216);
  not g82923 (n_38016, n36208);
  and g82924 (n36409, n_38017, n_38018, n_38019, n_162);
  not g82925 (n_38017, n36406);
  not g82926 (n_38018, n36405);
  not g82927 (n_38019, n36404);
  and g82928 (n36278, n_38020, n_38021, n_38022, pi0299);
  not g82929 (n_38020, n36275);
  not g82930 (n_38021, n36274);
  not g82931 (n_38022, n36273);
  and g82932 (n36272, n_38023, n_38024, n_38025, n_234);
  not g82933 (n_38023, n36268);
  not g82934 (n_38024, n36267);
  not g82935 (n_38025, n36269);
  and g82936 (n36642, n_38026, n_38027, n_27156, pi0680);
  not g82937 (n_38026, n36637);
  not g82938 (n_38027, n36639);
  and g82939 (n37239, n_38028, n_27227, pi0223, n_27434);
  not g82940 (n_38028, n37236);
  and g82941 (n36899, n_38029, n_38030, n_38031, pi0299);
  not g82942 (n_38029, n36896);
  not g82943 (n_38030, n36895);
  not g82944 (n_38031, n36894);
  and g82945 (n36893, n_38032, n_38033, n_38034, n_234);
  not g82946 (n_38032, n36889);
  not g82947 (n_38033, n36888);
  not g82948 (n_38034, n36890);
  and g82949 (n37287, n_38035, n_38036, n_38037, pi0680);
  not g82950 (n_38035, n37283);
  not g82951 (n_38036, n37284);
  not g82952 (n_38037, n37281);
  and g82953 (n37261, n_38038, n_38039, pi0680, n_12002);
  not g82954 (n_38038, n37258);
  not g82955 (n_38039, n37257);
  and g82956 (n37307, n_38040, n_38041, n_38042, pi0680);
  not g82957 (n_38040, n37304);
  not g82958 (n_38041, n37303);
  not g82959 (n_38042, n37302);
  and g82960 (n37324, n_38043, n_38044, n_12083, pi0680);
  not g82961 (n_38043, n37321);
  not g82962 (n_38044, n37320);
  and g82963 (n37478, n_38045, n_38046, n_38047, pi0299);
  not g82964 (n_38045, n37475);
  not g82965 (n_38046, n37474);
  not g82966 (n_38047, n37473);
  and g82967 (n37472, n_38048, n_38049, n_38050, n_234);
  not g82968 (n_38048, n37468);
  not g82969 (n_38049, n37467);
  not g82970 (n_38050, n37469);
  and g82971 (n37841, n_38051, n_38052, n_38053, n_223);
  not g82972 (n_38051, n37838);
  not g82973 (n_38052, n37809);
  not g82974 (n_38053, n37787);
  and g82975 (n37499, n_38054, n_38055, n_38056, n_223);
  not g82976 (n_38054, n37490);
  not g82977 (n_38055, n37496);
  not g82978 (n_38056, n37481);
  and g82979 (n37701, n_38057, n_38058, n_38059, n_223);
  not g82980 (n_38057, n37698);
  not g82981 (n_38058, n37694);
  not g82982 (n_38059, n37690);
  and g82983 (n37878, n_38060, n_38061, n_12108, pi0680);
  not g82984 (n_38060, n37875);
  not g82985 (n_38061, n37874);
  and g82986 (n_38063, n_38062, n_7437);
  not g82987 (n_38062, n38261);
  and g82988 (n38265, n2967, n_142, n10235, n_38063);
  and g82989 (n38715, n_38064, n_38065, n_38066, n_4226);
  not g82990 (n_38064, n38640);
  not g82991 (n_38065, n38667);
  not g82992 (n_38066, n38712);
  and g82993 (n38712, n_38067, n_38068, n_6933, n_28735);
  not g82994 (n_38067, n38709);
  not g82995 (n_38068, n38679);
  and g82996 (n39153, n_38069, n38416, pi0213, n_29079);
  not g82997 (n_38069, n39150);
  and g82998 (n39136, n_38070, n_38071, n_38072, n_6791);
  not g82999 (n_38070, n39120);
  not g83000 (n_38071, n39133);
  not g83001 (n_38072, n39109);
  and g83002 (n39168, n_38073, po1038, n_29089, n_29090);
  not g83003 (n_38073, n39165);
  and g83004 (n39820, n_38074, n_38075, n_4226, n_29607);
  not g83005 (n_38074, n39817);
  not g83006 (n_38075, n39791);
  and g83007 (n39902, n_38076, n_38077, n_38078, n_6791);
  not g83008 (n_38076, n39897);
  not g83009 (n_38077, n39898);
  not g83010 (n_38078, n39899);
  and g83011 (n39767, n_38079, n_38080, n_38081, n_6791);
  not g83012 (n_38079, n39761);
  not g83013 (n_38080, n39764);
  not g83014 (n_38081, n39751);
  and g83015 (n39815, n_38082, n_38083, n_38084, pi0212);
  not g83016 (n_38082, n39812);
  not g83017 (n_38083, n39811);
  not g83018 (n_38084, n39810);
  and g83019 (n39839, n_38085, n_38086, n39834, n_29471);
  not g83020 (n_38085, n39835);
  not g83021 (n_38086, n39836);
  and g83022 (n39691, n_38087, n_38088, n_38089, pi0212);
  not g83023 (n_38087, n39681);
  not g83024 (n_38088, n39688);
  not g83025 (n_38089, n39680);
  and g83026 (n40027, n_38090, n_38091, n_38092, pi0213);
  not g83027 (n_38090, n39997);
  not g83028 (n_38091, n40024);
  not g83029 (n_38092, n39999);
  and g83030 (n39997, n_38093, n_38094, n_26372, n39971);
  not g83031 (n_38093, n39988);
  not g83032 (n_38094, n39994);
  and g83033 (n40024, n_38095, n_38096, pi0209, n40015);
  not g83034 (n_38095, n40013);
  not g83035 (n_38096, n40021);
  and g83036 (n40645, n_30245, n_29518, n_6791, n_29977);
  and g83037 (n41166, n_38097, n_38098, n16479, n_28836);
  not g83038 (n_38097, n41163);
  not g83039 (n_38098, n40946);
  and g83040 (n40976, n_38099, n_38100, n_38101, pi0219);
  not g83041 (n_38099, n40964);
  not g83042 (n_38100, n40967);
  not g83043 (n_38101, n40973);
  and g83044 (n40896, n_38102, n_38103, n_38104, n_6791);
  not g83045 (n_38102, n40892);
  not g83046 (n_38103, n40893);
  not g83047 (n_38104, n40883);
  and g83048 (n41067, n_38105, n_38106, n_38107, n_11794);
  not g83049 (n_38105, n41061);
  not g83050 (n_38106, n41056);
  not g83051 (n_38107, n41064);
  and g83052 (n41201, n_38108, n_38109, n_26557, n_29304);
  not g83053 (n_38108, n41189);
  not g83054 (n_38109, n41198);
  and g83055 (n41198, n_38110, n_38111, n40410, pi1147);
  not g83056 (n_38110, n41195);
  not g83057 (n_38111, n41190);
  and g83058 (n41212, n_38112, n_38113, n_38114, n38665);
  not g83059 (n_38112, n41209);
  not g83060 (n_38113, n41208);
  not g83061 (n_38114, n41207);
  and g83062 (n41461, n_38115, n_38116, n_29904, n_30383);
  not g83063 (n_38115, n41458);
  not g83064 (n_38116, n41444);
  and g83065 (n41432, n_38117, n_38118, pi1148, n_30383);
  not g83066 (n_38117, n41429);
  not g83067 (n_38118, n41417);
  and g83068 (n41700, n_38119, n_38120, pi1150, n_29872);
  not g83069 (n_38119, n41691);
  not g83070 (n_38120, n41697);
  and g83071 (n41686, n_38121, n_38122, n_30133, n_29646);
  not g83072 (n_38121, n41683);
  not g83073 (n_38122, n41679);
  and g83074 (n41731, n_38123, n_38124, n_30133, n_29848);
  not g83075 (n_38123, n41726);
  not g83076 (n_38124, n41728);
  nor g83077 (n_38125, n41525, n41526);
  and g83078 (n41530, n_30734, n_30826, n_6791, n_38125);
  and g83079 (n41635, n_38126, n_38127, n_30133, n_29842);
  not g83080 (n_38126, n41632);
  not g83081 (n_38127, n41620);
  and g83082 (n41710, n_38128, n_31076, n_796, pi1147);
  not g83083 (n_38128, n41707);
  nor g83084 (n_38129, n41712, n41713);
  and g83085 (n41717, n_31076, n_796, n_29810, n_38129);
  and g83086 (n41571, n_38130, n41567, n_29796, n_29958);
  not g83087 (n_38130, n41568);
  and g83088 (n42212, n_38131, n_38132, n38922, n_31422);
  not g83089 (n_38131, n42205);
  not g83090 (n_38132, n42206);
  and g83091 (n42171, n_38133, n_31385, n_796, n_29468);
  not g83092 (n_38133, n42168);
  and g83093 (n42155, n_38134, n_31385, n_796, pi1151);
  not g83094 (n_38134, n42152);
  and g83095 (n42203, n_38135, n_38136, n_31409, n_6791);
  not g83096 (n_38135, n42200);
  not g83097 (n_38136, n42197);
  and g83098 (po0407, n_38137, n8881, n_172, n_3208);
  not g83099 (n_38137, n42329);
  and g83100 (n_38138, n6380, n_28488);
  and g83101 (n_38139, n6217, n21130);
  and g83102 (n42378, n10982, n42347, n_38138, n_38139);
  and g83103 (n42492, n_38140, n_38141, n_38142, pi1152);
  not g83104 (n_38140, n42482);
  not g83105 (n_38141, n42489);
  not g83106 (n_38142, n42457);
  and g83107 (n42407, n_38143, n_28715, n_29468, n_7410);
  not g83108 (n_38143, n42404);
  and g83109 (n42452, n_38144, n_38145, n_29468, n_31607);
  not g83110 (n_38144, n42447);
  not g83111 (n_38145, n42449);
  and g83112 (n42742, n_38146, n_31670, n_31763, n_31825);
  not g83113 (n_38146, n42739);
  and g83114 (n42738, n_38147, n42734, n_31825, pi0254);
  not g83115 (n_38147, n42735);
  and g83116 (n42787, n_38148, n_38149, n_38150, n_31763);
  not g83117 (n_38148, n42781);
  not g83118 (n_38149, n42776);
  not g83119 (n_38150, n42784);
  and g83120 (n42821, n_38151, n_38152, n_38153, pi0219);
  not g83121 (n_38151, n42818);
  not g83122 (n_38152, n42779);
  not g83123 (n_38153, n42775);
  and g83124 (n42833, n_38154, n_38155, n_38156, n_6791);
  not g83125 (n_38154, n42830);
  not g83126 (n_38155, n42827);
  not g83127 (n_38156, n42824);
  and g83128 (n42703, n_38157, n_38158, pi0219, n_31791);
  not g83129 (n_38157, n42697);
  not g83130 (n_38158, n42700);
  and g83131 (n42667, n_29000, n_28945, pi1091, n38488);
  and g83132 (n42984, n_38159, n_38160, pi0263, pi1091);
  not g83133 (n_38159, n42981);
  not g83134 (n_38160, n42968);
  and g83135 (n43083, n_38161, n_38162, n_38163, pi0219);
  not g83136 (n_38161, n43080);
  not g83137 (n_38162, n43078);
  not g83138 (n_38163, n43075);
  and g83139 (n43065, n_38164, n_38165, n_38166, pi0219);
  not g83140 (n_38164, n43058);
  not g83141 (n_38165, n43056);
  not g83142 (n_38166, n43062);
  and g83143 (n42942, n_38167, n_38168, n_38169, pi0219);
  not g83144 (n_38167, n42933);
  not g83145 (n_38168, n42939);
  not g83146 (n_38169, n42927);
  and g83147 (n42939, n_38170, n_38171, pi1091, n38483);
  not g83148 (n_38170, n42934);
  not g83149 (n_38171, n42936);
  and g83150 (n43395, n_38172, n_38173, n_38174, n_32322);
  not g83151 (n_38172, n43385);
  not g83152 (n_38173, n43389);
  not g83153 (n_38174, n43392);
  and g83154 (n43389, n_31840, n_32345, n38487, n_32101);
  and g83155 (n43433, n_38175, n_32373, pi1154, n_32124);
  not g83156 (n_38175, n43430);
  and g83157 (n43383, n_31855, n_30538, pi1154, pi1155);
  and g83158 (n43520, n_38176, n_38177, n_38178, n_30133);
  not g83159 (n_38176, n43517);
  not g83160 (n_38177, n43512);
  not g83161 (n_38178, n43507);
  nor g83162 (po0459, n44572, n44569, n44566, n44578);
  and g83163 (n44622, n_38179, n_38180, pi1147, n_33350);
  not g83164 (n_38179, n44619);
  not g83165 (n_38180, n44618);
  and g83166 (n45175, n_38181, n_38182, n_38183, po1038);
  not g83167 (n_38181, n45170);
  not g83168 (n_38182, n45171);
  not g83169 (n_38183, n45172);
  nor g83170 (po0623, n45184, n45191, n45181, n45188);
  and g83171 (n_38185, n_38184, n16845);
  not g83172 (n_38184, n45199);
  and g83173 (n45203, n16847, n8897, n10162, n_38185);
  and g83174 (n45228, n8962, n10197, pi0038, n_162);
  and g83175 (n45249, n_38186, n_38187, n_38188, po1038);
  not g83176 (n_38186, n45246);
  not g83177 (n_38187, n45244);
  not g83178 (n_38188, n45245);
  and g83179 (n45269, n_38189, n_38190, n_38191, po1038);
  not g83180 (n_38189, n45266);
  not g83181 (n_38190, n45264);
  not g83182 (n_38191, n45265);
  and g83183 (n45289, n_38192, n_38193, n_38194, po1038);
  not g83184 (n_38192, n45286);
  not g83185 (n_38193, n45284);
  not g83186 (n_38194, n45285);
  and g83187 (n45309, n_38195, n_38196, n_38197, po1038);
  not g83188 (n_38195, n45306);
  not g83189 (n_38196, n45304);
  not g83190 (n_38197, n45305);
  nor g83191 (po0630, n45315, n45318, n45312, n45316);
  nor g83192 (po0631, n45326, n45329, n45323, n45327);
  nor g83193 (po0632, n45337, n45340, n45334, n45338);
  and g83194 (n45352, n_38198, n13050, n2572, n10162);
  not g83195 (n_38198, n45349);
  and g83196 (n_38199, pi0603, n_11960);
  and g83197 (n45638, n_14295, n17182, n_14288, n_38199);
  and g83198 (n_38200, n30797, n20237);
  and g83199 (n_38201, n_26377, n_14288);
  and g83200 (n45805, pi0230, n17168, n_38200, n_38201);
  and g83201 (n46605, n_38202, n46596, n_34545, n46599);
  not g83202 (n_38202, n46602);
  and g83203 (n46609, n46596, n46599, pi0560, n_34545);
  nor g83204 (n_38205, n46591, n46584);
  nor g83205 (n_38206, n46590, n46587);
  and g83206 (n46596, n_38203, n_38204, n_38205, n_38206);
  not g83207 (n_38203, n46585);
  not g83208 (n_38204, n46586);
  nor g83209 (n_38207, n45856, n45846, n45849);
  nor g83210 (n_38208, n45850, n45851);
  nor g83211 (n_38209, n45852, n45855);
  nor g83212 (n_38210, n45847, n45848);
  and g83213 (n45864, n_38207, n_38208, n_38209, n_38210);
  nor g83214 (n_38214, n46370, n46360);
  and g83215 (n46374, n_38211, n_38212, n_38213, n_38214);
  not g83216 (n_38211, n46369);
  not g83217 (n_38212, n46363);
  not g83218 (n_38213, n46366);
  nor g83219 (n_38217, n45905, n45904);
  nor g83220 (n_38218, n45910, n45902);
  and g83221 (n45915, n_38215, n_38216, n_38217, n_38218);
  not g83222 (n_38215, n45906);
  not g83223 (n_38216, n45907);
  nor g83224 (n_38219, n46539, n46527, n46535);
  nor g83225 (n_38220, n46536, n46537, n46538);
  nor g83226 (n_38221, n46530, n46531, n46532);
  nor g83227 (n_38222, n46533, n46534);
  and g83228 (n46549, n_38219, n_38220, n_38221, n_38222);
  nor g83229 (n_38226, n46323, n46322);
  and g83230 (n46327, n_38223, n_38224, n_38225, n_38226);
  not g83231 (n_38223, n46321);
  not g83232 (n_38224, n46315);
  not g83233 (n_38225, n46318);
  nor g83234 (n_38227, n17856, n46768);
  and g83235 (n_38228, n19151, pi0230);
  and g83236 (n_38229, n16644, n_13449);
  and g83237 (n46774, n_13598, n_38227, n_38228, n_38229);
  nor g83238 (n_38230, pi0973, pi1054);
  and g83239 (n46888, pi0832, pi1088, pi1066, n_38230);
  and g83240 (n47095, n_38231, n_38232, n_38233, n47092);
  not g83241 (n_38231, n47087);
  not g83242 (n_38232, n47088);
  not g83243 (n_38233, n47089);
  and g83244 (n47160, n_38234, n_38235, n_38236, n47092);
  not g83245 (n_38234, n47155);
  not g83246 (n_38235, n47156);
  not g83247 (n_38236, n47157);
  and g83248 (n47233, n_38237, n_38238, n_38239, n47092);
  not g83249 (n_38237, n47228);
  not g83250 (n_38238, n47229);
  not g83251 (n_38239, n47230);
  and g83252 (n47281, n_38240, n_38241, n_38242, n47092);
  not g83253 (n_38240, n47278);
  not g83254 (n_38241, n47276);
  not g83255 (n_38242, n47277);
  and g83256 (n47287, n_38243, n_38244, n47283, n_2921);
  not g83257 (n_38243, n47284);
  not g83258 (n_38244, n47282);
  and g83259 (n47314, n_38245, n_38246, n_38247, n47092);
  not g83260 (n_38245, n47311);
  not g83261 (n_38246, n47309);
  not g83262 (n_38247, n47310);
  and g83263 (n47319, n_38248, n_38249, n47283, n_2921);
  not g83264 (n_38248, n47316);
  not g83265 (n_38249, n47315);
  and g83266 (n47338, n_38250, n_38251, n_38252, n47092);
  not g83267 (n_38250, n47333);
  not g83268 (n_38251, n47334);
  not g83269 (n_38252, n47335);
  and g83270 (n47374, n_38253, n_38254, n_38255, n47092);
  not g83271 (n_38253, n47369);
  not g83272 (n_38254, n47370);
  not g83273 (n_38255, n47371);
  and g83274 (n47484, n_38256, n_38257, n_38258, n47092);
  not g83275 (n_38256, n47479);
  not g83276 (n_38257, n47480);
  not g83277 (n_38258, n47481);
  and g83278 (n47528, n_38259, n_38260, n_38261, n47092);
  not g83279 (n_38259, n47525);
  not g83280 (n_38260, n47523);
  not g83281 (n_38261, n47524);
  and g83282 (n47533, n_38262, n_38263, n47283, n_2921);
  not g83283 (n_38262, n47530);
  not g83284 (n_38263, n47529);
  and g83285 (n47560, n_38264, n_38265, n_38266, n47092);
  not g83286 (n_38264, n47557);
  not g83287 (n_38265, n47555);
  not g83288 (n_38266, n47556);
  and g83289 (n47565, n_38267, n_38268, n47283, n_2921);
  not g83290 (n_38267, n47562);
  not g83291 (n_38268, n47561);
  and g83292 (n47602, n_38269, n_38270, n_38271, n47092);
  not g83293 (n_38269, n47597);
  not g83294 (n_38270, n47598);
  not g83295 (n_38271, n47599);
  and g83296 (n47637, n_38272, n_38273, n_38274, n47092);
  not g83297 (n_38272, n47634);
  not g83298 (n_38273, n47632);
  not g83299 (n_38274, n47633);
  and g83300 (n47642, n_38275, n_38276, n47283, n_2921);
  not g83301 (n_38275, n47639);
  not g83302 (n_38276, n47638);
  and g83303 (n47733, n_38277, n_38278, n_38279, n47092);
  not g83304 (n_38277, n47728);
  not g83305 (n_38278, n47729);
  not g83306 (n_38279, n47730);
  and g83307 (n47862, n_38280, n_38281, n47283, n_2921);
  not g83308 (n_38280, n47859);
  not g83309 (n_38281, n47858);
  and g83310 (n47868, n_38282, n_38283, n_38284, n47092);
  not g83311 (n_38282, n47865);
  not g83312 (n_38283, n47863);
  not g83313 (n_38284, n47864);
  and g83314 (n47895, n_38285, n_38286, n_38287, n7643);
  not g83315 (n_38285, n47885);
  not g83316 (n_38286, n47892);
  not g83317 (n_38287, n47874);
  nor g83318 (n_38289, n47904, n47903);
  and g83319 (n47908, n_38288, n47901, pi1134, n_38289);
  not g83320 (n_38288, n47902);
  and g83321 (n47900, n_38290, n_38291, n47283, n_2921);
  not g83322 (n_38290, n47897);
  not g83323 (n_38291, n47896);
  and g83324 (n47944, n_38292, n_38293, n47283, n_2921);
  not g83325 (n_38292, n47941);
  not g83326 (n_38293, n47940);
  and g83327 (n47950, n_38294, n_38295, n_38296, n47092);
  not g83328 (n_38294, n47947);
  not g83329 (n_38295, n47945);
  not g83330 (n_38296, n47946);
  and g83331 (n47973, n_38297, n_38298, n_38299, n_34961);
  not g83332 (n_38297, n47970);
  not g83333 (n_38298, n47969);
  not g83334 (n_38299, n47968);
  nor g83335 (n_38301, n47956, n47955);
  and g83336 (n47960, n_38300, n47901, pi1134, n_38301);
  not g83337 (n_38300, n47954);
  and g83338 (n47965, n_38302, n_38303, n47283, n_2921);
  not g83339 (n_38302, n47962);
  not g83340 (n_38303, n47961);
  and g83341 (n48013, n_38304, n_38305, n47283, n_2921);
  not g83342 (n_38304, n48010);
  not g83343 (n_38305, n48009);
  and g83344 (n48019, n_38306, n_38307, n_38308, n47092);
  not g83345 (n_38306, n48016);
  not g83346 (n_38307, n48014);
  not g83347 (n_38308, n48015);
  and g83348 (n48082, n_38309, n_38310, n_38311, n7643);
  not g83349 (n_38309, n48072);
  not g83350 (n_38310, n48079);
  not g83351 (n_38311, n48063);
  nor g83352 (n_38313, n48090, n48089);
  and g83353 (n48094, n_38312, n47901, pi1134, n_38313);
  not g83354 (n_38312, n48088);
  and g83355 (n48087, n_38314, n_38315, n47283, n_2921);
  not g83356 (n_38314, n48084);
  not g83357 (n_38315, n48083);
  nor g83358 (n_38317, n48116, n48117);
  and g83359 (n48121, n_38316, n47901, pi1134, n_38317);
  not g83360 (n_38316, n48115);
  and g83361 (n48152, n_38318, n_38319, n_38320, n7643);
  not g83362 (n_38318, n48142);
  not g83363 (n_38319, n48149);
  not g83364 (n_38320, n48133);
  nor g83365 (n_38322, n48160, n48159);
  and g83366 (n48164, n_38321, n47901, pi1134, n_38322);
  not g83367 (n_38321, n48158);
  and g83368 (n48157, n_38323, n_38324, n47283, n_2921);
  not g83369 (n_38323, n48154);
  not g83370 (n_38324, n48153);
  nor g83371 (n_38326, n48186, n48187);
  and g83372 (n48191, n_38325, n47901, pi1134, n_38326);
  not g83373 (n_38325, n48185);
  and g83374 (n48275, n48271, n48272, pi0794, pi0801);
  and g83375 (n48324, n_38327, n_38328, pi1135, pi1136);
  not g83376 (n_38327, n48321);
  not g83377 (n_38328, n48320);
  and g83378 (n_38329, n48271, n48367);
  and g83379 (n48371, n_35892, n_35921, pi0801, n_38329);
  and g83380 (n48401, n_38330, n_38331, n_38332, n7643);
  not g83381 (n_38330, n48391);
  not g83382 (n_38331, n48398);
  not g83383 (n_38332, n48382);
  nor g83384 (n_38334, n48409, n48408);
  and g83385 (n48413, n_38333, n47901, pi1134, n_38334);
  not g83386 (n_38333, n48407);
  and g83387 (n48406, n_38335, n_38336, n47283, n_2921);
  not g83388 (n_38335, n48403);
  not g83389 (n_38336, n48402);
  and g83390 (n48478, n_38337, n48471, n_35894, n_35892);
  not g83391 (n_38337, n48475);
  and g83392 (n48555, n_35890, n_35880, n_35882, n_35875);
  and g83393 (n_38338, n_35893, n48367);
  and g83394 (n48588, n_35894, pi0794, n_35895, n_38338);
  and g83395 (n_38339, n48256, n_35977);
  and g83396 (n_38340, pi0795, pi0800);
  and g83397 (n48640, pi0801, n_35896, n_38339, n_38340);
  nor g83398 (n_38341, pi1046, pi1083);
  and g83399 (n48660, pi0832, pi0956, pi1085, n_38341);
  and g83400 (n_38342, pi0266, n_34942);
  and g83401 (n48712, n_33067, pi0278, pi0279, n_38342);
  and g83402 (po0989, n8874, pi1162, n_12415, pi1091);
  and g83403 (po1080, n_33308, pi0301, pi0311, n_33305);
endmodule

